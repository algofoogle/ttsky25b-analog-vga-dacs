* NGSPICE file created from csdac255_parax.ext - technology: sky130A

.subckt csdac255_parax Iout VPWR VGND Vbias data[0] data[1] data[2] data[3] data[4]
+ data[5] data[6] data[7] bias[0] bias[1] bias[2]
X0 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout VGND.t1530 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1 VPWR.t1495 XThR.Tn[2].t12 XA.XIR[3].XIC[8].icell.PUM VPWR.t1494 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2 XA.XIR[12].XIC[10].icell.SM XA.XIR[12].XIC[10].icell.Ien Iout.t232 VGND.t2102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X3 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t381 VPWR.t383 VPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X4 VGND.t812 XThC.Tn[10].t12 XA.XIR[4].XIC[10].icell.PDM VGND.t811 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X5 VGND.t2390 XThR.XTBN.Y a_n997_2667# VGND.t2352 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t1578 XThR.Tn[6].t12 XA.XIR[7].XIC[8].icell.PUM VPWR.t1577 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X7 XA.XIR[14].XIC[5].icell.Ien XThR.Tn[14].t12 VPWR.t505 VPWR.t504 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X8 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12].t12 XA.XIR[12].XIC[6].icell.Ien VGND.t2681 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X9 XThC.Tn[6].t3 XThC.XTBN.Y.t4 VGND.t1140 VGND.t1139 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1926 VGND.t1506 VGND.t1505 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X11 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[9].t12 VGND.t435 VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X12 VGND.t36 XThC.XTBN.Y.t5 XThC.Tn[5].t3 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 XA.XIR[15].XIC[9].icell.PUM XThC.Tn[9].t12 XA.XIR[15].XIC[9].icell.Ien VPWR.t465 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X14 XA.XIR[9].XIC[0].icell.SM XA.XIR[9].XIC[0].icell.Ien Iout.t150 VGND.t1134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X15 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[12].t13 VGND.t2683 VGND.t2682 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X16 VGND.t2405 XThC.Tn[11].t12 XA.XIR[12].XIC[11].icell.PDM VGND.t2404 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X17 XA.XIR[12].XIC[1].icell.SM XA.XIR[12].XIC[1].icell.Ien Iout.t215 VGND.t1836 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X18 XA.XIR[8].XIC[12].icell.SM XA.XIR[8].XIC[12].icell.Ien Iout.t19 VGND.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X19 XThC.Tn[12].t3 XThC.XTB5.Y VPWR.t503 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 XA.XIR[8].XIC_15.icell.PDM VPWR.t1927 VGND.t1508 VGND.t1507 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X21 XA.XIR[7].XIC[13].icell.SM XA.XIR[7].XIC[13].icell.Ien Iout.t13 VGND.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X22 XA.XIR[14].XIC[13].icell.PUM XThC.Tn[13].t12 XA.XIR[14].XIC[13].icell.Ien VPWR.t902 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X23 a_2979_9615# XThC.XTBN.Y.t6 XThC.Tn[0].t10 VPWR.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t379 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t380 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X25 XA.XIR[10].XIC[14].icell.SM XA.XIR[10].XIC[14].icell.Ien Iout.t93 VGND.t688 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X26 a_4861_9615# XThC.XTB4.Y.t2 VPWR.t980 VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_5949_9615# XThC.XTBN.Y.t7 XThC.Tn[5].t7 VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6].t13 XA.XIR[6].XIC[10].icell.Ien VGND.t1666 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X29 XA.XIR[0].XIC[4].icell.PDM VGND.t1077 VGND.t1079 VGND.t1078 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X30 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[3].t12 VGND.t1441 VGND.t1440 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X31 XThR.Tn[5].t11 XThR.XTBN.Y a_n1049_5611# VPWR.t1756 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 XThC.Tn[4].t3 XThC.XTB5.Y VGND.t146 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND.t38 XThC.XTBN.Y.t8 XThC.Tn[2].t9 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 XThR.XTB2.Y XThR.XTB6.A VPWR.t448 VPWR.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[6].t14 VGND.t1668 VGND.t1667 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X36 XA.XIR[6].XIC[11].icell.SM XA.XIR[6].XIC[11].icell.Ien Iout.t18 VGND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X37 VGND.t1324 XThC.Tn[2].t12 XA.XIR[12].XIC[2].icell.PDM VGND.t1323 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X38 VPWR.t378 VPWR.t376 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t377 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X39 VGND.t1510 VPWR.t1928 XA.XIR[7].XIC_dummy_left.icell.PDM VGND.t1509 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X40 VPWR.t1391 XThR.Tn[3].t13 XA.XIR[4].XIC[11].icell.PUM VPWR.t1390 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X41 VGND.t789 Vbias.t6 XA.XIR[14].XIC[11].icell.SM VGND.t788 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X42 XA.XIR[2].XIC[1].icell.PUM XThC.Tn[1].t12 XA.XIR[2].XIC[1].icell.Ien VPWR.t763 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X43 VGND.t477 XThC.Tn[3].t12 XA.XIR[15].XIC[3].icell.PDM VGND.t476 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X44 VGND.t1512 VPWR.t1929 XA.XIR[10].XIC_15.icell.PDM VGND.t1511 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X45 VPWR.t879 XThR.Tn[10].t12 XA.XIR[11].XIC[9].icell.PUM VPWR.t878 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X46 XA.XIR[0].XIC[14].icell.PUM XThC.Tn[14].t12 XA.XIR[0].XIC[14].icell.Ien VPWR.t1038 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X47 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t373 VPWR.t375 VPWR.t374 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X48 a_7651_9569# XThC.XTB1.Y.t3 XThC.Tn[8].t11 VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 VGND.t791 Vbias.t7 XA.XIR[2].XIC[5].icell.SM VGND.t790 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X50 XA.XIR[1].XIC[6].icell.Ien XThR.Tn[1].t12 VPWR.t1598 VPWR.t1597 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X51 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t11 VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 VGND.t1802 XThC.Tn[4].t12 XA.XIR[2].XIC[4].icell.PDM VGND.t1801 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X53 XThC.XTB5.Y XThC.XTB7.B VGND.t1184 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 XThC.Tn[7].t3 XThC.XTBN.Y.t9 VPWR.t423 VPWR.t422 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X55 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[9].t13 VGND.t437 VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X56 VGND.t1369 XThR.XTB7.Y XThR.Tn[6].t3 VGND.t1368 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X57 XA.XIR[4].XIC[7].icell.Ien XThR.Tn[4].t12 VPWR.t1636 VPWR.t1635 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X58 VPWR.t1820 XThR.XTBN.Y XThR.Tn[9].t11 VPWR.t1807 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 XThR.XTB7.Y XThR.XTB7.A VGND.t1591 VGND.t1590 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 XA.XIR[3].XIC[8].icell.Ien XThR.Tn[3].t14 VPWR.t1393 VPWR.t1392 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X61 VPWR.t1395 XThR.Tn[3].t15 XA.XIR[4].XIC[2].icell.PUM VPWR.t1394 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X62 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[12].t14 VGND.t2685 VGND.t2684 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X63 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[1].t13 XA.XIR[1].XIC[9].icell.Ien VGND.t1705 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X64 VPWR.t1493 XThR.Tn[2].t13 XA.XIR[3].XIC[3].icell.PUM VPWR.t1492 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X65 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout VGND.t357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X66 VPWR.t1580 XThR.Tn[6].t15 XA.XIR[7].XIC[3].icell.PUM VPWR.t1579 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X67 VPWR.t372 VPWR.t370 XA.XIR[2].XIC_15.icell.PUM VPWR.t371 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X68 a_6243_9615# XThC.XTB7.Y VPWR.t1212 VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X69 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11].t12 XA.XIR[11].XIC[14].icell.Ien VGND.t1574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X70 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11].t13 XA.XIR[11].XIC[8].icell.Ien VGND.t1575 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X71 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[3].t16 VGND.t1443 VGND.t1442 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X72 XThR.Tn[7].t3 XThR.XTBN.Y VPWR.t1819 VPWR.t1818 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[0].t12 VGND.t753 VGND.t752 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X74 a_8963_9569# XThC.XTBN.Y.t10 VGND.t40 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X75 VGND.t793 Vbias.t8 XA.XIR[12].XIC[7].icell.SM VGND.t792 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X76 VGND.t2546 XThC.Tn[6].t12 XA.XIR[12].XIC[6].icell.PDM VGND.t2545 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X77 XA.XIR[6].XIC[9].icell.SM XA.XIR[6].XIC[9].icell.Ien Iout.t111 VGND.t781 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X78 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout VGND.t639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X79 XA.XIR[3].XIC[11].icell.SM XA.XIR[3].XIC[11].icell.Ien Iout.t176 VGND.t1372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X80 VGND.t1514 VPWR.t1930 XA.XIR[4].XIC_dummy_left.icell.PDM VGND.t1513 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X81 VGND.t2389 XThR.XTBN.Y XThR.Tn[5].t7 VGND.t2372 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 VGND.t795 Vbias.t9 XA.XIR[15].XIC[8].icell.SM VGND.t794 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X83 VGND.t797 Vbias.t10 XA.XIR[14].XIC[9].icell.SM VGND.t796 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X84 VGND.t775 XThC.Tn[7].t8 XA.XIR[15].XIC[7].icell.PDM VGND.t774 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X85 VGND.t2407 XThC.Tn[11].t13 XA.XIR[6].XIC[11].icell.PDM VGND.t2406 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X86 VGND.t471 XThC.Tn[1].t13 XA.XIR[3].XIC[1].icell.PDM VGND.t470 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X87 XA.XIR[4].XIC[11].icell.Ien XThR.Tn[4].t13 VPWR.t1638 VPWR.t1637 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X88 VPWR.t1102 XThR.XTB6.Y a_n1049_5611# VPWR.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X89 XA.XIR[14].XIC[6].icell.PUM XThC.Tn[6].t13 XA.XIR[14].XIC[6].icell.Ien VPWR.t1874 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X90 VGND.t799 Vbias.t11 XA.XIR[9].XIC[7].icell.SM VGND.t798 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X91 VGND.t1326 XThC.Tn[2].t13 XA.XIR[6].XIC[2].icell.PDM VGND.t1325 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X92 XA.XIR[11].XIC[9].icell.Ien XThR.Tn[11].t14 VPWR.t1533 VPWR.t1532 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X93 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t1931 XA.XIR[6].XIC_dummy_left.icell.Ien VGND.t1515 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X94 VGND.t304 Vbias.t0 Vbias.t1 VGND.t303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X95 a_n1049_7787# XThR.XTB2.Y VPWR.t464 VPWR.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X96 VGND.t121 XThC.Tn[9].t13 XA.XIR[14].XIC[9].icell.PDM VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X97 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8].t12 XA.XIR[8].XIC[11].icell.Ien VGND.t1583 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X98 VGND.t801 Vbias.t12 XA.XIR[2].XIC[0].icell.SM VGND.t800 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X99 XA.XIR[1].XIC[1].icell.Ien XThR.Tn[1].t14 VPWR.t1562 VPWR.t1561 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X100 XA.XIR[13].XIC[4].icell.PUM XThC.Tn[4].t13 XA.XIR[13].XIC[4].icell.Ien VPWR.t1657 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X101 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t368 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t369 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X102 VGND.t803 Vbias.t13 XA.XIR[0].XIC[13].icell.SM VGND.t802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X103 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[0].t13 VGND.t755 VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X104 XA.XIR[4].XIC[2].icell.Ien XThR.Tn[4].t14 VPWR.t1640 VPWR.t1639 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X105 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[8].t13 VGND.t1585 VGND.t1584 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X106 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[8].t14 VGND.t1587 VGND.t1586 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X107 XA.XIR[3].XIC[3].icell.Ien XThR.Tn[3].t17 VPWR.t1397 VPWR.t1396 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X108 VGND.t2450 XThC.Tn[12].t12 XA.XIR[0].XIC[12].icell.PDM VGND.t2449 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X109 VPWR.t581 XThC.XTB3.Y.t3 a_4067_9615# VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[1].t15 XA.XIR[1].XIC[4].icell.Ien VGND.t1605 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X111 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5].t12 XA.XIR[5].XIC[1].icell.Ien VGND.t431 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X112 VPWR.t1671 data[4].t0 a_n1335_4229# VPWR.t1670 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X113 XA.XIR[2].XIC_15.icell.Ien XThR.Tn[2].t14 VPWR.t1491 VPWR.t1490 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X114 XA.XIR[3].XIC[9].icell.SM XA.XIR[3].XIC[9].icell.Ien Iout.t140 VGND.t931 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X115 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9].t14 XA.XIR[9].XIC[1].icell.Ien VGND.t438 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X116 VGND.t2388 XThR.XTBN.Y XThR.Tn[7].t7 VGND.t2387 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X117 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[4].t15 XA.XIR[4].XIC[5].icell.Ien VGND.t1770 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X118 a_n1319_5317# XThR.XTB7.A VPWR.t1535 VPWR.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X119 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8].t15 XA.XIR[8].XIC[2].icell.Ien VGND.t596 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X120 VPWR.t403 XThR.Tn[13].t12 XA.XIR[14].XIC[14].icell.PUM VPWR.t402 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X121 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11].t15 XA.XIR[11].XIC[3].icell.Ien VGND.t1239 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X122 XA.XIR[7].XIC[8].icell.PUM XThC.Tn[8].t12 XA.XIR[7].XIC[8].icell.Ien VPWR.t1144 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X123 XThC.Tn[9].t7 XThC.XTB2.Y VPWR.t1741 VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X124 XA.XIR[15].XIC[4].icell.Ien VPWR.t365 VPWR.t367 VPWR.t366 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X125 VGND.t805 Vbias.t14 XA.XIR[12].XIC[2].icell.SM VGND.t804 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X126 XA.XIR[6].XIC[4].icell.SM XA.XIR[6].XIC[4].icell.Ien Iout.t159 VGND.t1188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X127 VGND.t2051 Vbias.t15 XA.XIR[11].XIC_15.icell.SM VGND.t2050 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X128 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t362 VPWR.t364 VPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X129 XThC.Tn[5].t2 XThC.XTBN.Y.t11 VGND.t41 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X130 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout VGND.t1596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X131 VGND.t2053 Vbias.t16 XA.XIR[15].XIC[3].icell.SM VGND.t2052 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X132 VGND.t2055 Vbias.t17 XA.XIR[14].XIC[4].icell.SM VGND.t2054 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X133 VGND.t2548 XThC.Tn[6].t14 XA.XIR[6].XIC[6].icell.PDM VGND.t2547 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X134 VPWR.t840 XThR.Tn[8].t16 XA.XIR[9].XIC[4].icell.PUM VPWR.t839 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X135 VPWR.t1909 XThR.Tn[12].t15 XA.XIR[13].XIC[12].icell.PUM VPWR.t1908 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X136 VGND.t1076 VGND.t1074 XA.XIR[13].XIC_dummy_right.icell.SM VGND.t1075 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X137 XThR.Tn[9].t7 XThR.XTB2.Y a_n997_3755# VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X138 XThC.Tn[0].t9 XThC.XTBN.Y.t12 a_2979_9615# VPWR.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X139 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1932 VGND.t1517 VGND.t1516 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X140 XThC.Tn[5].t6 XThC.XTBN.Y.t13 a_5949_9615# VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X141 VGND.t145 XThC.XTB5.Y XThC.Tn[4].t2 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X142 XA.XIR[14].XIC[1].icell.PUM XThC.Tn[1].t14 XA.XIR[14].XIC[1].icell.Ien VPWR.t764 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X143 VGND.t2057 Vbias.t18 XA.XIR[9].XIC[2].icell.SM VGND.t2056 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X144 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t7 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X145 XA.XIR[13].XIC[0].icell.PUM XThC.Tn[0].t12 XA.XIR[13].XIC[0].icell.Ien VPWR.t987 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X146 XThC.Tn[7].t7 XThC.XTBN.Y.t14 VGND.t43 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X147 XThC.Tn[2].t8 XThC.XTBN.Y.t15 VGND.t44 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X148 VGND.t814 XThC.Tn[10].t13 XA.XIR[0].XIC[10].icell.PDM VGND.t813 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X149 a_n997_1579# XThR.XTBN.Y VGND.t2386 VGND.t2370 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X150 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[5].t13 VGND.t433 VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X151 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[5].t14 VGND.t691 VGND.t690 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X152 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t360 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X153 XA.XIR[9].XIC[14].icell.SM XA.XIR[9].XIC[14].icell.Ien Iout.t124 VGND.t886 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X154 VGND.t1804 XThC.Tn[4].t14 XA.XIR[14].XIC[4].icell.PDM VGND.t1803 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X155 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8].t17 XA.XIR[8].XIC[6].icell.Ien VGND.t597 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X156 XA.XIR[1].XIC[7].icell.PUM XThC.Tn[7].t9 XA.XIR[1].XIC[7].icell.Ien VPWR.t982 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X157 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[6].t16 VGND.t1670 VGND.t1669 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X158 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[1].t16 VGND.t1607 VGND.t1606 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X159 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11].t16 XA.XIR[11].XIC[7].icell.Ien VGND.t1240 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X160 XA.XIR[4].XIC[8].icell.PUM XThC.Tn[8].t13 XA.XIR[4].XIC[8].icell.Ien VPWR.t632 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X161 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[8].t18 VGND.t599 VGND.t598 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X162 XA.XIR[0].XIC_15.icell.SM XA.XIR[0].XIC_15.icell.Ien Iout.t75 VGND.t558 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X163 XA.XIR[4].XIC[12].icell.SM XA.XIR[4].XIC[12].icell.Ien Iout.t179 VGND.t1415 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X164 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[13].t13 VGND.t23 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X165 XA.XIR[11].XIC[12].icell.PUM XThC.Tn[12].t13 XA.XIR[11].XIC[12].icell.Ien VPWR.t1859 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X166 XA.XIR[12].XIC[4].icell.Ien XThR.Tn[12].t16 VPWR.t1911 VPWR.t1910 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X167 XA.XIR[3].XIC[4].icell.SM XA.XIR[3].XIC[4].icell.Ien Iout.t106 VGND.t772 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X168 XA.XIR[15].XIC[0].icell.Ien VPWR.t357 VPWR.t359 VPWR.t358 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X169 VGND.t2059 Vbias.t19 XA.XIR[8].XIC_15.icell.SM VGND.t2058 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X170 VGND.t853 XThC.Tn[14].t13 XA.XIR[8].XIC[14].icell.PDM VGND.t852 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X171 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t354 VPWR.t356 VPWR.t355 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X172 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[4].t16 XA.XIR[4].XIC[0].icell.Ien VGND.t1771 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X173 VGND.t306 XThC.Tn[8].t14 XA.XIR[8].XIC[8].icell.PDM VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X174 XA.XIR[14].XIC[14].icell.Ien XThR.Tn[14].t13 VPWR.t521 VPWR.t520 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X175 VGND.t46 XThC.XTBN.Y.t16 XThC.Tn[1].t7 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X176 VGND.t2061 Vbias.t20 XA.XIR[1].XIC[5].icell.SM VGND.t2060 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X177 VPWR.t1913 XThR.Tn[12].t17 XA.XIR[13].XIC[10].icell.PUM VPWR.t1912 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X178 XA.XIR[7].XIC[3].icell.PUM XThC.Tn[3].t13 XA.XIR[7].XIC[3].icell.Ien VPWR.t767 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X179 XA.XIR[2].XIC_15.icell.PUM VPWR.t352 XA.XIR[2].XIC_15.icell.Ien VPWR.t353 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X180 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[2].t15 XA.XIR[2].XIC[13].icell.Ien VGND.t810 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X181 VPWR.t720 XThR.Tn[9].t15 XA.XIR[10].XIC[12].icell.PUM VPWR.t719 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X182 VPWR.t842 XThR.Tn[8].t19 XA.XIR[9].XIC[0].icell.PUM VPWR.t841 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X183 VGND.t2063 Vbias.t21 XA.XIR[4].XIC[6].icell.SM VGND.t2062 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X184 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1933 VGND.t1519 VGND.t1518 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X185 VPWR.t351 VPWR.t349 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t350 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X186 VPWR.t426 XThC.XTBN.Y.t17 XThC.Tn[10].t0 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X187 VGND.t2385 XThR.XTBN.Y XThR.Tn[3].t8 VGND.t2348 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X188 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[2].t16 VGND.t809 VGND.t808 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X189 XA.XIR[6].XIC[8].icell.Ien XThR.Tn[6].t17 VPWR.t1582 VPWR.t1581 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X190 XThR.Tn[0].t5 XThR.XTBN.Y a_n1049_8581# VPWR.t1817 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X191 XA.XIR[13].XIC[12].icell.Ien XThR.Tn[13].t14 VPWR.t405 VPWR.t404 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X192 XA.XIR[13].XIC[7].icell.SM XA.XIR[13].XIC[7].icell.Ien Iout.t44 VGND.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X193 VPWR.t1133 VGND.t2688 XA.XIR[0].XIC[8].icell.PUM VPWR.t1132 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X194 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10].t13 XA.XIR[10].XIC[14].icell.Ien VGND.t657 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X195 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10].t14 XA.XIR[10].XIC[8].icell.Ien VGND.t1807 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X196 XThC.Tn[12].t2 XThC.XTB5.Y VPWR.t502 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 XA.XIR[1].XIC[11].icell.PUM XThC.Tn[11].t14 XA.XIR[1].XIC[11].icell.Ien VPWR.t1824 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X198 XThR.Tn[11].t7 XThR.XTBN.Y VPWR.t1816 VPWR.t1805 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 XA.XIR[0].XIC[7].icell.Ien XThR.Tn[0].t14 VPWR.t970 VPWR.t969 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X200 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[2].t17 VGND.t606 VGND.t605 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X201 XA.XIR[8].XIC[9].icell.PUM XThC.Tn[9].t14 XA.XIR[8].XIC[9].icell.Ien VPWR.t466 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X202 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[8].t20 VGND.t601 VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X203 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout VGND.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X204 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[5].t15 VGND.t693 VGND.t692 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X205 VGND.t2409 XThC.Tn[11].t15 XA.XIR[5].XIC[11].icell.PDM VGND.t2408 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X206 XA.XIR[11].XIC[10].icell.PUM XThC.Tn[10].t14 XA.XIR[11].XIC[10].icell.Ien VPWR.t1001 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X207 XThR.Tn[2].t7 XThR.XTBN.Y VGND.t2384 VGND.t2337 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X208 VGND.t2411 XThC.Tn[11].t16 XA.XIR[9].XIC[11].icell.PDM VGND.t2410 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X209 VGND.t1073 VGND.t1071 XA.XIR[13].XIC_dummy_left.icell.SM VGND.t1072 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X210 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12].t18 VPWR.t1915 VPWR.t1914 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X211 XA.XIR[1].XIC[2].icell.PUM XThC.Tn[2].t14 XA.XIR[1].XIC[2].icell.Ien VPWR.t1347 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X212 VPWR.t1815 XThR.XTBN.Y XThR.Tn[12].t11 VPWR.t1766 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X213 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[1].t17 VGND.t1609 VGND.t1608 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X214 XThC.XTB7.A data[0].t0 VPWR.t1374 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X215 VPWR.t722 XThR.Tn[9].t16 XA.XIR[10].XIC[10].icell.PUM VPWR.t721 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X216 XA.XIR[4].XIC[3].icell.PUM XThC.Tn[3].t14 XA.XIR[4].XIC[3].icell.Ien VPWR.t768 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X217 VGND.t2065 Vbias.t22 XA.XIR[4].XIC[10].icell.SM VGND.t2064 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X218 XA.XIR[0].XIC[13].icell.PDM VGND.t1068 VGND.t1070 VGND.t1069 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X219 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[13].t15 VGND.t25 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X220 VGND.t1521 VPWR.t1934 XA.XIR[0].XIC_dummy_left.icell.PDM VGND.t1520 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X221 VGND.t1328 XThC.Tn[2].t15 XA.XIR[5].XIC[2].icell.PDM VGND.t1327 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X222 VGND.t2067 Vbias.t23 XA.XIR[11].XIC[8].icell.SM VGND.t2066 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X223 XThC.Tn[9].t11 XThC.XTB2.Y a_7875_9569# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X224 VGND.t1774 XThC.Tn[5].t12 XA.XIR[1].XIC[5].icell.PDM VGND.t1773 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X225 XA.XIR[10].XIC[9].icell.Ien XThR.Tn[10].t15 VPWR.t1663 VPWR.t1662 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X226 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1935 VGND.t2140 VGND.t2139 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X227 VGND.t1330 XThC.Tn[2].t16 XA.XIR[9].XIC[2].icell.PDM VGND.t1329 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X228 VGND.t479 XThC.Tn[3].t15 XA.XIR[8].XIC[3].icell.PDM VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X229 VGND.t2142 VPWR.t1936 XA.XIR[3].XIC_15.icell.PDM VGND.t2141 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X230 a_n1319_5611# XThR.XTB6.A VPWR.t446 VPWR.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X231 XA.XIR[13].XIC[10].icell.Ien XThR.Tn[13].t16 VPWR.t407 VPWR.t406 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X232 VGND.t2383 XThR.XTBN.Y a_n997_3979# VGND.t2299 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X233 XA.XIR[15].XIC_15.icell.SM XA.XIR[15].XIC_15.icell.Ien Iout.t64 VGND.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X234 VPWR.t428 XThC.XTBN.Y.t18 XThC.Tn[14].t3 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X235 VGND.t2069 Vbias.t24 XA.XIR[1].XIC[0].icell.SM VGND.t2068 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X236 VPWR.t1917 XThR.Tn[12].t19 XA.XIR[13].XIC[5].icell.PUM VPWR.t1916 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X237 XA.XIR[12].XIC[4].icell.PUM XThC.Tn[4].t15 XA.XIR[12].XIC[4].icell.Ien VPWR.t1658 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X238 VGND.t2071 Vbias.t25 XA.XIR[4].XIC[1].icell.SM VGND.t2070 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X239 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7].t8 XA.XIR[7].XIC[14].icell.Ien VGND.t584 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X240 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7].t9 XA.XIR[7].XIC[8].icell.Ien VGND.t585 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X241 XA.XIR[0].XIC[11].icell.Ien XThR.Tn[0].t15 VPWR.t972 VPWR.t971 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X242 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[2].t18 VGND.t604 VGND.t603 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X243 XA.XIR[6].XIC[3].icell.Ien XThR.Tn[6].t18 VPWR.t1584 VPWR.t1583 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X244 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14].t14 XA.XIR[14].XIC[12].icell.Ien VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X245 XA.XIR[11].XIC[6].icell.SM XA.XIR[11].XIC[6].icell.Ien Iout.t161 VGND.t1249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X246 XA.XIR[1].XIC_15.icell.Ien XThR.Tn[1].t18 VPWR.t1564 VPWR.t1563 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X247 VGND.t2073 Vbias.t26 XA.XIR[2].XIC[14].icell.SM VGND.t2072 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X248 VGND.t683 XThC.Tn[13].t13 XA.XIR[2].XIC[13].icell.PDM VGND.t682 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X249 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[5].t16 VGND.t695 VGND.t694 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X250 VPWR.t1862 XThR.XTB4.Y.t2 a_n1049_6699# VPWR.t680 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X251 VGND.t2144 VPWR.t1937 XA.XIR[15].XIC_dummy_right.icell.PDM VGND.t2143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X252 XA.XIR[13].XIC[2].icell.SM XA.XIR[13].XIC[2].icell.Ien Iout.t147 VGND.t1121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X253 VPWR.t1131 VGND.t2689 XA.XIR[0].XIC[3].icell.PUM VPWR.t1130 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X254 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10].t16 XA.XIR[10].XIC[3].icell.Ien VGND.t1808 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X255 VPWR.t1412 XThC.XTB6.Y a_5949_9615# VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X256 VPWR.t559 XThR.XTB1.Y.t3 a_n1049_8581# VPWR.t558 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X257 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5].t17 XA.XIR[5].XIC_15.icell.Ien VGND.t696 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X258 VPWR.t1283 XThR.Tn[11].t17 XA.XIR[12].XIC[7].icell.PUM VPWR.t1282 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X259 XA.XIR[0].XIC[2].icell.Ien XThR.Tn[0].t16 VPWR.t974 VPWR.t973 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X260 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9].t17 XA.XIR[9].XIC_15.icell.Ien VGND.t439 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X261 XA.XIR[0].XIC[8].icell.SM XA.XIR[0].XIC[8].icell.Ien Iout.t81 VGND.t609 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X262 VGND.t485 Vbias.t27 XA.XIR[5].XIC[7].icell.SM VGND.t484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X263 XA.XIR[11].XIC[5].icell.PUM XThC.Tn[5].t13 XA.XIR[11].XIC[5].icell.Ien VPWR.t1641 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X264 VGND.t2550 XThC.Tn[6].t15 XA.XIR[5].XIC[6].icell.PDM VGND.t2549 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X265 VGND.t2294 XThR.XTB7.B a_n1335_8107# VGND.t2288 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X266 VPWR.t832 XThR.Tn[7].t10 XA.XIR[8].XIC[4].icell.PUM VPWR.t831 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X267 XA.XIR[0].XIC[5].icell.PDM XThR.Tn[0].t17 XA.XIR[0].XIC[5].icell.Ien VGND.t756 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X268 VPWR.t348 VPWR.t346 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t347 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X269 VGND.t2552 XThC.Tn[6].t16 XA.XIR[9].XIC[6].icell.PDM VGND.t2551 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X270 VGND.t487 Vbias.t28 XA.XIR[8].XIC[8].icell.SM VGND.t486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X271 XA.XIR[7].XIC[9].icell.Ien XThR.Tn[7].t11 VPWR.t834 VPWR.t833 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X272 XThC.XTB4.Y.t0 XThC.XTB7.B VPWR.t1217 VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X273 VGND.t1067 VGND.t1065 XA.XIR[12].XIC_dummy_right.icell.SM VGND.t1066 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X274 VGND.t777 XThC.Tn[7].t10 XA.XIR[8].XIC[7].icell.PDM VGND.t776 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X275 VPWR.t345 VPWR.t343 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X276 XThR.Tn[2].t1 XThR.XTB3.Y.t3 VGND.t376 VGND.t375 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X277 VGND.t2382 XThR.XTBN.Y a_n997_2891# VGND.t2333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X278 VPWR.t724 XThR.Tn[9].t18 XA.XIR[10].XIC[5].icell.PUM VPWR.t723 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X279 XA.XIR[5].XIC[5].icell.SM XA.XIR[5].XIC[5].icell.Ien Iout.t104 VGND.t770 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X280 VPWR.t682 XThR.XTB5.Y XThR.Tn[12].t3 VPWR.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X281 XA.XIR[12].XIC[0].icell.PUM XThC.Tn[0].t13 XA.XIR[12].XIC[0].icell.Ien VPWR.t988 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X282 VGND.t783 XThC.Tn[0].t14 XA.XIR[1].XIC[0].icell.PDM VGND.t782 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X283 VGND.t489 Vbias.t29 XA.XIR[11].XIC[3].icell.SM VGND.t488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X284 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14].t15 XA.XIR[14].XIC[10].icell.Ien VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X285 XA.XIR[11].XIC[10].icell.SM XA.XIR[11].XIC[10].icell.Ien Iout.t89 VGND.t661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X286 VGND.t2381 XThR.XTBN.Y XThR.Tn[6].t11 VGND.t2380 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X287 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[11].t18 VGND.t1242 VGND.t1241 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X288 VPWR.t1814 XThR.XTBN.Y XThR.Tn[9].t10 VPWR.t1800 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X289 XA.XIR[8].XIC[6].icell.SM XA.XIR[8].XIC[6].icell.Ien Iout.t32 VGND.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X290 XA.XIR[13].XIC[5].icell.Ien XThR.Tn[13].t17 VPWR.t409 VPWR.t408 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X291 VGND.t1064 VGND.t1062 XA.XIR[9].XIC_dummy_right.icell.SM VGND.t1063 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X292 XA.XIR[14].XIC_15.icell.PUM VPWR.t341 XA.XIR[14].XIC_15.icell.Ien VPWR.t342 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X293 a_n997_715# XThR.XTBN.Y VGND.t2379 VGND.t2378 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X294 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10].t17 XA.XIR[10].XIC[7].icell.Ien VGND.t1809 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X295 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7].t12 XA.XIR[7].XIC[3].icell.Ien VGND.t586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X296 XThC.Tn[1].t6 XThC.XTBN.Y.t19 VGND.t47 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X297 VPWR.t1285 XThR.Tn[11].t19 XA.XIR[12].XIC[11].icell.PUM VPWR.t1284 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X298 XA.XIR[6].XIC[4].icell.PUM XThC.Tn[4].t16 XA.XIR[6].XIC[4].icell.Ien VPWR.t1659 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X299 XThR.Tn[14].t3 XThR.XTB7.Y VPWR.t1369 VPWR.t1087 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X300 XA.XIR[10].XIC[12].icell.PUM XThC.Tn[12].t14 XA.XIR[10].XIC[12].icell.Ien VPWR.t1860 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X301 XA.XIR[2].XIC[5].icell.SM XA.XIR[2].XIC[5].icell.Ien Iout.t109 VGND.t779 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X302 XA.XIR[11].XIC[1].icell.SM XA.XIR[11].XIC[1].icell.Ien Iout.t127 VGND.t897 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X303 XA.XIR[7].XIC_15.icell.PDM VPWR.t1938 VGND.t2146 VGND.t2145 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X304 XA.XIR[6].XIC[13].icell.SM XA.XIR[6].XIC[13].icell.Ien Iout.t182 VGND.t1419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X305 XA.XIR[13].XIC[13].icell.PUM XThC.Tn[13].t14 XA.XIR[13].XIC[13].icell.Ien VPWR.t903 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X306 VGND.t491 Vbias.t30 XA.XIR[15].XIC[12].icell.SM VGND.t490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X307 VGND.t493 Vbias.t31 XA.XIR[14].XIC[13].icell.SM VGND.t492 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X308 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[2].t19 XA.XIR[2].XIC[1].icell.Ien VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X309 VPWR.t836 XThR.Tn[7].t13 XA.XIR[8].XIC[0].icell.PUM VPWR.t835 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X310 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[1].t19 XA.XIR[1].XIC[13].icell.Ien VGND.t1610 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X311 VPWR.t681 XThR.XTB5.Y a_n1049_6405# VPWR.t680 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X312 VPWR.t1287 XThR.Tn[11].t20 XA.XIR[12].XIC[2].icell.PUM VPWR.t1286 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X313 XThR.XTB7.B data[6].t0 VPWR.t976 VPWR.t975 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X314 XA.XIR[0].XIC[8].icell.PUM XThC.Tn[8].t15 XA.XIR[0].XIC[8].icell.Ien VPWR.t633 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X315 VPWR.t981 XThC.XTB4.Y.t3 a_4861_9615# VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X316 XA.XIR[0].XIC[3].icell.SM XA.XIR[0].XIC[3].icell.Ien Iout.t51 VGND.t264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X317 VGND.t495 Vbias.t32 XA.XIR[5].XIC[2].icell.SM VGND.t494 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X318 XA.XIR[8].XIC[4].icell.Ien XThR.Tn[8].t21 VPWR.t844 VPWR.t843 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X319 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t338 VPWR.t340 VPWR.t339 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X320 VGND.t106 XThR.XTB2.Y XThR.Tn[1].t3 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X321 XA.XIR[0].XIC[0].icell.PDM XThR.Tn[0].t18 XA.XIR[0].XIC[0].icell.Ien VGND.t757 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X322 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[11].t21 VGND.t1244 VGND.t1243 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X323 XA.XIR[12].XIC[7].icell.SM XA.XIR[12].XIC[7].icell.Ien Iout.t34 VGND.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X324 XThR.XTB7.A data[4].t1 a_n1331_2891# VGND.t1815 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X325 XA.XIR[8].XIC[10].icell.SM XA.XIR[8].XIC[10].icell.Ien Iout.t190 VGND.t1501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X326 VGND.t497 Vbias.t33 XA.XIR[8].XIC[3].icell.SM VGND.t496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X327 XA.XIR[15].XIC[13].icell.Ien VPWR.t335 VPWR.t337 VPWR.t336 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X328 XA.XIR[15].XIC[8].icell.SM XA.XIR[15].XIC[8].icell.Ien Iout.t201 VGND.t1580 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X329 VPWR.t908 XThR.Tn[5].t18 XA.XIR[6].XIC[12].icell.PUM VPWR.t907 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X330 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1939 XA.XIR[11].XIC_dummy_right.icell.Ien VGND.t2147 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X331 VPWR.t942 XThR.Tn[8].t22 XA.XIR[9].XIC[13].icell.PUM VPWR.t941 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X332 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7].t14 XA.XIR[7].XIC[7].icell.Ien VGND.t587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X333 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t7 VPWR.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X334 XA.XIR[5].XIC[0].icell.SM XA.XIR[5].XIC[0].icell.Ien Iout.t146 VGND.t1120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X335 XA.XIR[10].XIC[10].icell.PUM XThC.Tn[10].t15 XA.XIR[10].XIC[10].icell.Ien VPWR.t1002 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X336 VGND.t1202 XThC.XTBN.Y.t20 XThC.Tn[4].t11 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X337 XA.XIR[6].XIC[0].icell.PUM XThC.Tn[0].t15 XA.XIR[6].XIC[0].icell.Ien VPWR.t989 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X338 XA.XIR[8].XIC[1].icell.SM XA.XIR[8].XIC[1].icell.Ien Iout.t60 VGND.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X339 XA.XIR[3].XIC[13].icell.SM XA.XIR[3].XIC[13].icell.Ien Iout.t114 VGND.t827 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X340 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t333 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t334 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X341 VGND.t1061 VGND.t1059 XA.XIR[12].XIC_dummy_left.icell.SM VGND.t1060 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X342 XThC.XTB5.A data[1].t0 a_7331_10587# VPWR.t1047 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X343 VGND.t1843 data[1].t1 a_8739_10571# VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X344 XA.XIR[0].XIC[1].icell.PDM VGND.t1056 VGND.t1058 VGND.t1057 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X345 VPWR.t462 XThR.XTB2.Y XThR.Tn[9].t3 VPWR.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X346 VGND.t2377 XThR.XTBN.Y XThR.Tn[7].t6 VGND.t2376 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X347 VGND.t685 XThC.Tn[13].t15 XA.XIR[14].XIC[13].icell.PDM VGND.t684 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X348 XA.XIR[2].XIC[0].icell.SM XA.XIR[2].XIC[0].icell.Ien Iout.t158 VGND.t1187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X349 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1940 XA.XIR[14].XIC_dummy_left.icell.Ien VGND.t2148 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X350 XThR.Tn[13].t11 XThR.XTBN.Y VPWR.t1813 VPWR.t1776 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X351 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[10].t18 VGND.t1811 VGND.t1810 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X352 XA.XIR[14].XIC_15.icell.SM XA.XIR[14].XIC_15.icell.Ien Iout.t33 VGND.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X353 VGND.t499 Vbias.t34 XA.XIR[10].XIC[11].icell.SM VGND.t498 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X354 VGND.t1055 VGND.t1053 XA.XIR[9].XIC_dummy_left.icell.SM VGND.t1054 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X355 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8].t23 VPWR.t944 VPWR.t943 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X356 VPWR.t1489 XThR.Tn[2].t20 XA.XIR[3].XIC[9].icell.PUM VPWR.t1488 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X357 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t330 VPWR.t332 VPWR.t331 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X358 XA.XIR[12].XIC[13].icell.Ien XThR.Tn[12].t20 VPWR.t1919 VPWR.t1918 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X359 VPWR.t1586 XThR.Tn[6].t19 XA.XIR[7].XIC[9].icell.PUM VPWR.t1585 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X360 XA.XIR[0].XIC[3].icell.PUM XThC.Tn[3].t16 XA.XIR[0].XIC[3].icell.Ien VPWR.t769 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X361 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t327 VPWR.t329 VPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X362 VPWR.t910 XThR.Tn[5].t19 XA.XIR[6].XIC[10].icell.PUM VPWR.t909 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X363 VGND.t473 XThC.Tn[1].t15 XA.XIR[2].XIC[1].icell.PDM VGND.t472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X364 VGND.t937 XThR.XTB6.Y XThR.Tn[5].t3 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X365 XA.XIR[13].XIC[6].icell.PUM XThC.Tn[6].t17 XA.XIR[13].XIC[6].icell.Ien VPWR.t1875 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X366 XThR.Tn[9].t6 XThR.XTB2.Y a_n997_3755# VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X367 VGND.t501 Vbias.t35 XA.XIR[1].XIC[14].icell.SM VGND.t500 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X368 XThR.XTB6.Y XThR.XTB6.A VGND.t95 VGND.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X369 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t1941 VGND.t2150 VGND.t2149 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X370 XA.XIR[12].XIC[2].icell.SM XA.XIR[12].XIC[2].icell.Ien Iout.t197 VGND.t1576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X371 a_n997_1579# XThR.XTBN.Y VGND.t2375 VGND.t2365 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X372 VGND.t123 XThC.Tn[9].t15 XA.XIR[13].XIC[9].icell.PDM VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X373 XA.XIR[15].XIC[3].icell.SM XA.XIR[15].XIC[3].icell.Ien Iout.t50 VGND.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X374 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[3].t18 XA.XIR[3].XIC[14].icell.Ien VGND.t1444 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X375 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[3].t19 XA.XIR[3].XIC[8].icell.Ien VGND.t1445 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X376 VPWR.t523 XThR.Tn[14].t16 XA.XIR[15].XIC[7].icell.PUM VPWR.t522 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X377 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t325 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t326 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X378 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout VGND.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X379 VPWR.t411 XThR.Tn[13].t18 XA.XIR[14].XIC[8].icell.PUM VPWR.t410 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X380 XA.XIR[10].XIC[5].icell.PUM XThC.Tn[5].t14 XA.XIR[10].XIC[5].icell.Ien VPWR.t1642 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X381 XA.XIR[15].XIC[6].icell.Ien VPWR.t322 VPWR.t324 VPWR.t323 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X382 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t1942 VGND.t2152 VGND.t2151 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X383 VGND.t503 Vbias.t36 XA.XIR[10].XIC[9].icell.SM VGND.t502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X384 VPWR.t1921 XThR.Tn[12].t21 XA.XIR[13].XIC[14].icell.PUM VPWR.t1920 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X385 VPWR.t946 XThR.Tn[8].t24 XA.XIR[9].XIC[6].icell.PUM VPWR.t945 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X386 XA.XIR[15].XIC[9].icell.PDM VPWR.t1943 XA.XIR[15].XIC[9].icell.Ien VGND.t2153 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X387 XA.XIR[3].XIC[9].icell.Ien XThR.Tn[3].t20 VPWR.t389 VPWR.t388 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X388 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[10].t19 VGND.t1813 VGND.t1812 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X389 XA.XIR[15].XIC[12].icell.PDM XThR.Tn[14].t17 VGND.t170 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X390 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1944 VGND.t2155 VGND.t2154 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X391 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[13].t19 VGND.t27 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X392 VPWR.t1293 XThR.XTBN.A XThR.XTBN.Y VPWR.t1292 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X393 VPWR.t912 XThR.Tn[5].t20 XA.XIR[6].XIC[5].icell.PUM VPWR.t911 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X394 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[4].t17 XA.XIR[4].XIC[11].icell.Ien VGND.t1772 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X395 XA.XIR[5].XIC[4].icell.PUM XThC.Tn[4].t17 XA.XIR[5].XIC[4].icell.Ien VPWR.t1660 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X396 VPWR.t525 XThR.Tn[14].t18 XA.XIR[15].XIC[11].icell.PUM VPWR.t524 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X397 XA.XIR[1].XIC[5].icell.SM XA.XIR[1].XIC[5].icell.Ien Iout.t208 VGND.t1805 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X398 XA.XIR[13].XIC[1].icell.PUM XThC.Tn[1].t16 XA.XIR[13].XIC[1].icell.Ien VPWR.t765 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X399 XA.XIR[9].XIC[4].icell.PUM XThC.Tn[4].t18 XA.XIR[9].XIC[4].icell.Ien VPWR.t1661 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X400 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t320 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t321 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X401 a_3523_10575# XThC.XTB7.B VGND.t1183 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X402 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[4].t18 VGND.t1310 VGND.t1309 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X403 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[4].t19 VGND.t1312 VGND.t1311 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X404 XA.XIR[12].XIC[13].icell.PUM XThC.Tn[13].t16 XA.XIR[12].XIC[13].icell.Ien VPWR.t904 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X405 XA.XIR[4].XIC[6].icell.SM XA.XIR[4].XIC[6].icell.Ien Iout.t17 VGND.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X406 XA.XIR[11].XIC[14].icell.PUM XThC.Tn[14].t14 XA.XIR[11].XIC[14].icell.Ien VPWR.t1039 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X407 VPWR.t1222 XThC.XTBN.Y.t21 XThC.Tn[13].t3 VPWR.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[1].t20 XA.XIR[1].XIC[1].icell.Ien VGND.t1611 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X409 VGND.t505 Vbias.t37 XA.XIR[13].XIC[5].icell.SM VGND.t504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X410 VGND.t759 XThC.Tn[4].t19 XA.XIR[13].XIC[4].icell.PDM VGND.t758 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X411 XA.XIR[12].XIC[6].icell.Ien XThR.Tn[12].t22 VPWR.t1923 VPWR.t1922 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X412 XThC.Tn[5].t11 XThC.XTB6.Y VGND.t1460 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 XThC.Tn[4].t1 XThC.XTB5.Y VGND.t144 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X414 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[4].t20 XA.XIR[4].XIC[2].icell.Ien VGND.t1313 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X415 VGND.t2157 VPWR.t1945 XA.XIR[8].XIC_dummy_right.icell.PDM VGND.t2156 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X416 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[3].t21 XA.XIR[3].XIC[3].icell.Ien VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X417 XA.XIR[14].XIC[8].icell.Ien XThR.Tn[14].t19 VPWR.t527 VPWR.t526 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X418 VPWR.t529 XThR.Tn[14].t20 XA.XIR[15].XIC[2].icell.PUM VPWR.t528 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X419 XA.XIR[2].XIC_15.icell.PDM XThR.Tn[2].t21 XA.XIR[2].XIC_15.icell.Ien VGND.t112 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X420 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t7 VGND.t351 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X421 VPWR.t413 XThR.Tn[13].t20 XA.XIR[14].XIC[3].icell.PUM VPWR.t412 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X422 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12].t23 XA.XIR[12].XIC[9].icell.Ien VGND.t2686 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X423 VPWR.t726 XThR.Tn[9].t19 XA.XIR[10].XIC[14].icell.PUM VPWR.t725 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X424 XA.XIR[15].XIC[1].icell.Ien VPWR.t314 VPWR.t316 VPWR.t315 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X425 VGND.t507 Vbias.t38 XA.XIR[11].XIC[12].icell.SM VGND.t506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X426 VGND.t51 Vbias.t39 XA.XIR[7].XIC_15.icell.SM VGND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X427 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t317 VPWR.t319 VPWR.t318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X428 VGND.t855 XThC.Tn[14].t15 XA.XIR[7].XIC[14].icell.PDM VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X429 VGND.t308 XThC.Tn[8].t16 XA.XIR[7].XIC[8].icell.PDM VGND.t307 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X430 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t10 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X431 XThC.Tn[4].t10 XThC.XTBN.Y.t22 VGND.t1203 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X432 VPWR.t1202 XThR.Tn[0].t19 XA.XIR[1].XIC[4].icell.PUM VPWR.t1201 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X433 a_n1049_5317# XThR.XTB7.Y VPWR.t1368 VPWR.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X434 XA.XIR[13].XIC[14].icell.Ien XThR.Tn[13].t21 VPWR.t415 VPWR.t414 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X435 XA.XIR[14].XIC[8].icell.SM XA.XIR[14].XIC[8].icell.Ien Iout.t240 VGND.t2418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X436 XA.XIR[15].XIC[10].icell.PDM XThR.Tn[14].t21 VGND.t172 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X437 VGND.t53 Vbias.t40 XA.XIR[10].XIC[4].icell.SM VGND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X438 VGND.t1052 VGND.t1050 XA.XIR[5].XIC_dummy_right.icell.SM VGND.t1051 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X439 VPWR.t948 XThR.Tn[8].t25 XA.XIR[9].XIC[1].icell.PUM VPWR.t947 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X440 VPWR.t1336 XThR.Tn[4].t21 XA.XIR[5].XIC[4].icell.PUM VPWR.t1335 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X441 XThC.XTB6.Y XThC.XTB7.B VGND.t1182 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X442 VPWR.t313 VPWR.t311 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t312 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X443 XA.XIR[15].XIC[4].icell.PDM VPWR.t1946 XA.XIR[15].XIC[4].icell.Ien VGND.t2158 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X444 VPWR.t931 XThR.Tn[7].t15 XA.XIR[8].XIC[13].icell.PUM VPWR.t930 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X445 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t1947 XA.XIR[10].XIC_dummy_right.icell.Ien VGND.t2159 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X446 a_6243_9615# XThC.XTBN.Y.t23 XThC.Tn[6].t7 VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X447 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout VGND.t1111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X448 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[1].t21 VGND.t1981 VGND.t1980 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X449 XA.XIR[5].XIC[0].icell.PUM XThC.Tn[0].t16 XA.XIR[5].XIC[0].icell.Ien VPWR.t990 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X450 XA.XIR[4].XIC[10].icell.SM XA.XIR[4].XIC[10].icell.Ien Iout.t14 VGND.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X451 XA.XIR[9].XIC[0].icell.PUM XThC.Tn[0].t17 XA.XIR[9].XIC[0].icell.Ien VPWR.t991 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X452 XThC.Tn[13].t7 XThC.XTB6.Y VPWR.t1411 VPWR.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X453 XA.XIR[5].XIC[14].icell.SM XA.XIR[5].XIC[14].icell.Ien Iout.t42 VGND.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X454 VGND.t1204 XThC.XTBN.Y.t24 XThC.Tn[0].t6 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X455 XThR.Tn[3].t4 XThR.XTBN.Y a_n1049_6699# VPWR.t1812 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X456 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[4].t22 XA.XIR[4].XIC[6].icell.Ien VGND.t1314 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X457 VGND.t475 XThC.Tn[1].t17 XA.XIR[14].XIC[1].icell.PDM VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X458 VGND.t2494 XThR.XTB4.Y.t3 XThR.Tn[3].t9 VGND.t858 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X459 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[3].t22 XA.XIR[3].XIC[7].icell.Ien VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X460 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[1].t22 VGND.t1983 VGND.t1982 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X461 XA.XIR[7].XIC[9].icell.PUM XThC.Tn[9].t16 XA.XIR[7].XIC[9].icell.Ien VPWR.t467 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X462 XA.XIR[1].XIC[0].icell.SM XA.XIR[1].XIC[0].icell.Ien Iout.t254 VGND.t2673 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X463 XA.XIR[3].XIC[12].icell.PUM XThC.Tn[12].t15 XA.XIR[3].XIC[12].icell.Ien VPWR.t1861 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X464 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[4].t23 VGND.t1316 VGND.t1315 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X465 XA.XIR[0].XIC[12].icell.SM XA.XIR[0].XIC[12].icell.Ien Iout.t2 VGND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X466 XA.XIR[0].XIC_15.icell.PDM VPWR.t1948 VGND.t2161 VGND.t2160 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X467 XA.XIR[4].XIC[1].icell.SM XA.XIR[4].XIC[1].icell.Ien Iout.t149 VGND.t1133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X468 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[9].t20 VGND.t441 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X469 VGND.t55 Vbias.t41 XA.XIR[13].XIC[0].icell.SM VGND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X470 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12].t24 VPWR.t1925 VPWR.t1924 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X471 XA.XIR[6].XIC[13].icell.PUM XThC.Tn[13].t17 XA.XIR[6].XIC[13].icell.Ien VPWR.t905 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X472 VGND.t57 Vbias.t42 XA.XIR[8].XIC[12].icell.SM VGND.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X473 XA.XIR[2].XIC[14].icell.SM XA.XIR[2].XIC[14].icell.Ien Iout.t3 VGND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X474 XThR.Tn[11].t8 XThR.XTB4.Y.t4 VPWR.t1863 VPWR.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X475 VGND.t310 XThC.Tn[8].t17 XA.XIR[4].XIC[8].icell.PDM VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X476 VGND.t857 XThC.Tn[14].t16 XA.XIR[4].XIC[14].icell.PDM VGND.t856 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X477 XThC.Tn[14].t11 XThC.XTB7.Y a_10915_9569# VGND.t1176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X478 VPWR.t1204 XThR.Tn[0].t20 XA.XIR[1].XIC[0].icell.PUM VPWR.t1203 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X479 XA.XIR[14].XIC[3].icell.Ien XThR.Tn[14].t22 VPWR.t531 VPWR.t530 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X480 VGND.t2452 XThC.Tn[12].t16 XA.XIR[11].XIC[12].icell.PDM VGND.t2451 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X481 VPWR.t1338 XThR.Tn[4].t24 XA.XIR[5].XIC[0].icell.PUM VPWR.t1337 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X482 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12].t25 XA.XIR[12].XIC[4].icell.Ien VGND.t911 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X483 XA.XIR[12].XIC[6].icell.PUM XThC.Tn[6].t18 XA.XIR[12].XIC[6].icell.Ien VPWR.t1876 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X484 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t1949 XA.XIR[7].XIC_dummy_right.icell.Ien VGND.t2162 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X485 VPWR.t310 VPWR.t308 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t309 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X486 XA.XIR[15].XIC[7].icell.PUM XThC.Tn[7].t11 XA.XIR[15].XIC[7].icell.Ien VPWR.t983 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X487 VGND.t2074 XThC.XTB4.Y.t4 XThC.Tn[3].t11 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X488 VPWR.t1740 XThC.XTB2.Y XThC.Tn[9].t6 VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X489 XA.XIR[5].XIC[12].icell.Ien XThR.Tn[5].t21 VPWR.t914 VPWR.t913 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X490 VGND.t481 XThC.Tn[3].t17 XA.XIR[7].XIC[3].icell.PDM VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X491 VGND.t59 Vbias.t43 XA.XIR[6].XIC[11].icell.SM VGND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X492 VGND.t2164 VPWR.t1950 XA.XIR[2].XIC_15.icell.PDM VGND.t2163 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X493 VPWR.t679 XThR.XTB5.Y XThR.Tn[12].t2 VPWR.t576 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 VGND.t125 XThC.Tn[9].t17 XA.XIR[12].XIC[9].icell.PDM VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X495 XA.XIR[14].XIC[3].icell.SM XA.XIR[14].XIC[3].icell.Ien Iout.t155 VGND.t1145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X496 XA.XIR[9].XIC[12].icell.Ien XThR.Tn[9].t21 VPWR.t728 VPWR.t727 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X497 XA.XIR[8].XIC[13].icell.Ien XThR.Tn[8].t26 VPWR.t950 VPWR.t949 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X498 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout VGND.t1338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X499 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6].t20 XA.XIR[6].XIC[14].icell.Ien VGND.t1671 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X500 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6].t21 XA.XIR[6].XIC[8].icell.Ien VGND.t1672 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X501 VPWR.t1367 XThR.XTB7.Y XThR.Tn[14].t2 VPWR.t1093 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X502 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[1].t23 VGND.t1985 VGND.t1984 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X503 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13].t22 XA.XIR[13].XIC[12].icell.Ien VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X504 XA.XIR[4].XIC[9].icell.PUM XThC.Tn[9].t18 XA.XIR[4].XIC[9].icell.Ien VPWR.t468 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X505 XThR.Tn[8].t3 XThR.XTB1.Y.t4 a_n997_3979# VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X506 XA.XIR[3].XIC[10].icell.PUM XThC.Tn[10].t16 XA.XIR[3].XIC[10].icell.Ien VPWR.t1003 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X507 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[4].t25 VGND.t1600 VGND.t1599 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X508 VGND.t2413 XThC.Tn[11].t17 XA.XIR[1].XIC[11].icell.PDM VGND.t2412 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X509 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1951 VGND.t2166 VGND.t2165 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X510 VPWR.t933 XThR.Tn[7].t16 XA.XIR[8].XIC[6].icell.PUM VPWR.t932 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X511 VPWR.t1072 data[2].t0 XThC.XTB7.B VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X512 VGND.t1049 VGND.t1047 XA.XIR[5].XIC_dummy_left.icell.SM VGND.t1048 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X513 VPWR.t1665 XThR.Tn[10].t20 XA.XIR[11].XIC[7].icell.PUM VPWR.t1664 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X514 VGND.t816 XThC.Tn[10].t17 XA.XIR[11].XIC[10].icell.PDM VGND.t815 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X515 XThC.Tn[13].t10 XThC.XTB6.Y a_10051_9569# VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X516 XThR.Tn[4].t7 XThR.XTBN.Y a_n1049_6405# VPWR.t1812 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X517 XThR.XTB5.Y XThR.XTB7.B a_n1319_6405# VPWR.t1752 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X518 VGND.t61 Vbias.t44 XA.XIR[4].XIC[7].icell.SM VGND.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X519 XThC.Tn[8].t3 XThC.XTBN.Y.t25 VPWR.t1224 VPWR.t1223 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X520 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[13].t23 VGND.t33 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X521 XA.XIR[15].XIC[11].icell.PUM XThC.Tn[11].t18 XA.XIR[15].XIC[11].icell.Ien VPWR.t1825 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X522 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[9].t22 VGND.t443 VGND.t442 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X523 a_n1335_4229# data[5].t0 XThR.XTB5.A VPWR.t1536 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X524 VGND.t1523 XThC.Tn[2].t17 XA.XIR[1].XIC[2].icell.PDM VGND.t1522 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X525 VGND.t63 Vbias.t45 XA.XIR[7].XIC[8].icell.SM VGND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X526 XA.XIR[6].XIC[9].icell.Ien XThR.Tn[6].t22 VPWR.t1588 VPWR.t1587 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X527 XA.XIR[5].XIC[10].icell.Ien XThR.Tn[5].t22 VPWR.t916 VPWR.t915 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X528 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[12].t26 VGND.t913 VGND.t912 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X529 VGND.t649 XThC.Tn[7].t12 XA.XIR[7].XIC[7].icell.PDM VGND.t648 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X530 VGND.t65 Vbias.t46 XA.XIR[6].XIC[9].icell.SM VGND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X531 VGND.t67 Vbias.t47 XA.XIR[3].XIC[11].icell.SM VGND.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X532 XThC.Tn[8].t10 XThC.XTB1.Y.t4 a_7651_9569# VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X533 XThC.Tn[13].t2 XThC.XTBN.Y.t26 VPWR.t1225 VPWR.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X534 VGND.t483 XThC.Tn[3].t18 XA.XIR[4].XIC[3].icell.PDM VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X535 XA.XIR[9].XIC[10].icell.Ien XThR.Tn[9].t23 VPWR.t730 VPWR.t729 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X536 XA.XIR[7].XIC_15.icell.SM XA.XIR[7].XIC_15.icell.Ien Iout.t20 VGND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X537 XA.XIR[15].XIC[12].icell.SM XA.XIR[15].XIC[12].icell.Ien Iout.t21 VGND.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X538 VPWR.t1129 VGND.t2690 XA.XIR[0].XIC[9].icell.PUM VPWR.t1128 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X539 VGND.t1459 XThC.XTB6.Y XThC.Tn[5].t10 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X540 XA.XIR[12].XIC[1].icell.PUM XThC.Tn[1].t18 XA.XIR[12].XIC[1].icell.Ien VPWR.t766 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X541 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t305 VPWR.t307 VPWR.t306 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X542 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[3].t23 VGND.t6 VGND.t5 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X543 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[3].t24 VGND.t8 VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X544 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13].t24 XA.XIR[13].XIC[10].icell.Ien VGND.t34 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X545 XA.XIR[15].XIC[2].icell.PUM XThC.Tn[2].t18 XA.XIR[15].XIC[2].icell.Ien VPWR.t1429 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X546 XA.XIR[6].XIC[6].icell.PUM XThC.Tn[6].t19 XA.XIR[6].XIC[6].icell.Ien VPWR.t1877 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X547 XA.XIR[10].XIC[14].icell.PUM XThC.Tn[14].t17 XA.XIR[10].XIC[14].icell.Ien VPWR.t1040 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X548 VGND.t69 Vbias.t48 XA.XIR[12].XIC[5].icell.SM VGND.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X549 VGND.t761 XThC.Tn[4].t20 XA.XIR[12].XIC[4].icell.PDM VGND.t760 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X550 a_n1049_5611# XThR.XTB6.Y VPWR.t1100 VPWR.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X551 XA.XIR[13].XIC_15.icell.PUM VPWR.t303 XA.XIR[13].XIC_15.icell.Ien VPWR.t304 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X552 XThR.Tn[10].t6 XThR.XTB3.Y.t4 a_n997_2891# VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X553 VGND.t71 Vbias.t49 XA.XIR[15].XIC[6].icell.SM VGND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X554 XA.XIR[0].XIC[11].icell.PDM XThR.Tn[0].t21 XA.XIR[0].XIC[11].icell.Ien VGND.t1158 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X555 VGND.t1776 XThC.Tn[5].t15 XA.XIR[15].XIC[5].icell.PDM VGND.t1775 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X556 VGND.t127 XThC.Tn[9].t19 XA.XIR[6].XIC[9].icell.PDM VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X557 VPWR.t1227 XThC.XTBN.Y.t27 XThC.Tn[7].t2 VPWR.t1226 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X558 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6].t23 XA.XIR[6].XIC[3].icell.Ien VGND.t1673 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X559 XA.XIR[1].XIC_15.icell.PDM XThR.Tn[1].t24 XA.XIR[1].XIC_15.icell.Ien VGND.t1986 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X560 VPWR.t1667 XThR.Tn[10].t21 XA.XIR[11].XIC[11].icell.PUM VPWR.t1666 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X561 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t301 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t302 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X562 VPWR.t460 XThR.XTB2.Y XThR.Tn[9].t2 VPWR.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X563 VPWR.t1127 VGND.t2691 Vbias.t4 VPWR.t570 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X564 XThC.Tn[6].t6 XThC.XTBN.Y.t28 a_6243_9615# VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X565 XA.XIR[3].XIC[5].icell.PUM XThC.Tn[5].t16 XA.XIR[3].XIC[5].icell.Ien VPWR.t1643 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X566 VGND.t73 Vbias.t50 XA.XIR[9].XIC[5].icell.SM VGND.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X567 XA.XIR[8].XIC[6].icell.Ien XThR.Tn[8].t27 VPWR.t952 VPWR.t951 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X568 VGND.t2554 XThC.Tn[6].t20 XA.XIR[1].XIC[6].icell.PDM VGND.t2553 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X569 VPWR.t391 XThR.Tn[3].t25 XA.XIR[4].XIC[4].icell.PUM VPWR.t390 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X570 VPWR.t935 XThR.Tn[7].t17 XA.XIR[8].XIC[1].icell.PUM VPWR.t934 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X571 XA.XIR[0].XIC[2].icell.PDM XThR.Tn[0].t22 XA.XIR[0].XIC[2].icell.Ien VGND.t1159 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X572 XA.XIR[11].XIC[7].icell.Ien XThR.Tn[11].t22 VPWR.t1353 VPWR.t1352 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X573 VGND.t2260 Vbias.t51 XA.XIR[3].XIC[9].icell.SM VGND.t2259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X574 VGND.t651 XThC.Tn[7].t13 XA.XIR[4].XIC[7].icell.PDM VGND.t650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X575 XA.XIR[15].XIC_15.icell.Ien VPWR.t298 VPWR.t300 VPWR.t299 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X576 VPWR.t1669 XThR.Tn[10].t22 XA.XIR[11].XIC[2].icell.PUM VPWR.t1668 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X577 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout VGND.t1340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X578 VPWR.t918 XThR.Tn[5].t23 XA.XIR[6].XIC[14].icell.PUM VPWR.t917 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X579 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t11 VPWR.t1759 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X580 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8].t28 XA.XIR[8].XIC[9].icell.Ien VGND.t729 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X581 XThC.Tn[0].t5 XThC.XTBN.Y.t29 VGND.t1205 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X582 VGND.t2262 Vbias.t52 XA.XIR[4].XIC[2].icell.SM VGND.t2261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X583 VPWR.t297 VPWR.t295 XA.XIR[9].XIC_15.icell.PUM VPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X584 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[0].t23 VGND.t1161 VGND.t1160 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X585 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[0].t24 VGND.t1163 VGND.t1162 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X586 VGND.t2264 Vbias.t53 XA.XIR[7].XIC[3].icell.SM VGND.t2263 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X587 a_4067_9615# XThC.XTBN.Y.t30 XThC.Tn[2].t5 VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X588 XThR.Tn[0].t0 XThR.XTB1.Y.t5 VGND.t207 VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X589 VGND.t2374 XThR.XTBN.Y XThR.Tn[5].t6 VGND.t2360 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X590 XA.XIR[11].XIC[7].icell.SM XA.XIR[11].XIC[7].icell.Ien Iout.t169 VGND.t1339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X591 XA.XIR[5].XIC[5].icell.Ien XThR.Tn[5].t24 VPWR.t954 VPWR.t953 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X592 VGND.t2266 Vbias.t54 XA.XIR[6].XIC[4].icell.SM VGND.t2265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X593 XThR.Tn[14].t7 XThR.XTB7.Y a_n997_715# VGND.t1367 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X594 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[12].t27 VGND.t915 VGND.t914 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X595 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[7].t18 VGND.t720 VGND.t719 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X596 VGND.t2268 Vbias.t55 XA.XIR[15].XIC[10].icell.SM VGND.t2267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X597 XA.XIR[9].XIC[5].icell.Ien XThR.Tn[9].t24 VPWR.t732 VPWR.t731 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X598 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[10].t23 VGND.t708 VGND.t707 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X599 XA.XIR[10].XIC[11].icell.SM XA.XIR[10].XIC[11].icell.Ien Iout.t173 VGND.t1344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X600 VGND.t2168 VPWR.t1952 XA.XIR[11].XIC_dummy_left.icell.PDM VGND.t2167 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X601 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6].t24 XA.XIR[6].XIC[7].icell.Ien VGND.t1674 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X602 VGND.t2373 XThR.XTBN.Y XThR.Tn[4].t11 VGND.t2372 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X603 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[3].t26 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X604 XA.XIR[6].XIC[1].icell.PUM XThC.Tn[1].t19 XA.XIR[6].XIC[1].icell.Ien VPWR.t1218 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X605 VGND.t2170 VPWR.t1953 XA.XIR[14].XIC_15.icell.PDM VGND.t2169 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X606 a_8963_9569# XThC.XTB4.Y.t5 XThC.Tn[11].t8 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X607 XA.XIR[5].XIC[13].icell.PUM XThC.Tn[13].t18 XA.XIR[5].XIC[13].icell.Ien VPWR.t906 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X608 VGND.t2270 Vbias.t56 XA.XIR[12].XIC[0].icell.SM VGND.t2269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X609 XA.XIR[1].XIC[14].icell.SM XA.XIR[1].XIC[14].icell.Ien Iout.t72 VGND.t468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X610 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t293 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X611 XA.XIR[9].XIC[13].icell.PUM XThC.Tn[13].t19 XA.XIR[9].XIC[13].icell.Ien VPWR.t1854 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X612 VGND.t2272 Vbias.t57 XA.XIR[15].XIC[1].icell.SM VGND.t2271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X613 XA.XIR[0].XIC[6].icell.PDM XThR.Tn[0].t25 XA.XIR[0].XIC[6].icell.Ien VGND.t1164 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X614 VGND.t763 XThC.Tn[4].t21 XA.XIR[6].XIC[4].icell.PDM VGND.t762 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X615 VGND.t1429 XThC.Tn[0].t18 XA.XIR[15].XIC[0].icell.PDM VGND.t1428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X616 VGND.t2274 Vbias.t58 XA.XIR[10].XIC[13].icell.SM VGND.t2273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X617 XA.XIR[11].XIC[11].icell.Ien XThR.Tn[11].t23 VPWR.t1355 VPWR.t1354 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X618 VGND.t2454 XThC.Tn[12].t17 XA.XIR[10].XIC[12].icell.PDM VGND.t2453 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X619 VPWR.t393 XThR.Tn[3].t27 XA.XIR[4].XIC[0].icell.PUM VPWR.t392 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X620 VGND.t2276 Vbias.t59 XA.XIR[13].XIC[14].icell.SM VGND.t2275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X621 XA.XIR[12].XIC_15.icell.Ien XThR.Tn[12].t28 VPWR.t1074 VPWR.t1073 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X622 VGND.t1206 XThC.XTBN.Y.t31 a_8739_9569# VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X623 VGND.t2436 XThC.Tn[13].t20 XA.XIR[13].XIC[13].icell.PDM VGND.t2435 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X624 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t1954 XA.XIR[13].XIC_dummy_left.icell.Ien VGND.t2171 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X625 VPWR.t571 bias[0].t0 Vbias.t2 VPWR.t570 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X626 VGND.t2278 Vbias.t60 XA.XIR[9].XIC[0].icell.SM VGND.t2277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X627 XA.XIR[4].XIC[4].icell.Ien XThR.Tn[4].t26 VPWR.t1540 VPWR.t1539 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X628 XA.XIR[8].XIC[1].icell.Ien XThR.Tn[8].t29 VPWR.t555 VPWR.t554 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X629 VGND.t2280 Vbias.t61 XA.XIR[0].XIC_15.icell.SM VGND.t2279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X630 VGND.t312 XThC.Tn[8].t18 XA.XIR[0].XIC[8].icell.PDM VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X631 VGND.t863 XThC.Tn[14].t18 XA.XIR[0].XIC[14].icell.PDM VGND.t862 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X632 XA.XIR[11].XIC[2].icell.Ien XThR.Tn[11].t24 VPWR.t1357 VPWR.t1356 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X633 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[7].t19 VGND.t722 VGND.t721 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X634 XA.XIR[8].XIC[7].icell.SM XA.XIR[8].XIC[7].icell.Ien Iout.t138 VGND.t929 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X635 a_9827_9569# XThC.XTBN.Y.t32 VGND.t1207 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X636 VGND.t2282 Vbias.t62 XA.XIR[3].XIC[4].icell.SM VGND.t2281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X637 XA.XIR[7].XIC[8].icell.SM XA.XIR[7].XIC[8].icell.Ien Iout.t40 VGND.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X638 VPWR.t1706 XThR.Tn[1].t25 XA.XIR[2].XIC[12].icell.PUM VPWR.t1705 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X639 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8].t30 XA.XIR[8].XIC[4].icell.Ien VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X640 VPWR.t1017 XThR.Tn[0].t26 XA.XIR[1].XIC[13].icell.PUM VPWR.t1016 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X641 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t1955 XA.XIR[3].XIC_dummy_right.icell.Ien VGND.t2172 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X642 XA.XIR[10].XIC[9].icell.SM XA.XIR[10].XIC[9].icell.Ien Iout.t112 VGND.t825 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X643 VPWR.t1542 XThR.Tn[4].t27 XA.XIR[5].XIC[13].icell.PUM VPWR.t1541 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X644 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11].t25 XA.XIR[11].XIC[5].icell.Ien VGND.t1345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X645 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[3].t28 VGND.t12 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X646 VPWR.t292 VPWR.t290 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t291 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X647 XA.XIR[15].XIC[13].icell.PDM VPWR.t1956 XA.XIR[15].XIC[13].icell.Ien VGND.t2173 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X648 VGND.t2687 XThC.XTB1.Y.t5 XThC.Tn[0].t11 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[0].t27 VGND.t837 VGND.t836 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X650 XA.XIR[11].XIC[2].icell.SM XA.XIR[11].XIC[2].icell.Ien Iout.t27 VGND.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X651 XThR.XTB7.A data[5].t1 VPWR.t1402 VPWR.t1401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X652 VGND.t818 XThC.Tn[10].t18 XA.XIR[10].XIC[10].icell.PDM VGND.t817 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X653 VPWR.t1076 XThR.Tn[12].t29 XA.XIR[13].XIC[8].icell.PUM VPWR.t1075 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X654 VGND.t2080 XThC.XTBN.A XThC.XTBN.Y.t3 VGND.t2079 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X655 XA.XIR[0].XIC[9].icell.PUM XThC.Tn[9].t20 XA.XIR[0].XIC[9].icell.Ien VPWR.t1629 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X656 VPWR.t1751 XThR.XTB7.B XThR.XTB1.Y.t2 VPWR.t1750 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X657 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t6 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X658 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[2].t22 VGND.t111 VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X659 XA.XIR[4].XIC[0].icell.Ien XThR.Tn[4].t28 VPWR.t1544 VPWR.t1543 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X660 XA.XIR[14].XIC[12].icell.SM XA.XIR[14].XIC[12].icell.Ien Iout.t213 VGND.t1829 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X661 XA.XIR[14].XIC_15.icell.PDM VPWR.t1957 VGND.t2175 VGND.t2174 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X662 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t287 VPWR.t289 VPWR.t288 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X663 XA.XIR[13].XIC[5].icell.SM XA.XIR[13].XIC[5].icell.Ien Iout.t59 VGND.t356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X664 VPWR.t1708 XThR.Tn[1].t26 XA.XIR[2].XIC[10].icell.PUM VPWR.t1707 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X665 XA.XIR[5].XIC[6].icell.PUM XThC.Tn[6].t21 XA.XIR[5].XIC[6].icell.Ien VPWR.t1878 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X666 XThC.Tn[7].t1 XThC.XTBN.Y.t33 VPWR.t1229 VPWR.t1228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X667 VGND.t2293 XThR.XTB7.B a_n1335_7243# VGND.t2292 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X668 XA.XIR[9].XIC[6].icell.PUM XThC.Tn[6].t22 XA.XIR[9].XIC[6].icell.Ien VPWR.t1422 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X669 XA.XIR[8].XIC[7].icell.PUM XThC.Tn[7].t14 XA.XIR[8].XIC[7].icell.Ien VPWR.t875 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X670 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[0].t28 VGND.t839 VGND.t838 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X671 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1958 VGND.t2177 VGND.t2176 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X672 XA.XIR[12].XIC_15.icell.PUM VPWR.t285 XA.XIR[12].XIC_15.icell.Ien VPWR.t286 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X673 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[8].t31 VGND.t216 VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X674 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12].t30 XA.XIR[12].XIC[13].icell.Ien VGND.t916 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X675 VGND.t1272 XThC.Tn[3].t19 XA.XIR[0].XIC[3].icell.PDM VGND.t1271 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X676 XA.XIR[11].XIC[8].icell.PUM XThC.Tn[8].t19 XA.XIR[11].XIC[8].icell.Ien VPWR.t634 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X677 VGND.t1755 XThC.Tn[9].t21 XA.XIR[5].XIC[9].icell.PDM VGND.t1754 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X678 XA.XIR[8].XIC[2].icell.SM XA.XIR[8].XIC[2].icell.Ien Iout.t131 VGND.t908 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X679 XA.XIR[2].XIC[12].icell.Ien XThR.Tn[2].t23 VPWR.t1487 VPWR.t1486 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X680 XA.XIR[7].XIC[3].icell.SM XA.XIR[7].XIC[3].icell.Ien Iout.t170 VGND.t1341 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X681 XThC.Tn[11].t9 XThC.XTB4.Y.t6 VPWR.t1725 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X682 VGND.t1757 XThC.Tn[9].t22 XA.XIR[9].XIC[9].icell.PDM VGND.t1756 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X683 XA.XIR[10].XIC[4].icell.SM XA.XIR[10].XIC[4].icell.Ien Iout.t37 VGND.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X684 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t282 VPWR.t284 VPWR.t283 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X685 a_n997_1803# XThR.XTBN.Y VGND.t2371 VGND.t2370 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X686 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11].t26 XA.XIR[11].XIC[0].icell.Ien VGND.t1346 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X687 XThR.Tn[3].t3 XThR.XTBN.Y a_n1049_6699# VPWR.t1811 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X688 VPWR.t744 XThR.Tn[9].t25 XA.XIR[10].XIC[8].icell.PUM VPWR.t743 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X689 VGND.t2369 XThR.XTBN.Y XThR.Tn[3].t7 VGND.t2335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X690 VGND.t2027 Vbias.t63 XA.XIR[11].XIC[6].icell.SM VGND.t2026 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X691 XA.XIR[10].XIC[7].icell.Ien XThR.Tn[10].t24 VPWR.t923 VPWR.t922 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X692 VGND.t2179 VPWR.t1959 XA.XIR[7].XIC_dummy_right.icell.PDM VGND.t2178 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X693 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1960 VGND.t2181 VGND.t2180 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X694 XThC.Tn[2].t4 XThC.XTBN.Y.t34 a_4067_9615# VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X695 VPWR.t1019 XThR.Tn[0].t29 XA.XIR[1].XIC[6].icell.PUM VPWR.t1018 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X696 XA.XIR[13].XIC[8].icell.Ien XThR.Tn[13].t25 VPWR.t417 VPWR.t416 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X697 VPWR.t1546 XThR.Tn[4].t29 XA.XIR[5].XIC[6].icell.PUM VPWR.t1545 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X698 VPWR.t1078 XThR.Tn[12].t31 XA.XIR[13].XIC[3].icell.PUM VPWR.t1077 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X699 XThR.Tn[11].t9 XThR.XTB4.Y.t5 VPWR.t1864 VPWR.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X700 VPWR.t281 VPWR.t279 XA.XIR[8].XIC_15.icell.PUM VPWR.t280 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X701 VPWR.t1739 XThC.XTB2.Y a_3773_9615# VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X702 a_n1049_8581# XThR.XTB1.Y.t6 VPWR.t694 VPWR.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X703 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t277 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t278 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X704 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[2].t24 VGND.t109 VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X705 XA.XIR[8].XIC[11].icell.PUM XThC.Tn[11].t19 XA.XIR[8].XIC[11].icell.Ien VPWR.t1826 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X706 VGND.t2029 Vbias.t64 XA.XIR[0].XIC[8].icell.SM VGND.t2028 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X707 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[10].t25 VGND.t710 VGND.t709 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X708 VGND.t653 XThC.Tn[7].t15 XA.XIR[0].XIC[7].icell.PDM VGND.t652 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X709 VGND.t1046 VGND.t1044 XA.XIR[4].XIC_dummy_right.icell.SM VGND.t1045 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X710 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[5].t25 VGND.t731 VGND.t730 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X711 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[9].t26 VGND.t454 VGND.t453 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X712 XA.XIR[9].XIC[11].icell.SM XA.XIR[9].XIC[11].icell.Ien Iout.t73 VGND.t469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X713 XA.XIR[2].XIC[10].icell.Ien XThR.Tn[2].t25 VPWR.t1469 VPWR.t1468 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X714 XA.XIR[13].XIC[0].icell.SM XA.XIR[13].XIC[0].icell.Ien Iout.t0 VGND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X715 VGND.t2183 VPWR.t1961 XA.XIR[10].XIC_dummy_left.icell.PDM VGND.t2182 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X716 VPWR.t568 XThC.XTB6.A a_5949_10571# VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X717 VPWR.t1710 XThR.Tn[1].t27 XA.XIR[2].XIC[5].icell.PUM VPWR.t1709 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X718 XA.XIR[1].XIC[4].icell.PUM XThC.Tn[4].t22 XA.XIR[1].XIC[4].icell.Ien VPWR.t977 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X719 XA.XIR[5].XIC[1].icell.PUM XThC.Tn[1].t20 XA.XIR[5].XIC[1].icell.Ien VPWR.t1219 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X720 VGND.t277 XThR.XTB3.Y.t5 XThR.Tn[2].t0 VGND.t244 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X721 VPWR.t419 XThR.Tn[13].t26 XA.XIR[14].XIC[9].icell.PUM VPWR.t418 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X722 XA.XIR[9].XIC[1].icell.PUM XThC.Tn[1].t21 XA.XIR[9].XIC[1].icell.Ien VPWR.t1220 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X723 XA.XIR[8].XIC[2].icell.PUM XThC.Tn[2].t19 XA.XIR[8].XIC[2].icell.Ien VPWR.t1430 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X724 XA.XIR[3].XIC[14].icell.PUM XThC.Tn[14].t19 XA.XIR[3].XIC[14].icell.Ien VPWR.t1043 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X725 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[8].t32 VGND.t218 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X726 XA.XIR[0].XIC[6].icell.SM XA.XIR[0].XIC[6].icell.Ien Iout.t164 VGND.t1264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X727 XThC.XTBN.Y.t1 XThC.XTBN.A VPWR.t1730 VPWR.t1729 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X728 VGND.t2031 Vbias.t65 XA.XIR[5].XIC[5].icell.SM VGND.t2030 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X729 XA.XIR[11].XIC[3].icell.PUM XThC.Tn[3].t20 XA.XIR[11].XIC[3].icell.Ien VPWR.t1324 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X730 VGND.t765 XThC.Tn[4].t23 XA.XIR[5].XIC[4].icell.PDM VGND.t764 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X731 VGND.t2033 Vbias.t66 XA.XIR[11].XIC[10].icell.SM VGND.t2032 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X732 XA.XIR[10].XIC[11].icell.Ien XThR.Tn[10].t26 VPWR.t925 VPWR.t924 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X733 XThR.Tn[8].t4 XThR.XTB1.Y.t7 a_n997_3979# VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X734 XA.XIR[6].XIC_15.icell.PUM VPWR.t275 XA.XIR[6].XIC_15.icell.Ien VPWR.t276 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X735 VGND.t1190 XThC.Tn[1].t22 XA.XIR[13].XIC[1].icell.PDM VGND.t1189 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X736 VGND.t2035 Vbias.t67 XA.XIR[12].XIC[14].icell.SM VGND.t2034 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X737 VGND.t767 XThC.Tn[4].t24 XA.XIR[9].XIC[4].icell.PDM VGND.t766 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X738 VGND.t2037 Vbias.t68 XA.XIR[8].XIC[6].icell.SM VGND.t2036 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X739 XA.XIR[7].XIC[7].icell.Ien XThR.Tn[7].t20 VPWR.t937 VPWR.t936 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X740 VGND.t2185 VPWR.t1962 XA.XIR[4].XIC_dummy_right.icell.PDM VGND.t2184 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X741 VGND.t1778 XThC.Tn[5].t17 XA.XIR[8].XIC[5].icell.PDM VGND.t1777 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X742 VGND.t2438 XThC.Tn[13].t21 XA.XIR[12].XIC[13].icell.PDM VGND.t2437 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X743 VGND.t1563 XThC.XTBN.Y.t35 a_9827_9569# VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X744 XA.XIR[2].XIC[12].icell.PUM XThC.Tn[12].t18 XA.XIR[2].XIC[12].icell.Ien VPWR.t845 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X745 VPWR.t746 XThR.Tn[9].t27 XA.XIR[10].XIC[3].icell.PUM VPWR.t745 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X746 VPWR.t1211 XThC.XTB7.Y XThC.Tn[14].t7 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X747 XThR.Tn[4].t6 XThR.XTBN.Y a_n1049_6405# VPWR.t1811 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X748 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14].t23 XA.XIR[14].XIC[8].icell.Ien VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X749 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14].t24 XA.XIR[14].XIC[14].icell.Ien VGND.t174 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X750 VGND.t2039 Vbias.t69 XA.XIR[11].XIC[1].icell.SM VGND.t2038 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X751 XA.XIR[10].XIC[2].icell.Ien XThR.Tn[10].t27 VPWR.t927 VPWR.t926 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X752 VGND.t2041 Vbias.t70 XA.XIR[7].XIC[12].icell.SM VGND.t2040 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X753 VPWR.t1906 XThR.XTB4.Y.t6 a_n1049_6699# VPWR.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X754 XA.XIR[5].XIC[14].icell.Ien XThR.Tn[5].t26 VPWR.t956 VPWR.t955 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X755 VGND.t2043 Vbias.t71 XA.XIR[6].XIC[13].icell.SM VGND.t2042 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X756 VPWR.t1021 XThR.Tn[0].t30 XA.XIR[1].XIC[1].icell.PUM VPWR.t1020 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X757 XA.XIR[13].XIC[3].icell.Ien XThR.Tn[13].t27 VPWR.t1880 VPWR.t1879 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X758 XA.XIR[9].XIC[14].icell.Ien XThR.Tn[9].t28 VPWR.t748 VPWR.t747 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X759 VGND.t2045 Vbias.t72 XA.XIR[9].XIC[14].icell.SM VGND.t2044 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X760 VPWR.t1548 XThR.Tn[4].t30 XA.XIR[5].XIC[1].icell.PUM VPWR.t1547 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X761 XA.XIR[9].XIC[9].icell.SM XA.XIR[9].XIC[9].icell.Ien Iout.t247 VGND.t2536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X762 XA.XIR[8].XIC_15.icell.Ien XThR.Tn[8].t33 VPWR.t557 VPWR.t556 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X763 XA.XIR[15].XIC[1].icell.PDM VPWR.t1963 XA.XIR[15].XIC[1].icell.Ien VGND.t2186 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X764 VPWR.t395 XThR.Tn[3].t29 XA.XIR[4].XIC[13].icell.PUM VPWR.t394 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X765 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10].t28 XA.XIR[10].XIC[5].icell.Ien VGND.t711 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X766 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1964 XA.XIR[6].XIC_dummy_right.icell.Ien VGND.t2187 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X767 XA.XIR[0].XIC[4].icell.Ien XThR.Tn[0].t31 VPWR.t1023 VPWR.t1022 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X768 XA.XIR[1].XIC[0].icell.PUM XThC.Tn[0].t19 XA.XIR[1].XIC[0].icell.Ien VPWR.t1384 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X769 VGND.t2047 Vbias.t73 XA.XIR[0].XIC[3].icell.SM VGND.t2046 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X770 XA.XIR[4].XIC[7].icell.SM XA.XIR[4].XIC[7].icell.Ien Iout.t79 VGND.t562 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X771 XA.XIR[0].XIC[10].icell.SM XA.XIR[0].XIC[10].icell.Ien Iout.t25 VGND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X772 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[5].t27 VGND.t733 VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X773 XA.XIR[2].XIC[5].icell.Ien XThR.Tn[2].t26 VPWR.t1485 VPWR.t1484 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X774 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout VGND.t680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X775 VGND.t2049 Vbias.t74 XA.XIR[8].XIC[10].icell.SM VGND.t2048 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X776 VPWR.t1810 XThR.XTBN.Y XThR.Tn[8].t8 VPWR.t1809 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X777 XA.XIR[7].XIC[11].icell.Ien XThR.Tn[7].t21 VPWR.t939 VPWR.t938 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X778 XThR.Tn[10].t3 XThR.XTB3.Y.t6 a_n997_2891# VGND.t246 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X779 XA.XIR[14].XIC[9].icell.Ien XThR.Tn[14].t25 VPWR.t533 VPWR.t532 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X780 XA.XIR[2].XIC[10].icell.PUM XThC.Tn[10].t19 XA.XIR[2].XIC[10].icell.Ien VPWR.t1004 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X781 XThC.XTB3.Y.t2 XThC.XTB7.B VPWR.t1216 VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X782 XA.XIR[0].XIC[1].icell.SM XA.XIR[0].XIC[1].icell.Ien Iout.t116 VGND.t829 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X783 VGND.t2496 Vbias.t75 XA.XIR[5].XIC[0].icell.SM VGND.t2495 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X784 VGND.t1043 VGND.t1041 XA.XIR[4].XIC_dummy_left.icell.SM VGND.t1042 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X785 VGND.t2498 Vbias.t76 XA.XIR[8].XIC[1].icell.SM VGND.t2497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X786 VPWR.t567 XThC.XTB6.A XThC.XTB2.Y VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X787 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[11].t27 VGND.t1348 VGND.t1347 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X788 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[11].t28 VGND.t1350 VGND.t1349 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X789 XA.XIR[12].XIC[5].icell.SM XA.XIR[12].XIC[5].icell.Ien Iout.t229 VGND.t2099 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X790 XA.XIR[7].XIC[2].icell.Ien XThR.Tn[7].t22 VPWR.t401 VPWR.t400 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X791 VGND.t2500 Vbias.t77 XA.XIR[3].XIC[13].icell.SM VGND.t2499 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X792 VGND.t1431 XThC.Tn[0].t20 XA.XIR[8].XIC[0].icell.PDM VGND.t1430 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X793 VGND.t611 XThC.Tn[12].t19 XA.XIR[3].XIC[12].icell.PDM VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X794 XThR.XTB3.Y.t0 XThR.XTB7.A VPWR.t1534 VPWR.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X795 XA.XIR[15].XIC[6].icell.SM XA.XIR[15].XIC[6].icell.Ien Iout.t157 VGND.t1186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X796 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12].t32 XA.XIR[12].XIC[1].icell.Ien VGND.t917 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X797 VGND.t2440 XThC.Tn[13].t22 XA.XIR[6].XIC[13].icell.PDM VGND.t2439 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X798 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7].t23 XA.XIR[7].XIC[5].icell.Ien VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X799 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1965 VGND.t2189 VGND.t2188 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X800 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t6 VGND.t1366 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X801 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14].t26 XA.XIR[14].XIC[3].icell.Ien VGND.t175 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X802 XA.XIR[10].XIC[8].icell.PUM XThC.Tn[8].t20 XA.XIR[10].XIC[8].icell.Ien VPWR.t1348 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X803 XA.XIR[1].XIC[12].icell.Ien XThR.Tn[1].t28 VPWR.t1897 VPWR.t1896 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X804 VGND.t2502 Vbias.t78 XA.XIR[2].XIC[11].icell.SM VGND.t2501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X805 XA.XIR[6].XIC_15.icell.SM XA.XIR[6].XIC_15.icell.Ien Iout.t35 VGND.t228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X806 XA.XIR[0].XIC[0].icell.Ien XThR.Tn[0].t32 VPWR.t1025 VPWR.t1024 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X807 XThR.Tn[0].t9 XThR.XTBN.Y VGND.t2368 VGND.t2311 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X808 VPWR.t678 XThR.XTB5.Y a_n1049_6405# VPWR.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X809 XA.XIR[4].XIC[13].icell.Ien XThR.Tn[4].t31 VPWR.t1550 VPWR.t1549 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X810 VGND.t2504 Vbias.t79 XA.XIR[14].XIC_15.icell.SM VGND.t2503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X811 XA.XIR[9].XIC[4].icell.SM XA.XIR[9].XIC[4].icell.Ien Iout.t242 VGND.t2531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X812 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10].t29 XA.XIR[10].XIC[0].icell.Ien VGND.t712 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X813 XThC.Tn[10].t1 XThC.XTB3.Y.t4 VPWR.t582 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X814 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5].t28 XA.XIR[5].XIC[12].icell.Ien VGND.t734 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X815 VPWR.t1808 XThR.XTBN.Y XThR.Tn[10].t11 VPWR.t1807 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X816 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout VGND.t662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X817 VPWR.t1259 XThR.Tn[11].t29 XA.XIR[12].XIC[4].icell.PUM VPWR.t1258 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X818 VPWR.t1520 XThC.XTBN.Y.t36 XThC.Tn[13].t1 VPWR.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X819 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9].t29 XA.XIR[9].XIC[12].icell.Ien VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X820 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8].t34 XA.XIR[8].XIC[13].icell.Ien VGND.t219 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X821 a_3773_9615# XThC.XTB2.Y VPWR.t1738 VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X822 XThC.Tn[5].t9 XThC.XTB6.Y VGND.t1458 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X823 XA.XIR[4].XIC[2].icell.SM XA.XIR[4].XIC[2].icell.Ien Iout.t228 VGND.t2098 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X824 XThC.Tn[2].t0 XThC.XTB3.Y.t5 VGND.t248 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X825 VPWR.t397 XThR.Tn[3].t30 XA.XIR[4].XIC[6].icell.PUM VPWR.t396 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X826 VPWR.t1483 XThR.Tn[2].t27 XA.XIR[3].XIC[7].icell.PUM VPWR.t1482 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X827 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[12].t33 VGND.t919 VGND.t918 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X828 VGND.t820 XThC.Tn[10].t20 XA.XIR[3].XIC[10].icell.PDM VGND.t819 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X829 VPWR.t1590 XThR.Tn[6].t25 XA.XIR[7].XIC[7].icell.PUM VPWR.t1589 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X830 XA.XIR[15].XIC[10].icell.SM XA.XIR[15].XIC[10].icell.Ien Iout.t8 VGND.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X831 VPWR.t958 XThR.Tn[5].t29 XA.XIR[6].XIC[8].icell.PUM VPWR.t957 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X832 VGND.t2367 XThR.XTBN.Y a_n997_3755# VGND.t2356 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X833 XA.XIR[2].XIC[5].icell.PUM XThC.Tn[5].t18 XA.XIR[2].XIC[5].icell.Ien VPWR.t1644 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X834 VPWR.t436 XThC.XTB1.Y.t6 a_2979_9615# VPWR.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X835 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[9].t30 VGND.t457 VGND.t456 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X836 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1966 VGND.t2191 VGND.t2190 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X837 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14].t27 XA.XIR[14].XIC[7].icell.Ien VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X838 XA.XIR[1].XIC[10].icell.Ien XThR.Tn[1].t29 VPWR.t1899 VPWR.t1898 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X839 VGND.t2506 Vbias.t80 XA.XIR[2].XIC[9].icell.SM VGND.t2505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X840 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[12].t34 VGND.t921 VGND.t920 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X841 XA.XIR[12].XIC[0].icell.SM XA.XIR[12].XIC[0].icell.Ien Iout.t251 VGND.t2560 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X842 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[11].t30 VGND.t1221 VGND.t1220 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X843 XA.XIR[3].XIC_15.icell.SM XA.XIR[3].XIC_15.icell.Ien Iout.t62 VGND.t385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X844 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout VGND.t1504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X845 XA.XIR[7].XIC[12].icell.SM XA.XIR[7].XIC[12].icell.Ien Iout.t248 VGND.t2537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X846 XA.XIR[14].XIC[12].icell.PUM XThC.Tn[12].t20 XA.XIR[14].XIC[12].icell.Ien VPWR.t846 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X847 XA.XIR[15].XIC[1].icell.SM XA.XIR[15].XIC[1].icell.Ien Iout.t1 VGND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X848 VGND.t2415 XThC.Tn[11].t20 XA.XIR[15].XIC[11].icell.PDM VGND.t2414 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X849 XA.XIR[11].XIC_15.icell.PDM VPWR.t1967 VGND.t2193 VGND.t2192 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X850 XA.XIR[10].XIC[13].icell.SM XA.XIR[10].XIC[13].icell.Ien Iout.t143 VGND.t1080 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X851 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5].t30 XA.XIR[5].XIC[10].icell.Ien VGND.t735 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X852 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7].t24 XA.XIR[7].XIC[0].icell.Ien VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X853 XA.XIR[13].XIC[14].icell.SM XA.XIR[13].XIC[14].icell.Ien Iout.t153 VGND.t1143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X854 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9].t31 XA.XIR[9].XIC[10].icell.Ien VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X855 XA.XIR[10].XIC[3].icell.PUM XThC.Tn[3].t21 XA.XIR[10].XIC[3].icell.Ien VPWR.t1325 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X856 a_5155_9615# XThC.XTB5.Y VPWR.t501 VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X857 XA.XIR[5].XIC_15.icell.PUM VPWR.t273 XA.XIR[5].XIC_15.icell.Ien VPWR.t274 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X858 VPWR.t1261 XThR.Tn[11].t31 XA.XIR[12].XIC[0].icell.PUM VPWR.t1260 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X859 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[6].t26 VGND.t538 VGND.t537 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X860 a_n1049_7493# XThR.XTB3.Y.t7 VPWR.t985 VPWR.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X861 VGND.t1192 XThC.Tn[1].t23 XA.XIR[12].XIC[1].icell.PDM VGND.t1191 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X862 XA.XIR[9].XIC_15.icell.PUM VPWR.t271 XA.XIR[9].XIC_15.icell.Ien VPWR.t272 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X863 VGND.t1525 XThC.Tn[2].t20 XA.XIR[15].XIC[2].icell.PDM VGND.t1524 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X864 VPWR.t1481 XThR.Tn[2].t28 XA.XIR[3].XIC[11].icell.PUM VPWR.t1480 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X865 VPWR.t791 XThR.Tn[6].t27 XA.XIR[7].XIC[11].icell.PUM VPWR.t790 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X866 VGND.t2195 VPWR.t1968 XA.XIR[13].XIC_15.icell.PDM VGND.t2194 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X867 XThC.Tn[8].t7 XThC.XTB1.Y.t7 VPWR.t438 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X868 Vbias.t3 bias[2].t0 VPWR.t1042 VPWR.t1041 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X869 XA.XIR[4].XIC[6].icell.Ien XThR.Tn[4].t32 VPWR.t587 VPWR.t586 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X870 XA.XIR[3].XIC[7].icell.Ien XThR.Tn[3].t31 VPWR.t399 VPWR.t398 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X871 VGND.t353 XThR.XTB5.Y XThR.Tn[4].t3 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X872 a_5155_9615# XThC.XTBN.Y.t37 XThC.Tn[4].t7 VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X873 VGND.t2197 VPWR.t1969 XA.XIR[0].XIC_dummy_right.icell.PDM VGND.t2196 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X874 VPWR.t1515 XThR.Tn[3].t32 XA.XIR[4].XIC[1].icell.PUM VPWR.t1514 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X875 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[12].t35 VGND.t923 VGND.t922 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X876 VPWR.t1479 XThR.Tn[2].t29 XA.XIR[3].XIC[2].icell.PUM VPWR.t1478 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X877 XThR.XTB5.Y XThR.XTB5.A VGND.t2 VGND.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X878 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[11].t32 VGND.t1223 VGND.t1222 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X879 VPWR.t793 XThR.Tn[6].t28 XA.XIR[7].XIC[2].icell.PUM VPWR.t792 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X880 VPWR.t1901 XThR.Tn[1].t30 XA.XIR[2].XIC[14].icell.PUM VPWR.t1900 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X881 VPWR.t960 XThR.Tn[5].t31 XA.XIR[6].XIC[3].icell.PUM VPWR.t959 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X882 XA.XIR[14].XIC[10].icell.PUM XThC.Tn[10].t21 XA.XIR[14].XIC[10].icell.Ien VPWR.t1005 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X883 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout VGND.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X884 VPWR.t270 VPWR.t268 XA.XIR[1].XIC_15.icell.PUM VPWR.t269 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X885 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[4].t33 XA.XIR[4].XIC[9].icell.Ien VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X886 VPWR.t267 VPWR.t265 XA.XIR[5].XIC_15.icell.PUM VPWR.t266 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X887 XA.XIR[15].XIC_15.icell.PDM VPWR.t1970 XA.XIR[15].XIC_15.icell.Ien VGND.t2198 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X888 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[6].t29 VGND.t540 VGND.t539 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X889 XA.XIR[1].XIC[5].icell.Ien XThR.Tn[1].t31 VPWR.t1903 VPWR.t1902 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X890 VGND.t2508 Vbias.t81 XA.XIR[2].XIC[4].icell.SM VGND.t2507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X891 XA.XIR[6].XIC[8].icell.SM XA.XIR[6].XIC[8].icell.Ien Iout.t107 VGND.t773 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X892 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[2].t30 VGND.t579 VGND.t578 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X893 VGND.t2510 Vbias.t82 XA.XIR[15].XIC[7].icell.SM VGND.t2509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X894 VGND.t2200 VPWR.t1971 XA.XIR[3].XIC_dummy_left.icell.PDM VGND.t2199 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X895 VGND.t2512 Vbias.t83 XA.XIR[14].XIC[8].icell.SM VGND.t2511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X896 VGND.t1486 XThC.Tn[6].t23 XA.XIR[15].XIC[6].icell.PDM VGND.t1485 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X897 VPWR.t264 VPWR.t262 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t263 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X898 XThC.Tn[14].t10 XThC.XTB7.Y a_10915_9569# VGND.t1175 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X899 XThC.XTB3.Y.t1 XThC.XTB7.A a_4387_10575# VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X900 a_n997_1803# XThR.XTBN.Y VGND.t2366 VGND.t2365 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X901 XA.XIR[1].XIC[13].icell.PUM XThC.Tn[13].t23 XA.XIR[1].XIC[13].icell.Ien VPWR.t1855 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X902 XA.XIR[3].XIC[11].icell.Ien XThR.Tn[3].t33 VPWR.t1517 VPWR.t1516 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X903 XA.XIR[15].XIC[14].icell.PDM XThR.Tn[14].t28 VGND.t178 VGND.t177 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X904 a_3773_9615# XThC.XTBN.Y.t38 XThC.Tn[1].t3 VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X905 VGND.t1194 XThC.Tn[1].t24 XA.XIR[6].XIC[1].icell.PDM VGND.t1193 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X906 XA.XIR[14].XIC[6].icell.SM XA.XIR[14].XIC[6].icell.Ien Iout.t142 VGND.t938 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X907 XA.XIR[15].XIC[8].icell.PDM XThR.Tn[14].t29 VGND.t180 VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X908 VGND.t2514 Vbias.t84 XA.XIR[5].XIC[14].icell.SM VGND.t2513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X909 VGND.t2442 XThC.Tn[13].t24 XA.XIR[5].XIC[13].icell.PDM VGND.t2441 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X910 VPWR.t1415 XThC.XTB5.A XThC.XTB1.Y.t1 VPWR.t1414 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X911 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1972 XA.XIR[5].XIC_dummy_left.icell.Ien VGND.t2201 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X912 VGND.t2444 XThC.Tn[13].t25 XA.XIR[9].XIC[13].icell.PDM VGND.t2443 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X913 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t1973 XA.XIR[9].XIC_dummy_left.icell.Ien VGND.t2202 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X914 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[1].t32 VGND.t2676 VGND.t2675 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X915 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11].t33 XA.XIR[11].XIC[11].icell.Ien VGND.t1224 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X916 VGND.t2516 Vbias.t85 XA.XIR[1].XIC[11].icell.SM VGND.t2515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X917 XA.XIR[4].XIC[1].icell.Ien XThR.Tn[4].t34 VPWR.t589 VPWR.t588 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X918 VGND.t2518 Vbias.t86 XA.XIR[0].XIC[12].icell.SM VGND.t2517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X919 XA.XIR[3].XIC[2].icell.Ien XThR.Tn[3].t34 VPWR.t1519 VPWR.t1518 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X920 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12].t36 XA.XIR[12].XIC_15.icell.Ien VGND.t924 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X921 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t260 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t261 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X922 XA.XIR[2].XIC[14].icell.Ien XThR.Tn[2].t31 VPWR.t1477 VPWR.t1476 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X923 XA.XIR[3].XIC[8].icell.SM XA.XIR[3].XIC[8].icell.Ien Iout.t204 VGND.t1592 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X924 VGND.t249 XThC.XTB3.Y.t6 XThC.Tn[2].t1 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X925 XA.XIR[14].XIC[5].icell.PUM XThC.Tn[5].t19 XA.XIR[14].XIC[5].icell.Ien VPWR.t1645 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X926 a_8739_9569# XThC.XTB3.Y.t7 XThC.Tn[10].t2 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X927 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8].t35 XA.XIR[8].XIC[1].icell.Ien VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X928 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[4].t35 XA.XIR[4].XIC[4].icell.Ien VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X929 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[3].t35 XA.XIR[3].XIC[5].icell.Ien VGND.t1550 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X930 a_n1319_6405# XThR.XTB5.A VPWR.t387 VPWR.t386 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X931 VPWR.t599 XThR.Tn[14].t30 XA.XIR[15].XIC[4].icell.PUM VPWR.t598 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X932 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11].t34 XA.XIR[11].XIC[2].icell.Ien VGND.t1225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X933 XA.XIR[7].XIC[7].icell.PUM XThC.Tn[7].t16 XA.XIR[7].XIC[7].icell.Ien VPWR.t876 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X934 VPWR.t259 VPWR.t257 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t258 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X935 XA.XIR[6].XIC[3].icell.SM XA.XIR[6].XIC[3].icell.Ien Iout.t137 VGND.t928 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X936 a_2979_9615# XThC.XTB1.Y.t8 VPWR.t440 VPWR.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X937 XA.XIR[0].XIC[13].icell.Ien XThR.Tn[0].t33 VPWR.t1196 VPWR.t1195 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X938 VGND.t1619 Vbias.t87 XA.XIR[15].XIC[2].icell.SM VGND.t1618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X939 VGND.t1621 Vbias.t88 XA.XIR[14].XIC[3].icell.SM VGND.t1620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X940 XThR.Tn[12].t10 XThR.XTBN.Y VPWR.t1806 VPWR.t1805 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X941 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout VGND.t1110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X942 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t254 VPWR.t256 VPWR.t255 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X943 XA.XIR[14].XIC[10].icell.SM XA.XIR[14].XIC[10].icell.Ien Iout.t250 VGND.t2559 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X944 XThC.Tn[11].t3 XThC.XTBN.Y.t39 VPWR.t1521 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X945 VGND.t1817 data[4].t2 XThR.XTB5.A VGND.t1816 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X946 XThR.XTBN.Y XThR.XTBN.A VGND.t1248 VGND.t1247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X947 VGND.t1847 data[3].t0 XThC.XTBN.A VGND.t1846 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X948 VGND.t1623 Vbias.t89 XA.XIR[1].XIC[9].icell.SM VGND.t1622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X949 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1974 VGND.t2204 VGND.t2203 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X950 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[8].t36 VGND.t665 VGND.t664 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X951 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t7 VGND.t351 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X952 XA.XIR[15].XIC[3].icell.PDM XThR.Tn[14].t31 VGND.t282 VGND.t281 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X953 XA.XIR[14].XIC[1].icell.SM XA.XIR[14].XIC[1].icell.Ien Iout.t4 VGND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X954 XA.XIR[10].XIC_15.icell.PDM VPWR.t1975 VGND.t2206 VGND.t2205 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X955 XA.XIR[9].XIC[13].icell.SM XA.XIR[9].XIC[13].icell.Ien Iout.t26 VGND.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X956 a_n997_2667# XThR.XTBN.Y VGND.t2364 VGND.t2323 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X957 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t252 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t253 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X958 XA.XIR[12].XIC[14].icell.SM XA.XIR[12].XIC[14].icell.Ien Iout.t95 VGND.t697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X959 XA.XIR[1].XIC[6].icell.PUM XThC.Tn[6].t24 XA.XIR[1].XIC[6].icell.Ien VPWR.t1423 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X960 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[1].t33 VGND.t2678 VGND.t2677 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X961 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11].t35 XA.XIR[11].XIC[6].icell.Ien VGND.t1226 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X962 XA.XIR[7].XIC[11].icell.PUM XThC.Tn[11].t21 XA.XIR[7].XIC[11].icell.Ien VPWR.t1827 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X963 XA.XIR[4].XIC[7].icell.PUM XThC.Tn[7].t17 XA.XIR[4].XIC[7].icell.Ien VPWR.t877 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X964 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[4].t36 VGND.t261 VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X965 VPWR.t601 XThR.Tn[14].t32 XA.XIR[15].XIC[0].icell.PUM VPWR.t600 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X966 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[8].t37 VGND.t667 VGND.t666 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X967 XA.XIR[3].XIC[8].icell.PUM XThC.Tn[8].t21 XA.XIR[3].XIC[8].icell.Ien VPWR.t1349 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X968 VGND.t1759 XThC.Tn[9].t23 XA.XIR[1].XIC[9].icell.PDM VGND.t1758 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X969 XA.XIR[3].XIC[3].icell.SM XA.XIR[3].XIC[3].icell.Ien Iout.t199 VGND.t1578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X970 XThC.Tn[4].t6 XThC.XTBN.Y.t40 a_5155_9615# VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X971 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[3].t36 XA.XIR[3].XIC[0].icell.Ien VGND.t1551 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X972 VGND.t2208 VPWR.t1976 XA.XIR[12].XIC_15.icell.PDM VGND.t2207 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X973 VPWR.t1080 XThR.Tn[12].t37 XA.XIR[13].XIC[9].icell.PUM VPWR.t1079 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X974 VPWR.t1804 XThR.XTBN.Y XThR.Tn[8].t7 VPWR.t1803 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X975 VGND.t865 XThC.Tn[14].t20 XA.XIR[11].XIC[14].icell.PDM VGND.t864 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X976 VGND.t1332 XThC.Tn[8].t22 XA.XIR[11].XIC[8].icell.PDM VGND.t1331 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X977 XA.XIR[7].XIC[2].icell.PUM XThC.Tn[2].t21 XA.XIR[7].XIC[2].icell.Ien VPWR.t1431 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X978 XA.XIR[2].XIC[14].icell.PUM XThC.Tn[14].t21 XA.XIR[2].XIC[14].icell.Ien VPWR.t1044 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X979 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t249 VPWR.t251 VPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X980 a_7651_9569# XThC.XTB1.Y.t9 XThC.Tn[8].t9 VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X981 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[2].t32 XA.XIR[2].XIC[12].icell.Ien VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X982 VGND.t1625 Vbias.t90 XA.XIR[4].XIC[5].icell.SM VGND.t1624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X983 VPWR.t500 XThC.XTB5.Y XThC.Tn[12].t1 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X984 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t1977 XA.XIR[14].XIC_dummy_right.icell.Ien VGND.t2209 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X985 VPWR.t1247 XThR.Tn[11].t36 XA.XIR[12].XIC[13].icell.PUM VPWR.t1246 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X986 VPWR.t248 VPWR.t246 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t247 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X987 VGND.t1627 Vbias.t91 XA.XIR[7].XIC[6].icell.SM VGND.t1626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X988 XA.XIR[6].XIC[7].icell.Ien XThR.Tn[6].t30 VPWR.t795 VPWR.t794 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X989 XA.XIR[5].XIC[8].icell.Ien XThR.Tn[5].t32 VPWR.t962 VPWR.t961 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X990 VGND.t1780 XThC.Tn[5].t20 XA.XIR[7].XIC[5].icell.PDM VGND.t1779 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X991 VGND.t2363 XThR.XTBN.Y XThR.Tn[1].t11 VGND.t2321 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X992 XA.XIR[15].XIC[7].icell.PDM XThR.Tn[14].t33 VGND.t284 VGND.t283 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X993 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[5].t33 VGND.t737 VGND.t736 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X994 XA.XIR[9].XIC[8].icell.Ien XThR.Tn[9].t32 VPWR.t750 VPWR.t749 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X995 VPWR.t1126 VGND.t2692 XA.XIR[0].XIC[7].icell.PUM VPWR.t1125 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X996 VPWR.t245 VPWR.t243 XA.XIR[4].XIC_15.icell.PUM VPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X997 XA.XIR[0].XIC[6].icell.Ien XThR.Tn[0].t34 VPWR.t1198 VPWR.t1197 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X998 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13].t28 XA.XIR[13].XIC[14].icell.Ien VGND.t2555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X999 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13].t29 XA.XIR[13].XIC[8].icell.Ien VGND.t2556 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1000 VGND.t1629 Vbias.t92 XA.XIR[1].XIC[4].icell.SM VGND.t1628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1001 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[2].t33 VGND.t115 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1002 XThR.Tn[6].t2 XThR.XTB7.Y VGND.t1365 VGND.t1364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1003 a_9827_9569# XThC.XTBN.Y.t41 VGND.t1564 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1004 XA.XIR[4].XIC[11].icell.PUM XThC.Tn[11].t22 XA.XIR[4].XIC[11].icell.Ien VPWR.t712 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1005 XThR.Tn[9].t9 XThR.XTBN.Y VPWR.t1802 VPWR.t1784 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1006 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[8].t38 VGND.t669 VGND.t668 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1007 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[5].t34 VGND.t321 VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1008 XA.XIR[11].XIC[9].icell.PUM XThC.Tn[9].t24 XA.XIR[11].XIC[9].icell.Ien VPWR.t1630 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1009 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout VGND.t840 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1010 XA.XIR[5].XIC[11].icell.SM XA.XIR[5].XIC[11].icell.Ien Iout.t165 VGND.t1265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1011 XA.XIR[0].XIC[9].icell.PDM XThR.Tn[0].t35 XA.XIR[0].XIC[9].icell.Ien VGND.t1152 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1012 XThC.Tn[1].t2 XThC.XTBN.Y.t42 a_3773_9615# VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1013 VGND.t418 XThC.Tn[11].t23 XA.XIR[8].XIC[11].icell.PDM VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1014 XThR.Tn[0].t8 XThR.XTBN.Y VGND.t2362 VGND.t2303 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1015 XThC.Tn[13].t9 XThC.XTB6.Y a_10051_9569# VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1016 XA.XIR[1].XIC[1].icell.PUM XThC.Tn[1].t25 XA.XIR[1].XIC[1].icell.Ien VPWR.t1221 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1017 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[2].t34 XA.XIR[2].XIC[10].icell.Ien VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1018 XA.XIR[4].XIC[2].icell.PUM XThC.Tn[2].t22 XA.XIR[4].XIC[2].icell.Ien VPWR.t1432 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1019 VPWR.t1801 XThR.XTBN.Y XThR.Tn[10].t10 VPWR.t1800 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1020 VPWR.t752 XThR.Tn[9].t33 XA.XIR[10].XIC[9].icell.PUM VPWR.t751 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1021 XA.XIR[3].XIC[3].icell.PUM XThC.Tn[3].t22 XA.XIR[3].XIC[3].icell.Ien VPWR.t1326 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1022 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[4].t37 VGND.t263 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1023 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t240 VPWR.t242 VPWR.t241 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1024 XA.XIR[0].XIC[12].icell.PDM VGND.t1038 VGND.t1040 VGND.t1039 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1025 VGND.t769 XThC.Tn[4].t25 XA.XIR[1].XIC[4].icell.PDM VGND.t768 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1026 VGND.t1196 XThC.Tn[1].t26 XA.XIR[5].XIC[1].icell.PDM VGND.t1195 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1027 VGND.t1631 Vbias.t93 XA.XIR[11].XIC[7].icell.SM VGND.t1630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1028 VGND.t1633 Vbias.t94 XA.XIR[7].XIC[10].icell.SM VGND.t1632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1029 XA.XIR[6].XIC[11].icell.Ien XThR.Tn[6].t31 VPWR.t797 VPWR.t796 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1030 VPWR.t1210 XThC.XTB7.Y a_6243_9615# VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1031 XA.XIR[2].XIC[11].icell.SM XA.XIR[2].XIC[11].icell.Ien Iout.t186 VGND.t1455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1032 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1978 VGND.t2211 VGND.t2210 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1033 VGND.t1198 XThC.Tn[1].t27 XA.XIR[9].XIC[1].icell.PDM VGND.t1197 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1034 VGND.t1782 XThC.Tn[5].t21 XA.XIR[4].XIC[5].icell.PDM VGND.t1781 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1035 XA.XIR[13].XIC[9].icell.Ien XThR.Tn[13].t30 VPWR.t1882 VPWR.t1881 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1036 VGND.t1527 XThC.Tn[2].t23 XA.XIR[8].XIC[2].icell.PDM VGND.t1526 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1037 VPWR.t1124 VGND.t2693 XA.XIR[0].XIC[11].icell.PUM VPWR.t1123 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1038 VGND.t1274 XThC.Tn[3].t23 XA.XIR[11].XIC[3].icell.PDM VGND.t1273 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1039 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10].t30 XA.XIR[10].XIC[11].icell.Ien VGND.t713 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1040 VGND.t2213 VPWR.t1979 XA.XIR[6].XIC_15.icell.PDM VGND.t2212 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1041 VGND.t1565 XThC.XTBN.Y.t43 a_8963_9569# VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1042 VGND.t1635 Vbias.t95 XA.XIR[4].XIC[0].icell.SM VGND.t1634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1043 XA.XIR[15].XIC[4].icell.PUM XThC.Tn[4].t26 XA.XIR[15].XIC[4].icell.Ien VPWR.t978 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1044 VPWR.t579 XThR.XTB1.Y.t8 XThR.Tn[8].t0 VPWR.t578 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1045 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t238 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t239 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1046 VGND.t1637 Vbias.t96 XA.XIR[7].XIC[1].icell.SM VGND.t1636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1047 VGND.t1639 Vbias.t97 XA.XIR[2].XIC[13].icell.SM VGND.t1638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1048 XA.XIR[6].XIC[2].icell.Ien XThR.Tn[6].t32 VPWR.t799 VPWR.t798 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1049 XA.XIR[11].XIC[5].icell.SM XA.XIR[11].XIC[5].icell.Ien Iout.t151 VGND.t1141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1050 VGND.t1433 XThC.Tn[0].t21 XA.XIR[7].XIC[0].icell.PDM VGND.t1432 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1051 XA.XIR[1].XIC[14].icell.Ien XThR.Tn[1].t34 VPWR.t1905 VPWR.t1904 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1052 XA.XIR[5].XIC[3].icell.Ien XThR.Tn[5].t35 VPWR.t653 VPWR.t652 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1053 VGND.t613 XThC.Tn[12].t21 XA.XIR[2].XIC[12].icell.PDM VGND.t612 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1054 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[5].t36 VGND.t323 VGND.t322 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1055 XThR.XTBN.A data[7].t0 VPWR.t1869 VPWR.t975 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1056 XA.XIR[9].XIC[3].icell.Ien XThR.Tn[9].t34 VPWR.t754 VPWR.t753 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1057 XA.XIR[4].XIC_15.icell.Ien XThR.Tn[4].t38 VPWR.t591 VPWR.t590 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1058 XA.XIR[5].XIC[9].icell.SM XA.XIR[5].XIC[9].icell.Ien Iout.t206 VGND.t1594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1059 a_6243_10571# XThC.XTB7.B XThC.XTB7.Y VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1060 VPWR.t1122 VGND.t2694 XA.XIR[0].XIC[2].icell.PUM VPWR.t1121 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1061 VPWR.t458 XThR.XTB2.Y a_n1049_7787# VPWR.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1062 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10].t31 XA.XIR[10].XIC[2].icell.Ien VGND.t714 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1063 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6].t33 XA.XIR[6].XIC[5].icell.Ien VGND.t541 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1064 XA.XIR[0].XIC[1].icell.Ien XThR.Tn[0].t36 VPWR.t1200 VPWR.t1199 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1065 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13].t31 XA.XIR[13].XIC[3].icell.Ien VGND.t2557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1066 VPWR.t1249 XThR.Tn[11].t37 XA.XIR[12].XIC[6].icell.PUM VPWR.t1248 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1067 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8].t39 XA.XIR[8].XIC_15.icell.Ien VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1068 XA.XIR[0].XIC[7].icell.SM XA.XIR[0].XIC[7].icell.Ien Iout.t77 VGND.t560 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1069 XA.XIR[0].XIC[10].icell.PDM VGND.t1035 VGND.t1037 VGND.t1036 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1070 XA.XIR[0].XIC[4].icell.PDM XThR.Tn[0].t37 XA.XIR[0].XIC[4].icell.Ien VGND.t1153 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1071 VGND.t1641 Vbias.t98 XA.XIR[8].XIC[7].icell.SM VGND.t1640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1072 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t10 VPWR.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1073 XA.XIR[2].XIC[9].icell.SM XA.XIR[2].XIC[9].icell.Ien Iout.t113 VGND.t826 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1074 VGND.t1488 XThC.Tn[6].t25 XA.XIR[8].XIC[6].icell.PDM VGND.t1487 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1075 XThC.Tn[8].t6 XThC.XTB1.Y.t10 VPWR.t442 VPWR.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1076 VPWR.t1311 XThR.Tn[10].t32 XA.XIR[11].XIC[4].icell.PUM VPWR.t1310 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1077 VPWR.t237 VPWR.t235 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1078 VGND.t1034 VGND.t1032 XA.XIR[15].XIC_dummy_right.icell.SM VGND.t1033 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1079 VGND.t655 XThC.Tn[7].t18 XA.XIR[11].XIC[7].icell.PDM VGND.t654 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1080 XThR.Tn[0].t10 XThR.XTB1.Y.t9 VGND.t2577 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1081 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7].t25 XA.XIR[7].XIC[11].icell.Ien VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1082 VGND.t1280 Vbias.t99 XA.XIR[11].XIC[2].icell.SM VGND.t1279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1083 XA.XIR[15].XIC[0].icell.PUM XThC.Tn[0].t22 XA.XIR[15].XIC[0].icell.Ien VPWR.t1385 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1084 VPWR.t595 XThR.XTB3.Y.t8 XThR.Tn[10].t1 VPWR.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1085 VGND.t822 XThC.Tn[10].t22 XA.XIR[2].XIC[10].icell.PDM VGND.t821 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1086 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[7].t26 VGND.t18 VGND.t17 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1087 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[7].t27 VGND.t20 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1088 XA.XIR[8].XIC[5].icell.SM XA.XIR[8].XIC[5].icell.Ien Iout.t156 VGND.t1185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1089 VPWR.t1737 XThC.XTB2.Y a_3773_9615# VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1090 VGND.t1435 XThC.Tn[0].t23 XA.XIR[4].XIC[0].icell.PDM VGND.t1434 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1091 VGND.t2361 XThR.XTBN.Y XThR.Tn[4].t10 VGND.t2360 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1092 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t233 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1093 XA.XIR[7].XIC[6].icell.SM XA.XIR[7].XIC[6].icell.Ien Iout.t188 VGND.t1461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1094 XA.XIR[14].XIC[14].icell.PUM XThC.Tn[14].t22 XA.XIR[14].XIC[14].icell.Ien VPWR.t1045 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1095 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10].t33 XA.XIR[10].XIC[6].icell.Ien VGND.t1266 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1096 VPWR.t1522 XThC.XTBN.Y.t44 XThC.Tn[9].t3 VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1097 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t1980 XA.XIR[2].XIC_dummy_left.icell.Ien VGND.t2214 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1098 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7].t28 XA.XIR[7].XIC[2].icell.Ien VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1099 VGND.t1566 XThC.XTBN.Y.t45 XThC.Tn[5].t1 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1100 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[3].t37 VGND.t1553 VGND.t1552 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1101 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13].t32 XA.XIR[13].XIC[7].icell.Ien VGND.t2558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1102 XA.XIR[11].XIC[0].icell.SM XA.XIR[11].XIC[0].icell.Ien Iout.t120 VGND.t860 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1103 XA.XIR[6].XIC[12].icell.SM XA.XIR[6].XIC[12].icell.Ien Iout.t210 VGND.t1814 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1104 VGND.t2359 XThR.XTBN.Y a_n997_1579# VGND.t2342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1105 XA.XIR[13].XIC[12].icell.PUM XThC.Tn[12].t22 XA.XIR[13].XIC[12].icell.Ien VPWR.t847 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1106 XA.XIR[5].XIC[4].icell.SM XA.XIR[5].XIC[4].icell.Ien Iout.t130 VGND.t907 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1107 VGND.t1282 Vbias.t100 XA.XIR[14].XIC[12].icell.SM VGND.t1281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1108 VGND.t1284 Vbias.t101 XA.XIR[10].XIC_15.icell.SM VGND.t1283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1109 a_2979_9615# XThC.XTBN.Y.t46 XThC.Tn[0].t8 VPWR.t1523 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1110 VGND.t867 XThC.Tn[14].t23 XA.XIR[10].XIC[14].icell.PDM VGND.t866 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1111 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6].t34 XA.XIR[6].XIC[0].icell.Ien VGND.t542 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1112 VGND.t1334 XThC.Tn[8].t23 XA.XIR[10].XIC[8].icell.PDM VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1113 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[1].t35 XA.XIR[1].XIC[12].icell.Ien VGND.t369 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1114 VPWR.t1251 XThR.Tn[11].t38 XA.XIR[12].XIC[1].icell.PUM VPWR.t1250 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1115 XA.XIR[0].XIC[7].icell.PUM XThC.Tn[7].t19 XA.XIR[0].XIC[7].icell.Ien VPWR.t1061 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1116 XThC.Tn[12].t6 XThC.XTB5.Y a_9827_9569# VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1117 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[4].t39 XA.XIR[4].XIC[13].icell.Ien VGND.t1820 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1118 VPWR.t1313 XThR.Tn[10].t34 XA.XIR[11].XIC[0].icell.PUM VPWR.t1312 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1119 XThR.XTB6.A data[5].t2 VPWR.t597 VPWR.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1120 XA.XIR[0].XIC[2].icell.SM XA.XIR[0].XIC[2].icell.Ien Iout.t233 VGND.t2233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1121 VPWR.t232 VPWR.t230 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t231 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1122 XThR.Tn[14].t5 XThR.XTB7.Y a_n997_715# VGND.t1363 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1123 VPWR.t603 XThR.Tn[14].t34 XA.XIR[15].XIC[13].icell.PUM VPWR.t602 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1124 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t7 VPWR.t1797 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1125 XA.XIR[11].XIC[4].icell.Ien XThR.Tn[11].t39 VPWR.t1253 VPWR.t1252 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1126 VGND.t1286 Vbias.t102 XA.XIR[8].XIC[2].icell.SM VGND.t1285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1127 XA.XIR[2].XIC[4].icell.SM XA.XIR[2].XIC[4].icell.Ien Iout.t67 VGND.t447 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1128 XA.XIR[15].XIC[12].icell.Ien VPWR.t227 VPWR.t229 VPWR.t228 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1129 XA.XIR[7].XIC[10].icell.SM XA.XIR[7].XIC[10].icell.Ien Iout.t207 VGND.t1595 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1130 XA.XIR[15].XIC[7].icell.SM XA.XIR[15].XIC[7].icell.Ien Iout.t172 VGND.t1343 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1131 VPWR.t688 XThR.Tn[1].t36 XA.XIR[2].XIC[8].icell.PUM VPWR.t687 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1132 VPWR.t881 XThR.Tn[8].t40 XA.XIR[9].XIC[12].icell.PUM VPWR.t880 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1133 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7].t29 XA.XIR[7].XIC[6].icell.Ien VGND.t315 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1134 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1981 VGND.t2216 VGND.t2215 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1135 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[0].t38 VGND.t1155 VGND.t1154 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1136 XA.XIR[10].XIC[9].icell.PUM XThC.Tn[9].t25 XA.XIR[10].XIC[9].icell.Ien VPWR.t1631 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1137 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[7].t30 VGND.t317 VGND.t316 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1138 XA.XIR[8].XIC[0].icell.SM XA.XIR[8].XIC[0].icell.Ien Iout.t68 VGND.t448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1139 XA.XIR[3].XIC[12].icell.SM XA.XIR[3].XIC[12].icell.Ien Iout.t255 VGND.t2674 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1140 XA.XIR[3].XIC_15.icell.PDM VPWR.t1982 VGND.t2218 VGND.t2217 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1141 XA.XIR[13].XIC[10].icell.PUM XThC.Tn[10].t23 XA.XIR[13].XIC[10].icell.Ien VPWR.t1006 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1142 XA.XIR[7].XIC[1].icell.SM XA.XIR[7].XIC[1].icell.Ien Iout.t175 VGND.t1371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1143 a_6243_9615# XThC.XTB7.Y VPWR.t1209 VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1144 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t225 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t226 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1145 VGND.t1031 VGND.t1029 XA.XIR[15].XIC_dummy_left.icell.SM VGND.t1030 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1146 XThC.Tn[10].t9 XThC.XTBN.Y.t47 VPWR.t1524 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1147 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[1].t37 XA.XIR[1].XIC[10].icell.Ien VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1148 XA.XIR[0].XIC[11].icell.PUM XThC.Tn[11].t24 XA.XIR[0].XIC[11].icell.Ien VPWR.t713 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1149 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[3].t38 VGND.t1555 VGND.t1554 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1150 VGND.t615 XThC.Tn[12].t23 XA.XIR[14].XIC[12].icell.PDM VGND.t614 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1151 XA.XIR[1].XIC_15.icell.PUM VPWR.t223 XA.XIR[1].XIC_15.icell.Ien VPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1152 XThC.Tn[10].t3 XThC.XTB3.Y.t8 a_8739_9569# VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1153 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[1].t38 VGND.t372 VGND.t371 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1154 VGND.t1174 XThC.XTB7.Y XThC.Tn[6].t11 VGND.t1173 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1155 XA.XIR[1].XIC[11].icell.SM XA.XIR[1].XIC[11].icell.Ien Iout.t171 VGND.t1342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1156 VGND.t2220 VPWR.t1983 XA.XIR[2].XIC_dummy_left.icell.PDM VGND.t2219 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1157 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1984 VGND.t2222 VGND.t2221 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1158 XThR.Tn[11].t6 XThR.XTBN.Y VPWR.t1798 VPWR.t1779 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1159 VGND.t1276 XThC.Tn[3].t24 XA.XIR[10].XIC[3].icell.PDM VGND.t1275 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1160 VPWR.t1525 XThC.XTBN.Y.t48 XThC.Tn[12].t11 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1161 VGND.t2224 VPWR.t1985 XA.XIR[5].XIC_15.icell.PDM VGND.t2223 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1162 XA.XIR[15].XIC[10].icell.Ien VPWR.t220 VPWR.t222 VPWR.t221 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1163 VGND.t1288 Vbias.t103 XA.XIR[13].XIC[11].icell.SM VGND.t1287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1164 XA.XIR[12].XIC[12].icell.Ien XThR.Tn[12].t38 VPWR.t1082 VPWR.t1081 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1165 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11].t40 VPWR.t1255 VPWR.t1254 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1166 VGND.t2226 VPWR.t1986 XA.XIR[9].XIC_15.icell.PDM VGND.t2225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1167 VPWR.t655 XThR.Tn[5].t37 XA.XIR[6].XIC[9].icell.PUM VPWR.t654 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1168 XA.XIR[0].XIC[2].icell.PUM XThC.Tn[2].t24 XA.XIR[0].XIC[2].icell.Ien VPWR.t1433 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1169 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t217 VPWR.t219 VPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1170 VPWR.t883 XThR.Tn[8].t41 XA.XIR[9].XIC[10].icell.PUM VPWR.t882 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1171 VGND.t1290 Vbias.t104 XA.XIR[1].XIC[13].icell.SM VGND.t1289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1172 VGND.t1292 Vbias.t105 XA.XIR[0].XIC[6].icell.SM VGND.t1291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1173 VGND.t1784 XThC.Tn[5].t22 XA.XIR[0].XIC[5].icell.PDM VGND.t1783 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1174 VGND.t1294 Vbias.t106 XA.XIR[4].XIC[14].icell.SM VGND.t1293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1175 VGND.t255 XThC.XTB7.A XThC.XTB7.Y VGND.t254 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1176 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[7].t31 VGND.t319 VGND.t318 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1177 XA.XIR[2].XIC[8].icell.Ien XThR.Tn[2].t35 VPWR.t1475 VPWR.t1474 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1178 VPWR.t690 XThR.Tn[1].t39 XA.XIR[2].XIC[3].icell.PUM VPWR.t689 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1179 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t6 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1180 XA.XIR[15].XIC[2].icell.SM XA.XIR[15].XIC[2].icell.Ien Iout.t221 VGND.t1987 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1181 a_n997_2667# XThR.XTBN.Y VGND.t2358 VGND.t2313 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1182 VPWR.t605 XThR.Tn[14].t35 XA.XIR[15].XIC[6].icell.PUM VPWR.t604 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1183 VPWR.t1497 XThR.Tn[13].t33 XA.XIR[14].XIC[7].icell.PUM VPWR.t1496 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1184 a_7875_9569# XThC.XTBN.Y.t49 VGND.t1567 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1185 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[0].t39 VGND.t1157 VGND.t1156 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1186 VGND.t824 XThC.Tn[10].t24 XA.XIR[14].XIC[10].icell.PDM VGND.t823 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1187 VGND.t2357 XThR.XTBN.Y a_n997_3979# VGND.t2356 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1188 XA.XIR[0].XIC_15.icell.Ien XThR.Tn[0].t40 VPWR.t430 VPWR.t429 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1189 XA.XIR[1].XIC[9].icell.SM XA.XIR[1].XIC[9].icell.Ien Iout.t97 VGND.t715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1190 XA.XIR[13].XIC[5].icell.PUM XThC.Tn[5].t23 XA.XIR[13].XIC[5].icell.Ien VPWR.t1646 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1191 XThC.Tn[14].t2 XThC.XTBN.Y.t50 VPWR.t1526 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1192 a_n1049_6699# XThR.XTB4.Y.t7 VPWR.t1907 VPWR.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1193 a_4861_9615# XThC.XTBN.Y.t51 XThC.Tn[3].t7 VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1194 VGND.t1296 Vbias.t107 XA.XIR[10].XIC[8].icell.SM VGND.t1295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1195 VGND.t890 XThC.Tn[7].t20 XA.XIR[10].XIC[7].icell.PDM VGND.t889 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1196 VGND.t1298 Vbias.t108 XA.XIR[13].XIC[9].icell.SM VGND.t1297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1197 XA.XIR[12].XIC[10].icell.Ien XThR.Tn[12].t39 VPWR.t1084 VPWR.t1083 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1198 XThC.Tn[2].t10 XThC.XTB3.Y.t9 VGND.t884 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1199 XThC.Tn[9].t2 XThC.XTBN.Y.t52 VPWR.t1416 VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1200 XThC.Tn[5].t0 XThC.XTBN.Y.t53 VGND.t1463 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1201 a_n1335_8107# XThR.XTB6.A XThR.XTB2.Y VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1202 VGND.t1300 Vbias.t109 XA.XIR[0].XIC[10].icell.SM VGND.t1299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1203 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[13].t34 VGND.t1534 VGND.t1533 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1204 VGND.t2446 XThC.Tn[13].t26 XA.XIR[1].XIC[13].icell.PDM VGND.t2445 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1205 XA.XIR[15].XIC[5].icell.Ien VPWR.t214 VPWR.t216 VPWR.t215 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1206 VGND.t1028 VGND.t1026 XA.XIR[11].XIC_dummy_right.icell.SM VGND.t1027 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1207 VPWR.t444 XThC.XTB1.Y.t11 a_2979_9615# VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1208 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1987 XA.XIR[1].XIC_dummy_left.icell.Ien VGND.t2227 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1209 XThC.Tn[0].t7 XThC.XTBN.Y.t54 a_2979_9615# VPWR.t1417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1210 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[3].t39 XA.XIR[3].XIC[11].icell.Ien VGND.t1556 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1211 VPWR.t885 XThR.Tn[8].t42 XA.XIR[9].XIC[5].icell.PUM VPWR.t884 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1212 VPWR.t1499 XThR.Tn[13].t35 XA.XIR[14].XIC[11].icell.PUM VPWR.t1498 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1213 XThR.Tn[12].t1 XThR.XTB5.Y VPWR.t676 VPWR.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1214 XA.XIR[8].XIC[4].icell.PUM XThC.Tn[4].t27 XA.XIR[8].XIC[4].icell.Ien VPWR.t979 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1215 XA.XIR[12].XIC[12].icell.PUM XThC.Tn[12].t24 XA.XIR[12].XIC[12].icell.Ien VPWR.t848 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1216 VGND.t1302 Vbias.t110 XA.XIR[0].XIC[1].icell.SM VGND.t1301 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1217 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t212 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t213 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1218 XA.XIR[4].XIC[5].icell.SM XA.XIR[4].XIC[5].icell.Ien Iout.t71 VGND.t452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1219 VGND.t1437 XThC.Tn[0].t24 XA.XIR[0].XIC[0].icell.PDM VGND.t1436 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1220 XThR.Tn[6].t10 XThR.XTBN.Y VGND.t2355 VGND.t2354 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1221 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t10 VPWR.t1797 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1222 XA.XIR[15].XIC[13].icell.PUM XThC.Tn[13].t27 XA.XIR[15].XIC[13].icell.Ien VPWR.t1856 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1223 VGND.t2353 XThR.XTBN.Y a_n997_2891# VGND.t2352 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1224 VGND.t2291 XThR.XTB7.B XThR.XTB7.Y VGND.t2290 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1225 XA.XIR[2].XIC[3].icell.Ien XThR.Tn[2].t36 VPWR.t1473 VPWR.t1472 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1226 XA.XIR[11].XIC[14].icell.SM XA.XIR[11].XIC[14].icell.Ien Iout.t203 VGND.t1588 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1227 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[4].t40 XA.XIR[4].XIC[1].icell.Ien VGND.t1821 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1228 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[3].t40 XA.XIR[3].XIC[2].icell.Ien VGND.t1557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1229 XA.XIR[14].XIC[7].icell.Ien XThR.Tn[14].t36 VPWR.t607 VPWR.t606 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1230 VPWR.t609 XThR.Tn[14].t37 XA.XIR[15].XIC[1].icell.PUM VPWR.t608 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1231 VGND.t2229 VPWR.t1988 XA.XIR[11].XIC_dummy_right.icell.PDM VGND.t2228 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1232 XA.XIR[2].XIC[8].icell.PUM XThC.Tn[8].t24 XA.XIR[2].XIC[8].icell.Ien VPWR.t1350 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1233 VPWR.t1501 XThR.Tn[13].t36 XA.XIR[14].XIC[2].icell.PUM VPWR.t1500 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1234 a_n997_2667# XThR.XTB4.Y.t8 XThR.Tn[11].t10 VGND.t1848 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1235 VPWR.t211 VPWR.t209 XA.XIR[12].XIC_15.icell.PUM VPWR.t210 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1236 XA.XIR[1].XIC[4].icell.SM XA.XIR[1].XIC[4].icell.Ien Iout.t41 VGND.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1237 XA.XIR[10].XIC[4].icell.Ien XThR.Tn[10].t35 VPWR.t1315 VPWR.t1314 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1238 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t206 VPWR.t208 VPWR.t207 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1239 VGND.t1878 Vbias.t111 XA.XIR[6].XIC_15.icell.SM VGND.t1877 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1240 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout VGND.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1241 XA.XIR[14].XIC[7].icell.SM XA.XIR[14].XIC[7].icell.Ien Iout.t10 VGND.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1242 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[13].t37 VGND.t1536 VGND.t1535 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1243 VGND.t1880 Vbias.t112 XA.XIR[10].XIC[3].icell.SM VGND.t1879 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1244 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t203 VPWR.t205 VPWR.t204 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1245 VGND.t1464 XThC.XTBN.Y.t55 XThC.Tn[1].t5 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1246 a_n1049_6405# XThR.XTB5.Y VPWR.t674 VPWR.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1247 VGND.t1882 Vbias.t113 XA.XIR[13].XIC[4].icell.SM VGND.t1881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1248 XA.XIR[12].XIC[5].icell.Ien XThR.Tn[12].t40 VPWR.t1086 VPWR.t1085 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1249 VPWR.t645 XThR.Tn[7].t32 XA.XIR[8].XIC[12].icell.PUM VPWR.t644 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1250 XA.XIR[0].XIC[13].icell.PDM XThR.Tn[0].t41 XA.XIR[0].XIC[13].icell.Ien VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1251 VGND.t1025 VGND.t1023 XA.XIR[8].XIC_dummy_right.icell.SM VGND.t1024 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1252 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1989 XA.XIR[13].XIC_dummy_right.icell.Ien VGND.t2230 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1253 VGND.t2232 VPWR.t1990 XA.XIR[14].XIC_dummy_left.icell.PDM VGND.t2231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1254 VPWR.t1317 XThR.Tn[10].t36 XA.XIR[11].XIC[13].icell.PUM VPWR.t1316 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1255 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[4].t41 VGND.t1823 VGND.t1822 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1256 XA.XIR[12].XIC[10].icell.PUM XThC.Tn[10].t25 XA.XIR[12].XIC[10].icell.Ien VPWR.t1007 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1257 VPWR.t1889 XThR.XTB1.Y.t10 XThR.Tn[8].t9 VPWR.t1888 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1258 XA.XIR[8].XIC[0].icell.PUM XThC.Tn[0].t25 XA.XIR[8].XIC[0].icell.Ien VPWR.t1386 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1259 XA.XIR[5].XIC[13].icell.SM XA.XIR[5].XIC[13].icell.Ien Iout.t243 VGND.t2532 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1260 VPWR.t1796 XThR.XTBN.Y XThR.Tn[7].t2 VPWR.t1795 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1261 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t201 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t202 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1262 VGND.t2096 XThC.XTB2.Y XThC.Tn[1].t11 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1263 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t199 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1264 XA.XIR[8].XIC[14].icell.SM XA.XIR[8].XIC[14].icell.Ien Iout.t121 VGND.t861 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1265 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[3].t41 XA.XIR[3].XIC[6].icell.Ien VGND.t1558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1266 XThC.Tn[12].t10 XThC.XTBN.Y.t56 VPWR.t1418 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1267 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[1].t40 VGND.t374 VGND.t373 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1268 XA.XIR[14].XIC[11].icell.Ien XThR.Tn[14].t38 VPWR.t611 VPWR.t610 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1269 VGND.t103 XThR.XTB2.Y XThR.Tn[1].t2 VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1270 XThR.Tn[1].t6 XThR.XTBN.Y a_n1049_7787# VPWR.t1775 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1271 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[4].t42 VGND.t1825 VGND.t1824 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1272 XA.XIR[4].XIC[0].icell.SM XA.XIR[4].XIC[0].icell.Ien Iout.t43 VGND.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1273 XA.XIR[6].XIC[12].icell.PUM XThC.Tn[12].t25 XA.XIR[6].XIC[12].icell.Ien VPWR.t849 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1274 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[12].t41 VGND.t1253 VGND.t1252 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1275 VGND.t420 XThC.Tn[11].t25 XA.XIR[7].XIC[11].icell.PDM VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1276 XA.XIR[2].XIC[13].icell.SM XA.XIR[2].XIC[13].icell.Ien Iout.t76 VGND.t559 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1277 XA.XIR[7].XIC[4].icell.Ien XThR.Tn[7].t33 VPWR.t647 VPWR.t646 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1278 VGND.t1884 Vbias.t114 XA.XIR[3].XIC_15.icell.SM VGND.t1883 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1279 VGND.t1886 Vbias.t115 XA.XIR[12].XIC[11].icell.SM VGND.t1885 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1280 VGND.t1022 VGND.t1020 XA.XIR[11].XIC_dummy_left.icell.SM VGND.t1021 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1281 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10].t37 VPWR.t1319 VPWR.t1318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1282 VGND.t1336 XThC.Tn[8].t25 XA.XIR[3].XIC[8].icell.PDM VGND.t1335 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1283 VGND.t869 XThC.Tn[14].t24 XA.XIR[3].XIC[14].icell.PDM VGND.t868 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1284 XA.XIR[14].XIC[2].icell.Ien XThR.Tn[14].t39 VPWR.t613 VPWR.t612 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1285 XThR.Tn[9].t1 XThR.XTB2.Y VPWR.t456 VPWR.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1286 XThR.Tn[7].t5 XThR.XTBN.Y VGND.t2351 VGND.t2350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1287 VPWR.t984 data[1].t2 XThC.XTB6.A VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1288 XA.XIR[2].XIC[3].icell.PUM XThC.Tn[3].t25 XA.XIR[2].XIC[3].icell.Ien VPWR.t1327 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1289 VPWR.t649 XThR.Tn[7].t34 XA.XIR[8].XIC[10].icell.PUM VPWR.t648 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1290 XA.XIR[15].XIC[6].icell.PUM XThC.Tn[6].t26 XA.XIR[15].XIC[6].icell.Ien VPWR.t1424 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1291 VPWR.t198 VPWR.t196 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1292 VGND.t1465 XThC.XTBN.Y.t57 a_7875_9569# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1293 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14].t40 XA.XIR[14].XIC[5].icell.Ien VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1294 VPWR.t1794 XThR.XTBN.Y XThR.Tn[13].t10 VPWR.t1782 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1295 XA.XIR[1].XIC[8].icell.Ien XThR.Tn[1].t41 VPWR.t692 VPWR.t691 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1296 VPWR.t195 VPWR.t193 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t194 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1297 VGND.t1529 XThC.Tn[2].t25 XA.XIR[7].XIC[2].icell.PDM VGND.t1528 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1298 a_8739_10571# data[0].t1 XThC.XTB7.A VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1299 XA.XIR[14].XIC[2].icell.SM XA.XIR[14].XIC[2].icell.Ien Iout.t53 VGND.t276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1300 VGND.t1888 Vbias.t116 XA.XIR[9].XIC[11].icell.SM VGND.t1887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1301 VPWR.t1000 XThR.XTB3.Y.t9 XThR.Tn[10].t4 VPWR.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1302 XA.XIR[8].XIC[12].icell.Ien XThR.Tn[8].t43 VPWR.t1180 VPWR.t1179 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1303 VGND.t1761 XThC.Tn[9].t26 XA.XIR[15].XIC[9].icell.PDM VGND.t1760 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1304 XThC.Tn[3].t6 XThC.XTBN.Y.t58 a_4861_9615# VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1305 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5].t38 XA.XIR[5].XIC[8].icell.Ien VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1306 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5].t39 XA.XIR[5].XIC[14].icell.Ien VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1307 XA.XIR[11].XIC[13].icell.Ien XThR.Tn[11].t41 VPWR.t1257 VPWR.t1256 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1308 XThR.Tn[5].t2 XThR.XTB6.Y VGND.t936 VGND.t348 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1309 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9].t35 XA.XIR[9].XIC[14].icell.Ien VGND.t459 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1310 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9].t36 XA.XIR[9].XIC[8].icell.Ien VGND.t460 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1311 VPWR.t1749 XThR.XTB7.B XThR.XTB4.Y.t0 VPWR.t1748 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1312 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout VGND.t727 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1313 XA.XIR[3].XIC[9].icell.PUM XThC.Tn[9].t27 XA.XIR[3].XIC[9].icell.Ien VPWR.t1632 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1314 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[4].t43 VGND.t1827 VGND.t1826 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1315 XA.XIR[12].XIC[5].icell.PUM XThC.Tn[5].t24 XA.XIR[12].XIC[5].icell.Ien VPWR.t1049 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1316 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1991 VGND.t2580 VGND.t2579 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1317 XA.XIR[6].XIC[10].icell.PUM XThC.Tn[10].t26 XA.XIR[6].XIC[10].icell.Ien VPWR.t1008 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1318 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout VGND.t686 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1319 VGND.t1890 Vbias.t117 XA.XIR[12].XIC[9].icell.SM VGND.t1889 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1320 VGND.t422 XThC.Tn[11].t26 XA.XIR[4].XIC[11].icell.PDM VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1321 VPWR.t1321 XThR.Tn[10].t38 XA.XIR[11].XIC[6].icell.PUM VPWR.t1320 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1322 VGND.t1019 VGND.t1017 XA.XIR[8].XIC_dummy_left.icell.SM VGND.t1018 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1323 XA.XIR[7].XIC[0].icell.Ien XThR.Tn[7].t35 VPWR.t651 VPWR.t650 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1324 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t4 VGND.t1362 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1325 VGND.t1113 XThC.Tn[1].t28 XA.XIR[1].XIC[1].icell.PDM VGND.t1112 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1326 VGND.t1892 Vbias.t118 XA.XIR[7].XIC[7].icell.SM VGND.t1891 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1327 XA.XIR[5].XIC[9].icell.Ien XThR.Tn[5].t40 VPWR.t657 VPWR.t656 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1328 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[12].t42 VGND.t1255 VGND.t1254 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1329 VGND.t1490 XThC.Tn[6].t27 XA.XIR[7].XIC[6].icell.PDM VGND.t1489 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1330 VGND.t1894 Vbias.t119 XA.XIR[6].XIC[8].icell.SM VGND.t1893 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1331 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[11].t42 VGND.t1219 VGND.t1218 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1332 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t1992 VGND.t2582 VGND.t2581 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1333 VGND.t1786 XThC.Tn[2].t26 XA.XIR[4].XIC[2].icell.PDM VGND.t1785 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1334 XA.XIR[9].XIC[9].icell.Ien XThR.Tn[9].t37 VPWR.t756 VPWR.t755 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1335 VGND.t1278 XThC.Tn[3].t26 XA.XIR[3].XIC[3].icell.PDM VGND.t1277 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1336 XA.XIR[14].XIC[8].icell.PUM XThC.Tn[8].t26 XA.XIR[14].XIC[8].icell.Ien VPWR.t1351 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1337 VGND.t1896 Vbias.t120 XA.XIR[9].XIC[9].icell.SM VGND.t1895 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1338 XA.XIR[8].XIC[10].icell.Ien XThR.Tn[8].t44 VPWR.t1182 VPWR.t1181 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1339 XA.XIR[10].XIC_15.icell.SM XA.XIR[10].XIC_15.icell.Ien Iout.t249 VGND.t2538 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1340 VPWR.t887 XThR.Tn[7].t36 XA.XIR[8].XIC[5].icell.PUM VPWR.t886 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1341 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6].t35 XA.XIR[6].XIC[11].icell.Ien VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1342 XA.XIR[15].XIC[1].icell.PUM XThC.Tn[1].t29 XA.XIR[15].XIC[1].icell.Ien VPWR.t1165 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1343 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14].t41 XA.XIR[14].XIC[0].icell.Ien VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1344 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[6].t36 VGND.t545 VGND.t544 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1345 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[6].t37 VGND.t547 VGND.t546 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1346 XA.XIR[1].XIC[3].icell.Ien XThR.Tn[1].t42 VPWR.t1027 VPWR.t1026 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1347 XA.XIR[6].XIC[6].icell.SM XA.XIR[6].XIC[6].icell.Ien Iout.t11 VGND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1348 XA.XIR[13].XIC[14].icell.PUM XThC.Tn[14].t25 XA.XIR[13].XIC[14].icell.Ien VPWR.t1046 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1349 VGND.t1898 Vbias.t121 XA.XIR[15].XIC[5].icell.SM VGND.t1897 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1350 VGND.t1900 Vbias.t122 XA.XIR[14].XIC[6].icell.SM VGND.t1899 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1351 VGND.t2520 XThC.Tn[4].t28 XA.XIR[15].XIC[4].icell.PDM VGND.t2519 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1352 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6].t38 XA.XIR[6].XIC[2].icell.Ien VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1353 VGND.t2584 VPWR.t1993 XA.XIR[10].XIC_dummy_right.icell.PDM VGND.t2583 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1354 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5].t41 XA.XIR[5].XIC[3].icell.Ien VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1355 XThC.Tn[1].t4 XThC.XTBN.Y.t59 VGND.t1466 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1356 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9].t38 XA.XIR[9].XIC[3].icell.Ien VGND.t461 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1357 XA.XIR[4].XIC_15.icell.PDM XThR.Tn[4].t44 XA.XIR[4].XIC_15.icell.Ien VGND.t1828 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1358 VPWR.t192 VPWR.t190 XA.XIR[15].XIC_15.icell.PUM VPWR.t191 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1359 XA.XIR[6].XIC[5].icell.PUM XThC.Tn[5].t25 XA.XIR[6].XIC[5].icell.Ien VPWR.t1050 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1360 XA.XIR[0].XIC[1].icell.PDM XThR.Tn[0].t42 XA.XIR[0].XIC[1].icell.Ien VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1361 XA.XIR[11].XIC[6].icell.Ien XThR.Tn[11].t43 VPWR.t1839 VPWR.t1838 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1362 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t9 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1363 VPWR.t1471 XThR.Tn[2].t37 XA.XIR[3].XIC[4].icell.PUM VPWR.t1470 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1364 VGND.t1854 Vbias.t123 XA.XIR[3].XIC[8].icell.SM VGND.t1853 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1365 VGND.t1492 XThC.Tn[6].t28 XA.XIR[4].XIC[6].icell.PDM VGND.t1491 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1366 XA.XIR[15].XIC[14].icell.Ien VPWR.t187 VPWR.t189 VPWR.t188 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1367 VGND.t1856 Vbias.t124 XA.XIR[12].XIC[4].icell.SM VGND.t1855 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1368 VPWR.t1323 XThR.Tn[10].t39 XA.XIR[11].XIC[1].icell.PUM VPWR.t1322 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1369 VGND.t892 XThC.Tn[7].t21 XA.XIR[3].XIC[7].icell.PDM VGND.t891 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1370 VPWR.t801 XThR.Tn[6].t39 XA.XIR[7].XIC[4].icell.PUM VPWR.t800 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1371 VPWR.t183 VPWR.t181 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t182 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1372 XThR.Tn[13].t5 XThR.XTB6.Y a_n997_1579# VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1373 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t4 VPWR.t1793 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1374 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout VGND.t1850 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1375 VPWR.t1184 XThR.Tn[8].t45 XA.XIR[9].XIC[14].icell.PUM VPWR.t1183 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1376 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11].t44 XA.XIR[11].XIC[9].icell.Ien VGND.t2423 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1377 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[3].t42 VGND.t1560 VGND.t1559 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1378 VGND.t1858 Vbias.t125 XA.XIR[7].XIC[2].icell.SM VGND.t1857 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1379 VGND.t1860 Vbias.t126 XA.XIR[6].XIC[3].icell.SM VGND.t1859 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1380 XA.XIR[6].XIC[10].icell.SM XA.XIR[6].XIC[10].icell.Ien Iout.t185 VGND.t1452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1381 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[11].t45 VGND.t2425 VGND.t2424 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1382 XA.XIR[3].XIC[6].icell.SM XA.XIR[3].XIC[6].icell.Ien Iout.t52 VGND.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1383 XA.XIR[14].XIC[3].icell.PUM XThC.Tn[3].t27 XA.XIR[14].XIC[3].icell.Ien VPWR.t1328 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1384 VGND.t1862 Vbias.t127 XA.XIR[9].XIC[4].icell.SM VGND.t1861 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1385 XA.XIR[8].XIC[5].icell.Ien XThR.Tn[8].t46 VPWR.t1186 VPWR.t1185 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1386 VGND.t1864 Vbias.t128 XA.XIR[14].XIC[10].icell.SM VGND.t1863 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1387 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[10].t40 VGND.t1268 VGND.t1267 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1388 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6].t40 XA.XIR[6].XIC[6].icell.Ien VGND.t549 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1389 VGND.t2076 data[2].t1 XThC.XTB7.B VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1390 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5].t42 XA.XIR[5].XIC[7].icell.Ien VGND.t327 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1391 VGND.t2349 XThR.XTBN.Y XThR.Tn[2].t6 VGND.t2348 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1392 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[3].t43 VGND.t1562 VGND.t1561 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1393 XA.XIR[13].XIC[11].icell.SM XA.XIR[13].XIC[11].icell.Ien Iout.t55 VGND.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1394 a_n1049_5317# XThR.XTB7.Y VPWR.t1366 VPWR.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1395 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9].t39 XA.XIR[9].XIC[7].icell.Ien VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1396 VGND.t1467 XThC.XTBN.Y.t60 XThC.Tn[4].t9 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1397 XA.XIR[5].XIC[12].icell.PUM XThC.Tn[12].t26 XA.XIR[5].XIC[12].icell.Ien VPWR.t850 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1398 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[6].t41 VGND.t551 VGND.t550 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1399 XA.XIR[2].XIC_15.icell.PDM VPWR.t1994 VGND.t2586 VGND.t2585 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1400 XA.XIR[6].XIC[1].icell.SM XA.XIR[6].XIC[1].icell.Ien Iout.t241 VGND.t2493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1401 XA.XIR[1].XIC[13].icell.SM XA.XIR[1].XIC[13].icell.Ien Iout.t181 VGND.t1418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1402 XA.XIR[9].XIC[12].icell.PUM XThC.Tn[12].t27 XA.XIR[9].XIC[12].icell.Ien VPWR.t851 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1403 VGND.t1866 Vbias.t129 XA.XIR[15].XIC[0].icell.SM VGND.t1865 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1404 XA.XIR[8].XIC[13].icell.PUM XThC.Tn[13].t28 XA.XIR[8].XIC[13].icell.Ien VPWR.t1857 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1405 VGND.t1868 Vbias.t130 XA.XIR[14].XIC[1].icell.SM VGND.t1867 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1406 VGND.t1870 Vbias.t131 XA.XIR[10].XIC[12].icell.SM VGND.t1869 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1407 XA.XIR[4].XIC[14].icell.SM XA.XIR[4].XIC[14].icell.Ien Iout.t216 VGND.t1844 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1408 XThR.Tn[3].t10 XThR.XTB4.Y.t9 VGND.t2679 VGND.t1200 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1409 VGND.t1872 Vbias.t132 XA.XIR[13].XIC[13].icell.SM VGND.t1871 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1410 VPWR.t1467 XThR.Tn[2].t38 XA.XIR[3].XIC[0].icell.PUM VPWR.t1466 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1411 VGND.t617 XThC.Tn[12].t28 XA.XIR[13].XIC[12].icell.PDM VGND.t616 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1412 XA.XIR[12].XIC[14].icell.Ien XThR.Tn[12].t43 VPWR.t1295 VPWR.t1294 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1413 VPWR.t803 XThR.Tn[6].t42 XA.XIR[7].XIC[0].icell.PUM VPWR.t802 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1414 VPWR.t1208 XThC.XTB7.Y a_6243_9615# VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1415 VPWR.t1410 XThC.XTB6.Y XThC.Tn[13].t6 VPWR.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1416 VPWR.t186 VPWR.t184 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1417 VGND.t1582 data[1].t3 XThC.XTB5.A VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1418 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[0].t43 VGND.t80 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1419 XA.XIR[3].XIC[4].icell.Ien XThR.Tn[3].t44 VPWR.t1265 VPWR.t1264 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1420 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[8].t47 VGND.t1136 VGND.t1135 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1421 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11].t46 VPWR.t1841 VPWR.t1840 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1422 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t178 VPWR.t180 VPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1423 VGND.t1874 Vbias.t133 XA.XIR[3].XIC[3].icell.SM VGND.t1873 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1424 XA.XIR[7].XIC[7].icell.SM XA.XIR[7].XIC[7].icell.Ien Iout.t99 VGND.t717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1425 XA.XIR[3].XIC[10].icell.SM XA.XIR[3].XIC[10].icell.Ien Iout.t7 VGND.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1426 XA.XIR[10].XIC[13].icell.Ien XThR.Tn[10].t41 VPWR.t1340 VPWR.t1339 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1427 VPWR.t432 XThR.Tn[0].t44 XA.XIR[1].XIC[12].icell.PUM VPWR.t431 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1428 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[10].t42 VGND.t1318 VGND.t1317 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1429 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout VGND.t467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1430 XA.XIR[10].XIC[8].icell.SM XA.XIR[10].XIC[8].icell.Ien Iout.t83 VGND.t646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1431 VGND.t1469 XThC.XTBN.Y.t61 XThC.Tn[7].t6 VGND.t1468 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1432 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[3].t45 VGND.t1236 VGND.t1235 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1433 VPWR.t1673 XThR.Tn[4].t45 XA.XIR[5].XIC[12].icell.PUM VPWR.t1672 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1434 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11].t47 XA.XIR[11].XIC[4].icell.Ien VGND.t2426 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1435 XA.XIR[13].XIC[9].icell.SM XA.XIR[13].XIC[9].icell.Ien Iout.t49 VGND.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1436 XA.XIR[15].XIC[12].icell.PDM VPWR.t1995 XA.XIR[15].XIC[12].icell.Ien VGND.t2587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1437 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[0].t45 VGND.t82 VGND.t81 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1438 XA.XIR[5].XIC[10].icell.PUM XThC.Tn[10].t27 XA.XIR[5].XIC[10].icell.Ien VPWR.t1009 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1439 XThR.Tn[12].t0 XThR.XTB5.Y VPWR.t672 VPWR.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1440 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[6].t43 VGND.t565 VGND.t564 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1441 a_10915_9569# XThC.XTBN.Y.t62 VGND.t1471 VGND.t1470 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1442 XA.XIR[3].XIC[1].icell.SM XA.XIR[3].XIC[1].icell.Ien Iout.t217 VGND.t1845 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1443 XA.XIR[9].XIC[10].icell.PUM XThC.Tn[10].t28 XA.XIR[9].XIC[10].icell.Ien VPWR.t701 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1444 XThR.Tn[6].t9 XThR.XTBN.Y VGND.t2347 VGND.t2346 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1445 VPWR.t1297 XThR.Tn[12].t44 XA.XIR[13].XIC[7].icell.PUM VPWR.t1296 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1446 XThC.Tn[3].t10 XThC.XTB4.Y.t7 VGND.t2075 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1447 XThC.Tn[9].t5 XThC.XTB2.Y VPWR.t1736 VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1448 VGND.t390 XThC.Tn[10].t29 XA.XIR[13].XIC[10].icell.PDM VGND.t389 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1449 a_n997_2667# XThR.XTB4.Y.t10 XThR.Tn[11].t11 VGND.t607 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1450 VGND.t424 XThC.Tn[11].t27 XA.XIR[0].XIC[11].icell.PDM VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1451 XA.XIR[15].XIC[5].icell.PDM XThR.Tn[14].t42 VGND.t288 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1452 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[5].t43 VGND.t329 VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1453 VGND.t1876 Vbias.t134 XA.XIR[5].XIC[11].icell.SM VGND.t1875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1454 XA.XIR[3].XIC[0].icell.Ien XThR.Tn[3].t46 VPWR.t1267 VPWR.t1266 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1455 XA.XIR[9].XIC_15.icell.SM XA.XIR[9].XIC_15.icell.Ien Iout.t234 VGND.t2234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1456 VGND.t2589 VPWR.t1996 XA.XIR[1].XIC_15.icell.PDM VGND.t2588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1457 VPWR.t1029 XThR.Tn[1].t43 XA.XIR[2].XIC[9].icell.PUM VPWR.t1028 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1458 VPWR.t434 XThR.Tn[0].t46 XA.XIR[1].XIC[10].icell.PUM VPWR.t433 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1459 XA.XIR[7].XIC[13].icell.Ien XThR.Tn[7].t37 VPWR.t889 VPWR.t888 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1460 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t175 VPWR.t177 VPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1461 VPWR.t1694 XThR.Tn[4].t46 XA.XIR[5].XIC[10].icell.PUM VPWR.t1693 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1462 XA.XIR[15].XIC[10].icell.PDM VPWR.t1997 XA.XIR[15].XIC[10].icell.Ien VGND.t2590 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1463 XA.XIR[12].XIC[14].icell.PUM XThC.Tn[14].t26 XA.XIR[12].XIC[14].icell.Ien VPWR.t1379 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1464 XA.XIR[8].XIC[6].icell.PUM XThC.Tn[6].t29 XA.XIR[8].XIC[6].icell.Ien VPWR.t1425 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1465 VGND.t2289 XThR.XTB7.B a_n1335_8331# VGND.t2288 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1466 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[0].t47 VGND.t623 VGND.t622 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1467 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12].t45 XA.XIR[12].XIC[12].icell.Ien VGND.t1256 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1468 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[8].t48 VGND.t1138 VGND.t1137 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1469 VGND.t1788 XThC.Tn[2].t27 XA.XIR[0].XIC[2].icell.PDM VGND.t1787 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1470 XA.XIR[11].XIC[7].icell.PUM XThC.Tn[7].t22 XA.XIR[11].XIC[7].icell.Ien VPWR.t1062 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1471 VPWR.t1419 XThC.XTBN.Y.t63 XThC.Tn[9].t1 VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1472 XA.XIR[15].XIC_15.icell.PUM VPWR.t173 XA.XIR[15].XIC_15.icell.Ien VPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1473 XA.XIR[7].XIC[2].icell.SM XA.XIR[7].XIC[2].icell.Ien Iout.t230 VGND.t2100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1474 a_10051_9569# XThC.XTBN.Y.t64 VGND.t1472 VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1475 VGND.t1763 XThC.Tn[9].t28 XA.XIR[8].XIC[9].icell.PDM VGND.t1762 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1476 XA.XIR[10].XIC[3].icell.SM XA.XIR[10].XIC[3].icell.Ien Iout.t46 VGND.t242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1477 VPWR.t1792 XThR.XTBN.Y XThR.Tn[7].t1 VPWR.t1791 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1478 VPWR.t1299 XThR.Tn[12].t46 XA.XIR[13].XIC[11].icell.PUM VPWR.t1298 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1479 XA.XIR[7].XIC[4].icell.PUM XThC.Tn[4].t29 XA.XIR[7].XIC[4].icell.Ien VPWR.t1865 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1480 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t171 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t172 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1481 XA.XIR[13].XIC[4].icell.SM XA.XIR[13].XIC[4].icell.Ien Iout.t101 VGND.t725 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1482 VPWR.t507 XThR.Tn[9].t40 XA.XIR[10].XIC[7].icell.PUM VPWR.t506 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1483 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[2].t39 XA.XIR[2].XIC[8].icell.Ien VGND.t582 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1484 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[2].t40 XA.XIR[2].XIC[14].icell.Ien VGND.t581 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1485 XThC.Tn[11].t10 XThC.XTB4.Y.t8 VPWR.t1726 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1486 VGND.t2345 XThR.XTBN.Y XThR.Tn[1].t10 VGND.t2301 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1487 XThR.Tn[1].t5 XThR.XTBN.Y a_n1049_7787# VPWR.t1772 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1488 a_7651_9569# XThC.XTBN.Y.t65 VGND.t1473 VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1489 XA.XIR[5].XIC[5].icell.PUM XThC.Tn[5].t26 XA.XIR[5].XIC[5].icell.Ien VPWR.t1051 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1490 VGND.t2470 Vbias.t135 XA.XIR[11].XIC[5].icell.SM VGND.t2469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1491 XA.XIR[10].XIC[6].icell.Ien XThR.Tn[10].t43 VPWR.t1342 VPWR.t1341 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1492 XA.XIR[9].XIC[5].icell.PUM XThC.Tn[5].t27 XA.XIR[9].XIC[5].icell.Ien VPWR.t1052 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1493 XA.XIR[13].XIC[7].icell.Ien XThR.Tn[13].t38 VPWR.t1503 VPWR.t1502 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1494 VGND.t2472 Vbias.t136 XA.XIR[5].XIC[9].icell.SM VGND.t2471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1495 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t1998 VGND.t2592 VGND.t2591 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1496 VPWR.t1301 XThR.Tn[12].t47 XA.XIR[13].XIC[2].icell.PUM VPWR.t1300 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1497 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout VGND.t1370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1498 VPWR.t891 XThR.Tn[7].t38 XA.XIR[8].XIC[14].icell.PUM VPWR.t890 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1499 XA.XIR[0].XIC_15.icell.PDM XThR.Tn[0].t48 XA.XIR[0].XIC_15.icell.Ien VGND.t624 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1500 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10].t44 XA.XIR[10].XIC[9].icell.Ien VGND.t1319 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1501 XThR.Tn[6].t1 XThR.XTB7.Y VGND.t1361 VGND.t1360 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1502 a_n1049_5611# XThR.XTB6.Y VPWR.t1098 VPWR.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1503 XThR.Tn[9].t0 XThR.XTB2.Y VPWR.t454 VPWR.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1504 VPWR.t170 VPWR.t168 XA.XIR[11].XIC_15.icell.PUM VPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1505 VGND.t2474 Vbias.t137 XA.XIR[0].XIC[7].icell.SM VGND.t2473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1506 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12].t48 XA.XIR[12].XIC[10].icell.Ien VGND.t1257 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1507 XThC.Tn[4].t8 XThC.XTBN.Y.t66 VGND.t1474 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1508 VGND.t1494 XThC.Tn[6].t30 XA.XIR[0].XIC[6].icell.PDM VGND.t1493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1509 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[5].t44 VGND.t297 VGND.t296 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1510 XA.XIR[15].XIC[0].icell.PDM XThR.Tn[14].t43 VGND.t290 VGND.t289 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1511 XA.XIR[11].XIC[11].icell.PUM XThC.Tn[11].t28 XA.XIR[11].XIC[11].icell.Ien VPWR.t714 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1512 VPWR.t1790 XThR.XTBN.Y XThR.Tn[13].t9 VPWR.t1768 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1513 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[9].t41 VGND.t155 VGND.t154 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1514 XA.XIR[2].XIC[9].icell.Ien XThR.Tn[2].t41 VPWR.t1465 VPWR.t1464 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1515 VGND.t1016 VGND.t1014 XA.XIR[7].XIC_dummy_right.icell.SM VGND.t1015 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1516 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[12].t49 VGND.t1259 VGND.t1258 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1517 XA.XIR[12].XIC[11].icell.SM XA.XIR[12].XIC[11].icell.Ien Iout.t16 VGND.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1518 VPWR.t853 XThR.Tn[0].t49 XA.XIR[1].XIC[5].icell.PUM VPWR.t852 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1519 VGND.t2594 VPWR.t1999 XA.XIR[13].XIC_dummy_left.icell.PDM VGND.t2593 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1520 VPWR.t1696 XThR.Tn[4].t47 XA.XIR[5].XIC[5].icell.PUM VPWR.t1695 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1521 VPWR.t509 XThR.Tn[9].t42 XA.XIR[10].XIC[11].icell.PUM VPWR.t508 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1522 XA.XIR[8].XIC[1].icell.PUM XThC.Tn[1].t30 XA.XIR[8].XIC[1].icell.Ien VPWR.t1166 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1523 XA.XIR[4].XIC[4].icell.PUM XThC.Tn[4].t30 XA.XIR[4].XIC[4].icell.Ien VPWR.t1866 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1524 VGND.t2578 XThR.XTB1.Y.t11 XThR.Tn[0].t11 VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1525 XA.XIR[0].XIC[5].icell.SM XA.XIR[0].XIC[5].icell.Ien Iout.t235 VGND.t2391 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1526 XThR.Tn[5].t5 XThR.XTBN.Y VGND.t2344 VGND.t2328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1527 XA.XIR[7].XIC[0].icell.PUM XThC.Tn[0].t26 XA.XIR[7].XIC[0].icell.Ien VPWR.t1387 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1528 XA.XIR[0].XIC[8].icell.PDM VGND.t1011 VGND.t1013 VGND.t1012 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1529 XA.XIR[0].XIC[14].icell.PDM VGND.t1008 VGND.t1010 VGND.t1009 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1530 VGND.t2287 XThR.XTB7.B XThR.XTB6.Y VGND.t2285 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 XA.XIR[11].XIC[2].icell.PUM XThC.Tn[2].t28 XA.XIR[11].XIC[2].icell.Ien VPWR.t1647 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1532 XA.XIR[6].XIC[14].icell.PUM XThC.Tn[14].t27 XA.XIR[6].XIC[14].icell.Ien VPWR.t1380 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1533 VGND.t625 XThC.XTBN.Y.t67 XThC.Tn[0].t4 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1534 VGND.t2476 Vbias.t138 XA.XIR[8].XIC[5].icell.SM VGND.t2475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1535 XA.XIR[7].XIC[6].icell.Ien XThR.Tn[7].t39 VPWR.t893 VPWR.t892 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1536 XA.XIR[13].XIC[11].icell.Ien XThR.Tn[13].t39 VPWR.t1371 VPWR.t1370 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1537 VGND.t2478 Vbias.t139 XA.XIR[12].XIC[13].icell.SM VGND.t2477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1538 VGND.t2522 XThC.Tn[4].t31 XA.XIR[8].XIC[4].icell.PDM VGND.t2521 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1539 VGND.t2596 VPWR.t2000 XA.XIR[3].XIC_dummy_right.icell.PDM VGND.t2595 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1540 VGND.t619 XThC.Tn[12].t29 XA.XIR[12].XIC[12].icell.PDM VGND.t618 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1541 VGND.t626 XThC.XTBN.Y.t68 XThC.Tn[3].t3 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1542 VGND.t2480 Vbias.t140 XA.XIR[15].XIC[14].icell.SM VGND.t2479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1543 VGND.t871 XThC.Tn[5].t28 XA.XIR[11].XIC[5].icell.PDM VGND.t870 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1544 VGND.t2448 XThC.Tn[13].t29 XA.XIR[15].XIC[13].icell.PDM VGND.t2447 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1545 VPWR.t511 XThR.Tn[9].t43 XA.XIR[10].XIC[2].icell.PUM VPWR.t510 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1546 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[2].t42 XA.XIR[2].XIC[3].icell.Ien VGND.t580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1547 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t2001 XA.XIR[15].XIC_dummy_left.icell.Ien VGND.t2597 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1548 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7].t40 XA.XIR[7].XIC[9].icell.Ien VGND.t672 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1549 XThC.Tn[7].t5 XThC.XTBN.Y.t69 VGND.t628 VGND.t627 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1550 VPWR.t862 XThC.XTBN.Y.t70 XThC.Tn[12].t9 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1551 VGND.t2482 Vbias.t141 XA.XIR[11].XIC[0].icell.SM VGND.t2481 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1552 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10].t45 VPWR.t1344 VPWR.t1343 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1553 XA.XIR[6].XIC[4].icell.Ien XThR.Tn[6].t44 VPWR.t805 VPWR.t804 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1554 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t165 VPWR.t167 VPWR.t166 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1555 VGND.t2484 Vbias.t142 XA.XIR[2].XIC_15.icell.SM VGND.t2483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1556 VGND.t2486 Vbias.t143 XA.XIR[6].XIC[12].icell.SM VGND.t2485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1557 VGND.t900 XThC.Tn[8].t27 XA.XIR[2].XIC[8].icell.PDM VGND.t899 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1558 VGND.t1423 XThC.Tn[14].t28 XA.XIR[2].XIC[14].icell.PDM VGND.t1422 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1559 VPWR.t452 XThR.XTB2.Y a_n1049_7787# VPWR.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1560 XA.XIR[13].XIC[2].icell.Ien XThR.Tn[13].t40 VPWR.t1373 VPWR.t1372 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1561 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[9].t44 VGND.t157 VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1562 VGND.t2488 Vbias.t144 XA.XIR[5].XIC[4].icell.SM VGND.t2487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1563 VGND.t2490 Vbias.t145 XA.XIR[9].XIC[13].icell.SM VGND.t2489 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1564 XA.XIR[9].XIC[8].icell.SM XA.XIR[9].XIC[8].icell.Ien Iout.t28 VGND.t205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1565 XA.XIR[8].XIC[14].icell.Ien XThR.Tn[8].t49 VPWR.t1188 VPWR.t1187 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1566 VGND.t630 XThC.XTBN.Y.t71 a_10915_9569# VGND.t629 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1567 VPWR.t1120 VGND.t2695 XA.XIR[0].XIC[4].icell.PUM VPWR.t1119 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1568 VPWR.t1269 XThR.Tn[3].t47 XA.XIR[4].XIC[12].icell.PUM VPWR.t1268 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1569 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10].t46 XA.XIR[10].XIC[4].icell.Ien VGND.t1320 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1570 VPWR.t1463 XThR.Tn[2].t43 XA.XIR[3].XIC[13].icell.PUM VPWR.t1462 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1571 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t2002 XA.XIR[5].XIC_dummy_right.icell.Ien VGND.t2598 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1572 XA.XIR[12].XIC[9].icell.SM XA.XIR[12].XIC[9].icell.Ien Iout.t166 VGND.t1269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1573 XA.XIR[11].XIC_15.icell.Ien XThR.Tn[11].t48 VPWR.t1843 VPWR.t1842 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1574 XThC.Tn[11].t11 XThC.XTB4.Y.t9 a_8963_9569# VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1575 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13].t41 XA.XIR[13].XIC[5].icell.Ien VGND.t1375 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1576 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t2003 XA.XIR[9].XIC_dummy_right.icell.Ien VGND.t2599 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1577 VPWR.t807 XThR.Tn[6].t45 XA.XIR[7].XIC[13].icell.PUM VPWR.t806 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1578 VGND.t1597 XThC.XTB4.Y.t10 XThC.Tn[3].t9 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1579 VGND.t2492 Vbias.t146 XA.XIR[0].XIC[2].icell.SM VGND.t2491 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1580 XThR.Tn[14].t11 XThR.XTBN.Y VPWR.t1789 VPWR.t1770 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1581 XA.XIR[4].XIC[0].icell.PUM XThC.Tn[0].t27 XA.XIR[4].XIC[0].icell.Ien VPWR.t1388 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1582 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t163 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t164 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1583 a_7875_9569# XThC.XTBN.Y.t72 VGND.t631 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1584 VPWR.t1096 XThR.XTB6.Y XThR.Tn[13].t3 VPWR.t1095 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1585 VGND.t392 XThC.Tn[10].t30 XA.XIR[12].XIC[10].icell.PDM VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1586 XA.XIR[2].XIC[9].icell.PUM XThC.Tn[9].t29 XA.XIR[2].XIC[9].icell.Ien VPWR.t1633 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1587 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[2].t44 XA.XIR[2].XIC[7].icell.Ien VGND.t583 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1588 XA.XIR[0].XIC[0].icell.SM XA.XIR[0].XIC[0].icell.Ien Iout.t163 VGND.t1251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1589 XA.XIR[0].XIC[3].icell.PDM VGND.t1005 VGND.t1007 VGND.t1006 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1590 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t2004 XA.XIR[12].XIC_dummy_left.icell.Ien VGND.t2600 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1591 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14].t44 XA.XIR[14].XIC[11].icell.Ien VGND.t291 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1592 XThC.Tn[11].t5 XThC.XTB4.Y.t11 a_8963_9569# VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1593 VGND.t1954 Vbias.t147 XA.XIR[8].XIC[0].icell.SM VGND.t1953 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1594 XA.XIR[7].XIC[1].icell.Ien XThR.Tn[7].t41 VPWR.t895 VPWR.t894 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1595 VGND.t1956 Vbias.t148 XA.XIR[3].XIC[12].icell.SM VGND.t1955 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1596 XA.XIR[6].XIC[0].icell.Ien XThR.Tn[6].t46 VPWR.t809 VPWR.t808 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1597 VGND.t1004 VGND.t1002 XA.XIR[7].XIC_dummy_left.icell.SM VGND.t1003 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1598 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t161 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t162 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1599 XThC.Tn[0].t0 XThC.XTB1.Y.t12 VGND.t89 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1600 XA.XIR[15].XIC[5].icell.SM XA.XIR[15].XIC[5].icell.Ien Iout.t36 VGND.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1601 VGND.t633 XThC.XTBN.Y.t73 a_10051_9569# VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1602 VGND.t1439 XThC.Tn[0].t28 XA.XIR[11].XIC[0].icell.PDM VGND.t1438 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1603 VPWR.t1271 XThR.Tn[3].t48 XA.XIR[4].XIC[10].icell.PUM VPWR.t1270 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1604 VGND.t621 XThC.Tn[12].t30 XA.XIR[6].XIC[12].icell.PDM VGND.t620 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1605 XThR.XTB1.Y.t0 XThR.XTB5.A VPWR.t385 VPWR.t384 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1606 VPWR.t1118 VGND.t2696 XA.XIR[0].XIC[0].icell.PUM VPWR.t1117 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1607 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7].t42 XA.XIR[7].XIC[4].icell.Ien VGND.t673 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1608 XThR.Tn[13].t4 XThR.XTB6.Y a_n997_1579# VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1609 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14].t45 XA.XIR[14].XIC[2].icell.Ien VGND.t292 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1610 XA.XIR[10].XIC[7].icell.PUM XThC.Tn[7].t23 XA.XIR[10].XIC[7].icell.Ien VPWR.t1063 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1611 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2005 VGND.t2602 VGND.t2601 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1612 VGND.t1103 XThC.Tn[3].t28 XA.XIR[2].XIC[3].icell.PDM VGND.t1102 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1613 XA.XIR[13].XIC[8].icell.PUM XThC.Tn[8].t28 XA.XIR[13].XIC[8].icell.Ien VPWR.t1064 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1614 VGND.t634 XThC.XTBN.Y.t74 a_7651_9569# VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1615 XA.XIR[4].XIC[12].icell.Ien XThR.Tn[4].t48 VPWR.t1698 VPWR.t1697 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1616 XA.XIR[9].XIC[3].icell.SM XA.XIR[9].XIC[3].icell.Ien Iout.t65 VGND.t445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1617 XThC.XTBN.Y.t2 XThC.XTBN.A VGND.t2078 VGND.t2077 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1618 XA.XIR[3].XIC[13].icell.Ien XThR.Tn[3].t49 VPWR.t1273 VPWR.t1272 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1619 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t158 VPWR.t160 VPWR.t159 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1620 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[1].t44 XA.XIR[1].XIC[14].icell.Ien VGND.t844 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1621 XA.XIR[12].XIC[4].icell.SM XA.XIR[12].XIC[4].icell.Ien Iout.t105 VGND.t771 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1622 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[1].t45 XA.XIR[1].XIC[8].icell.Ien VGND.t845 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1623 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout VGND.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1624 a_n1335_7243# XThR.XTB7.A XThR.XTB3.Y.t1 VGND.t1589 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1625 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13].t42 XA.XIR[13].XIC[0].icell.Ien VGND.t1376 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1626 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8].t50 XA.XIR[8].XIC[12].icell.Ien VGND.t1837 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1627 XA.XIR[0].XIC[7].icell.PDM VGND.t999 VGND.t1001 VGND.t1000 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1628 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t6 VPWR.t1786 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1629 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11].t49 XA.XIR[11].XIC[13].icell.Ien VGND.t2427 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1630 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2006 VGND.t2604 VGND.t2603 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1631 a_4067_9615# XThC.XTB3.Y.t10 VPWR.t1057 VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1632 VPWR.t864 XThC.XTBN.Y.t75 XThC.Tn[7].t0 VPWR.t863 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1633 VPWR.t1461 XThR.Tn[2].t45 XA.XIR[3].XIC[6].icell.PUM VPWR.t1460 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1634 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[11].t50 VGND.t184 VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1635 XA.XIR[15].XIC[8].icell.Ien VPWR.t155 VPWR.t157 VPWR.t156 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1636 VPWR.t811 XThR.Tn[6].t47 XA.XIR[7].XIC[6].icell.PUM VPWR.t810 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1637 VGND.t2343 XThR.XTBN.Y a_n997_1803# VGND.t2342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1638 VPWR.t621 XThR.Tn[5].t45 XA.XIR[6].XIC[7].icell.PUM VPWR.t620 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1639 XThR.Tn[3].t6 XThR.XTBN.Y VGND.t2341 VGND.t2295 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1640 VGND.t394 XThC.Tn[10].t31 XA.XIR[6].XIC[10].icell.PDM VGND.t393 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1641 VPWR.t1683 XThR.Tn[8].t51 XA.XIR[9].XIC[8].icell.PUM VPWR.t1682 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1642 VPWR.t1537 XThC.XTB4.Y.t12 XThC.Tn[11].t6 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14].t46 XA.XIR[14].XIC[6].icell.Ien VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1644 XA.XIR[10].XIC[11].icell.PUM XThC.Tn[11].t29 XA.XIR[10].XIC[11].icell.Ien VPWR.t715 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1645 VGND.t1958 Vbias.t149 XA.XIR[2].XIC[8].icell.SM VGND.t1957 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1646 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[12].t50 VGND.t1261 VGND.t1260 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1647 XA.XIR[1].XIC[9].icell.Ien XThR.Tn[1].t46 VPWR.t1031 VPWR.t1030 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1648 VGND.t894 XThC.Tn[7].t24 XA.XIR[2].XIC[7].icell.PDM VGND.t893 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1649 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[11].t51 VGND.t186 VGND.t185 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1650 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[7].t43 VGND.t675 VGND.t674 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1651 XA.XIR[4].XIC[10].icell.Ien XThR.Tn[4].t49 VPWR.t1700 VPWR.t1699 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1652 XA.XIR[15].XIC[0].icell.SM XA.XIR[15].XIC[0].icell.Ien Iout.t57 VGND.t354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1653 VGND.t2606 VPWR.t2007 XA.XIR[12].XIC_dummy_left.icell.PDM VGND.t2605 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1654 XThC.Tn[0].t3 XThC.XTBN.Y.t76 VGND.t635 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1655 XA.XIR[10].XIC[12].icell.SM XA.XIR[10].XIC[12].icell.Ien Iout.t108 VGND.t778 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1656 VPWR.t1275 XThR.Tn[3].t50 XA.XIR[4].XIC[5].icell.PUM VPWR.t1274 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1657 XA.XIR[13].XIC[13].icell.SM XA.XIR[13].XIC[13].icell.Ien Iout.t135 VGND.t926 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1658 XThC.Tn[3].t2 XThC.XTBN.Y.t77 VGND.t636 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1659 VGND.t902 XThC.Tn[8].t29 XA.XIR[14].XIC[8].icell.PDM VGND.t901 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1660 VGND.t1425 XThC.Tn[14].t29 XA.XIR[14].XIC[14].icell.PDM VGND.t1424 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1661 XA.XIR[10].XIC[2].icell.PUM XThC.Tn[2].t29 XA.XIR[10].XIC[2].icell.Ien VPWR.t1648 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1662 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8].t52 XA.XIR[8].XIC[10].icell.Ien VGND.t1838 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1663 XA.XIR[5].XIC[14].icell.PUM XThC.Tn[14].t30 XA.XIR[5].XIC[14].icell.Ien VPWR.t1381 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1664 XA.XIR[13].XIC[3].icell.PUM XThC.Tn[3].t29 XA.XIR[13].XIC[3].icell.Ien VPWR.t1160 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1665 XA.XIR[9].XIC[14].icell.PUM XThC.Tn[14].t31 XA.XIR[9].XIC[14].icell.Ien VPWR.t1382 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1666 XA.XIR[8].XIC_15.icell.PUM VPWR.t153 XA.XIR[8].XIC_15.icell.Ien VPWR.t154 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1667 a_n1049_8581# XThR.XTB1.Y.t12 VPWR.t1891 VPWR.t1890 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1668 VGND.t1115 XThC.Tn[1].t31 XA.XIR[15].XIC[1].icell.PDM VGND.t1114 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1669 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[8].t53 VGND.t1840 VGND.t1839 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1670 VPWR.t152 VPWR.t150 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1671 VGND.t1960 Vbias.t150 XA.XIR[10].XIC[6].icell.SM VGND.t1959 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1672 VGND.t873 XThC.Tn[5].t29 XA.XIR[10].XIC[5].icell.PDM VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1673 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[1].t47 XA.XIR[1].XIC[3].icell.Ien VGND.t846 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1674 XA.XIR[12].XIC[8].icell.Ien XThR.Tn[12].t51 VPWR.t1303 VPWR.t1302 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1675 VPWR.t623 XThR.Tn[5].t46 XA.XIR[6].XIC[11].icell.PUM VPWR.t622 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1676 XA.XIR[0].XIC[4].icell.PUM XThC.Tn[4].t32 XA.XIR[0].XIC[4].icell.Ien VPWR.t1867 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1677 VGND.t1962 Vbias.t151 XA.XIR[1].XIC_15.icell.SM VGND.t1961 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1678 XA.XIR[7].XIC[13].icell.PUM XThC.Tn[13].t30 XA.XIR[7].XIC[13].icell.Ien VPWR.t1858 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1679 XThC.XTB1.Y.t2 XThC.XTB5.A a_3299_10575# VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1680 XA.XIR[3].XIC[6].icell.Ien XThR.Tn[3].t51 VPWR.t1277 VPWR.t1276 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1681 VPWR.t1459 XThR.Tn[2].t46 XA.XIR[3].XIC[1].icell.PUM VPWR.t1458 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1682 VGND.t859 XThR.XTB3.Y.t10 XThR.Tn[2].t2 VGND.t858 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1683 XA.XIR[15].XIC[3].icell.Ien VPWR.t147 VPWR.t149 VPWR.t148 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1684 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[11].t52 VGND.t188 VGND.t187 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1685 VGND.t1964 Vbias.t152 XA.XIR[11].XIC[14].icell.SM VGND.t1963 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1686 XA.XIR[10].XIC_15.icell.Ien XThR.Tn[10].t47 VPWR.t1346 VPWR.t1345 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1687 XA.XIR[14].XIC[9].icell.PUM XThC.Tn[9].t30 XA.XIR[14].XIC[9].icell.Ien VPWR.t1634 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1688 VPWR.t813 XThR.Tn[6].t48 XA.XIR[7].XIC[1].icell.PUM VPWR.t812 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1689 VPWR.t625 XThR.Tn[5].t47 XA.XIR[6].XIC[2].icell.PUM VPWR.t624 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1690 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout VGND.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1691 VPWR.t855 XThR.Tn[0].t50 XA.XIR[1].XIC[14].icell.PUM VPWR.t854 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1692 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[3].t52 XA.XIR[3].XIC[9].icell.Ien VGND.t1237 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1693 VPWR.t1702 XThR.Tn[4].t50 XA.XIR[5].XIC[14].icell.PUM VPWR.t1701 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1694 VPWR.t1685 XThR.Tn[8].t54 XA.XIR[9].XIC[3].icell.PUM VPWR.t1684 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1695 VGND.t638 XThC.XTBN.Y.t78 XThC.Tn[6].t2 VGND.t637 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1696 VGND.t1966 Vbias.t153 XA.XIR[2].XIC[3].icell.SM VGND.t1965 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1697 XA.XIR[6].XIC[7].icell.SM XA.XIR[6].XIC[7].icell.Ien Iout.t48 VGND.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1698 XThC.Tn[10].t5 XThC.XTB3.Y.t11 VPWR.t1058 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1699 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[7].t44 VGND.t677 VGND.t676 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1700 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[2].t47 VGND.t523 VGND.t522 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1701 XA.XIR[4].XIC[5].icell.Ien XThR.Tn[4].t51 VPWR.t1704 VPWR.t1703 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1702 VGND.t998 VGND.t996 XA.XIR[0].XIC_dummy_right.icell.SM VGND.t997 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1703 VGND.t1968 Vbias.t154 XA.XIR[14].XIC[7].icell.SM VGND.t1967 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1704 VGND.t1970 Vbias.t155 XA.XIR[10].XIC[10].icell.SM VGND.t1969 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1705 XThC.Tn[14].t6 XThC.XTB7.Y VPWR.t1207 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1706 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[5].t48 VGND.t299 VGND.t298 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1707 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[1].t48 XA.XIR[1].XIC[7].icell.Ien VGND.t847 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1708 VGND.t2608 VPWR.t2008 XA.XIR[6].XIC_dummy_left.icell.PDM VGND.t2607 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1709 VGND.t294 XThC.XTB1.Y.t13 XThC.Tn[0].t1 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1710 VGND.t1105 XThC.Tn[3].t30 XA.XIR[14].XIC[3].icell.PDM VGND.t1104 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1711 XA.XIR[0].XIC[0].icell.PUM XThC.Tn[0].t29 XA.XIR[0].XIC[0].icell.Ien VPWR.t1389 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1712 XA.XIR[1].XIC[12].icell.PUM XThC.Tn[12].t31 XA.XIR[1].XIC[12].icell.Ien VPWR.t963 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1713 XA.XIR[4].XIC[13].icell.PUM XThC.Tn[13].t31 XA.XIR[4].XIC[13].icell.Ien VPWR.t538 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1714 VGND.t1972 Vbias.t156 XA.XIR[10].XIC[1].icell.SM VGND.t1971 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1715 XThR.Tn[8].t6 XThR.XTBN.Y VPWR.t1788 VPWR.t1787 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1716 XA.XIR[0].XIC[14].icell.SM XA.XIR[0].XIC[14].icell.Ien Iout.t117 VGND.t841 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1717 VGND.t1974 Vbias.t157 XA.XIR[5].XIC[13].icell.SM VGND.t1973 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1718 XA.XIR[14].XIC[5].icell.SM XA.XIR[14].XIC[5].icell.Ien Iout.t193 VGND.t1531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1719 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[13].t43 VGND.t1378 VGND.t1377 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1720 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[13].t44 VGND.t1380 VGND.t1379 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1721 VGND.t2564 XThC.Tn[0].t30 XA.XIR[10].XIC[0].icell.PDM VGND.t2563 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1722 VGND.t739 XThC.Tn[12].t32 XA.XIR[5].XIC[12].icell.PDM VGND.t738 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1723 XA.XIR[12].XIC[3].icell.Ien XThR.Tn[12].t52 VPWR.t1305 VPWR.t1304 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1724 VGND.t741 XThC.Tn[12].t33 XA.XIR[9].XIC[12].icell.PDM VGND.t740 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1725 VGND.t1976 Vbias.t158 XA.XIR[8].XIC[14].icell.SM VGND.t1975 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1726 XA.XIR[7].XIC_15.icell.Ien XThR.Tn[7].t45 VPWR.t897 VPWR.t896 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1727 VGND.t192 XThC.Tn[13].t32 XA.XIR[8].XIC[13].icell.PDM VGND.t191 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1728 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t2009 XA.XIR[8].XIC_dummy_left.icell.Ien VGND.t2609 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1729 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t9 VPWR.t1786 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1730 XA.XIR[3].XIC[1].icell.Ien XThR.Tn[3].t53 VPWR.t1279 VPWR.t1278 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1731 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[4].t52 VGND.t1978 VGND.t1977 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1732 XA.XIR[12].XIC[8].icell.PUM XThC.Tn[8].t30 XA.XIR[12].XIC[8].icell.Ien VPWR.t1065 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1733 VGND.t1643 Vbias.t159 XA.XIR[4].XIC[11].icell.SM VGND.t1642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1734 XA.XIR[3].XIC[7].icell.SM XA.XIR[3].XIC[7].icell.Ien Iout.t129 VGND.t905 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1735 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[2].t48 VGND.t521 VGND.t520 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1736 XThR.XTBN.A data[7].t1 VGND.t1454 VGND.t1453 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1737 XA.XIR[6].XIC[13].icell.Ien XThR.Tn[6].t49 VPWR.t815 VPWR.t814 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1738 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[3].t54 XA.XIR[3].XIC[4].icell.Ien VGND.t1238 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1739 XThC.Tn[14].t5 XThC.XTB7.Y VPWR.t1206 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1740 VPWR.t1359 XThR.Tn[13].t45 XA.XIR[14].XIC[4].icell.PUM VPWR.t1358 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1741 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11].t53 XA.XIR[11].XIC[1].icell.Ien VGND.t189 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1742 XA.XIR[7].XIC[6].icell.PUM XThC.Tn[6].t31 XA.XIR[7].XIC[6].icell.Ien VPWR.t1426 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1743 VPWR.t1116 VGND.t2697 XA.XIR[0].XIC[13].icell.PUM VPWR.t1115 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1744 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2010 XA.XIR[2].XIC_dummy_right.icell.Ien VGND.t2610 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1745 VGND.t896 XThC.Tn[7].t25 XA.XIR[14].XIC[7].icell.PDM VGND.t895 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1746 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10].t48 XA.XIR[10].XIC[13].icell.Ien VGND.t1321 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1747 XThC.XTB2.Y XThC.XTB7.B VPWR.t1215 VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1748 XA.XIR[1].XIC[10].icell.PUM XThC.Tn[10].t32 XA.XIR[1].XIC[10].icell.Ien VPWR.t702 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1749 XA.XIR[6].XIC[2].icell.SM XA.XIR[6].XIC[2].icell.Ien Iout.t122 VGND.t882 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1750 XA.XIR[0].XIC[12].icell.Ien XThR.Tn[0].t51 VPWR.t857 VPWR.t856 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1751 XThR.Tn[5].t4 XThR.XTBN.Y VGND.t2340 VGND.t2319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1752 VGND.t1765 XThC.Tn[9].t31 XA.XIR[7].XIC[9].icell.PDM VGND.t1764 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1753 XA.XIR[15].XIC[11].icell.PDM XThR.Tn[14].t47 VGND.t509 VGND.t508 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1754 VGND.t1645 Vbias.t160 XA.XIR[14].XIC[2].icell.SM VGND.t1644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1755 VGND.t396 XThC.Tn[10].t33 XA.XIR[5].XIC[10].icell.PDM VGND.t395 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1756 XThR.Tn[10].t9 XThR.XTBN.Y VPWR.t1785 VPWR.t1784 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1757 VPWR.t899 XThR.Tn[7].t46 XA.XIR[8].XIC[8].icell.PUM VPWR.t898 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1758 VGND.t398 XThC.Tn[10].t34 XA.XIR[9].XIC[10].icell.PDM VGND.t397 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1759 a_5949_9615# XThC.XTB6.Y VPWR.t1409 VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1760 VGND.t1647 Vbias.t161 XA.XIR[1].XIC[8].icell.SM VGND.t1646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1761 VGND.t1649 Vbias.t162 XA.XIR[4].XIC[9].icell.SM VGND.t1648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1762 XA.XIR[14].XIC[0].icell.SM XA.XIR[14].XIC[0].icell.Ien Iout.t90 VGND.t663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1763 XA.XIR[15].XIC[2].icell.PDM XThR.Tn[14].t48 VGND.t511 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1764 VPWR.t1059 XThC.XTB3.Y.t12 XThC.Tn[10].t6 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1765 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[13].t46 VGND.t1352 VGND.t1351 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1766 VGND.t995 VGND.t993 XA.XIR[0].XIC_dummy_left.icell.SM VGND.t994 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1767 XA.XIR[5].XIC_15.icell.SM XA.XIR[5].XIC_15.icell.Ien Iout.t61 VGND.t359 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1768 XA.XIR[9].XIC[12].icell.SM XA.XIR[9].XIC[12].icell.Ien Iout.t74 VGND.t536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1769 XThC.Tn[13].t0 XThC.XTBN.Y.t79 VPWR.t866 VPWR.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1770 XA.XIR[13].XIC_15.icell.PDM VPWR.t2011 VGND.t2612 VGND.t2611 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1771 a_n997_3755# XThR.XTBN.Y VGND.t2339 VGND.t2325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1772 XA.XIR[12].XIC[13].icell.SM XA.XIR[12].XIC[13].icell.Ien Iout.t91 VGND.t681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1773 VPWR.t1783 XThR.XTBN.Y XThR.Tn[14].t10 VPWR.t1782 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 XA.XIR[15].XIC[14].icell.SM XA.XIR[15].XIC[14].icell.Ien Iout.t54 VGND.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1775 XA.XIR[4].XIC[6].icell.PUM XThC.Tn[6].t32 XA.XIR[4].XIC[6].icell.Ien VPWR.t1427 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1776 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[8].t55 VGND.t1842 VGND.t1841 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1777 XA.XIR[3].XIC[7].icell.PUM XThC.Tn[7].t26 XA.XIR[3].XIC[7].icell.Ien VPWR.t1157 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1778 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[4].t53 VGND.t1700 VGND.t1699 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1779 XA.XIR[12].XIC[3].icell.PUM XThC.Tn[3].t31 XA.XIR[12].XIC[3].icell.Ien VPWR.t1161 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1780 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2012 VGND.t2614 VGND.t2613 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1781 VPWR.t1361 XThR.Tn[13].t47 XA.XIR[14].XIC[0].icell.PUM VPWR.t1360 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1782 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7].t47 XA.XIR[7].XIC[13].icell.Ien VGND.t678 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1783 XA.XIR[0].XIC[10].icell.Ien XThR.Tn[0].t52 VPWR.t859 VPWR.t858 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1784 XA.XIR[3].XIC[2].icell.SM XA.XIR[3].XIC[2].icell.Ien Iout.t47 VGND.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1785 XA.XIR[6].XIC[8].icell.PUM XThC.Tn[8].t31 XA.XIR[6].XIC[8].icell.Ien VPWR.t1066 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1786 XA.XIR[11].XIC[11].icell.SM XA.XIR[11].XIC[11].icell.Ien Iout.t136 VGND.t927 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1787 XThR.Tn[7].t4 XThR.XTBN.Y VGND.t2331 VGND.t2330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1788 XA.XIR[2].XIC_15.icell.SM XA.XIR[2].XIC_15.icell.Ien Iout.t160 VGND.t1199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1789 VPWR.t146 VPWR.t144 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1790 VGND.t1767 XThC.Tn[9].t32 XA.XIR[4].XIC[9].icell.PDM VGND.t1766 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1791 XA.XIR[14].XIC[4].icell.Ien XThR.Tn[14].t49 VPWR.t771 VPWR.t770 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1792 XA.XIR[7].XIC[1].icell.PUM XThC.Tn[1].t32 XA.XIR[7].XIC[1].icell.Ien VPWR.t1167 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1793 VGND.t2616 VPWR.t2013 XA.XIR[15].XIC_15.icell.PDM VGND.t2615 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1794 XThC.XTB4.Y.t1 XThC.XTB7.B VGND.t1181 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1795 VPWR.t1094 XThR.XTB6.Y XThR.Tn[13].t2 VPWR.t1093 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VPWR.t1048 XThR.XTB3.Y.t11 a_n1049_7493# VPWR.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1797 XA.XIR[1].XIC[5].icell.PUM XThC.Tn[5].t30 XA.XIR[1].XIC[5].icell.Ien VPWR.t1053 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1798 VPWR.t535 XThR.Tn[11].t54 XA.XIR[12].XIC[12].icell.PUM VPWR.t534 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1799 VGND.t1651 Vbias.t163 XA.XIR[7].XIC[5].icell.SM VGND.t1650 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1800 XA.XIR[6].XIC[6].icell.Ien XThR.Tn[6].t50 VPWR.t817 VPWR.t816 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1801 XA.XIR[5].XIC[7].icell.Ien XThR.Tn[5].t49 VPWR.t627 VPWR.t626 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1802 VPWR.t929 data[4].t3 XThR.XTB7.A VPWR.t928 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1803 VGND.t2524 XThC.Tn[4].t33 XA.XIR[7].XIC[4].icell.PDM VGND.t2523 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1804 VGND.t1653 Vbias.t164 XA.XIR[6].XIC[6].icell.SM VGND.t1652 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1805 VGND.t2618 VPWR.t2014 XA.XIR[2].XIC_dummy_right.icell.PDM VGND.t2617 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1806 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2015 VGND.t2620 VGND.t2619 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1807 XA.XIR[15].XIC[6].icell.PDM XThR.Tn[14].t50 VGND.t513 VGND.t512 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1808 XThC.Tn[6].t1 XThC.XTBN.Y.t80 VGND.t1476 VGND.t1475 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1809 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[13].t48 VGND.t1354 VGND.t1353 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1810 XA.XIR[9].XIC[7].icell.Ien XThR.Tn[9].t45 VPWR.t513 VPWR.t512 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1811 XA.XIR[8].XIC[8].icell.Ien XThR.Tn[8].t56 VPWR.t1687 VPWR.t1686 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1812 VPWR.t1114 VGND.t2698 XA.XIR[0].XIC[6].icell.PUM VPWR.t1113 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1813 VPWR.t1281 XThR.Tn[3].t55 XA.XIR[4].XIC[14].icell.PUM VPWR.t1280 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1814 XThR.Tn[5].t1 XThR.XTB6.Y VGND.t935 VGND.t344 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1815 VPWR.t901 XThR.Tn[7].t48 XA.XIR[8].XIC[3].icell.PUM VPWR.t900 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1816 VPWR.t499 XThC.XTB5.Y a_5155_9615# VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1817 VPWR.t143 VPWR.t141 XA.XIR[3].XIC_15.icell.PUM VPWR.t142 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1818 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6].t51 XA.XIR[6].XIC[9].icell.Ien VGND.t566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1819 VPWR.t140 VPWR.t138 XA.XIR[7].XIC_15.icell.PUM VPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1820 VGND.t1655 Vbias.t165 XA.XIR[1].XIC[3].icell.SM VGND.t1654 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1821 XA.XIR[3].XIC[11].icell.PUM XThC.Tn[11].t30 XA.XIR[3].XIC[11].icell.Ien VPWR.t716 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1822 XThR.Tn[4].t2 XThR.XTB5.Y VGND.t349 VGND.t348 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1823 a_4861_9615# XThC.XTB4.Y.t13 VPWR.t1538 VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1824 a_5949_9615# XThC.XTBN.Y.t81 XThC.Tn[5].t5 VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1825 VGND.t1657 Vbias.t166 XA.XIR[4].XIC[4].icell.SM VGND.t1656 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1826 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[5].t50 VGND.t301 VGND.t300 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1827 VGND.t2622 VPWR.t2016 XA.XIR[5].XIC_dummy_left.icell.PDM VGND.t2621 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1828 XA.XIR[11].XIC[9].icell.SM XA.XIR[11].XIC[9].icell.Ien Iout.t184 VGND.t1421 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1829 VGND.t1477 XThC.XTBN.Y.t82 XThC.Tn[2].t7 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1830 VGND.t2624 VPWR.t2017 XA.XIR[9].XIC_dummy_left.icell.PDM VGND.t2623 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1831 XA.XIR[8].XIC[11].icell.SM XA.XIR[8].XIC[11].icell.Ien Iout.t183 VGND.t1420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1832 VPWR.t615 XThC.XTB1.Y.t14 XThC.Tn[8].t5 VPWR.t614 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1833 VGND.t426 XThC.Tn[11].t31 XA.XIR[11].XIC[11].icell.PDM VGND.t425 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1834 a_5155_10571# XThC.XTB7.B XThC.XTB5.Y VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1835 a_10915_9569# XThC.XTBN.Y.t83 VGND.t1479 VGND.t1478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1836 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14].t51 VPWR.t773 VPWR.t772 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1837 XA.XIR[4].XIC[1].icell.PUM XThC.Tn[1].t33 XA.XIR[4].XIC[1].icell.Ien VPWR.t1168 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1838 XA.XIR[3].XIC[2].icell.PUM XThC.Tn[2].t30 XA.XIR[3].XIC[2].icell.Ien VPWR.t1649 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1839 VPWR.t537 XThR.Tn[11].t55 XA.XIR[12].XIC[10].icell.PUM VPWR.t536 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1840 XA.XIR[0].XIC[5].icell.Ien XThR.Tn[0].t53 VPWR.t861 VPWR.t860 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1841 XA.XIR[6].XIC[3].icell.PUM XThC.Tn[3].t32 XA.XIR[6].XIC[3].icell.Ien VPWR.t1162 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1842 VGND.t1659 Vbias.t167 XA.XIR[6].XIC[10].icell.SM VGND.t1658 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1843 XA.XIR[5].XIC[11].icell.Ien XThR.Tn[5].t51 VPWR.t629 VPWR.t628 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1844 XThC.Tn[3].t8 XThC.XTB4.Y.t14 VGND.t1598 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1845 VGND.t1661 Vbias.t168 XA.XIR[3].XIC[6].icell.SM VGND.t1660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1846 VGND.t2526 XThC.Tn[4].t34 XA.XIR[4].XIC[4].icell.PDM VGND.t2525 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1847 VGND.t1117 XThC.Tn[1].t34 XA.XIR[8].XIC[1].icell.PDM VGND.t1116 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1848 VGND.t875 XThC.Tn[5].t31 XA.XIR[3].XIC[5].icell.PDM VGND.t874 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1849 XA.XIR[9].XIC[11].icell.Ien XThR.Tn[9].t46 VPWR.t515 VPWR.t514 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1850 VGND.t1790 XThC.Tn[2].t31 XA.XIR[11].XIC[2].icell.PDM VGND.t1789 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1851 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[3].t56 VGND.t1538 VGND.t1537 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1852 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13].t49 XA.XIR[13].XIC[11].icell.Ien VGND.t1355 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1853 XThR.Tn[3].t5 XThR.XTBN.Y VGND.t2338 VGND.t2337 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1854 XA.XIR[0].XIC[13].icell.PUM XThC.Tn[13].t33 XA.XIR[0].XIC[13].icell.Ien VPWR.t539 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1855 XA.XIR[6].XIC[1].icell.Ien XThR.Tn[6].t52 VPWR.t819 VPWR.t818 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1856 VGND.t1663 Vbias.t169 XA.XIR[7].XIC[0].icell.SM VGND.t1662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1857 VGND.t1665 Vbias.t170 XA.XIR[2].XIC[12].icell.SM VGND.t1664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1858 XA.XIR[5].XIC[2].icell.Ien XThR.Tn[5].t52 VPWR.t631 VPWR.t630 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1859 VGND.t1382 Vbias.t171 XA.XIR[6].XIC[1].icell.SM VGND.t1381 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1860 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t136 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1861 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t9 VGND.t1172 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1862 XA.XIR[9].XIC[2].icell.Ien XThR.Tn[9].t47 VPWR.t517 VPWR.t516 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1863 a_4387_10575# XThC.XTB7.B VGND.t1180 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1864 XA.XIR[4].XIC[14].icell.Ien XThR.Tn[4].t54 VPWR.t1592 VPWR.t1591 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1865 XA.XIR[5].XIC[8].icell.SM XA.XIR[5].XIC[8].icell.Ien Iout.t96 VGND.t706 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1866 XA.XIR[8].XIC[3].icell.Ien XThR.Tn[8].t57 VPWR.t1033 VPWR.t1032 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1867 VPWR.t1112 VGND.t2699 XA.XIR[0].XIC[1].icell.PUM VPWR.t1111 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1868 XA.XIR[3].XIC_15.icell.Ien XThR.Tn[3].t57 VPWR.t1505 VPWR.t1504 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1869 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10].t49 XA.XIR[10].XIC[1].icell.Ien VGND.t1322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1870 XA.XIR[8].XIC[9].icell.SM XA.XIR[8].XIC[9].icell.Ien Iout.t126 VGND.t888 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1871 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6].t53 XA.XIR[6].XIC[4].icell.Ien VGND.t567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1872 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t2018 XA.XIR[1].XIC_dummy_right.icell.Ien VGND.t2625 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1873 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5].t53 XA.XIR[5].XIC[5].icell.Ien VGND.t302 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1874 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13].t50 XA.XIR[13].XIC[2].icell.Ien VGND.t1356 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1875 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9].t48 XA.XIR[9].XIC[5].icell.Ien VGND.t158 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1876 a_10051_9569# XThC.XTBN.Y.t84 VGND.t1480 VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1877 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11].t56 XA.XIR[11].XIC_15.icell.Ien VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1878 XThC.XTB1.Y.t0 XThC.XTB7.B VPWR.t1214 VPWR.t1213 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1879 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t2 VPWR.t1778 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1880 XA.XIR[2].XIC[8].icell.SM XA.XIR[2].XIC[8].icell.Ien Iout.t212 VGND.t1819 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1881 XA.XIR[11].XIC[4].icell.SM XA.XIR[11].XIC[4].icell.Ien Iout.t98 VGND.t716 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1882 VGND.t1384 Vbias.t172 XA.XIR[3].XIC[10].icell.SM VGND.t1383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1883 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t133 VPWR.t135 VPWR.t134 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1884 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout VGND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1885 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t3 VPWR.t1781 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1886 a_7651_9569# XThC.XTBN.Y.t85 VGND.t1481 VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1887 VGND.t992 VGND.t990 XA.XIR[14].XIC_dummy_right.icell.SM VGND.t991 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1888 VGND.t1496 XThC.Tn[6].t33 XA.XIR[11].XIC[6].icell.PDM VGND.t1495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1889 VPWR.t585 XThC.XTB7.A a_6243_10571# VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1890 VPWR.t132 VPWR.t130 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t131 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1891 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[0].t54 VGND.t1147 VGND.t1146 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1892 VPWR.t1829 XThR.Tn[11].t57 XA.XIR[12].XIC[5].icell.PUM VPWR.t1828 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1893 XThC.Tn[10].t7 XThC.XTB3.Y.t13 a_8739_9569# VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1894 VGND.t1386 Vbias.t173 XA.XIR[3].XIC[1].icell.SM VGND.t1385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1895 XA.XIR[7].XIC[5].icell.SM XA.XIR[7].XIC[5].icell.Ien Iout.t56 VGND.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1896 VGND.t2566 XThC.Tn[0].t31 XA.XIR[3].XIC[0].icell.PDM VGND.t2565 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1897 VGND.t2336 XThR.XTBN.Y XThR.Tn[2].t5 VGND.t2335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1898 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[10].t50 VGND.t1123 VGND.t1122 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1899 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[10].t51 VGND.t1125 VGND.t1124 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1900 XA.XIR[10].XIC[6].icell.SM XA.XIR[10].XIC[6].icell.Ien Iout.t66 VGND.t446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1901 XThR.XTB5.A data[5].t3 VGND.t2540 VGND.t2539 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1902 XA.XIR[14].XIC[14].icell.SM XA.XIR[14].XIC[14].icell.Ien Iout.t145 VGND.t1089 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1903 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t128 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t129 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1904 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[3].t58 VGND.t1540 VGND.t1539 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1905 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7].t49 XA.XIR[7].XIC[1].icell.Ien VGND.t679 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1906 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13].t51 XA.XIR[13].XIC[6].icell.Ien VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1907 XThR.Tn[12].t9 XThR.XTBN.Y VPWR.t1780 VPWR.t1779 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1908 VGND.t2627 VPWR.t2019 XA.XIR[14].XIC_dummy_right.icell.PDM VGND.t2626 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1909 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[6].t54 VGND.t569 VGND.t568 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1910 XA.XIR[5].XIC[8].icell.PUM XThC.Tn[8].t32 XA.XIR[5].XIC[8].icell.Ien VPWR.t1067 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1911 XThR.Tn[12].t5 XThR.XTB5.Y a_n997_1803# VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1912 XA.XIR[1].XIC_15.icell.SM XA.XIR[1].XIC_15.icell.Ien Iout.t139 VGND.t930 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1913 XA.XIR[9].XIC[8].icell.PUM XThC.Tn[8].t33 XA.XIR[9].XIC[8].icell.Ien VPWR.t1068 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1914 XThR.Tn[3].t11 XThR.XTB4.Y.t11 VGND.t2680 VGND.t375 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1915 XA.XIR[5].XIC[3].icell.SM XA.XIR[5].XIC[3].icell.Ien Iout.t123 VGND.t883 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1916 VGND.t2334 XThR.XTBN.Y a_n997_2667# VGND.t2333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1917 XA.XIR[9].XIC_15.icell.PDM VPWR.t2020 VGND.t2629 VGND.t2628 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1918 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5].t54 XA.XIR[5].XIC[0].icell.Ien VGND.t1090 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1919 XA.XIR[8].XIC[4].icell.SM XA.XIR[8].XIC[4].icell.Ien Iout.t198 VGND.t1577 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1920 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout VGND.t671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1921 VGND.t1388 Vbias.t174 XA.XIR[13].XIC_15.icell.SM VGND.t1387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1922 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t125 VPWR.t127 VPWR.t126 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1923 XA.XIR[0].XIC[6].icell.PUM XThC.Tn[6].t34 XA.XIR[0].XIC[6].icell.Ien VPWR.t1428 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1924 VGND.t1427 XThC.Tn[14].t32 XA.XIR[13].XIC[14].icell.PDM VGND.t1426 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1925 VGND.t904 XThC.Tn[8].t34 XA.XIR[13].XIC[8].icell.PDM VGND.t903 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1926 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9].t49 XA.XIR[9].XIC[0].icell.Ien VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1927 a_5155_9615# XThC.XTB5.Y VPWR.t498 VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1928 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[4].t55 XA.XIR[4].XIC[12].icell.Ien VGND.t1701 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1929 VPWR.t497 XThC.XTB5.Y XThC.Tn[12].t0 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1930 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[3].t59 XA.XIR[3].XIC[13].icell.Ien VGND.t1541 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1931 VPWR.t775 XThR.Tn[14].t52 XA.XIR[15].XIC[12].icell.PUM VPWR.t774 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1932 XA.XIR[7].XIC_15.icell.PUM VPWR.t123 XA.XIR[7].XIC_15.icell.Ien VPWR.t124 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1933 VPWR.t734 XThR.Tn[13].t52 XA.XIR[14].XIC[13].icell.PUM VPWR.t733 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1934 VPWR.t122 VPWR.t120 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t121 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1935 VGND.t1769 XThC.Tn[9].t33 XA.XIR[0].XIC[9].icell.PDM VGND.t1768 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1936 XThC.Tn[5].t4 XThC.XTBN.Y.t86 a_5949_9615# VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1937 XA.XIR[2].XIC[3].icell.SM XA.XIR[2].XIC[3].icell.Ien Iout.t100 VGND.t718 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1938 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[7].t50 VGND.t336 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1939 VGND.t143 XThC.XTB5.Y XThC.Tn[4].t0 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1940 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t5 VPWR.t1778 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1941 VPWR.t1552 XThR.Tn[1].t49 XA.XIR[2].XIC[7].icell.PUM VPWR.t1551 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1942 VPWR.t1190 XThR.Tn[0].t55 XA.XIR[1].XIC[8].icell.PUM VPWR.t1189 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1943 XA.XIR[10].XIC[10].icell.SM XA.XIR[10].XIC[10].icell.Ien Iout.t45 VGND.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1944 XThC.Tn[2].t6 XThC.XTBN.Y.t87 VGND.t1482 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1945 VPWR.t1594 XThR.Tn[4].t56 XA.XIR[5].XIC[8].icell.PUM VPWR.t1593 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1946 XA.XIR[15].XIC[14].icell.PDM VPWR.t2021 XA.XIR[15].XIC[14].icell.Ien VGND.t2630 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1947 XA.XIR[15].XIC[8].icell.PDM VPWR.t2022 XA.XIR[15].XIC[8].icell.Ien VGND.t2631 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1948 a_5155_9615# XThC.XTBN.Y.t88 XThC.Tn[4].t5 VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1949 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[0].t56 VGND.t1149 VGND.t1148 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1950 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[7].t51 VGND.t338 VGND.t337 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1951 XA.XIR[13].XIC[9].icell.PUM XThC.Tn[9].t34 XA.XIR[13].XIC[9].icell.Ien VPWR.t1599 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1952 XA.XIR[7].XIC[0].icell.SM XA.XIR[7].XIC[0].icell.Ien Iout.t82 VGND.t645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1953 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout VGND.t933 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1954 VPWR.t1747 XThR.XTB7.B XThR.XTB2.Y VPWR.t1744 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1955 XThC.Tn[8].t8 XThC.XTB1.Y.t15 a_7651_9569# VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1956 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[10].t52 VGND.t1127 VGND.t1126 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1957 VGND.t428 XThC.Tn[11].t32 XA.XIR[10].XIC[11].icell.PDM VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1958 XA.XIR[10].XIC[1].icell.SM XA.XIR[10].XIC[1].icell.Ien Iout.t38 VGND.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1959 XA.XIR[6].XIC_15.icell.PDM VPWR.t2023 VGND.t2633 VGND.t2632 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1960 VGND.t1462 XThC.XTB5.A XThC.XTB5.Y VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1961 VGND.t989 VGND.t987 XA.XIR[14].XIC_dummy_left.icell.SM VGND.t988 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1962 VGND.t1359 XThR.XTB7.Y XThR.Tn[6].t0 VGND.t1358 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1963 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[4].t57 XA.XIR[4].XIC[10].icell.Ien VGND.t1702 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1964 XA.XIR[1].XIC[14].icell.PUM XThC.Tn[14].t33 XA.XIR[1].XIC[14].icell.Ien VPWR.t1383 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1965 XA.XIR[5].XIC[3].icell.PUM XThC.Tn[3].t33 XA.XIR[5].XIC[3].icell.Ien VPWR.t1163 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1966 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[6].t55 VGND.t571 VGND.t570 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1967 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[1].t50 VGND.t1602 VGND.t1601 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1968 VPWR.t777 XThR.Tn[14].t53 XA.XIR[15].XIC[10].icell.PUM VPWR.t776 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1969 XA.XIR[9].XIC[3].icell.PUM XThC.Tn[3].t34 XA.XIR[9].XIC[3].icell.Ien VPWR.t1164 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1970 XA.XIR[4].XIC_15.icell.PUM VPWR.t118 XA.XIR[4].XIC_15.icell.Ien VPWR.t119 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1971 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[4].t58 VGND.t1704 VGND.t1703 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1972 XA.XIR[4].XIC[11].icell.SM XA.XIR[4].XIC[11].icell.Ien Iout.t191 VGND.t1502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1973 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2024 VGND.t2635 VGND.t2634 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1974 XA.XIR[15].XIC[9].icell.Ien VPWR.t115 VPWR.t117 VPWR.t116 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1975 VGND.t1792 XThC.Tn[2].t32 XA.XIR[10].XIC[2].icell.PDM VGND.t1791 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1976 XThR.Tn[9].t8 XThR.XTBN.Y VPWR.t1774 VPWR.t1757 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1977 VGND.t1483 XThC.XTBN.Y.t89 a_9827_9569# VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1978 XA.XIR[0].XIC[1].icell.PUM XThC.Tn[1].t35 XA.XIR[0].XIC[1].icell.Ien VPWR.t1169 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1979 VPWR.t1554 XThR.Tn[1].t51 XA.XIR[2].XIC[11].icell.PUM VPWR.t1553 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1980 VGND.t1107 XThC.Tn[3].t35 XA.XIR[13].XIC[3].icell.PDM VGND.t1106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1981 VGND.t2637 VPWR.t2025 XA.XIR[8].XIC_15.icell.PDM VGND.t2636 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1982 VPWR.t1035 XThR.Tn[8].t58 XA.XIR[9].XIC[9].icell.PUM VPWR.t1034 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1983 VGND.t1390 Vbias.t175 XA.XIR[1].XIC[12].icell.SM VGND.t1389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1984 XA.XIR[14].XIC[13].icell.Ien XThR.Tn[14].t54 VPWR.t779 VPWR.t778 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1985 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t112 VPWR.t114 VPWR.t113 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1986 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12].t53 XA.XIR[12].XIC[14].icell.Ien VGND.t1262 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1987 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t110 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t111 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1988 XThC.Tn[0].t2 XThC.XTB1.Y.t16 VGND.t295 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1989 VGND.t1392 Vbias.t176 XA.XIR[0].XIC[5].icell.SM VGND.t1391 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1990 VGND.t1394 Vbias.t177 XA.XIR[4].XIC[13].icell.SM VGND.t1393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1991 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12].t54 XA.XIR[12].XIC[8].icell.Ien VGND.t1263 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1992 VGND.t2528 XThC.Tn[4].t35 XA.XIR[0].XIC[4].icell.PDM VGND.t2527 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1993 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t8 VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1994 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[7].t52 VGND.t340 VGND.t339 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1995 XA.XIR[2].XIC[7].icell.Ien XThR.Tn[2].t49 VPWR.t1457 VPWR.t1456 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1996 VGND.t1396 Vbias.t178 XA.XIR[7].XIC[14].icell.SM VGND.t1395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1997 XA.XIR[6].XIC_15.icell.Ien XThR.Tn[6].t56 VPWR.t821 VPWR.t820 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1998 VPWR.t1556 XThR.Tn[1].t52 XA.XIR[2].XIC[2].icell.PUM VPWR.t1555 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1999 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[10].t53 VGND.t1129 VGND.t1128 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2000 VGND.t194 XThC.Tn[13].t34 XA.XIR[7].XIC[13].icell.PDM VGND.t193 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2001 VPWR.t1192 XThR.Tn[0].t57 XA.XIR[1].XIC[3].icell.PUM VPWR.t1191 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2002 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout VGND.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2003 XThR.Tn[14].t9 XThR.XTBN.Y VPWR.t1777 VPWR.t1776 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2004 VPWR.t1596 XThR.Tn[4].t59 XA.XIR[5].XIC[3].icell.PUM VPWR.t1595 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2005 VPWR.t109 VPWR.t107 XA.XIR[0].XIC_15.icell.PUM VPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2006 VPWR.t736 XThR.Tn[13].t53 XA.XIR[14].XIC[6].icell.PUM VPWR.t735 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2007 XA.XIR[15].XIC[3].icell.PDM VPWR.t2026 XA.XIR[15].XIC[3].icell.Ien VGND.t2638 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2008 a_n997_3755# XThR.XTBN.Y VGND.t2332 VGND.t2317 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2009 XThR.Tn[8].t10 XThR.XTB1.Y.t13 VPWR.t1893 VPWR.t1892 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2010 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10].t54 XA.XIR[10].XIC_15.icell.Ien VGND.t1130 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2011 XA.XIR[0].XIC[14].icell.Ien XThR.Tn[0].t58 VPWR.t1194 VPWR.t1193 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2012 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[1].t53 VGND.t1604 VGND.t1603 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2013 XA.XIR[1].XIC[8].icell.SM XA.XIR[1].XIC[8].icell.Ien Iout.t102 VGND.t726 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2014 VGND.t1398 Vbias.t179 XA.XIR[10].XIC[7].icell.SM VGND.t1397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2015 a_n1049_7787# XThR.XTB2.Y VPWR.t450 VPWR.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2016 XA.XIR[4].XIC[9].icell.SM XA.XIR[4].XIC[9].icell.Ien Iout.t6 VGND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2017 VGND.t1498 XThC.Tn[6].t35 XA.XIR[10].XIC[6].icell.PDM VGND.t1497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2018 VPWR.t1307 XThR.Tn[12].t55 XA.XIR[13].XIC[4].icell.PUM VPWR.t1306 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2019 a_n1331_2891# data[5].t4 VGND.t384 VGND.t383 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2020 VGND.t1400 Vbias.t180 XA.XIR[13].XIC[8].icell.SM VGND.t1399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2021 XA.XIR[12].XIC[9].icell.Ien XThR.Tn[12].t56 VPWR.t1309 VPWR.t1308 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2022 VPWR.t106 VPWR.t104 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t105 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2023 VGND.t1095 XThC.Tn[7].t27 XA.XIR[13].XIC[7].icell.PDM VGND.t1094 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2024 VPWR.t781 XThR.Tn[14].t55 XA.XIR[15].XIC[5].icell.PUM VPWR.t780 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2025 XThR.XTB7.B data[6].t1 VGND.t787 VGND.t786 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2026 XThR.Tn[2].t9 XThR.XTBN.Y a_n1049_7493# VPWR.t1775 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2027 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[9].t50 VGND.t161 VGND.t160 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2028 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[9].t51 VGND.t163 VGND.t162 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2029 XA.XIR[2].XIC[11].icell.Ien XThR.Tn[2].t50 VPWR.t1455 VPWR.t1454 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2030 XA.XIR[9].XIC[6].icell.SM XA.XIR[9].XIC[6].icell.Ien Iout.t239 VGND.t2417 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2031 VGND.t743 XThC.Tn[12].t34 XA.XIR[1].XIC[12].icell.PDM VGND.t742 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2032 VGND.t196 XThC.Tn[13].t35 XA.XIR[4].XIC[13].icell.PDM VGND.t195 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2033 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t2027 XA.XIR[4].XIC_dummy_left.icell.Ien VGND.t2639 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2034 XA.XIR[15].XIC[7].icell.PDM VPWR.t2028 XA.XIR[15].XIC[7].icell.Ien VGND.t2640 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2035 VGND.t1402 Vbias.t181 XA.XIR[0].XIC[0].icell.SM VGND.t1401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2036 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12].t57 XA.XIR[12].XIC[3].icell.Ien VGND.t1988 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2037 VPWR.t1421 XThC.XTBN.Y.t90 XThC.Tn[8].t2 VPWR.t1420 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2038 XThR.Tn[10].t0 XThR.XTB3.Y.t12 VPWR.t477 VPWR.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2039 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7].t53 XA.XIR[7].XIC_15.icell.Ien VGND.t341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2040 XA.XIR[11].XIC[4].icell.PUM XThC.Tn[4].t36 XA.XIR[11].XIC[4].icell.Ien VPWR.t1868 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2041 XThR.Tn[4].t9 XThR.XTBN.Y VGND.t2329 VGND.t2328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2042 XA.XIR[15].XIC[12].icell.PUM XThC.Tn[12].t35 XA.XIR[15].XIC[12].icell.Ien VPWR.t964 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2043 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t102 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2044 XA.XIR[2].XIC[2].icell.Ien XThR.Tn[2].t51 VPWR.t1453 VPWR.t1452 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2045 XA.XIR[11].XIC[13].icell.SM XA.XIR[11].XIC[13].icell.Ien Iout.t214 VGND.t1830 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2046 VGND.t2286 XThR.XTB7.B XThR.XTB5.Y VGND.t2285 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2047 VGND.t1404 Vbias.t182 XA.XIR[12].XIC_15.icell.SM VGND.t1403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2048 VGND.t266 XThC.Tn[14].t34 XA.XIR[12].XIC[14].icell.PDM VGND.t265 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2049 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[3].t60 XA.XIR[3].XIC[1].icell.Ien VGND.t1542 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2050 XA.XIR[14].XIC[6].icell.Ien XThR.Tn[14].t56 VPWR.t783 VPWR.t782 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2051 VGND.t2394 XThC.Tn[8].t35 XA.XIR[12].XIC[8].icell.PDM VGND.t2393 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2052 VPWR.t738 XThR.Tn[13].t54 XA.XIR[14].XIC[1].icell.PUM VPWR.t737 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2053 XA.XIR[2].XIC[7].icell.PUM XThC.Tn[7].t28 XA.XIR[2].XIC[7].icell.Ien VPWR.t1158 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2054 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[2].t52 XA.XIR[2].XIC[5].icell.Ien VGND.t524 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2055 VPWR.t1712 XThR.Tn[12].t58 XA.XIR[13].XIC[0].icell.PUM VPWR.t1711 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2056 VPWR.t519 XThR.Tn[9].t52 XA.XIR[10].XIC[4].icell.PUM VPWR.t518 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2057 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6].t57 XA.XIR[6].XIC[13].icell.Ien VGND.t572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2058 XA.XIR[1].XIC[3].icell.SM XA.XIR[1].XIC[3].icell.Ien Iout.t103 VGND.t728 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2059 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14].t57 XA.XIR[14].XIC[9].icell.Ien VGND.t514 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2060 VPWR.t1831 XThR.Tn[11].t58 XA.XIR[12].XIC[14].icell.PUM VPWR.t1830 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2061 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t5 VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2062 XThC.Tn[4].t4 XThC.XTBN.Y.t91 a_5155_9615# VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2063 XA.XIR[13].XIC[4].icell.Ien XThR.Tn[13].t55 VPWR.t740 VPWR.t739 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2064 VGND.t1715 Vbias.t183 XA.XIR[10].XIC[2].icell.SM VGND.t1714 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2065 XA.XIR[4].XIC[4].icell.SM XA.XIR[4].XIC[4].icell.Ien Iout.t218 VGND.t1849 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2066 VGND.t1717 Vbias.t184 XA.XIR[9].XIC_15.icell.SM VGND.t1716 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2067 XA.XIR[9].XIC[10].icell.SM XA.XIR[9].XIC[10].icell.Ien Iout.t152 VGND.t1142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2068 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t99 VPWR.t101 VPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2069 VGND.t400 XThC.Tn[10].t35 XA.XIR[1].XIC[10].icell.PDM VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2070 VGND.t1719 Vbias.t185 XA.XIR[13].XIC[3].icell.SM VGND.t1718 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2071 XA.XIR[0].XIC[12].icell.PDM XThR.Tn[0].t59 XA.XIR[0].XIC[12].icell.Ien VGND.t1150 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2072 VPWR.t1507 XThR.Tn[3].t61 XA.XIR[4].XIC[8].icell.PUM VPWR.t1506 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2073 VGND.t2327 XThR.XTBN.Y a_n997_1579# VGND.t2309 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2074 VPWR.t1171 XThR.Tn[10].t55 XA.XIR[11].XIC[12].icell.PUM VPWR.t1170 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2075 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2029 VGND.t2642 VGND.t2641 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2076 XA.XIR[12].XIC[9].icell.PUM XThC.Tn[9].t35 XA.XIR[12].XIC[9].icell.Ien VPWR.t1600 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2077 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12].t59 XA.XIR[12].XIC[7].icell.Ien VGND.t1989 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2078 XA.XIR[15].XIC[10].icell.PUM XThC.Tn[10].t36 XA.XIR[15].XIC[10].icell.Ien VPWR.t703 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2079 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[9].t53 VGND.t165 VGND.t164 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2080 XA.XIR[5].XIC[12].icell.SM XA.XIR[5].XIC[12].icell.Ien Iout.t5 VGND.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2081 XA.XIR[9].XIC[1].icell.SM XA.XIR[9].XIC[1].icell.Ien Iout.t94 VGND.t689 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2082 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t5 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2083 XA.XIR[11].XIC[0].icell.PUM XThC.Tn[0].t32 XA.XIR[11].XIC[0].icell.Ien VPWR.t1883 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2084 XA.XIR[8].XIC[13].icell.SM XA.XIR[8].XIC[13].icell.Ien Iout.t168 VGND.t1337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2085 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t97 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2086 XA.XIR[7].XIC[14].icell.SM XA.XIR[7].XIC[14].icell.Ien Iout.t110 VGND.t780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2087 XA.XIR[2].XIC[11].icell.PUM XThC.Tn[11].t33 XA.XIR[2].XIC[11].icell.Ien VPWR.t717 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2088 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[4].t60 VGND.t1751 VGND.t1750 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2089 XA.XIR[0].XIC[5].icell.PDM VGND.t984 VGND.t986 VGND.t985 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2090 VPWR.t1231 XThR.Tn[9].t54 XA.XIR[10].XIC[0].icell.PUM VPWR.t1230 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2091 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[3].t62 VGND.t1544 VGND.t1543 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2092 XA.XIR[2].XIC[12].icell.SM XA.XIR[2].XIC[12].icell.Ien Iout.t226 VGND.t2092 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2093 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[11].t59 VGND.t2420 VGND.t2419 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2094 VGND.t1109 XThC.Tn[3].t36 XA.XIR[12].XIC[3].icell.PDM VGND.t1108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2095 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14].t58 VPWR.t785 VPWR.t784 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2096 XThR.XTBN.Y XThR.XTBN.A VPWR.t1291 VPWR.t1290 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2097 VGND.t1721 Vbias.t186 XA.XIR[15].XIC[11].icell.SM VGND.t1720 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2098 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13].t56 VPWR.t742 VPWR.t741 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2099 VPWR.t665 XThR.Tn[7].t54 XA.XIR[8].XIC[9].icell.PUM VPWR.t664 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2100 VGND.t268 XThC.Tn[14].t35 XA.XIR[6].XIC[14].icell.PDM VGND.t267 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2101 XA.XIR[0].XIC[10].icell.PDM XThR.Tn[0].t60 XA.XIR[0].XIC[10].icell.Ien VGND.t1151 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2102 XA.XIR[2].XIC[2].icell.PUM XThC.Tn[2].t33 XA.XIR[2].XIC[2].icell.Ien VPWR.t1650 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2103 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[2].t53 XA.XIR[2].XIC[0].icell.Ien VGND.t535 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2104 VGND.t2396 XThC.Tn[8].t36 XA.XIR[6].XIC[8].icell.PDM VGND.t2395 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2105 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t94 VPWR.t96 VPWR.t95 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2106 VPWR.t1173 XThR.Tn[10].t56 XA.XIR[11].XIC[10].icell.PUM VPWR.t1172 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2107 XA.XIR[0].XIC_15.icell.PUM VPWR.t92 XA.XIR[0].XIC_15.icell.Ien VPWR.t93 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2108 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14].t59 XA.XIR[14].XIC[4].icell.Ien VGND.t515 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2109 XA.XIR[1].XIC[7].icell.Ien XThR.Tn[1].t54 VPWR.t1558 VPWR.t1557 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2110 VGND.t1723 Vbias.t187 XA.XIR[2].XIC[6].icell.SM VGND.t1722 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2111 VGND.t1119 XThC.Tn[1].t36 XA.XIR[7].XIC[1].icell.PDM VGND.t1118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2112 VGND.t877 XThC.Tn[5].t32 XA.XIR[2].XIC[5].icell.PDM VGND.t876 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2113 VPWR.t1773 XThR.XTBN.Y XThR.Tn[11].t5 VPWR.t1753 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2114 XA.XIR[4].XIC[8].icell.Ien XThR.Tn[4].t61 VPWR.t1622 VPWR.t1621 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2115 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[9].t55 VGND.t1209 VGND.t1208 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2116 VPWR.t569 data[1].t4 XThC.XTB7.A VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2117 VPWR.t1509 XThR.Tn[3].t63 XA.XIR[4].XIC[3].icell.PUM VPWR.t1508 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2118 XA.XIR[11].XIC[12].icell.Ien XThR.Tn[11].t60 VPWR.t1833 VPWR.t1832 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2119 a_8739_9569# XThC.XTBN.Y.t92 VGND.t313 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2120 VGND.t1246 XThR.XTBN.A XThR.XTBN.Y VGND.t1245 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 XThC.Tn[6].t10 XThC.XTB7.Y VGND.t1171 VGND.t1170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2122 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8].t59 XA.XIR[8].XIC[14].icell.Ien VGND.t848 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2123 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8].t60 XA.XIR[8].XIC[8].icell.Ien VGND.t849 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2124 XA.XIR[15].XIC[5].icell.PUM XThC.Tn[5].t33 XA.XIR[15].XIC[5].icell.Ien VPWR.t1054 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2125 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[0].t61 VGND.t831 VGND.t830 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2126 XA.XIR[6].XIC[9].icell.PUM XThC.Tn[9].t36 XA.XIR[6].XIC[9].icell.Ien VPWR.t1601 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2127 XThR.Tn[12].t4 XThR.XTB5.Y a_n997_1803# VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2128 VGND.t2644 VPWR.t2030 XA.XIR[1].XIC_dummy_left.icell.PDM VGND.t2643 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2129 VGND.t1725 Vbias.t188 XA.XIR[12].XIC[8].icell.SM VGND.t1724 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2130 VGND.t430 XThC.Tn[11].t34 XA.XIR[3].XIC[11].icell.PDM VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2131 VGND.t1097 XThC.Tn[7].t29 XA.XIR[12].XIC[7].icell.PDM VGND.t1096 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2132 VGND.t1727 Vbias.t189 XA.XIR[15].XIC[9].icell.SM VGND.t1726 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2133 a_n997_3979# XThR.XTBN.Y VGND.t2326 VGND.t2325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2134 XThC.XTB7.Y XThC.XTB7.B VGND.t1179 VGND.t1178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2135 XA.XIR[0].XIC[0].icell.PDM VGND.t981 VGND.t983 VGND.t982 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2136 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t89 VPWR.t91 VPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2137 VGND.t1729 Vbias.t190 XA.XIR[6].XIC[7].icell.SM VGND.t1728 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2138 XA.XIR[1].XIC[11].icell.Ien XThR.Tn[1].t55 VPWR.t1560 VPWR.t1559 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2139 VGND.t1731 Vbias.t191 XA.XIR[2].XIC[10].icell.SM VGND.t1730 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2140 XThC.Tn[8].t1 XThC.XTBN.Y.t93 VPWR.t636 VPWR.t635 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2141 VGND.t699 XThC.Tn[1].t37 XA.XIR[4].XIC[1].icell.PDM VGND.t698 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2142 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[11].t61 VGND.t2422 VGND.t2421 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2143 VGND.t1794 XThC.Tn[2].t34 XA.XIR[3].XIC[2].icell.PDM VGND.t1793 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2144 VGND.t1733 Vbias.t192 XA.XIR[9].XIC[8].icell.SM VGND.t1732 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2145 XA.XIR[14].XIC[7].icell.PUM XThC.Tn[7].t30 XA.XIR[14].XIC[7].icell.Ien VPWR.t1159 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2146 XA.XIR[8].XIC[9].icell.Ien XThR.Tn[8].t61 VPWR.t1037 VPWR.t1036 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2147 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t2031 VGND.t2646 VGND.t2645 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2148 VGND.t2084 XThC.Tn[3].t37 XA.XIR[6].XIC[3].icell.PDM VGND.t2083 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2149 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5].t55 XA.XIR[5].XIC[11].icell.Ien VGND.t1091 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2150 XA.XIR[11].XIC[10].icell.Ien XThR.Tn[11].t62 VPWR.t1835 VPWR.t1834 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2151 a_n1049_6699# XThR.XTB4.Y.t12 VPWR.t573 VPWR.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2152 XA.XIR[13].XIC_15.icell.SM XA.XIR[13].XIC_15.icell.Ien Iout.t9 VGND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2153 VPWR.t1175 XThR.Tn[10].t57 XA.XIR[11].XIC[5].icell.PUM VPWR.t1174 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2154 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9].t56 XA.XIR[9].XIC[11].icell.Ien VGND.t1210 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2155 XA.XIR[10].XIC[4].icell.PUM XThC.Tn[4].t37 XA.XIR[10].XIC[4].icell.Ien VPWR.t1375 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2156 XA.XIR[1].XIC[2].icell.Ien XThR.Tn[1].t56 VPWR.t838 VPWR.t837 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2157 VGND.t1735 Vbias.t193 XA.XIR[2].XIC[1].icell.SM VGND.t1734 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2158 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t87 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2159 XA.XIR[6].XIC[5].icell.SM XA.XIR[6].XIC[5].icell.Ien Iout.t224 VGND.t2082 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2160 VGND.t2568 XThC.Tn[0].t33 XA.XIR[2].XIC[0].icell.PDM VGND.t2567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2161 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t85 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2162 XA.XIR[4].XIC[3].icell.Ien XThR.Tn[4].t62 VPWR.t1624 VPWR.t1623 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2163 VGND.t1737 Vbias.t194 XA.XIR[0].XIC[14].icell.SM VGND.t1736 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2164 VGND.t1906 Vbias.t195 XA.XIR[14].XIC[5].icell.SM VGND.t1905 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2165 VGND.t198 XThC.Tn[13].t36 XA.XIR[0].XIC[13].icell.PDM VGND.t197 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2166 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6].t58 XA.XIR[6].XIC[1].icell.Ien VGND.t573 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2167 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t2032 XA.XIR[0].XIC_dummy_left.icell.Ien VGND.t2647 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2168 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[1].t57 XA.XIR[1].XIC[5].icell.Ien VGND.t588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2169 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5].t56 XA.XIR[5].XIC[2].icell.Ien VGND.t1092 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2170 VGND.t2649 VPWR.t2033 XA.XIR[13].XIC_dummy_right.icell.PDM VGND.t2648 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2171 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9].t57 XA.XIR[9].XIC[2].icell.Ien VGND.t1211 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2172 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8].t62 XA.XIR[8].XIC[3].icell.Ien VGND.t850 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2173 XA.XIR[3].XIC_15.icell.PDM XThR.Tn[3].t64 XA.XIR[3].XIC_15.icell.Ien VGND.t1545 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2174 VGND.t1852 data[1].t5 XThC.XTB6.A VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2175 VPWR.t787 XThR.Tn[14].t60 XA.XIR[15].XIC[14].icell.PUM VPWR.t786 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2176 VPWR.t84 VPWR.t82 XA.XIR[14].XIC_15.icell.PUM VPWR.t83 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2177 a_n997_2891# XThR.XTBN.Y VGND.t2324 VGND.t2323 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2178 VGND.t1908 Vbias.t196 XA.XIR[12].XIC[3].icell.SM VGND.t1907 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2179 VGND.t1910 Vbias.t197 XA.XIR[3].XIC[7].icell.SM VGND.t1909 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2180 VGND.t1500 XThC.Tn[6].t36 XA.XIR[3].XIC[6].icell.PDM VGND.t1499 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2181 XA.XIR[14].XIC[11].icell.PUM XThC.Tn[11].t35 XA.XIR[14].XIC[11].icell.Ien VPWR.t718 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2182 VPWR.t1146 XThR.Tn[5].t57 XA.XIR[6].XIC[4].icell.PUM VPWR.t1145 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2183 VPWR.t81 VPWR.t79 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t80 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2184 VGND.t1912 Vbias.t198 XA.XIR[15].XIC[4].icell.SM VGND.t1911 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2185 VGND.t980 VGND.t978 XA.XIR[10].XIC_dummy_right.icell.SM VGND.t979 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2186 VGND.t1099 XThC.Tn[7].t31 XA.XIR[6].XIC[7].icell.PDM VGND.t1098 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2187 VPWR.t78 VPWR.t76 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2188 VPWR.t1714 XThR.Tn[12].t60 XA.XIR[13].XIC[13].icell.PUM VPWR.t1713 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2189 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t2034 XA.XIR[15].XIC_dummy_right.icell.Ien VGND.t2650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2190 XThR.Tn[11].t0 XThR.XTB4.Y.t13 a_n997_2667# VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2191 VGND.t1914 Vbias.t199 XA.XIR[6].XIC[2].icell.SM VGND.t1913 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2192 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[6].t59 VGND.t575 VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2193 VPWR.t495 XThC.XTB5.Y a_5155_9615# VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2194 XA.XIR[10].XIC[0].icell.PUM XThC.Tn[0].t34 XA.XIR[10].XIC[0].icell.Ien VPWR.t1884 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2195 XA.XIR[3].XIC[5].icell.SM XA.XIR[3].XIC[5].icell.Ien Iout.t12 VGND.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2196 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[2].t54 VGND.t534 VGND.t533 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2197 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[2].t55 VGND.t532 VGND.t531 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2198 VGND.t1916 Vbias.t200 XA.XIR[9].XIC[3].icell.SM VGND.t1915 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2199 XA.XIR[14].XIC[2].icell.PUM XThC.Tn[2].t35 XA.XIR[14].XIC[2].icell.Ien VPWR.t1651 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2200 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5].t58 XA.XIR[5].XIC[6].icell.Ien VGND.t1093 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2201 XA.XIR[11].XIC[5].icell.Ien XThR.Tn[11].t63 VPWR.t1837 VPWR.t1836 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2202 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[3].t65 VGND.t1547 VGND.t1546 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2203 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9].t58 XA.XIR[9].XIC[6].icell.Ien VGND.t1212 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2204 VGND.t879 XThC.Tn[5].t34 XA.XIR[14].XIC[5].icell.PDM VGND.t878 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2205 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8].t63 XA.XIR[8].XIC[7].icell.Ien VGND.t851 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2206 VGND.t2322 XThR.XTBN.Y XThR.Tn[0].t7 VGND.t2321 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2207 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[6].t60 VGND.t130 VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2208 XA.XIR[1].XIC[8].icell.PUM XThC.Tn[8].t37 XA.XIR[1].XIC[8].icell.Ien VPWR.t1821 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2209 a_n1049_6405# XThR.XTB5.Y VPWR.t670 VPWR.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2210 XA.XIR[6].XIC[0].icell.SM XA.XIR[6].XIC[0].icell.Ien Iout.t253 VGND.t2562 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2211 XThR.Tn[8].t11 XThR.XTB1.Y.t14 VPWR.t1895 VPWR.t1894 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2212 XA.XIR[1].XIC[12].icell.SM XA.XIR[1].XIC[12].icell.Ien Iout.t80 VGND.t608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2213 XA.XIR[8].XIC[12].icell.PUM XThC.Tn[12].t36 XA.XIR[8].XIC[12].icell.Ien VPWR.t965 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2214 VGND.t1918 Vbias.t201 XA.XIR[14].XIC[0].icell.SM VGND.t1917 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2215 XA.XIR[15].XIC[9].icell.PDM XThR.Tn[14].t61 VGND.t517 VGND.t516 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2216 XA.XIR[4].XIC[13].icell.SM XA.XIR[4].XIC[13].icell.Ien Iout.t245 VGND.t2534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2217 XA.XIR[5].XIC_15.icell.PDM VPWR.t2035 VGND.t2652 VGND.t2651 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2218 VGND.t1920 Vbias.t202 XA.XIR[5].XIC_15.icell.SM VGND.t1919 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2219 XA.XIR[11].XIC[13].icell.PUM XThC.Tn[13].t37 XA.XIR[11].XIC[13].icell.Ien VPWR.t540 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2220 VGND.t2398 XThC.Tn[8].t38 XA.XIR[5].XIC[8].icell.PDM VGND.t2397 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2221 VGND.t270 XThC.Tn[14].t36 XA.XIR[5].XIC[14].icell.PDM VGND.t269 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2222 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[1].t58 XA.XIR[1].XIC[0].icell.Ien VGND.t589 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2223 VGND.t1922 Vbias.t203 XA.XIR[13].XIC[12].icell.SM VGND.t1921 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2224 XThR.Tn[1].t1 XThR.XTB2.Y VGND.t100 VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2225 VGND.t272 XThC.Tn[14].t37 XA.XIR[9].XIC[14].icell.PDM VGND.t271 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2226 VGND.t2400 XThC.Tn[8].t39 XA.XIR[9].XIC[8].icell.PDM VGND.t2399 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2227 VPWR.t1148 XThR.Tn[5].t59 XA.XIR[6].XIC[0].icell.PUM VPWR.t1147 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2228 VGND.t314 XThC.XTBN.Y.t94 a_8739_9569# VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2229 XA.XIR[14].XIC_15.icell.Ien XThR.Tn[14].t62 VPWR.t789 VPWR.t788 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2230 VGND.t1924 Vbias.t204 XA.XIR[1].XIC[6].icell.SM VGND.t1923 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2231 VPWR.t75 VPWR.t73 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t74 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2232 XThC.Tn[1].t10 XThC.XTB2.Y VGND.t2095 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2233 VGND.t1169 XThC.XTB7.Y XThC.Tn[6].t9 VGND.t1168 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2234 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t2036 XA.XIR[12].XIC_dummy_right.icell.Ien VGND.t2653 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2235 VPWR.t1233 XThR.Tn[9].t59 XA.XIR[10].XIC[13].icell.PUM VPWR.t1232 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2236 VPWR.t72 VPWR.t70 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2237 a_6243_9615# XThC.XTBN.Y.t95 XThC.Tn[6].t5 VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2238 VGND.t1926 Vbias.t205 XA.XIR[3].XIC[2].icell.SM VGND.t1925 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2239 VGND.t1928 Vbias.t206 XA.XIR[11].XIC[11].icell.SM VGND.t1927 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2240 XA.XIR[10].XIC[12].icell.Ien XThR.Tn[10].t58 VPWR.t1177 VPWR.t1176 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2241 XThR.Tn[2].t8 XThR.XTBN.Y a_n1049_7493# VPWR.t1772 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2242 VGND.t2655 VPWR.t2037 XA.XIR[7].XIC_15.icell.PDM VGND.t2654 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2243 XA.XIR[10].XIC[7].icell.SM XA.XIR[10].XIC[7].icell.Ien Iout.t84 VGND.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2244 XA.XIR[13].XIC[13].icell.Ien XThR.Tn[13].t57 VPWR.t758 VPWR.t757 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2245 XA.XIR[13].XIC[8].icell.SM XA.XIR[13].XIC[8].icell.Ien Iout.t148 VGND.t1132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2246 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[0].t62 VGND.t833 VGND.t832 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2247 XThR.Tn[13].t8 XThR.XTBN.Y VPWR.t1771 VPWR.t1770 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2248 XA.XIR[5].XIC[9].icell.PUM XThC.Tn[9].t37 XA.XIR[5].XIC[9].icell.Ien VPWR.t1602 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2249 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[6].t61 VGND.t132 VGND.t131 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2250 XA.XIR[0].XIC[8].icell.Ien XThR.Tn[0].t63 VPWR.t1011 VPWR.t1010 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2251 XA.XIR[3].XIC[0].icell.SM XA.XIR[3].XIC[0].icell.Ien Iout.t87 VGND.t659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2252 XA.XIR[9].XIC[9].icell.PUM XThC.Tn[9].t38 XA.XIR[9].XIC[9].icell.Ien VPWR.t1603 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2253 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[2].t56 VGND.t530 VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2254 XThR.Tn[10].t5 XThR.XTB3.Y.t13 VPWR.t1178 VPWR.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2255 XA.XIR[8].XIC[10].icell.PUM XThC.Tn[10].t37 XA.XIR[8].XIC[10].icell.Ien VPWR.t704 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2256 XThR.Tn[4].t8 XThR.XTBN.Y VGND.t2320 VGND.t2319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2257 VPWR.t1716 XThR.Tn[12].t61 XA.XIR[13].XIC[6].icell.PUM VPWR.t1715 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2258 VGND.t977 VGND.t975 XA.XIR[10].XIC_dummy_left.icell.SM VGND.t976 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2259 VGND.t934 XThR.XTB6.Y XThR.Tn[5].t0 VGND.t342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2260 VGND.t2570 XThC.Tn[0].t35 XA.XIR[14].XIC[0].icell.PDM VGND.t2569 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2261 XA.XIR[1].XIC[3].icell.PUM XThC.Tn[3].t38 XA.XIR[1].XIC[3].icell.Ien VPWR.t1731 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2262 VGND.t2236 Vbias.t207 XA.XIR[1].XIC[10].icell.SM VGND.t2235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2263 a_4861_9615# XThC.XTBN.Y.t96 XThC.Tn[3].t5 VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2264 XA.XIR[15].XIC[4].icell.PDM XThR.Tn[14].t63 VGND.t519 VGND.t518 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2265 XA.XIR[0].XIC[11].icell.SM XA.XIR[0].XIC[11].icell.Ien Iout.t128 VGND.t898 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2266 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[13].t58 VGND.t463 VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2267 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2038 VGND.t2657 VGND.t2656 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2268 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t4 VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2269 VGND.t2086 XThC.Tn[3].t39 XA.XIR[5].XIC[3].icell.PDM VGND.t2085 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2270 VGND.t2238 Vbias.t208 XA.XIR[11].XIC[9].icell.SM VGND.t2237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2271 XA.XIR[10].XIC[10].icell.Ien XThR.Tn[10].t59 VPWR.t1612 VPWR.t1611 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2272 XA.XIR[12].XIC_15.icell.SM XA.XIR[12].XIC_15.icell.Ien Iout.t86 VGND.t658 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2273 VGND.t2088 XThC.Tn[3].t40 XA.XIR[9].XIC[3].icell.PDM VGND.t2087 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2274 VGND.t2240 Vbias.t209 XA.XIR[8].XIC[11].icell.SM VGND.t2239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2275 XA.XIR[7].XIC[12].icell.Ien XThR.Tn[7].t55 VPWR.t667 VPWR.t666 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2276 VPWR.t1013 XThR.Tn[0].t64 XA.XIR[1].XIC[9].icell.PUM VPWR.t1012 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2277 VGND.t2659 VPWR.t2039 XA.XIR[4].XIC_15.icell.PDM VGND.t2658 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2278 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t67 VPWR.t69 VPWR.t68 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2279 VGND.t2242 Vbias.t210 XA.XIR[1].XIC[1].icell.SM VGND.t2241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2280 VPWR.t1626 XThR.Tn[4].t63 XA.XIR[5].XIC[9].icell.PUM VPWR.t1625 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2281 VGND.t701 XThC.Tn[1].t38 XA.XIR[0].XIC[1].icell.PDM VGND.t700 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2282 XA.XIR[11].XIC[6].icell.PUM XThC.Tn[6].t37 XA.XIR[11].XIC[6].icell.Ien VPWR.t695 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2283 XA.XIR[15].XIC[14].icell.PUM XThC.Tn[14].t38 XA.XIR[15].XIC[14].icell.Ien VPWR.t592 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2284 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[2].t57 VGND.t528 VGND.t527 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2285 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14].t64 XA.XIR[14].XIC[13].icell.Ien VGND.t2428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2286 VGND.t2661 VPWR.t2040 XA.XIR[12].XIC_dummy_right.icell.PDM VGND.t2660 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2287 XA.XIR[10].XIC[2].icell.SM XA.XIR[10].XIC[2].icell.Ien Iout.t22 VGND.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2288 VGND.t1707 XThC.Tn[9].t39 XA.XIR[11].XIC[9].icell.PDM VGND.t1706 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2289 VPWR.t830 XThR.XTB3.Y.t14 a_n1049_7493# VPWR.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2290 XA.XIR[13].XIC[3].icell.SM XA.XIR[13].XIC[3].icell.Ien Iout.t132 VGND.t909 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2291 VPWR.t1235 XThR.Tn[9].t60 XA.XIR[10].XIC[6].icell.PUM VPWR.t1234 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2292 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6].t62 XA.XIR[6].XIC_15.icell.Ien VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2293 VPWR.t1572 XThR.Tn[11].t64 XA.XIR[12].XIC[8].icell.PUM VPWR.t1571 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2294 XA.XIR[0].XIC[3].icell.Ien XThR.Tn[0].t65 VPWR.t1015 VPWR.t1014 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2295 XA.XIR[8].XIC[5].icell.PUM XThC.Tn[5].t35 XA.XIR[8].XIC[5].icell.Ien VPWR.t1055 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2296 XA.XIR[13].XIC[6].icell.Ien XThR.Tn[13].t59 VPWR.t760 VPWR.t759 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2297 XA.XIR[0].XIC[9].icell.SM XA.XIR[0].XIC[9].icell.Ien Iout.t223 VGND.t2081 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2298 VGND.t2244 Vbias.t211 XA.XIR[5].XIC[8].icell.SM VGND.t2243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2299 VGND.t1101 XThC.Tn[7].t32 XA.XIR[5].XIC[7].icell.PDM VGND.t1100 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2300 VPWR.t1718 XThR.Tn[12].t62 XA.XIR[13].XIC[1].icell.PUM VPWR.t1717 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2301 XThC.XTB2.Y XThC.XTB6.A a_3523_10575# VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2302 VPWR.t66 VPWR.t64 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2303 VGND.t1902 XThC.Tn[7].t33 XA.XIR[9].XIC[7].icell.PDM VGND.t1901 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2304 VGND.t2246 Vbias.t212 XA.XIR[8].XIC[9].icell.SM VGND.t2245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2305 XA.XIR[7].XIC[10].icell.Ien XThR.Tn[7].t56 VPWR.t669 VPWR.t668 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2306 XThR.Tn[4].t1 XThR.XTB5.Y VGND.t345 VGND.t344 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2307 VPWR.t1769 XThR.XTBN.Y XThR.Tn[14].t8 VPWR.t1768 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2308 VPWR.t1614 XThR.Tn[10].t60 XA.XIR[11].XIC[14].icell.PUM VPWR.t1613 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2309 XThC.Tn[13].t5 XThC.XTB6.Y VPWR.t1408 VPWR.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2310 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13].t60 XA.XIR[13].XIC[9].icell.Ien VGND.t464 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2311 VGND.t1457 XThC.XTB6.Y XThC.Tn[5].t8 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2312 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[13].t61 VGND.t466 VGND.t465 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2313 XA.XIR[5].XIC[6].icell.SM XA.XIR[5].XIC[6].icell.Ien Iout.t238 VGND.t2416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2314 VPWR.t1767 XThR.XTBN.Y XThR.Tn[11].t4 VPWR.t1766 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2315 VGND.t2248 Vbias.t213 XA.XIR[11].XIC[4].icell.SM VGND.t2247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2316 XA.XIR[10].XIC[5].icell.Ien XThR.Tn[10].t61 VPWR.t1616 VPWR.t1615 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2317 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[12].t63 VGND.t1991 VGND.t1990 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2318 VGND.t974 VGND.t972 XA.XIR[6].XIC_dummy_right.icell.SM VGND.t973 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2319 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[11].t65 VGND.t1613 VGND.t1612 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2320 XA.XIR[15].XIC[11].icell.SM XA.XIR[15].XIC[11].icell.Ien Iout.t236 VGND.t2392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2321 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[2].t58 XA.XIR[2].XIC[11].icell.Ien VGND.t526 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2322 XA.XIR[3].XIC[4].icell.PUM XThC.Tn[4].t38 XA.XIR[3].XIC[4].icell.Ien VPWR.t1376 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2323 XThC.Tn[9].t8 XThC.XTB2.Y a_7875_9569# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2324 XA.XIR[4].XIC_15.icell.PDM VPWR.t2041 VGND.t2663 VGND.t2662 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2325 XA.XIR[11].XIC[1].icell.PUM XThC.Tn[1].t39 XA.XIR[11].XIC[1].icell.Ien VPWR.t919 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2326 VGND.t227 XThC.XTB6.A XThC.XTB6.Y VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2327 VGND.t2094 XThC.XTB2.Y XThC.Tn[1].t9 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 XA.XIR[10].XIC[13].icell.PUM XThC.Tn[13].t38 XA.XIR[10].XIC[13].icell.Ien VPWR.t541 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2329 XA.XIR[2].XIC[6].icell.SM XA.XIR[2].XIC[6].icell.Ien Iout.t29 VGND.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2330 VGND.t2250 Vbias.t214 XA.XIR[12].XIC[12].icell.SM VGND.t2249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2331 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t62 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2332 XThC.Tn[6].t4 XThC.XTBN.Y.t97 a_6243_9615# VPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2333 XA.XIR[6].XIC[14].icell.SM XA.XIR[6].XIC[14].icell.Ien Iout.t178 VGND.t1374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2334 VGND.t2252 Vbias.t215 XA.XIR[15].XIC[13].icell.SM VGND.t2251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2335 VGND.t2254 Vbias.t216 XA.XIR[14].XIC[14].icell.SM VGND.t2253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2336 VGND.t745 XThC.Tn[12].t37 XA.XIR[15].XIC[12].icell.PDM VGND.t744 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2337 VGND.t1406 XThC.Tn[4].t39 XA.XIR[11].XIC[4].icell.PDM VGND.t1405 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2338 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[2].t59 XA.XIR[2].XIC[2].icell.Ien VGND.t525 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2339 VPWR.t1365 XThR.XTB7.Y a_n1049_5317# VPWR.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2340 VPWR.t1237 XThR.Tn[9].t61 XA.XIR[10].XIC[1].icell.PUM VPWR.t1236 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2341 VGND.t2665 VPWR.t2042 XA.XIR[6].XIC_dummy_right.icell.PDM VGND.t2664 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2342 VPWR.t1407 XThC.XTB6.Y XThC.Tn[13].t4 VPWR.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2343 VPWR.t1574 XThR.Tn[11].t66 XA.XIR[12].XIC[3].icell.PUM VPWR.t1573 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2344 a_n997_3979# XThR.XTBN.Y VGND.t2318 VGND.t2317 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2345 XA.XIR[5].XIC[4].icell.Ien XThR.Tn[5].t60 VPWR.t1150 VPWR.t1149 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2346 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13].t62 VPWR.t762 VPWR.t761 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2347 XA.XIR[9].XIC[4].icell.Ien XThR.Tn[9].t62 VPWR.t1239 VPWR.t1238 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2348 XA.XIR[0].XIC[4].icell.SM XA.XIR[0].XIC[4].icell.Ien Iout.t244 VGND.t2533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2349 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t59 VPWR.t61 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2350 VGND.t2256 Vbias.t217 XA.XIR[5].XIC[3].icell.SM VGND.t2255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2351 VGND.t2258 Vbias.t218 XA.XIR[9].XIC[12].icell.SM VGND.t2257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2352 XA.XIR[9].XIC[7].icell.SM XA.XIR[9].XIC[7].icell.Ien Iout.t219 VGND.t1851 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2353 VGND.t245 XThR.XTB4.Y.t14 XThR.Tn[3].t0 VGND.t244 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2354 XA.XIR[5].XIC[10].icell.SM XA.XIR[5].XIC[10].icell.Ien Iout.t154 VGND.t1144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2355 a_7331_10587# data[0].t2 VPWR.t1070 VPWR.t1069 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2356 a_4067_9615# XThC.XTBN.Y.t98 XThC.Tn[2].t3 VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2357 VPWR.t1451 XThR.Tn[2].t60 XA.XIR[3].XIC[12].icell.PUM VPWR.t1450 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2358 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[12].t64 VGND.t1993 VGND.t1992 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2359 XA.XIR[12].XIC[8].icell.SM XA.XIR[12].XIC[8].icell.Ien Iout.t24 VGND.t181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2360 XA.XIR[11].XIC[14].icell.Ien XThR.Tn[11].t67 VPWR.t1576 VPWR.t1575 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2361 VGND.t1676 Vbias.t219 XA.XIR[8].XIC[4].icell.SM VGND.t1675 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2362 VGND.t971 VGND.t969 XA.XIR[3].XIC_dummy_right.icell.SM VGND.t970 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2363 XA.XIR[7].XIC[5].icell.Ien XThR.Tn[7].t57 VPWR.t868 VPWR.t867 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2364 VPWR.t479 XThR.Tn[6].t63 XA.XIR[7].XIC[12].icell.PUM VPWR.t478 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2365 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13].t63 XA.XIR[13].XIC[4].icell.Ien VGND.t361 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2366 XA.XIR[15].XIC[9].icell.SM XA.XIR[15].XIC[9].icell.Ien Iout.t31 VGND.t213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2367 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t2043 XA.XIR[8].XIC_dummy_right.icell.Ien VGND.t2666 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2368 VPWR.t1152 XThR.Tn[5].t61 XA.XIR[6].XIC[13].icell.PUM VPWR.t1151 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2369 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t1 VPWR.t1765 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2370 XA.XIR[0].XIC[11].icell.PDM VGND.t966 VGND.t968 VGND.t967 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2371 XA.XIR[3].XIC[0].icell.PUM XThC.Tn[0].t36 XA.XIR[3].XIC[0].icell.Ien VPWR.t1885 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2372 XA.XIR[1].XIC_15.icell.PDM VPWR.t2044 VGND.t2668 VGND.t2667 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2373 XA.XIR[5].XIC[1].icell.SM XA.XIR[5].XIC[1].icell.Ien Iout.t119 VGND.t843 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2374 XA.XIR[2].XIC[10].icell.SM XA.XIR[2].XIC[10].icell.Ien Iout.t30 VGND.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2375 XThC.Tn[3].t4 XThC.XTBN.Y.t99 a_4861_9615# VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2376 XA.XIR[3].XIC[14].icell.SM XA.XIR[3].XIC[14].icell.Ien Iout.t118 VGND.t842 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2377 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t57 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t58 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2378 XThC.XTB5.A data[0].t3 VGND.t906 VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2379 VGND.t402 XThC.Tn[10].t38 XA.XIR[15].XIC[10].icell.PDM VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2380 VPWR.t575 XThR.XTB4.Y.t15 XThR.Tn[11].t1 VPWR.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2381 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[2].t61 XA.XIR[2].XIC[6].icell.Ien VGND.t552 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2382 XA.XIR[0].XIC[2].icell.PDM VGND.t963 VGND.t965 VGND.t964 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2383 XA.XIR[2].XIC[1].icell.SM XA.XIR[2].XIC[1].icell.Ien Iout.t70 VGND.t450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2384 VGND.t1569 XThC.Tn[11].t36 XA.XIR[2].XIC[11].icell.PDM VGND.t1568 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2385 VGND.t2316 XThR.XTBN.Y a_n997_715# VGND.t2315 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2386 a_n997_2891# XThR.XTBN.Y VGND.t2314 VGND.t2313 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2387 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[7].t58 VGND.t641 VGND.t640 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2388 VGND.t962 VGND.t960 XA.XIR[6].XIC_dummy_left.icell.SM VGND.t961 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2389 XA.XIR[5].XIC[0].icell.Ien XThR.Tn[5].t62 VPWR.t1154 VPWR.t1153 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2390 VPWR.t1511 XThR.Tn[3].t66 XA.XIR[4].XIC[9].icell.PUM VPWR.t1510 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2391 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9].t63 VPWR.t1241 VPWR.t1240 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2392 VPWR.t1449 XThR.Tn[2].t62 XA.XIR[3].XIC[10].icell.PUM VPWR.t1448 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2393 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t54 VPWR.t56 VPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2394 VPWR.t481 XThR.Tn[6].t64 XA.XIR[7].XIC[10].icell.PUM VPWR.t480 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2395 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14].t65 XA.XIR[14].XIC[1].icell.Ien VGND.t2429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2396 XA.XIR[10].XIC[6].icell.PUM XThC.Tn[6].t38 XA.XIR[10].XIC[6].icell.Ien VPWR.t696 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2397 XThR.Tn[11].t2 XThR.XTB4.Y.t16 a_n997_2667# VGND.t246 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2398 VPWR.t53 VPWR.t51 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t52 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2399 VGND.t1796 XThC.Tn[2].t36 XA.XIR[2].XIC[2].icell.PDM VGND.t1795 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2400 XA.XIR[13].XIC[7].icell.PUM XThC.Tn[7].t34 XA.XIR[13].XIC[7].icell.Ien VPWR.t1688 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2401 XA.XIR[9].XIC[2].icell.SM XA.XIR[9].XIC[2].icell.Ien Iout.t174 VGND.t1357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2402 VPWR.t1735 XThC.XTB2.Y XThC.Tn[9].t4 VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2403 XA.XIR[3].XIC[12].icell.Ien XThR.Tn[3].t67 VPWR.t1513 VPWR.t1512 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2404 a_n997_3979# XThR.XTB1.Y.t15 XThR.Tn[8].t1 VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2405 VGND.t2670 VPWR.t2045 XA.XIR[0].XIC_15.icell.PDM VGND.t2669 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2406 VGND.t1709 XThC.Tn[9].t40 XA.XIR[10].XIC[9].icell.PDM VGND.t1708 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2407 XA.XIR[12].XIC[3].icell.SM XA.XIR[12].XIC[3].icell.Ien Iout.t23 VGND.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2408 VPWR.t639 XThC.XTBN.Y.t100 XThC.Tn[8].t0 VPWR.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2409 XA.XIR[15].XIC[4].icell.SM XA.XIR[15].XIC[4].icell.Ien Iout.t227 VGND.t2097 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2410 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[4].t64 XA.XIR[4].XIC[8].icell.Ien VGND.t1752 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2411 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[4].t65 XA.XIR[4].XIC[14].icell.Ien VGND.t1753 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2412 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout VGND.t563 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2413 a_n1335_8331# XThR.XTB5.A XThR.XTB1.Y.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2414 VPWR.t1845 XThR.Tn[14].t66 XA.XIR[15].XIC[8].icell.PUM VPWR.t1844 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2415 XA.XIR[0].XIC[6].icell.PDM VGND.t957 VGND.t959 VGND.t958 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2416 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11].t68 XA.XIR[11].XIC[12].icell.Ien VGND.t1614 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2417 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t4 VPWR.t1765 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2418 XA.XIR[15].XIC[7].icell.Ien VPWR.t48 VPWR.t50 VPWR.t49 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2419 XThR.Tn[7].t0 XThR.XTBN.Y VPWR.t1764 VPWR.t1763 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2420 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2046 VGND.t2672 VGND.t2671 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2421 VPWR.t1156 XThR.Tn[5].t63 XA.XIR[6].XIC[6].icell.PUM VPWR.t1155 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2422 VGND.t956 VGND.t954 XA.XIR[3].XIC_dummy_left.icell.SM VGND.t955 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2423 VPWR.t545 XThR.Tn[8].t64 XA.XIR[9].XIC[7].icell.PUM VPWR.t544 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2424 XThC.Tn[9].t0 XThC.XTBN.Y.t101 VPWR.t641 VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2425 XThR.Tn[1].t9 XThR.XTBN.Y VGND.t2312 VGND.t2311 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2426 VPWR.t34 VPWR.t32 XA.XIR[13].XIC_15.icell.PUM VPWR.t33 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2427 VGND.t1678 Vbias.t220 XA.XIR[2].XIC[7].icell.SM VGND.t1677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2428 VGND.t378 XThC.Tn[6].t39 XA.XIR[2].XIC[6].icell.PDM VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2429 XA.XIR[13].XIC[11].icell.PUM XThC.Tn[11].t37 XA.XIR[13].XIC[11].icell.Ien VPWR.t1527 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2430 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[11].t69 VGND.t1616 VGND.t1615 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2431 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[7].t59 VGND.t643 VGND.t642 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2432 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2047 VGND.t2105 VGND.t2104 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2433 XA.XIR[4].XIC[9].icell.Ien XThR.Tn[4].t66 VPWR.t1628 VPWR.t1627 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2434 XA.XIR[3].XIC[10].icell.Ien XThR.Tn[3].t68 VPWR.t993 VPWR.t992 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2435 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[10].t62 VGND.t1745 VGND.t1744 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2436 XA.XIR[14].XIC[11].icell.SM XA.XIR[14].XIC[11].icell.Ien Iout.t220 VGND.t1979 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2437 XA.XIR[15].XIC[13].icell.PDM XThR.Tn[14].t67 VGND.t2431 VGND.t2430 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2438 VPWR.t643 XThC.XTBN.Y.t102 XThC.Tn[11].t2 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2439 VPWR.t1447 XThR.Tn[2].t63 XA.XIR[3].XIC[5].icell.PUM VPWR.t1446 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2440 VPWR.t1092 XThR.XTB6.Y a_n1049_5611# VPWR.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2441 VGND.t2107 VPWR.t2048 XA.XIR[15].XIC_dummy_left.icell.PDM VGND.t2106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2442 a_n997_2891# XThR.XTB3.Y.t15 XThR.Tn[10].t7 VGND.t1848 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2443 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[1].t59 XA.XIR[1].XIC[11].icell.Ien VGND.t590 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2444 XA.XIR[13].XIC[12].icell.SM XA.XIR[13].XIC[12].icell.Ien Iout.t58 VGND.t355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2445 VPWR.t483 XThR.Tn[6].t65 XA.XIR[7].XIC[5].icell.PUM VPWR.t482 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2446 XA.XIR[10].XIC[1].icell.PUM XThC.Tn[1].t40 XA.XIR[10].XIC[1].icell.Ien VPWR.t920 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2447 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t46 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t47 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2448 XA.XIR[1].XIC[6].icell.SM XA.XIR[1].XIC[6].icell.Ien Iout.t187 VGND.t1456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2449 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[1].t60 VGND.t592 VGND.t591 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2450 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[1].t61 VGND.t594 VGND.t593 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2451 XA.XIR[13].XIC[2].icell.PUM XThC.Tn[2].t37 XA.XIR[13].XIC[2].icell.Ien VPWR.t1652 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2452 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11].t70 XA.XIR[11].XIC[10].icell.Ien VGND.t1617 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2453 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[8].t65 VGND.t209 VGND.t208 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2454 XA.XIR[8].XIC[14].icell.PUM XThC.Tn[14].t39 XA.XIR[8].XIC[14].icell.Ien VPWR.t593 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2455 VGND.t1680 Vbias.t221 XA.XIR[10].XIC[5].icell.SM VGND.t1679 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2456 XA.XIR[15].XIC[11].icell.Ien VPWR.t43 VPWR.t45 VPWR.t44 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2457 VGND.t1408 XThC.Tn[4].t40 XA.XIR[10].XIC[4].icell.PDM VGND.t1407 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2458 VGND.t2109 VPWR.t2049 XA.XIR[5].XIC_dummy_right.icell.PDM VGND.t2108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2459 XA.XIR[11].XIC_15.icell.PUM VPWR.t41 XA.XIR[11].XIC_15.icell.Ien VPWR.t42 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2460 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[1].t62 XA.XIR[1].XIC[2].icell.Ien VGND.t595 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2461 VGND.t1682 Vbias.t222 XA.XIR[13].XIC[6].icell.SM VGND.t1681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2462 XA.XIR[12].XIC[7].icell.Ien XThR.Tn[12].t65 VPWR.t1720 VPWR.t1719 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2463 VGND.t881 XThC.Tn[5].t36 XA.XIR[13].XIC[5].icell.PDM VGND.t880 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2464 VGND.t2111 VPWR.t2050 XA.XIR[9].XIC_dummy_right.icell.PDM VGND.t2110 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2465 XThC.Tn[2].t2 XThC.XTBN.Y.t103 a_4067_9615# VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2466 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[4].t67 XA.XIR[4].XIC[3].icell.Ien VGND.t1303 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2467 VPWR.t547 XThR.Tn[8].t66 XA.XIR[9].XIC[11].icell.PUM VPWR.t546 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2468 VPWR.t1847 XThR.Tn[14].t68 XA.XIR[15].XIC[3].icell.PUM VPWR.t1846 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2469 XA.XIR[7].XIC[12].icell.PUM XThC.Tn[12].t38 XA.XIR[7].XIC[12].icell.Ien VPWR.t966 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2470 VGND.t2284 XThR.XTB7.B XThR.XTB4.Y.t1 VGND.t2283 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2471 VPWR.t40 VPWR.t38 XA.XIR[10].XIC_15.icell.PUM VPWR.t39 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2472 VGND.t1684 Vbias.t223 XA.XIR[4].XIC_15.icell.SM VGND.t1683 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2473 XA.XIR[15].XIC[2].icell.Ien VPWR.t35 VPWR.t37 VPWR.t36 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2474 VGND.t1686 Vbias.t224 XA.XIR[11].XIC[13].icell.SM VGND.t1685 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2475 XA.XIR[10].XIC[14].icell.Ien XThR.Tn[10].t63 VPWR.t1618 VPWR.t1617 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2476 VGND.t360 XThR.XTB1.Y.t16 XThR.Tn[0].t1 VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2477 VPWR.t1675 XThR.Tn[1].t63 XA.XIR[2].XIC[4].icell.PUM VPWR.t1674 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2478 VPWR.t1135 XThR.Tn[5].t64 XA.XIR[6].XIC[1].icell.PUM VPWR.t1134 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2479 XA.XIR[13].XIC_15.icell.Ien XThR.Tn[13].t64 VPWR.t686 VPWR.t685 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2480 XA.XIR[14].XIC[9].icell.SM XA.XIR[14].XIC[9].icell.Ien Iout.t195 VGND.t1548 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2481 VPWR.t549 XThR.Tn[8].t67 XA.XIR[9].XIC[2].icell.PUM VPWR.t548 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2482 XA.XIR[15].XIC[5].icell.PDM VPWR.t2051 XA.XIR[15].XIC[5].icell.Ien VGND.t2112 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2483 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout VGND.t885 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2484 VGND.t1571 XThC.Tn[11].t38 XA.XIR[14].XIC[11].icell.PDM VGND.t1570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2485 VGND.t1688 Vbias.t225 XA.XIR[2].XIC[2].icell.SM VGND.t1687 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2486 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t29 VPWR.t31 VPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2487 XA.XIR[1].XIC[10].icell.SM XA.XIR[1].XIC[10].icell.Ien Iout.t237 VGND.t2403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2488 a_8739_9569# XThC.XTBN.Y.t104 VGND.t407 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2489 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[8].t68 VGND.t211 VGND.t210 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2490 XThC.Tn[6].t8 XThC.XTB7.Y VGND.t1167 VGND.t1166 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2491 XA.XIR[3].XIC[5].icell.Ien XThR.Tn[3].t69 VPWR.t995 VPWR.t994 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2492 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[10].t64 VGND.t1747 VGND.t1746 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2493 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[5].t65 VGND.t1082 VGND.t1081 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2494 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[1].t64 XA.XIR[1].XIC[6].icell.Ien VGND.t1831 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2495 VGND.t1690 Vbias.t226 XA.XIR[13].XIC[10].icell.SM VGND.t1689 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2496 VGND.t409 XThC.XTBN.Y.t105 XThC.Tn[7].t4 VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2497 XThC.Tn[12].t8 XThC.XTBN.Y.t106 VPWR.t708 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2498 XA.XIR[12].XIC[11].icell.Ien XThR.Tn[12].t66 VPWR.t1722 VPWR.t1721 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2499 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[4].t68 XA.XIR[4].XIC[7].icell.Ien VGND.t1304 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2500 VGND.t1798 XThC.Tn[2].t38 XA.XIR[14].XIC[2].icell.PDM VGND.t1797 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2501 XThC.Tn[12].t4 XThC.XTB5.Y a_9827_9569# VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2502 XA.XIR[1].XIC[1].icell.SM XA.XIR[1].XIC[1].icell.Ien Iout.t141 VGND.t932 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2503 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[1].t65 VGND.t1833 VGND.t1832 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2504 XA.XIR[7].XIC[10].icell.PUM XThC.Tn[10].t39 XA.XIR[7].XIC[10].icell.Ien VPWR.t705 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2505 XA.XIR[4].XIC[12].icell.PUM XThC.Tn[12].t39 XA.XIR[4].XIC[12].icell.Ien VPWR.t967 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2506 a_8963_9569# XThC.XTB4.Y.t15 XThC.Tn[11].t7 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2507 XA.XIR[0].XIC[13].icell.SM XA.XIR[0].XIC[13].icell.Ien Iout.t134 VGND.t925 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2508 XA.XIR[3].XIC[13].icell.PUM XThC.Tn[13].t39 XA.XIR[3].XIC[13].icell.Ien VPWR.t542 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2509 VGND.t1692 Vbias.t227 XA.XIR[10].XIC[0].icell.SM VGND.t1691 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2510 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t27 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2511 VGND.t1694 Vbias.t228 XA.XIR[5].XIC[12].icell.SM VGND.t1693 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2512 VGND.t2402 XThC.Tn[8].t40 XA.XIR[1].XIC[8].icell.PDM VGND.t2401 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2513 VGND.t274 XThC.Tn[14].t40 XA.XIR[1].XIC[14].icell.PDM VGND.t273 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2514 XThR.Tn[13].t1 XThR.XTB6.Y VPWR.t1090 VPWR.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2515 VGND.t1696 Vbias.t229 XA.XIR[13].XIC[1].icell.SM VGND.t1695 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2516 XA.XIR[12].XIC[2].icell.Ien XThR.Tn[12].t67 VPWR.t1724 VPWR.t1723 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2517 VGND.t2572 XThC.Tn[0].t37 XA.XIR[13].XIC[0].icell.PDM VGND.t2571 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2518 VGND.t1698 Vbias.t230 XA.XIR[8].XIC[13].icell.SM VGND.t1697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2519 XA.XIR[7].XIC[14].icell.Ien XThR.Tn[7].t60 VPWR.t870 VPWR.t869 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2520 VGND.t747 XThC.Tn[12].t40 XA.XIR[8].XIC[12].icell.PDM VGND.t746 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2521 VPWR.t1677 XThR.Tn[1].t66 XA.XIR[2].XIC[0].icell.PUM VPWR.t1676 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2522 VGND.t200 XThC.Tn[13].t40 XA.XIR[11].XIC[13].icell.PDM VGND.t199 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2523 XA.XIR[12].XIC[7].icell.PUM XThC.Tn[7].t35 XA.XIR[12].XIC[7].icell.Ien VPWR.t1689 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2524 VGND.t411 XThC.XTBN.Y.t107 a_7875_9569# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2525 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12].t68 XA.XIR[12].XIC[5].icell.Ien VGND.t1994 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2526 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2052 XA.XIR[11].XIC_dummy_left.icell.Ien VGND.t2113 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2527 XA.XIR[15].XIC[8].icell.PUM XThC.Tn[8].t41 XA.XIR[15].XIC[8].icell.Ien VPWR.t1822 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2528 XA.XIR[2].XIC[4].icell.Ien XThR.Tn[2].t64 VPWR.t1445 VPWR.t1444 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2529 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14].t69 XA.XIR[14].XIC_15.icell.Ien VGND.t2432 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2530 XA.XIR[11].XIC_15.icell.SM XA.XIR[11].XIC_15.icell.Ien Iout.t39 VGND.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2531 VGND.t2003 Vbias.t231 XA.XIR[7].XIC[11].icell.SM VGND.t2002 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2532 XA.XIR[6].XIC[12].icell.Ien XThR.Tn[6].t66 VPWR.t485 VPWR.t484 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2533 XA.XIR[5].XIC[13].icell.Ien XThR.Tn[5].t66 VPWR.t1137 VPWR.t1136 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2534 XA.XIR[14].XIC[4].icell.SM XA.XIR[14].XIC[4].icell.Ien Iout.t196 VGND.t1549 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2535 XA.XIR[9].XIC[13].icell.Ien XThR.Tn[9].t64 VPWR.t1243 VPWR.t1242 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2536 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[5].t67 VGND.t1084 VGND.t1083 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2537 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout VGND.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2538 VPWR.t1110 VGND.t2700 XA.XIR[0].XIC[12].icell.PUM VPWR.t1109 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2539 XA.XIR[15].XIC[0].icell.PDM VPWR.t2053 XA.XIR[15].XIC[0].icell.Ien VGND.t2114 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2540 a_8963_9569# XThC.XTBN.Y.t108 VGND.t412 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2541 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10].t65 XA.XIR[10].XIC[12].icell.Ien VGND.t1748 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2542 VGND.t380 XThC.Tn[6].t40 XA.XIR[14].XIC[6].icell.PDM VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2543 XA.XIR[1].XIC[9].icell.PUM XThC.Tn[9].t41 XA.XIR[1].XIC[9].icell.Ien VPWR.t1604 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2544 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[1].t67 VGND.t1835 VGND.t1834 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2545 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13].t65 XA.XIR[13].XIC[13].icell.Ien VGND.t362 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2546 VPWR.t26 VPWR.t24 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t25 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2547 XA.XIR[4].XIC[10].icell.PUM XThC.Tn[10].t40 XA.XIR[4].XIC[10].icell.Ien VPWR.t706 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2548 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[13].t66 VGND.t364 VGND.t363 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2549 XA.XIR[0].XIC[8].icell.PDM XThR.Tn[0].t66 XA.XIR[0].XIC[8].icell.Ien VGND.t834 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2550 XA.XIR[0].XIC[14].icell.PDM XThR.Tn[0].t67 XA.XIR[0].XIC[14].icell.Ien VGND.t835 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2551 VPWR.t872 XThR.Tn[7].t61 XA.XIR[8].XIC[7].icell.PUM VPWR.t871 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2552 VGND.t404 XThC.Tn[10].t41 XA.XIR[8].XIC[10].icell.PDM VGND.t403 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2553 XThC.Tn[11].t1 XThC.XTBN.Y.t109 VPWR.t709 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2554 VPWR.t1620 XThR.Tn[10].t66 XA.XIR[11].XIC[8].icell.PUM VPWR.t1619 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2555 VGND.t2005 Vbias.t232 XA.XIR[1].XIC[7].icell.SM VGND.t2004 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2556 XThR.Tn[6].t5 XThR.XTBN.Y a_n1049_5317# VPWR.t1760 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2557 XA.XIR[7].XIC[5].icell.PUM XThC.Tn[5].t37 XA.XIR[7].XIC[5].icell.Ien VPWR.t1056 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2558 VPWR.t1288 XThC.XTB4.Y.t16 XThC.Tn[11].t4 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2559 XThR.XTB7.Y XThR.XTB7.B a_n1319_5317# VPWR.t1746 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2560 XA.XIR[12].XIC[11].icell.PUM XThC.Tn[11].t39 XA.XIR[12].XIC[11].icell.Ien VPWR.t1528 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2561 VGND.t2007 Vbias.t233 XA.XIR[4].XIC[8].icell.SM VGND.t2006 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2562 XA.XIR[15].XIC[1].icell.PDM XThR.Tn[14].t70 VGND.t2434 VGND.t2433 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2563 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[13].t67 VGND.t366 VGND.t365 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2564 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[9].t65 VGND.t1214 VGND.t1213 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2565 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2054 VGND.t2116 VGND.t2115 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2566 VGND.t2090 XThC.Tn[3].t41 XA.XIR[1].XIC[3].icell.PDM VGND.t2089 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2567 VGND.t2009 Vbias.t234 XA.XIR[7].XIC[9].icell.SM VGND.t2008 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2568 XA.XIR[6].XIC[10].icell.Ien XThR.Tn[6].t67 VPWR.t487 VPWR.t486 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2569 XA.XIR[2].XIC[0].icell.Ien XThR.Tn[2].t65 VPWR.t1443 VPWR.t1442 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2570 XA.XIR[12].XIC_15.icell.PDM VPWR.t2055 VGND.t2118 VGND.t2117 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2571 XA.XIR[12].XIC[12].icell.SM XA.XIR[12].XIC[12].icell.Ien Iout.t69 VGND.t449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2572 XA.XIR[8].XIC_15.icell.SM XA.XIR[8].XIC_15.icell.Ien Iout.t133 VGND.t910 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2573 XA.XIR[15].XIC[13].icell.SM XA.XIR[15].XIC[13].icell.Ien Iout.t200 VGND.t1579 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2574 VPWR.t1108 VGND.t2701 XA.XIR[0].XIC[10].icell.PUM VPWR.t1107 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2575 VPWR.t1060 XThC.XTB3.Y.t14 a_4067_9615# VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2576 XA.XIR[3].XIC[6].icell.PUM XThC.Tn[6].t41 XA.XIR[3].XIC[6].icell.Ien VPWR.t697 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2577 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12].t69 XA.XIR[12].XIC[0].icell.Ien VGND.t1995 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2578 XA.XIR[12].XIC[2].icell.PUM XThC.Tn[2].t39 XA.XIR[12].XIC[2].icell.Ien VPWR.t1653 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2579 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10].t67 XA.XIR[10].XIC[10].icell.Ien VGND.t1749 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2580 VGND.t2310 XThR.XTBN.Y a_n997_1803# VGND.t2309 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2581 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7].t62 XA.XIR[7].XIC[12].icell.Ien VGND.t644 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2582 XA.XIR[0].XIC[9].icell.Ien XThR.Tn[0].t68 VPWR.t823 VPWR.t822 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2583 XA.XIR[15].XIC[3].icell.PUM XThC.Tn[3].t42 XA.XIR[15].XIC[3].icell.Ien VPWR.t1732 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2584 XA.XIR[6].XIC[7].icell.PUM XThC.Tn[7].t36 XA.XIR[6].XIC[7].icell.Ien VPWR.t1690 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2585 XA.XIR[10].XIC_15.icell.PUM VPWR.t22 XA.XIR[10].XIC_15.icell.Ien VPWR.t23 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2586 a_3773_9615# XThC.XTB2.Y VPWR.t1734 VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2587 VPWR.t21 VPWR.t19 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2588 VGND.t2011 Vbias.t235 XA.XIR[12].XIC[6].icell.SM VGND.t2010 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2589 VGND.t1711 XThC.Tn[9].t42 XA.XIR[3].XIC[9].icell.PDM VGND.t1710 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2590 VGND.t1228 XThC.Tn[5].t38 XA.XIR[12].XIC[5].icell.PDM VGND.t1227 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2591 VPWR.t874 XThR.Tn[7].t63 XA.XIR[8].XIC[11].icell.PUM VPWR.t873 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2592 XA.XIR[2].XIC[4].icell.PUM XThC.Tn[4].t41 XA.XIR[2].XIC[4].icell.Ien VPWR.t1377 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2593 VPWR.t577 XThR.XTB4.Y.t17 XThR.Tn[11].t3 VPWR.t576 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2594 a_n997_715# XThR.XTBN.Y VGND.t2308 VGND.t2307 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2595 VGND.t2013 Vbias.t236 XA.XIR[6].XIC[5].icell.SM VGND.t2012 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2596 VPWR.t684 XThR.XTB1.Y.t17 a_n1049_8581# VPWR.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2597 XA.XIR[4].XIC[5].icell.PUM XThC.Tn[5].t39 XA.XIR[4].XIC[5].icell.Ien VPWR.t1262 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2598 XA.XIR[5].XIC[6].icell.Ien XThR.Tn[5].t68 VPWR.t1139 VPWR.t1138 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2599 XThR.Tn[14].t1 XThR.XTB7.Y VPWR.t1364 VPWR.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2600 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[13].t68 VGND.t368 VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2601 XA.XIR[9].XIC[6].icell.Ien XThR.Tn[9].t66 VPWR.t1245 VPWR.t1244 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2602 VGND.t2015 Vbias.t237 XA.XIR[9].XIC[6].icell.SM VGND.t2014 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2603 VGND.t414 XThC.XTBN.Y.t110 XThC.Tn[3].t1 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2604 XA.XIR[8].XIC[7].icell.Ien XThR.Tn[8].t69 VPWR.t551 VPWR.t550 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2605 VGND.t1904 XThC.Tn[7].t37 XA.XIR[1].XIC[7].icell.PDM VGND.t1903 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2606 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2056 VGND.t2120 VGND.t2119 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2607 XA.XIR[0].XIC[3].icell.PDM XThR.Tn[0].t69 XA.XIR[0].XIC[3].icell.Ien VGND.t576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2608 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout VGND.t1417 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2609 VPWR.t659 XThR.Tn[7].t64 XA.XIR[8].XIC[2].icell.PUM VPWR.t658 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2610 XThC.Tn[1].t8 XThC.XTB2.Y VGND.t2093 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2611 VPWR.t1441 XThR.Tn[2].t66 XA.XIR[3].XIC[14].icell.PUM VPWR.t1440 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2612 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5].t69 XA.XIR[5].XIC[9].icell.Ien VGND.t1085 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2613 XA.XIR[11].XIC[8].icell.Ien XThR.Tn[11].t71 VPWR.t1566 VPWR.t1565 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2614 VPWR.t1728 XThC.XTBN.A XThC.XTBN.Y.t0 VPWR.t1727 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2615 VPWR.t1606 XThR.Tn[10].t68 XA.XIR[11].XIC[3].icell.PUM VPWR.t1605 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2616 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9].t67 XA.XIR[9].XIC[9].icell.Ien VGND.t1215 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2617 VPWR.t489 XThR.Tn[6].t68 XA.XIR[7].XIC[14].icell.PUM VPWR.t488 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2618 VGND.t2017 Vbias.t238 XA.XIR[1].XIC[2].icell.SM VGND.t2016 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2619 VPWR.t18 VPWR.t16 XA.XIR[6].XIC_15.icell.PUM VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2620 VGND.t2019 Vbias.t239 XA.XIR[4].XIC[3].icell.SM VGND.t2018 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2621 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7].t65 XA.XIR[7].XIC[10].icell.Ien VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2622 XThR.Tn[2].t3 XThR.XTB3.Y.t16 VGND.t1201 VGND.t1200 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2623 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[9].t68 VGND.t1217 VGND.t1216 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2624 XA.XIR[6].XIC[11].icell.PUM XThC.Tn[11].t40 XA.XIR[6].XIC[11].icell.Ien VPWR.t1529 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2625 XA.XIR[11].XIC[8].icell.SM XA.XIR[11].XIC[8].icell.Ien Iout.t180 VGND.t1416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2626 VGND.t2021 Vbias.t240 XA.XIR[7].XIC[4].icell.SM VGND.t2020 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2627 XA.XIR[6].XIC[5].icell.Ien XThR.Tn[6].t69 VPWR.t491 VPWR.t490 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2628 VGND.t953 VGND.t951 XA.XIR[2].XIC_dummy_right.icell.SM VGND.t952 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2629 VGND.t2023 Vbias.t241 XA.XIR[12].XIC[10].icell.SM VGND.t2022 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2630 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[7].t66 VGND.t332 VGND.t331 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2631 a_n997_3979# XThR.XTB1.Y.t18 XThR.Tn[8].t2 VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2632 XA.XIR[7].XIC[11].icell.SM XA.XIR[7].XIC[11].icell.Ien Iout.t194 VGND.t1532 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2633 a_3299_10575# XThC.XTB7.B VGND.t1177 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2634 VGND.t2122 VPWR.t2057 XA.XIR[8].XIC_dummy_left.icell.PDM VGND.t2121 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2635 VGND.t2306 XThR.XTBN.Y XThR.Tn[6].t8 VGND.t2305 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2636 VPWR.t1106 VGND.t2702 XA.XIR[0].XIC[5].icell.PUM VPWR.t1105 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2637 XA.XIR[3].XIC[1].icell.PUM XThC.Tn[1].t41 XA.XIR[3].XIC[1].icell.Ien VPWR.t921 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2638 XA.XIR[2].XIC[0].icell.PUM XThC.Tn[0].t38 XA.XIR[2].XIC[0].icell.Ien VPWR.t1886 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2639 VPWR.t1568 XThR.Tn[11].t72 XA.XIR[12].XIC[9].icell.PUM VPWR.t1567 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2640 XA.XIR[6].XIC[2].icell.PUM XThC.Tn[2].t40 XA.XIR[6].XIC[2].icell.Ien VPWR.t1654 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2641 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t6 VPWR.t8 VPWR.t7 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2642 VGND.t2025 Vbias.t242 XA.XIR[12].XIC[1].icell.SM VGND.t2024 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2643 VGND.t1930 Vbias.t243 XA.XIR[3].XIC[5].icell.SM VGND.t1929 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2644 VGND.t2574 XThC.Tn[0].t39 XA.XIR[12].XIC[0].icell.PDM VGND.t2573 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2645 VGND.t1410 XThC.Tn[4].t42 XA.XIR[3].XIC[4].icell.PDM VGND.t1409 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2646 VGND.t1932 Vbias.t244 XA.XIR[9].XIC[10].icell.SM VGND.t1931 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2647 XA.XIR[8].XIC[11].icell.Ien XThR.Tn[8].t70 VPWR.t553 VPWR.t552 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2648 VGND.t703 XThC.Tn[1].t42 XA.XIR[11].XIC[1].icell.PDM VGND.t702 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2649 VGND.t1934 Vbias.t245 XA.XIR[10].XIC[14].icell.SM VGND.t1933 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2650 XA.XIR[0].XIC[7].icell.PDM XThR.Tn[0].t70 XA.XIR[0].XIC[7].icell.Ien VGND.t577 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2651 VGND.t1230 XThC.Tn[5].t40 XA.XIR[6].XIC[5].icell.PDM VGND.t1229 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2652 VPWR.t710 XThC.XTBN.Y.t111 XThC.Tn[10].t4 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2653 VGND.t202 XThC.Tn[13].t41 XA.XIR[10].XIC[13].icell.PDM VGND.t201 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2654 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2058 XA.XIR[10].XIC_dummy_left.icell.Ien VGND.t2123 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2655 XA.XIR[0].XIC[12].icell.PUM XThC.Tn[12].t41 XA.XIR[0].XIC[12].icell.Ien VPWR.t968 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2656 VGND.t415 XThC.XTBN.Y.t112 a_8963_9569# VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2657 XA.XIR[5].XIC[1].icell.Ien XThR.Tn[5].t70 VPWR.t1141 VPWR.t1140 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2658 VGND.t1936 Vbias.t246 XA.XIR[6].XIC[0].icell.SM VGND.t1935 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2659 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[6].t70 VGND.t135 VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2660 VPWR.t1413 XThC.XTB5.A a_5155_10571# VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2661 VPWR.t1205 XThC.XTB7.Y XThC.Tn[14].t4 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2662 XThR.Tn[1].t8 XThR.XTBN.Y VGND.t2304 VGND.t2303 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2663 XA.XIR[1].XIC[4].icell.Ien XThR.Tn[1].t68 VPWR.t1679 VPWR.t1678 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2664 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9].t69 VPWR.t1871 VPWR.t1870 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2665 VGND.t1938 Vbias.t247 XA.XIR[9].XIC[1].icell.SM VGND.t1937 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2666 XA.XIR[8].XIC[2].icell.Ien XThR.Tn[8].t71 VPWR.t700 VPWR.t699 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2667 XA.XIR[3].XIC[14].icell.Ien XThR.Tn[3].t70 VPWR.t997 VPWR.t996 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2668 XA.XIR[5].XIC[7].icell.SM XA.XIR[5].XIC[7].icell.Ien Iout.t177 VGND.t1373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2669 VPWR.t583 XThC.XTB7.A XThC.XTB3.Y.t0 VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2670 XA.XIR[11].XIC[3].icell.Ien XThR.Tn[11].t73 VPWR.t1570 VPWR.t1569 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2671 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5].t71 XA.XIR[5].XIC[4].icell.Ien VGND.t1086 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2672 XA.XIR[8].XIC[8].icell.SM XA.XIR[8].XIC[8].icell.Ien Iout.t115 VGND.t828 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2673 XA.XIR[7].XIC[9].icell.SM XA.XIR[7].XIC[9].icell.Ien Iout.t15 VGND.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2674 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13].t69 XA.XIR[13].XIC[1].icell.Ien VGND.t223 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2675 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9].t70 XA.XIR[9].XIC[4].icell.Ien VGND.t2541 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2676 XThR.Tn[8].t5 XThR.XTBN.Y VPWR.t1762 VPWR.t1761 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2677 VPWR.t1681 XThR.Tn[1].t69 XA.XIR[2].XIC[13].icell.PUM VPWR.t1680 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2678 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t2059 XA.XIR[4].XIC_dummy_right.icell.Ien VGND.t2124 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2679 XThR.Tn[5].t8 XThR.XTBN.Y a_n1049_5611# VPWR.t1760 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2680 a_n997_2891# XThR.XTB3.Y.t17 XThR.Tn[10].t2 VGND.t607 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2681 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8].t72 XA.XIR[8].XIC[5].icell.Ien VGND.t386 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2682 XThR.XTB6.Y XThR.XTB7.B a_n1319_5611# VPWR.t1746 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2683 VPWR.t11 VPWR.t9 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2684 XA.XIR[2].XIC[7].icell.SM XA.XIR[2].XIC[7].icell.Ien Iout.t192 VGND.t1503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2685 XA.XIR[11].XIC[3].icell.SM XA.XIR[11].XIC[3].icell.Ien Iout.t211 VGND.t1818 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2686 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t4 VPWR.t1759 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2687 a_3773_9615# XThC.XTBN.Y.t113 XThC.Tn[1].t1 VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2688 VPWR.t1745 XThR.XTB7.B XThR.XTB3.Y.t2 VPWR.t1744 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2689 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t2060 XA.XIR[7].XIC_dummy_left.icell.Ien VGND.t2125 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2690 XA.XIR[0].XIC[10].icell.PUM XThC.Tn[10].t42 XA.XIR[0].XIC[10].icell.Ien VPWR.t707 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2691 a_4067_9615# XThC.XTB3.Y.t15 VPWR.t1742 VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2692 VGND.t1940 Vbias.t248 XA.XIR[3].XIC[0].icell.SM VGND.t1939 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2693 VPWR.t1743 XThC.XTB3.Y.t16 XThC.Tn[10].t10 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2694 VPWR.t711 XThC.XTBN.Y.t114 XThC.Tn[14].t1 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2695 XA.XIR[1].XIC[0].icell.Ien XThR.Tn[1].t70 VPWR.t470 VPWR.t469 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2696 VGND.t950 VGND.t948 XA.XIR[2].XIC_dummy_left.icell.SM VGND.t949 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2697 XA.XIR[14].XIC[4].icell.PUM XThC.Tn[4].t43 XA.XIR[14].XIC[4].icell.Ien VPWR.t1378 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2698 XA.XIR[15].XIC_15.icell.PDM VPWR.t2061 VGND.t2127 VGND.t2126 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2699 XA.XIR[10].XIC[5].icell.SM XA.XIR[10].XIC[5].icell.Ien Iout.t225 VGND.t2091 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2700 VGND.t2576 XThC.Tn[0].t40 XA.XIR[6].XIC[0].icell.PDM VGND.t2575 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2701 XA.XIR[14].XIC[13].icell.SM XA.XIR[14].XIC[13].icell.Ien Iout.t63 VGND.t388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2702 VGND.t2302 XThR.XTBN.Y XThR.Tn[0].t6 VGND.t2301 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2703 XA.XIR[13].XIC[6].icell.SM XA.XIR[13].XIC[6].icell.Ien Iout.t162 VGND.t1250 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2704 VGND.t2103 XThC.XTB3.Y.t17 XThC.Tn[2].t11 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2705 XA.XIR[5].XIC[7].icell.PUM XThC.Tn[7].t38 XA.XIR[5].XIC[7].icell.Ien VPWR.t1691 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2706 XThR.Tn[10].t8 XThR.XTBN.Y VPWR.t1758 VPWR.t1757 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2707 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[6].t71 VGND.t137 VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2708 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2062 VGND.t2129 VGND.t2128 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2709 XA.XIR[9].XIC[7].icell.PUM XThC.Tn[7].t39 XA.XIR[9].XIC[7].icell.Ien VPWR.t1692 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2710 XA.XIR[5].XIC[2].icell.SM XA.XIR[5].XIC[2].icell.Ien Iout.t189 VGND.t1484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2711 XA.XIR[8].XIC[8].icell.PUM XThC.Tn[8].t42 XA.XIR[8].XIC[8].icell.Ien VPWR.t1823 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2712 VGND.t1942 Vbias.t249 XA.XIR[0].XIC[11].icell.SM VGND.t1941 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2713 VPWR.t1406 XThC.XTB6.Y a_5949_9615# VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2714 XThR.Tn[1].t0 XThR.XTB2.Y VGND.t97 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2715 XA.XIR[4].XIC_15.icell.SM XA.XIR[4].XIC_15.icell.Ien Iout.t205 VGND.t1593 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2716 VGND.t2300 XThR.XTBN.Y a_n997_3755# VGND.t2299 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2717 VPWR.t1071 data[3].t1 XThC.XTBN.A VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2718 XA.XIR[8].XIC[3].icell.SM XA.XIR[8].XIC[3].icell.Ien Iout.t231 VGND.t2101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2719 a_2979_9615# XThC.XTB1.Y.t17 VPWR.t617 VPWR.t616 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2720 XThC.Tn[3].t0 XThC.XTBN.Y.t115 VGND.t416 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2721 XA.XIR[2].XIC[13].icell.Ien XThR.Tn[2].t67 VPWR.t1439 VPWR.t1438 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2722 XA.XIR[7].XIC[4].icell.SM XA.XIR[7].XIC[4].icell.Ien Iout.t202 VGND.t1581 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2723 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8].t73 XA.XIR[8].XIC[0].icell.Ien VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2724 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[3].t71 XA.XIR[3].XIC[12].icell.Ien VGND.t784 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2725 XA.XIR[7].XIC[14].icell.PUM XThC.Tn[14].t41 XA.XIR[7].XIC[14].icell.Ien VPWR.t594 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2726 VPWR.t561 XThR.Tn[13].t70 XA.XIR[14].XIC[12].icell.PUM VPWR.t560 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2727 XA.XIR[2].XIC[2].icell.SM XA.XIR[2].XIC[2].icell.Ien Iout.t92 VGND.t687 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2728 XA.XIR[10].XIC[8].icell.Ien XThR.Tn[10].t69 VPWR.t1608 VPWR.t1607 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2729 a_5949_10571# XThC.XTB7.B XThC.XTB6.Y VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2730 VPWR.t472 XThR.Tn[1].t71 XA.XIR[2].XIC[6].icell.PUM VPWR.t471 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2731 VPWR.t825 XThR.Tn[0].t71 XA.XIR[1].XIC[7].icell.PUM VPWR.t824 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2732 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[10].t70 VGND.t1739 VGND.t1738 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2733 XA.XIR[14].XIC[0].icell.PUM XThC.Tn[0].t41 XA.XIR[14].XIC[0].icell.Ien VPWR.t1887 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2734 XThR.Tn[13].t0 XThR.XTB6.Y VPWR.t1088 VPWR.t1087 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2735 VPWR.t1330 XThR.Tn[4].t69 XA.XIR[5].XIC[7].icell.PUM VPWR.t1329 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2736 XA.XIR[13].XIC[10].icell.SM XA.XIR[13].XIC[10].icell.Ien Iout.t78 VGND.t561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2737 a_n1049_7493# XThR.XTB3.Y.t18 VPWR.t986 VPWR.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2738 XA.XIR[0].XIC[5].icell.PUM XThC.Tn[5].t41 XA.XIR[0].XIC[5].icell.Ien VPWR.t1263 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2739 XA.XIR[5].XIC[11].icell.PUM XThC.Tn[11].t41 XA.XIR[5].XIC[11].icell.Ien VPWR.t1530 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2740 XA.XIR[9].XIC[11].icell.PUM XThC.Tn[11].t42 XA.XIR[9].XIC[11].icell.Ien VPWR.t1531 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2741 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[7].t67 VGND.t334 VGND.t333 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2742 VGND.t947 VGND.t945 XA.XIR[1].XIC_dummy_right.icell.SM VGND.t946 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2743 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[2].t68 VGND.t554 VGND.t553 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2744 VGND.t1944 Vbias.t250 XA.XIR[0].XIC[9].icell.SM VGND.t1943 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2745 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[10].t71 VGND.t1741 VGND.t1740 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2746 XA.XIR[10].XIC[0].icell.SM XA.XIR[10].XIC[0].icell.Ien Iout.t246 VGND.t2535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2747 VPWR.t619 XThC.XTB1.Y.t18 XThC.Tn[8].t4 VPWR.t618 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2748 VGND.t1573 XThC.Tn[11].t43 XA.XIR[13].XIC[11].icell.PDM VGND.t1572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2749 XA.XIR[13].XIC[1].icell.SM XA.XIR[13].XIC[1].icell.Ien Iout.t209 VGND.t1806 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2750 VGND.t343 XThR.XTB5.Y XThR.Tn[4].t0 VGND.t342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2751 XThC.Tn[10].t8 XThC.XTBN.Y.t116 VPWR.t1398 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2752 VGND.t1447 XThC.XTBN.Y.t117 XThC.Tn[6].t0 VGND.t1446 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2753 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[3].t72 XA.XIR[3].XIC[10].icell.Ien VGND.t785 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2754 XA.XIR[5].XIC[2].icell.PUM XThC.Tn[2].t41 XA.XIR[5].XIC[2].icell.Ien VPWR.t1655 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2755 VPWR.t1849 XThR.Tn[14].t71 XA.XIR[15].XIC[9].icell.PUM VPWR.t1848 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2756 VPWR.t563 XThR.Tn[13].t71 XA.XIR[14].XIC[10].icell.PUM VPWR.t562 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2757 XA.XIR[9].XIC[2].icell.PUM XThC.Tn[2].t42 XA.XIR[9].XIC[2].icell.Ien VPWR.t1656 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2758 XA.XIR[4].XIC[14].icell.PUM XThC.Tn[14].t42 XA.XIR[4].XIC[14].icell.Ien VPWR.t940 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2759 XA.XIR[8].XIC[3].icell.PUM XThC.Tn[3].t43 XA.XIR[8].XIC[3].icell.Ien VPWR.t1733 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2760 XA.XIR[3].XIC_15.icell.PUM VPWR.t14 XA.XIR[3].XIC_15.icell.Ien VPWR.t15 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2761 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[4].t70 VGND.t1306 VGND.t1305 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2762 VGND.t1946 Vbias.t251 XA.XIR[5].XIC[6].icell.SM VGND.t1945 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2763 VGND.t705 XThC.Tn[1].t43 XA.XIR[10].XIC[1].icell.PDM VGND.t704 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2764 VGND.t2131 VPWR.t2063 XA.XIR[1].XIC_dummy_right.icell.PDM VGND.t2130 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2765 VGND.t1232 XThC.Tn[5].t42 XA.XIR[5].XIC[5].icell.PDM VGND.t1231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2766 VGND.t1800 XThC.Tn[2].t43 XA.XIR[13].XIC[2].icell.PDM VGND.t1799 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2767 VGND.t1234 XThC.Tn[5].t43 XA.XIR[9].XIC[5].icell.PDM VGND.t1233 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2768 VPWR.t827 XThR.Tn[0].t72 XA.XIR[1].XIC[11].icell.PUM VPWR.t826 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2769 XA.XIR[7].XIC[8].icell.Ien XThR.Tn[7].t68 VPWR.t661 VPWR.t660 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2770 VPWR.t1289 XThC.XTB4.Y.t17 a_4861_9615# VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2771 VPWR.t1332 XThR.Tn[4].t71 XA.XIR[5].XIC[11].icell.PUM VPWR.t1331 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2772 XA.XIR[14].XIC[12].icell.Ien XThR.Tn[14].t72 VPWR.t1851 VPWR.t1850 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2773 XA.XIR[15].XIC[11].icell.PDM VPWR.t2064 XA.XIR[15].XIC[11].icell.Ien VGND.t2132 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2774 VGND.t2134 VPWR.t2065 XA.XIR[11].XIC_15.icell.PDM VGND.t2133 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2775 XA.XIR[2].XIC[13].icell.PUM XThC.Tn[13].t42 XA.XIR[2].XIC[13].icell.Ien VPWR.t543 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2776 VGND.t1948 Vbias.t252 XA.XIR[4].XIC[12].icell.SM VGND.t1947 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2777 XThR.Tn[6].t4 XThR.XTBN.Y a_n1049_5317# VPWR.t1756 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2778 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t12 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t13 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2779 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t8 VGND.t1165 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2780 XA.XIR[2].XIC[6].icell.Ien XThR.Tn[2].t69 VPWR.t1437 VPWR.t1436 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2781 XA.XIR[10].XIC[3].icell.Ien XThR.Tn[10].t72 VPWR.t1610 VPWR.t1609 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2782 VGND.t1950 Vbias.t253 XA.XIR[7].XIC[13].icell.SM VGND.t1949 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2783 XA.XIR[6].XIC[14].icell.Ien XThR.Tn[6].t72 VPWR.t493 VPWR.t492 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2784 VGND.t1449 XThC.XTBN.Y.t118 a_10915_9569# VGND.t1448 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2785 VPWR.t474 XThR.Tn[1].t72 XA.XIR[2].XIC[1].icell.PUM VPWR.t473 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2786 XA.XIR[5].XIC_15.icell.Ien XThR.Tn[5].t72 VPWR.t1143 VPWR.t1142 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2787 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[10].t73 VGND.t1743 VGND.t1742 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2788 VGND.t749 XThC.Tn[12].t42 XA.XIR[7].XIC[12].icell.PDM VGND.t748 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2789 VGND.t1952 Vbias.t254 XA.XIR[6].XIC[14].icell.SM VGND.t1951 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2790 VPWR.t829 XThR.Tn[0].t73 XA.XIR[1].XIC[2].icell.PUM VPWR.t828 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2791 XA.XIR[9].XIC_15.icell.Ien XThR.Tn[9].t71 VPWR.t1873 VPWR.t1872 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2792 VPWR.t1334 XThR.Tn[4].t72 XA.XIR[5].XIC[2].icell.PUM VPWR.t1333 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2793 VPWR.t1104 VGND.t2703 XA.XIR[0].XIC[14].icell.PUM VPWR.t1103 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2794 XA.XIR[15].XIC[2].icell.PDM VPWR.t2066 XA.XIR[15].XIC[2].icell.Ien VGND.t2135 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2795 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[2].t70 XA.XIR[2].XIC[9].icell.Ien VGND.t152 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2796 XThC.Tn[1].t0 XThC.XTBN.Y.t119 a_3773_9615# VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2797 XA.XIR[1].XIC[7].icell.SM XA.XIR[1].XIC[7].icell.Ien Iout.t144 VGND.t1088 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2798 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13].t72 XA.XIR[13].XIC_15.icell.Ien VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2799 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[2].t71 VGND.t557 VGND.t556 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2800 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[4].t73 VGND.t1308 VGND.t1307 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2801 VGND.t2456 Vbias.t255 XA.XIR[0].XIC[4].icell.SM VGND.t2455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2802 XA.XIR[4].XIC[8].icell.SM XA.XIR[4].XIC[8].icell.Ien Iout.t222 VGND.t2001 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2803 XThC.Tn[14].t0 XThC.XTBN.Y.t120 VPWR.t1399 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2804 VGND.t2458 Vbias.t256 XA.XIR[5].XIC[10].icell.SM VGND.t2457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2805 VGND.t2460 Vbias.t257 XA.XIR[13].XIC[7].icell.SM VGND.t2459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2806 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2067 XA.XIR[0].XIC_dummy_right.icell.Ien VGND.t2136 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2807 VGND.t382 XThC.Tn[6].t42 XA.XIR[13].XIC[6].icell.PDM VGND.t381 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2808 VGND.t2298 XThR.XTBN.Y a_n997_715# VGND.t2297 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2809 VPWR.t5 VPWR.t3 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2810 XA.XIR[14].XIC[10].icell.Ien XThR.Tn[14].t73 VPWR.t1853 VPWR.t1852 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2811 VPWR.t565 XThR.Tn[13].t73 XA.XIR[14].XIC[5].icell.PUM VPWR.t564 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2812 VPWR.t1363 XThR.XTB7.Y XThR.Tn[14].t0 VPWR.t1095 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2813 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12].t70 XA.XIR[12].XIC[11].icell.Ien VGND.t1996 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2814 VGND.t944 VGND.t942 XA.XIR[1].XIC_dummy_left.icell.SM VGND.t943 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2815 VGND.t2462 Vbias.t258 XA.XIR[5].XIC[1].icell.SM VGND.t2461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2816 XA.XIR[9].XIC[5].icell.SM XA.XIR[9].XIC[5].icell.Ien Iout.t85 VGND.t656 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2817 XThR.XTB6.A data[5].t5 VGND.t807 VGND.t806 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2818 XThR.Tn[0].t2 XThR.XTBN.Y a_n1049_8581# VPWR.t1755 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2819 VGND.t1412 XThC.Tn[0].t42 XA.XIR[5].XIC[0].icell.PDM VGND.t1411 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2820 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[12].t71 VGND.t1998 VGND.t1997 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2821 a_5949_9615# XThC.XTB6.Y VPWR.t1405 VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2822 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[12].t72 VGND.t2000 VGND.t1999 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2823 XA.XIR[12].XIC[6].icell.SM XA.XIR[12].XIC[6].icell.Ien Iout.t167 VGND.t1270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2824 VGND.t1414 XThC.Tn[0].t43 XA.XIR[9].XIC[0].icell.PDM VGND.t1413 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2825 VGND.t406 XThC.Tn[10].t43 XA.XIR[7].XIC[10].icell.PDM VGND.t405 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2826 XA.XIR[7].XIC[3].icell.Ien XThR.Tn[7].t69 VPWR.t663 VPWR.t662 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2827 VGND.t1450 XThC.XTBN.Y.t121 a_10051_9569# VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2828 VGND.t2464 Vbias.t259 XA.XIR[3].XIC[14].icell.SM VGND.t2463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2829 VGND.t751 XThC.Tn[12].t43 XA.XIR[4].XIC[12].icell.PDM VGND.t750 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2830 VGND.t49 XThC.Tn[13].t43 XA.XIR[3].XIC[13].icell.PDM VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2831 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2068 XA.XIR[3].XIC_dummy_left.icell.Ien VGND.t2137 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2832 XA.XIR[15].XIC[6].icell.PDM VPWR.t2069 XA.XIR[15].XIC[6].icell.Ien VGND.t2138 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2833 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12].t73 XA.XIR[12].XIC[2].icell.Ien VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2834 XA.XIR[0].XIC[9].icell.PDM VGND.t939 VGND.t941 VGND.t940 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2835 VPWR.t1400 XThC.XTBN.Y.t122 XThC.Tn[11].t0 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2836 VGND.t1451 XThC.XTBN.Y.t123 a_7651_9569# VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2837 XA.XIR[2].XIC[1].icell.Ien XThR.Tn[2].t72 VPWR.t1435 VPWR.t1434 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2838 Vbias.t5 bias[1].t0 VPWR.t1404 VPWR.t1403 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
X2839 XA.XIR[11].XIC[12].icell.SM XA.XIR[11].XIC[12].icell.Ien Iout.t125 VGND.t887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2840 XA.XIR[1].XIC[13].icell.Ien XThR.Tn[1].t73 VPWR.t476 VPWR.t475 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2841 XThR.Tn[2].t4 XThR.XTBN.Y VGND.t2296 VGND.t2295 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2842 VPWR.t1362 XThR.XTB7.Y a_n1049_5317# VPWR.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2843 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout VGND.t1131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2844 VGND.t2466 Vbias.t260 XA.XIR[15].XIC_15.icell.SM VGND.t2465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2845 a_8739_9569# XThC.XTB3.Y.t18 XThC.Tn[10].t11 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2846 XA.XIR[2].XIC[6].icell.PUM XThC.Tn[6].t43 XA.XIR[2].XIC[6].icell.Ien VPWR.t698 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2847 VGND.t724 XThC.Tn[14].t43 XA.XIR[15].XIC[14].icell.PDM VGND.t723 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2848 VGND.t2530 XThC.Tn[8].t43 XA.XIR[15].XIC[8].icell.PDM VGND.t2529 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2849 VPWR.t1754 XThR.XTBN.Y XThR.Tn[12].t8 VPWR.t1753 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2850 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[2].t73 XA.XIR[2].XIC[4].icell.Ien VGND.t555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2851 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6].t73 XA.XIR[6].XIC[12].icell.Ien VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2852 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5].t73 XA.XIR[5].XIC[13].icell.Ien VGND.t1087 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2853 XA.XIR[1].XIC[2].icell.SM XA.XIR[1].XIC[2].icell.Ien Iout.t252 VGND.t2561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2854 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9].t72 XA.XIR[9].XIC[13].icell.Ien VGND.t2542 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2855 VPWR.t2 VPWR.t0 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2856 VGND.t1713 XThC.Tn[9].t43 XA.XIR[2].XIC[9].icell.PDM VGND.t1712 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2857 XA.XIR[4].XIC[3].icell.SM XA.XIR[4].XIC[3].icell.Ien Iout.t88 VGND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2858 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[9].t73 VGND.t2544 VGND.t2543 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2859 VGND.t2468 Vbias.t261 XA.XIR[13].XIC[2].icell.SM VGND.t2467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2860 VPWR.t999 XThR.Tn[3].t73 XA.XIR[4].XIC[7].icell.PUM VPWR.t998 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
R0 VGND.n3019 VGND.n3018 15660.6
R1 VGND.n196 VGND.n195 13477
R2 VGND.n3018 VGND.n7 11578
R3 VGND.n195 VGND.n7 10429.6
R4 VGND.n3012 VGND.n8 9309.26
R5 VGND.n200 VGND.n199 9223.7
R6 VGND.n198 VGND.n197 9223.7
R7 VGND.n197 VGND.n196 9223.7
R8 VGND.n2969 VGND.n200 9223.7
R9 VGND.n2969 VGND.n2968 7447.41
R10 VGND.n2249 VGND.n2248 7387.65
R11 VGND.n2250 VGND.n2249 7387.65
R12 VGND.n2285 VGND.n2284 7387.65
R13 VGND.n3017 VGND.n3016 7387.65
R14 VGND.n3016 VGND.n3015 7387.65
R15 VGND.n3015 VGND.n3014 7387.65
R16 VGND.n3014 VGND.n3013 7387.65
R17 VGND.n3013 VGND.n3012 7387.65
R18 VGND.n2351 VGND.n2285 6674.35
R19 VGND.n1386 VGND.t1846 6324.96
R20 VGND.n199 VGND.n198 5231.11
R21 VGND.n1336 VGND.t2613 5168.13
R22 VGND.n2967 VGND.n8 5074.71
R23 VGND.n3018 VGND.n3017 5063.19
R24 VGND.n1154 VGND.n806 4539.15
R25 VGND VGND.n8 4240.58
R26 VGND.t943 VGND.t686 4212.19
R27 VGND.t949 VGND.t240 4212.19
R28 VGND.t955 VGND.t639 4212.19
R29 VGND.t1042 VGND.t257 4212.19
R30 VGND.t1048 VGND.t840 4212.19
R31 VGND.t961 VGND.t357 4212.19
R32 VGND.t1003 VGND.t933 4212.19
R33 VGND.t247 VGND.t1054 4212.19
R34 VGND.t1417 VGND.t976 4212.19
R35 VGND.t885 VGND.t1021 4212.19
R36 VGND.t1504 VGND.t1060 4212.19
R37 VGND.t1340 VGND.t1072 4212.19
R38 VGND.t1111 VGND.t988 4212.19
R39 VGND.t1370 VGND.t1030 4212.19
R40 VGND.n2919 VGND.n222 4077.12
R41 VGND.n1340 VGND.n1338 3417.39
R42 VGND.n1340 VGND.n1339 3417.39
R43 VGND.n1388 VGND.n1387 3417.39
R44 VGND.n2180 VGND.n504 3417.39
R45 VGND.n503 VGND.n473 3417.39
R46 VGND.n2353 VGND.n2352 3417.39
R47 VGND.n2920 VGND.n2919 3331.79
R48 VGND.n2921 VGND.n2920 3331.79
R49 VGND.n2922 VGND.n2921 3331.79
R50 VGND.n2923 VGND.n2922 3331.79
R51 VGND.n2924 VGND.n2923 3331.79
R52 VGND.n2925 VGND.n2924 3331.79
R53 VGND.n2926 VGND.n2925 3331.79
R54 VGND.n2927 VGND.n2926 3331.79
R55 VGND.n2928 VGND.n2927 3331.79
R56 VGND.n2929 VGND.n2928 3331.79
R57 VGND.n2930 VGND.n2929 3331.79
R58 VGND.n2931 VGND.n2930 3331.79
R59 VGND.n2932 VGND.n2931 3331.79
R60 VGND.n2933 VGND.n2932 3331.79
R61 VGND.n2934 VGND.n2933 3331.79
R62 VGND.n1339 VGND.n806 3273.91
R63 VGND.n2181 VGND.n539 3265.22
R64 VGND.n2934 VGND.n201 2725.63
R65 VGND.n197 VGND.t2372 2655.17
R66 VGND.n196 VGND.t2348 2655.17
R67 VGND.n2353 VGND.n2285 2517.39
R68 VGND.t1850 VGND.n201 2334.15
R69 VGND.t2647 VGND.n2701 2307.69
R70 VGND.n359 VGND.t2227 2307.69
R71 VGND.n360 VGND.t2214 2307.69
R72 VGND.n370 VGND.t2137 2307.69
R73 VGND.n371 VGND.t2639 2307.69
R74 VGND.n381 VGND.t2201 2307.69
R75 VGND.n382 VGND.t1515 2307.69
R76 VGND.t2125 VGND.n327 2307.69
R77 VGND.n2705 VGND.t2609 2307.69
R78 VGND.n2728 VGND.t2202 2307.69
R79 VGND.n2738 VGND.t2123 2307.69
R80 VGND.t2113 VGND.n2737 2307.69
R81 VGND.n2731 VGND.t2600 2307.69
R82 VGND.n2776 VGND.t2171 2307.69
R83 VGND.t2148 VGND.n2775 2307.69
R84 VGND.n2943 VGND.t2597 2307.69
R85 VGND.t994 VGND.n2703 2280.49
R86 VGND.n3020 VGND.n5 2229.43
R87 VGND.n3020 VGND.n6 2229.43
R88 VGND.n2348 VGND.n6 2229.43
R89 VGND.n2348 VGND.n5 2229.43
R90 VGND.n1338 VGND.n1337 2173.91
R91 VGND.n2704 VGND.t148 2132.93
R92 VGND.n2701 VGND.t1518 2123.08
R93 VGND.t2641 VGND.n359 2123.08
R94 VGND.n360 VGND.t2619 2123.08
R95 VGND.t1516 VGND.n370 2123.08
R96 VGND.n371 VGND.t1505 2123.08
R97 VGND.t2119 VGND.n381 2123.08
R98 VGND.n382 VGND.t2203 2123.08
R99 VGND.n2705 VGND.t2115 2123.08
R100 VGND.t2603 VGND.n2728 2123.08
R101 VGND.n2738 VGND.t2591 2123.08
R102 VGND.n2737 VGND.t2151 2123.08
R103 VGND.n2731 VGND.t2671 2123.08
R104 VGND.n2776 VGND.t2579 2123.08
R105 VGND.n2775 VGND.t2165 2123.08
R106 VGND.n2704 VGND.t1018 2079.27
R107 VGND.t686 VGND.t994 2012.2
R108 VGND.t240 VGND.t943 2012.2
R109 VGND.t639 VGND.t949 2012.2
R110 VGND.t257 VGND.t955 2012.2
R111 VGND.t840 VGND.t1042 2012.2
R112 VGND.t357 VGND.t1048 2012.2
R113 VGND.t933 VGND.t961 2012.2
R114 VGND.t148 VGND.t1003 2012.2
R115 VGND.t1018 VGND.t247 2012.2
R116 VGND.t1054 VGND.t1417 2012.2
R117 VGND.t976 VGND.t885 2012.2
R118 VGND.t1021 VGND.t1504 2012.2
R119 VGND.t1060 VGND.t1340 2012.2
R120 VGND.t1072 VGND.t1111 2012.2
R121 VGND.t988 VGND.t1370 2012.2
R122 VGND.t1030 VGND.t1850 2012.2
R123 VGND.n199 VGND 1997.7
R124 VGND.n200 VGND 1997.7
R125 VGND VGND.n2969 1997.7
R126 VGND.n2968 VGND.n2944 1907.51
R127 VGND.n2284 VGND.n2251 1831.57
R128 VGND.n198 VGND.t2305 1807.04
R129 VGND.n2970 VGND.t1453 1785.51
R130 VGND.n2352 VGND.n2351 1760.87
R131 VGND.n2702 VGND.t2215 1738.46
R132 VGND.n2250 VGND.n504 1691.3
R133 VGND.n2351 VGND.n2350 1656.52
R134 VGND.t107 VGND.n66 1618.39
R135 VGND.n3011 VGND.t243 1618.39
R136 VGND.n2971 VGND.t347 1618.39
R137 VGND.n2702 VGND.n7 1604.17
R138 VGND.n2350 VGND.n328 1517.39
R139 VGND.n195 VGND.t2321 1517.24
R140 VGND.n2248 VGND.n540 1513.49
R141 VGND.t2180 VGND.n2704 1507.69
R142 VGND.n2703 VGND.n2702 1441.28
R143 VGND.n1386 VGND.n540 1370.36
R144 VGND.t2215 VGND.t1520 1353.85
R145 VGND.t1520 VGND.t2647 1353.85
R146 VGND.t2643 VGND.t1518 1353.85
R147 VGND.t2227 VGND.t2643 1353.85
R148 VGND.t2219 VGND.t2641 1353.85
R149 VGND.t2214 VGND.t2219 1353.85
R150 VGND.t2619 VGND.t2199 1353.85
R151 VGND.t2199 VGND.t2137 1353.85
R152 VGND.t1513 VGND.t1516 1353.85
R153 VGND.t2639 VGND.t1513 1353.85
R154 VGND.t1505 VGND.t2621 1353.85
R155 VGND.t2621 VGND.t2201 1353.85
R156 VGND.t2607 VGND.t2119 1353.85
R157 VGND.t1515 VGND.t2607 1353.85
R158 VGND.t2203 VGND.t1509 1353.85
R159 VGND.t1509 VGND.t2125 1353.85
R160 VGND.t2121 VGND.t2180 1353.85
R161 VGND.t2609 VGND.t2121 1353.85
R162 VGND.t2115 VGND.t2623 1353.85
R163 VGND.t2623 VGND.t2202 1353.85
R164 VGND.t2182 VGND.t2603 1353.85
R165 VGND.t2123 VGND.t2182 1353.85
R166 VGND.t2591 VGND.t2167 1353.85
R167 VGND.t2167 VGND.t2113 1353.85
R168 VGND.t2605 VGND.t2151 1353.85
R169 VGND.t2600 VGND.t2605 1353.85
R170 VGND.t2671 VGND.t2593 1353.85
R171 VGND.t2593 VGND.t2171 1353.85
R172 VGND.t2579 VGND.t2231 1353.85
R173 VGND.t2231 VGND.t2148 1353.85
R174 VGND.t2165 VGND.t2106 1353.85
R175 VGND.t2106 VGND.t2597 1353.85
R176 VGND.n2944 VGND.n201 1301.35
R177 VGND.n2703 VGND.n328 1278.26
R178 VGND.t940 VGND.n540 1270.28
R179 VGND.n1127 VGND.t632 1268.93
R180 VGND.n1127 VGND.t141 1268.93
R181 VGND.n502 VGND.t45 1253.59
R182 VGND.t88 VGND.n502 1253.59
R183 VGND.n2283 VGND.t413 1253.59
R184 VGND.t37 VGND.n2283 1253.59
R185 VGND.n538 VGND.t35 1253.59
R186 VGND.t142 VGND.n538 1253.59
R187 VGND.n2247 VGND.t410 1253.59
R188 VGND.t87 VGND.n2247 1253.59
R189 VGND.n1385 VGND.t39 1253.59
R190 VGND.t250 VGND.n1385 1253.59
R191 VGND.n1337 VGND.n1336 1243.48
R192 VGND.n2251 VGND.t985 1237.71
R193 VGND.n66 VGND.t1816 1213.79
R194 VGND.n2967 VGND.n2966 1198.25
R195 VGND.n1155 VGND.n1154 1198.25
R196 VGND.n2943 VGND.n2942 1180.79
R197 VGND.n2936 VGND.n2935 1180.79
R198 VGND.n2534 VGND.n208 1180.79
R199 VGND.n2529 VGND.n209 1180.79
R200 VGND.n2817 VGND.n210 1180.79
R201 VGND.n1989 VGND.n211 1180.79
R202 VGND.n1996 VGND.n212 1180.79
R203 VGND.n2842 VGND.n213 1180.79
R204 VGND.n1829 VGND.n214 1180.79
R205 VGND.n1836 VGND.n215 1180.79
R206 VGND.n2867 VGND.n216 1180.79
R207 VGND.n1655 VGND.n217 1180.79
R208 VGND.n1650 VGND.n218 1180.79
R209 VGND.n2892 VGND.n219 1180.79
R210 VGND.n1607 VGND.n220 1180.79
R211 VGND.n2912 VGND.n221 1180.79
R212 VGND.n1282 VGND.n222 1180.79
R213 VGND.n2918 VGND.n2917 1180.79
R214 VGND.n1335 VGND.n1334 1180.46
R215 VGND.n929 VGND.n890 1180.46
R216 VGND.n934 VGND.n933 1180.46
R217 VGND.n939 VGND.n938 1180.46
R218 VGND.n944 VGND.n943 1180.46
R219 VGND.n949 VGND.n948 1180.46
R220 VGND.n954 VGND.n953 1180.46
R221 VGND.n959 VGND.n958 1180.46
R222 VGND.n964 VGND.n963 1180.46
R223 VGND.n969 VGND.n968 1180.46
R224 VGND.n974 VGND.n973 1180.46
R225 VGND.n979 VGND.n978 1180.46
R226 VGND.n984 VGND.n983 1180.46
R227 VGND.n989 VGND.n988 1180.46
R228 VGND.n991 VGND.n990 1180.46
R229 VGND.n1279 VGND.n1278 1180.46
R230 VGND.n1277 VGND.n1276 1180.46
R231 VGND.n1234 VGND.n1233 1180.46
R232 VGND.n1239 VGND.n1238 1180.46
R233 VGND.n1241 VGND.n1240 1180.46
R234 VGND.n1246 VGND.n1245 1180.46
R235 VGND.n1248 VGND.n1247 1180.46
R236 VGND.n1220 VGND.n1219 1180.46
R237 VGND.n1209 VGND.n1208 1180.46
R238 VGND.n1207 VGND.n1206 1180.46
R239 VGND.n1190 VGND.n1189 1180.46
R240 VGND.n1188 VGND.n1187 1180.46
R241 VGND.n1177 VGND.n1176 1180.46
R242 VGND.n1175 VGND.n1174 1180.46
R243 VGND.n1167 VGND.n1166 1180.46
R244 VGND.n2775 VGND.n2774 1180.46
R245 VGND.n2777 VGND.n2776 1180.46
R246 VGND.n2732 VGND.n2731 1180.46
R247 VGND.n2737 VGND.n2736 1180.46
R248 VGND.n2739 VGND.n2738 1180.46
R249 VGND.n2728 VGND.n2727 1180.46
R250 VGND.n2706 VGND.n2705 1180.46
R251 VGND.n388 VGND.n327 1180.46
R252 VGND.n383 VGND.n382 1180.46
R253 VGND.n381 VGND.n380 1180.46
R254 VGND.n372 VGND.n371 1180.46
R255 VGND.n370 VGND.n369 1180.46
R256 VGND.n361 VGND.n360 1180.46
R257 VGND.n359 VGND.n333 1180.46
R258 VGND.n2701 VGND.n2700 1180.46
R259 VGND.n2641 VGND.n2640 1180.46
R260 VGND.n2646 VGND.n2645 1180.46
R261 VGND.n2651 VGND.n2650 1180.46
R262 VGND.n2656 VGND.n2655 1180.46
R263 VGND.n2661 VGND.n2660 1180.46
R264 VGND.n2666 VGND.n2665 1180.46
R265 VGND.n2671 VGND.n2670 1180.46
R266 VGND.n2673 VGND.n2672 1180.46
R267 VGND.n2717 VGND.n2716 1180.46
R268 VGND.n2719 VGND.n2718 1180.46
R269 VGND.n2750 VGND.n2749 1180.46
R270 VGND.n2757 VGND.n2756 1180.46
R271 VGND.n2755 VGND.n2754 1180.46
R272 VGND.n2790 VGND.n2789 1180.46
R273 VGND.n2792 VGND.n2791 1180.46
R274 VGND.n2345 VGND.n2344 1180.46
R275 VGND.n2340 VGND.n2339 1180.46
R276 VGND.n2335 VGND.n2334 1180.46
R277 VGND.n2330 VGND.n2329 1180.46
R278 VGND.n2325 VGND.n2324 1180.46
R279 VGND.n2320 VGND.n2319 1180.46
R280 VGND.n2315 VGND.n2314 1180.46
R281 VGND.n2310 VGND.n2309 1180.46
R282 VGND.n2305 VGND.n2304 1180.46
R283 VGND.n2300 VGND.n2299 1180.46
R284 VGND.n2295 VGND.n2294 1180.46
R285 VGND.n2290 VGND.n2289 1180.46
R286 VGND.n2545 VGND.n2544 1180.46
R287 VGND.n2543 VGND.n2542 1180.46
R288 VGND.n2538 VGND.n2537 1180.46
R289 VGND.n2355 VGND.n2354 1180.46
R290 VGND.n2379 VGND.n2378 1180.46
R291 VGND.n2381 VGND.n2380 1180.46
R292 VGND.n2405 VGND.n2404 1180.46
R293 VGND.n2407 VGND.n2406 1180.46
R294 VGND.n2431 VGND.n2430 1180.46
R295 VGND.n2433 VGND.n2432 1180.46
R296 VGND.n2457 VGND.n2456 1180.46
R297 VGND.n2459 VGND.n2458 1180.46
R298 VGND.n2483 VGND.n2482 1180.46
R299 VGND.n2485 VGND.n2484 1180.46
R300 VGND.n2514 VGND.n2513 1180.46
R301 VGND.n2519 VGND.n2518 1180.46
R302 VGND.n2524 VGND.n2523 1180.46
R303 VGND.n2526 VGND.n2525 1180.46
R304 VGND.n2366 VGND.n2365 1180.46
R305 VGND.n2368 VGND.n2367 1180.46
R306 VGND.n2392 VGND.n2391 1180.46
R307 VGND.n2394 VGND.n2393 1180.46
R308 VGND.n2418 VGND.n2417 1180.46
R309 VGND.n2420 VGND.n2419 1180.46
R310 VGND.n2444 VGND.n2443 1180.46
R311 VGND.n2446 VGND.n2445 1180.46
R312 VGND.n2470 VGND.n2469 1180.46
R313 VGND.n2472 VGND.n2471 1180.46
R314 VGND.n2496 VGND.n2495 1180.46
R315 VGND.n2503 VGND.n2502 1180.46
R316 VGND.n2501 VGND.n2500 1180.46
R317 VGND.n2812 VGND.n2811 1180.46
R318 VGND.n2814 VGND.n2813 1180.46
R319 VGND.n1913 VGND.n1912 1180.46
R320 VGND.n1915 VGND.n1914 1180.46
R321 VGND.n1924 VGND.n1923 1180.46
R322 VGND.n1926 VGND.n1925 1180.46
R323 VGND.n1935 VGND.n1934 1180.46
R324 VGND.n1937 VGND.n1936 1180.46
R325 VGND.n1946 VGND.n1945 1180.46
R326 VGND.n1948 VGND.n1947 1180.46
R327 VGND.n1957 VGND.n1956 1180.46
R328 VGND.n1959 VGND.n1958 1180.46
R329 VGND.n1968 VGND.n1967 1180.46
R330 VGND.n1970 VGND.n1969 1180.46
R331 VGND.n1979 VGND.n1978 1180.46
R332 VGND.n1984 VGND.n1983 1180.46
R333 VGND.n1986 VGND.n1985 1180.46
R334 VGND.n599 VGND.n598 1180.46
R335 VGND.n2060 VGND.n2059 1180.46
R336 VGND.n2058 VGND.n2057 1180.46
R337 VGND.n2053 VGND.n2052 1180.46
R338 VGND.n2048 VGND.n2047 1180.46
R339 VGND.n2043 VGND.n2042 1180.46
R340 VGND.n2038 VGND.n2037 1180.46
R341 VGND.n2033 VGND.n2032 1180.46
R342 VGND.n2028 VGND.n2027 1180.46
R343 VGND.n2023 VGND.n2022 1180.46
R344 VGND.n2018 VGND.n2017 1180.46
R345 VGND.n2013 VGND.n2012 1180.46
R346 VGND.n2008 VGND.n2007 1180.46
R347 VGND.n2003 VGND.n2002 1180.46
R348 VGND.n602 VGND.n601 1180.46
R349 VGND.n2072 VGND.n2071 1180.46
R350 VGND.n2077 VGND.n2076 1180.46
R351 VGND.n2082 VGND.n2081 1180.46
R352 VGND.n2087 VGND.n2086 1180.46
R353 VGND.n2092 VGND.n2091 1180.46
R354 VGND.n2097 VGND.n2096 1180.46
R355 VGND.n2102 VGND.n2101 1180.46
R356 VGND.n2107 VGND.n2106 1180.46
R357 VGND.n2112 VGND.n2111 1180.46
R358 VGND.n2117 VGND.n2116 1180.46
R359 VGND.n2122 VGND.n2121 1180.46
R360 VGND.n2129 VGND.n2128 1180.46
R361 VGND.n2127 VGND.n2126 1180.46
R362 VGND.n2837 VGND.n2836 1180.46
R363 VGND.n2839 VGND.n2838 1180.46
R364 VGND.n2179 VGND.n2178 1180.46
R365 VGND.n1754 VGND.n550 1180.46
R366 VGND.n1764 VGND.n1763 1180.46
R367 VGND.n1766 VGND.n1765 1180.46
R368 VGND.n1775 VGND.n1774 1180.46
R369 VGND.n1777 VGND.n1776 1180.46
R370 VGND.n1786 VGND.n1785 1180.46
R371 VGND.n1788 VGND.n1787 1180.46
R372 VGND.n1797 VGND.n1796 1180.46
R373 VGND.n1799 VGND.n1798 1180.46
R374 VGND.n1808 VGND.n1807 1180.46
R375 VGND.n1810 VGND.n1809 1180.46
R376 VGND.n1819 VGND.n1818 1180.46
R377 VGND.n1824 VGND.n1823 1180.46
R378 VGND.n1826 VGND.n1825 1180.46
R379 VGND.n1681 VGND.n1680 1180.46
R380 VGND.n1683 VGND.n1682 1180.46
R381 VGND.n1692 VGND.n1691 1180.46
R382 VGND.n1697 VGND.n1696 1180.46
R383 VGND.n1702 VGND.n1701 1180.46
R384 VGND.n1707 VGND.n1706 1180.46
R385 VGND.n1712 VGND.n1711 1180.46
R386 VGND.n1717 VGND.n1716 1180.46
R387 VGND.n1722 VGND.n1721 1180.46
R388 VGND.n1727 VGND.n1726 1180.46
R389 VGND.n1732 VGND.n1731 1180.46
R390 VGND.n1850 VGND.n1849 1180.46
R391 VGND.n1848 VGND.n1847 1180.46
R392 VGND.n1843 VGND.n1842 1180.46
R393 VGND.n1735 VGND.n1734 1180.46
R394 VGND.n672 VGND.n671 1180.46
R395 VGND.n677 VGND.n676 1180.46
R396 VGND.n682 VGND.n681 1180.46
R397 VGND.n687 VGND.n686 1180.46
R398 VGND.n692 VGND.n691 1180.46
R399 VGND.n697 VGND.n696 1180.46
R400 VGND.n702 VGND.n701 1180.46
R401 VGND.n707 VGND.n706 1180.46
R402 VGND.n712 VGND.n711 1180.46
R403 VGND.n717 VGND.n716 1180.46
R404 VGND.n722 VGND.n721 1180.46
R405 VGND.n729 VGND.n728 1180.46
R406 VGND.n727 VGND.n726 1180.46
R407 VGND.n2862 VGND.n2861 1180.46
R408 VGND.n2864 VGND.n2863 1180.46
R409 VGND.n1355 VGND.n1354 1180.46
R410 VGND.n877 VGND.n876 1180.46
R411 VGND.n872 VGND.n871 1180.46
R412 VGND.n821 VGND.n808 1180.46
R413 VGND.n826 VGND.n825 1180.46
R414 VGND.n831 VGND.n830 1180.46
R415 VGND.n836 VGND.n835 1180.46
R416 VGND.n841 VGND.n840 1180.46
R417 VGND.n846 VGND.n845 1180.46
R418 VGND.n851 VGND.n850 1180.46
R419 VGND.n858 VGND.n857 1180.46
R420 VGND.n856 VGND.n855 1180.46
R421 VGND.n1666 VGND.n1665 1180.46
R422 VGND.n1664 VGND.n1663 1180.46
R423 VGND.n1659 VGND.n1658 1180.46
R424 VGND.n1393 VGND.n1392 1180.46
R425 VGND.n1398 VGND.n1397 1180.46
R426 VGND.n1400 VGND.n1399 1180.46
R427 VGND.n1493 VGND.n1492 1180.46
R428 VGND.n1495 VGND.n1494 1180.46
R429 VGND.n1519 VGND.n1518 1180.46
R430 VGND.n1521 VGND.n1520 1180.46
R431 VGND.n1545 VGND.n1544 1180.46
R432 VGND.n1550 VGND.n1549 1180.46
R433 VGND.n1557 VGND.n1556 1180.46
R434 VGND.n1555 VGND.n1554 1180.46
R435 VGND.n1635 VGND.n1634 1180.46
R436 VGND.n1640 VGND.n1639 1180.46
R437 VGND.n1645 VGND.n1644 1180.46
R438 VGND.n1647 VGND.n1646 1180.46
R439 VGND.n1413 VGND.n1412 1180.46
R440 VGND.n1415 VGND.n1414 1180.46
R441 VGND.n1480 VGND.n1479 1180.46
R442 VGND.n1482 VGND.n1481 1180.46
R443 VGND.n1506 VGND.n1505 1180.46
R444 VGND.n1508 VGND.n1507 1180.46
R445 VGND.n1532 VGND.n1531 1180.46
R446 VGND.n1534 VGND.n1533 1180.46
R447 VGND.n1569 VGND.n1568 1180.46
R448 VGND.n1586 VGND.n1585 1180.46
R449 VGND.n1584 VGND.n1583 1180.46
R450 VGND.n1579 VGND.n1578 1180.46
R451 VGND.n1574 VGND.n1573 1180.46
R452 VGND.n2887 VGND.n2886 1180.46
R453 VGND.n2889 VGND.n2888 1180.46
R454 VGND.n1342 VGND.n1341 1180.46
R455 VGND.n1426 VGND.n1425 1180.46
R456 VGND.n1431 VGND.n1430 1180.46
R457 VGND.n1436 VGND.n1435 1180.46
R458 VGND.n1441 VGND.n1440 1180.46
R459 VGND.n1446 VGND.n1445 1180.46
R460 VGND.n1451 VGND.n1450 1180.46
R461 VGND.n1456 VGND.n1455 1180.46
R462 VGND.n1463 VGND.n1462 1180.46
R463 VGND.n1461 VGND.n1460 1180.46
R464 VGND.n1598 VGND.n1597 1180.46
R465 VGND.n1603 VGND.n1602 1180.46
R466 VGND.n1618 VGND.n1617 1180.46
R467 VGND.n1616 VGND.n1615 1180.46
R468 VGND.n1611 VGND.n1610 1180.46
R469 VGND.n1034 VGND.n1033 1180.46
R470 VGND.n1039 VGND.n1038 1180.46
R471 VGND.n1099 VGND.n1098 1180.46
R472 VGND.n1097 VGND.n1096 1180.46
R473 VGND.n1092 VGND.n1091 1180.46
R474 VGND.n1087 VGND.n1086 1180.46
R475 VGND.n1082 VGND.n1081 1180.46
R476 VGND.n1077 VGND.n1076 1180.46
R477 VGND.n1072 VGND.n1071 1180.46
R478 VGND.n1050 VGND.n1041 1180.46
R479 VGND.n1055 VGND.n1054 1180.46
R480 VGND.n1060 VGND.n1059 1180.46
R481 VGND.n1062 VGND.n1061 1180.46
R482 VGND.n2907 VGND.n2906 1180.46
R483 VGND.n2909 VGND.n2908 1180.46
R484 VGND.t1815 VGND.n3011 1180.08
R485 VGND.n1387 VGND.n1386 1169.57
R486 VGND.n3015 VGND.t1 1146.36
R487 VGND.n3017 VGND.t0 1112.64
R488 VGND.n3016 VGND.t1589 1112.64
R489 VGND.n2351 VGND.n2349 1070.21
R490 VGND.n2968 VGND 1055.35
R491 VGND.n2251 VGND.n2250 1052.29
R492 VGND.t1139 VGND.n2181 1032.59
R493 VGND.t1156 VGND.n2641 988.926
R494 VGND.t1608 VGND.n2646 988.926
R495 VGND.t556 VGND.n2651 988.926
R496 VGND.t1554 VGND.n2656 988.926
R497 VGND.t262 VGND.n2661 988.926
R498 VGND.t732 VGND.n2666 988.926
R499 VGND.t570 VGND.n2671 988.926
R500 VGND.n2672 VGND.t676 988.926
R501 VGND.t217 VGND.n2717 988.926
R502 VGND.n2718 VGND.t1216 988.926
R503 VGND.t1746 VGND.n2750 988.926
R504 VGND.n2756 VGND.t2424 988.926
R505 VGND.n2755 VGND.t914 988.926
R506 VGND.t465 VGND.n2790 988.926
R507 VGND.n2791 VGND.t289 988.926
R508 VGND.n2345 VGND.t832 988.926
R509 VGND.n2340 VGND.t373 988.926
R510 VGND.n2335 VGND.t114 988.926
R511 VGND.n2330 VGND.t1546 988.926
R512 VGND.n2325 VGND.t1750 988.926
R513 VGND.n2320 VGND.t300 988.926
R514 VGND.n2315 VGND.t1669 988.926
R515 VGND.n2310 VGND.t333 988.926
R516 VGND.n2305 VGND.t1841 988.926
R517 VGND.n2300 VGND.t456 988.926
R518 VGND.n2295 VGND.t709 988.926
R519 VGND.n2290 VGND.t1615 988.926
R520 VGND.n2544 VGND.t1260 988.926
R521 VGND.n2543 VGND.t32 988.926
R522 VGND.n2538 VGND.t2433 988.926
R523 VGND.n2354 VGND.t81 988.926
R524 VGND.t1982 VGND.n2379 988.926
R525 VGND.n2380 VGND.t605 988.926
R526 VGND.t1561 VGND.n2405 988.926
R527 VGND.n2406 VGND.t1824 988.926
R528 VGND.t320 VGND.n2431 988.926
R529 VGND.n2432 VGND.t129 988.926
R530 VGND.t337 VGND.n2457 988.926
R531 VGND.n2458 VGND.t666 988.926
R532 VGND.t434 VGND.n2483 988.926
R533 VGND.n2484 VGND.t1740 988.926
R534 VGND.t185 VGND.n2514 988.926
R535 VGND.t920 VGND.n2519 988.926
R536 VGND.t365 VGND.n2524 988.926
R537 VGND.n2525 VGND.t510 988.926
R538 VGND.t836 VGND.n2366 988.926
R539 VGND.n2367 VGND.t1832 988.926
R540 VGND.t529 VGND.n2392 988.926
R541 VGND.n2393 VGND.t9 988.926
R542 VGND.t1315 VGND.n2418 988.926
R543 VGND.n2419 VGND.t692 988.926
R544 VGND.t550 VGND.n2444 988.926
R545 VGND.n2445 VGND.t316 988.926
R546 VGND.t598 VGND.n2470 988.926
R547 VGND.n2471 VGND.t164 988.926
R548 VGND.t1126 VGND.n2496 988.926
R549 VGND.n2502 VGND.t1220 988.926
R550 VGND.n2501 VGND.t2682 988.926
R551 VGND.t1351 VGND.n2812 988.926
R552 VGND.n2813 VGND.t281 988.926
R553 VGND.t1148 VGND.n1913 988.926
R554 VGND.n1914 VGND.t2677 988.926
R555 VGND.t108 VGND.n1924 988.926
R556 VGND.n1925 VGND.t1539 988.926
R557 VGND.t1699 VGND.n1935 988.926
R558 VGND.n1936 VGND.t296 988.926
R559 VGND.t136 VGND.n1946 988.926
R560 VGND.n1947 VGND.t642 988.926
R561 VGND.t1137 VGND.n1957 988.926
R562 VGND.n1958 VGND.t442 988.926
R563 VGND.t1812 VGND.n1968 988.926
R564 VGND.n1969 VGND.t2421 988.926
R565 VGND.t1254 VGND.n1979 988.926
R566 VGND.t24 VGND.n1984 988.926
R567 VGND.n1985 VGND.t518 988.926
R568 VGND.t1154 VGND.n599 988.926
R569 VGND.n2059 VGND.t1606 988.926
R570 VGND.n2058 VGND.t553 988.926
R571 VGND.n2053 VGND.t1552 988.926
R572 VGND.n2048 VGND.t260 988.926
R573 VGND.n2043 VGND.t730 988.926
R574 VGND.n2038 VGND.t568 988.926
R575 VGND.n2033 VGND.t674 988.926
R576 VGND.n2028 VGND.t215 988.926
R577 VGND.n2023 VGND.t1213 988.926
R578 VGND.n2018 VGND.t1744 988.926
R579 VGND.n2013 VGND.t1218 988.926
R580 VGND.n2008 VGND.t912 988.926
R581 VGND.n2003 VGND.t462 988.926
R582 VGND.n601 VGND.t287 988.926
R583 VGND.t622 VGND.n2072 988.926
R584 VGND.t1984 VGND.n2077 988.926
R585 VGND.t603 VGND.n2082 988.926
R586 VGND.t1235 VGND.n2087 988.926
R587 VGND.t1826 VGND.n2092 988.926
R588 VGND.t322 VGND.n2097 988.926
R589 VGND.t131 VGND.n2102 988.926
R590 VGND.t339 VGND.n2107 988.926
R591 VGND.t668 VGND.n2112 988.926
R592 VGND.t436 VGND.n2117 988.926
R593 VGND.t1742 VGND.n2122 988.926
R594 VGND.n2128 VGND.t187 988.926
R595 VGND.n2127 VGND.t922 988.926
R596 VGND.t367 VGND.n2837 988.926
R597 VGND.n2838 VGND.t512 988.926
R598 VGND.n2179 VGND.t838 988.926
R599 VGND.t1834 VGND.n1754 988.926
R600 VGND.t527 VGND.n1764 988.926
R601 VGND.n1765 VGND.t11 988.926
R602 VGND.t1599 VGND.n1775 988.926
R603 VGND.n1776 VGND.t694 988.926
R604 VGND.t564 VGND.n1786 988.926
R605 VGND.n1787 VGND.t318 988.926
R606 VGND.t600 VGND.n1797 988.926
R607 VGND.n1798 VGND.t1208 988.926
R608 VGND.t1128 VGND.n1808 988.926
R609 VGND.n1809 VGND.t1222 988.926
R610 VGND.t2684 VGND.n1819 988.926
R611 VGND.t1353 VGND.n1824 988.926
R612 VGND.n1825 VGND.t283 988.926
R613 VGND.t1160 VGND.n1681 988.926
R614 VGND.n1682 VGND.t591 988.926
R615 VGND.t533 VGND.n1692 988.926
R616 VGND.t5 VGND.n1697 988.926
R617 VGND.t1309 VGND.n1702 988.926
R618 VGND.t690 VGND.n1707 988.926
R619 VGND.t546 VGND.n1712 988.926
R620 VGND.t19 VGND.n1717 988.926
R621 VGND.t1586 VGND.n1722 988.926
R622 VGND.t162 VGND.n1727 988.926
R623 VGND.t1124 VGND.n1732 988.926
R624 VGND.n1849 VGND.t1349 988.926
R625 VGND.n1848 VGND.t1999 988.926
R626 VGND.n1843 VGND.t1377 988.926
R627 VGND.n1734 VGND.t179 988.926
R628 VGND.t1146 VGND.n672 988.926
R629 VGND.t2675 VGND.n677 988.926
R630 VGND.t110 VGND.n682 988.926
R631 VGND.t1537 VGND.n687 988.926
R632 VGND.t1977 VGND.n692 988.926
R633 VGND.t328 VGND.n697 988.926
R634 VGND.t134 VGND.n702 988.926
R635 VGND.t640 VGND.n707 988.926
R636 VGND.t1135 VGND.n712 988.926
R637 VGND.t440 VGND.n717 988.926
R638 VGND.t1810 VGND.n722 988.926
R639 VGND.n728 VGND.t2419 988.926
R640 VGND.n727 VGND.t1252 988.926
R641 VGND.t22 VGND.n2862 988.926
R642 VGND.n2863 VGND.t516 988.926
R643 VGND.n1355 VGND.t754 988.926
R644 VGND.n877 VGND.t1603 988.926
R645 VGND.n872 VGND.t520 988.926
R646 VGND.t1442 VGND.n821 988.926
R647 VGND.t1307 VGND.n826 988.926
R648 VGND.t1083 VGND.n831 988.926
R649 VGND.t539 VGND.n836 988.926
R650 VGND.t721 VGND.n841 988.926
R651 VGND.t210 VGND.n846 988.926
R652 VGND.t156 VGND.n851 988.926
R653 VGND.n857 VGND.t1317 988.926
R654 VGND.n856 VGND.t1243 988.926
R655 VGND.n1665 VGND.t1992 988.926
R656 VGND.n1664 VGND.t1535 988.926
R657 VGND.n1659 VGND.t171 988.926
R658 VGND.t79 VGND.n1393 988.926
R659 VGND.t1980 VGND.n1398 988.926
R660 VGND.n1399 VGND.t808 988.926
R661 VGND.t1559 VGND.n1493 988.926
R662 VGND.n1494 VGND.t1822 988.926
R663 VGND.t736 VGND.n1519 988.926
R664 VGND.n1520 VGND.t574 988.926
R665 VGND.t335 VGND.n1545 988.926
R666 VGND.t664 VGND.n1550 988.926
R667 VGND.n1556 VGND.t2543 988.926
R668 VGND.n1555 VGND.t1738 988.926
R669 VGND.t183 VGND.n1635 988.926
R670 VGND.t918 VGND.n1640 988.926
R671 VGND.t363 VGND.n1645 988.926
R672 VGND.n1646 VGND.t508 988.926
R673 VGND.t752 VGND.n1413 988.926
R674 VGND.n1414 VGND.t1601 988.926
R675 VGND.t522 VGND.n1480 988.926
R676 VGND.n1481 VGND.t1440 988.926
R677 VGND.t1305 VGND.n1506 988.926
R678 VGND.n1507 VGND.t1081 988.926
R679 VGND.t537 VGND.n1532 988.926
R680 VGND.n1533 VGND.t719 988.926
R681 VGND.t208 VGND.n1569 988.926
R682 VGND.n1585 VGND.t154 988.926
R683 VGND.n1584 VGND.t1267 988.926
R684 VGND.n1579 VGND.t1241 988.926
R685 VGND.n1574 VGND.t1990 988.926
R686 VGND.t1533 VGND.n2887 988.926
R687 VGND.n2888 VGND.t169 988.926
R688 VGND.n1341 VGND.t830 988.926
R689 VGND.t371 VGND.n1426 988.926
R690 VGND.t578 VGND.n1431 988.926
R691 VGND.t1543 VGND.n1436 988.926
R692 VGND.t1703 VGND.n1441 988.926
R693 VGND.t298 VGND.n1446 988.926
R694 VGND.t1667 VGND.n1451 988.926
R695 VGND.t331 VGND.n1456 988.926
R696 VGND.n1462 VGND.t1839 988.926
R697 VGND.n1461 VGND.t453 988.926
R698 VGND.t707 VGND.n1598 988.926
R699 VGND.t1612 VGND.n1603 988.926
R700 VGND.n1617 VGND.t1258 988.926
R701 VGND.n1616 VGND.t26 988.926
R702 VGND.n1611 VGND.t2430 988.926
R703 VGND.t1162 VGND.n1034 988.926
R704 VGND.t593 VGND.n1039 988.926
R705 VGND.n1098 VGND.t531 988.926
R706 VGND.n1097 VGND.t7 988.926
R707 VGND.n1092 VGND.t1311 988.926
R708 VGND.n1087 VGND.t432 988.926
R709 VGND.n1082 VGND.t544 988.926
R710 VGND.n1077 VGND.t17 988.926
R711 VGND.n1072 VGND.t1584 988.926
R712 VGND.t160 VGND.n1050 988.926
R713 VGND.t1122 VGND.n1055 988.926
R714 VGND.t1347 VGND.n1060 988.926
R715 VGND.n1061 VGND.t1997 988.926
R716 VGND.t1379 VGND.n2907 988.926
R717 VGND.n2908 VGND.t177 988.926
R718 VGND.n1335 VGND.t2667 988.926
R719 VGND.t2585 VGND.n929 988.926
R720 VGND.t2217 VGND.n934 988.926
R721 VGND.t2662 VGND.n939 988.926
R722 VGND.t2651 VGND.n944 988.926
R723 VGND.t2632 VGND.n949 988.926
R724 VGND.t2145 VGND.n954 988.926
R725 VGND.t1507 VGND.n959 988.926
R726 VGND.t2628 VGND.n964 988.926
R727 VGND.t2205 VGND.n969 988.926
R728 VGND.t2192 VGND.n974 988.926
R729 VGND.t2117 VGND.n979 988.926
R730 VGND.t2611 VGND.n984 988.926
R731 VGND.t2174 VGND.n989 988.926
R732 VGND.n990 VGND.t2126 988.926
R733 VGND.n2248 VGND.n539 934.784
R734 VGND.n116 VGND 927.203
R735 VGND.n134 VGND 927.203
R736 VGND.n2182 VGND 918.774
R737 VGND.n194 VGND 910.346
R738 VGND.n165 VGND 910.346
R739 VGND.t1367 VGND.n2967 909.365
R740 VGND.n2285 VGND.n473 900
R741 VGND.n2641 VGND.t1251 852.769
R742 VGND.n2646 VGND.t2673 852.769
R743 VGND.n2651 VGND.t1187 852.769
R744 VGND.n2656 VGND.t659 852.769
R745 VGND.n2661 VGND.t238 852.769
R746 VGND.n2666 VGND.t1120 852.769
R747 VGND.n2671 VGND.t2562 852.769
R748 VGND.n2672 VGND.t645 852.769
R749 VGND.n2717 VGND.t448 852.769
R750 VGND.n2718 VGND.t1134 852.769
R751 VGND.n2750 VGND.t2535 852.769
R752 VGND.n2756 VGND.t860 852.769
R753 VGND.t2560 VGND.n2755 852.769
R754 VGND.n2790 VGND.t13 852.769
R755 VGND.n2791 VGND.t663 852.769
R756 VGND.n2935 VGND.t354 852.769
R757 VGND.t829 VGND.n2345 852.769
R758 VGND.t932 VGND.n2340 852.769
R759 VGND.t450 VGND.n2335 852.769
R760 VGND.t1845 VGND.n2330 852.769
R761 VGND.t1133 VGND.n2325 852.769
R762 VGND.t843 VGND.n2320 852.769
R763 VGND.t2493 VGND.n2315 852.769
R764 VGND.t1371 VGND.n2310 852.769
R765 VGND.t358 VGND.n2305 852.769
R766 VGND.t689 VGND.n2300 852.769
R767 VGND.t232 VGND.n2295 852.769
R768 VGND.t897 VGND.n2290 852.769
R769 VGND.n2544 VGND.t1836 852.769
R770 VGND.t1806 VGND.n2543 852.769
R771 VGND.t75 VGND.n2538 852.769
R772 VGND.t28 VGND.n208 852.769
R773 VGND.n2354 VGND.t2233 852.769
R774 VGND.n2379 VGND.t2561 852.769
R775 VGND.n2380 VGND.t687 852.769
R776 VGND.n2405 VGND.t251 852.769
R777 VGND.n2406 VGND.t2098 852.769
R778 VGND.n2431 VGND.t1484 852.769
R779 VGND.n2432 VGND.t882 852.769
R780 VGND.n2457 VGND.t2100 852.769
R781 VGND.n2458 VGND.t908 852.769
R782 VGND.n2483 VGND.t1357 852.769
R783 VGND.n2484 VGND.t151 852.769
R784 VGND.n2514 VGND.t204 852.769
R785 VGND.n2519 VGND.t1576 852.769
R786 VGND.n2524 VGND.t1121 852.769
R787 VGND.n2525 VGND.t276 852.769
R788 VGND.t1987 VGND.n209 852.769
R789 VGND.n2366 VGND.t264 852.769
R790 VGND.n2367 VGND.t728 852.769
R791 VGND.n2392 VGND.t718 852.769
R792 VGND.n2393 VGND.t1578 852.769
R793 VGND.n2418 VGND.t660 852.769
R794 VGND.n2419 VGND.t883 852.769
R795 VGND.n2444 VGND.t928 852.769
R796 VGND.n2445 VGND.t1341 852.769
R797 VGND.n2470 VGND.t2101 852.769
R798 VGND.n2471 VGND.t445 852.769
R799 VGND.n2496 VGND.t242 852.769
R800 VGND.n2502 VGND.t1818 852.769
R801 VGND.t166 VGND.n2501 852.769
R802 VGND.n2812 VGND.t909 852.769
R803 VGND.n2813 VGND.t1145 852.769
R804 VGND.t256 VGND.n210 852.769
R805 VGND.n1913 VGND.t2533 852.769
R806 VGND.n1914 VGND.t235 852.769
R807 VGND.n1924 VGND.t447 852.769
R808 VGND.n1925 VGND.t772 852.769
R809 VGND.n1935 VGND.t1849 852.769
R810 VGND.n1936 VGND.t907 852.769
R811 VGND.n1946 VGND.t1188 852.769
R812 VGND.n1947 VGND.t1581 852.769
R813 VGND.n1957 VGND.t1577 852.769
R814 VGND.n1958 VGND.t2531 852.769
R815 VGND.n1968 VGND.t231 852.769
R816 VGND.n1969 VGND.t716 852.769
R817 VGND.n1979 VGND.t771 852.769
R818 VGND.n1984 VGND.t725 852.769
R819 VGND.n1985 VGND.t1549 852.769
R820 VGND.t2097 VGND.n211 852.769
R821 VGND.n599 VGND.t2391 852.769
R822 VGND.n2059 VGND.t1805 852.769
R823 VGND.t779 VGND.n2058 852.769
R824 VGND.t94 VGND.n2053 852.769
R825 VGND.t452 VGND.n2048 852.769
R826 VGND.t770 VGND.n2043 852.769
R827 VGND.t2082 VGND.n2038 852.769
R828 VGND.t280 VGND.n2033 852.769
R829 VGND.t1185 VGND.n2028 852.769
R830 VGND.t656 VGND.n2023 852.769
R831 VGND.t2091 VGND.n2018 852.769
R832 VGND.t1141 VGND.n2013 852.769
R833 VGND.t2099 VGND.n2008 852.769
R834 VGND.t356 VGND.n2003 852.769
R835 VGND.n601 VGND.t1531 852.769
R836 VGND.t230 VGND.n212 852.769
R837 VGND.n2072 VGND.t1264 852.769
R838 VGND.n2077 VGND.t1456 852.769
R839 VGND.n2082 VGND.t206 852.769
R840 VGND.n2087 VGND.t275 852.769
R841 VGND.n2092 VGND.t139 852.769
R842 VGND.n2097 VGND.t2416 852.769
R843 VGND.n2102 VGND.t92 852.769
R844 VGND.n2107 VGND.t1461 852.769
R845 VGND.n2112 VGND.t221 852.769
R846 VGND.n2117 VGND.t2417 852.769
R847 VGND.n2122 VGND.t446 852.769
R848 VGND.n2128 VGND.t1249 852.769
R849 VGND.t1270 VGND.n2127 852.769
R850 VGND.n2837 VGND.t1250 852.769
R851 VGND.n2838 VGND.t938 852.769
R852 VGND.t1186 VGND.n213 852.769
R853 VGND.t560 VGND.n2179 852.769
R854 VGND.n1754 VGND.t1088 852.769
R855 VGND.n1764 VGND.t1503 852.769
R856 VGND.n1765 VGND.t905 852.769
R857 VGND.n1775 VGND.t562 852.769
R858 VGND.n1776 VGND.t1373 852.769
R859 VGND.n1786 VGND.t252 852.769
R860 VGND.n1787 VGND.t717 852.769
R861 VGND.n1797 VGND.t929 852.769
R862 VGND.n1798 VGND.t1851 852.769
R863 VGND.n1808 VGND.t647 852.769
R864 VGND.n1809 VGND.t1339 852.769
R865 VGND.n1819 VGND.t225 852.769
R866 VGND.n1824 VGND.t239 852.769
R867 VGND.n1825 VGND.t91 852.769
R868 VGND.t1343 VGND.n214 852.769
R869 VGND.n1681 VGND.t609 852.769
R870 VGND.n1682 VGND.t726 852.769
R871 VGND.n1692 VGND.t1819 852.769
R872 VGND.n1697 VGND.t1592 852.769
R873 VGND.n1702 VGND.t2001 852.769
R874 VGND.n1707 VGND.t706 852.769
R875 VGND.n1712 VGND.t773 852.769
R876 VGND.n1717 VGND.t234 852.769
R877 VGND.n1722 VGND.t828 852.769
R878 VGND.n1727 VGND.t205 852.769
R879 VGND.n1732 VGND.t646 852.769
R880 VGND.n1849 VGND.t1416 852.769
R881 VGND.t181 VGND.n1848 852.769
R882 VGND.t1132 VGND.n1843 852.769
R883 VGND.n1734 VGND.t2418 852.769
R884 VGND.t1580 VGND.n215 852.769
R885 VGND.n672 VGND.t2081 852.769
R886 VGND.n677 VGND.t715 852.769
R887 VGND.n682 VGND.t826 852.769
R888 VGND.n687 VGND.t931 852.769
R889 VGND.n692 VGND.t84 852.769
R890 VGND.n697 VGND.t1594 852.769
R891 VGND.n702 VGND.t781 852.769
R892 VGND.n707 VGND.t119 852.769
R893 VGND.n712 VGND.t888 852.769
R894 VGND.n717 VGND.t2536 852.769
R895 VGND.n722 VGND.t825 852.769
R896 VGND.n728 VGND.t1421 852.769
R897 VGND.t1269 VGND.n727 852.769
R898 VGND.n2862 VGND.t253 852.769
R899 VGND.n2863 VGND.t1548 852.769
R900 VGND.t213 VGND.n216 852.769
R901 VGND.t182 VGND.n1355 852.769
R902 VGND.t2403 VGND.n877 852.769
R903 VGND.t212 VGND.n872 852.769
R904 VGND.n821 VGND.t85 852.769
R905 VGND.n826 VGND.t118 852.769
R906 VGND.n831 VGND.t1144 852.769
R907 VGND.n836 VGND.t1452 852.769
R908 VGND.n841 VGND.t1595 852.769
R909 VGND.n846 VGND.t1501 852.769
R910 VGND.n851 VGND.t1142 852.769
R911 VGND.n857 VGND.t241 852.769
R912 VGND.t661 VGND.n856 852.769
R913 VGND.n1665 VGND.t2102 852.769
R914 VGND.t561 VGND.n1664 852.769
R915 VGND.t2559 VGND.n1659 852.769
R916 VGND.t86 VGND.n217 852.769
R917 VGND.n1393 VGND.t898 852.769
R918 VGND.n1398 VGND.t1342 852.769
R919 VGND.n1399 VGND.t1455 852.769
R920 VGND.n1493 VGND.t1372 852.769
R921 VGND.n1494 VGND.t1502 852.769
R922 VGND.n1519 VGND.t1265 852.769
R923 VGND.n1520 VGND.t140 852.769
R924 VGND.n1545 VGND.t1532 852.769
R925 VGND.n1550 VGND.t1420 852.769
R926 VGND.n1556 VGND.t469 852.769
R927 VGND.t1344 VGND.n1555 852.769
R928 VGND.n1635 VGND.t927 852.769
R929 VGND.n1640 VGND.t128 852.769
R930 VGND.n1645 VGND.t279 852.769
R931 VGND.n1646 VGND.t1979 852.769
R932 VGND.t2392 VGND.n218 852.769
R933 VGND.n1413 VGND.t30 852.769
R934 VGND.n1414 VGND.t608 852.769
R935 VGND.n1480 VGND.t2092 852.769
R936 VGND.n1481 VGND.t2674 852.769
R937 VGND.n1506 VGND.t1415 852.769
R938 VGND.n1507 VGND.t76 852.769
R939 VGND.n1532 VGND.t1814 852.769
R940 VGND.n1533 VGND.t2537 852.769
R941 VGND.n1569 VGND.t147 852.769
R942 VGND.n1585 VGND.t536 852.769
R943 VGND.t778 VGND.n1584 852.769
R944 VGND.t887 VGND.n1579 852.769
R945 VGND.t449 VGND.n1574 852.769
R946 VGND.n2887 VGND.t355 852.769
R947 VGND.n2888 VGND.t1829 852.769
R948 VGND.t150 VGND.n219 852.769
R949 VGND.n1341 VGND.t925 852.769
R950 VGND.n1426 VGND.t1418 852.769
R951 VGND.n1431 VGND.t559 852.769
R952 VGND.n1436 VGND.t827 852.769
R953 VGND.n1441 VGND.t2534 852.769
R954 VGND.n1446 VGND.t2532 852.769
R955 VGND.n1451 VGND.t1419 852.769
R956 VGND.n1456 VGND.t117 852.769
R957 VGND.n1462 VGND.t1337 852.769
R958 VGND.t203 VGND.n1461 852.769
R959 VGND.n1598 VGND.t1080 852.769
R960 VGND.n1603 VGND.t1830 852.769
R961 VGND.n1617 VGND.t681 852.769
R962 VGND.t926 VGND.n1616 852.769
R963 VGND.t388 VGND.n1611 852.769
R964 VGND.t1579 VGND.n220 852.769
R965 VGND.n1034 VGND.t841 852.769
R966 VGND.n1039 VGND.t468 852.769
R967 VGND.n1098 VGND.t74 852.769
R968 VGND.t842 VGND.n1097 852.769
R969 VGND.t1844 VGND.n1092 852.769
R970 VGND.t236 VGND.n1087 852.769
R971 VGND.t1374 VGND.n1082 852.769
R972 VGND.t780 VGND.n1077 852.769
R973 VGND.t861 VGND.n1072 852.769
R974 VGND.n1050 VGND.t886 852.769
R975 VGND.n1055 VGND.t688 852.769
R976 VGND.n1060 VGND.t1588 852.769
R977 VGND.n1061 VGND.t697 852.769
R978 VGND.n2907 VGND.t1143 852.769
R979 VGND.n2908 VGND.t1089 852.769
R980 VGND.t278 VGND.n221 852.769
R981 VGND.t558 VGND.n1335 852.769
R982 VGND.n929 VGND.t930 852.769
R983 VGND.n934 VGND.t1199 852.769
R984 VGND.n939 VGND.t385 852.769
R985 VGND.n944 VGND.t1593 852.769
R986 VGND.n949 VGND.t359 852.769
R987 VGND.n954 VGND.t228 852.769
R988 VGND.n959 VGND.t149 852.769
R989 VGND.n964 VGND.t910 852.769
R990 VGND.n969 VGND.t2234 852.769
R991 VGND.n974 VGND.t2538 852.769
R992 VGND.n979 VGND.t233 852.769
R993 VGND.n984 VGND.t658 852.769
R994 VGND.n989 VGND.t90 852.769
R995 VGND.n990 VGND.t222 852.769
R996 VGND.n2918 VGND.t444 852.769
R997 VGND.n2249 VGND 851.341
R998 VGND.n2944 VGND.n2943 846.154
R999 VGND.n2350 VGND.t982 809.773
R1000 VGND.n2352 VGND.t1057 809.773
R1001 VGND.t964 VGND.n2353 809.773
R1002 VGND.n473 VGND.t1006 809.773
R1003 VGND.t1078 VGND.n503 809.773
R1004 VGND.t958 VGND.n504 809.773
R1005 VGND.n2180 VGND.t1000 809.773
R1006 VGND.t1012 VGND.n539 809.773
R1007 VGND.n1387 VGND.t1036 809.773
R1008 VGND.t967 VGND.n1388 809.773
R1009 VGND.n1339 VGND.t1039 809.773
R1010 VGND.t1069 VGND.n1340 809.773
R1011 VGND.n1338 VGND.t1009 809.773
R1012 VGND.n1336 VGND.t2160 809.773
R1013 VGND.t2321 VGND.t2303 708.047
R1014 VGND.t2303 VGND.t2301 708.047
R1015 VGND.t2301 VGND.t2311 708.047
R1016 VGND.t2311 VGND.t102 708.047
R1017 VGND.t102 VGND.t99 708.047
R1018 VGND.t99 VGND.t105 708.047
R1019 VGND.t105 VGND.t96 708.047
R1020 VGND.t2288 VGND.t0 708.047
R1021 VGND.t2317 VGND.t2356 708.047
R1022 VGND.t2356 VGND.t2325 708.047
R1023 VGND.t2325 VGND.t2299 708.047
R1024 VGND.t2299 VGND.t98 708.047
R1025 VGND.t98 VGND.t104 708.047
R1026 VGND.t104 VGND.t101 708.047
R1027 VGND.t101 VGND.t107 708.047
R1028 VGND.t2372 VGND.t2319 708.047
R1029 VGND.t2319 VGND.t2360 708.047
R1030 VGND.t2360 VGND.t2328 708.047
R1031 VGND.t2328 VGND.t352 708.047
R1032 VGND.t352 VGND.t348 708.047
R1033 VGND.t348 VGND.t342 708.047
R1034 VGND.t342 VGND.t344 708.047
R1035 VGND.t2285 VGND.t1 708.047
R1036 VGND.t2348 VGND.t2337 708.047
R1037 VGND.t2337 VGND.t2335 708.047
R1038 VGND.t2335 VGND.t2295 708.047
R1039 VGND.t2295 VGND.t858 708.047
R1040 VGND.t858 VGND.t1200 708.047
R1041 VGND.t1200 VGND.t244 708.047
R1042 VGND.t244 VGND.t375 708.047
R1043 VGND.t2313 VGND.t2352 708.047
R1044 VGND.t2352 VGND.t2323 708.047
R1045 VGND.t2323 VGND.t2333 708.047
R1046 VGND.t2333 VGND.t607 708.047
R1047 VGND.t607 VGND.t246 708.047
R1048 VGND.t246 VGND.t1848 708.047
R1049 VGND.t1848 VGND.t243 708.047
R1050 VGND.t2309 VGND.t2365 708.047
R1051 VGND.t2370 VGND.t2309 708.047
R1052 VGND.t2342 VGND.t2370 708.047
R1053 VGND.t350 VGND.t2342 708.047
R1054 VGND.t346 VGND.t350 708.047
R1055 VGND.t351 VGND.t346 708.047
R1056 VGND.t347 VGND.t351 708.047
R1057 VGND.n2971 VGND.n2970 708.047
R1058 VGND.t1245 VGND.t1590 691.188
R1059 VGND.t2077 VGND.t254 691.188
R1060 VGND.t2376 VGND.t2354 657.471
R1061 VGND.t2350 VGND.t1368 657.471
R1062 VGND.t2387 VGND.t1364 657.471
R1063 VGND.t2330 VGND.t1358 657.471
R1064 VGND.t1468 VGND.t1170 657.471
R1065 VGND.t627 VGND.t1168 657.471
R1066 VGND.t408 VGND.t1166 657.471
R1067 VGND.t42 VGND.t637 657.471
R1068 VGND.t2354 VGND.t2380 654.197
R1069 VGND.t637 VGND.t1475 654.197
R1070 VGND VGND.n194 640.614
R1071 VGND VGND.n134 640.614
R1072 VGND VGND.n165 640.614
R1073 VGND.n2182 VGND 640.614
R1074 VGND.n116 VGND 632.184
R1075 VGND.t1436 VGND.t757 630.62
R1076 VGND.t589 VGND.t782 630.62
R1077 VGND.t535 VGND.t2567 630.62
R1078 VGND.t1551 VGND.t2565 630.62
R1079 VGND.t1771 VGND.t1434 630.62
R1080 VGND.t1090 VGND.t1411 630.62
R1081 VGND.t542 VGND.t2575 630.62
R1082 VGND.t15 VGND.t1432 630.62
R1083 VGND.t1430 VGND.t387 630.62
R1084 VGND.t159 VGND.t1413 630.62
R1085 VGND.t2563 VGND.t712 630.62
R1086 VGND.t1346 VGND.t1438 630.62
R1087 VGND.t2573 VGND.t1995 630.62
R1088 VGND.t2571 VGND.t1376 630.62
R1089 VGND.t286 VGND.t2569 630.62
R1090 VGND.t1428 VGND.t2114 630.62
R1091 VGND.t700 VGND.t78 630.62
R1092 VGND.t1112 VGND.t1611 630.62
R1093 VGND.t472 VGND.t602 630.62
R1094 VGND.t470 VGND.t1542 630.62
R1095 VGND.t698 VGND.t1821 630.62
R1096 VGND.t1195 VGND.t431 630.62
R1097 VGND.t1193 VGND.t573 630.62
R1098 VGND.t1118 VGND.t679 630.62
R1099 VGND.t1116 VGND.t220 630.62
R1100 VGND.t1197 VGND.t438 630.62
R1101 VGND.t704 VGND.t1322 630.62
R1102 VGND.t702 VGND.t189 630.62
R1103 VGND.t1191 VGND.t917 630.62
R1104 VGND.t1189 VGND.t223 630.62
R1105 VGND.t474 VGND.t2429 630.62
R1106 VGND.t1114 VGND.t2186 630.62
R1107 VGND.t1159 VGND.t1787 630.62
R1108 VGND.t1522 VGND.t595 630.62
R1109 VGND.t525 VGND.t1795 630.62
R1110 VGND.t1793 VGND.t1557 630.62
R1111 VGND.t1313 VGND.t1785 630.62
R1112 VGND.t1327 VGND.t1092 630.62
R1113 VGND.t548 VGND.t1325 630.62
R1114 VGND.t1528 VGND.t21 630.62
R1115 VGND.t596 VGND.t1526 630.62
R1116 VGND.t1329 VGND.t1211 630.62
R1117 VGND.t714 VGND.t1791 630.62
R1118 VGND.t1789 VGND.t1225 630.62
R1119 VGND.t83 VGND.t1323 630.62
R1120 VGND.t1356 VGND.t1799 630.62
R1121 VGND.t292 VGND.t1797 630.62
R1122 VGND.t1524 VGND.t2135 630.62
R1123 VGND.t1271 VGND.t576 630.62
R1124 VGND.t846 VGND.t2089 630.62
R1125 VGND.t1102 VGND.t580 630.62
R1126 VGND.t3 VGND.t1277 630.62
R1127 VGND.t482 VGND.t1303 630.62
R1128 VGND.t326 VGND.t2085 630.62
R1129 VGND.t2083 VGND.t1673 630.62
R1130 VGND.t586 VGND.t480 630.62
R1131 VGND.t478 VGND.t850 630.62
R1132 VGND.t461 VGND.t2087 630.62
R1133 VGND.t1275 VGND.t1808 630.62
R1134 VGND.t1239 VGND.t1273 630.62
R1135 VGND.t1108 VGND.t1988 630.62
R1136 VGND.t1106 VGND.t2557 630.62
R1137 VGND.t175 VGND.t1104 630.62
R1138 VGND.t476 VGND.t2638 630.62
R1139 VGND.t1153 VGND.t2527 630.62
R1140 VGND.t1605 VGND.t768 630.62
R1141 VGND.t1801 VGND.t555 630.62
R1142 VGND.t1238 VGND.t1409 630.62
R1143 VGND.t2525 VGND.t259 630.62
R1144 VGND.t1086 VGND.t764 630.62
R1145 VGND.t762 VGND.t567 630.62
R1146 VGND.t673 VGND.t2523 630.62
R1147 VGND.t2521 VGND.t214 630.62
R1148 VGND.t2541 VGND.t766 630.62
R1149 VGND.t1407 VGND.t1320 630.62
R1150 VGND.t2426 VGND.t1405 630.62
R1151 VGND.t760 VGND.t911 630.62
R1152 VGND.t361 VGND.t758 630.62
R1153 VGND.t515 VGND.t1803 630.62
R1154 VGND.t2519 VGND.t2158 630.62
R1155 VGND.t756 VGND.t1783 630.62
R1156 VGND.t588 VGND.t1773 630.62
R1157 VGND.t876 VGND.t524 630.62
R1158 VGND.t874 VGND.t1550 630.62
R1159 VGND.t1781 VGND.t1770 630.62
R1160 VGND.t1231 VGND.t302 630.62
R1161 VGND.t1229 VGND.t541 630.62
R1162 VGND.t1779 VGND.t14 630.62
R1163 VGND.t1777 VGND.t386 630.62
R1164 VGND.t1233 VGND.t158 630.62
R1165 VGND.t872 VGND.t711 630.62
R1166 VGND.t870 VGND.t1345 630.62
R1167 VGND.t1227 VGND.t1994 630.62
R1168 VGND.t880 VGND.t1375 630.62
R1169 VGND.t285 VGND.t878 630.62
R1170 VGND.t1775 VGND.t2112 630.62
R1171 VGND.t1164 VGND.t1493 630.62
R1172 VGND.t1831 VGND.t2553 630.62
R1173 VGND.t552 VGND.t377 630.62
R1174 VGND.t1558 VGND.t1499 630.62
R1175 VGND.t1314 VGND.t1491 630.62
R1176 VGND.t1093 VGND.t2549 630.62
R1177 VGND.t549 VGND.t2547 630.62
R1178 VGND.t315 VGND.t1489 630.62
R1179 VGND.t597 VGND.t1487 630.62
R1180 VGND.t1212 VGND.t2551 630.62
R1181 VGND.t1266 VGND.t1497 630.62
R1182 VGND.t1226 VGND.t1495 630.62
R1183 VGND.t2545 VGND.t2681 630.62
R1184 VGND.t381 VGND.t451 630.62
R1185 VGND.t293 VGND.t379 630.62
R1186 VGND.t1485 VGND.t2138 630.62
R1187 VGND.t652 VGND.t577 630.62
R1188 VGND.t847 VGND.t1903 630.62
R1189 VGND.t583 VGND.t893 630.62
R1190 VGND.t4 VGND.t891 630.62
R1191 VGND.t650 VGND.t1304 630.62
R1192 VGND.t327 VGND.t1100 630.62
R1193 VGND.t1098 VGND.t1674 630.62
R1194 VGND.t587 VGND.t648 630.62
R1195 VGND.t776 VGND.t851 630.62
R1196 VGND.t153 VGND.t1901 630.62
R1197 VGND.t889 VGND.t1809 630.62
R1198 VGND.t1240 VGND.t654 630.62
R1199 VGND.t1096 VGND.t1989 630.62
R1200 VGND.t2558 VGND.t1094 630.62
R1201 VGND.t176 VGND.t895 630.62
R1202 VGND.t774 VGND.t2640 630.62
R1203 VGND.t834 VGND.t311 630.62
R1204 VGND.t845 VGND.t2401 630.62
R1205 VGND.t899 VGND.t582 630.62
R1206 VGND.t1445 VGND.t1335 630.62
R1207 VGND.t1752 VGND.t309 630.62
R1208 VGND.t324 VGND.t2397 630.62
R1209 VGND.t1672 VGND.t2395 630.62
R1210 VGND.t585 VGND.t307 630.62
R1211 VGND.t849 VGND.t305 630.62
R1212 VGND.t460 VGND.t2399 630.62
R1213 VGND.t1807 VGND.t1333 630.62
R1214 VGND.t1575 VGND.t1331 630.62
R1215 VGND.t2393 VGND.t1263 630.62
R1216 VGND.t903 VGND.t2556 630.62
R1217 VGND.t173 VGND.t901 630.62
R1218 VGND.t2529 VGND.t2631 630.62
R1219 VGND.t1152 VGND.t1768 630.62
R1220 VGND.t1705 VGND.t1758 630.62
R1221 VGND.t152 VGND.t1712 630.62
R1222 VGND.t1237 VGND.t1710 630.62
R1223 VGND.t258 VGND.t1766 630.62
R1224 VGND.t1085 VGND.t1754 630.62
R1225 VGND.t566 VGND.t126 630.62
R1226 VGND.t672 VGND.t1764 630.62
R1227 VGND.t729 VGND.t1762 630.62
R1228 VGND.t1215 VGND.t1756 630.62
R1229 VGND.t1319 VGND.t1708 630.62
R1230 VGND.t2423 VGND.t1706 630.62
R1231 VGND.t124 VGND.t2686 630.62
R1232 VGND.t122 VGND.t464 630.62
R1233 VGND.t514 VGND.t120 630.62
R1234 VGND.t1760 VGND.t2153 630.62
R1235 VGND.t813 VGND.t1151 630.62
R1236 VGND.t399 VGND.t370 630.62
R1237 VGND.t821 VGND.t113 630.62
R1238 VGND.t785 VGND.t819 630.62
R1239 VGND.t1702 VGND.t811 630.62
R1240 VGND.t735 VGND.t395 630.62
R1241 VGND.t1666 VGND.t393 630.62
R1242 VGND.t330 VGND.t405 630.62
R1243 VGND.t1838 VGND.t403 630.62
R1244 VGND.t458 VGND.t397 630.62
R1245 VGND.t1749 VGND.t817 630.62
R1246 VGND.t815 VGND.t1617 630.62
R1247 VGND.t391 VGND.t1257 630.62
R1248 VGND.t389 VGND.t34 630.62
R1249 VGND.t823 VGND.t168 630.62
R1250 VGND.t401 VGND.t2590 630.62
R1251 VGND.t1158 VGND.t423 630.62
R1252 VGND.t590 VGND.t2412 630.62
R1253 VGND.t526 VGND.t1568 630.62
R1254 VGND.t429 VGND.t1556 630.62
R1255 VGND.t1772 VGND.t421 630.62
R1256 VGND.t2408 VGND.t1091 630.62
R1257 VGND.t543 VGND.t2406 630.62
R1258 VGND.t419 VGND.t16 630.62
R1259 VGND.t1583 VGND.t417 630.62
R1260 VGND.t1210 VGND.t2410 630.62
R1261 VGND.t427 VGND.t713 630.62
R1262 VGND.t425 VGND.t1224 630.62
R1263 VGND.t1996 VGND.t2404 630.62
R1264 VGND.t1355 VGND.t1572 630.62
R1265 VGND.t291 VGND.t1570 630.62
R1266 VGND.t2414 VGND.t2132 630.62
R1267 VGND.t2449 VGND.t1150 630.62
R1268 VGND.t369 VGND.t742 630.62
R1269 VGND.t612 VGND.t116 630.62
R1270 VGND.t784 VGND.t610 630.62
R1271 VGND.t750 VGND.t1701 630.62
R1272 VGND.t734 VGND.t738 630.62
R1273 VGND.t620 VGND.t138 630.62
R1274 VGND.t644 VGND.t748 630.62
R1275 VGND.t746 VGND.t1837 630.62
R1276 VGND.t455 VGND.t740 630.62
R1277 VGND.t2453 VGND.t1748 630.62
R1278 VGND.t2451 VGND.t1614 630.62
R1279 VGND.t618 VGND.t1256 630.62
R1280 VGND.t616 VGND.t31 630.62
R1281 VGND.t167 VGND.t614 630.62
R1282 VGND.t744 VGND.t2587 630.62
R1283 VGND.t77 VGND.t197 630.62
R1284 VGND.t2445 VGND.t1610 630.62
R1285 VGND.t810 VGND.t682 630.62
R1286 VGND.t1541 VGND.t48 630.62
R1287 VGND.t1820 VGND.t195 630.62
R1288 VGND.t1087 VGND.t2441 630.62
R1289 VGND.t572 VGND.t2439 630.62
R1290 VGND.t678 VGND.t193 630.62
R1291 VGND.t219 VGND.t191 630.62
R1292 VGND.t2443 VGND.t2542 630.62
R1293 VGND.t201 VGND.t1321 630.62
R1294 VGND.t2427 VGND.t199 630.62
R1295 VGND.t916 VGND.t2437 630.62
R1296 VGND.t2435 VGND.t362 630.62
R1297 VGND.t684 VGND.t2428 630.62
R1298 VGND.t2447 VGND.t2173 630.62
R1299 VGND.t835 VGND.t862 630.62
R1300 VGND.t844 VGND.t273 630.62
R1301 VGND.t581 VGND.t1422 630.62
R1302 VGND.t868 VGND.t1444 630.62
R1303 VGND.t856 VGND.t1753 630.62
R1304 VGND.t269 VGND.t325 630.62
R1305 VGND.t267 VGND.t1671 630.62
R1306 VGND.t854 VGND.t584 630.62
R1307 VGND.t852 VGND.t848 630.62
R1308 VGND.t459 VGND.t271 630.62
R1309 VGND.t657 VGND.t866 630.62
R1310 VGND.t1574 VGND.t864 630.62
R1311 VGND.t1262 VGND.t265 630.62
R1312 VGND.t1426 VGND.t2555 630.62
R1313 VGND.t174 VGND.t1424 630.62
R1314 VGND.t723 VGND.t2630 630.62
R1315 VGND.t2669 VGND.t624 630.62
R1316 VGND.t1986 VGND.t2588 630.62
R1317 VGND.t112 VGND.t2163 630.62
R1318 VGND.t1545 VGND.t2141 630.62
R1319 VGND.t1828 VGND.t2658 630.62
R1320 VGND.t696 VGND.t2223 630.62
R1321 VGND.t133 VGND.t2212 630.62
R1322 VGND.t341 VGND.t2654 630.62
R1323 VGND.t670 VGND.t2636 630.62
R1324 VGND.t439 VGND.t2225 630.62
R1325 VGND.t1130 VGND.t1511 630.62
R1326 VGND.t190 VGND.t2133 630.62
R1327 VGND.t924 VGND.t2207 630.62
R1328 VGND.t224 VGND.t2194 630.62
R1329 VGND.t2432 VGND.t2169 630.62
R1330 VGND.t2615 VGND.t2198 630.62
R1331 VGND.n2704 VGND.n327 615.385
R1332 VGND.n2349 VGND.t303 602.708
R1333 VGND.n3019 VGND.t303 602.708
R1334 VGND.n3011 VGND.n3010 599.125
R1335 VGND.n194 VGND.n193 599.125
R1336 VGND.n66 VGND.n65 599.125
R1337 VGND.n117 VGND.n116 599.125
R1338 VGND.n134 VGND.n133 599.125
R1339 VGND.n165 VGND.n164 599.125
R1340 VGND.n2210 VGND.n2182 599.125
R1341 VGND.n2972 VGND.n2971 599.125
R1342 VGND VGND.t383 581.61
R1343 VGND.t96 VGND 573.181
R1344 VGND VGND.t1360 573.181
R1345 VGND.t344 VGND 573.181
R1346 VGND.t375 VGND 573.181
R1347 VGND.n3013 VGND 564.751
R1348 VGND.t1247 VGND 564.751
R1349 VGND.n3014 VGND 564.751
R1350 VGND.n3012 VGND 556.322
R1351 VGND.t2539 VGND 539.465
R1352 VGND VGND.t1178 539.465
R1353 VGND.t632 VGND.n806 494.779
R1354 VGND.n1166 VGND.t2190 492.058
R1355 VGND.t2128 VGND.n1175 492.058
R1356 VGND.n1176 VGND.t2104 492.058
R1357 VGND.t2188 VGND.n1188 492.058
R1358 VGND.n1189 VGND.t2176 492.058
R1359 VGND.t2154 VGND.n1207 492.058
R1360 VGND.n1208 VGND.t2601 492.058
R1361 VGND.t2581 VGND.n1220 492.058
R1362 VGND.n1247 VGND.t2149 492.058
R1363 VGND.n1246 VGND.t2656 492.058
R1364 VGND.n1240 VGND.t2645 492.058
R1365 VGND.n1239 VGND.t2210 492.058
R1366 VGND.n1233 VGND.t2139 492.058
R1367 VGND.t2634 VGND.n1277 492.058
R1368 VGND.n1278 VGND.t2221 492.058
R1369 VGND.t2346 VGND.t2305 481.877
R1370 VGND.t2380 VGND.t2346 481.877
R1371 VGND.t1475 VGND.t1446 481.877
R1372 VGND.t1446 VGND.t1139 481.877
R1373 VGND.t1846 VGND 452.382
R1374 VGND.n1166 VGND.t93 424.312
R1375 VGND.n1175 VGND.t1596 424.312
R1376 VGND.n1176 VGND.t1530 424.312
R1377 VGND.n1188 VGND.t671 424.312
R1378 VGND.n1189 VGND.t1110 424.312
R1379 VGND.n1207 VGND.t1131 424.312
R1380 VGND.n1208 VGND.t29 424.312
R1381 VGND.n1220 VGND.t237 424.312
R1382 VGND.n1247 VGND.t662 424.312
R1383 VGND.t226 VGND.n1246 424.312
R1384 VGND.n1240 VGND.t563 424.312
R1385 VGND.t680 VGND.n1239 424.312
R1386 VGND.n1233 VGND.t1338 424.312
R1387 VGND.n1277 VGND.t229 424.312
R1388 VGND.n1278 VGND.t467 424.312
R1389 VGND.t727 VGND.n222 424.312
R1390 VGND.t141 VGND 419.68
R1391 VGND.n2284 VGND.n503 413.043
R1392 VGND.t982 VGND.t1401 408.469
R1393 VGND.t2068 VGND.t1156 408.469
R1394 VGND.t800 VGND.t1608 408.469
R1395 VGND.t1939 VGND.t556 408.469
R1396 VGND.t1634 VGND.t1554 408.469
R1397 VGND.t2495 VGND.t262 408.469
R1398 VGND.t1935 VGND.t732 408.469
R1399 VGND.t1662 VGND.t570 408.469
R1400 VGND.t676 VGND.t1953 408.469
R1401 VGND.t2277 VGND.t217 408.469
R1402 VGND.t1216 VGND.t1691 408.469
R1403 VGND.t2481 VGND.t1746 408.469
R1404 VGND.t2424 VGND.t2269 408.469
R1405 VGND.t914 VGND.t54 408.469
R1406 VGND.t1917 VGND.t465 408.469
R1407 VGND.t289 VGND.t1865 408.469
R1408 VGND.t1057 VGND.t1301 408.469
R1409 VGND.t832 VGND.t2241 408.469
R1410 VGND.t373 VGND.t1734 408.469
R1411 VGND.t114 VGND.t1385 408.469
R1412 VGND.t1546 VGND.t2070 408.469
R1413 VGND.t1750 VGND.t2461 408.469
R1414 VGND.t300 VGND.t1381 408.469
R1415 VGND.t1669 VGND.t1636 408.469
R1416 VGND.t333 VGND.t2497 408.469
R1417 VGND.t1841 VGND.t1937 408.469
R1418 VGND.t456 VGND.t1971 408.469
R1419 VGND.t709 VGND.t2038 408.469
R1420 VGND.t1615 VGND.t2024 408.469
R1421 VGND.t1260 VGND.t1695 408.469
R1422 VGND.t32 VGND.t1867 408.469
R1423 VGND.t2433 VGND.t2271 408.469
R1424 VGND.t2491 VGND.t964 408.469
R1425 VGND.t81 VGND.t2016 408.469
R1426 VGND.t1687 VGND.t1982 408.469
R1427 VGND.t605 VGND.t1925 408.469
R1428 VGND.t2261 VGND.t1561 408.469
R1429 VGND.t1824 VGND.t494 408.469
R1430 VGND.t1913 VGND.t320 408.469
R1431 VGND.t129 VGND.t1857 408.469
R1432 VGND.t1285 VGND.t337 408.469
R1433 VGND.t666 VGND.t2056 408.469
R1434 VGND.t1714 VGND.t434 408.469
R1435 VGND.t1740 VGND.t1279 408.469
R1436 VGND.t804 VGND.t185 408.469
R1437 VGND.t2467 VGND.t920 408.469
R1438 VGND.t1644 VGND.t365 408.469
R1439 VGND.t510 VGND.t1618 408.469
R1440 VGND.t1006 VGND.t2046 408.469
R1441 VGND.t1654 VGND.t836 408.469
R1442 VGND.t1832 VGND.t1965 408.469
R1443 VGND.t1873 VGND.t529 408.469
R1444 VGND.t9 VGND.t2018 408.469
R1445 VGND.t2255 VGND.t1315 408.469
R1446 VGND.t692 VGND.t1859 408.469
R1447 VGND.t2263 VGND.t550 408.469
R1448 VGND.t316 VGND.t496 408.469
R1449 VGND.t1915 VGND.t598 408.469
R1450 VGND.t164 VGND.t1879 408.469
R1451 VGND.t488 VGND.t1126 408.469
R1452 VGND.t1220 VGND.t1907 408.469
R1453 VGND.t2682 VGND.t1718 408.469
R1454 VGND.t1620 VGND.t1351 408.469
R1455 VGND.t281 VGND.t2052 408.469
R1456 VGND.t2455 VGND.t1078 408.469
R1457 VGND.t1628 VGND.t1148 408.469
R1458 VGND.t2677 VGND.t2507 408.469
R1459 VGND.t2281 VGND.t108 408.469
R1460 VGND.t1539 VGND.t1656 408.469
R1461 VGND.t2487 VGND.t1699 408.469
R1462 VGND.t296 VGND.t2265 408.469
R1463 VGND.t2020 VGND.t136 408.469
R1464 VGND.t642 VGND.t1675 408.469
R1465 VGND.t1861 VGND.t1137 408.469
R1466 VGND.t442 VGND.t52 408.469
R1467 VGND.t2247 VGND.t1812 408.469
R1468 VGND.t2421 VGND.t1855 408.469
R1469 VGND.t1881 VGND.t1254 408.469
R1470 VGND.t2054 VGND.t24 408.469
R1471 VGND.t518 VGND.t1911 408.469
R1472 VGND.t1391 VGND.t985 408.469
R1473 VGND.t2060 VGND.t1154 408.469
R1474 VGND.t1606 VGND.t790 408.469
R1475 VGND.t553 VGND.t1929 408.469
R1476 VGND.t1552 VGND.t1624 408.469
R1477 VGND.t260 VGND.t2030 408.469
R1478 VGND.t730 VGND.t2012 408.469
R1479 VGND.t568 VGND.t1650 408.469
R1480 VGND.t674 VGND.t2475 408.469
R1481 VGND.t215 VGND.t72 408.469
R1482 VGND.t1213 VGND.t1679 408.469
R1483 VGND.t1744 VGND.t2469 408.469
R1484 VGND.t1218 VGND.t68 408.469
R1485 VGND.t912 VGND.t504 408.469
R1486 VGND.t1905 VGND.t462 408.469
R1487 VGND.t287 VGND.t1897 408.469
R1488 VGND.t1291 VGND.t958 408.469
R1489 VGND.t1923 VGND.t622 408.469
R1490 VGND.t1722 VGND.t1984 408.469
R1491 VGND.t1660 VGND.t603 408.469
R1492 VGND.t2062 VGND.t1235 408.469
R1493 VGND.t1945 VGND.t1826 408.469
R1494 VGND.t1652 VGND.t322 408.469
R1495 VGND.t1626 VGND.t131 408.469
R1496 VGND.t2036 VGND.t339 408.469
R1497 VGND.t2014 VGND.t668 408.469
R1498 VGND.t1959 VGND.t436 408.469
R1499 VGND.t2026 VGND.t1742 408.469
R1500 VGND.t187 VGND.t2010 408.469
R1501 VGND.t922 VGND.t1681 408.469
R1502 VGND.t1899 VGND.t367 408.469
R1503 VGND.t512 VGND.t70 408.469
R1504 VGND.t1000 VGND.t2473 408.469
R1505 VGND.t2004 VGND.t838 408.469
R1506 VGND.t1677 VGND.t1834 408.469
R1507 VGND.t1909 VGND.t527 408.469
R1508 VGND.t11 VGND.t60 408.469
R1509 VGND.t484 VGND.t1599 408.469
R1510 VGND.t694 VGND.t1728 408.469
R1511 VGND.t1891 VGND.t564 408.469
R1512 VGND.t318 VGND.t1640 408.469
R1513 VGND.t798 VGND.t600 408.469
R1514 VGND.t1208 VGND.t1397 408.469
R1515 VGND.t1630 VGND.t1128 408.469
R1516 VGND.t1222 VGND.t792 408.469
R1517 VGND.t2459 VGND.t2684 408.469
R1518 VGND.t1967 VGND.t1353 408.469
R1519 VGND.t283 VGND.t2509 408.469
R1520 VGND.t2028 VGND.t1012 408.469
R1521 VGND.t1646 VGND.t1160 408.469
R1522 VGND.t591 VGND.t1957 408.469
R1523 VGND.t1853 VGND.t533 408.469
R1524 VGND.t2006 VGND.t5 408.469
R1525 VGND.t2243 VGND.t1309 408.469
R1526 VGND.t1893 VGND.t690 408.469
R1527 VGND.t62 VGND.t546 408.469
R1528 VGND.t486 VGND.t19 408.469
R1529 VGND.t1732 VGND.t1586 408.469
R1530 VGND.t1295 VGND.t162 408.469
R1531 VGND.t2066 VGND.t1124 408.469
R1532 VGND.t1349 VGND.t1724 408.469
R1533 VGND.t1999 VGND.t1399 408.469
R1534 VGND.t2511 VGND.t1377 408.469
R1535 VGND.t179 VGND.t794 408.469
R1536 VGND.t1943 VGND.t940 408.469
R1537 VGND.t1622 VGND.t1146 408.469
R1538 VGND.t2505 VGND.t2675 408.469
R1539 VGND.t2259 VGND.t110 408.469
R1540 VGND.t1648 VGND.t1537 408.469
R1541 VGND.t2471 VGND.t1977 408.469
R1542 VGND.t64 VGND.t328 408.469
R1543 VGND.t2008 VGND.t134 408.469
R1544 VGND.t2245 VGND.t640 408.469
R1545 VGND.t1895 VGND.t1135 408.469
R1546 VGND.t502 VGND.t440 408.469
R1547 VGND.t2237 VGND.t1810 408.469
R1548 VGND.t2419 VGND.t1889 408.469
R1549 VGND.t1252 VGND.t1297 408.469
R1550 VGND.t796 VGND.t22 408.469
R1551 VGND.t516 VGND.t1726 408.469
R1552 VGND.t1036 VGND.t1299 408.469
R1553 VGND.t754 VGND.t2235 408.469
R1554 VGND.t1603 VGND.t1730 408.469
R1555 VGND.t1383 VGND.t520 408.469
R1556 VGND.t2064 VGND.t1442 408.469
R1557 VGND.t2457 VGND.t1307 408.469
R1558 VGND.t1658 VGND.t1083 408.469
R1559 VGND.t1632 VGND.t539 408.469
R1560 VGND.t2048 VGND.t721 408.469
R1561 VGND.t1931 VGND.t210 408.469
R1562 VGND.t1969 VGND.t156 408.469
R1563 VGND.t1317 VGND.t2032 408.469
R1564 VGND.t1243 VGND.t2022 408.469
R1565 VGND.t1992 VGND.t1689 408.469
R1566 VGND.t1535 VGND.t1863 408.469
R1567 VGND.t171 VGND.t2267 408.469
R1568 VGND.t1941 VGND.t967 408.469
R1569 VGND.t2515 VGND.t79 408.469
R1570 VGND.t2501 VGND.t1980 408.469
R1571 VGND.t808 VGND.t66 408.469
R1572 VGND.t1642 VGND.t1559 408.469
R1573 VGND.t1822 VGND.t1875 408.469
R1574 VGND.t58 VGND.t736 408.469
R1575 VGND.t574 VGND.t2002 408.469
R1576 VGND.t2239 VGND.t335 408.469
R1577 VGND.t1887 VGND.t664 408.469
R1578 VGND.t2543 VGND.t498 408.469
R1579 VGND.t1738 VGND.t1927 408.469
R1580 VGND.t1885 VGND.t183 408.469
R1581 VGND.t1287 VGND.t918 408.469
R1582 VGND.t788 VGND.t363 408.469
R1583 VGND.t508 VGND.t1720 408.469
R1584 VGND.t1039 VGND.t2517 408.469
R1585 VGND.t1389 VGND.t752 408.469
R1586 VGND.t1601 VGND.t1664 408.469
R1587 VGND.t1955 VGND.t522 408.469
R1588 VGND.t1440 VGND.t1947 408.469
R1589 VGND.t1693 VGND.t1305 408.469
R1590 VGND.t1081 VGND.t2485 408.469
R1591 VGND.t2040 VGND.t537 408.469
R1592 VGND.t719 VGND.t56 408.469
R1593 VGND.t2257 VGND.t208 408.469
R1594 VGND.t154 VGND.t1869 408.469
R1595 VGND.t1267 VGND.t506 408.469
R1596 VGND.t1241 VGND.t2249 408.469
R1597 VGND.t1990 VGND.t1921 408.469
R1598 VGND.t1281 VGND.t1533 408.469
R1599 VGND.t169 VGND.t490 408.469
R1600 VGND.t802 VGND.t1069 408.469
R1601 VGND.t830 VGND.t1289 408.469
R1602 VGND.t1638 VGND.t371 408.469
R1603 VGND.t2499 VGND.t578 408.469
R1604 VGND.t1393 VGND.t1543 408.469
R1605 VGND.t1973 VGND.t1703 408.469
R1606 VGND.t2042 VGND.t298 408.469
R1607 VGND.t1949 VGND.t1667 408.469
R1608 VGND.t1697 VGND.t331 408.469
R1609 VGND.t1839 VGND.t2489 408.469
R1610 VGND.t453 VGND.t2273 408.469
R1611 VGND.t1685 VGND.t707 408.469
R1612 VGND.t2477 VGND.t1612 408.469
R1613 VGND.t1258 VGND.t1871 408.469
R1614 VGND.t26 VGND.t492 408.469
R1615 VGND.t2430 VGND.t2251 408.469
R1616 VGND.t1736 VGND.t1009 408.469
R1617 VGND.t500 VGND.t1162 408.469
R1618 VGND.t2072 VGND.t593 408.469
R1619 VGND.t531 VGND.t2463 408.469
R1620 VGND.t7 VGND.t1293 408.469
R1621 VGND.t1311 VGND.t2513 408.469
R1622 VGND.t432 VGND.t1951 408.469
R1623 VGND.t544 VGND.t1395 408.469
R1624 VGND.t17 VGND.t1975 408.469
R1625 VGND.t2044 VGND.t1584 408.469
R1626 VGND.t1933 VGND.t160 408.469
R1627 VGND.t1963 VGND.t1122 408.469
R1628 VGND.t2034 VGND.t1347 408.469
R1629 VGND.t1997 VGND.t2275 408.469
R1630 VGND.t2253 VGND.t1379 408.469
R1631 VGND.t177 VGND.t2479 408.469
R1632 VGND.t2160 VGND.t2279 408.469
R1633 VGND.t1961 VGND.t2667 408.469
R1634 VGND.t2483 VGND.t2585 408.469
R1635 VGND.t1883 VGND.t2217 408.469
R1636 VGND.t1683 VGND.t2662 408.469
R1637 VGND.t1919 VGND.t2651 408.469
R1638 VGND.t1877 VGND.t2632 408.469
R1639 VGND.t50 VGND.t2145 408.469
R1640 VGND.t2058 VGND.t1507 408.469
R1641 VGND.t1716 VGND.t2628 408.469
R1642 VGND.t1283 VGND.t2205 408.469
R1643 VGND.t2050 VGND.t2192 408.469
R1644 VGND.t1403 VGND.t2117 408.469
R1645 VGND.t1387 VGND.t2611 408.469
R1646 VGND.t2503 VGND.t2174 408.469
R1647 VGND.t2126 VGND.t2465 408.469
R1648 VGND.t2378 VGND.t2297 397.848
R1649 VGND.t2297 VGND.t2307 397.848
R1650 VGND.t2307 VGND.t2315 397.848
R1651 VGND.t2315 VGND.t1362 397.848
R1652 VGND.t1362 VGND.t1363 397.848
R1653 VGND.t1363 VGND.t1366 397.848
R1654 VGND.t1366 VGND.t1367 397.848
R1655 VGND.t2283 VGND.t1589 396.17
R1656 VGND.t786 VGND.t1815 396.17
R1657 VGND.n2935 VGND.n2934 394.137
R1658 VGND.n2933 VGND.n208 394.137
R1659 VGND.n2932 VGND.n209 394.137
R1660 VGND.n2931 VGND.n210 394.137
R1661 VGND.n2930 VGND.n211 394.137
R1662 VGND.n2929 VGND.n212 394.137
R1663 VGND.n2928 VGND.n213 394.137
R1664 VGND.n2927 VGND.n214 394.137
R1665 VGND.n2926 VGND.n215 394.137
R1666 VGND.n2925 VGND.n216 394.137
R1667 VGND.n2924 VGND.n217 394.137
R1668 VGND.n2923 VGND.n218 394.137
R1669 VGND.n2922 VGND.n219 394.137
R1670 VGND.n2921 VGND.n220 394.137
R1671 VGND.n2920 VGND.n221 394.137
R1672 VGND.n2919 VGND.n2918 394.137
R1673 VGND.n2285 VGND.t45 387.421
R1674 VGND.n2284 VGND.t413 387.421
R1675 VGND.n2250 VGND.t35 387.421
R1676 VGND.n2248 VGND.t410 387.421
R1677 VGND.n1386 VGND.t39 387.421
R1678 VGND.t1816 VGND.t806 362.452
R1679 VGND.t806 VGND.t2539 345.594
R1680 VGND VGND.t88 328.616
R1681 VGND VGND.t37 328.616
R1682 VGND VGND.t142 328.616
R1683 VGND VGND.t87 328.616
R1684 VGND VGND.t250 328.616
R1685 VGND.t2136 VGND.t2196 313.776
R1686 VGND.t2130 VGND.t2625 313.776
R1687 VGND.t2610 VGND.t2617 313.776
R1688 VGND.t2595 VGND.t2172 313.776
R1689 VGND.t2124 VGND.t2184 313.776
R1690 VGND.t2108 VGND.t2598 313.776
R1691 VGND.t2187 VGND.t2664 313.776
R1692 VGND.t2178 VGND.t2162 313.776
R1693 VGND.t2666 VGND.t2156 313.776
R1694 VGND.t2110 VGND.t2599 313.776
R1695 VGND.t2159 VGND.t2583 313.776
R1696 VGND.t2228 VGND.t2147 313.776
R1697 VGND.t2653 VGND.t2660 313.776
R1698 VGND.t2648 VGND.t2230 313.776
R1699 VGND.t2209 VGND.t2626 313.776
R1700 VGND.t2143 VGND.t2650 313.776
R1701 VGND.t2292 VGND.t2283 311.877
R1702 VGND.t383 VGND.t786 311.877
R1703 VGND VGND.t2288 303.449
R1704 VGND VGND.t2292 295.019
R1705 VGND.n101 VGND.t2306 287.832
R1706 VGND VGND.t1173 286.591
R1707 VGND.n93 VGND.t2331 282.327
R1708 VGND.n2184 VGND.t1469 282.327
R1709 VGND.n104 VGND.t2377 281.13
R1710 VGND.n2189 VGND.t43 281.13
R1711 VGND.n177 VGND.t2322 280.978
R1712 VGND.n177 VGND.t2363 280.978
R1713 VGND.n78 VGND.t2373 280.978
R1714 VGND.n78 VGND.t2389 280.978
R1715 VGND.n146 VGND.t2349 280.978
R1716 VGND.n146 VGND.t2385 280.978
R1717 VGND.n482 VGND.t635 280.978
R1718 VGND.n482 VGND.t1466 280.978
R1719 VGND.n2263 VGND.t44 280.978
R1720 VGND.n2263 VGND.t416 280.978
R1721 VGND.n518 VGND.t1474 280.978
R1722 VGND.n518 VGND.t1463 280.978
R1723 VGND.n2194 VGND.t1140 280.978
R1724 VGND.t2079 VGND 278.161
R1725 VGND.n2970 VGND 271.014
R1726 VGND.n3021 VGND.n4 259.389
R1727 VGND.n2347 VGND.n4 259.389
R1728 VGND.n3022 VGND.n3 252.988
R1729 VGND VGND.t2317 252.875
R1730 VGND VGND.t2290 252.875
R1731 VGND VGND.t2285 252.875
R1732 VGND VGND.t2313 252.875
R1733 VGND.t2365 VGND 252.875
R1734 VGND.n887 VGND.t2280 241.393
R1735 VGND.n330 VGND.t995 241.393
R1736 VGND.n396 VGND.t1402 241.393
R1737 VGND.n400 VGND.t1302 241.393
R1738 VGND.n469 VGND.t2492 241.393
R1739 VGND.n466 VGND.t2047 241.393
R1740 VGND.n625 VGND.t2456 241.393
R1741 VGND.n590 VGND.t1392 241.393
R1742 VGND.n587 VGND.t1292 241.393
R1743 VGND.n547 VGND.t2474 241.393
R1744 VGND.n628 VGND.t2029 241.393
R1745 VGND.n632 VGND.t1944 241.393
R1746 VGND.n879 VGND.t1300 241.393
R1747 VGND.n800 VGND.t1942 241.393
R1748 VGND.n797 VGND.t2518 241.393
R1749 VGND.n882 VGND.t803 241.393
R1750 VGND.n1024 VGND.t1737 241.393
R1751 VGND.n1014 VGND.t998 241.393
R1752 VGND.n1333 VGND.t1962 241.284
R1753 VGND.n894 VGND.t2484 241.284
R1754 VGND.n932 VGND.t1884 241.284
R1755 VGND.n937 VGND.t1684 241.284
R1756 VGND.n942 VGND.t1920 241.284
R1757 VGND.n947 VGND.t1878 241.284
R1758 VGND.n952 VGND.t51 241.284
R1759 VGND.n957 VGND.t2059 241.284
R1760 VGND.n962 VGND.t1717 241.284
R1761 VGND.n967 VGND.t1284 241.284
R1762 VGND.n972 VGND.t2051 241.284
R1763 VGND.n977 VGND.t1404 241.284
R1764 VGND.n982 VGND.t1388 241.284
R1765 VGND.n987 VGND.t2504 241.284
R1766 VGND.n1280 VGND.t1034 241.284
R1767 VGND.n1275 VGND.t992 241.284
R1768 VGND.n1232 VGND.t1076 241.284
R1769 VGND.n1237 VGND.t1067 241.284
R1770 VGND.n1225 VGND.t1028 241.284
R1771 VGND.n1244 VGND.t980 241.284
R1772 VGND.n1001 VGND.t1064 241.284
R1773 VGND.n1218 VGND.t1025 241.284
R1774 VGND.n1210 VGND.t1016 241.284
R1775 VGND.n1205 VGND.t974 241.284
R1776 VGND.n1009 VGND.t1052 241.284
R1777 VGND.n1186 VGND.t1046 241.284
R1778 VGND.n1178 VGND.t971 241.284
R1779 VGND.n1173 VGND.t953 241.284
R1780 VGND.n1168 VGND.t947 241.284
R1781 VGND.n2773 VGND.t1031 241.284
R1782 VGND.n294 VGND.t989 241.284
R1783 VGND.n2730 VGND.t1073 241.284
R1784 VGND.n2735 VGND.t1061 241.284
R1785 VGND.n312 VGND.t1022 241.284
R1786 VGND.n2726 VGND.t977 241.284
R1787 VGND.n326 VGND.t1055 241.284
R1788 VGND.n387 VGND.t1019 241.284
R1789 VGND.n384 VGND.t1004 241.284
R1790 VGND.n379 VGND.t962 241.284
R1791 VGND.n373 VGND.t1049 241.284
R1792 VGND.n368 VGND.t1043 241.284
R1793 VGND.n362 VGND.t956 241.284
R1794 VGND.n355 VGND.t950 241.284
R1795 VGND.n2699 VGND.t944 241.284
R1796 VGND.n2639 VGND.t2069 241.284
R1797 VGND.n2644 VGND.t801 241.284
R1798 VGND.n2649 VGND.t1940 241.284
R1799 VGND.n2654 VGND.t1635 241.284
R1800 VGND.n2659 VGND.t2496 241.284
R1801 VGND.n2664 VGND.t1936 241.284
R1802 VGND.n2669 VGND.t1663 241.284
R1803 VGND.n394 VGND.t1954 241.284
R1804 VGND.n2715 VGND.t2278 241.284
R1805 VGND.n320 VGND.t1692 241.284
R1806 VGND.n2748 VGND.t2482 241.284
R1807 VGND.n304 VGND.t2270 241.284
R1808 VGND.n2753 VGND.t55 241.284
R1809 VGND.n2788 VGND.t1918 241.284
R1810 VGND.n287 VGND.t1866 241.284
R1811 VGND.n2343 VGND.t2242 241.284
R1812 VGND.n2338 VGND.t1735 241.284
R1813 VGND.n2333 VGND.t1386 241.284
R1814 VGND.n2328 VGND.t2071 241.284
R1815 VGND.n2323 VGND.t2462 241.284
R1816 VGND.n2318 VGND.t1382 241.284
R1817 VGND.n2313 VGND.t1637 241.284
R1818 VGND.n2308 VGND.t2498 241.284
R1819 VGND.n2303 VGND.t1938 241.284
R1820 VGND.n2298 VGND.t1972 241.284
R1821 VGND.n2293 VGND.t2039 241.284
R1822 VGND.n2288 VGND.t2025 241.284
R1823 VGND.n415 VGND.t1696 241.284
R1824 VGND.n2541 VGND.t1868 241.284
R1825 VGND.n2536 VGND.t2272 241.284
R1826 VGND.n472 VGND.t2017 241.284
R1827 VGND.n2377 VGND.t1688 241.284
R1828 VGND.n460 VGND.t1926 241.284
R1829 VGND.n2403 VGND.t2262 241.284
R1830 VGND.n452 VGND.t495 241.284
R1831 VGND.n2429 VGND.t1914 241.284
R1832 VGND.n444 VGND.t1858 241.284
R1833 VGND.n2455 VGND.t1286 241.284
R1834 VGND.n436 VGND.t2057 241.284
R1835 VGND.n2481 VGND.t1715 241.284
R1836 VGND.n428 VGND.t1280 241.284
R1837 VGND.n2512 VGND.t805 241.284
R1838 VGND.n2517 VGND.t2468 241.284
R1839 VGND.n2522 VGND.t1645 241.284
R1840 VGND.n2527 VGND.t1619 241.284
R1841 VGND.n2364 VGND.t1655 241.284
R1842 VGND.n464 VGND.t1966 241.284
R1843 VGND.n2390 VGND.t1874 241.284
R1844 VGND.n456 VGND.t2019 241.284
R1845 VGND.n2416 VGND.t2256 241.284
R1846 VGND.n448 VGND.t1860 241.284
R1847 VGND.n2442 VGND.t2264 241.284
R1848 VGND.n440 VGND.t497 241.284
R1849 VGND.n2468 VGND.t1916 241.284
R1850 VGND.n432 VGND.t1880 241.284
R1851 VGND.n2494 VGND.t489 241.284
R1852 VGND.n424 VGND.t1908 241.284
R1853 VGND.n2499 VGND.t1719 241.284
R1854 VGND.n2810 VGND.t1621 241.284
R1855 VGND.n2815 VGND.t2053 241.284
R1856 VGND.n1911 VGND.t1629 241.284
R1857 VGND.n623 VGND.t2508 241.284
R1858 VGND.n1922 VGND.t2282 241.284
R1859 VGND.n620 VGND.t1657 241.284
R1860 VGND.n1933 VGND.t2488 241.284
R1861 VGND.n617 VGND.t2266 241.284
R1862 VGND.n1944 VGND.t2021 241.284
R1863 VGND.n614 VGND.t1676 241.284
R1864 VGND.n1955 VGND.t1862 241.284
R1865 VGND.n611 VGND.t53 241.284
R1866 VGND.n1966 VGND.t2248 241.284
R1867 VGND.n608 VGND.t1856 241.284
R1868 VGND.n1977 VGND.t1882 241.284
R1869 VGND.n1982 VGND.t2055 241.284
R1870 VGND.n1987 VGND.t1912 241.284
R1871 VGND.n597 VGND.t2061 241.284
R1872 VGND.n594 VGND.t791 241.284
R1873 VGND.n2056 VGND.t1930 241.284
R1874 VGND.n2051 VGND.t1625 241.284
R1875 VGND.n2046 VGND.t2031 241.284
R1876 VGND.n2041 VGND.t2013 241.284
R1877 VGND.n2036 VGND.t1651 241.284
R1878 VGND.n2031 VGND.t2476 241.284
R1879 VGND.n2026 VGND.t73 241.284
R1880 VGND.n2021 VGND.t1680 241.284
R1881 VGND.n2016 VGND.t2470 241.284
R1882 VGND.n2011 VGND.t69 241.284
R1883 VGND.n2006 VGND.t505 241.284
R1884 VGND.n2001 VGND.t1906 241.284
R1885 VGND.n1994 VGND.t1898 241.284
R1886 VGND.n2070 VGND.t1924 241.284
R1887 VGND.n2075 VGND.t1723 241.284
R1888 VGND.n2080 VGND.t1661 241.284
R1889 VGND.n2085 VGND.t2063 241.284
R1890 VGND.n2090 VGND.t1946 241.284
R1891 VGND.n2095 VGND.t1653 241.284
R1892 VGND.n2100 VGND.t1627 241.284
R1893 VGND.n2105 VGND.t2037 241.284
R1894 VGND.n2110 VGND.t2015 241.284
R1895 VGND.n2115 VGND.t1960 241.284
R1896 VGND.n2120 VGND.t2027 241.284
R1897 VGND.n585 VGND.t2011 241.284
R1898 VGND.n2125 VGND.t1682 241.284
R1899 VGND.n2835 VGND.t1900 241.284
R1900 VGND.n2840 VGND.t71 241.284
R1901 VGND.n2177 VGND.t2005 241.284
R1902 VGND.n1756 VGND.t1678 241.284
R1903 VGND.n1762 VGND.t1910 241.284
R1904 VGND.n1753 VGND.t61 241.284
R1905 VGND.n1773 VGND.t485 241.284
R1906 VGND.n1750 VGND.t1729 241.284
R1907 VGND.n1784 VGND.t1892 241.284
R1908 VGND.n1747 VGND.t1641 241.284
R1909 VGND.n1795 VGND.t799 241.284
R1910 VGND.n1744 VGND.t1398 241.284
R1911 VGND.n1806 VGND.t1631 241.284
R1912 VGND.n1741 VGND.t793 241.284
R1913 VGND.n1817 VGND.t2460 241.284
R1914 VGND.n1822 VGND.t1968 241.284
R1915 VGND.n1827 VGND.t2510 241.284
R1916 VGND.n1679 VGND.t1647 241.284
R1917 VGND.n1676 VGND.t1958 241.284
R1918 VGND.n1690 VGND.t1854 241.284
R1919 VGND.n1695 VGND.t2007 241.284
R1920 VGND.n1700 VGND.t2244 241.284
R1921 VGND.n1705 VGND.t1894 241.284
R1922 VGND.n1710 VGND.t63 241.284
R1923 VGND.n1715 VGND.t487 241.284
R1924 VGND.n1720 VGND.t1733 241.284
R1925 VGND.n1725 VGND.t1296 241.284
R1926 VGND.n1730 VGND.t2067 241.284
R1927 VGND.n1673 VGND.t1725 241.284
R1928 VGND.n1846 VGND.t1400 241.284
R1929 VGND.n1841 VGND.t2512 241.284
R1930 VGND.n1834 VGND.t795 241.284
R1931 VGND.n670 VGND.t1623 241.284
R1932 VGND.n675 VGND.t2506 241.284
R1933 VGND.n680 VGND.t2260 241.284
R1934 VGND.n685 VGND.t1649 241.284
R1935 VGND.n690 VGND.t2472 241.284
R1936 VGND.n695 VGND.t65 241.284
R1937 VGND.n700 VGND.t2009 241.284
R1938 VGND.n705 VGND.t2246 241.284
R1939 VGND.n710 VGND.t1896 241.284
R1940 VGND.n715 VGND.t503 241.284
R1941 VGND.n720 VGND.t2238 241.284
R1942 VGND.n667 VGND.t1890 241.284
R1943 VGND.n725 VGND.t1298 241.284
R1944 VGND.n2860 VGND.t797 241.284
R1945 VGND.n2865 VGND.t1727 241.284
R1946 VGND.n1353 VGND.t2236 241.284
R1947 VGND.n875 VGND.t1731 241.284
R1948 VGND.n870 VGND.t1384 241.284
R1949 VGND.n810 VGND.t2065 241.284
R1950 VGND.n824 VGND.t2458 241.284
R1951 VGND.n829 VGND.t1659 241.284
R1952 VGND.n834 VGND.t1633 241.284
R1953 VGND.n839 VGND.t2049 241.284
R1954 VGND.n844 VGND.t1932 241.284
R1955 VGND.n849 VGND.t1970 241.284
R1956 VGND.n820 VGND.t2033 241.284
R1957 VGND.n854 VGND.t2023 241.284
R1958 VGND.n735 VGND.t1690 241.284
R1959 VGND.n1662 VGND.t1864 241.284
R1960 VGND.n1657 VGND.t2268 241.284
R1961 VGND.n1391 VGND.t2516 241.284
R1962 VGND.n1396 VGND.t2502 241.284
R1963 VGND.n805 VGND.t67 241.284
R1964 VGND.n1491 VGND.t1643 241.284
R1965 VGND.n777 VGND.t1876 241.284
R1966 VGND.n1517 VGND.t59 241.284
R1967 VGND.n769 VGND.t2003 241.284
R1968 VGND.n1543 VGND.t2240 241.284
R1969 VGND.n1548 VGND.t1888 241.284
R1970 VGND.n761 VGND.t499 241.284
R1971 VGND.n1553 VGND.t1928 241.284
R1972 VGND.n1633 VGND.t1886 241.284
R1973 VGND.n1638 VGND.t1288 241.284
R1974 VGND.n1643 VGND.t789 241.284
R1975 VGND.n1648 VGND.t1721 241.284
R1976 VGND.n1411 VGND.t1390 241.284
R1977 VGND.n795 VGND.t1665 241.284
R1978 VGND.n1478 VGND.t1956 241.284
R1979 VGND.n781 VGND.t1948 241.284
R1980 VGND.n1504 VGND.t1694 241.284
R1981 VGND.n773 VGND.t2486 241.284
R1982 VGND.n1530 VGND.t2041 241.284
R1983 VGND.n765 VGND.t57 241.284
R1984 VGND.n1567 VGND.t2258 241.284
R1985 VGND.n756 VGND.t1870 241.284
R1986 VGND.n1582 VGND.t507 241.284
R1987 VGND.n1577 VGND.t2250 241.284
R1988 VGND.n1572 VGND.t1922 241.284
R1989 VGND.n2885 VGND.t1282 241.284
R1990 VGND.n2890 VGND.t491 241.284
R1991 VGND.n885 VGND.t1290 241.284
R1992 VGND.n1424 VGND.t1639 241.284
R1993 VGND.n1429 VGND.t2500 241.284
R1994 VGND.n1434 VGND.t1394 241.284
R1995 VGND.n1439 VGND.t1974 241.284
R1996 VGND.n1444 VGND.t2043 241.284
R1997 VGND.n1449 VGND.t1950 241.284
R1998 VGND.n1454 VGND.t1698 241.284
R1999 VGND.n791 VGND.t2490 241.284
R2000 VGND.n1459 VGND.t2274 241.284
R2001 VGND.n1596 VGND.t1686 241.284
R2002 VGND.n1601 VGND.t2478 241.284
R2003 VGND.n750 VGND.t1872 241.284
R2004 VGND.n1614 VGND.t493 241.284
R2005 VGND.n1609 VGND.t2252 241.284
R2006 VGND.n1032 VGND.t501 241.284
R2007 VGND.n1037 VGND.t2073 241.284
R2008 VGND.n1029 VGND.t2464 241.284
R2009 VGND.n1095 VGND.t1294 241.284
R2010 VGND.n1090 VGND.t2514 241.284
R2011 VGND.n1085 VGND.t1952 241.284
R2012 VGND.n1080 VGND.t1396 241.284
R2013 VGND.n1075 VGND.t1976 241.284
R2014 VGND.n1070 VGND.t2045 241.284
R2015 VGND.n1043 VGND.t1934 241.284
R2016 VGND.n1053 VGND.t1964 241.284
R2017 VGND.n1058 VGND.t2035 241.284
R2018 VGND.n1049 VGND.t2276 241.284
R2019 VGND.n2905 VGND.t2254 241.284
R2020 VGND.n2910 VGND.t2480 241.284
R2021 VGND.n928 VGND.t2466 241.284
R2022 VGND.t1401 VGND.t1436 222.15
R2023 VGND.t757 VGND.t1251 222.15
R2024 VGND.t782 VGND.t2068 222.15
R2025 VGND.t2673 VGND.t589 222.15
R2026 VGND.t2567 VGND.t800 222.15
R2027 VGND.t1187 VGND.t535 222.15
R2028 VGND.t2565 VGND.t1939 222.15
R2029 VGND.t659 VGND.t1551 222.15
R2030 VGND.t1434 VGND.t1634 222.15
R2031 VGND.t238 VGND.t1771 222.15
R2032 VGND.t1411 VGND.t2495 222.15
R2033 VGND.t1120 VGND.t1090 222.15
R2034 VGND.t2575 VGND.t1935 222.15
R2035 VGND.t2562 VGND.t542 222.15
R2036 VGND.t1432 VGND.t1662 222.15
R2037 VGND.t645 VGND.t15 222.15
R2038 VGND.t1953 VGND.t1430 222.15
R2039 VGND.t387 VGND.t448 222.15
R2040 VGND.t1413 VGND.t2277 222.15
R2041 VGND.t1134 VGND.t159 222.15
R2042 VGND.t1691 VGND.t2563 222.15
R2043 VGND.t712 VGND.t2535 222.15
R2044 VGND.t1438 VGND.t2481 222.15
R2045 VGND.t860 VGND.t1346 222.15
R2046 VGND.t2269 VGND.t2573 222.15
R2047 VGND.t1995 VGND.t2560 222.15
R2048 VGND.t54 VGND.t2571 222.15
R2049 VGND.t1376 VGND.t13 222.15
R2050 VGND.t2569 VGND.t1917 222.15
R2051 VGND.t663 VGND.t286 222.15
R2052 VGND.t1865 VGND.t1428 222.15
R2053 VGND.t2114 VGND.t354 222.15
R2054 VGND.t1301 VGND.t700 222.15
R2055 VGND.t78 VGND.t829 222.15
R2056 VGND.t2241 VGND.t1112 222.15
R2057 VGND.t1611 VGND.t932 222.15
R2058 VGND.t1734 VGND.t472 222.15
R2059 VGND.t602 VGND.t450 222.15
R2060 VGND.t1385 VGND.t470 222.15
R2061 VGND.t1542 VGND.t1845 222.15
R2062 VGND.t2070 VGND.t698 222.15
R2063 VGND.t1821 VGND.t1133 222.15
R2064 VGND.t2461 VGND.t1195 222.15
R2065 VGND.t431 VGND.t843 222.15
R2066 VGND.t1381 VGND.t1193 222.15
R2067 VGND.t573 VGND.t2493 222.15
R2068 VGND.t1636 VGND.t1118 222.15
R2069 VGND.t679 VGND.t1371 222.15
R2070 VGND.t2497 VGND.t1116 222.15
R2071 VGND.t220 VGND.t358 222.15
R2072 VGND.t1937 VGND.t1197 222.15
R2073 VGND.t438 VGND.t689 222.15
R2074 VGND.t1971 VGND.t704 222.15
R2075 VGND.t1322 VGND.t232 222.15
R2076 VGND.t2038 VGND.t702 222.15
R2077 VGND.t189 VGND.t897 222.15
R2078 VGND.t2024 VGND.t1191 222.15
R2079 VGND.t917 VGND.t1836 222.15
R2080 VGND.t1695 VGND.t1189 222.15
R2081 VGND.t223 VGND.t1806 222.15
R2082 VGND.t1867 VGND.t474 222.15
R2083 VGND.t2429 VGND.t75 222.15
R2084 VGND.t2271 VGND.t1114 222.15
R2085 VGND.t2186 VGND.t28 222.15
R2086 VGND.t1787 VGND.t2491 222.15
R2087 VGND.t2233 VGND.t1159 222.15
R2088 VGND.t2016 VGND.t1522 222.15
R2089 VGND.t595 VGND.t2561 222.15
R2090 VGND.t1795 VGND.t1687 222.15
R2091 VGND.t687 VGND.t525 222.15
R2092 VGND.t1925 VGND.t1793 222.15
R2093 VGND.t1557 VGND.t251 222.15
R2094 VGND.t1785 VGND.t2261 222.15
R2095 VGND.t2098 VGND.t1313 222.15
R2096 VGND.t494 VGND.t1327 222.15
R2097 VGND.t1092 VGND.t1484 222.15
R2098 VGND.t1325 VGND.t1913 222.15
R2099 VGND.t882 VGND.t548 222.15
R2100 VGND.t1857 VGND.t1528 222.15
R2101 VGND.t21 VGND.t2100 222.15
R2102 VGND.t1526 VGND.t1285 222.15
R2103 VGND.t908 VGND.t596 222.15
R2104 VGND.t2056 VGND.t1329 222.15
R2105 VGND.t1211 VGND.t1357 222.15
R2106 VGND.t1791 VGND.t1714 222.15
R2107 VGND.t151 VGND.t714 222.15
R2108 VGND.t1279 VGND.t1789 222.15
R2109 VGND.t1225 VGND.t204 222.15
R2110 VGND.t1323 VGND.t804 222.15
R2111 VGND.t1576 VGND.t83 222.15
R2112 VGND.t1799 VGND.t2467 222.15
R2113 VGND.t1121 VGND.t1356 222.15
R2114 VGND.t1797 VGND.t1644 222.15
R2115 VGND.t276 VGND.t292 222.15
R2116 VGND.t1618 VGND.t1524 222.15
R2117 VGND.t2135 VGND.t1987 222.15
R2118 VGND.t2046 VGND.t1271 222.15
R2119 VGND.t576 VGND.t264 222.15
R2120 VGND.t2089 VGND.t1654 222.15
R2121 VGND.t728 VGND.t846 222.15
R2122 VGND.t1965 VGND.t1102 222.15
R2123 VGND.t580 VGND.t718 222.15
R2124 VGND.t1277 VGND.t1873 222.15
R2125 VGND.t1578 VGND.t3 222.15
R2126 VGND.t2018 VGND.t482 222.15
R2127 VGND.t1303 VGND.t660 222.15
R2128 VGND.t2085 VGND.t2255 222.15
R2129 VGND.t883 VGND.t326 222.15
R2130 VGND.t1859 VGND.t2083 222.15
R2131 VGND.t1673 VGND.t928 222.15
R2132 VGND.t480 VGND.t2263 222.15
R2133 VGND.t1341 VGND.t586 222.15
R2134 VGND.t496 VGND.t478 222.15
R2135 VGND.t850 VGND.t2101 222.15
R2136 VGND.t2087 VGND.t1915 222.15
R2137 VGND.t445 VGND.t461 222.15
R2138 VGND.t1879 VGND.t1275 222.15
R2139 VGND.t1808 VGND.t242 222.15
R2140 VGND.t1273 VGND.t488 222.15
R2141 VGND.t1818 VGND.t1239 222.15
R2142 VGND.t1907 VGND.t1108 222.15
R2143 VGND.t1988 VGND.t166 222.15
R2144 VGND.t1718 VGND.t1106 222.15
R2145 VGND.t2557 VGND.t909 222.15
R2146 VGND.t1104 VGND.t1620 222.15
R2147 VGND.t1145 VGND.t175 222.15
R2148 VGND.t2052 VGND.t476 222.15
R2149 VGND.t2638 VGND.t256 222.15
R2150 VGND.t2527 VGND.t2455 222.15
R2151 VGND.t2533 VGND.t1153 222.15
R2152 VGND.t768 VGND.t1628 222.15
R2153 VGND.t235 VGND.t1605 222.15
R2154 VGND.t2507 VGND.t1801 222.15
R2155 VGND.t555 VGND.t447 222.15
R2156 VGND.t1409 VGND.t2281 222.15
R2157 VGND.t772 VGND.t1238 222.15
R2158 VGND.t1656 VGND.t2525 222.15
R2159 VGND.t259 VGND.t1849 222.15
R2160 VGND.t764 VGND.t2487 222.15
R2161 VGND.t907 VGND.t1086 222.15
R2162 VGND.t2265 VGND.t762 222.15
R2163 VGND.t567 VGND.t1188 222.15
R2164 VGND.t2523 VGND.t2020 222.15
R2165 VGND.t1581 VGND.t673 222.15
R2166 VGND.t1675 VGND.t2521 222.15
R2167 VGND.t214 VGND.t1577 222.15
R2168 VGND.t766 VGND.t1861 222.15
R2169 VGND.t2531 VGND.t2541 222.15
R2170 VGND.t52 VGND.t1407 222.15
R2171 VGND.t1320 VGND.t231 222.15
R2172 VGND.t1405 VGND.t2247 222.15
R2173 VGND.t716 VGND.t2426 222.15
R2174 VGND.t1855 VGND.t760 222.15
R2175 VGND.t911 VGND.t771 222.15
R2176 VGND.t758 VGND.t1881 222.15
R2177 VGND.t725 VGND.t361 222.15
R2178 VGND.t1803 VGND.t2054 222.15
R2179 VGND.t1549 VGND.t515 222.15
R2180 VGND.t1911 VGND.t2519 222.15
R2181 VGND.t2158 VGND.t2097 222.15
R2182 VGND.t1783 VGND.t1391 222.15
R2183 VGND.t2391 VGND.t756 222.15
R2184 VGND.t1773 VGND.t2060 222.15
R2185 VGND.t1805 VGND.t588 222.15
R2186 VGND.t790 VGND.t876 222.15
R2187 VGND.t524 VGND.t779 222.15
R2188 VGND.t1929 VGND.t874 222.15
R2189 VGND.t1550 VGND.t94 222.15
R2190 VGND.t1624 VGND.t1781 222.15
R2191 VGND.t1770 VGND.t452 222.15
R2192 VGND.t2030 VGND.t1231 222.15
R2193 VGND.t302 VGND.t770 222.15
R2194 VGND.t2012 VGND.t1229 222.15
R2195 VGND.t541 VGND.t2082 222.15
R2196 VGND.t1650 VGND.t1779 222.15
R2197 VGND.t14 VGND.t280 222.15
R2198 VGND.t2475 VGND.t1777 222.15
R2199 VGND.t386 VGND.t1185 222.15
R2200 VGND.t72 VGND.t1233 222.15
R2201 VGND.t158 VGND.t656 222.15
R2202 VGND.t1679 VGND.t872 222.15
R2203 VGND.t711 VGND.t2091 222.15
R2204 VGND.t2469 VGND.t870 222.15
R2205 VGND.t1345 VGND.t1141 222.15
R2206 VGND.t68 VGND.t1227 222.15
R2207 VGND.t1994 VGND.t2099 222.15
R2208 VGND.t504 VGND.t880 222.15
R2209 VGND.t1375 VGND.t356 222.15
R2210 VGND.t878 VGND.t1905 222.15
R2211 VGND.t1531 VGND.t285 222.15
R2212 VGND.t1897 VGND.t1775 222.15
R2213 VGND.t2112 VGND.t230 222.15
R2214 VGND.t1493 VGND.t1291 222.15
R2215 VGND.t1264 VGND.t1164 222.15
R2216 VGND.t2553 VGND.t1923 222.15
R2217 VGND.t1456 VGND.t1831 222.15
R2218 VGND.t377 VGND.t1722 222.15
R2219 VGND.t206 VGND.t552 222.15
R2220 VGND.t1499 VGND.t1660 222.15
R2221 VGND.t275 VGND.t1558 222.15
R2222 VGND.t1491 VGND.t2062 222.15
R2223 VGND.t139 VGND.t1314 222.15
R2224 VGND.t2549 VGND.t1945 222.15
R2225 VGND.t2416 VGND.t1093 222.15
R2226 VGND.t2547 VGND.t1652 222.15
R2227 VGND.t92 VGND.t549 222.15
R2228 VGND.t1489 VGND.t1626 222.15
R2229 VGND.t1461 VGND.t315 222.15
R2230 VGND.t1487 VGND.t2036 222.15
R2231 VGND.t221 VGND.t597 222.15
R2232 VGND.t2551 VGND.t2014 222.15
R2233 VGND.t2417 VGND.t1212 222.15
R2234 VGND.t1497 VGND.t1959 222.15
R2235 VGND.t446 VGND.t1266 222.15
R2236 VGND.t1495 VGND.t2026 222.15
R2237 VGND.t1249 VGND.t1226 222.15
R2238 VGND.t2010 VGND.t2545 222.15
R2239 VGND.t2681 VGND.t1270 222.15
R2240 VGND.t1681 VGND.t381 222.15
R2241 VGND.t451 VGND.t1250 222.15
R2242 VGND.t379 VGND.t1899 222.15
R2243 VGND.t938 VGND.t293 222.15
R2244 VGND.t70 VGND.t1485 222.15
R2245 VGND.t2138 VGND.t1186 222.15
R2246 VGND.t2473 VGND.t652 222.15
R2247 VGND.t577 VGND.t560 222.15
R2248 VGND.t1903 VGND.t2004 222.15
R2249 VGND.t1088 VGND.t847 222.15
R2250 VGND.t893 VGND.t1677 222.15
R2251 VGND.t1503 VGND.t583 222.15
R2252 VGND.t891 VGND.t1909 222.15
R2253 VGND.t905 VGND.t4 222.15
R2254 VGND.t60 VGND.t650 222.15
R2255 VGND.t1304 VGND.t562 222.15
R2256 VGND.t1100 VGND.t484 222.15
R2257 VGND.t1373 VGND.t327 222.15
R2258 VGND.t1728 VGND.t1098 222.15
R2259 VGND.t1674 VGND.t252 222.15
R2260 VGND.t648 VGND.t1891 222.15
R2261 VGND.t717 VGND.t587 222.15
R2262 VGND.t1640 VGND.t776 222.15
R2263 VGND.t851 VGND.t929 222.15
R2264 VGND.t1901 VGND.t798 222.15
R2265 VGND.t1851 VGND.t153 222.15
R2266 VGND.t1397 VGND.t889 222.15
R2267 VGND.t1809 VGND.t647 222.15
R2268 VGND.t654 VGND.t1630 222.15
R2269 VGND.t1339 VGND.t1240 222.15
R2270 VGND.t792 VGND.t1096 222.15
R2271 VGND.t1989 VGND.t225 222.15
R2272 VGND.t1094 VGND.t2459 222.15
R2273 VGND.t239 VGND.t2558 222.15
R2274 VGND.t895 VGND.t1967 222.15
R2275 VGND.t91 VGND.t176 222.15
R2276 VGND.t2509 VGND.t774 222.15
R2277 VGND.t2640 VGND.t1343 222.15
R2278 VGND.t311 VGND.t2028 222.15
R2279 VGND.t609 VGND.t834 222.15
R2280 VGND.t2401 VGND.t1646 222.15
R2281 VGND.t726 VGND.t845 222.15
R2282 VGND.t1957 VGND.t899 222.15
R2283 VGND.t582 VGND.t1819 222.15
R2284 VGND.t1335 VGND.t1853 222.15
R2285 VGND.t1592 VGND.t1445 222.15
R2286 VGND.t309 VGND.t2006 222.15
R2287 VGND.t2001 VGND.t1752 222.15
R2288 VGND.t2397 VGND.t2243 222.15
R2289 VGND.t706 VGND.t324 222.15
R2290 VGND.t2395 VGND.t1893 222.15
R2291 VGND.t773 VGND.t1672 222.15
R2292 VGND.t307 VGND.t62 222.15
R2293 VGND.t234 VGND.t585 222.15
R2294 VGND.t305 VGND.t486 222.15
R2295 VGND.t828 VGND.t849 222.15
R2296 VGND.t2399 VGND.t1732 222.15
R2297 VGND.t205 VGND.t460 222.15
R2298 VGND.t1333 VGND.t1295 222.15
R2299 VGND.t646 VGND.t1807 222.15
R2300 VGND.t1331 VGND.t2066 222.15
R2301 VGND.t1416 VGND.t1575 222.15
R2302 VGND.t1724 VGND.t2393 222.15
R2303 VGND.t1263 VGND.t181 222.15
R2304 VGND.t1399 VGND.t903 222.15
R2305 VGND.t2556 VGND.t1132 222.15
R2306 VGND.t901 VGND.t2511 222.15
R2307 VGND.t2418 VGND.t173 222.15
R2308 VGND.t794 VGND.t2529 222.15
R2309 VGND.t2631 VGND.t1580 222.15
R2310 VGND.t1768 VGND.t1943 222.15
R2311 VGND.t2081 VGND.t1152 222.15
R2312 VGND.t1758 VGND.t1622 222.15
R2313 VGND.t715 VGND.t1705 222.15
R2314 VGND.t1712 VGND.t2505 222.15
R2315 VGND.t826 VGND.t152 222.15
R2316 VGND.t1710 VGND.t2259 222.15
R2317 VGND.t931 VGND.t1237 222.15
R2318 VGND.t1766 VGND.t1648 222.15
R2319 VGND.t84 VGND.t258 222.15
R2320 VGND.t1754 VGND.t2471 222.15
R2321 VGND.t1594 VGND.t1085 222.15
R2322 VGND.t126 VGND.t64 222.15
R2323 VGND.t781 VGND.t566 222.15
R2324 VGND.t1764 VGND.t2008 222.15
R2325 VGND.t119 VGND.t672 222.15
R2326 VGND.t1762 VGND.t2245 222.15
R2327 VGND.t888 VGND.t729 222.15
R2328 VGND.t1756 VGND.t1895 222.15
R2329 VGND.t2536 VGND.t1215 222.15
R2330 VGND.t1708 VGND.t502 222.15
R2331 VGND.t825 VGND.t1319 222.15
R2332 VGND.t1706 VGND.t2237 222.15
R2333 VGND.t1421 VGND.t2423 222.15
R2334 VGND.t1889 VGND.t124 222.15
R2335 VGND.t2686 VGND.t1269 222.15
R2336 VGND.t1297 VGND.t122 222.15
R2337 VGND.t464 VGND.t253 222.15
R2338 VGND.t120 VGND.t796 222.15
R2339 VGND.t1548 VGND.t514 222.15
R2340 VGND.t1726 VGND.t1760 222.15
R2341 VGND.t2153 VGND.t213 222.15
R2342 VGND.t1299 VGND.t813 222.15
R2343 VGND.t1151 VGND.t182 222.15
R2344 VGND.t2235 VGND.t399 222.15
R2345 VGND.t370 VGND.t2403 222.15
R2346 VGND.t1730 VGND.t821 222.15
R2347 VGND.t113 VGND.t212 222.15
R2348 VGND.t819 VGND.t1383 222.15
R2349 VGND.t85 VGND.t785 222.15
R2350 VGND.t811 VGND.t2064 222.15
R2351 VGND.t118 VGND.t1702 222.15
R2352 VGND.t395 VGND.t2457 222.15
R2353 VGND.t1144 VGND.t735 222.15
R2354 VGND.t393 VGND.t1658 222.15
R2355 VGND.t1452 VGND.t1666 222.15
R2356 VGND.t405 VGND.t1632 222.15
R2357 VGND.t1595 VGND.t330 222.15
R2358 VGND.t403 VGND.t2048 222.15
R2359 VGND.t1501 VGND.t1838 222.15
R2360 VGND.t397 VGND.t1931 222.15
R2361 VGND.t1142 VGND.t458 222.15
R2362 VGND.t817 VGND.t1969 222.15
R2363 VGND.t241 VGND.t1749 222.15
R2364 VGND.t2032 VGND.t815 222.15
R2365 VGND.t1617 VGND.t661 222.15
R2366 VGND.t2022 VGND.t391 222.15
R2367 VGND.t1257 VGND.t2102 222.15
R2368 VGND.t1689 VGND.t389 222.15
R2369 VGND.t34 VGND.t561 222.15
R2370 VGND.t1863 VGND.t823 222.15
R2371 VGND.t168 VGND.t2559 222.15
R2372 VGND.t2267 VGND.t401 222.15
R2373 VGND.t2590 VGND.t86 222.15
R2374 VGND.t423 VGND.t1941 222.15
R2375 VGND.t898 VGND.t1158 222.15
R2376 VGND.t2412 VGND.t2515 222.15
R2377 VGND.t1342 VGND.t590 222.15
R2378 VGND.t1568 VGND.t2501 222.15
R2379 VGND.t1455 VGND.t526 222.15
R2380 VGND.t66 VGND.t429 222.15
R2381 VGND.t1556 VGND.t1372 222.15
R2382 VGND.t421 VGND.t1642 222.15
R2383 VGND.t1502 VGND.t1772 222.15
R2384 VGND.t1875 VGND.t2408 222.15
R2385 VGND.t1091 VGND.t1265 222.15
R2386 VGND.t2406 VGND.t58 222.15
R2387 VGND.t140 VGND.t543 222.15
R2388 VGND.t2002 VGND.t419 222.15
R2389 VGND.t16 VGND.t1532 222.15
R2390 VGND.t417 VGND.t2239 222.15
R2391 VGND.t1420 VGND.t1583 222.15
R2392 VGND.t2410 VGND.t1887 222.15
R2393 VGND.t469 VGND.t1210 222.15
R2394 VGND.t498 VGND.t427 222.15
R2395 VGND.t713 VGND.t1344 222.15
R2396 VGND.t1927 VGND.t425 222.15
R2397 VGND.t1224 VGND.t927 222.15
R2398 VGND.t2404 VGND.t1885 222.15
R2399 VGND.t128 VGND.t1996 222.15
R2400 VGND.t1572 VGND.t1287 222.15
R2401 VGND.t279 VGND.t1355 222.15
R2402 VGND.t1570 VGND.t788 222.15
R2403 VGND.t1979 VGND.t291 222.15
R2404 VGND.t1720 VGND.t2414 222.15
R2405 VGND.t2132 VGND.t2392 222.15
R2406 VGND.t2517 VGND.t2449 222.15
R2407 VGND.t1150 VGND.t30 222.15
R2408 VGND.t742 VGND.t1389 222.15
R2409 VGND.t608 VGND.t369 222.15
R2410 VGND.t1664 VGND.t612 222.15
R2411 VGND.t116 VGND.t2092 222.15
R2412 VGND.t610 VGND.t1955 222.15
R2413 VGND.t2674 VGND.t784 222.15
R2414 VGND.t1947 VGND.t750 222.15
R2415 VGND.t1701 VGND.t1415 222.15
R2416 VGND.t738 VGND.t1693 222.15
R2417 VGND.t76 VGND.t734 222.15
R2418 VGND.t2485 VGND.t620 222.15
R2419 VGND.t138 VGND.t1814 222.15
R2420 VGND.t748 VGND.t2040 222.15
R2421 VGND.t2537 VGND.t644 222.15
R2422 VGND.t56 VGND.t746 222.15
R2423 VGND.t1837 VGND.t147 222.15
R2424 VGND.t740 VGND.t2257 222.15
R2425 VGND.t536 VGND.t455 222.15
R2426 VGND.t1869 VGND.t2453 222.15
R2427 VGND.t1748 VGND.t778 222.15
R2428 VGND.t506 VGND.t2451 222.15
R2429 VGND.t1614 VGND.t887 222.15
R2430 VGND.t2249 VGND.t618 222.15
R2431 VGND.t1256 VGND.t449 222.15
R2432 VGND.t1921 VGND.t616 222.15
R2433 VGND.t31 VGND.t355 222.15
R2434 VGND.t614 VGND.t1281 222.15
R2435 VGND.t1829 VGND.t167 222.15
R2436 VGND.t490 VGND.t744 222.15
R2437 VGND.t2587 VGND.t150 222.15
R2438 VGND.t197 VGND.t802 222.15
R2439 VGND.t925 VGND.t77 222.15
R2440 VGND.t1289 VGND.t2445 222.15
R2441 VGND.t1610 VGND.t1418 222.15
R2442 VGND.t682 VGND.t1638 222.15
R2443 VGND.t559 VGND.t810 222.15
R2444 VGND.t48 VGND.t2499 222.15
R2445 VGND.t827 VGND.t1541 222.15
R2446 VGND.t195 VGND.t1393 222.15
R2447 VGND.t2534 VGND.t1820 222.15
R2448 VGND.t2441 VGND.t1973 222.15
R2449 VGND.t2532 VGND.t1087 222.15
R2450 VGND.t2439 VGND.t2042 222.15
R2451 VGND.t1419 VGND.t572 222.15
R2452 VGND.t193 VGND.t1949 222.15
R2453 VGND.t117 VGND.t678 222.15
R2454 VGND.t191 VGND.t1697 222.15
R2455 VGND.t1337 VGND.t219 222.15
R2456 VGND.t2489 VGND.t2443 222.15
R2457 VGND.t2542 VGND.t203 222.15
R2458 VGND.t2273 VGND.t201 222.15
R2459 VGND.t1321 VGND.t1080 222.15
R2460 VGND.t199 VGND.t1685 222.15
R2461 VGND.t1830 VGND.t2427 222.15
R2462 VGND.t2437 VGND.t2477 222.15
R2463 VGND.t681 VGND.t916 222.15
R2464 VGND.t1871 VGND.t2435 222.15
R2465 VGND.t362 VGND.t926 222.15
R2466 VGND.t492 VGND.t684 222.15
R2467 VGND.t2428 VGND.t388 222.15
R2468 VGND.t2251 VGND.t2447 222.15
R2469 VGND.t2173 VGND.t1579 222.15
R2470 VGND.t862 VGND.t1736 222.15
R2471 VGND.t841 VGND.t835 222.15
R2472 VGND.t273 VGND.t500 222.15
R2473 VGND.t468 VGND.t844 222.15
R2474 VGND.t1422 VGND.t2072 222.15
R2475 VGND.t74 VGND.t581 222.15
R2476 VGND.t2463 VGND.t868 222.15
R2477 VGND.t1444 VGND.t842 222.15
R2478 VGND.t1293 VGND.t856 222.15
R2479 VGND.t1753 VGND.t1844 222.15
R2480 VGND.t2513 VGND.t269 222.15
R2481 VGND.t325 VGND.t236 222.15
R2482 VGND.t1951 VGND.t267 222.15
R2483 VGND.t1671 VGND.t1374 222.15
R2484 VGND.t1395 VGND.t854 222.15
R2485 VGND.t584 VGND.t780 222.15
R2486 VGND.t1975 VGND.t852 222.15
R2487 VGND.t848 VGND.t861 222.15
R2488 VGND.t271 VGND.t2044 222.15
R2489 VGND.t886 VGND.t459 222.15
R2490 VGND.t866 VGND.t1933 222.15
R2491 VGND.t688 VGND.t657 222.15
R2492 VGND.t864 VGND.t1963 222.15
R2493 VGND.t1588 VGND.t1574 222.15
R2494 VGND.t265 VGND.t2034 222.15
R2495 VGND.t697 VGND.t1262 222.15
R2496 VGND.t2275 VGND.t1426 222.15
R2497 VGND.t2555 VGND.t1143 222.15
R2498 VGND.t1424 VGND.t2253 222.15
R2499 VGND.t1089 VGND.t174 222.15
R2500 VGND.t2479 VGND.t723 222.15
R2501 VGND.t2630 VGND.t278 222.15
R2502 VGND.t2279 VGND.t2669 222.15
R2503 VGND.t624 VGND.t558 222.15
R2504 VGND.t2588 VGND.t1961 222.15
R2505 VGND.t930 VGND.t1986 222.15
R2506 VGND.t2163 VGND.t2483 222.15
R2507 VGND.t1199 VGND.t112 222.15
R2508 VGND.t2141 VGND.t1883 222.15
R2509 VGND.t385 VGND.t1545 222.15
R2510 VGND.t2658 VGND.t1683 222.15
R2511 VGND.t1593 VGND.t1828 222.15
R2512 VGND.t2223 VGND.t1919 222.15
R2513 VGND.t359 VGND.t696 222.15
R2514 VGND.t2212 VGND.t1877 222.15
R2515 VGND.t228 VGND.t133 222.15
R2516 VGND.t2654 VGND.t50 222.15
R2517 VGND.t149 VGND.t341 222.15
R2518 VGND.t2636 VGND.t2058 222.15
R2519 VGND.t910 VGND.t670 222.15
R2520 VGND.t2225 VGND.t1716 222.15
R2521 VGND.t2234 VGND.t439 222.15
R2522 VGND.t1511 VGND.t1283 222.15
R2523 VGND.t2538 VGND.t1130 222.15
R2524 VGND.t2133 VGND.t2050 222.15
R2525 VGND.t233 VGND.t190 222.15
R2526 VGND.t2207 VGND.t1403 222.15
R2527 VGND.t658 VGND.t924 222.15
R2528 VGND.t2194 VGND.t1387 222.15
R2529 VGND.t90 VGND.t224 222.15
R2530 VGND.t2169 VGND.t2503 222.15
R2531 VGND.t222 VGND.t2432 222.15
R2532 VGND.t2465 VGND.t2615 222.15
R2533 VGND.t2198 VGND.t444 222.15
R2534 VGND.n2346 VGND.n3 218.73
R2535 VGND.n489 VGND.n487 214.365
R2536 VGND.n489 VGND.n488 214.365
R2537 VGND.n479 VGND.n477 214.365
R2538 VGND.n479 VGND.n478 214.365
R2539 VGND.n497 VGND.n495 214.365
R2540 VGND.n497 VGND.n496 214.365
R2541 VGND.n2270 VGND.n2268 214.365
R2542 VGND.n2270 VGND.n2269 214.365
R2543 VGND.n2260 VGND.n2258 214.365
R2544 VGND.n2260 VGND.n2259 214.365
R2545 VGND.n2278 VGND.n2276 214.365
R2546 VGND.n2278 VGND.n2277 214.365
R2547 VGND.n525 VGND.n523 214.365
R2548 VGND.n525 VGND.n524 214.365
R2549 VGND.n515 VGND.n513 214.365
R2550 VGND.n515 VGND.n514 214.365
R2551 VGND.n533 VGND.n531 214.365
R2552 VGND.n533 VGND.n532 214.365
R2553 VGND.n2191 VGND.n2190 214.365
R2554 VGND.n1140 VGND.n1139 213.613
R2555 VGND.n1142 VGND.n1141 213.613
R2556 VGND.n1112 VGND.n1110 213.613
R2557 VGND.n1112 VGND.n1111 213.613
R2558 VGND.n1115 VGND.n1113 213.613
R2559 VGND.n1115 VGND.n1114 213.613
R2560 VGND.n2236 VGND.n2229 213.613
R2561 VGND.n2236 VGND.n2230 213.613
R2562 VGND.n2234 VGND.n2231 213.613
R2563 VGND.n2234 VGND.n2233 213.613
R2564 VGND.n1374 VGND.n1367 213.613
R2565 VGND.n1374 VGND.n1368 213.613
R2566 VGND.n1372 VGND.n1369 213.613
R2567 VGND.n1372 VGND.n1371 213.613
R2568 VGND.n1154 VGND.t1165 211.359
R2569 VGND.n179 VGND.n175 207.965
R2570 VGND.n179 VGND.n176 207.965
R2571 VGND.n173 VGND.n171 207.965
R2572 VGND.n173 VGND.n172 207.965
R2573 VGND.n186 VGND.n169 207.965
R2574 VGND.n186 VGND.n170 207.965
R2575 VGND.n98 VGND.n97 207.965
R2576 VGND.n110 VGND.n95 207.965
R2577 VGND.n102 VGND.n100 207.965
R2578 VGND.n80 VGND.n76 207.965
R2579 VGND.n80 VGND.n77 207.965
R2580 VGND.n74 VGND.n72 207.965
R2581 VGND.n74 VGND.n73 207.965
R2582 VGND.n87 VGND.n70 207.965
R2583 VGND.n87 VGND.n71 207.965
R2584 VGND.n148 VGND.n144 207.965
R2585 VGND.n148 VGND.n145 207.965
R2586 VGND.n142 VGND.n140 207.965
R2587 VGND.n142 VGND.n141 207.965
R2588 VGND.n155 VGND.n138 207.965
R2589 VGND.n155 VGND.n139 207.965
R2590 VGND.n2188 VGND.n2187 207.965
R2591 VGND.n2205 VGND.n2185 207.965
R2592 VGND.n2981 VGND.n2979 207.213
R2593 VGND.n2981 VGND.n2980 207.213
R2594 VGND.n2985 VGND.n2976 207.213
R2595 VGND.n2985 VGND.n2977 207.213
R2596 VGND.n18 VGND.n16 207.213
R2597 VGND.n18 VGND.n17 207.213
R2598 VGND.n22 VGND.n14 207.213
R2599 VGND.n22 VGND.n15 207.213
R2600 VGND.n2951 VGND.n2950 207.213
R2601 VGND.n2955 VGND.n2949 207.213
R2602 VGND.n44 VGND.n42 207.213
R2603 VGND.n44 VGND.n43 207.213
R2604 VGND.n48 VGND.n40 207.213
R2605 VGND.n48 VGND.n41 207.213
R2606 VGND.n109 VGND.n96 207.213
R2607 VGND.n2204 VGND.n2186 207.213
R2608 VGND.t997 VGND.t2613 203.242
R2609 VGND.t2190 VGND.t946 203.242
R2610 VGND.t952 VGND.t2128 203.242
R2611 VGND.t2104 VGND.t970 203.242
R2612 VGND.t1045 VGND.t2188 203.242
R2613 VGND.t2176 VGND.t1051 203.242
R2614 VGND.t973 VGND.t2154 203.242
R2615 VGND.t2601 VGND.t1015 203.242
R2616 VGND.t1024 VGND.t2581 203.242
R2617 VGND.t2149 VGND.t1063 203.242
R2618 VGND.t979 VGND.t2656 203.242
R2619 VGND.t2645 VGND.t1027 203.242
R2620 VGND.t1066 VGND.t2210 203.242
R2621 VGND.t2139 VGND.t1075 203.242
R2622 VGND.t991 VGND.t2634 203.242
R2623 VGND.t2221 VGND.t1033 203.242
R2624 VGND VGND.n332 194.419
R2625 VGND VGND.n356 194.419
R2626 VGND VGND.n363 194.419
R2627 VGND VGND.n366 194.419
R2628 VGND VGND.n374 194.419
R2629 VGND VGND.n377 194.419
R2630 VGND VGND.n385 194.419
R2631 VGND VGND.n324 194.419
R2632 VGND VGND.n313 194.419
R2633 VGND VGND.n308 194.419
R2634 VGND VGND.n310 194.419
R2635 VGND VGND.n2729 194.419
R2636 VGND VGND.n292 194.419
R2637 VGND VGND.n295 194.419
R2638 VGND VGND.n202 194.419
R2639 VGND.n887 VGND.n886 194.391
R2640 VGND.n1332 VGND.n889 194.391
R2641 VGND.n895 VGND.n893 194.391
R2642 VGND.n931 VGND.n930 194.391
R2643 VGND.n936 VGND.n935 194.391
R2644 VGND.n941 VGND.n940 194.391
R2645 VGND.n946 VGND.n945 194.391
R2646 VGND.n951 VGND.n950 194.391
R2647 VGND.n956 VGND.n955 194.391
R2648 VGND.n961 VGND.n960 194.391
R2649 VGND.n966 VGND.n965 194.391
R2650 VGND.n971 VGND.n970 194.391
R2651 VGND.n976 VGND.n975 194.391
R2652 VGND.n981 VGND.n980 194.391
R2653 VGND.n986 VGND.n985 194.391
R2654 VGND.n1281 VGND.n996 194.391
R2655 VGND.n1274 VGND.n1273 194.391
R2656 VGND.n1231 VGND.n1230 194.391
R2657 VGND.n1236 VGND.n1229 194.391
R2658 VGND.n1227 VGND.n1226 194.391
R2659 VGND.n1243 VGND.n1224 194.391
R2660 VGND.n1222 VGND.n1221 194.391
R2661 VGND.n1217 VGND.n1216 194.391
R2662 VGND.n1211 VGND.n1002 194.391
R2663 VGND.n1204 VGND.n1203 194.391
R2664 VGND.n1008 VGND.n1007 194.391
R2665 VGND.n1185 VGND.n1184 194.391
R2666 VGND.n1179 VGND.n1010 194.391
R2667 VGND.n1172 VGND.n1171 194.391
R2668 VGND.n1169 VGND.n1012 194.391
R2669 VGND.n330 VGND.n329 194.391
R2670 VGND.n396 VGND.n395 194.391
R2671 VGND.n2638 VGND.n2637 194.391
R2672 VGND.n2643 VGND.n2642 194.391
R2673 VGND.n2648 VGND.n2647 194.391
R2674 VGND.n2653 VGND.n2652 194.391
R2675 VGND.n2658 VGND.n2657 194.391
R2676 VGND.n2663 VGND.n2662 194.391
R2677 VGND.n2668 VGND.n2667 194.391
R2678 VGND.n393 VGND.n392 194.391
R2679 VGND.n2714 VGND.n2713 194.391
R2680 VGND.n319 VGND.n318 194.391
R2681 VGND.n2747 VGND.n2746 194.391
R2682 VGND.n303 VGND.n302 194.391
R2683 VGND.n2752 VGND.n2751 194.391
R2684 VGND.n2787 VGND.n2786 194.391
R2685 VGND.n286 VGND.n285 194.391
R2686 VGND.n400 VGND.n399 194.391
R2687 VGND.n2342 VGND.n2341 194.391
R2688 VGND.n2337 VGND.n2336 194.391
R2689 VGND.n2332 VGND.n2331 194.391
R2690 VGND.n2327 VGND.n2326 194.391
R2691 VGND.n2322 VGND.n2321 194.391
R2692 VGND.n2317 VGND.n2316 194.391
R2693 VGND.n2312 VGND.n2311 194.391
R2694 VGND.n2307 VGND.n2306 194.391
R2695 VGND.n2302 VGND.n2301 194.391
R2696 VGND.n2297 VGND.n2296 194.391
R2697 VGND.n2292 VGND.n2291 194.391
R2698 VGND.n2287 VGND.n2286 194.391
R2699 VGND.n414 VGND.n413 194.391
R2700 VGND.n2540 VGND.n2539 194.391
R2701 VGND.n2535 VGND.n416 194.391
R2702 VGND.n469 VGND.n468 194.391
R2703 VGND.n471 VGND.n470 194.391
R2704 VGND.n2376 VGND.n2375 194.391
R2705 VGND.n459 VGND.n458 194.391
R2706 VGND.n2402 VGND.n2401 194.391
R2707 VGND.n451 VGND.n450 194.391
R2708 VGND.n2428 VGND.n2427 194.391
R2709 VGND.n443 VGND.n442 194.391
R2710 VGND.n2454 VGND.n2453 194.391
R2711 VGND.n435 VGND.n434 194.391
R2712 VGND.n2480 VGND.n2479 194.391
R2713 VGND.n427 VGND.n426 194.391
R2714 VGND.n2511 VGND.n2510 194.391
R2715 VGND.n2516 VGND.n2515 194.391
R2716 VGND.n2521 VGND.n2520 194.391
R2717 VGND.n2528 VGND.n418 194.391
R2718 VGND.n466 VGND.n465 194.391
R2719 VGND.n2363 VGND.n2362 194.391
R2720 VGND.n463 VGND.n462 194.391
R2721 VGND.n2389 VGND.n2388 194.391
R2722 VGND.n455 VGND.n454 194.391
R2723 VGND.n2415 VGND.n2414 194.391
R2724 VGND.n447 VGND.n446 194.391
R2725 VGND.n2441 VGND.n2440 194.391
R2726 VGND.n439 VGND.n438 194.391
R2727 VGND.n2467 VGND.n2466 194.391
R2728 VGND.n431 VGND.n430 194.391
R2729 VGND.n2493 VGND.n2492 194.391
R2730 VGND.n423 VGND.n422 194.391
R2731 VGND.n2498 VGND.n2497 194.391
R2732 VGND.n2809 VGND.n2808 194.391
R2733 VGND.n2816 VGND.n276 194.391
R2734 VGND.n625 VGND.n624 194.391
R2735 VGND.n1910 VGND.n1909 194.391
R2736 VGND.n622 VGND.n621 194.391
R2737 VGND.n1921 VGND.n1920 194.391
R2738 VGND.n619 VGND.n618 194.391
R2739 VGND.n1932 VGND.n1931 194.391
R2740 VGND.n616 VGND.n615 194.391
R2741 VGND.n1943 VGND.n1942 194.391
R2742 VGND.n613 VGND.n612 194.391
R2743 VGND.n1954 VGND.n1953 194.391
R2744 VGND.n610 VGND.n609 194.391
R2745 VGND.n1965 VGND.n1964 194.391
R2746 VGND.n607 VGND.n606 194.391
R2747 VGND.n1976 VGND.n1975 194.391
R2748 VGND.n1981 VGND.n1980 194.391
R2749 VGND.n1988 VGND.n605 194.391
R2750 VGND.n590 VGND.n589 194.391
R2751 VGND.n596 VGND.n595 194.391
R2752 VGND.n593 VGND.n592 194.391
R2753 VGND.n2055 VGND.n2054 194.391
R2754 VGND.n2050 VGND.n2049 194.391
R2755 VGND.n2045 VGND.n2044 194.391
R2756 VGND.n2040 VGND.n2039 194.391
R2757 VGND.n2035 VGND.n2034 194.391
R2758 VGND.n2030 VGND.n2029 194.391
R2759 VGND.n2025 VGND.n2024 194.391
R2760 VGND.n2020 VGND.n2019 194.391
R2761 VGND.n2015 VGND.n2014 194.391
R2762 VGND.n2010 VGND.n2009 194.391
R2763 VGND.n2005 VGND.n2004 194.391
R2764 VGND.n2000 VGND.n600 194.391
R2765 VGND.n1995 VGND.n1993 194.391
R2766 VGND.n587 VGND.n586 194.391
R2767 VGND.n2069 VGND.n2068 194.391
R2768 VGND.n2074 VGND.n2073 194.391
R2769 VGND.n2079 VGND.n2078 194.391
R2770 VGND.n2084 VGND.n2083 194.391
R2771 VGND.n2089 VGND.n2088 194.391
R2772 VGND.n2094 VGND.n2093 194.391
R2773 VGND.n2099 VGND.n2098 194.391
R2774 VGND.n2104 VGND.n2103 194.391
R2775 VGND.n2109 VGND.n2108 194.391
R2776 VGND.n2114 VGND.n2113 194.391
R2777 VGND.n2119 VGND.n2118 194.391
R2778 VGND.n584 VGND.n583 194.391
R2779 VGND.n2124 VGND.n2123 194.391
R2780 VGND.n2834 VGND.n2833 194.391
R2781 VGND.n2841 VGND.n264 194.391
R2782 VGND.n547 VGND.n546 194.391
R2783 VGND.n2176 VGND.n549 194.391
R2784 VGND.n1757 VGND.n1755 194.391
R2785 VGND.n1761 VGND.n1760 194.391
R2786 VGND.n1752 VGND.n1751 194.391
R2787 VGND.n1772 VGND.n1771 194.391
R2788 VGND.n1749 VGND.n1748 194.391
R2789 VGND.n1783 VGND.n1782 194.391
R2790 VGND.n1746 VGND.n1745 194.391
R2791 VGND.n1794 VGND.n1793 194.391
R2792 VGND.n1743 VGND.n1742 194.391
R2793 VGND.n1805 VGND.n1804 194.391
R2794 VGND.n1740 VGND.n1739 194.391
R2795 VGND.n1816 VGND.n1815 194.391
R2796 VGND.n1821 VGND.n1820 194.391
R2797 VGND.n1828 VGND.n1738 194.391
R2798 VGND.n628 VGND.n627 194.391
R2799 VGND.n1678 VGND.n1677 194.391
R2800 VGND.n1675 VGND.n1674 194.391
R2801 VGND.n1689 VGND.n1688 194.391
R2802 VGND.n1694 VGND.n1693 194.391
R2803 VGND.n1699 VGND.n1698 194.391
R2804 VGND.n1704 VGND.n1703 194.391
R2805 VGND.n1709 VGND.n1708 194.391
R2806 VGND.n1714 VGND.n1713 194.391
R2807 VGND.n1719 VGND.n1718 194.391
R2808 VGND.n1724 VGND.n1723 194.391
R2809 VGND.n1729 VGND.n1728 194.391
R2810 VGND.n1672 VGND.n1671 194.391
R2811 VGND.n1845 VGND.n1844 194.391
R2812 VGND.n1840 VGND.n1733 194.391
R2813 VGND.n1835 VGND.n1833 194.391
R2814 VGND.n632 VGND.n631 194.391
R2815 VGND.n669 VGND.n668 194.391
R2816 VGND.n674 VGND.n673 194.391
R2817 VGND.n679 VGND.n678 194.391
R2818 VGND.n684 VGND.n683 194.391
R2819 VGND.n689 VGND.n688 194.391
R2820 VGND.n694 VGND.n693 194.391
R2821 VGND.n699 VGND.n698 194.391
R2822 VGND.n704 VGND.n703 194.391
R2823 VGND.n709 VGND.n708 194.391
R2824 VGND.n714 VGND.n713 194.391
R2825 VGND.n719 VGND.n718 194.391
R2826 VGND.n666 VGND.n665 194.391
R2827 VGND.n724 VGND.n723 194.391
R2828 VGND.n2859 VGND.n2858 194.391
R2829 VGND.n2866 VGND.n252 194.391
R2830 VGND.n879 VGND.n878 194.391
R2831 VGND.n1352 VGND.n1351 194.391
R2832 VGND.n874 VGND.n873 194.391
R2833 VGND.n869 VGND.n807 194.391
R2834 VGND.n811 VGND.n809 194.391
R2835 VGND.n823 VGND.n822 194.391
R2836 VGND.n828 VGND.n827 194.391
R2837 VGND.n833 VGND.n832 194.391
R2838 VGND.n838 VGND.n837 194.391
R2839 VGND.n843 VGND.n842 194.391
R2840 VGND.n848 VGND.n847 194.391
R2841 VGND.n819 VGND.n818 194.391
R2842 VGND.n853 VGND.n852 194.391
R2843 VGND.n734 VGND.n733 194.391
R2844 VGND.n1661 VGND.n1660 194.391
R2845 VGND.n1656 VGND.n736 194.391
R2846 VGND.n800 VGND.n799 194.391
R2847 VGND.n1390 VGND.n1389 194.391
R2848 VGND.n1395 VGND.n1394 194.391
R2849 VGND.n804 VGND.n803 194.391
R2850 VGND.n1490 VGND.n1489 194.391
R2851 VGND.n776 VGND.n775 194.391
R2852 VGND.n1516 VGND.n1515 194.391
R2853 VGND.n768 VGND.n767 194.391
R2854 VGND.n1542 VGND.n1541 194.391
R2855 VGND.n1547 VGND.n1546 194.391
R2856 VGND.n760 VGND.n759 194.391
R2857 VGND.n1552 VGND.n1551 194.391
R2858 VGND.n1632 VGND.n1631 194.391
R2859 VGND.n1637 VGND.n1636 194.391
R2860 VGND.n1642 VGND.n1641 194.391
R2861 VGND.n1649 VGND.n739 194.391
R2862 VGND.n797 VGND.n796 194.391
R2863 VGND.n1410 VGND.n1409 194.391
R2864 VGND.n794 VGND.n793 194.391
R2865 VGND.n1477 VGND.n1476 194.391
R2866 VGND.n780 VGND.n779 194.391
R2867 VGND.n1503 VGND.n1502 194.391
R2868 VGND.n772 VGND.n771 194.391
R2869 VGND.n1529 VGND.n1528 194.391
R2870 VGND.n764 VGND.n763 194.391
R2871 VGND.n1566 VGND.n1565 194.391
R2872 VGND.n755 VGND.n754 194.391
R2873 VGND.n1581 VGND.n1580 194.391
R2874 VGND.n1576 VGND.n1575 194.391
R2875 VGND.n1571 VGND.n1570 194.391
R2876 VGND.n2884 VGND.n2883 194.391
R2877 VGND.n2891 VGND.n239 194.391
R2878 VGND.n882 VGND.n881 194.391
R2879 VGND.n884 VGND.n883 194.391
R2880 VGND.n1423 VGND.n1422 194.391
R2881 VGND.n1428 VGND.n1427 194.391
R2882 VGND.n1433 VGND.n1432 194.391
R2883 VGND.n1438 VGND.n1437 194.391
R2884 VGND.n1443 VGND.n1442 194.391
R2885 VGND.n1448 VGND.n1447 194.391
R2886 VGND.n1453 VGND.n1452 194.391
R2887 VGND.n790 VGND.n789 194.391
R2888 VGND.n1458 VGND.n1457 194.391
R2889 VGND.n1595 VGND.n1594 194.391
R2890 VGND.n1600 VGND.n1599 194.391
R2891 VGND.n749 VGND.n748 194.391
R2892 VGND.n1613 VGND.n1612 194.391
R2893 VGND.n1608 VGND.n1604 194.391
R2894 VGND.n1024 VGND.n1023 194.391
R2895 VGND.n1031 VGND.n1030 194.391
R2896 VGND.n1036 VGND.n1035 194.391
R2897 VGND.n1028 VGND.n1027 194.391
R2898 VGND.n1094 VGND.n1093 194.391
R2899 VGND.n1089 VGND.n1088 194.391
R2900 VGND.n1084 VGND.n1083 194.391
R2901 VGND.n1079 VGND.n1078 194.391
R2902 VGND.n1074 VGND.n1073 194.391
R2903 VGND.n1069 VGND.n1040 194.391
R2904 VGND.n1044 VGND.n1042 194.391
R2905 VGND.n1052 VGND.n1051 194.391
R2906 VGND.n1057 VGND.n1056 194.391
R2907 VGND.n1048 VGND.n1047 194.391
R2908 VGND.n2904 VGND.n2903 194.391
R2909 VGND.n2911 VGND.n227 194.391
R2910 VGND.n1014 VGND.n1013 194.391
R2911 VGND.n927 VGND.n926 194.391
R2912 VGND.n2606 VGND.n2605 161.308
R2913 VGND.n2603 VGND.n2602 161.308
R2914 VGND.n2600 VGND.n2599 161.308
R2915 VGND.n2597 VGND.n2596 161.308
R2916 VGND.n2594 VGND.n2593 161.308
R2917 VGND.n2591 VGND.n2590 161.308
R2918 VGND.n2588 VGND.n2587 161.308
R2919 VGND.n2585 VGND.n2584 161.308
R2920 VGND.n2582 VGND.n2581 161.308
R2921 VGND.n2579 VGND.n2578 161.308
R2922 VGND.n2576 VGND.n2575 161.308
R2923 VGND.n2573 VGND.n2572 161.308
R2924 VGND.n2570 VGND.n2569 161.308
R2925 VGND.n2567 VGND.n2566 161.308
R2926 VGND.n2564 VGND.n2563 161.308
R2927 VGND.n2605 VGND.t2696 159.978
R2928 VGND.n2602 VGND.t2699 159.978
R2929 VGND.n2599 VGND.t2694 159.978
R2930 VGND.n2596 VGND.t2689 159.978
R2931 VGND.n2593 VGND.t2695 159.978
R2932 VGND.n2590 VGND.t2702 159.978
R2933 VGND.n2587 VGND.t2698 159.978
R2934 VGND.n2584 VGND.t2692 159.978
R2935 VGND.n2581 VGND.t2688 159.978
R2936 VGND.n2578 VGND.t2690 159.978
R2937 VGND.n2575 VGND.t2701 159.978
R2938 VGND.n2572 VGND.t2693 159.978
R2939 VGND.n2569 VGND.t2700 159.978
R2940 VGND.n2566 VGND.t2697 159.978
R2941 VGND.n2563 VGND.t2703 159.978
R2942 VGND.n123 VGND.t1248 159.315
R2943 VGND.n2216 VGND.t2080 159.315
R2944 VGND.n1132 VGND.t1847 158.361
R2945 VGND.n2999 VGND.t1454 158.361
R2946 VGND.n121 VGND.t1246 157.291
R2947 VGND.n544 VGND.t2078 157.291
R2948 VGND.n68 VGND.t2286 156.915
R2949 VGND.n506 VGND.t1184 156.915
R2950 VGND.n68 VGND.t2287 156.915
R2951 VGND.n506 VGND.t1182 156.915
R2952 VGND.n36 VGND.t1817 154.131
R2953 VGND.n123 VGND.t1591 154.131
R2954 VGND.n128 VGND.t95 154.131
R2955 VGND.n128 VGND.t2 154.131
R2956 VGND.n508 VGND.t1462 154.131
R2957 VGND.n508 VGND.t227 154.131
R2958 VGND.n2216 VGND.t255 154.131
R2959 VGND.n541 VGND.t906 154.131
R2960 VGND.n3005 VGND.t787 153.631
R2961 VGND.n60 VGND.t807 153.631
R2962 VGND.n160 VGND.t2284 153.631
R2963 VGND.n2255 VGND.t1181 153.631
R2964 VGND.n2222 VGND.t1852 153.631
R2965 VGND.n1360 VGND.t2076 153.631
R2966 VGND.n59 VGND.t2540 152.757
R2967 VGND.n2221 VGND.t1582 152.757
R2968 VGND.n92 VGND.t2291 152.381
R2969 VGND.n2211 VGND.t1179 152.381
R2970 VGND.n2181 VGND.n2180 152.174
R2971 VGND.n167 VGND.t2294 150.922
R2972 VGND.n167 VGND.t2289 150.922
R2973 VGND.n475 VGND.t1183 150.922
R2974 VGND.n475 VGND.t1177 150.922
R2975 VGND.n166 VGND.t97 150.922
R2976 VGND.n67 VGND.t935 150.922
R2977 VGND.n135 VGND.t2680 150.922
R2978 VGND.n474 VGND.t2096 150.922
R2979 VGND.n2253 VGND.t2074 150.922
R2980 VGND.n505 VGND.t1457 150.922
R2981 VGND.n166 VGND.t2577 150.922
R2982 VGND.n67 VGND.t345 150.922
R2983 VGND.n135 VGND.t376 150.922
R2984 VGND.n474 VGND.t2687 150.922
R2985 VGND.n2253 VGND.t2103 150.922
R2986 VGND.n505 VGND.t143 150.922
R2987 VGND.n3004 VGND.t384 147.411
R2988 VGND.n159 VGND.t2293 147.411
R2989 VGND.n2254 VGND.t1180 147.411
R2990 VGND.n1359 VGND.t1843 147.411
R2991 VGND.n115 VGND.t1361 146.964
R2992 VGND.n545 VGND.t1174 146.964
R2993 VGND.n2605 VGND.t981 143.911
R2994 VGND.n2602 VGND.t1056 143.911
R2995 VGND.n2599 VGND.t963 143.911
R2996 VGND.n2596 VGND.t1005 143.911
R2997 VGND.n2593 VGND.t1077 143.911
R2998 VGND.n2590 VGND.t984 143.911
R2999 VGND.n2587 VGND.t957 143.911
R3000 VGND.n2584 VGND.t999 143.911
R3001 VGND.n2581 VGND.t1011 143.911
R3002 VGND.n2578 VGND.t939 143.911
R3003 VGND.n2575 VGND.t1035 143.911
R3004 VGND.n2572 VGND.t966 143.911
R3005 VGND.n2569 VGND.t1038 143.911
R3006 VGND.n2566 VGND.t1068 143.911
R3007 VGND.n2563 VGND.t1008 143.911
R3008 VGND.n1388 VGND.n806 143.478
R3009 VGND VGND.t2378 142.089
R3010 VGND.n1021 VGND.t996 119.309
R3011 VGND.n994 VGND.t1032 119.309
R3012 VGND.n2630 VGND.t993 119.309
R3013 VGND.n204 VGND.t1029 119.309
R3014 VGND.n334 VGND.t942 119.309
R3015 VGND.n2626 VGND.t948 119.309
R3016 VGND.n2623 VGND.t954 119.309
R3017 VGND.n2620 VGND.t1041 119.309
R3018 VGND.n2617 VGND.t1047 119.309
R3019 VGND.n2614 VGND.t960 119.309
R3020 VGND.n2611 VGND.t1002 119.309
R3021 VGND.n322 VGND.t1017 119.309
R3022 VGND.n315 VGND.t1053 119.309
R3023 VGND.n306 VGND.t975 119.309
R3024 VGND.n299 VGND.t1020 119.309
R3025 VGND.n2765 VGND.t1059 119.309
R3026 VGND.n290 VGND.t1071 119.309
R3027 VGND.n297 VGND.t987 119.309
R3028 VGND.n1018 VGND.t945 119.309
R3029 VGND.n1015 VGND.t951 119.309
R3030 VGND.n1180 VGND.t969 119.309
R3031 VGND.n1006 VGND.t1044 119.309
R3032 VGND.n1004 VGND.t1050 119.309
R3033 VGND.n1195 VGND.t972 119.309
R3034 VGND.n1212 VGND.t1014 119.309
R3035 VGND.n1000 VGND.t1023 119.309
R3036 VGND.n1253 VGND.t1062 119.309
R3037 VGND.n1256 VGND.t978 119.309
R3038 VGND.n1259 VGND.t1026 119.309
R3039 VGND.n1262 VGND.t1065 119.309
R3040 VGND.n998 VGND.t1074 119.309
R3041 VGND.n1265 VGND.t990 119.309
R3042 VGND.n5 VGND.n3 117.001
R3043 VGND.t303 VGND.n5 117.001
R3044 VGND.n6 VGND.n4 117.001
R3045 VGND.n328 VGND.n6 117.001
R3046 VGND.t2196 VGND.t997 110.535
R3047 VGND.t93 VGND.t2136 110.535
R3048 VGND.t946 VGND.t2130 110.535
R3049 VGND.t2625 VGND.t1596 110.535
R3050 VGND.t2617 VGND.t952 110.535
R3051 VGND.t1530 VGND.t2610 110.535
R3052 VGND.t970 VGND.t2595 110.535
R3053 VGND.t2172 VGND.t671 110.535
R3054 VGND.t2184 VGND.t1045 110.535
R3055 VGND.t1110 VGND.t2124 110.535
R3056 VGND.t1051 VGND.t2108 110.535
R3057 VGND.t2598 VGND.t1131 110.535
R3058 VGND.t2664 VGND.t973 110.535
R3059 VGND.t29 VGND.t2187 110.535
R3060 VGND.t1015 VGND.t2178 110.535
R3061 VGND.t2162 VGND.t237 110.535
R3062 VGND.t2156 VGND.t1024 110.535
R3063 VGND.t662 VGND.t2666 110.535
R3064 VGND.t1063 VGND.t2110 110.535
R3065 VGND.t2599 VGND.t226 110.535
R3066 VGND.t2583 VGND.t979 110.535
R3067 VGND.t563 VGND.t2159 110.535
R3068 VGND.t1027 VGND.t2228 110.535
R3069 VGND.t2147 VGND.t680 110.535
R3070 VGND.t2660 VGND.t1066 110.535
R3071 VGND.t1338 VGND.t2653 110.535
R3072 VGND.t1075 VGND.t2648 110.535
R3073 VGND.t2230 VGND.t229 110.535
R3074 VGND.t2626 VGND.t991 110.535
R3075 VGND.t467 VGND.t2209 110.535
R3076 VGND.t1033 VGND.t2143 110.535
R3077 VGND.t2650 VGND.t727 110.535
R3078 VGND.t1165 VGND.t1175 92.4699
R3079 VGND.t1175 VGND.t1172 92.4699
R3080 VGND.t1172 VGND.t1176 92.4699
R3081 VGND.t1176 VGND.t1470 92.4699
R3082 VGND.t1470 VGND.t629 92.4699
R3083 VGND.t629 VGND.t1478 92.4699
R3084 VGND.t1478 VGND.t1448 92.4699
R3085 VGND VGND.n806 80.9529
R3086 VGND VGND.n806 75.1009
R3087 VGND.n1337 VGND 74.8566
R3088 VGND.t1448 VGND 70.4533
R3089 VGND.n2285 VGND 58.8055
R3090 VGND.n2284 VGND 58.8055
R3091 VGND.n2250 VGND 58.8055
R3092 VGND.n2248 VGND 58.8055
R3093 VGND.n1386 VGND 58.8055
R3094 VGND.n2348 VGND.n2347 53.1823
R3095 VGND.n2349 VGND.n2348 53.1823
R3096 VGND.n3021 VGND.n3020 53.1823
R3097 VGND.n3020 VGND.n3019 53.1823
R3098 VGND.t1368 VGND.t2376 50.5752
R3099 VGND.t1364 VGND.t2350 50.5752
R3100 VGND.t1358 VGND.t2387 50.5752
R3101 VGND.t1360 VGND.t2330 50.5752
R3102 VGND.t1173 VGND.t1468 50.5752
R3103 VGND.t1170 VGND.t627 50.5752
R3104 VGND.t1168 VGND.t408 50.5752
R3105 VGND.t1166 VGND.t42 50.5752
R3106 VGND VGND.n2981 43.2063
R3107 VGND VGND.n18 43.2063
R3108 VGND VGND.n2951 43.2063
R3109 VGND VGND.n44 43.2063
R3110 VGND.n2347 VGND.n2346 40.6593
R3111 VGND.n886 VGND.t2161 34.8005
R3112 VGND.n886 VGND.t2670 34.8005
R3113 VGND.n889 VGND.t2668 34.8005
R3114 VGND.n889 VGND.t2589 34.8005
R3115 VGND.n893 VGND.t2586 34.8005
R3116 VGND.n893 VGND.t2164 34.8005
R3117 VGND.n930 VGND.t2218 34.8005
R3118 VGND.n930 VGND.t2142 34.8005
R3119 VGND.n935 VGND.t2663 34.8005
R3120 VGND.n935 VGND.t2659 34.8005
R3121 VGND.n940 VGND.t2652 34.8005
R3122 VGND.n940 VGND.t2224 34.8005
R3123 VGND.n945 VGND.t2633 34.8005
R3124 VGND.n945 VGND.t2213 34.8005
R3125 VGND.n950 VGND.t2146 34.8005
R3126 VGND.n950 VGND.t2655 34.8005
R3127 VGND.n955 VGND.t1508 34.8005
R3128 VGND.n955 VGND.t2637 34.8005
R3129 VGND.n960 VGND.t2629 34.8005
R3130 VGND.n960 VGND.t2226 34.8005
R3131 VGND.n965 VGND.t2206 34.8005
R3132 VGND.n965 VGND.t1512 34.8005
R3133 VGND.n970 VGND.t2193 34.8005
R3134 VGND.n970 VGND.t2134 34.8005
R3135 VGND.n975 VGND.t2118 34.8005
R3136 VGND.n975 VGND.t2208 34.8005
R3137 VGND.n980 VGND.t2612 34.8005
R3138 VGND.n980 VGND.t2195 34.8005
R3139 VGND.n985 VGND.t2175 34.8005
R3140 VGND.n985 VGND.t2170 34.8005
R3141 VGND.n996 VGND.t2222 34.8005
R3142 VGND.n996 VGND.t2144 34.8005
R3143 VGND.n1273 VGND.t2635 34.8005
R3144 VGND.n1273 VGND.t2627 34.8005
R3145 VGND.n1230 VGND.t2140 34.8005
R3146 VGND.n1230 VGND.t2649 34.8005
R3147 VGND.n1229 VGND.t2211 34.8005
R3148 VGND.n1229 VGND.t2661 34.8005
R3149 VGND.n1226 VGND.t2646 34.8005
R3150 VGND.n1226 VGND.t2229 34.8005
R3151 VGND.n1224 VGND.t2657 34.8005
R3152 VGND.n1224 VGND.t2584 34.8005
R3153 VGND.n1221 VGND.t2150 34.8005
R3154 VGND.n1221 VGND.t2111 34.8005
R3155 VGND.n1216 VGND.t2582 34.8005
R3156 VGND.n1216 VGND.t2157 34.8005
R3157 VGND.n1002 VGND.t2602 34.8005
R3158 VGND.n1002 VGND.t2179 34.8005
R3159 VGND.n1203 VGND.t2155 34.8005
R3160 VGND.n1203 VGND.t2665 34.8005
R3161 VGND.n1007 VGND.t2177 34.8005
R3162 VGND.n1007 VGND.t2109 34.8005
R3163 VGND.n1184 VGND.t2189 34.8005
R3164 VGND.n1184 VGND.t2185 34.8005
R3165 VGND.n1010 VGND.t2105 34.8005
R3166 VGND.n1010 VGND.t2596 34.8005
R3167 VGND.n1171 VGND.t2129 34.8005
R3168 VGND.n1171 VGND.t2618 34.8005
R3169 VGND.n1012 VGND.t2191 34.8005
R3170 VGND.n1012 VGND.t2131 34.8005
R3171 VGND.n329 VGND.t2216 34.8005
R3172 VGND.n329 VGND.t1521 34.8005
R3173 VGND.n332 VGND.t1519 34.8005
R3174 VGND.n332 VGND.t2644 34.8005
R3175 VGND.n356 VGND.t2642 34.8005
R3176 VGND.n356 VGND.t2220 34.8005
R3177 VGND.n363 VGND.t2620 34.8005
R3178 VGND.n363 VGND.t2200 34.8005
R3179 VGND.n366 VGND.t1517 34.8005
R3180 VGND.n366 VGND.t1514 34.8005
R3181 VGND.n374 VGND.t1506 34.8005
R3182 VGND.n374 VGND.t2622 34.8005
R3183 VGND.n377 VGND.t2120 34.8005
R3184 VGND.n377 VGND.t2608 34.8005
R3185 VGND.n385 VGND.t2204 34.8005
R3186 VGND.n385 VGND.t1510 34.8005
R3187 VGND.n324 VGND.t2181 34.8005
R3188 VGND.n324 VGND.t2122 34.8005
R3189 VGND.n313 VGND.t2116 34.8005
R3190 VGND.n313 VGND.t2624 34.8005
R3191 VGND.n308 VGND.t2604 34.8005
R3192 VGND.n308 VGND.t2183 34.8005
R3193 VGND.n310 VGND.t2592 34.8005
R3194 VGND.n310 VGND.t2168 34.8005
R3195 VGND.n2729 VGND.t2152 34.8005
R3196 VGND.n2729 VGND.t2606 34.8005
R3197 VGND.n292 VGND.t2672 34.8005
R3198 VGND.n292 VGND.t2594 34.8005
R3199 VGND.n295 VGND.t2580 34.8005
R3200 VGND.n295 VGND.t2232 34.8005
R3201 VGND.n202 VGND.t2166 34.8005
R3202 VGND.n202 VGND.t2107 34.8005
R3203 VGND.n395 VGND.t983 34.8005
R3204 VGND.n395 VGND.t1437 34.8005
R3205 VGND.n2637 VGND.t1157 34.8005
R3206 VGND.n2637 VGND.t783 34.8005
R3207 VGND.n2642 VGND.t1609 34.8005
R3208 VGND.n2642 VGND.t2568 34.8005
R3209 VGND.n2647 VGND.t557 34.8005
R3210 VGND.n2647 VGND.t2566 34.8005
R3211 VGND.n2652 VGND.t1555 34.8005
R3212 VGND.n2652 VGND.t1435 34.8005
R3213 VGND.n2657 VGND.t263 34.8005
R3214 VGND.n2657 VGND.t1412 34.8005
R3215 VGND.n2662 VGND.t733 34.8005
R3216 VGND.n2662 VGND.t2576 34.8005
R3217 VGND.n2667 VGND.t571 34.8005
R3218 VGND.n2667 VGND.t1433 34.8005
R3219 VGND.n392 VGND.t677 34.8005
R3220 VGND.n392 VGND.t1431 34.8005
R3221 VGND.n2713 VGND.t218 34.8005
R3222 VGND.n2713 VGND.t1414 34.8005
R3223 VGND.n318 VGND.t1217 34.8005
R3224 VGND.n318 VGND.t2564 34.8005
R3225 VGND.n2746 VGND.t1747 34.8005
R3226 VGND.n2746 VGND.t1439 34.8005
R3227 VGND.n302 VGND.t2425 34.8005
R3228 VGND.n302 VGND.t2574 34.8005
R3229 VGND.n2751 VGND.t915 34.8005
R3230 VGND.n2751 VGND.t2572 34.8005
R3231 VGND.n2786 VGND.t466 34.8005
R3232 VGND.n2786 VGND.t2570 34.8005
R3233 VGND.n285 VGND.t290 34.8005
R3234 VGND.n285 VGND.t1429 34.8005
R3235 VGND.n399 VGND.t1058 34.8005
R3236 VGND.n399 VGND.t701 34.8005
R3237 VGND.n2341 VGND.t833 34.8005
R3238 VGND.n2341 VGND.t1113 34.8005
R3239 VGND.n2336 VGND.t374 34.8005
R3240 VGND.n2336 VGND.t473 34.8005
R3241 VGND.n2331 VGND.t115 34.8005
R3242 VGND.n2331 VGND.t471 34.8005
R3243 VGND.n2326 VGND.t1547 34.8005
R3244 VGND.n2326 VGND.t699 34.8005
R3245 VGND.n2321 VGND.t1751 34.8005
R3246 VGND.n2321 VGND.t1196 34.8005
R3247 VGND.n2316 VGND.t301 34.8005
R3248 VGND.n2316 VGND.t1194 34.8005
R3249 VGND.n2311 VGND.t1670 34.8005
R3250 VGND.n2311 VGND.t1119 34.8005
R3251 VGND.n2306 VGND.t334 34.8005
R3252 VGND.n2306 VGND.t1117 34.8005
R3253 VGND.n2301 VGND.t1842 34.8005
R3254 VGND.n2301 VGND.t1198 34.8005
R3255 VGND.n2296 VGND.t457 34.8005
R3256 VGND.n2296 VGND.t705 34.8005
R3257 VGND.n2291 VGND.t710 34.8005
R3258 VGND.n2291 VGND.t703 34.8005
R3259 VGND.n2286 VGND.t1616 34.8005
R3260 VGND.n2286 VGND.t1192 34.8005
R3261 VGND.n413 VGND.t1261 34.8005
R3262 VGND.n413 VGND.t1190 34.8005
R3263 VGND.n2539 VGND.t33 34.8005
R3264 VGND.n2539 VGND.t475 34.8005
R3265 VGND.n416 VGND.t2434 34.8005
R3266 VGND.n416 VGND.t1115 34.8005
R3267 VGND.n468 VGND.t965 34.8005
R3268 VGND.n468 VGND.t1788 34.8005
R3269 VGND.n470 VGND.t82 34.8005
R3270 VGND.n470 VGND.t1523 34.8005
R3271 VGND.n2375 VGND.t1983 34.8005
R3272 VGND.n2375 VGND.t1796 34.8005
R3273 VGND.n458 VGND.t606 34.8005
R3274 VGND.n458 VGND.t1794 34.8005
R3275 VGND.n2401 VGND.t1562 34.8005
R3276 VGND.n2401 VGND.t1786 34.8005
R3277 VGND.n450 VGND.t1825 34.8005
R3278 VGND.n450 VGND.t1328 34.8005
R3279 VGND.n2427 VGND.t321 34.8005
R3280 VGND.n2427 VGND.t1326 34.8005
R3281 VGND.n442 VGND.t130 34.8005
R3282 VGND.n442 VGND.t1529 34.8005
R3283 VGND.n2453 VGND.t338 34.8005
R3284 VGND.n2453 VGND.t1527 34.8005
R3285 VGND.n434 VGND.t667 34.8005
R3286 VGND.n434 VGND.t1330 34.8005
R3287 VGND.n2479 VGND.t435 34.8005
R3288 VGND.n2479 VGND.t1792 34.8005
R3289 VGND.n426 VGND.t1741 34.8005
R3290 VGND.n426 VGND.t1790 34.8005
R3291 VGND.n2510 VGND.t186 34.8005
R3292 VGND.n2510 VGND.t1324 34.8005
R3293 VGND.n2515 VGND.t921 34.8005
R3294 VGND.n2515 VGND.t1800 34.8005
R3295 VGND.n2520 VGND.t366 34.8005
R3296 VGND.n2520 VGND.t1798 34.8005
R3297 VGND.n418 VGND.t511 34.8005
R3298 VGND.n418 VGND.t1525 34.8005
R3299 VGND.n465 VGND.t1007 34.8005
R3300 VGND.n465 VGND.t1272 34.8005
R3301 VGND.n2362 VGND.t837 34.8005
R3302 VGND.n2362 VGND.t2090 34.8005
R3303 VGND.n462 VGND.t1833 34.8005
R3304 VGND.n462 VGND.t1103 34.8005
R3305 VGND.n2388 VGND.t530 34.8005
R3306 VGND.n2388 VGND.t1278 34.8005
R3307 VGND.n454 VGND.t10 34.8005
R3308 VGND.n454 VGND.t483 34.8005
R3309 VGND.n2414 VGND.t1316 34.8005
R3310 VGND.n2414 VGND.t2086 34.8005
R3311 VGND.n446 VGND.t693 34.8005
R3312 VGND.n446 VGND.t2084 34.8005
R3313 VGND.n2440 VGND.t551 34.8005
R3314 VGND.n2440 VGND.t481 34.8005
R3315 VGND.n438 VGND.t317 34.8005
R3316 VGND.n438 VGND.t479 34.8005
R3317 VGND.n2466 VGND.t599 34.8005
R3318 VGND.n2466 VGND.t2088 34.8005
R3319 VGND.n430 VGND.t165 34.8005
R3320 VGND.n430 VGND.t1276 34.8005
R3321 VGND.n2492 VGND.t1127 34.8005
R3322 VGND.n2492 VGND.t1274 34.8005
R3323 VGND.n422 VGND.t1221 34.8005
R3324 VGND.n422 VGND.t1109 34.8005
R3325 VGND.n2497 VGND.t2683 34.8005
R3326 VGND.n2497 VGND.t1107 34.8005
R3327 VGND.n2808 VGND.t1352 34.8005
R3328 VGND.n2808 VGND.t1105 34.8005
R3329 VGND.n276 VGND.t282 34.8005
R3330 VGND.n276 VGND.t477 34.8005
R3331 VGND.n624 VGND.t1079 34.8005
R3332 VGND.n624 VGND.t2528 34.8005
R3333 VGND.n1909 VGND.t1149 34.8005
R3334 VGND.n1909 VGND.t769 34.8005
R3335 VGND.n621 VGND.t2678 34.8005
R3336 VGND.n621 VGND.t1802 34.8005
R3337 VGND.n1920 VGND.t109 34.8005
R3338 VGND.n1920 VGND.t1410 34.8005
R3339 VGND.n618 VGND.t1540 34.8005
R3340 VGND.n618 VGND.t2526 34.8005
R3341 VGND.n1931 VGND.t1700 34.8005
R3342 VGND.n1931 VGND.t765 34.8005
R3343 VGND.n615 VGND.t297 34.8005
R3344 VGND.n615 VGND.t763 34.8005
R3345 VGND.n1942 VGND.t137 34.8005
R3346 VGND.n1942 VGND.t2524 34.8005
R3347 VGND.n612 VGND.t643 34.8005
R3348 VGND.n612 VGND.t2522 34.8005
R3349 VGND.n1953 VGND.t1138 34.8005
R3350 VGND.n1953 VGND.t767 34.8005
R3351 VGND.n609 VGND.t443 34.8005
R3352 VGND.n609 VGND.t1408 34.8005
R3353 VGND.n1964 VGND.t1813 34.8005
R3354 VGND.n1964 VGND.t1406 34.8005
R3355 VGND.n606 VGND.t2422 34.8005
R3356 VGND.n606 VGND.t761 34.8005
R3357 VGND.n1975 VGND.t1255 34.8005
R3358 VGND.n1975 VGND.t759 34.8005
R3359 VGND.n1980 VGND.t25 34.8005
R3360 VGND.n1980 VGND.t1804 34.8005
R3361 VGND.n605 VGND.t519 34.8005
R3362 VGND.n605 VGND.t2520 34.8005
R3363 VGND.n589 VGND.t986 34.8005
R3364 VGND.n589 VGND.t1784 34.8005
R3365 VGND.n595 VGND.t1155 34.8005
R3366 VGND.n595 VGND.t1774 34.8005
R3367 VGND.n592 VGND.t1607 34.8005
R3368 VGND.n592 VGND.t877 34.8005
R3369 VGND.n2054 VGND.t554 34.8005
R3370 VGND.n2054 VGND.t875 34.8005
R3371 VGND.n2049 VGND.t1553 34.8005
R3372 VGND.n2049 VGND.t1782 34.8005
R3373 VGND.n2044 VGND.t261 34.8005
R3374 VGND.n2044 VGND.t1232 34.8005
R3375 VGND.n2039 VGND.t731 34.8005
R3376 VGND.n2039 VGND.t1230 34.8005
R3377 VGND.n2034 VGND.t569 34.8005
R3378 VGND.n2034 VGND.t1780 34.8005
R3379 VGND.n2029 VGND.t675 34.8005
R3380 VGND.n2029 VGND.t1778 34.8005
R3381 VGND.n2024 VGND.t216 34.8005
R3382 VGND.n2024 VGND.t1234 34.8005
R3383 VGND.n2019 VGND.t1214 34.8005
R3384 VGND.n2019 VGND.t873 34.8005
R3385 VGND.n2014 VGND.t1745 34.8005
R3386 VGND.n2014 VGND.t871 34.8005
R3387 VGND.n2009 VGND.t1219 34.8005
R3388 VGND.n2009 VGND.t1228 34.8005
R3389 VGND.n2004 VGND.t913 34.8005
R3390 VGND.n2004 VGND.t881 34.8005
R3391 VGND.n600 VGND.t463 34.8005
R3392 VGND.n600 VGND.t879 34.8005
R3393 VGND.n1993 VGND.t288 34.8005
R3394 VGND.n1993 VGND.t1776 34.8005
R3395 VGND.n586 VGND.t959 34.8005
R3396 VGND.n586 VGND.t1494 34.8005
R3397 VGND.n2068 VGND.t623 34.8005
R3398 VGND.n2068 VGND.t2554 34.8005
R3399 VGND.n2073 VGND.t1985 34.8005
R3400 VGND.n2073 VGND.t378 34.8005
R3401 VGND.n2078 VGND.t604 34.8005
R3402 VGND.n2078 VGND.t1500 34.8005
R3403 VGND.n2083 VGND.t1236 34.8005
R3404 VGND.n2083 VGND.t1492 34.8005
R3405 VGND.n2088 VGND.t1827 34.8005
R3406 VGND.n2088 VGND.t2550 34.8005
R3407 VGND.n2093 VGND.t323 34.8005
R3408 VGND.n2093 VGND.t2548 34.8005
R3409 VGND.n2098 VGND.t132 34.8005
R3410 VGND.n2098 VGND.t1490 34.8005
R3411 VGND.n2103 VGND.t340 34.8005
R3412 VGND.n2103 VGND.t1488 34.8005
R3413 VGND.n2108 VGND.t669 34.8005
R3414 VGND.n2108 VGND.t2552 34.8005
R3415 VGND.n2113 VGND.t437 34.8005
R3416 VGND.n2113 VGND.t1498 34.8005
R3417 VGND.n2118 VGND.t1743 34.8005
R3418 VGND.n2118 VGND.t1496 34.8005
R3419 VGND.n583 VGND.t188 34.8005
R3420 VGND.n583 VGND.t2546 34.8005
R3421 VGND.n2123 VGND.t923 34.8005
R3422 VGND.n2123 VGND.t382 34.8005
R3423 VGND.n2833 VGND.t368 34.8005
R3424 VGND.n2833 VGND.t380 34.8005
R3425 VGND.n264 VGND.t513 34.8005
R3426 VGND.n264 VGND.t1486 34.8005
R3427 VGND.n546 VGND.t1001 34.8005
R3428 VGND.n546 VGND.t653 34.8005
R3429 VGND.n549 VGND.t839 34.8005
R3430 VGND.n549 VGND.t1904 34.8005
R3431 VGND.n1755 VGND.t1835 34.8005
R3432 VGND.n1755 VGND.t894 34.8005
R3433 VGND.n1760 VGND.t528 34.8005
R3434 VGND.n1760 VGND.t892 34.8005
R3435 VGND.n1751 VGND.t12 34.8005
R3436 VGND.n1751 VGND.t651 34.8005
R3437 VGND.n1771 VGND.t1600 34.8005
R3438 VGND.n1771 VGND.t1101 34.8005
R3439 VGND.n1748 VGND.t695 34.8005
R3440 VGND.n1748 VGND.t1099 34.8005
R3441 VGND.n1782 VGND.t565 34.8005
R3442 VGND.n1782 VGND.t649 34.8005
R3443 VGND.n1745 VGND.t319 34.8005
R3444 VGND.n1745 VGND.t777 34.8005
R3445 VGND.n1793 VGND.t601 34.8005
R3446 VGND.n1793 VGND.t1902 34.8005
R3447 VGND.n1742 VGND.t1209 34.8005
R3448 VGND.n1742 VGND.t890 34.8005
R3449 VGND.n1804 VGND.t1129 34.8005
R3450 VGND.n1804 VGND.t655 34.8005
R3451 VGND.n1739 VGND.t1223 34.8005
R3452 VGND.n1739 VGND.t1097 34.8005
R3453 VGND.n1815 VGND.t2685 34.8005
R3454 VGND.n1815 VGND.t1095 34.8005
R3455 VGND.n1820 VGND.t1354 34.8005
R3456 VGND.n1820 VGND.t896 34.8005
R3457 VGND.n1738 VGND.t284 34.8005
R3458 VGND.n1738 VGND.t775 34.8005
R3459 VGND.n627 VGND.t1013 34.8005
R3460 VGND.n627 VGND.t312 34.8005
R3461 VGND.n1677 VGND.t1161 34.8005
R3462 VGND.n1677 VGND.t2402 34.8005
R3463 VGND.n1674 VGND.t592 34.8005
R3464 VGND.n1674 VGND.t900 34.8005
R3465 VGND.n1688 VGND.t534 34.8005
R3466 VGND.n1688 VGND.t1336 34.8005
R3467 VGND.n1693 VGND.t6 34.8005
R3468 VGND.n1693 VGND.t310 34.8005
R3469 VGND.n1698 VGND.t1310 34.8005
R3470 VGND.n1698 VGND.t2398 34.8005
R3471 VGND.n1703 VGND.t691 34.8005
R3472 VGND.n1703 VGND.t2396 34.8005
R3473 VGND.n1708 VGND.t547 34.8005
R3474 VGND.n1708 VGND.t308 34.8005
R3475 VGND.n1713 VGND.t20 34.8005
R3476 VGND.n1713 VGND.t306 34.8005
R3477 VGND.n1718 VGND.t1587 34.8005
R3478 VGND.n1718 VGND.t2400 34.8005
R3479 VGND.n1723 VGND.t163 34.8005
R3480 VGND.n1723 VGND.t1334 34.8005
R3481 VGND.n1728 VGND.t1125 34.8005
R3482 VGND.n1728 VGND.t1332 34.8005
R3483 VGND.n1671 VGND.t1350 34.8005
R3484 VGND.n1671 VGND.t2394 34.8005
R3485 VGND.n1844 VGND.t2000 34.8005
R3486 VGND.n1844 VGND.t904 34.8005
R3487 VGND.n1733 VGND.t1378 34.8005
R3488 VGND.n1733 VGND.t902 34.8005
R3489 VGND.n1833 VGND.t180 34.8005
R3490 VGND.n1833 VGND.t2530 34.8005
R3491 VGND.n631 VGND.t941 34.8005
R3492 VGND.n631 VGND.t1769 34.8005
R3493 VGND.n668 VGND.t1147 34.8005
R3494 VGND.n668 VGND.t1759 34.8005
R3495 VGND.n673 VGND.t2676 34.8005
R3496 VGND.n673 VGND.t1713 34.8005
R3497 VGND.n678 VGND.t111 34.8005
R3498 VGND.n678 VGND.t1711 34.8005
R3499 VGND.n683 VGND.t1538 34.8005
R3500 VGND.n683 VGND.t1767 34.8005
R3501 VGND.n688 VGND.t1978 34.8005
R3502 VGND.n688 VGND.t1755 34.8005
R3503 VGND.n693 VGND.t329 34.8005
R3504 VGND.n693 VGND.t127 34.8005
R3505 VGND.n698 VGND.t135 34.8005
R3506 VGND.n698 VGND.t1765 34.8005
R3507 VGND.n703 VGND.t641 34.8005
R3508 VGND.n703 VGND.t1763 34.8005
R3509 VGND.n708 VGND.t1136 34.8005
R3510 VGND.n708 VGND.t1757 34.8005
R3511 VGND.n713 VGND.t441 34.8005
R3512 VGND.n713 VGND.t1709 34.8005
R3513 VGND.n718 VGND.t1811 34.8005
R3514 VGND.n718 VGND.t1707 34.8005
R3515 VGND.n665 VGND.t2420 34.8005
R3516 VGND.n665 VGND.t125 34.8005
R3517 VGND.n723 VGND.t1253 34.8005
R3518 VGND.n723 VGND.t123 34.8005
R3519 VGND.n2858 VGND.t23 34.8005
R3520 VGND.n2858 VGND.t121 34.8005
R3521 VGND.n252 VGND.t517 34.8005
R3522 VGND.n252 VGND.t1761 34.8005
R3523 VGND.n878 VGND.t1037 34.8005
R3524 VGND.n878 VGND.t814 34.8005
R3525 VGND.n1351 VGND.t755 34.8005
R3526 VGND.n1351 VGND.t400 34.8005
R3527 VGND.n873 VGND.t1604 34.8005
R3528 VGND.n873 VGND.t822 34.8005
R3529 VGND.n807 VGND.t521 34.8005
R3530 VGND.n807 VGND.t820 34.8005
R3531 VGND.n809 VGND.t1443 34.8005
R3532 VGND.n809 VGND.t812 34.8005
R3533 VGND.n822 VGND.t1308 34.8005
R3534 VGND.n822 VGND.t396 34.8005
R3535 VGND.n827 VGND.t1084 34.8005
R3536 VGND.n827 VGND.t394 34.8005
R3537 VGND.n832 VGND.t540 34.8005
R3538 VGND.n832 VGND.t406 34.8005
R3539 VGND.n837 VGND.t722 34.8005
R3540 VGND.n837 VGND.t404 34.8005
R3541 VGND.n842 VGND.t211 34.8005
R3542 VGND.n842 VGND.t398 34.8005
R3543 VGND.n847 VGND.t157 34.8005
R3544 VGND.n847 VGND.t818 34.8005
R3545 VGND.n818 VGND.t1318 34.8005
R3546 VGND.n818 VGND.t816 34.8005
R3547 VGND.n852 VGND.t1244 34.8005
R3548 VGND.n852 VGND.t392 34.8005
R3549 VGND.n733 VGND.t1993 34.8005
R3550 VGND.n733 VGND.t390 34.8005
R3551 VGND.n1660 VGND.t1536 34.8005
R3552 VGND.n1660 VGND.t824 34.8005
R3553 VGND.n736 VGND.t172 34.8005
R3554 VGND.n736 VGND.t402 34.8005
R3555 VGND.n799 VGND.t968 34.8005
R3556 VGND.n799 VGND.t424 34.8005
R3557 VGND.n1389 VGND.t80 34.8005
R3558 VGND.n1389 VGND.t2413 34.8005
R3559 VGND.n1394 VGND.t1981 34.8005
R3560 VGND.n1394 VGND.t1569 34.8005
R3561 VGND.n803 VGND.t809 34.8005
R3562 VGND.n803 VGND.t430 34.8005
R3563 VGND.n1489 VGND.t1560 34.8005
R3564 VGND.n1489 VGND.t422 34.8005
R3565 VGND.n775 VGND.t1823 34.8005
R3566 VGND.n775 VGND.t2409 34.8005
R3567 VGND.n1515 VGND.t737 34.8005
R3568 VGND.n1515 VGND.t2407 34.8005
R3569 VGND.n767 VGND.t575 34.8005
R3570 VGND.n767 VGND.t420 34.8005
R3571 VGND.n1541 VGND.t336 34.8005
R3572 VGND.n1541 VGND.t418 34.8005
R3573 VGND.n1546 VGND.t665 34.8005
R3574 VGND.n1546 VGND.t2411 34.8005
R3575 VGND.n759 VGND.t2544 34.8005
R3576 VGND.n759 VGND.t428 34.8005
R3577 VGND.n1551 VGND.t1739 34.8005
R3578 VGND.n1551 VGND.t426 34.8005
R3579 VGND.n1631 VGND.t184 34.8005
R3580 VGND.n1631 VGND.t2405 34.8005
R3581 VGND.n1636 VGND.t919 34.8005
R3582 VGND.n1636 VGND.t1573 34.8005
R3583 VGND.n1641 VGND.t364 34.8005
R3584 VGND.n1641 VGND.t1571 34.8005
R3585 VGND.n739 VGND.t509 34.8005
R3586 VGND.n739 VGND.t2415 34.8005
R3587 VGND.n796 VGND.t1040 34.8005
R3588 VGND.n796 VGND.t2450 34.8005
R3589 VGND.n1409 VGND.t753 34.8005
R3590 VGND.n1409 VGND.t743 34.8005
R3591 VGND.n793 VGND.t1602 34.8005
R3592 VGND.n793 VGND.t613 34.8005
R3593 VGND.n1476 VGND.t523 34.8005
R3594 VGND.n1476 VGND.t611 34.8005
R3595 VGND.n779 VGND.t1441 34.8005
R3596 VGND.n779 VGND.t751 34.8005
R3597 VGND.n1502 VGND.t1306 34.8005
R3598 VGND.n1502 VGND.t739 34.8005
R3599 VGND.n771 VGND.t1082 34.8005
R3600 VGND.n771 VGND.t621 34.8005
R3601 VGND.n1528 VGND.t538 34.8005
R3602 VGND.n1528 VGND.t749 34.8005
R3603 VGND.n763 VGND.t720 34.8005
R3604 VGND.n763 VGND.t747 34.8005
R3605 VGND.n1565 VGND.t209 34.8005
R3606 VGND.n1565 VGND.t741 34.8005
R3607 VGND.n754 VGND.t155 34.8005
R3608 VGND.n754 VGND.t2454 34.8005
R3609 VGND.n1580 VGND.t1268 34.8005
R3610 VGND.n1580 VGND.t2452 34.8005
R3611 VGND.n1575 VGND.t1242 34.8005
R3612 VGND.n1575 VGND.t619 34.8005
R3613 VGND.n1570 VGND.t1991 34.8005
R3614 VGND.n1570 VGND.t617 34.8005
R3615 VGND.n2883 VGND.t1534 34.8005
R3616 VGND.n2883 VGND.t615 34.8005
R3617 VGND.n239 VGND.t170 34.8005
R3618 VGND.n239 VGND.t745 34.8005
R3619 VGND.n881 VGND.t1070 34.8005
R3620 VGND.n881 VGND.t198 34.8005
R3621 VGND.n883 VGND.t831 34.8005
R3622 VGND.n883 VGND.t2446 34.8005
R3623 VGND.n1422 VGND.t372 34.8005
R3624 VGND.n1422 VGND.t683 34.8005
R3625 VGND.n1427 VGND.t579 34.8005
R3626 VGND.n1427 VGND.t49 34.8005
R3627 VGND.n1432 VGND.t1544 34.8005
R3628 VGND.n1432 VGND.t196 34.8005
R3629 VGND.n1437 VGND.t1704 34.8005
R3630 VGND.n1437 VGND.t2442 34.8005
R3631 VGND.n1442 VGND.t299 34.8005
R3632 VGND.n1442 VGND.t2440 34.8005
R3633 VGND.n1447 VGND.t1668 34.8005
R3634 VGND.n1447 VGND.t194 34.8005
R3635 VGND.n1452 VGND.t332 34.8005
R3636 VGND.n1452 VGND.t192 34.8005
R3637 VGND.n789 VGND.t1840 34.8005
R3638 VGND.n789 VGND.t2444 34.8005
R3639 VGND.n1457 VGND.t454 34.8005
R3640 VGND.n1457 VGND.t202 34.8005
R3641 VGND.n1594 VGND.t708 34.8005
R3642 VGND.n1594 VGND.t200 34.8005
R3643 VGND.n1599 VGND.t1613 34.8005
R3644 VGND.n1599 VGND.t2438 34.8005
R3645 VGND.n748 VGND.t1259 34.8005
R3646 VGND.n748 VGND.t2436 34.8005
R3647 VGND.n1612 VGND.t27 34.8005
R3648 VGND.n1612 VGND.t685 34.8005
R3649 VGND.n1604 VGND.t2431 34.8005
R3650 VGND.n1604 VGND.t2448 34.8005
R3651 VGND.n1023 VGND.t1010 34.8005
R3652 VGND.n1023 VGND.t863 34.8005
R3653 VGND.n1030 VGND.t1163 34.8005
R3654 VGND.n1030 VGND.t274 34.8005
R3655 VGND.n1035 VGND.t594 34.8005
R3656 VGND.n1035 VGND.t1423 34.8005
R3657 VGND.n1027 VGND.t532 34.8005
R3658 VGND.n1027 VGND.t869 34.8005
R3659 VGND.n1093 VGND.t8 34.8005
R3660 VGND.n1093 VGND.t857 34.8005
R3661 VGND.n1088 VGND.t1312 34.8005
R3662 VGND.n1088 VGND.t270 34.8005
R3663 VGND.n1083 VGND.t433 34.8005
R3664 VGND.n1083 VGND.t268 34.8005
R3665 VGND.n1078 VGND.t545 34.8005
R3666 VGND.n1078 VGND.t855 34.8005
R3667 VGND.n1073 VGND.t18 34.8005
R3668 VGND.n1073 VGND.t853 34.8005
R3669 VGND.n1040 VGND.t1585 34.8005
R3670 VGND.n1040 VGND.t272 34.8005
R3671 VGND.n1042 VGND.t161 34.8005
R3672 VGND.n1042 VGND.t867 34.8005
R3673 VGND.n1051 VGND.t1123 34.8005
R3674 VGND.n1051 VGND.t865 34.8005
R3675 VGND.n1056 VGND.t1348 34.8005
R3676 VGND.n1056 VGND.t266 34.8005
R3677 VGND.n1047 VGND.t1998 34.8005
R3678 VGND.n1047 VGND.t1427 34.8005
R3679 VGND.n2903 VGND.t1380 34.8005
R3680 VGND.n2903 VGND.t1425 34.8005
R3681 VGND.n227 VGND.t178 34.8005
R3682 VGND.n227 VGND.t724 34.8005
R3683 VGND.n1013 VGND.t2614 34.8005
R3684 VGND.n1013 VGND.t2197 34.8005
R3685 VGND.n926 VGND.t2127 34.8005
R3686 VGND.n926 VGND.t2616 34.8005
R3687 VGND.n105 VGND.n103 34.6358
R3688 VGND.n2984 VGND.n2978 34.6358
R3689 VGND.n2987 VGND.n2986 34.6358
R3690 VGND.n2987 VGND.n2974 34.6358
R3691 VGND.n2991 VGND.n2974 34.6358
R3692 VGND.n2992 VGND.n2991 34.6358
R3693 VGND.n2993 VGND.n2992 34.6358
R3694 VGND.n21 VGND.n20 34.6358
R3695 VGND.n23 VGND.n12 34.6358
R3696 VGND.n27 VGND.n12 34.6358
R3697 VGND.n28 VGND.n27 34.6358
R3698 VGND.n29 VGND.n28 34.6358
R3699 VGND.n29 VGND.n9 34.6358
R3700 VGND.n3006 VGND.n10 34.6358
R3701 VGND.n181 VGND.n180 34.6358
R3702 VGND.n185 VGND.n184 34.6358
R3703 VGND.n2954 VGND.n2953 34.6358
R3704 VGND.n2956 VGND.n2947 34.6358
R3705 VGND.n2960 VGND.n2947 34.6358
R3706 VGND.n2961 VGND.n2960 34.6358
R3707 VGND.n2962 VGND.n2961 34.6358
R3708 VGND.n2962 VGND.n2945 34.6358
R3709 VGND.n47 VGND.n46 34.6358
R3710 VGND.n49 VGND.n38 34.6358
R3711 VGND.n53 VGND.n38 34.6358
R3712 VGND.n54 VGND.n53 34.6358
R3713 VGND.n55 VGND.n54 34.6358
R3714 VGND.n55 VGND.n35 34.6358
R3715 VGND.n109 VGND.n108 34.6358
R3716 VGND.n82 VGND.n81 34.6358
R3717 VGND.n86 VGND.n85 34.6358
R3718 VGND.n150 VGND.n149 34.6358
R3719 VGND.n154 VGND.n153 34.6358
R3720 VGND.n1153 VGND.n1135 34.6358
R3721 VGND.n1149 VGND.n1135 34.6358
R3722 VGND.n1149 VGND.n1148 34.6358
R3723 VGND.n1148 VGND.n1147 34.6358
R3724 VGND.n1147 VGND.n1137 34.6358
R3725 VGND.n1131 VGND.n1105 34.6358
R3726 VGND.n1126 VGND.n1106 34.6358
R3727 VGND.n1122 VGND.n1106 34.6358
R3728 VGND.n1122 VGND.n1121 34.6358
R3729 VGND.n1121 VGND.n1120 34.6358
R3730 VGND.n1120 VGND.n1108 34.6358
R3731 VGND.n486 VGND.n481 34.6358
R3732 VGND.n491 VGND.n490 34.6358
R3733 VGND.n2267 VGND.n2262 34.6358
R3734 VGND.n2272 VGND.n2271 34.6358
R3735 VGND.n522 VGND.n517 34.6358
R3736 VGND.n527 VGND.n526 34.6358
R3737 VGND.n2196 VGND.n2195 34.6358
R3738 VGND.n2204 VGND.n2203 34.6358
R3739 VGND.n2200 VGND.n2199 34.6358
R3740 VGND.n2243 VGND.n542 34.6358
R3741 VGND.n2243 VGND.n2242 34.6358
R3742 VGND.n2242 VGND.n2241 34.6358
R3743 VGND.n2241 VGND.n2227 34.6358
R3744 VGND.n2237 VGND.n2227 34.6358
R3745 VGND.n1361 VGND.n1356 34.6358
R3746 VGND.n1381 VGND.n1357 34.6358
R3747 VGND.n1381 VGND.n1380 34.6358
R3748 VGND.n1380 VGND.n1379 34.6358
R3749 VGND.n1379 VGND.n1365 34.6358
R3750 VGND.n1375 VGND.n1365 34.6358
R3751 VGND.n2998 VGND.n2997 34.6358
R3752 VGND.n2 VGND.t304 34.4422
R3753 VGND.n122 VGND.n121 33.1299
R3754 VGND.n2215 VGND.n544 33.1299
R3755 VGND.n111 VGND.n93 32.377
R3756 VGND.n187 VGND.n186 32.377
R3757 VGND.n111 VGND.n110 32.377
R3758 VGND.n88 VGND.n87 32.377
R3759 VGND.n156 VGND.n155 32.377
R3760 VGND.n2206 VGND.n2205 32.377
R3761 VGND.n2206 VGND.n2184 32.0005
R3762 VGND.n497 VGND.n494 30.4946
R3763 VGND.n2278 VGND.n2275 30.4946
R3764 VGND.n533 VGND.n530 30.4946
R3765 VGND.n190 VGND.n167 29.8709
R3766 VGND.n1143 VGND.n1142 28.9887
R3767 VGND.n1116 VGND.n1115 28.9887
R3768 VGND.n2235 VGND.n2234 28.9887
R3769 VGND.n1373 VGND.n1372 28.9887
R3770 VGND.n2985 VGND.n2984 27.8593
R3771 VGND.n22 VGND.n21 27.8593
R3772 VGND.n2955 VGND.n2954 27.8593
R3773 VGND.n48 VGND.n47 27.8593
R3774 VGND.n2256 VGND.n2255 27.0003
R3775 VGND.n161 VGND.n160 26.8591
R3776 VGND.n184 VGND.n173 26.3534
R3777 VGND.n108 VGND.n98 26.3534
R3778 VGND.n85 VGND.n74 26.3534
R3779 VGND.n153 VGND.n142 26.3534
R3780 VGND.n2203 VGND.n2188 26.3534
R3781 VGND.n129 VGND.n68 25.977
R3782 VGND.n498 VGND.n497 25.977
R3783 VGND.n2279 VGND.n2278 25.977
R3784 VGND.n534 VGND.n533 25.977
R3785 VGND.n509 VGND.n506 25.977
R3786 VGND.n2980 VGND.t2375 24.9236
R3787 VGND.n2980 VGND.t2327 24.9236
R3788 VGND.n2979 VGND.t2366 24.9236
R3789 VGND.n2979 VGND.t2310 24.9236
R3790 VGND.n2977 VGND.t2386 24.9236
R3791 VGND.n2977 VGND.t2359 24.9236
R3792 VGND.n2976 VGND.t2371 24.9236
R3793 VGND.n2976 VGND.t2343 24.9236
R3794 VGND.n17 VGND.t2358 24.9236
R3795 VGND.n17 VGND.t2390 24.9236
R3796 VGND.n16 VGND.t2314 24.9236
R3797 VGND.n16 VGND.t2353 24.9236
R3798 VGND.n15 VGND.t2364 24.9236
R3799 VGND.n15 VGND.t2334 24.9236
R3800 VGND.n14 VGND.t2324 24.9236
R3801 VGND.n14 VGND.t2382 24.9236
R3802 VGND.n176 VGND.t2304 24.9236
R3803 VGND.n176 VGND.t2345 24.9236
R3804 VGND.n175 VGND.t2362 24.9236
R3805 VGND.n175 VGND.t2302 24.9236
R3806 VGND.n172 VGND.t2312 24.9236
R3807 VGND.n172 VGND.t103 24.9236
R3808 VGND.n171 VGND.t2368 24.9236
R3809 VGND.n171 VGND.t360 24.9236
R3810 VGND.n170 VGND.t100 24.9236
R3811 VGND.n170 VGND.t106 24.9236
R3812 VGND.n169 VGND.t207 24.9236
R3813 VGND.n169 VGND.t2578 24.9236
R3814 VGND.n2950 VGND.t2379 24.9236
R3815 VGND.n2950 VGND.t2298 24.9236
R3816 VGND.n2949 VGND.t2308 24.9236
R3817 VGND.n2949 VGND.t2316 24.9236
R3818 VGND.n43 VGND.t2332 24.9236
R3819 VGND.n43 VGND.t2367 24.9236
R3820 VGND.n42 VGND.t2318 24.9236
R3821 VGND.n42 VGND.t2357 24.9236
R3822 VGND.n41 VGND.t2339 24.9236
R3823 VGND.n41 VGND.t2300 24.9236
R3824 VGND.n40 VGND.t2326 24.9236
R3825 VGND.n40 VGND.t2383 24.9236
R3826 VGND.n96 VGND.t2351 24.9236
R3827 VGND.n96 VGND.t2388 24.9236
R3828 VGND.n97 VGND.t2355 24.9236
R3829 VGND.n97 VGND.t1369 24.9236
R3830 VGND.n95 VGND.t1365 24.9236
R3831 VGND.n95 VGND.t1359 24.9236
R3832 VGND.n100 VGND.t2347 24.9236
R3833 VGND.n100 VGND.t2381 24.9236
R3834 VGND.n77 VGND.t2340 24.9236
R3835 VGND.n77 VGND.t2374 24.9236
R3836 VGND.n76 VGND.t2320 24.9236
R3837 VGND.n76 VGND.t2361 24.9236
R3838 VGND.n73 VGND.t2344 24.9236
R3839 VGND.n73 VGND.t937 24.9236
R3840 VGND.n72 VGND.t2329 24.9236
R3841 VGND.n72 VGND.t353 24.9236
R3842 VGND.n71 VGND.t936 24.9236
R3843 VGND.n71 VGND.t934 24.9236
R3844 VGND.n70 VGND.t349 24.9236
R3845 VGND.n70 VGND.t343 24.9236
R3846 VGND.n145 VGND.t2338 24.9236
R3847 VGND.n145 VGND.t2369 24.9236
R3848 VGND.n144 VGND.t2384 24.9236
R3849 VGND.n144 VGND.t2336 24.9236
R3850 VGND.n141 VGND.t2341 24.9236
R3851 VGND.n141 VGND.t2494 24.9236
R3852 VGND.n140 VGND.t2296 24.9236
R3853 VGND.n140 VGND.t859 24.9236
R3854 VGND.n139 VGND.t2679 24.9236
R3855 VGND.n139 VGND.t245 24.9236
R3856 VGND.n138 VGND.t1201 24.9236
R3857 VGND.n138 VGND.t277 24.9236
R3858 VGND.n1139 VGND.t1471 24.9236
R3859 VGND.n1139 VGND.t630 24.9236
R3860 VGND.n1141 VGND.t1479 24.9236
R3861 VGND.n1141 VGND.t1449 24.9236
R3862 VGND.n1111 VGND.t1207 24.9236
R3863 VGND.n1111 VGND.t1563 24.9236
R3864 VGND.n1110 VGND.t1472 24.9236
R3865 VGND.n1110 VGND.t633 24.9236
R3866 VGND.n1114 VGND.t1564 24.9236
R3867 VGND.n1114 VGND.t1483 24.9236
R3868 VGND.n1113 VGND.t1480 24.9236
R3869 VGND.n1113 VGND.t1450 24.9236
R3870 VGND.n488 VGND.t1205 24.9236
R3871 VGND.n488 VGND.t625 24.9236
R3872 VGND.n487 VGND.t47 24.9236
R3873 VGND.n487 VGND.t1464 24.9236
R3874 VGND.n478 VGND.t295 24.9236
R3875 VGND.n478 VGND.t1204 24.9236
R3876 VGND.n477 VGND.t2093 24.9236
R3877 VGND.n477 VGND.t46 24.9236
R3878 VGND.n496 VGND.t89 24.9236
R3879 VGND.n496 VGND.t294 24.9236
R3880 VGND.n495 VGND.t2095 24.9236
R3881 VGND.n495 VGND.t2094 24.9236
R3882 VGND.n2269 VGND.t1482 24.9236
R3883 VGND.n2269 VGND.t38 24.9236
R3884 VGND.n2268 VGND.t636 24.9236
R3885 VGND.n2268 VGND.t414 24.9236
R3886 VGND.n2259 VGND.t884 24.9236
R3887 VGND.n2259 VGND.t1477 24.9236
R3888 VGND.n2258 VGND.t1598 24.9236
R3889 VGND.n2258 VGND.t626 24.9236
R3890 VGND.n2277 VGND.t248 24.9236
R3891 VGND.n2277 VGND.t249 24.9236
R3892 VGND.n2276 VGND.t2075 24.9236
R3893 VGND.n2276 VGND.t1597 24.9236
R3894 VGND.n524 VGND.t1203 24.9236
R3895 VGND.n524 VGND.t1467 24.9236
R3896 VGND.n523 VGND.t41 24.9236
R3897 VGND.n523 VGND.t1566 24.9236
R3898 VGND.n514 VGND.t144 24.9236
R3899 VGND.n514 VGND.t1202 24.9236
R3900 VGND.n513 VGND.t1458 24.9236
R3901 VGND.n513 VGND.t36 24.9236
R3902 VGND.n532 VGND.t146 24.9236
R3903 VGND.n532 VGND.t145 24.9236
R3904 VGND.n531 VGND.t1460 24.9236
R3905 VGND.n531 VGND.t1459 24.9236
R3906 VGND.n2186 VGND.t628 24.9236
R3907 VGND.n2186 VGND.t409 24.9236
R3908 VGND.n2187 VGND.t1167 24.9236
R3909 VGND.n2187 VGND.t638 24.9236
R3910 VGND.n2185 VGND.t1171 24.9236
R3911 VGND.n2185 VGND.t1169 24.9236
R3912 VGND.n2190 VGND.t1476 24.9236
R3913 VGND.n2190 VGND.t1447 24.9236
R3914 VGND.n2230 VGND.t1473 24.9236
R3915 VGND.n2230 VGND.t634 24.9236
R3916 VGND.n2229 VGND.t1567 24.9236
R3917 VGND.n2229 VGND.t1465 24.9236
R3918 VGND.n2233 VGND.t1481 24.9236
R3919 VGND.n2233 VGND.t1451 24.9236
R3920 VGND.n2231 VGND.t631 24.9236
R3921 VGND.n2231 VGND.t411 24.9236
R3922 VGND.n1368 VGND.t313 24.9236
R3923 VGND.n1368 VGND.t314 24.9236
R3924 VGND.n1367 VGND.t412 24.9236
R3925 VGND.n1367 VGND.t415 24.9236
R3926 VGND.n1371 VGND.t407 24.9236
R3927 VGND.n1371 VGND.t1206 24.9236
R3928 VGND.n1369 VGND.t40 24.9236
R3929 VGND.n1369 VGND.t1565 24.9236
R3930 VGND.n187 VGND.n166 24.4711
R3931 VGND.n61 VGND.n36 24.4711
R3932 VGND.n123 VGND.n122 24.4711
R3933 VGND.n88 VGND.n67 24.4711
R3934 VGND.n129 VGND.n128 24.4711
R3935 VGND.n156 VGND.n135 24.4711
R3936 VGND.n498 VGND.n474 24.4711
R3937 VGND.n2279 VGND.n2253 24.4711
R3938 VGND.n534 VGND.n505 24.4711
R3939 VGND.n509 VGND.n508 24.4711
R3940 VGND.n2216 VGND.n2215 24.4711
R3941 VGND.n2223 VGND.n541 24.4711
R3942 VGND.n164 VGND.n136 23.7181
R3943 VGND.n2993 VGND.n2972 23.7181
R3944 VGND.n3010 VGND.n9 23.7181
R3945 VGND.n3010 VGND.n10 23.7181
R3946 VGND.n2966 VGND.n2945 23.7181
R3947 VGND.n65 VGND.n35 23.7181
R3948 VGND.n1155 VGND.n1153 23.7181
R3949 VGND.n1127 VGND.n1105 23.7181
R3950 VGND.n1127 VGND.n1126 23.7181
R3951 VGND.n2283 VGND.n2252 23.7181
R3952 VGND.n2210 VGND.n545 23.7181
R3953 VGND.n2247 VGND.n542 23.7181
R3954 VGND.n1385 VGND.n1356 23.7181
R3955 VGND.n1385 VGND.n1357 23.7181
R3956 VGND.n2997 VGND.n2972 23.7181
R3957 VGND.n117 VGND.n115 23.3417
R3958 VGND.n117 VGND.n92 23.3417
R3959 VGND.n2211 VGND.n2210 23.3417
R3960 VGND.n1143 VGND.n1140 21.4593
R3961 VGND.n1116 VGND.n1112 21.4593
R3962 VGND.n2236 VGND.n2235 21.4593
R3963 VGND.n1374 VGND.n1373 21.4593
R3964 VGND.n179 VGND.n178 21.0905
R3965 VGND.n102 VGND.n101 21.0905
R3966 VGND.n80 VGND.n79 21.0905
R3967 VGND.n148 VGND.n147 21.0905
R3968 VGND.n180 VGND.n179 20.3299
R3969 VGND.n103 VGND.n102 20.3299
R3970 VGND.n81 VGND.n80 20.3299
R3971 VGND.n149 VGND.n148 20.3299
R3972 VGND.n494 VGND.n479 19.9534
R3973 VGND.n2275 VGND.n2260 19.9534
R3974 VGND.n530 VGND.n515 19.9534
R3975 VGND.n3006 VGND.n3005 19.2005
R3976 VGND.n61 VGND.n60 19.2005
R3977 VGND.n2223 VGND.n2222 19.2005
R3978 VGND.n1361 VGND.n1360 19.2005
R3979 VGND.t2290 VGND.t1245 16.8587
R3980 VGND.t1590 VGND.t1247 16.8587
R3981 VGND.t254 VGND.t2079 16.8587
R3982 VGND.t1178 VGND.t2077 16.8587
R3983 VGND.n1133 VGND.n1132 16.077
R3984 VGND.n3000 VGND.n2999 16.077
R3985 VGND.n60 VGND.n59 15.4358
R3986 VGND.n2222 VGND.n2221 15.4358
R3987 VGND.n3005 VGND.n3004 14.6829
R3988 VGND.n160 VGND.n159 14.6829
R3989 VGND.n2255 VGND.n2254 14.6829
R3990 VGND.n1360 VGND.n1359 14.6829
R3991 VGND.n483 VGND.n482 14.5711
R3992 VGND.n2264 VGND.n2263 14.5711
R3993 VGND.n519 VGND.n518 14.5711
R3994 VGND.n2194 VGND.n2193 14.5711
R3995 VGND.n133 VGND.n68 14.3064
R3996 VGND.n538 VGND.n506 14.3064
R3997 VGND.n490 VGND.n489 13.9299
R3998 VGND.n2271 VGND.n2270 13.9299
R3999 VGND.n526 VGND.n525 13.9299
R4000 VGND.n2199 VGND.n2191 13.9299
R4001 VGND.n65 VGND.n36 13.5534
R4002 VGND.n2247 VGND.n541 13.5534
R4003 VGND.n193 VGND.n166 13.177
R4004 VGND.n133 VGND.n67 13.177
R4005 VGND.n164 VGND.n135 13.177
R4006 VGND.n502 VGND.n474 13.177
R4007 VGND.n2283 VGND.n2253 13.177
R4008 VGND.n538 VGND.n505 13.177
R4009 VGND.n193 VGND.n167 12.8005
R4010 VGND.n502 VGND.n475 12.8005
R4011 VGND.n3023 VGND.t2691 12.5645
R4012 VGND.n1132 VGND.n1131 10.5417
R4013 VGND.n2999 VGND.n2998 10.5417
R4014 VGND.n3004 VGND.n3003 10.0534
R4015 VGND.n1359 VGND.n1358 10.0534
R4016 VGND.n20 VGND.n19 9.3005
R4017 VGND.n21 VGND.n13 9.3005
R4018 VGND.n24 VGND.n23 9.3005
R4019 VGND.n25 VGND.n12 9.3005
R4020 VGND.n27 VGND.n26 9.3005
R4021 VGND.n28 VGND.n11 9.3005
R4022 VGND.n30 VGND.n29 9.3005
R4023 VGND.n31 VGND.n9 9.3005
R4024 VGND.n3008 VGND.n10 9.3005
R4025 VGND.n3007 VGND.n3006 9.3005
R4026 VGND.n3010 VGND.n3009 9.3005
R4027 VGND.n191 VGND.n167 9.3005
R4028 VGND.n180 VGND.n174 9.3005
R4029 VGND.n182 VGND.n181 9.3005
R4030 VGND.n184 VGND.n183 9.3005
R4031 VGND.n185 VGND.n168 9.3005
R4032 VGND.n188 VGND.n187 9.3005
R4033 VGND.n189 VGND.n166 9.3005
R4034 VGND.n193 VGND.n192 9.3005
R4035 VGND.n2953 VGND.n2952 9.3005
R4036 VGND.n2954 VGND.n2948 9.3005
R4037 VGND.n2957 VGND.n2956 9.3005
R4038 VGND.n2958 VGND.n2947 9.3005
R4039 VGND.n2960 VGND.n2959 9.3005
R4040 VGND.n2961 VGND.n2946 9.3005
R4041 VGND.n2963 VGND.n2962 9.3005
R4042 VGND.n2964 VGND.n2945 9.3005
R4043 VGND.n2966 VGND.n2965 9.3005
R4044 VGND.n59 VGND.n58 9.3005
R4045 VGND.n46 VGND.n45 9.3005
R4046 VGND.n47 VGND.n39 9.3005
R4047 VGND.n50 VGND.n49 9.3005
R4048 VGND.n51 VGND.n38 9.3005
R4049 VGND.n53 VGND.n52 9.3005
R4050 VGND.n54 VGND.n37 9.3005
R4051 VGND.n56 VGND.n55 9.3005
R4052 VGND.n57 VGND.n35 9.3005
R4053 VGND.n63 VGND.n36 9.3005
R4054 VGND.n62 VGND.n61 9.3005
R4055 VGND.n65 VGND.n64 9.3005
R4056 VGND.n124 VGND.n123 9.3005
R4057 VGND.n103 VGND.n99 9.3005
R4058 VGND.n106 VGND.n105 9.3005
R4059 VGND.n108 VGND.n107 9.3005
R4060 VGND.n109 VGND.n94 9.3005
R4061 VGND.n112 VGND.n111 9.3005
R4062 VGND.n114 VGND.n113 9.3005
R4063 VGND.n120 VGND.n119 9.3005
R4064 VGND.n122 VGND.n91 9.3005
R4065 VGND.n118 VGND.n117 9.3005
R4066 VGND.n128 VGND.n127 9.3005
R4067 VGND.n81 VGND.n75 9.3005
R4068 VGND.n83 VGND.n82 9.3005
R4069 VGND.n85 VGND.n84 9.3005
R4070 VGND.n86 VGND.n69 9.3005
R4071 VGND.n89 VGND.n88 9.3005
R4072 VGND.n90 VGND.n67 9.3005
R4073 VGND.n131 VGND.n68 9.3005
R4074 VGND.n130 VGND.n129 9.3005
R4075 VGND.n133 VGND.n132 9.3005
R4076 VGND.n162 VGND.n136 9.3005
R4077 VGND.n149 VGND.n143 9.3005
R4078 VGND.n151 VGND.n150 9.3005
R4079 VGND.n153 VGND.n152 9.3005
R4080 VGND.n154 VGND.n137 9.3005
R4081 VGND.n157 VGND.n156 9.3005
R4082 VGND.n158 VGND.n135 9.3005
R4083 VGND.n164 VGND.n163 9.3005
R4084 VGND.n1144 VGND.n1143 9.3005
R4085 VGND.n1145 VGND.n1137 9.3005
R4086 VGND.n1147 VGND.n1146 9.3005
R4087 VGND.n1148 VGND.n1136 9.3005
R4088 VGND.n1150 VGND.n1149 9.3005
R4089 VGND.n1151 VGND.n1135 9.3005
R4090 VGND.n1153 VGND.n1152 9.3005
R4091 VGND.n1156 VGND.n1155 9.3005
R4092 VGND.n1117 VGND.n1116 9.3005
R4093 VGND.n1118 VGND.n1108 9.3005
R4094 VGND.n1120 VGND.n1119 9.3005
R4095 VGND.n1121 VGND.n1107 9.3005
R4096 VGND.n1123 VGND.n1122 9.3005
R4097 VGND.n1124 VGND.n1106 9.3005
R4098 VGND.n1126 VGND.n1125 9.3005
R4099 VGND.n1129 VGND.n1105 9.3005
R4100 VGND.n1131 VGND.n1130 9.3005
R4101 VGND.n1128 VGND.n1127 9.3005
R4102 VGND.n500 VGND.n474 9.3005
R4103 VGND.n484 VGND.n481 9.3005
R4104 VGND.n486 VGND.n485 9.3005
R4105 VGND.n490 VGND.n480 9.3005
R4106 VGND.n492 VGND.n491 9.3005
R4107 VGND.n494 VGND.n493 9.3005
R4108 VGND.n497 VGND.n476 9.3005
R4109 VGND.n499 VGND.n498 9.3005
R4110 VGND.n502 VGND.n501 9.3005
R4111 VGND.n2281 VGND.n2253 9.3005
R4112 VGND.n2265 VGND.n2262 9.3005
R4113 VGND.n2267 VGND.n2266 9.3005
R4114 VGND.n2271 VGND.n2261 9.3005
R4115 VGND.n2273 VGND.n2272 9.3005
R4116 VGND.n2275 VGND.n2274 9.3005
R4117 VGND.n2278 VGND.n2257 9.3005
R4118 VGND.n2280 VGND.n2279 9.3005
R4119 VGND.n2256 VGND.n2252 9.3005
R4120 VGND.n2283 VGND.n2282 9.3005
R4121 VGND.n508 VGND.n507 9.3005
R4122 VGND.n511 VGND.n506 9.3005
R4123 VGND.n536 VGND.n505 9.3005
R4124 VGND.n520 VGND.n517 9.3005
R4125 VGND.n522 VGND.n521 9.3005
R4126 VGND.n526 VGND.n516 9.3005
R4127 VGND.n528 VGND.n527 9.3005
R4128 VGND.n530 VGND.n529 9.3005
R4129 VGND.n533 VGND.n512 9.3005
R4130 VGND.n535 VGND.n534 9.3005
R4131 VGND.n510 VGND.n509 9.3005
R4132 VGND.n538 VGND.n537 9.3005
R4133 VGND.n2217 VGND.n2216 9.3005
R4134 VGND.n2208 VGND.n545 9.3005
R4135 VGND.n2195 VGND.n2192 9.3005
R4136 VGND.n2197 VGND.n2196 9.3005
R4137 VGND.n2199 VGND.n2198 9.3005
R4138 VGND.n2201 VGND.n2200 9.3005
R4139 VGND.n2203 VGND.n2202 9.3005
R4140 VGND.n2204 VGND.n2183 9.3005
R4141 VGND.n2207 VGND.n2206 9.3005
R4142 VGND.n2213 VGND.n2212 9.3005
R4143 VGND.n2215 VGND.n2214 9.3005
R4144 VGND.n2210 VGND.n2209 9.3005
R4145 VGND.n2235 VGND.n2228 9.3005
R4146 VGND.n2238 VGND.n2237 9.3005
R4147 VGND.n2239 VGND.n2227 9.3005
R4148 VGND.n2241 VGND.n2240 9.3005
R4149 VGND.n2242 VGND.n2226 9.3005
R4150 VGND.n2244 VGND.n2243 9.3005
R4151 VGND.n2245 VGND.n542 9.3005
R4152 VGND.n2225 VGND.n541 9.3005
R4153 VGND.n2224 VGND.n2223 9.3005
R4154 VGND.n2221 VGND.n2220 9.3005
R4155 VGND.n2247 VGND.n2246 9.3005
R4156 VGND.n1373 VGND.n1366 9.3005
R4157 VGND.n1376 VGND.n1375 9.3005
R4158 VGND.n1377 VGND.n1365 9.3005
R4159 VGND.n1379 VGND.n1378 9.3005
R4160 VGND.n1380 VGND.n1364 9.3005
R4161 VGND.n1382 VGND.n1381 9.3005
R4162 VGND.n1383 VGND.n1357 9.3005
R4163 VGND.n1363 VGND.n1356 9.3005
R4164 VGND.n1362 VGND.n1361 9.3005
R4165 VGND.n1385 VGND.n1384 9.3005
R4166 VGND.n2982 VGND.n2978 9.3005
R4167 VGND.n2984 VGND.n2983 9.3005
R4168 VGND.n2986 VGND.n2975 9.3005
R4169 VGND.n2988 VGND.n2987 9.3005
R4170 VGND.n2989 VGND.n2974 9.3005
R4171 VGND.n2991 VGND.n2990 9.3005
R4172 VGND.n2992 VGND.n2973 9.3005
R4173 VGND.n2994 VGND.n2993 9.3005
R4174 VGND.n2995 VGND.n2972 9.3005
R4175 VGND.n2997 VGND.n2996 9.3005
R4176 VGND.n2998 VGND.n34 9.3005
R4177 VGND.n181 VGND.n173 8.28285
R4178 VGND.n82 VGND.n74 8.28285
R4179 VGND.n150 VGND.n142 8.28285
R4180 VGND.n2636 VGND.n2635 7.9105
R4181 VGND.n2693 VGND.n337 7.9105
R4182 VGND.n2692 VGND.n338 7.9105
R4183 VGND.n2687 VGND.n343 7.9105
R4184 VGND.n2686 VGND.n344 7.9105
R4185 VGND.n2681 VGND.n349 7.9105
R4186 VGND.n2680 VGND.n350 7.9105
R4187 VGND.n2675 VGND.n2674 7.9105
R4188 VGND.n2712 VGND.n2711 7.9105
R4189 VGND.n2721 VGND.n2720 7.9105
R4190 VGND.n2745 VGND.n2744 7.9105
R4191 VGND.n2759 VGND.n2758 7.9105
R4192 VGND.n2783 VGND.n288 7.9105
R4193 VGND.n2785 VGND.n2784 7.9105
R4194 VGND.n2794 VGND.n2793 7.9105
R4195 VGND.n2937 VGND.n2936 7.9105
R4196 VGND.n2559 VGND.n401 7.9105
R4197 VGND.n2558 VGND.n402 7.9105
R4198 VGND.n2557 VGND.n403 7.9105
R4199 VGND.n2556 VGND.n404 7.9105
R4200 VGND.n2555 VGND.n405 7.9105
R4201 VGND.n2554 VGND.n406 7.9105
R4202 VGND.n2553 VGND.n407 7.9105
R4203 VGND.n2552 VGND.n408 7.9105
R4204 VGND.n2551 VGND.n409 7.9105
R4205 VGND.n2550 VGND.n410 7.9105
R4206 VGND.n2549 VGND.n411 7.9105
R4207 VGND.n2548 VGND.n412 7.9105
R4208 VGND.n2547 VGND.n2546 7.9105
R4209 VGND.n2798 VGND.n282 7.9105
R4210 VGND.n2797 VGND.n283 7.9105
R4211 VGND.n2534 VGND.n2533 7.9105
R4212 VGND.n2357 VGND.n2356 7.9105
R4213 VGND.n2374 VGND.n2373 7.9105
R4214 VGND.n2383 VGND.n2382 7.9105
R4215 VGND.n2400 VGND.n2399 7.9105
R4216 VGND.n2409 VGND.n2408 7.9105
R4217 VGND.n2426 VGND.n2425 7.9105
R4218 VGND.n2435 VGND.n2434 7.9105
R4219 VGND.n2452 VGND.n2451 7.9105
R4220 VGND.n2461 VGND.n2460 7.9105
R4221 VGND.n2478 VGND.n2477 7.9105
R4222 VGND.n2487 VGND.n2486 7.9105
R4223 VGND.n2509 VGND.n2508 7.9105
R4224 VGND.n2802 VGND.n279 7.9105
R4225 VGND.n2801 VGND.n280 7.9105
R4226 VGND.n420 VGND.n419 7.9105
R4227 VGND.n2530 VGND.n2529 7.9105
R4228 VGND.n2361 VGND.n2360 7.9105
R4229 VGND.n2370 VGND.n2369 7.9105
R4230 VGND.n2387 VGND.n2386 7.9105
R4231 VGND.n2396 VGND.n2395 7.9105
R4232 VGND.n2413 VGND.n2412 7.9105
R4233 VGND.n2422 VGND.n2421 7.9105
R4234 VGND.n2439 VGND.n2438 7.9105
R4235 VGND.n2448 VGND.n2447 7.9105
R4236 VGND.n2465 VGND.n2464 7.9105
R4237 VGND.n2474 VGND.n2473 7.9105
R4238 VGND.n2491 VGND.n2490 7.9105
R4239 VGND.n2505 VGND.n2504 7.9105
R4240 VGND.n2805 VGND.n277 7.9105
R4241 VGND.n2807 VGND.n2806 7.9105
R4242 VGND.n2819 VGND.n273 7.9105
R4243 VGND.n2818 VGND.n2817 7.9105
R4244 VGND.n1908 VGND.n1907 7.9105
R4245 VGND.n1917 VGND.n1916 7.9105
R4246 VGND.n1919 VGND.n1918 7.9105
R4247 VGND.n1928 VGND.n1927 7.9105
R4248 VGND.n1930 VGND.n1929 7.9105
R4249 VGND.n1939 VGND.n1938 7.9105
R4250 VGND.n1941 VGND.n1940 7.9105
R4251 VGND.n1950 VGND.n1949 7.9105
R4252 VGND.n1952 VGND.n1951 7.9105
R4253 VGND.n1961 VGND.n1960 7.9105
R4254 VGND.n1963 VGND.n1962 7.9105
R4255 VGND.n1972 VGND.n1971 7.9105
R4256 VGND.n1974 VGND.n1973 7.9105
R4257 VGND.n2823 VGND.n270 7.9105
R4258 VGND.n2822 VGND.n271 7.9105
R4259 VGND.n1990 VGND.n1989 7.9105
R4260 VGND.n2063 VGND.n591 7.9105
R4261 VGND.n2062 VGND.n2061 7.9105
R4262 VGND.n2167 VGND.n556 7.9105
R4263 VGND.n2166 VGND.n557 7.9105
R4264 VGND.n2159 VGND.n562 7.9105
R4265 VGND.n2158 VGND.n563 7.9105
R4266 VGND.n2151 VGND.n568 7.9105
R4267 VGND.n2150 VGND.n569 7.9105
R4268 VGND.n2143 VGND.n574 7.9105
R4269 VGND.n2142 VGND.n575 7.9105
R4270 VGND.n2135 VGND.n580 7.9105
R4271 VGND.n2134 VGND.n581 7.9105
R4272 VGND.n2827 VGND.n267 7.9105
R4273 VGND.n2826 VGND.n268 7.9105
R4274 VGND.n1999 VGND.n1998 7.9105
R4275 VGND.n1997 VGND.n1996 7.9105
R4276 VGND.n2067 VGND.n2066 7.9105
R4277 VGND.n2171 VGND.n553 7.9105
R4278 VGND.n2170 VGND.n554 7.9105
R4279 VGND.n2163 VGND.n559 7.9105
R4280 VGND.n2162 VGND.n560 7.9105
R4281 VGND.n2155 VGND.n565 7.9105
R4282 VGND.n2154 VGND.n566 7.9105
R4283 VGND.n2147 VGND.n571 7.9105
R4284 VGND.n2146 VGND.n572 7.9105
R4285 VGND.n2139 VGND.n577 7.9105
R4286 VGND.n2138 VGND.n578 7.9105
R4287 VGND.n2131 VGND.n2130 7.9105
R4288 VGND.n2830 VGND.n265 7.9105
R4289 VGND.n2832 VGND.n2831 7.9105
R4290 VGND.n2844 VGND.n261 7.9105
R4291 VGND.n2843 VGND.n2842 7.9105
R4292 VGND.n1901 VGND.n548 7.9105
R4293 VGND.n2175 VGND.n2174 7.9105
R4294 VGND.n1759 VGND.n1758 7.9105
R4295 VGND.n1768 VGND.n1767 7.9105
R4296 VGND.n1770 VGND.n1769 7.9105
R4297 VGND.n1779 VGND.n1778 7.9105
R4298 VGND.n1781 VGND.n1780 7.9105
R4299 VGND.n1790 VGND.n1789 7.9105
R4300 VGND.n1792 VGND.n1791 7.9105
R4301 VGND.n1801 VGND.n1800 7.9105
R4302 VGND.n1803 VGND.n1802 7.9105
R4303 VGND.n1812 VGND.n1811 7.9105
R4304 VGND.n1814 VGND.n1813 7.9105
R4305 VGND.n2848 VGND.n258 7.9105
R4306 VGND.n2847 VGND.n259 7.9105
R4307 VGND.n1830 VGND.n1829 7.9105
R4308 VGND.n1899 VGND.n629 7.9105
R4309 VGND.n1685 VGND.n1684 7.9105
R4310 VGND.n1687 VGND.n1686 7.9105
R4311 VGND.n1884 VGND.n643 7.9105
R4312 VGND.n1883 VGND.n644 7.9105
R4313 VGND.n1876 VGND.n649 7.9105
R4314 VGND.n1875 VGND.n650 7.9105
R4315 VGND.n1868 VGND.n655 7.9105
R4316 VGND.n1867 VGND.n656 7.9105
R4317 VGND.n1860 VGND.n661 7.9105
R4318 VGND.n1859 VGND.n662 7.9105
R4319 VGND.n1852 VGND.n1851 7.9105
R4320 VGND.n2852 VGND.n255 7.9105
R4321 VGND.n2851 VGND.n256 7.9105
R4322 VGND.n1839 VGND.n1838 7.9105
R4323 VGND.n1837 VGND.n1836 7.9105
R4324 VGND.n1896 VGND.n633 7.9105
R4325 VGND.n1895 VGND.n634 7.9105
R4326 VGND.n1888 VGND.n640 7.9105
R4327 VGND.n1887 VGND.n641 7.9105
R4328 VGND.n1880 VGND.n646 7.9105
R4329 VGND.n1879 VGND.n647 7.9105
R4330 VGND.n1872 VGND.n652 7.9105
R4331 VGND.n1871 VGND.n653 7.9105
R4332 VGND.n1864 VGND.n658 7.9105
R4333 VGND.n1863 VGND.n659 7.9105
R4334 VGND.n1856 VGND.n664 7.9105
R4335 VGND.n1855 VGND.n730 7.9105
R4336 VGND.n2855 VGND.n253 7.9105
R4337 VGND.n2857 VGND.n2856 7.9105
R4338 VGND.n2869 VGND.n249 7.9105
R4339 VGND.n2868 VGND.n2867 7.9105
R4340 VGND.n1350 VGND.n1349 7.9105
R4341 VGND.n1892 VGND.n636 7.9105
R4342 VGND.n1891 VGND.n637 7.9105
R4343 VGND.n868 VGND.n867 7.9105
R4344 VGND.n866 VGND.n812 7.9105
R4345 VGND.n865 VGND.n813 7.9105
R4346 VGND.n864 VGND.n814 7.9105
R4347 VGND.n863 VGND.n815 7.9105
R4348 VGND.n862 VGND.n816 7.9105
R4349 VGND.n861 VGND.n817 7.9105
R4350 VGND.n860 VGND.n859 7.9105
R4351 VGND.n1669 VGND.n732 7.9105
R4352 VGND.n1668 VGND.n1667 7.9105
R4353 VGND.n2873 VGND.n246 7.9105
R4354 VGND.n2872 VGND.n247 7.9105
R4355 VGND.n1655 VGND.n1654 7.9105
R4356 VGND.n1404 VGND.n801 7.9105
R4357 VGND.n1403 VGND.n802 7.9105
R4358 VGND.n1402 VGND.n1401 7.9105
R4359 VGND.n1488 VGND.n1487 7.9105
R4360 VGND.n1497 VGND.n1496 7.9105
R4361 VGND.n1514 VGND.n1513 7.9105
R4362 VGND.n1523 VGND.n1522 7.9105
R4363 VGND.n1540 VGND.n1539 7.9105
R4364 VGND.n1560 VGND.n758 7.9105
R4365 VGND.n1559 VGND.n1558 7.9105
R4366 VGND.n1628 VGND.n742 7.9105
R4367 VGND.n1630 VGND.n1629 7.9105
R4368 VGND.n2877 VGND.n243 7.9105
R4369 VGND.n2876 VGND.n244 7.9105
R4370 VGND.n741 VGND.n740 7.9105
R4371 VGND.n1651 VGND.n1650 7.9105
R4372 VGND.n1408 VGND.n1407 7.9105
R4373 VGND.n1417 VGND.n1416 7.9105
R4374 VGND.n1475 VGND.n1474 7.9105
R4375 VGND.n1484 VGND.n1483 7.9105
R4376 VGND.n1501 VGND.n1500 7.9105
R4377 VGND.n1510 VGND.n1509 7.9105
R4378 VGND.n1527 VGND.n1526 7.9105
R4379 VGND.n1536 VGND.n1535 7.9105
R4380 VGND.n1564 VGND.n1563 7.9105
R4381 VGND.n1588 VGND.n1587 7.9105
R4382 VGND.n1625 VGND.n744 7.9105
R4383 VGND.n1624 VGND.n745 7.9105
R4384 VGND.n2880 VGND.n240 7.9105
R4385 VGND.n2882 VGND.n2881 7.9105
R4386 VGND.n2894 VGND.n236 7.9105
R4387 VGND.n2893 VGND.n2892 7.9105
R4388 VGND.n1344 VGND.n1343 7.9105
R4389 VGND.n1421 VGND.n1420 7.9105
R4390 VGND.n1471 VGND.n783 7.9105
R4391 VGND.n1470 VGND.n784 7.9105
R4392 VGND.n1469 VGND.n785 7.9105
R4393 VGND.n1468 VGND.n786 7.9105
R4394 VGND.n1467 VGND.n787 7.9105
R4395 VGND.n1466 VGND.n788 7.9105
R4396 VGND.n1465 VGND.n1464 7.9105
R4397 VGND.n1591 VGND.n751 7.9105
R4398 VGND.n1593 VGND.n1592 7.9105
R4399 VGND.n1621 VGND.n747 7.9105
R4400 VGND.n1620 VGND.n1619 7.9105
R4401 VGND.n2898 VGND.n231 7.9105
R4402 VGND.n2897 VGND.n232 7.9105
R4403 VGND.n1607 VGND.n1606 7.9105
R4404 VGND.n1103 VGND.n1025 7.9105
R4405 VGND.n1102 VGND.n1026 7.9105
R4406 VGND.n1101 VGND.n1100 7.9105
R4407 VGND.n1321 VGND.n899 7.9105
R4408 VGND.n1320 VGND.n900 7.9105
R4409 VGND.n1313 VGND.n905 7.9105
R4410 VGND.n1312 VGND.n906 7.9105
R4411 VGND.n1305 VGND.n911 7.9105
R4412 VGND.n1304 VGND.n912 7.9105
R4413 VGND.n1068 VGND.n1067 7.9105
R4414 VGND.n1066 VGND.n1045 7.9105
R4415 VGND.n1065 VGND.n1046 7.9105
R4416 VGND.n1064 VGND.n1063 7.9105
R4417 VGND.n2902 VGND.n2901 7.9105
R4418 VGND.n233 VGND.n228 7.9105
R4419 VGND.n2913 VGND.n2912 7.9105
R4420 VGND.n1161 VGND.n888 7.9105
R4421 VGND.n1331 VGND.n1330 7.9105
R4422 VGND.n1325 VGND.n896 7.9105
R4423 VGND.n1324 VGND.n897 7.9105
R4424 VGND.n1317 VGND.n902 7.9105
R4425 VGND.n1316 VGND.n903 7.9105
R4426 VGND.n1309 VGND.n908 7.9105
R4427 VGND.n1308 VGND.n909 7.9105
R4428 VGND.n1301 VGND.n914 7.9105
R4429 VGND.n1300 VGND.n915 7.9105
R4430 VGND.n1295 VGND.n919 7.9105
R4431 VGND.n1294 VGND.n920 7.9105
R4432 VGND.n1289 VGND.n924 7.9105
R4433 VGND.n1288 VGND.n925 7.9105
R4434 VGND.n1287 VGND.n992 7.9105
R4435 VGND.n2917 VGND.n2916 7.9105
R4436 VGND.n489 VGND.n486 7.90638
R4437 VGND.n482 VGND.n481 7.90638
R4438 VGND.n2270 VGND.n2267 7.90638
R4439 VGND.n2263 VGND.n2262 7.90638
R4440 VGND.n525 VGND.n522 7.90638
R4441 VGND.n518 VGND.n517 7.90638
R4442 VGND.n2196 VGND.n2191 7.90638
R4443 VGND.n2195 VGND.n2194 7.90638
R4444 VGND.n1142 VGND.n1138 7.4049
R4445 VGND.n1115 VGND.n1109 7.4049
R4446 VGND.n2234 VGND.n2232 7.4049
R4447 VGND.n1372 VGND.n1370 7.4049
R4448 VGND VGND.n475 7.12482
R4449 VGND.n178 VGND.n177 6.85473
R4450 VGND.n79 VGND.n78 6.85473
R4451 VGND.n147 VGND.n146 6.85473
R4452 VGND.n2986 VGND.n2985 6.77697
R4453 VGND.n23 VGND.n22 6.77697
R4454 VGND.n2956 VGND.n2955 6.77697
R4455 VGND.n49 VGND.n48 6.77697
R4456 VGND.n3022 VGND.n3021 6.4005
R4457 VGND.n104 VGND.n98 5.27109
R4458 VGND.n2189 VGND.n2188 5.27109
R4459 VGND.n2565 VGND.n2564 4.5005
R4460 VGND.n2568 VGND.n2567 4.5005
R4461 VGND.n2571 VGND.n2570 4.5005
R4462 VGND.n2574 VGND.n2573 4.5005
R4463 VGND.n2577 VGND.n2576 4.5005
R4464 VGND.n2580 VGND.n2579 4.5005
R4465 VGND.n2583 VGND.n2582 4.5005
R4466 VGND.n2586 VGND.n2585 4.5005
R4467 VGND.n2589 VGND.n2588 4.5005
R4468 VGND.n2592 VGND.n2591 4.5005
R4469 VGND.n2595 VGND.n2594 4.5005
R4470 VGND.n2598 VGND.n2597 4.5005
R4471 VGND.n2601 VGND.n2600 4.5005
R4472 VGND.n2604 VGND.n2603 4.5005
R4473 VGND.n2607 VGND.n2606 4.5005
R4474 VGND.n335 VGND.n334 4.5005
R4475 VGND.n2627 VGND.n2626 4.5005
R4476 VGND.n2624 VGND.n2623 4.5005
R4477 VGND.n2621 VGND.n2620 4.5005
R4478 VGND.n2618 VGND.n2617 4.5005
R4479 VGND.n2615 VGND.n2614 4.5005
R4480 VGND.n2612 VGND.n2611 4.5005
R4481 VGND.n323 VGND.n322 4.5005
R4482 VGND.n316 VGND.n315 4.5005
R4483 VGND.n307 VGND.n306 4.5005
R4484 VGND.n2763 VGND.n299 4.5005
R4485 VGND.n2766 VGND.n2765 4.5005
R4486 VGND.n291 VGND.n290 4.5005
R4487 VGND.n2770 VGND.n297 4.5005
R4488 VGND.n205 VGND.n204 4.5005
R4489 VGND.n2631 VGND.n2630 4.5005
R4490 VGND.n2632 VGND.n331 4.5005
R4491 VGND.n2697 VGND.n2696 4.5005
R4492 VGND.n358 VGND.n340 4.5005
R4493 VGND.n365 VGND.n341 4.5005
R4494 VGND.n354 VGND.n346 4.5005
R4495 VGND.n376 VGND.n347 4.5005
R4496 VGND.n353 VGND.n352 4.5005
R4497 VGND.n390 VGND.n389 4.5005
R4498 VGND.n2708 VGND.n2707 4.5005
R4499 VGND.n2725 VGND.n2724 4.5005
R4500 VGND.n2741 VGND.n2740 4.5005
R4501 VGND.n2762 VGND.n300 4.5005
R4502 VGND.n2733 VGND.n289 4.5005
R4503 VGND.n2779 VGND.n2778 4.5005
R4504 VGND.n2772 VGND.n2771 4.5005
R4505 VGND.n2942 VGND.n2941 4.5005
R4506 VGND.n1019 VGND.n1018 4.5005
R4507 VGND.n1016 VGND.n1015 4.5005
R4508 VGND.n1181 VGND.n1180 4.5005
R4509 VGND.n1193 VGND.n1006 4.5005
R4510 VGND.n1200 VGND.n1004 4.5005
R4511 VGND.n1197 VGND.n1195 4.5005
R4512 VGND.n1213 VGND.n1212 4.5005
R4513 VGND.n1251 VGND.n1000 4.5005
R4514 VGND.n1254 VGND.n1253 4.5005
R4515 VGND.n1257 VGND.n1256 4.5005
R4516 VGND.n1260 VGND.n1259 4.5005
R4517 VGND.n1263 VGND.n1262 4.5005
R4518 VGND.n1269 VGND.n998 4.5005
R4519 VGND.n1266 VGND.n1265 4.5005
R4520 VGND.n995 VGND.n994 4.5005
R4521 VGND.n1022 VGND.n1021 4.5005
R4522 VGND.n1165 VGND.n1164 4.5005
R4523 VGND.n1170 VGND.n891 4.5005
R4524 VGND.n1011 VGND.n892 4.5005
R4525 VGND.n1183 VGND.n1182 4.5005
R4526 VGND.n1192 VGND.n1191 4.5005
R4527 VGND.n1202 VGND.n1201 4.5005
R4528 VGND.n1196 VGND.n1003 4.5005
R4529 VGND.n1215 VGND.n1214 4.5005
R4530 VGND.n1250 VGND.n1249 4.5005
R4531 VGND.n1223 VGND.n916 4.5005
R4532 VGND.n1242 VGND.n917 4.5005
R4533 VGND.n1228 VGND.n921 4.5005
R4534 VGND.n1235 VGND.n922 4.5005
R4535 VGND.n1272 VGND.n1271 4.5005
R4536 VGND.n997 VGND.n993 4.5005
R4537 VGND.n1283 VGND.n1282 4.5005
R4538 VGND.n1157 VGND.n1156 4.41365
R4539 VGND VGND.n33 4.35375
R4540 VGND.n1134 VGND.n1133 4.05427
R4541 VGND.n507 VGND.n0 4.05427
R4542 VGND.n2218 VGND.n2217 4.05427
R4543 VGND.n2220 VGND.n2219 4.05427
R4544 VGND.n1358 VGND.n543 4.05427
R4545 VGND VGND.n3002 3.99438
R4546 VGND VGND.n32 3.99438
R4547 VGND.n125 VGND 3.99438
R4548 VGND VGND.n126 3.99438
R4549 VGND.n3001 VGND 3.99437
R4550 VGND.n1284 VGND.n223 3.77268
R4551 VGND.n2940 VGND.n206 3.77268
R4552 VGND.n1163 VGND.n1162 3.77268
R4553 VGND.n2634 VGND.n2633 3.77268
R4554 VGND.n1327 VGND.n1326 3.77268
R4555 VGND.n2691 VGND.n2690 3.77268
R4556 VGND.n1323 VGND.n898 3.77268
R4557 VGND.n2689 VGND.n2688 3.77268
R4558 VGND.n1318 VGND.n901 3.77268
R4559 VGND.n2685 VGND.n2684 3.77268
R4560 VGND.n1315 VGND.n904 3.77268
R4561 VGND.n2683 VGND.n2682 3.77268
R4562 VGND.n1310 VGND.n907 3.77268
R4563 VGND.n2679 VGND.n2678 3.77268
R4564 VGND.n1307 VGND.n910 3.77268
R4565 VGND.n2677 VGND.n2676 3.77268
R4566 VGND.n1302 VGND.n913 3.77268
R4567 VGND.n2710 VGND.n2709 3.77268
R4568 VGND.n1299 VGND.n1298 3.77268
R4569 VGND.n2723 VGND.n2722 3.77268
R4570 VGND.n1297 VGND.n1296 3.77268
R4571 VGND.n2743 VGND.n2742 3.77268
R4572 VGND.n1293 VGND.n1292 3.77268
R4573 VGND.n2761 VGND.n2760 3.77268
R4574 VGND.n1291 VGND.n1290 3.77268
R4575 VGND.n2782 VGND.n2781 3.77268
R4576 VGND.n1270 VGND.n229 3.77268
R4577 VGND.n2780 VGND.n281 3.77268
R4578 VGND.n1286 VGND.n1285 3.77268
R4579 VGND.n2795 VGND.n284 3.77268
R4580 VGND.n1329 VGND.n1328 3.77268
R4581 VGND.n2695 VGND.n2694 3.77268
R4582 VGND.n2769 VGND.n205 3.75914
R4583 VGND.n2631 VGND.n2629 3.75914
R4584 VGND.n1267 VGND.n995 3.75914
R4585 VGND.n1022 VGND.n1020 3.75914
R4586 VGND.n2771 VGND.n284 3.4105
R4587 VGND.n2780 VGND.n2779 3.4105
R4588 VGND.n2781 VGND.n289 3.4105
R4589 VGND.n2762 VGND.n2761 3.4105
R4590 VGND.n2742 VGND.n2741 3.4105
R4591 VGND.n2724 VGND.n2723 3.4105
R4592 VGND.n2709 VGND.n2708 3.4105
R4593 VGND.n2677 VGND.n390 3.4105
R4594 VGND.n2678 VGND.n352 3.4105
R4595 VGND.n2683 VGND.n347 3.4105
R4596 VGND.n2684 VGND.n346 3.4105
R4597 VGND.n2689 VGND.n341 3.4105
R4598 VGND.n2690 VGND.n340 3.4105
R4599 VGND.n2696 VGND.n2695 3.4105
R4600 VGND.n2941 VGND.n2940 3.4105
R4601 VGND.n2770 VGND.n2769 3.4105
R4602 VGND.n2768 VGND.n291 3.4105
R4603 VGND.n2767 VGND.n2766 3.4105
R4604 VGND.n2764 VGND.n2763 3.4105
R4605 VGND.n307 VGND.n298 3.4105
R4606 VGND.n2609 VGND.n316 3.4105
R4607 VGND.n2610 VGND.n323 3.4105
R4608 VGND.n2613 VGND.n2612 3.4105
R4609 VGND.n2616 VGND.n2615 3.4105
R4610 VGND.n2619 VGND.n2618 3.4105
R4611 VGND.n2622 VGND.n2621 3.4105
R4612 VGND.n2625 VGND.n2624 3.4105
R4613 VGND.n2628 VGND.n2627 3.4105
R4614 VGND.n2629 VGND.n335 3.4105
R4615 VGND.n2633 VGND.n2632 3.4105
R4616 VGND.n2937 VGND.n206 3.4105
R4617 VGND.n2635 VGND.n2634 3.4105
R4618 VGND.n2559 VGND.n397 3.4105
R4619 VGND.n2533 VGND.n2532 3.4105
R4620 VGND.n2557 VGND.n339 3.4105
R4621 VGND.n2692 VGND.n2691 3.4105
R4622 VGND.n2384 VGND.n2383 3.4105
R4623 VGND.n2358 VGND.n2357 3.4105
R4624 VGND.n2531 VGND.n2530 3.4105
R4625 VGND.n2399 VGND.n2398 3.4105
R4626 VGND.n2556 VGND.n342 3.4105
R4627 VGND.n2688 VGND.n2687 3.4105
R4628 VGND.n2397 VGND.n2396 3.4105
R4629 VGND.n2386 VGND.n2385 3.4105
R4630 VGND.n2360 VGND.n2359 3.4105
R4631 VGND.n2818 VGND.n274 3.4105
R4632 VGND.n2412 VGND.n2411 3.4105
R4633 VGND.n2410 VGND.n2409 3.4105
R4634 VGND.n2555 VGND.n345 3.4105
R4635 VGND.n2686 VGND.n2685 3.4105
R4636 VGND.n1929 VGND.n449 3.4105
R4637 VGND.n1928 VGND.n453 3.4105
R4638 VGND.n1918 VGND.n457 3.4105
R4639 VGND.n1907 VGND.n467 3.4105
R4640 VGND.n1990 VGND.n604 3.4105
R4641 VGND.n1939 VGND.n445 3.4105
R4642 VGND.n2423 VGND.n2422 3.4105
R4643 VGND.n2425 VGND.n2424 3.4105
R4644 VGND.n2554 VGND.n348 3.4105
R4645 VGND.n2682 VGND.n2681 3.4105
R4646 VGND.n2158 VGND.n2157 3.4105
R4647 VGND.n2160 VGND.n2159 3.4105
R4648 VGND.n2166 VGND.n2165 3.4105
R4649 VGND.n2168 VGND.n2167 3.4105
R4650 VGND.n2064 VGND.n2063 3.4105
R4651 VGND.n1997 VGND.n603 3.4105
R4652 VGND.n2152 VGND.n2151 3.4105
R4653 VGND.n1940 VGND.n441 3.4105
R4654 VGND.n2438 VGND.n2437 3.4105
R4655 VGND.n2436 VGND.n2435 3.4105
R4656 VGND.n2553 VGND.n351 3.4105
R4657 VGND.n2680 VGND.n2679 3.4105
R4658 VGND.n2154 VGND.n2153 3.4105
R4659 VGND.n2156 VGND.n2155 3.4105
R4660 VGND.n2162 VGND.n2161 3.4105
R4661 VGND.n2164 VGND.n2163 3.4105
R4662 VGND.n2170 VGND.n2169 3.4105
R4663 VGND.n2066 VGND.n2065 3.4105
R4664 VGND.n2843 VGND.n262 3.4105
R4665 VGND.n2148 VGND.n2147 3.4105
R4666 VGND.n2150 VGND.n2149 3.4105
R4667 VGND.n1950 VGND.n437 3.4105
R4668 VGND.n2449 VGND.n2448 3.4105
R4669 VGND.n2451 VGND.n2450 3.4105
R4670 VGND.n2552 VGND.n391 3.4105
R4671 VGND.n2676 VGND.n2675 3.4105
R4672 VGND.n1790 VGND.n570 3.4105
R4673 VGND.n1780 VGND.n567 3.4105
R4674 VGND.n1779 VGND.n564 3.4105
R4675 VGND.n1769 VGND.n561 3.4105
R4676 VGND.n1768 VGND.n558 3.4105
R4677 VGND.n1758 VGND.n555 3.4105
R4678 VGND.n1901 VGND.n588 3.4105
R4679 VGND.n1830 VGND.n1737 3.4105
R4680 VGND.n1791 VGND.n573 3.4105
R4681 VGND.n2146 VGND.n2145 3.4105
R4682 VGND.n2144 VGND.n2143 3.4105
R4683 VGND.n1951 VGND.n433 3.4105
R4684 VGND.n2464 VGND.n2463 3.4105
R4685 VGND.n2462 VGND.n2461 3.4105
R4686 VGND.n2551 VGND.n321 3.4105
R4687 VGND.n2711 VGND.n2710 3.4105
R4688 VGND.n1867 VGND.n1866 3.4105
R4689 VGND.n1869 VGND.n1868 3.4105
R4690 VGND.n1875 VGND.n1874 3.4105
R4691 VGND.n1877 VGND.n1876 3.4105
R4692 VGND.n1883 VGND.n1882 3.4105
R4693 VGND.n1885 VGND.n1884 3.4105
R4694 VGND.n1686 VGND.n639 3.4105
R4695 VGND.n1899 VGND.n1898 3.4105
R4696 VGND.n1837 VGND.n1736 3.4105
R4697 VGND.n1861 VGND.n1860 3.4105
R4698 VGND.n1801 VGND.n576 3.4105
R4699 VGND.n2140 VGND.n2139 3.4105
R4700 VGND.n2142 VGND.n2141 3.4105
R4701 VGND.n1961 VGND.n429 3.4105
R4702 VGND.n2475 VGND.n2474 3.4105
R4703 VGND.n2477 VGND.n2476 3.4105
R4704 VGND.n2550 VGND.n317 3.4105
R4705 VGND.n2722 VGND.n2721 3.4105
R4706 VGND.n1863 VGND.n1862 3.4105
R4707 VGND.n1865 VGND.n1864 3.4105
R4708 VGND.n1871 VGND.n1870 3.4105
R4709 VGND.n1873 VGND.n1872 3.4105
R4710 VGND.n1879 VGND.n1878 3.4105
R4711 VGND.n1881 VGND.n1880 3.4105
R4712 VGND.n1887 VGND.n1886 3.4105
R4713 VGND.n1889 VGND.n1888 3.4105
R4714 VGND.n1897 VGND.n1896 3.4105
R4715 VGND.n2868 VGND.n250 3.4105
R4716 VGND.n1857 VGND.n1856 3.4105
R4717 VGND.n1859 VGND.n1858 3.4105
R4718 VGND.n1802 VGND.n579 3.4105
R4719 VGND.n2138 VGND.n2137 3.4105
R4720 VGND.n2136 VGND.n2135 3.4105
R4721 VGND.n1962 VGND.n425 3.4105
R4722 VGND.n2490 VGND.n2489 3.4105
R4723 VGND.n2488 VGND.n2487 3.4105
R4724 VGND.n2549 VGND.n305 3.4105
R4725 VGND.n2744 VGND.n2743 3.4105
R4726 VGND.n860 VGND.n663 3.4105
R4727 VGND.n861 VGND.n660 3.4105
R4728 VGND.n862 VGND.n657 3.4105
R4729 VGND.n863 VGND.n654 3.4105
R4730 VGND.n864 VGND.n651 3.4105
R4731 VGND.n865 VGND.n648 3.4105
R4732 VGND.n866 VGND.n645 3.4105
R4733 VGND.n867 VGND.n642 3.4105
R4734 VGND.n1891 VGND.n1890 3.4105
R4735 VGND.n1349 VGND.n630 3.4105
R4736 VGND.n1654 VGND.n737 3.4105
R4737 VGND.n1670 VGND.n1669 3.4105
R4738 VGND.n1855 VGND.n1854 3.4105
R4739 VGND.n1853 VGND.n1852 3.4105
R4740 VGND.n1812 VGND.n582 3.4105
R4741 VGND.n2132 VGND.n2131 3.4105
R4742 VGND.n2134 VGND.n2133 3.4105
R4743 VGND.n1972 VGND.n421 3.4105
R4744 VGND.n2506 VGND.n2505 3.4105
R4745 VGND.n2508 VGND.n2507 3.4105
R4746 VGND.n2548 VGND.n301 3.4105
R4747 VGND.n2760 VGND.n2759 3.4105
R4748 VGND.n1629 VGND.n731 3.4105
R4749 VGND.n1628 VGND.n1627 3.4105
R4750 VGND.n1559 VGND.n753 3.4105
R4751 VGND.n1561 VGND.n1560 3.4105
R4752 VGND.n1539 VGND.n1538 3.4105
R4753 VGND.n1524 VGND.n1523 3.4105
R4754 VGND.n1513 VGND.n1512 3.4105
R4755 VGND.n1498 VGND.n1497 3.4105
R4756 VGND.n1487 VGND.n1486 3.4105
R4757 VGND.n1402 VGND.n638 3.4105
R4758 VGND.n1405 VGND.n1404 3.4105
R4759 VGND.n1651 VGND.n738 3.4105
R4760 VGND.n2878 VGND.n2877 3.4105
R4761 VGND.n1668 VGND.n242 3.4105
R4762 VGND.n2855 VGND.n2854 3.4105
R4763 VGND.n2853 VGND.n2852 3.4105
R4764 VGND.n1813 VGND.n254 3.4105
R4765 VGND.n2830 VGND.n2829 3.4105
R4766 VGND.n2828 VGND.n2827 3.4105
R4767 VGND.n1973 VGND.n266 3.4105
R4768 VGND.n2805 VGND.n2804 3.4105
R4769 VGND.n2803 VGND.n2802 3.4105
R4770 VGND.n2547 VGND.n278 3.4105
R4771 VGND.n2783 VGND.n2782 3.4105
R4772 VGND.n2880 VGND.n2879 3.4105
R4773 VGND.n1624 VGND.n1623 3.4105
R4774 VGND.n1626 VGND.n1625 3.4105
R4775 VGND.n1589 VGND.n1588 3.4105
R4776 VGND.n1563 VGND.n1562 3.4105
R4777 VGND.n1537 VGND.n1536 3.4105
R4778 VGND.n1526 VGND.n1525 3.4105
R4779 VGND.n1511 VGND.n1510 3.4105
R4780 VGND.n1500 VGND.n1499 3.4105
R4781 VGND.n1485 VGND.n1484 3.4105
R4782 VGND.n1474 VGND.n1473 3.4105
R4783 VGND.n1407 VGND.n1406 3.4105
R4784 VGND.n2893 VGND.n237 3.4105
R4785 VGND.n2881 VGND.n230 3.4105
R4786 VGND.n2876 VGND.n2875 3.4105
R4787 VGND.n2874 VGND.n2873 3.4105
R4788 VGND.n2856 VGND.n245 3.4105
R4789 VGND.n2851 VGND.n2850 3.4105
R4790 VGND.n2849 VGND.n2848 3.4105
R4791 VGND.n2831 VGND.n257 3.4105
R4792 VGND.n2826 VGND.n2825 3.4105
R4793 VGND.n2824 VGND.n2823 3.4105
R4794 VGND.n2806 VGND.n269 3.4105
R4795 VGND.n2801 VGND.n2800 3.4105
R4796 VGND.n2799 VGND.n2798 3.4105
R4797 VGND.n2784 VGND.n281 3.4105
R4798 VGND.n2899 VGND.n2898 3.4105
R4799 VGND.n1620 VGND.n241 3.4105
R4800 VGND.n1622 VGND.n1621 3.4105
R4801 VGND.n1592 VGND.n743 3.4105
R4802 VGND.n1591 VGND.n1590 3.4105
R4803 VGND.n1465 VGND.n757 3.4105
R4804 VGND.n1466 VGND.n762 3.4105
R4805 VGND.n1467 VGND.n766 3.4105
R4806 VGND.n1468 VGND.n770 3.4105
R4807 VGND.n1469 VGND.n774 3.4105
R4808 VGND.n1470 VGND.n778 3.4105
R4809 VGND.n1472 VGND.n1471 3.4105
R4810 VGND.n1344 VGND.n798 3.4105
R4811 VGND.n1606 VGND.n1605 3.4105
R4812 VGND.n2897 VGND.n2896 3.4105
R4813 VGND.n2895 VGND.n2894 3.4105
R4814 VGND.n740 VGND.n235 3.4105
R4815 VGND.n2872 VGND.n2871 3.4105
R4816 VGND.n2870 VGND.n2869 3.4105
R4817 VGND.n1838 VGND.n248 3.4105
R4818 VGND.n2847 VGND.n2846 3.4105
R4819 VGND.n2845 VGND.n2844 3.4105
R4820 VGND.n1998 VGND.n260 3.4105
R4821 VGND.n2822 VGND.n2821 3.4105
R4822 VGND.n2820 VGND.n2819 3.4105
R4823 VGND.n419 VGND.n272 3.4105
R4824 VGND.n2797 VGND.n2796 3.4105
R4825 VGND.n2795 VGND.n2794 3.4105
R4826 VGND.n234 VGND.n233 3.4105
R4827 VGND.n2901 VGND.n2900 3.4105
R4828 VGND.n1064 VGND.n923 3.4105
R4829 VGND.n1065 VGND.n746 3.4105
R4830 VGND.n1066 VGND.n918 3.4105
R4831 VGND.n1067 VGND.n752 3.4105
R4832 VGND.n1304 VGND.n1303 3.4105
R4833 VGND.n1306 VGND.n1305 3.4105
R4834 VGND.n1312 VGND.n1311 3.4105
R4835 VGND.n1314 VGND.n1313 3.4105
R4836 VGND.n1320 VGND.n1319 3.4105
R4837 VGND.n1322 VGND.n1321 3.4105
R4838 VGND.n1101 VGND.n782 3.4105
R4839 VGND.n1104 VGND.n1103 3.4105
R4840 VGND.n2913 VGND.n226 3.4105
R4841 VGND.n1102 VGND.n792 3.4105
R4842 VGND.n1420 VGND.n1419 3.4105
R4843 VGND.n1418 VGND.n1417 3.4105
R4844 VGND.n1403 VGND.n635 3.4105
R4845 VGND.n1893 VGND.n1892 3.4105
R4846 VGND.n1895 VGND.n1894 3.4105
R4847 VGND.n1685 VGND.n551 3.4105
R4848 VGND.n2174 VGND.n2173 3.4105
R4849 VGND.n2172 VGND.n2171 3.4105
R4850 VGND.n2062 VGND.n552 3.4105
R4851 VGND.n1917 VGND.n461 3.4105
R4852 VGND.n2371 VGND.n2370 3.4105
R4853 VGND.n2373 VGND.n2372 3.4105
R4854 VGND.n2558 VGND.n336 3.4105
R4855 VGND.n2694 VGND.n2693 3.4105
R4856 VGND.n1285 VGND.n993 3.4105
R4857 VGND.n1271 VGND.n1270 3.4105
R4858 VGND.n1291 VGND.n922 3.4105
R4859 VGND.n1292 VGND.n921 3.4105
R4860 VGND.n1297 VGND.n917 3.4105
R4861 VGND.n1298 VGND.n916 3.4105
R4862 VGND.n1250 VGND.n913 3.4105
R4863 VGND.n1214 VGND.n910 3.4105
R4864 VGND.n1196 VGND.n907 3.4105
R4865 VGND.n1201 VGND.n904 3.4105
R4866 VGND.n1192 VGND.n901 3.4105
R4867 VGND.n1182 VGND.n898 3.4105
R4868 VGND.n1327 VGND.n892 3.4105
R4869 VGND.n1328 VGND.n891 3.4105
R4870 VGND.n1284 VGND.n1283 3.4105
R4871 VGND.n1267 VGND.n1266 3.4105
R4872 VGND.n1269 VGND.n1268 3.4105
R4873 VGND.n1264 VGND.n1263 3.4105
R4874 VGND.n1261 VGND.n1260 3.4105
R4875 VGND.n1258 VGND.n1257 3.4105
R4876 VGND.n1255 VGND.n1254 3.4105
R4877 VGND.n1252 VGND.n1251 3.4105
R4878 VGND.n1213 VGND.n999 3.4105
R4879 VGND.n1198 VGND.n1197 3.4105
R4880 VGND.n1200 VGND.n1199 3.4105
R4881 VGND.n1194 VGND.n1193 3.4105
R4882 VGND.n1181 VGND.n1005 3.4105
R4883 VGND.n1017 VGND.n1016 3.4105
R4884 VGND.n1020 VGND.n1019 3.4105
R4885 VGND.n1164 VGND.n1163 3.4105
R4886 VGND.n1287 VGND.n1286 3.4105
R4887 VGND.n1288 VGND.n229 3.4105
R4888 VGND.n1290 VGND.n1289 3.4105
R4889 VGND.n1294 VGND.n1293 3.4105
R4890 VGND.n1296 VGND.n1295 3.4105
R4891 VGND.n1300 VGND.n1299 3.4105
R4892 VGND.n1302 VGND.n1301 3.4105
R4893 VGND.n1308 VGND.n1307 3.4105
R4894 VGND.n1310 VGND.n1309 3.4105
R4895 VGND.n1316 VGND.n1315 3.4105
R4896 VGND.n1318 VGND.n1317 3.4105
R4897 VGND.n1324 VGND.n1323 3.4105
R4898 VGND.n1326 VGND.n1325 3.4105
R4899 VGND.n1330 VGND.n1329 3.4105
R4900 VGND.n1162 VGND.n1161 3.4105
R4901 VGND.n2916 VGND.n223 3.4105
R4902 VGND.n105 VGND.n104 3.01226
R4903 VGND.n2200 VGND.n2189 3.01226
R4904 VGND.n2184 VGND.n545 2.63579
R4905 VGND.n2565 VGND 2.52282
R4906 VGND.n2568 VGND 2.52282
R4907 VGND.n2571 VGND 2.52282
R4908 VGND.n2574 VGND 2.52282
R4909 VGND.n2577 VGND 2.52282
R4910 VGND.n2580 VGND 2.52282
R4911 VGND.n2583 VGND 2.52282
R4912 VGND.n2586 VGND 2.52282
R4913 VGND.n2589 VGND 2.52282
R4914 VGND.n2592 VGND 2.52282
R4915 VGND.n2595 VGND 2.52282
R4916 VGND.n2598 VGND 2.52282
R4917 VGND.n2601 VGND 2.52282
R4918 VGND.n2604 VGND 2.52282
R4919 VGND.n2607 VGND 2.52282
R4920 VGND.n186 VGND.n185 2.25932
R4921 VGND.n114 VGND.n93 2.25932
R4922 VGND.n110 VGND.n109 2.25932
R4923 VGND.n87 VGND.n86 2.25932
R4924 VGND.n155 VGND.n154 2.25932
R4925 VGND.n2205 VGND.n2204 2.25932
R4926 VGND.n491 VGND.n479 1.88285
R4927 VGND.n2272 VGND.n2260 1.88285
R4928 VGND.n527 VGND.n515 1.88285
R4929 VGND.n2608 VGND 1.79514
R4930 VGND.n1158 VGND.n224 1.76378
R4931 VGND.n2608 VGND 1.57193
R4932 VGND.n2940 VGND.n2939 1.54254
R4933 VGND.n2938 VGND.n2937 1.54254
R4934 VGND.n2533 VGND.n207 1.54254
R4935 VGND.n2530 VGND.n417 1.54254
R4936 VGND.n2818 VGND.n275 1.54254
R4937 VGND.n1991 VGND.n1990 1.54254
R4938 VGND.n1997 VGND.n1992 1.54254
R4939 VGND.n2843 VGND.n263 1.54254
R4940 VGND.n1831 VGND.n1830 1.54254
R4941 VGND.n1837 VGND.n1832 1.54254
R4942 VGND.n2868 VGND.n251 1.54254
R4943 VGND.n1654 VGND.n1653 1.54254
R4944 VGND.n1652 VGND.n1651 1.54254
R4945 VGND.n2893 VGND.n238 1.54254
R4946 VGND.n1606 VGND.n225 1.54254
R4947 VGND.n2914 VGND.n2913 1.54254
R4948 VGND.n1284 VGND.n224 1.54254
R4949 VGND.n2916 VGND.n2915 1.54254
R4950 VGND.n121 VGND.n120 1.50638
R4951 VGND.n2212 VGND.n544 1.50638
R4952 VGND VGND.n2562 1.3946
R4953 VGND.n2561 VGND 1.3946
R4954 VGND.n2560 VGND 1.3946
R4955 VGND VGND.n398 1.3946
R4956 VGND.n1905 VGND 1.3946
R4957 VGND VGND.n1906 1.3946
R4958 VGND.n1904 VGND 1.3946
R4959 VGND.n1903 VGND 1.3946
R4960 VGND.n1902 VGND 1.3946
R4961 VGND.n1900 VGND 1.3946
R4962 VGND VGND.n626 1.3946
R4963 VGND VGND.n1348 1.3946
R4964 VGND.n1347 VGND 1.3946
R4965 VGND.n1346 VGND 1.3946
R4966 VGND.n1345 VGND 1.3946
R4967 VGND VGND.n880 1.3946
R4968 VGND.n1159 VGND 1.3946
R4969 VGND VGND.n1160 1.3946
R4970 VGND.n1158 VGND.n1157 1.04899
R4971 VGND.n2696 VGND.n335 1.00149
R4972 VGND.n2627 VGND.n340 1.00149
R4973 VGND.n2624 VGND.n341 1.00149
R4974 VGND.n2621 VGND.n346 1.00149
R4975 VGND.n2618 VGND.n347 1.00149
R4976 VGND.n2615 VGND.n352 1.00149
R4977 VGND.n2612 VGND.n390 1.00149
R4978 VGND.n2708 VGND.n323 1.00149
R4979 VGND.n2724 VGND.n316 1.00149
R4980 VGND.n2741 VGND.n307 1.00149
R4981 VGND.n2763 VGND.n2762 1.00149
R4982 VGND.n2766 VGND.n289 1.00149
R4983 VGND.n2779 VGND.n291 1.00149
R4984 VGND.n2771 VGND.n2770 1.00149
R4985 VGND.n2941 VGND.n205 1.00149
R4986 VGND.n1019 VGND.n891 1.00149
R4987 VGND.n1016 VGND.n892 1.00149
R4988 VGND.n1182 VGND.n1181 1.00149
R4989 VGND.n1193 VGND.n1192 1.00149
R4990 VGND.n1201 VGND.n1200 1.00149
R4991 VGND.n1197 VGND.n1196 1.00149
R4992 VGND.n1214 VGND.n1213 1.00149
R4993 VGND.n1251 VGND.n1250 1.00149
R4994 VGND.n1254 VGND.n916 1.00149
R4995 VGND.n1257 VGND.n917 1.00149
R4996 VGND.n1260 VGND.n921 1.00149
R4997 VGND.n1263 VGND.n922 1.00149
R4998 VGND.n1271 VGND.n1269 1.00149
R4999 VGND.n1266 VGND.n993 1.00149
R5000 VGND.n1283 VGND.n995 1.00149
R5001 VGND.n1164 VGND.n1022 1.00149
R5002 VGND.n2632 VGND.n2631 0.973133
R5003 VGND.n2346 VGND.n2 0.9305
R5004 VGND.n178 VGND.n174 0.929432
R5005 VGND.n101 VGND.n99 0.929432
R5006 VGND.n79 VGND.n75 0.929432
R5007 VGND.n147 VGND.n143 0.929432
R5008 VGND.n126 VGND.n1 0.916608
R5009 VGND VGND.n2565 0.839786
R5010 VGND VGND.n2568 0.839786
R5011 VGND VGND.n2571 0.839786
R5012 VGND VGND.n2574 0.839786
R5013 VGND VGND.n2577 0.839786
R5014 VGND VGND.n2580 0.839786
R5015 VGND VGND.n2583 0.839786
R5016 VGND VGND.n2586 0.839786
R5017 VGND VGND.n2589 0.839786
R5018 VGND VGND.n2592 0.839786
R5019 VGND VGND.n2595 0.839786
R5020 VGND VGND.n2598 0.839786
R5021 VGND VGND.n2601 0.839786
R5022 VGND VGND.n2604 0.839786
R5023 VGND VGND.n2607 0.839786
R5024 VGND.n3023 VGND.n3022 0.7755
R5025 VGND.n3024 VGND.n3023 0.774207
R5026 VGND.n2981 VGND.n2978 0.753441
R5027 VGND.n20 VGND.n18 0.753441
R5028 VGND.n2953 VGND.n2951 0.753441
R5029 VGND.n46 VGND.n44 0.753441
R5030 VGND.n159 VGND.n136 0.753441
R5031 VGND.n2254 VGND.n2252 0.753441
R5032 VGND.n3025 VGND 0.706681
R5033 VGND VGND.n0 0.542567
R5034 VGND.n3025 VGND.n1 0.507317
R5035 VGND.n2939 VGND.n33 0.404308
R5036 VGND.n115 VGND.n114 0.376971
R5037 VGND.n120 VGND.n92 0.376971
R5038 VGND.n1140 VGND.n1137 0.376971
R5039 VGND.n1112 VGND.n1108 0.376971
R5040 VGND.n2212 VGND.n2211 0.376971
R5041 VGND.n2237 VGND.n2236 0.376971
R5042 VGND.n1375 VGND.n1374 0.376971
R5043 VGND VGND.n3025 0.37415
R5044 VGND.n226 VGND.n223 0.362676
R5045 VGND.n1605 VGND.n226 0.362676
R5046 VGND.n1605 VGND.n237 0.362676
R5047 VGND.n738 VGND.n237 0.362676
R5048 VGND.n738 VGND.n737 0.362676
R5049 VGND.n737 VGND.n250 0.362676
R5050 VGND.n1736 VGND.n250 0.362676
R5051 VGND.n1737 VGND.n1736 0.362676
R5052 VGND.n1737 VGND.n262 0.362676
R5053 VGND.n603 VGND.n262 0.362676
R5054 VGND.n604 VGND.n603 0.362676
R5055 VGND.n604 VGND.n274 0.362676
R5056 VGND.n2531 VGND.n274 0.362676
R5057 VGND.n2532 VGND.n2531 0.362676
R5058 VGND.n2532 VGND.n206 0.362676
R5059 VGND.n1162 VGND.n1104 0.362676
R5060 VGND.n1104 VGND.n798 0.362676
R5061 VGND.n1406 VGND.n798 0.362676
R5062 VGND.n1406 VGND.n1405 0.362676
R5063 VGND.n1405 VGND.n630 0.362676
R5064 VGND.n1897 VGND.n630 0.362676
R5065 VGND.n1898 VGND.n1897 0.362676
R5066 VGND.n1898 VGND.n588 0.362676
R5067 VGND.n2065 VGND.n588 0.362676
R5068 VGND.n2065 VGND.n2064 0.362676
R5069 VGND.n2064 VGND.n467 0.362676
R5070 VGND.n2359 VGND.n467 0.362676
R5071 VGND.n2359 VGND.n2358 0.362676
R5072 VGND.n2358 VGND.n397 0.362676
R5073 VGND.n2634 VGND.n397 0.362676
R5074 VGND.n1326 VGND.n782 0.362676
R5075 VGND.n1472 VGND.n782 0.362676
R5076 VGND.n1473 VGND.n1472 0.362676
R5077 VGND.n1473 VGND.n638 0.362676
R5078 VGND.n1890 VGND.n638 0.362676
R5079 VGND.n1890 VGND.n1889 0.362676
R5080 VGND.n1889 VGND.n639 0.362676
R5081 VGND.n639 VGND.n555 0.362676
R5082 VGND.n2169 VGND.n555 0.362676
R5083 VGND.n2169 VGND.n2168 0.362676
R5084 VGND.n2168 VGND.n457 0.362676
R5085 VGND.n2385 VGND.n457 0.362676
R5086 VGND.n2385 VGND.n2384 0.362676
R5087 VGND.n2384 VGND.n339 0.362676
R5088 VGND.n2691 VGND.n339 0.362676
R5089 VGND.n1323 VGND.n1322 0.362676
R5090 VGND.n1322 VGND.n778 0.362676
R5091 VGND.n1485 VGND.n778 0.362676
R5092 VGND.n1486 VGND.n1485 0.362676
R5093 VGND.n1486 VGND.n642 0.362676
R5094 VGND.n1886 VGND.n642 0.362676
R5095 VGND.n1886 VGND.n1885 0.362676
R5096 VGND.n1885 VGND.n558 0.362676
R5097 VGND.n2164 VGND.n558 0.362676
R5098 VGND.n2165 VGND.n2164 0.362676
R5099 VGND.n2165 VGND.n453 0.362676
R5100 VGND.n2397 VGND.n453 0.362676
R5101 VGND.n2398 VGND.n2397 0.362676
R5102 VGND.n2398 VGND.n342 0.362676
R5103 VGND.n2688 VGND.n342 0.362676
R5104 VGND.n1319 VGND.n1318 0.362676
R5105 VGND.n1319 VGND.n774 0.362676
R5106 VGND.n1499 VGND.n774 0.362676
R5107 VGND.n1499 VGND.n1498 0.362676
R5108 VGND.n1498 VGND.n645 0.362676
R5109 VGND.n1881 VGND.n645 0.362676
R5110 VGND.n1882 VGND.n1881 0.362676
R5111 VGND.n1882 VGND.n561 0.362676
R5112 VGND.n2161 VGND.n561 0.362676
R5113 VGND.n2161 VGND.n2160 0.362676
R5114 VGND.n2160 VGND.n449 0.362676
R5115 VGND.n2411 VGND.n449 0.362676
R5116 VGND.n2411 VGND.n2410 0.362676
R5117 VGND.n2410 VGND.n345 0.362676
R5118 VGND.n2685 VGND.n345 0.362676
R5119 VGND.n1315 VGND.n1314 0.362676
R5120 VGND.n1314 VGND.n770 0.362676
R5121 VGND.n1511 VGND.n770 0.362676
R5122 VGND.n1512 VGND.n1511 0.362676
R5123 VGND.n1512 VGND.n648 0.362676
R5124 VGND.n1878 VGND.n648 0.362676
R5125 VGND.n1878 VGND.n1877 0.362676
R5126 VGND.n1877 VGND.n564 0.362676
R5127 VGND.n2156 VGND.n564 0.362676
R5128 VGND.n2157 VGND.n2156 0.362676
R5129 VGND.n2157 VGND.n445 0.362676
R5130 VGND.n2423 VGND.n445 0.362676
R5131 VGND.n2424 VGND.n2423 0.362676
R5132 VGND.n2424 VGND.n348 0.362676
R5133 VGND.n2682 VGND.n348 0.362676
R5134 VGND.n1311 VGND.n1310 0.362676
R5135 VGND.n1311 VGND.n766 0.362676
R5136 VGND.n1525 VGND.n766 0.362676
R5137 VGND.n1525 VGND.n1524 0.362676
R5138 VGND.n1524 VGND.n651 0.362676
R5139 VGND.n1873 VGND.n651 0.362676
R5140 VGND.n1874 VGND.n1873 0.362676
R5141 VGND.n1874 VGND.n567 0.362676
R5142 VGND.n2153 VGND.n567 0.362676
R5143 VGND.n2153 VGND.n2152 0.362676
R5144 VGND.n2152 VGND.n441 0.362676
R5145 VGND.n2437 VGND.n441 0.362676
R5146 VGND.n2437 VGND.n2436 0.362676
R5147 VGND.n2436 VGND.n351 0.362676
R5148 VGND.n2679 VGND.n351 0.362676
R5149 VGND.n1307 VGND.n1306 0.362676
R5150 VGND.n1306 VGND.n762 0.362676
R5151 VGND.n1537 VGND.n762 0.362676
R5152 VGND.n1538 VGND.n1537 0.362676
R5153 VGND.n1538 VGND.n654 0.362676
R5154 VGND.n1870 VGND.n654 0.362676
R5155 VGND.n1870 VGND.n1869 0.362676
R5156 VGND.n1869 VGND.n570 0.362676
R5157 VGND.n2148 VGND.n570 0.362676
R5158 VGND.n2149 VGND.n2148 0.362676
R5159 VGND.n2149 VGND.n437 0.362676
R5160 VGND.n2449 VGND.n437 0.362676
R5161 VGND.n2450 VGND.n2449 0.362676
R5162 VGND.n2450 VGND.n391 0.362676
R5163 VGND.n2676 VGND.n391 0.362676
R5164 VGND.n1303 VGND.n1302 0.362676
R5165 VGND.n1303 VGND.n757 0.362676
R5166 VGND.n1562 VGND.n757 0.362676
R5167 VGND.n1562 VGND.n1561 0.362676
R5168 VGND.n1561 VGND.n657 0.362676
R5169 VGND.n1865 VGND.n657 0.362676
R5170 VGND.n1866 VGND.n1865 0.362676
R5171 VGND.n1866 VGND.n573 0.362676
R5172 VGND.n2145 VGND.n573 0.362676
R5173 VGND.n2145 VGND.n2144 0.362676
R5174 VGND.n2144 VGND.n433 0.362676
R5175 VGND.n2463 VGND.n433 0.362676
R5176 VGND.n2463 VGND.n2462 0.362676
R5177 VGND.n2462 VGND.n321 0.362676
R5178 VGND.n2710 VGND.n321 0.362676
R5179 VGND.n1299 VGND.n752 0.362676
R5180 VGND.n1590 VGND.n752 0.362676
R5181 VGND.n1590 VGND.n1589 0.362676
R5182 VGND.n1589 VGND.n753 0.362676
R5183 VGND.n753 VGND.n660 0.362676
R5184 VGND.n1862 VGND.n660 0.362676
R5185 VGND.n1862 VGND.n1861 0.362676
R5186 VGND.n1861 VGND.n576 0.362676
R5187 VGND.n2140 VGND.n576 0.362676
R5188 VGND.n2141 VGND.n2140 0.362676
R5189 VGND.n2141 VGND.n429 0.362676
R5190 VGND.n2475 VGND.n429 0.362676
R5191 VGND.n2476 VGND.n2475 0.362676
R5192 VGND.n2476 VGND.n317 0.362676
R5193 VGND.n2722 VGND.n317 0.362676
R5194 VGND.n1296 VGND.n918 0.362676
R5195 VGND.n918 VGND.n743 0.362676
R5196 VGND.n1626 VGND.n743 0.362676
R5197 VGND.n1627 VGND.n1626 0.362676
R5198 VGND.n1627 VGND.n663 0.362676
R5199 VGND.n1857 VGND.n663 0.362676
R5200 VGND.n1858 VGND.n1857 0.362676
R5201 VGND.n1858 VGND.n579 0.362676
R5202 VGND.n2137 VGND.n579 0.362676
R5203 VGND.n2137 VGND.n2136 0.362676
R5204 VGND.n2136 VGND.n425 0.362676
R5205 VGND.n2489 VGND.n425 0.362676
R5206 VGND.n2489 VGND.n2488 0.362676
R5207 VGND.n2488 VGND.n305 0.362676
R5208 VGND.n2743 VGND.n305 0.362676
R5209 VGND.n1293 VGND.n746 0.362676
R5210 VGND.n1622 VGND.n746 0.362676
R5211 VGND.n1623 VGND.n1622 0.362676
R5212 VGND.n1623 VGND.n731 0.362676
R5213 VGND.n1670 VGND.n731 0.362676
R5214 VGND.n1854 VGND.n1670 0.362676
R5215 VGND.n1854 VGND.n1853 0.362676
R5216 VGND.n1853 VGND.n582 0.362676
R5217 VGND.n2132 VGND.n582 0.362676
R5218 VGND.n2133 VGND.n2132 0.362676
R5219 VGND.n2133 VGND.n421 0.362676
R5220 VGND.n2506 VGND.n421 0.362676
R5221 VGND.n2507 VGND.n2506 0.362676
R5222 VGND.n2507 VGND.n301 0.362676
R5223 VGND.n2760 VGND.n301 0.362676
R5224 VGND.n1290 VGND.n923 0.362676
R5225 VGND.n923 VGND.n241 0.362676
R5226 VGND.n2879 VGND.n241 0.362676
R5227 VGND.n2879 VGND.n2878 0.362676
R5228 VGND.n2878 VGND.n242 0.362676
R5229 VGND.n2854 VGND.n242 0.362676
R5230 VGND.n2854 VGND.n2853 0.362676
R5231 VGND.n2853 VGND.n254 0.362676
R5232 VGND.n2829 VGND.n254 0.362676
R5233 VGND.n2829 VGND.n2828 0.362676
R5234 VGND.n2828 VGND.n266 0.362676
R5235 VGND.n2804 VGND.n266 0.362676
R5236 VGND.n2804 VGND.n2803 0.362676
R5237 VGND.n2803 VGND.n278 0.362676
R5238 VGND.n2782 VGND.n278 0.362676
R5239 VGND.n2900 VGND.n229 0.362676
R5240 VGND.n2900 VGND.n2899 0.362676
R5241 VGND.n2899 VGND.n230 0.362676
R5242 VGND.n2875 VGND.n230 0.362676
R5243 VGND.n2875 VGND.n2874 0.362676
R5244 VGND.n2874 VGND.n245 0.362676
R5245 VGND.n2850 VGND.n245 0.362676
R5246 VGND.n2850 VGND.n2849 0.362676
R5247 VGND.n2849 VGND.n257 0.362676
R5248 VGND.n2825 VGND.n257 0.362676
R5249 VGND.n2825 VGND.n2824 0.362676
R5250 VGND.n2824 VGND.n269 0.362676
R5251 VGND.n2800 VGND.n269 0.362676
R5252 VGND.n2800 VGND.n2799 0.362676
R5253 VGND.n2799 VGND.n281 0.362676
R5254 VGND.n1286 VGND.n234 0.362676
R5255 VGND.n2896 VGND.n234 0.362676
R5256 VGND.n2896 VGND.n2895 0.362676
R5257 VGND.n2895 VGND.n235 0.362676
R5258 VGND.n2871 VGND.n235 0.362676
R5259 VGND.n2871 VGND.n2870 0.362676
R5260 VGND.n2870 VGND.n248 0.362676
R5261 VGND.n2846 VGND.n248 0.362676
R5262 VGND.n2846 VGND.n2845 0.362676
R5263 VGND.n2845 VGND.n260 0.362676
R5264 VGND.n2821 VGND.n260 0.362676
R5265 VGND.n2821 VGND.n2820 0.362676
R5266 VGND.n2820 VGND.n272 0.362676
R5267 VGND.n2796 VGND.n272 0.362676
R5268 VGND.n2796 VGND.n2795 0.362676
R5269 VGND.n1329 VGND.n792 0.362676
R5270 VGND.n1419 VGND.n792 0.362676
R5271 VGND.n1419 VGND.n1418 0.362676
R5272 VGND.n1418 VGND.n635 0.362676
R5273 VGND.n1893 VGND.n635 0.362676
R5274 VGND.n1894 VGND.n1893 0.362676
R5275 VGND.n1894 VGND.n551 0.362676
R5276 VGND.n2173 VGND.n551 0.362676
R5277 VGND.n2173 VGND.n2172 0.362676
R5278 VGND.n2172 VGND.n552 0.362676
R5279 VGND.n552 VGND.n461 0.362676
R5280 VGND.n2371 VGND.n461 0.362676
R5281 VGND.n2372 VGND.n2371 0.362676
R5282 VGND.n2372 VGND.n336 0.362676
R5283 VGND.n2694 VGND.n336 0.362676
R5284 VGND.n2769 VGND.n2768 0.349144
R5285 VGND.n2768 VGND.n2767 0.349144
R5286 VGND.n2767 VGND.n2764 0.349144
R5287 VGND.n2764 VGND.n298 0.349144
R5288 VGND.n2609 VGND.n298 0.349144
R5289 VGND.n2610 VGND.n2609 0.349144
R5290 VGND.n2613 VGND.n2610 0.349144
R5291 VGND.n2616 VGND.n2613 0.349144
R5292 VGND.n2619 VGND.n2616 0.349144
R5293 VGND.n2622 VGND.n2619 0.349144
R5294 VGND.n2625 VGND.n2622 0.349144
R5295 VGND.n2628 VGND.n2625 0.349144
R5296 VGND.n2629 VGND.n2628 0.349144
R5297 VGND.n1268 VGND.n1267 0.349144
R5298 VGND.n1268 VGND.n1264 0.349144
R5299 VGND.n1264 VGND.n1261 0.349144
R5300 VGND.n1261 VGND.n1258 0.349144
R5301 VGND.n1258 VGND.n1255 0.349144
R5302 VGND.n1255 VGND.n1252 0.349144
R5303 VGND.n1252 VGND.n999 0.349144
R5304 VGND.n1198 VGND.n999 0.349144
R5305 VGND.n1199 VGND.n1198 0.349144
R5306 VGND.n1199 VGND.n1194 0.349144
R5307 VGND.n1194 VGND.n1005 0.349144
R5308 VGND.n1017 VGND.n1005 0.349144
R5309 VGND.n1020 VGND.n1017 0.349144
R5310 VGND.n2700 VGND.n331 0.327628
R5311 VGND.n2697 VGND.n333 0.327628
R5312 VGND.n361 VGND.n358 0.327628
R5313 VGND.n369 VGND.n365 0.327628
R5314 VGND.n372 VGND.n354 0.327628
R5315 VGND.n380 VGND.n376 0.327628
R5316 VGND.n383 VGND.n353 0.327628
R5317 VGND.n389 VGND.n388 0.327628
R5318 VGND.n2707 VGND.n2706 0.327628
R5319 VGND.n2727 VGND.n2725 0.327628
R5320 VGND.n2740 VGND.n2739 0.327628
R5321 VGND.n2736 VGND.n300 0.327628
R5322 VGND.n2733 VGND.n2732 0.327628
R5323 VGND.n2778 VGND.n2777 0.327628
R5324 VGND.n2774 VGND.n2772 0.327628
R5325 VGND.n2793 VGND.n2792 0.327628
R5326 VGND.n2789 VGND.n2785 0.327628
R5327 VGND.n2754 VGND.n288 0.327628
R5328 VGND.n2758 VGND.n2757 0.327628
R5329 VGND.n2749 VGND.n2745 0.327628
R5330 VGND.n2720 VGND.n2719 0.327628
R5331 VGND.n2716 VGND.n2712 0.327628
R5332 VGND.n2674 VGND.n2673 0.327628
R5333 VGND.n2670 VGND.n350 0.327628
R5334 VGND.n2665 VGND.n349 0.327628
R5335 VGND.n2660 VGND.n344 0.327628
R5336 VGND.n2655 VGND.n343 0.327628
R5337 VGND.n2650 VGND.n338 0.327628
R5338 VGND.n2645 VGND.n337 0.327628
R5339 VGND.n2640 VGND.n2636 0.327628
R5340 VGND.n2537 VGND.n283 0.327628
R5341 VGND.n2542 VGND.n282 0.327628
R5342 VGND.n2546 VGND.n2545 0.327628
R5343 VGND.n2289 VGND.n412 0.327628
R5344 VGND.n2294 VGND.n411 0.327628
R5345 VGND.n2299 VGND.n410 0.327628
R5346 VGND.n2304 VGND.n409 0.327628
R5347 VGND.n2309 VGND.n408 0.327628
R5348 VGND.n2314 VGND.n407 0.327628
R5349 VGND.n2319 VGND.n406 0.327628
R5350 VGND.n2324 VGND.n405 0.327628
R5351 VGND.n2329 VGND.n404 0.327628
R5352 VGND.n2334 VGND.n403 0.327628
R5353 VGND.n2339 VGND.n402 0.327628
R5354 VGND.n2344 VGND.n401 0.327628
R5355 VGND.n2526 VGND.n420 0.327628
R5356 VGND.n2523 VGND.n280 0.327628
R5357 VGND.n2518 VGND.n279 0.327628
R5358 VGND.n2513 VGND.n2509 0.327628
R5359 VGND.n2486 VGND.n2485 0.327628
R5360 VGND.n2482 VGND.n2478 0.327628
R5361 VGND.n2460 VGND.n2459 0.327628
R5362 VGND.n2456 VGND.n2452 0.327628
R5363 VGND.n2434 VGND.n2433 0.327628
R5364 VGND.n2430 VGND.n2426 0.327628
R5365 VGND.n2408 VGND.n2407 0.327628
R5366 VGND.n2404 VGND.n2400 0.327628
R5367 VGND.n2382 VGND.n2381 0.327628
R5368 VGND.n2378 VGND.n2374 0.327628
R5369 VGND.n2356 VGND.n2355 0.327628
R5370 VGND.n2814 VGND.n273 0.327628
R5371 VGND.n2811 VGND.n2807 0.327628
R5372 VGND.n2500 VGND.n277 0.327628
R5373 VGND.n2504 VGND.n2503 0.327628
R5374 VGND.n2495 VGND.n2491 0.327628
R5375 VGND.n2473 VGND.n2472 0.327628
R5376 VGND.n2469 VGND.n2465 0.327628
R5377 VGND.n2447 VGND.n2446 0.327628
R5378 VGND.n2443 VGND.n2439 0.327628
R5379 VGND.n2421 VGND.n2420 0.327628
R5380 VGND.n2417 VGND.n2413 0.327628
R5381 VGND.n2395 VGND.n2394 0.327628
R5382 VGND.n2391 VGND.n2387 0.327628
R5383 VGND.n2369 VGND.n2368 0.327628
R5384 VGND.n2365 VGND.n2361 0.327628
R5385 VGND.n1986 VGND.n271 0.327628
R5386 VGND.n1983 VGND.n270 0.327628
R5387 VGND.n1978 VGND.n1974 0.327628
R5388 VGND.n1971 VGND.n1970 0.327628
R5389 VGND.n1967 VGND.n1963 0.327628
R5390 VGND.n1960 VGND.n1959 0.327628
R5391 VGND.n1956 VGND.n1952 0.327628
R5392 VGND.n1949 VGND.n1948 0.327628
R5393 VGND.n1945 VGND.n1941 0.327628
R5394 VGND.n1938 VGND.n1937 0.327628
R5395 VGND.n1934 VGND.n1930 0.327628
R5396 VGND.n1927 VGND.n1926 0.327628
R5397 VGND.n1923 VGND.n1919 0.327628
R5398 VGND.n1916 VGND.n1915 0.327628
R5399 VGND.n1912 VGND.n1908 0.327628
R5400 VGND.n1999 VGND.n602 0.327628
R5401 VGND.n2002 VGND.n268 0.327628
R5402 VGND.n2007 VGND.n267 0.327628
R5403 VGND.n2012 VGND.n581 0.327628
R5404 VGND.n2017 VGND.n580 0.327628
R5405 VGND.n2022 VGND.n575 0.327628
R5406 VGND.n2027 VGND.n574 0.327628
R5407 VGND.n2032 VGND.n569 0.327628
R5408 VGND.n2037 VGND.n568 0.327628
R5409 VGND.n2042 VGND.n563 0.327628
R5410 VGND.n2047 VGND.n562 0.327628
R5411 VGND.n2052 VGND.n557 0.327628
R5412 VGND.n2057 VGND.n556 0.327628
R5413 VGND.n2061 VGND.n2060 0.327628
R5414 VGND.n598 VGND.n591 0.327628
R5415 VGND.n2839 VGND.n261 0.327628
R5416 VGND.n2836 VGND.n2832 0.327628
R5417 VGND.n2126 VGND.n265 0.327628
R5418 VGND.n2130 VGND.n2129 0.327628
R5419 VGND.n2121 VGND.n578 0.327628
R5420 VGND.n2116 VGND.n577 0.327628
R5421 VGND.n2111 VGND.n572 0.327628
R5422 VGND.n2106 VGND.n571 0.327628
R5423 VGND.n2101 VGND.n566 0.327628
R5424 VGND.n2096 VGND.n565 0.327628
R5425 VGND.n2091 VGND.n560 0.327628
R5426 VGND.n2086 VGND.n559 0.327628
R5427 VGND.n2081 VGND.n554 0.327628
R5428 VGND.n2076 VGND.n553 0.327628
R5429 VGND.n2071 VGND.n2067 0.327628
R5430 VGND.n1826 VGND.n259 0.327628
R5431 VGND.n1823 VGND.n258 0.327628
R5432 VGND.n1818 VGND.n1814 0.327628
R5433 VGND.n1811 VGND.n1810 0.327628
R5434 VGND.n1807 VGND.n1803 0.327628
R5435 VGND.n1800 VGND.n1799 0.327628
R5436 VGND.n1796 VGND.n1792 0.327628
R5437 VGND.n1789 VGND.n1788 0.327628
R5438 VGND.n1785 VGND.n1781 0.327628
R5439 VGND.n1778 VGND.n1777 0.327628
R5440 VGND.n1774 VGND.n1770 0.327628
R5441 VGND.n1767 VGND.n1766 0.327628
R5442 VGND.n1763 VGND.n1759 0.327628
R5443 VGND.n2175 VGND.n550 0.327628
R5444 VGND.n2178 VGND.n548 0.327628
R5445 VGND.n1839 VGND.n1735 0.327628
R5446 VGND.n1842 VGND.n256 0.327628
R5447 VGND.n1847 VGND.n255 0.327628
R5448 VGND.n1851 VGND.n1850 0.327628
R5449 VGND.n1731 VGND.n662 0.327628
R5450 VGND.n1726 VGND.n661 0.327628
R5451 VGND.n1721 VGND.n656 0.327628
R5452 VGND.n1716 VGND.n655 0.327628
R5453 VGND.n1711 VGND.n650 0.327628
R5454 VGND.n1706 VGND.n649 0.327628
R5455 VGND.n1701 VGND.n644 0.327628
R5456 VGND.n1696 VGND.n643 0.327628
R5457 VGND.n1691 VGND.n1687 0.327628
R5458 VGND.n1684 VGND.n1683 0.327628
R5459 VGND.n1680 VGND.n629 0.327628
R5460 VGND.n2864 VGND.n249 0.327628
R5461 VGND.n2861 VGND.n2857 0.327628
R5462 VGND.n726 VGND.n253 0.327628
R5463 VGND.n730 VGND.n729 0.327628
R5464 VGND.n721 VGND.n664 0.327628
R5465 VGND.n716 VGND.n659 0.327628
R5466 VGND.n711 VGND.n658 0.327628
R5467 VGND.n706 VGND.n653 0.327628
R5468 VGND.n701 VGND.n652 0.327628
R5469 VGND.n696 VGND.n647 0.327628
R5470 VGND.n691 VGND.n646 0.327628
R5471 VGND.n686 VGND.n641 0.327628
R5472 VGND.n681 VGND.n640 0.327628
R5473 VGND.n676 VGND.n634 0.327628
R5474 VGND.n671 VGND.n633 0.327628
R5475 VGND.n1658 VGND.n247 0.327628
R5476 VGND.n1663 VGND.n246 0.327628
R5477 VGND.n1667 VGND.n1666 0.327628
R5478 VGND.n855 VGND.n732 0.327628
R5479 VGND.n859 VGND.n858 0.327628
R5480 VGND.n850 VGND.n817 0.327628
R5481 VGND.n845 VGND.n816 0.327628
R5482 VGND.n840 VGND.n815 0.327628
R5483 VGND.n835 VGND.n814 0.327628
R5484 VGND.n830 VGND.n813 0.327628
R5485 VGND.n825 VGND.n812 0.327628
R5486 VGND.n868 VGND.n808 0.327628
R5487 VGND.n871 VGND.n637 0.327628
R5488 VGND.n876 VGND.n636 0.327628
R5489 VGND.n1354 VGND.n1350 0.327628
R5490 VGND.n1647 VGND.n741 0.327628
R5491 VGND.n1644 VGND.n244 0.327628
R5492 VGND.n1639 VGND.n243 0.327628
R5493 VGND.n1634 VGND.n1630 0.327628
R5494 VGND.n1554 VGND.n742 0.327628
R5495 VGND.n1558 VGND.n1557 0.327628
R5496 VGND.n1549 VGND.n758 0.327628
R5497 VGND.n1544 VGND.n1540 0.327628
R5498 VGND.n1522 VGND.n1521 0.327628
R5499 VGND.n1518 VGND.n1514 0.327628
R5500 VGND.n1496 VGND.n1495 0.327628
R5501 VGND.n1492 VGND.n1488 0.327628
R5502 VGND.n1401 VGND.n1400 0.327628
R5503 VGND.n1397 VGND.n802 0.327628
R5504 VGND.n1392 VGND.n801 0.327628
R5505 VGND.n2889 VGND.n236 0.327628
R5506 VGND.n2886 VGND.n2882 0.327628
R5507 VGND.n1573 VGND.n240 0.327628
R5508 VGND.n1578 VGND.n745 0.327628
R5509 VGND.n1583 VGND.n744 0.327628
R5510 VGND.n1587 VGND.n1586 0.327628
R5511 VGND.n1568 VGND.n1564 0.327628
R5512 VGND.n1535 VGND.n1534 0.327628
R5513 VGND.n1531 VGND.n1527 0.327628
R5514 VGND.n1509 VGND.n1508 0.327628
R5515 VGND.n1505 VGND.n1501 0.327628
R5516 VGND.n1483 VGND.n1482 0.327628
R5517 VGND.n1479 VGND.n1475 0.327628
R5518 VGND.n1416 VGND.n1415 0.327628
R5519 VGND.n1412 VGND.n1408 0.327628
R5520 VGND.n1610 VGND.n232 0.327628
R5521 VGND.n1615 VGND.n231 0.327628
R5522 VGND.n1619 VGND.n1618 0.327628
R5523 VGND.n1602 VGND.n747 0.327628
R5524 VGND.n1597 VGND.n1593 0.327628
R5525 VGND.n1460 VGND.n751 0.327628
R5526 VGND.n1464 VGND.n1463 0.327628
R5527 VGND.n1455 VGND.n788 0.327628
R5528 VGND.n1450 VGND.n787 0.327628
R5529 VGND.n1445 VGND.n786 0.327628
R5530 VGND.n1440 VGND.n785 0.327628
R5531 VGND.n1435 VGND.n784 0.327628
R5532 VGND.n1430 VGND.n783 0.327628
R5533 VGND.n1425 VGND.n1421 0.327628
R5534 VGND.n1343 VGND.n1342 0.327628
R5535 VGND.n2909 VGND.n228 0.327628
R5536 VGND.n2906 VGND.n2902 0.327628
R5537 VGND.n1063 VGND.n1062 0.327628
R5538 VGND.n1059 VGND.n1046 0.327628
R5539 VGND.n1054 VGND.n1045 0.327628
R5540 VGND.n1068 VGND.n1041 0.327628
R5541 VGND.n1071 VGND.n912 0.327628
R5542 VGND.n1076 VGND.n911 0.327628
R5543 VGND.n1081 VGND.n906 0.327628
R5544 VGND.n1086 VGND.n905 0.327628
R5545 VGND.n1091 VGND.n900 0.327628
R5546 VGND.n1096 VGND.n899 0.327628
R5547 VGND.n1100 VGND.n1099 0.327628
R5548 VGND.n1038 VGND.n1026 0.327628
R5549 VGND.n1033 VGND.n1025 0.327628
R5550 VGND.n1167 VGND.n1165 0.327628
R5551 VGND.n1174 VGND.n1170 0.327628
R5552 VGND.n1177 VGND.n1011 0.327628
R5553 VGND.n1187 VGND.n1183 0.327628
R5554 VGND.n1191 VGND.n1190 0.327628
R5555 VGND.n1206 VGND.n1202 0.327628
R5556 VGND.n1209 VGND.n1003 0.327628
R5557 VGND.n1219 VGND.n1215 0.327628
R5558 VGND.n1249 VGND.n1248 0.327628
R5559 VGND.n1245 VGND.n1223 0.327628
R5560 VGND.n1242 VGND.n1241 0.327628
R5561 VGND.n1238 VGND.n1228 0.327628
R5562 VGND.n1235 VGND.n1234 0.327628
R5563 VGND.n1276 VGND.n1272 0.327628
R5564 VGND.n1279 VGND.n997 0.327628
R5565 VGND.n992 VGND.n991 0.327628
R5566 VGND.n988 VGND.n925 0.327628
R5567 VGND.n983 VGND.n924 0.327628
R5568 VGND.n978 VGND.n920 0.327628
R5569 VGND.n973 VGND.n919 0.327628
R5570 VGND.n968 VGND.n915 0.327628
R5571 VGND.n963 VGND.n914 0.327628
R5572 VGND.n958 VGND.n909 0.327628
R5573 VGND.n953 VGND.n908 0.327628
R5574 VGND.n948 VGND.n903 0.327628
R5575 VGND.n943 VGND.n902 0.327628
R5576 VGND.n938 VGND.n897 0.327628
R5577 VGND.n933 VGND.n896 0.327628
R5578 VGND.n1331 VGND.n890 0.327628
R5579 VGND.n1334 VGND.n888 0.327628
R5580 VGND.n126 VGND.n125 0.213567
R5581 VGND.n125 VGND.n32 0.213567
R5582 VGND.n3002 VGND.n32 0.213567
R5583 VGND.n3002 VGND.n3001 0.213567
R5584 VGND.n1157 VGND.n1134 0.213567
R5585 VGND.n1134 VGND.n543 0.213567
R5586 VGND.n2219 VGND.n543 0.213567
R5587 VGND.n2219 VGND.n2218 0.213567
R5588 VGND.n2218 VGND.n0 0.213567
R5589 VGND.n3001 VGND.n33 0.2073
R5590 VGND.n3024 VGND.n2 0.18968
R5591 VGND.n1159 VGND.n1158 0.175967
R5592 VGND.n2633 VGND 0.169807
R5593 VGND.n2695 VGND 0.169807
R5594 VGND.n2690 VGND 0.169807
R5595 VGND.n2689 VGND 0.169807
R5596 VGND.n2684 VGND 0.169807
R5597 VGND.n2683 VGND 0.169807
R5598 VGND.n2678 VGND 0.169807
R5599 VGND.n2677 VGND 0.169807
R5600 VGND.n2709 VGND 0.169807
R5601 VGND.n2723 VGND 0.169807
R5602 VGND.n2742 VGND 0.169807
R5603 VGND.n2761 VGND 0.169807
R5604 VGND.n2781 VGND 0.169807
R5605 VGND.n2780 VGND 0.169807
R5606 VGND.n284 VGND 0.169807
R5607 VGND.n2635 VGND 0.169807
R5608 VGND.n2693 VGND 0.169807
R5609 VGND.n2692 VGND 0.169807
R5610 VGND.n2687 VGND 0.169807
R5611 VGND.n2686 VGND 0.169807
R5612 VGND.n2681 VGND 0.169807
R5613 VGND.n2680 VGND 0.169807
R5614 VGND.n2675 VGND 0.169807
R5615 VGND.n2711 VGND 0.169807
R5616 VGND.n2721 VGND 0.169807
R5617 VGND.n2744 VGND 0.169807
R5618 VGND.n2759 VGND 0.169807
R5619 VGND VGND.n2783 0.169807
R5620 VGND.n2784 VGND 0.169807
R5621 VGND.n2794 VGND 0.169807
R5622 VGND.n2559 VGND 0.169807
R5623 VGND.n2558 VGND 0.169807
R5624 VGND.n2557 VGND 0.169807
R5625 VGND.n2556 VGND 0.169807
R5626 VGND.n2555 VGND 0.169807
R5627 VGND.n2554 VGND 0.169807
R5628 VGND.n2553 VGND 0.169807
R5629 VGND.n2552 VGND 0.169807
R5630 VGND.n2551 VGND 0.169807
R5631 VGND.n2550 VGND 0.169807
R5632 VGND.n2549 VGND 0.169807
R5633 VGND.n2548 VGND 0.169807
R5634 VGND.n2547 VGND 0.169807
R5635 VGND.n2798 VGND 0.169807
R5636 VGND.n2797 VGND 0.169807
R5637 VGND.n2357 VGND 0.169807
R5638 VGND.n2373 VGND 0.169807
R5639 VGND.n2383 VGND 0.169807
R5640 VGND.n2399 VGND 0.169807
R5641 VGND.n2409 VGND 0.169807
R5642 VGND.n2425 VGND 0.169807
R5643 VGND.n2435 VGND 0.169807
R5644 VGND.n2451 VGND 0.169807
R5645 VGND.n2461 VGND 0.169807
R5646 VGND.n2477 VGND 0.169807
R5647 VGND.n2487 VGND 0.169807
R5648 VGND.n2508 VGND 0.169807
R5649 VGND.n2802 VGND 0.169807
R5650 VGND.n2801 VGND 0.169807
R5651 VGND.n419 VGND 0.169807
R5652 VGND.n2360 VGND 0.169807
R5653 VGND.n2370 VGND 0.169807
R5654 VGND.n2386 VGND 0.169807
R5655 VGND.n2396 VGND 0.169807
R5656 VGND.n2412 VGND 0.169807
R5657 VGND.n2422 VGND 0.169807
R5658 VGND.n2438 VGND 0.169807
R5659 VGND.n2448 VGND 0.169807
R5660 VGND.n2464 VGND 0.169807
R5661 VGND.n2474 VGND 0.169807
R5662 VGND.n2490 VGND 0.169807
R5663 VGND.n2505 VGND 0.169807
R5664 VGND VGND.n2805 0.169807
R5665 VGND.n2806 VGND 0.169807
R5666 VGND.n2819 VGND 0.169807
R5667 VGND.n1907 VGND 0.169807
R5668 VGND VGND.n1917 0.169807
R5669 VGND.n1918 VGND 0.169807
R5670 VGND VGND.n1928 0.169807
R5671 VGND.n1929 VGND 0.169807
R5672 VGND VGND.n1939 0.169807
R5673 VGND.n1940 VGND 0.169807
R5674 VGND VGND.n1950 0.169807
R5675 VGND.n1951 VGND 0.169807
R5676 VGND VGND.n1961 0.169807
R5677 VGND.n1962 VGND 0.169807
R5678 VGND VGND.n1972 0.169807
R5679 VGND.n1973 VGND 0.169807
R5680 VGND.n2823 VGND 0.169807
R5681 VGND.n2822 VGND 0.169807
R5682 VGND.n2063 VGND 0.169807
R5683 VGND.n2062 VGND 0.169807
R5684 VGND.n2167 VGND 0.169807
R5685 VGND.n2166 VGND 0.169807
R5686 VGND.n2159 VGND 0.169807
R5687 VGND.n2158 VGND 0.169807
R5688 VGND.n2151 VGND 0.169807
R5689 VGND.n2150 VGND 0.169807
R5690 VGND.n2143 VGND 0.169807
R5691 VGND.n2142 VGND 0.169807
R5692 VGND.n2135 VGND 0.169807
R5693 VGND.n2134 VGND 0.169807
R5694 VGND.n2827 VGND 0.169807
R5695 VGND.n2826 VGND 0.169807
R5696 VGND.n1998 VGND 0.169807
R5697 VGND.n2066 VGND 0.169807
R5698 VGND.n2171 VGND 0.169807
R5699 VGND.n2170 VGND 0.169807
R5700 VGND.n2163 VGND 0.169807
R5701 VGND.n2162 VGND 0.169807
R5702 VGND.n2155 VGND 0.169807
R5703 VGND.n2154 VGND 0.169807
R5704 VGND.n2147 VGND 0.169807
R5705 VGND.n2146 VGND 0.169807
R5706 VGND.n2139 VGND 0.169807
R5707 VGND.n2138 VGND 0.169807
R5708 VGND.n2131 VGND 0.169807
R5709 VGND VGND.n2830 0.169807
R5710 VGND.n2831 VGND 0.169807
R5711 VGND.n2844 VGND 0.169807
R5712 VGND.n1901 VGND 0.169807
R5713 VGND.n2174 VGND 0.169807
R5714 VGND.n1758 VGND 0.169807
R5715 VGND VGND.n1768 0.169807
R5716 VGND.n1769 VGND 0.169807
R5717 VGND VGND.n1779 0.169807
R5718 VGND.n1780 VGND 0.169807
R5719 VGND VGND.n1790 0.169807
R5720 VGND.n1791 VGND 0.169807
R5721 VGND VGND.n1801 0.169807
R5722 VGND.n1802 VGND 0.169807
R5723 VGND VGND.n1812 0.169807
R5724 VGND.n1813 VGND 0.169807
R5725 VGND.n2848 VGND 0.169807
R5726 VGND.n2847 VGND 0.169807
R5727 VGND.n1899 VGND 0.169807
R5728 VGND VGND.n1685 0.169807
R5729 VGND.n1686 VGND 0.169807
R5730 VGND.n1884 VGND 0.169807
R5731 VGND.n1883 VGND 0.169807
R5732 VGND.n1876 VGND 0.169807
R5733 VGND.n1875 VGND 0.169807
R5734 VGND.n1868 VGND 0.169807
R5735 VGND.n1867 VGND 0.169807
R5736 VGND.n1860 VGND 0.169807
R5737 VGND.n1859 VGND 0.169807
R5738 VGND.n1852 VGND 0.169807
R5739 VGND.n2852 VGND 0.169807
R5740 VGND.n2851 VGND 0.169807
R5741 VGND.n1838 VGND 0.169807
R5742 VGND.n1896 VGND 0.169807
R5743 VGND.n1895 VGND 0.169807
R5744 VGND.n1888 VGND 0.169807
R5745 VGND.n1887 VGND 0.169807
R5746 VGND.n1880 VGND 0.169807
R5747 VGND.n1879 VGND 0.169807
R5748 VGND.n1872 VGND 0.169807
R5749 VGND.n1871 VGND 0.169807
R5750 VGND.n1864 VGND 0.169807
R5751 VGND.n1863 VGND 0.169807
R5752 VGND.n1856 VGND 0.169807
R5753 VGND.n1855 VGND 0.169807
R5754 VGND VGND.n2855 0.169807
R5755 VGND.n2856 VGND 0.169807
R5756 VGND.n2869 VGND 0.169807
R5757 VGND.n1349 VGND 0.169807
R5758 VGND.n1892 VGND 0.169807
R5759 VGND.n1891 VGND 0.169807
R5760 VGND.n867 VGND 0.169807
R5761 VGND.n866 VGND 0.169807
R5762 VGND.n865 VGND 0.169807
R5763 VGND.n864 VGND 0.169807
R5764 VGND.n863 VGND 0.169807
R5765 VGND.n862 VGND 0.169807
R5766 VGND.n861 VGND 0.169807
R5767 VGND.n860 VGND 0.169807
R5768 VGND.n1669 VGND 0.169807
R5769 VGND.n1668 VGND 0.169807
R5770 VGND.n2873 VGND 0.169807
R5771 VGND.n2872 VGND 0.169807
R5772 VGND.n1404 VGND 0.169807
R5773 VGND.n1403 VGND 0.169807
R5774 VGND.n1402 VGND 0.169807
R5775 VGND.n1487 VGND 0.169807
R5776 VGND.n1497 VGND 0.169807
R5777 VGND.n1513 VGND 0.169807
R5778 VGND.n1523 VGND 0.169807
R5779 VGND.n1539 VGND 0.169807
R5780 VGND.n1560 VGND 0.169807
R5781 VGND.n1559 VGND 0.169807
R5782 VGND VGND.n1628 0.169807
R5783 VGND.n1629 VGND 0.169807
R5784 VGND.n2877 VGND 0.169807
R5785 VGND.n2876 VGND 0.169807
R5786 VGND.n740 VGND 0.169807
R5787 VGND.n1407 VGND 0.169807
R5788 VGND.n1417 VGND 0.169807
R5789 VGND.n1474 VGND 0.169807
R5790 VGND.n1484 VGND 0.169807
R5791 VGND.n1500 VGND 0.169807
R5792 VGND.n1510 VGND 0.169807
R5793 VGND.n1526 VGND 0.169807
R5794 VGND.n1536 VGND 0.169807
R5795 VGND.n1563 VGND 0.169807
R5796 VGND.n1588 VGND 0.169807
R5797 VGND.n1625 VGND 0.169807
R5798 VGND.n1624 VGND 0.169807
R5799 VGND VGND.n2880 0.169807
R5800 VGND.n2881 VGND 0.169807
R5801 VGND.n2894 VGND 0.169807
R5802 VGND.n1344 VGND 0.169807
R5803 VGND.n1420 VGND 0.169807
R5804 VGND.n1471 VGND 0.169807
R5805 VGND.n1470 VGND 0.169807
R5806 VGND.n1469 VGND 0.169807
R5807 VGND.n1468 VGND 0.169807
R5808 VGND.n1467 VGND 0.169807
R5809 VGND.n1466 VGND 0.169807
R5810 VGND.n1465 VGND 0.169807
R5811 VGND VGND.n1591 0.169807
R5812 VGND.n1592 VGND 0.169807
R5813 VGND.n1621 VGND 0.169807
R5814 VGND.n1620 VGND 0.169807
R5815 VGND.n2898 VGND 0.169807
R5816 VGND.n2897 VGND 0.169807
R5817 VGND.n1103 VGND 0.169807
R5818 VGND.n1102 VGND 0.169807
R5819 VGND.n1101 VGND 0.169807
R5820 VGND.n1321 VGND 0.169807
R5821 VGND.n1320 VGND 0.169807
R5822 VGND.n1313 VGND 0.169807
R5823 VGND.n1312 VGND 0.169807
R5824 VGND.n1305 VGND 0.169807
R5825 VGND.n1304 VGND 0.169807
R5826 VGND.n1067 VGND 0.169807
R5827 VGND.n1066 VGND 0.169807
R5828 VGND.n1065 VGND 0.169807
R5829 VGND.n1064 VGND 0.169807
R5830 VGND.n2901 VGND 0.169807
R5831 VGND.n233 VGND 0.169807
R5832 VGND.n1163 VGND 0.169807
R5833 VGND.n1328 VGND 0.169807
R5834 VGND.n1327 VGND 0.169807
R5835 VGND VGND.n898 0.169807
R5836 VGND VGND.n901 0.169807
R5837 VGND VGND.n904 0.169807
R5838 VGND VGND.n907 0.169807
R5839 VGND VGND.n910 0.169807
R5840 VGND VGND.n913 0.169807
R5841 VGND.n1298 VGND 0.169807
R5842 VGND.n1297 VGND 0.169807
R5843 VGND.n1292 VGND 0.169807
R5844 VGND.n1291 VGND 0.169807
R5845 VGND.n1270 VGND 0.169807
R5846 VGND.n1285 VGND 0.169807
R5847 VGND.n1161 VGND 0.169807
R5848 VGND.n1330 VGND 0.169807
R5849 VGND.n1325 VGND 0.169807
R5850 VGND.n1324 VGND 0.169807
R5851 VGND.n1317 VGND 0.169807
R5852 VGND.n1316 VGND 0.169807
R5853 VGND.n1309 VGND 0.169807
R5854 VGND.n1308 VGND 0.169807
R5855 VGND.n1301 VGND 0.169807
R5856 VGND.n1300 VGND 0.169807
R5857 VGND.n1295 VGND 0.169807
R5858 VGND.n1294 VGND 0.169807
R5859 VGND.n1289 VGND 0.169807
R5860 VGND.n1288 VGND 0.169807
R5861 VGND.n1287 VGND 0.169807
R5862 VGND.n190 VGND 0.159538
R5863 VGND.n161 VGND 0.159538
R5864 VGND.n2915 VGND.n224 0.154425
R5865 VGND.n2915 VGND.n2914 0.154425
R5866 VGND.n2914 VGND.n225 0.154425
R5867 VGND.n238 VGND.n225 0.154425
R5868 VGND.n1652 VGND.n238 0.154425
R5869 VGND.n1653 VGND.n1652 0.154425
R5870 VGND.n1653 VGND.n251 0.154425
R5871 VGND.n1832 VGND.n251 0.154425
R5872 VGND.n1832 VGND.n1831 0.154425
R5873 VGND.n1831 VGND.n263 0.154425
R5874 VGND.n1992 VGND.n263 0.154425
R5875 VGND.n1992 VGND.n1991 0.154425
R5876 VGND.n1991 VGND.n275 0.154425
R5877 VGND.n417 VGND.n275 0.154425
R5878 VGND.n417 VGND.n207 0.154425
R5879 VGND.n2938 VGND.n207 0.154425
R5880 VGND.n2939 VGND.n2938 0.154425
R5881 VGND.n1160 VGND.n1159 0.154425
R5882 VGND.n1160 VGND.n880 0.154425
R5883 VGND.n1345 VGND.n880 0.154425
R5884 VGND.n1346 VGND.n1345 0.154425
R5885 VGND.n1347 VGND.n1346 0.154425
R5886 VGND.n1348 VGND.n1347 0.154425
R5887 VGND.n1348 VGND.n626 0.154425
R5888 VGND.n1900 VGND.n626 0.154425
R5889 VGND.n1902 VGND.n1900 0.154425
R5890 VGND.n1903 VGND.n1902 0.154425
R5891 VGND.n1904 VGND.n1903 0.154425
R5892 VGND.n1906 VGND.n1904 0.154425
R5893 VGND.n1906 VGND.n1905 0.154425
R5894 VGND.n1905 VGND.n398 0.154425
R5895 VGND.n2560 VGND.n398 0.154425
R5896 VGND.n2561 VGND.n2560 0.154425
R5897 VGND.n2562 VGND.n2561 0.154425
R5898 VGND.n1144 VGND.n1138 0.144904
R5899 VGND.n1117 VGND.n1109 0.144904
R5900 VGND.n2232 VGND.n2228 0.144904
R5901 VGND.n1370 VGND.n1366 0.144904
R5902 VGND.n2632 VGND.n2608 0.138284
R5903 VGND.n2700 VGND.n2699 0.13638
R5904 VGND.n355 VGND.n333 0.13638
R5905 VGND.n362 VGND.n361 0.13638
R5906 VGND.n369 VGND.n368 0.13638
R5907 VGND.n373 VGND.n372 0.13638
R5908 VGND.n380 VGND.n379 0.13638
R5909 VGND.n384 VGND.n383 0.13638
R5910 VGND.n388 VGND.n387 0.13638
R5911 VGND.n2706 VGND.n326 0.13638
R5912 VGND.n2727 VGND.n2726 0.13638
R5913 VGND.n2739 VGND.n312 0.13638
R5914 VGND.n2736 VGND.n2735 0.13638
R5915 VGND.n2732 VGND.n2730 0.13638
R5916 VGND.n2777 VGND.n294 0.13638
R5917 VGND.n2774 VGND.n2773 0.13638
R5918 VGND.n2792 VGND.n287 0.13638
R5919 VGND.n2789 VGND.n2788 0.13638
R5920 VGND.n2754 VGND.n2753 0.13638
R5921 VGND.n2757 VGND.n304 0.13638
R5922 VGND.n2749 VGND.n2748 0.13638
R5923 VGND.n2719 VGND.n320 0.13638
R5924 VGND.n2716 VGND.n2715 0.13638
R5925 VGND.n2673 VGND.n394 0.13638
R5926 VGND.n2670 VGND.n2669 0.13638
R5927 VGND.n2665 VGND.n2664 0.13638
R5928 VGND.n2660 VGND.n2659 0.13638
R5929 VGND.n2655 VGND.n2654 0.13638
R5930 VGND.n2650 VGND.n2649 0.13638
R5931 VGND.n2645 VGND.n2644 0.13638
R5932 VGND.n2640 VGND.n2639 0.13638
R5933 VGND.n2537 VGND.n2536 0.13638
R5934 VGND.n2542 VGND.n2541 0.13638
R5935 VGND.n2545 VGND.n415 0.13638
R5936 VGND.n2289 VGND.n2288 0.13638
R5937 VGND.n2294 VGND.n2293 0.13638
R5938 VGND.n2299 VGND.n2298 0.13638
R5939 VGND.n2304 VGND.n2303 0.13638
R5940 VGND.n2309 VGND.n2308 0.13638
R5941 VGND.n2314 VGND.n2313 0.13638
R5942 VGND.n2319 VGND.n2318 0.13638
R5943 VGND.n2324 VGND.n2323 0.13638
R5944 VGND.n2329 VGND.n2328 0.13638
R5945 VGND.n2334 VGND.n2333 0.13638
R5946 VGND.n2339 VGND.n2338 0.13638
R5947 VGND.n2344 VGND.n2343 0.13638
R5948 VGND.n2527 VGND.n2526 0.13638
R5949 VGND.n2523 VGND.n2522 0.13638
R5950 VGND.n2518 VGND.n2517 0.13638
R5951 VGND.n2513 VGND.n2512 0.13638
R5952 VGND.n2485 VGND.n428 0.13638
R5953 VGND.n2482 VGND.n2481 0.13638
R5954 VGND.n2459 VGND.n436 0.13638
R5955 VGND.n2456 VGND.n2455 0.13638
R5956 VGND.n2433 VGND.n444 0.13638
R5957 VGND.n2430 VGND.n2429 0.13638
R5958 VGND.n2407 VGND.n452 0.13638
R5959 VGND.n2404 VGND.n2403 0.13638
R5960 VGND.n2381 VGND.n460 0.13638
R5961 VGND.n2378 VGND.n2377 0.13638
R5962 VGND.n2355 VGND.n472 0.13638
R5963 VGND.n2815 VGND.n2814 0.13638
R5964 VGND.n2811 VGND.n2810 0.13638
R5965 VGND.n2500 VGND.n2499 0.13638
R5966 VGND.n2503 VGND.n424 0.13638
R5967 VGND.n2495 VGND.n2494 0.13638
R5968 VGND.n2472 VGND.n432 0.13638
R5969 VGND.n2469 VGND.n2468 0.13638
R5970 VGND.n2446 VGND.n440 0.13638
R5971 VGND.n2443 VGND.n2442 0.13638
R5972 VGND.n2420 VGND.n448 0.13638
R5973 VGND.n2417 VGND.n2416 0.13638
R5974 VGND.n2394 VGND.n456 0.13638
R5975 VGND.n2391 VGND.n2390 0.13638
R5976 VGND.n2368 VGND.n464 0.13638
R5977 VGND.n2365 VGND.n2364 0.13638
R5978 VGND.n1987 VGND.n1986 0.13638
R5979 VGND.n1983 VGND.n1982 0.13638
R5980 VGND.n1978 VGND.n1977 0.13638
R5981 VGND.n1970 VGND.n608 0.13638
R5982 VGND.n1967 VGND.n1966 0.13638
R5983 VGND.n1959 VGND.n611 0.13638
R5984 VGND.n1956 VGND.n1955 0.13638
R5985 VGND.n1948 VGND.n614 0.13638
R5986 VGND.n1945 VGND.n1944 0.13638
R5987 VGND.n1937 VGND.n617 0.13638
R5988 VGND.n1934 VGND.n1933 0.13638
R5989 VGND.n1926 VGND.n620 0.13638
R5990 VGND.n1923 VGND.n1922 0.13638
R5991 VGND.n1915 VGND.n623 0.13638
R5992 VGND.n1912 VGND.n1911 0.13638
R5993 VGND.n1994 VGND.n602 0.13638
R5994 VGND.n2002 VGND.n2001 0.13638
R5995 VGND.n2007 VGND.n2006 0.13638
R5996 VGND.n2012 VGND.n2011 0.13638
R5997 VGND.n2017 VGND.n2016 0.13638
R5998 VGND.n2022 VGND.n2021 0.13638
R5999 VGND.n2027 VGND.n2026 0.13638
R6000 VGND.n2032 VGND.n2031 0.13638
R6001 VGND.n2037 VGND.n2036 0.13638
R6002 VGND.n2042 VGND.n2041 0.13638
R6003 VGND.n2047 VGND.n2046 0.13638
R6004 VGND.n2052 VGND.n2051 0.13638
R6005 VGND.n2057 VGND.n2056 0.13638
R6006 VGND.n2060 VGND.n594 0.13638
R6007 VGND.n598 VGND.n597 0.13638
R6008 VGND.n2840 VGND.n2839 0.13638
R6009 VGND.n2836 VGND.n2835 0.13638
R6010 VGND.n2126 VGND.n2125 0.13638
R6011 VGND.n2129 VGND.n585 0.13638
R6012 VGND.n2121 VGND.n2120 0.13638
R6013 VGND.n2116 VGND.n2115 0.13638
R6014 VGND.n2111 VGND.n2110 0.13638
R6015 VGND.n2106 VGND.n2105 0.13638
R6016 VGND.n2101 VGND.n2100 0.13638
R6017 VGND.n2096 VGND.n2095 0.13638
R6018 VGND.n2091 VGND.n2090 0.13638
R6019 VGND.n2086 VGND.n2085 0.13638
R6020 VGND.n2081 VGND.n2080 0.13638
R6021 VGND.n2076 VGND.n2075 0.13638
R6022 VGND.n2071 VGND.n2070 0.13638
R6023 VGND.n1827 VGND.n1826 0.13638
R6024 VGND.n1823 VGND.n1822 0.13638
R6025 VGND.n1818 VGND.n1817 0.13638
R6026 VGND.n1810 VGND.n1741 0.13638
R6027 VGND.n1807 VGND.n1806 0.13638
R6028 VGND.n1799 VGND.n1744 0.13638
R6029 VGND.n1796 VGND.n1795 0.13638
R6030 VGND.n1788 VGND.n1747 0.13638
R6031 VGND.n1785 VGND.n1784 0.13638
R6032 VGND.n1777 VGND.n1750 0.13638
R6033 VGND.n1774 VGND.n1773 0.13638
R6034 VGND.n1766 VGND.n1753 0.13638
R6035 VGND.n1763 VGND.n1762 0.13638
R6036 VGND.n1756 VGND.n550 0.13638
R6037 VGND.n2178 VGND.n2177 0.13638
R6038 VGND.n1834 VGND.n1735 0.13638
R6039 VGND.n1842 VGND.n1841 0.13638
R6040 VGND.n1847 VGND.n1846 0.13638
R6041 VGND.n1850 VGND.n1673 0.13638
R6042 VGND.n1731 VGND.n1730 0.13638
R6043 VGND.n1726 VGND.n1725 0.13638
R6044 VGND.n1721 VGND.n1720 0.13638
R6045 VGND.n1716 VGND.n1715 0.13638
R6046 VGND.n1711 VGND.n1710 0.13638
R6047 VGND.n1706 VGND.n1705 0.13638
R6048 VGND.n1701 VGND.n1700 0.13638
R6049 VGND.n1696 VGND.n1695 0.13638
R6050 VGND.n1691 VGND.n1690 0.13638
R6051 VGND.n1683 VGND.n1676 0.13638
R6052 VGND.n1680 VGND.n1679 0.13638
R6053 VGND.n2865 VGND.n2864 0.13638
R6054 VGND.n2861 VGND.n2860 0.13638
R6055 VGND.n726 VGND.n725 0.13638
R6056 VGND.n729 VGND.n667 0.13638
R6057 VGND.n721 VGND.n720 0.13638
R6058 VGND.n716 VGND.n715 0.13638
R6059 VGND.n711 VGND.n710 0.13638
R6060 VGND.n706 VGND.n705 0.13638
R6061 VGND.n701 VGND.n700 0.13638
R6062 VGND.n696 VGND.n695 0.13638
R6063 VGND.n691 VGND.n690 0.13638
R6064 VGND.n686 VGND.n685 0.13638
R6065 VGND.n681 VGND.n680 0.13638
R6066 VGND.n676 VGND.n675 0.13638
R6067 VGND.n671 VGND.n670 0.13638
R6068 VGND.n1658 VGND.n1657 0.13638
R6069 VGND.n1663 VGND.n1662 0.13638
R6070 VGND.n1666 VGND.n735 0.13638
R6071 VGND.n855 VGND.n854 0.13638
R6072 VGND.n858 VGND.n820 0.13638
R6073 VGND.n850 VGND.n849 0.13638
R6074 VGND.n845 VGND.n844 0.13638
R6075 VGND.n840 VGND.n839 0.13638
R6076 VGND.n835 VGND.n834 0.13638
R6077 VGND.n830 VGND.n829 0.13638
R6078 VGND.n825 VGND.n824 0.13638
R6079 VGND.n810 VGND.n808 0.13638
R6080 VGND.n871 VGND.n870 0.13638
R6081 VGND.n876 VGND.n875 0.13638
R6082 VGND.n1354 VGND.n1353 0.13638
R6083 VGND.n1648 VGND.n1647 0.13638
R6084 VGND.n1644 VGND.n1643 0.13638
R6085 VGND.n1639 VGND.n1638 0.13638
R6086 VGND.n1634 VGND.n1633 0.13638
R6087 VGND.n1554 VGND.n1553 0.13638
R6088 VGND.n1557 VGND.n761 0.13638
R6089 VGND.n1549 VGND.n1548 0.13638
R6090 VGND.n1544 VGND.n1543 0.13638
R6091 VGND.n1521 VGND.n769 0.13638
R6092 VGND.n1518 VGND.n1517 0.13638
R6093 VGND.n1495 VGND.n777 0.13638
R6094 VGND.n1492 VGND.n1491 0.13638
R6095 VGND.n1400 VGND.n805 0.13638
R6096 VGND.n1397 VGND.n1396 0.13638
R6097 VGND.n1392 VGND.n1391 0.13638
R6098 VGND.n2890 VGND.n2889 0.13638
R6099 VGND.n2886 VGND.n2885 0.13638
R6100 VGND.n1573 VGND.n1572 0.13638
R6101 VGND.n1578 VGND.n1577 0.13638
R6102 VGND.n1583 VGND.n1582 0.13638
R6103 VGND.n1586 VGND.n756 0.13638
R6104 VGND.n1568 VGND.n1567 0.13638
R6105 VGND.n1534 VGND.n765 0.13638
R6106 VGND.n1531 VGND.n1530 0.13638
R6107 VGND.n1508 VGND.n773 0.13638
R6108 VGND.n1505 VGND.n1504 0.13638
R6109 VGND.n1482 VGND.n781 0.13638
R6110 VGND.n1479 VGND.n1478 0.13638
R6111 VGND.n1415 VGND.n795 0.13638
R6112 VGND.n1412 VGND.n1411 0.13638
R6113 VGND.n1610 VGND.n1609 0.13638
R6114 VGND.n1615 VGND.n1614 0.13638
R6115 VGND.n1618 VGND.n750 0.13638
R6116 VGND.n1602 VGND.n1601 0.13638
R6117 VGND.n1597 VGND.n1596 0.13638
R6118 VGND.n1460 VGND.n1459 0.13638
R6119 VGND.n1463 VGND.n791 0.13638
R6120 VGND.n1455 VGND.n1454 0.13638
R6121 VGND.n1450 VGND.n1449 0.13638
R6122 VGND.n1445 VGND.n1444 0.13638
R6123 VGND.n1440 VGND.n1439 0.13638
R6124 VGND.n1435 VGND.n1434 0.13638
R6125 VGND.n1430 VGND.n1429 0.13638
R6126 VGND.n1425 VGND.n1424 0.13638
R6127 VGND.n1342 VGND.n885 0.13638
R6128 VGND.n2910 VGND.n2909 0.13638
R6129 VGND.n2906 VGND.n2905 0.13638
R6130 VGND.n1062 VGND.n1049 0.13638
R6131 VGND.n1059 VGND.n1058 0.13638
R6132 VGND.n1054 VGND.n1053 0.13638
R6133 VGND.n1043 VGND.n1041 0.13638
R6134 VGND.n1071 VGND.n1070 0.13638
R6135 VGND.n1076 VGND.n1075 0.13638
R6136 VGND.n1081 VGND.n1080 0.13638
R6137 VGND.n1086 VGND.n1085 0.13638
R6138 VGND.n1091 VGND.n1090 0.13638
R6139 VGND.n1096 VGND.n1095 0.13638
R6140 VGND.n1099 VGND.n1029 0.13638
R6141 VGND.n1038 VGND.n1037 0.13638
R6142 VGND.n1033 VGND.n1032 0.13638
R6143 VGND.n1168 VGND.n1167 0.13638
R6144 VGND.n1174 VGND.n1173 0.13638
R6145 VGND.n1178 VGND.n1177 0.13638
R6146 VGND.n1187 VGND.n1186 0.13638
R6147 VGND.n1190 VGND.n1009 0.13638
R6148 VGND.n1206 VGND.n1205 0.13638
R6149 VGND.n1210 VGND.n1209 0.13638
R6150 VGND.n1219 VGND.n1218 0.13638
R6151 VGND.n1248 VGND.n1001 0.13638
R6152 VGND.n1245 VGND.n1244 0.13638
R6153 VGND.n1241 VGND.n1225 0.13638
R6154 VGND.n1238 VGND.n1237 0.13638
R6155 VGND.n1234 VGND.n1232 0.13638
R6156 VGND.n1276 VGND.n1275 0.13638
R6157 VGND.n1280 VGND.n1279 0.13638
R6158 VGND.n991 VGND.n928 0.13638
R6159 VGND.n988 VGND.n987 0.13638
R6160 VGND.n983 VGND.n982 0.13638
R6161 VGND.n978 VGND.n977 0.13638
R6162 VGND.n973 VGND.n972 0.13638
R6163 VGND.n968 VGND.n967 0.13638
R6164 VGND.n963 VGND.n962 0.13638
R6165 VGND.n958 VGND.n957 0.13638
R6166 VGND.n953 VGND.n952 0.13638
R6167 VGND.n948 VGND.n947 0.13638
R6168 VGND.n943 VGND.n942 0.13638
R6169 VGND.n938 VGND.n937 0.13638
R6170 VGND.n933 VGND.n932 0.13638
R6171 VGND.n894 VGND.n890 0.13638
R6172 VGND.n1334 VGND.n1333 0.13638
R6173 VGND VGND.n190 0.120838
R6174 VGND.n19 VGND.n13 0.120292
R6175 VGND.n24 VGND.n13 0.120292
R6176 VGND.n25 VGND.n24 0.120292
R6177 VGND.n26 VGND.n25 0.120292
R6178 VGND.n26 VGND.n11 0.120292
R6179 VGND.n30 VGND.n11 0.120292
R6180 VGND.n31 VGND.n30 0.120292
R6181 VGND.n3008 VGND.n3007 0.120292
R6182 VGND.n3007 VGND.n3003 0.120292
R6183 VGND.n182 VGND.n174 0.120292
R6184 VGND.n183 VGND.n182 0.120292
R6185 VGND.n183 VGND.n168 0.120292
R6186 VGND.n188 VGND.n168 0.120292
R6187 VGND.n189 VGND.n188 0.120292
R6188 VGND.n2952 VGND.n2948 0.120292
R6189 VGND.n2957 VGND.n2948 0.120292
R6190 VGND.n2958 VGND.n2957 0.120292
R6191 VGND.n2959 VGND.n2958 0.120292
R6192 VGND.n2959 VGND.n2946 0.120292
R6193 VGND.n2963 VGND.n2946 0.120292
R6194 VGND.n2964 VGND.n2963 0.120292
R6195 VGND.n45 VGND.n39 0.120292
R6196 VGND.n50 VGND.n39 0.120292
R6197 VGND.n51 VGND.n50 0.120292
R6198 VGND.n52 VGND.n51 0.120292
R6199 VGND.n52 VGND.n37 0.120292
R6200 VGND.n56 VGND.n37 0.120292
R6201 VGND.n57 VGND.n56 0.120292
R6202 VGND.n63 VGND.n62 0.120292
R6203 VGND.n62 VGND.n58 0.120292
R6204 VGND.n106 VGND.n99 0.120292
R6205 VGND.n107 VGND.n106 0.120292
R6206 VGND.n107 VGND.n94 0.120292
R6207 VGND.n112 VGND.n94 0.120292
R6208 VGND.n113 VGND.n112 0.120292
R6209 VGND.n124 VGND.n91 0.120292
R6210 VGND.n83 VGND.n75 0.120292
R6211 VGND.n84 VGND.n83 0.120292
R6212 VGND.n84 VGND.n69 0.120292
R6213 VGND.n89 VGND.n69 0.120292
R6214 VGND.n90 VGND.n89 0.120292
R6215 VGND.n130 VGND.n127 0.120292
R6216 VGND.n151 VGND.n143 0.120292
R6217 VGND.n152 VGND.n151 0.120292
R6218 VGND.n152 VGND.n137 0.120292
R6219 VGND.n157 VGND.n137 0.120292
R6220 VGND.n158 VGND.n157 0.120292
R6221 VGND.n1152 VGND.n1151 0.120292
R6222 VGND.n1151 VGND.n1150 0.120292
R6223 VGND.n1150 VGND.n1136 0.120292
R6224 VGND.n1146 VGND.n1136 0.120292
R6225 VGND.n1146 VGND.n1145 0.120292
R6226 VGND.n1145 VGND.n1144 0.120292
R6227 VGND.n1130 VGND.n1129 0.120292
R6228 VGND.n1125 VGND.n1124 0.120292
R6229 VGND.n1124 VGND.n1123 0.120292
R6230 VGND.n1123 VGND.n1107 0.120292
R6231 VGND.n1119 VGND.n1107 0.120292
R6232 VGND.n1119 VGND.n1118 0.120292
R6233 VGND.n1118 VGND.n1117 0.120292
R6234 VGND.n499 VGND.n476 0.120292
R6235 VGND.n493 VGND.n476 0.120292
R6236 VGND.n493 VGND.n492 0.120292
R6237 VGND.n492 VGND.n480 0.120292
R6238 VGND.n485 VGND.n480 0.120292
R6239 VGND.n485 VGND.n484 0.120292
R6240 VGND.n484 VGND.n483 0.120292
R6241 VGND.n2280 VGND.n2257 0.120292
R6242 VGND.n2274 VGND.n2257 0.120292
R6243 VGND.n2274 VGND.n2273 0.120292
R6244 VGND.n2273 VGND.n2261 0.120292
R6245 VGND.n2266 VGND.n2261 0.120292
R6246 VGND.n2266 VGND.n2265 0.120292
R6247 VGND.n2265 VGND.n2264 0.120292
R6248 VGND.n510 VGND.n507 0.120292
R6249 VGND.n511 VGND.n510 0.120292
R6250 VGND.n535 VGND.n512 0.120292
R6251 VGND.n529 VGND.n512 0.120292
R6252 VGND.n529 VGND.n528 0.120292
R6253 VGND.n528 VGND.n516 0.120292
R6254 VGND.n521 VGND.n516 0.120292
R6255 VGND.n521 VGND.n520 0.120292
R6256 VGND.n520 VGND.n519 0.120292
R6257 VGND.n2214 VGND.n2213 0.120292
R6258 VGND.n2207 VGND.n2183 0.120292
R6259 VGND.n2202 VGND.n2183 0.120292
R6260 VGND.n2202 VGND.n2201 0.120292
R6261 VGND.n2198 VGND.n2197 0.120292
R6262 VGND.n2197 VGND.n2192 0.120292
R6263 VGND.n2193 VGND.n2192 0.120292
R6264 VGND.n2225 VGND.n2224 0.120292
R6265 VGND.n2245 VGND.n2244 0.120292
R6266 VGND.n2244 VGND.n2226 0.120292
R6267 VGND.n2240 VGND.n2226 0.120292
R6268 VGND.n2240 VGND.n2239 0.120292
R6269 VGND.n2239 VGND.n2238 0.120292
R6270 VGND.n2238 VGND.n2228 0.120292
R6271 VGND.n1363 VGND.n1362 0.120292
R6272 VGND.n1383 VGND.n1382 0.120292
R6273 VGND.n1382 VGND.n1364 0.120292
R6274 VGND.n1378 VGND.n1364 0.120292
R6275 VGND.n1378 VGND.n1377 0.120292
R6276 VGND.n1377 VGND.n1376 0.120292
R6277 VGND.n1376 VGND.n1366 0.120292
R6278 VGND.n2983 VGND.n2982 0.120292
R6279 VGND.n2983 VGND.n2975 0.120292
R6280 VGND.n2988 VGND.n2975 0.120292
R6281 VGND.n2989 VGND.n2988 0.120292
R6282 VGND.n2990 VGND.n2989 0.120292
R6283 VGND.n2990 VGND.n2973 0.120292
R6284 VGND.n2994 VGND.n2973 0.120292
R6285 VGND.n2996 VGND.n34 0.120292
R6286 VGND.n3000 VGND.n34 0.120292
R6287 VGND VGND.n161 0.119536
R6288 VGND.n1138 VGND 0.117202
R6289 VGND.n1109 VGND 0.117202
R6290 VGND.n2232 VGND 0.117202
R6291 VGND.n1370 VGND 0.117202
R6292 VGND.n287 VGND.n286 0.110872
R6293 VGND.n2788 VGND.n2787 0.110872
R6294 VGND.n2753 VGND.n2752 0.110872
R6295 VGND.n304 VGND.n303 0.110872
R6296 VGND.n2748 VGND.n2747 0.110872
R6297 VGND.n320 VGND.n319 0.110872
R6298 VGND.n2715 VGND.n2714 0.110872
R6299 VGND.n394 VGND.n393 0.110872
R6300 VGND.n2669 VGND.n2668 0.110872
R6301 VGND.n2664 VGND.n2663 0.110872
R6302 VGND.n2659 VGND.n2658 0.110872
R6303 VGND.n2654 VGND.n2653 0.110872
R6304 VGND.n2649 VGND.n2648 0.110872
R6305 VGND.n2644 VGND.n2643 0.110872
R6306 VGND.n2639 VGND.n2638 0.110872
R6307 VGND.n2536 VGND.n2535 0.110872
R6308 VGND.n2541 VGND.n2540 0.110872
R6309 VGND.n415 VGND.n414 0.110872
R6310 VGND.n2288 VGND.n2287 0.110872
R6311 VGND.n2293 VGND.n2292 0.110872
R6312 VGND.n2298 VGND.n2297 0.110872
R6313 VGND.n2303 VGND.n2302 0.110872
R6314 VGND.n2308 VGND.n2307 0.110872
R6315 VGND.n2313 VGND.n2312 0.110872
R6316 VGND.n2318 VGND.n2317 0.110872
R6317 VGND.n2323 VGND.n2322 0.110872
R6318 VGND.n2328 VGND.n2327 0.110872
R6319 VGND.n2333 VGND.n2332 0.110872
R6320 VGND.n2338 VGND.n2337 0.110872
R6321 VGND.n2343 VGND.n2342 0.110872
R6322 VGND.n2528 VGND.n2527 0.110872
R6323 VGND.n2522 VGND.n2521 0.110872
R6324 VGND.n2517 VGND.n2516 0.110872
R6325 VGND.n2512 VGND.n2511 0.110872
R6326 VGND.n428 VGND.n427 0.110872
R6327 VGND.n2481 VGND.n2480 0.110872
R6328 VGND.n436 VGND.n435 0.110872
R6329 VGND.n2455 VGND.n2454 0.110872
R6330 VGND.n444 VGND.n443 0.110872
R6331 VGND.n2429 VGND.n2428 0.110872
R6332 VGND.n452 VGND.n451 0.110872
R6333 VGND.n2403 VGND.n2402 0.110872
R6334 VGND.n460 VGND.n459 0.110872
R6335 VGND.n2377 VGND.n2376 0.110872
R6336 VGND.n472 VGND.n471 0.110872
R6337 VGND.n2816 VGND.n2815 0.110872
R6338 VGND.n2810 VGND.n2809 0.110872
R6339 VGND.n2499 VGND.n2498 0.110872
R6340 VGND.n424 VGND.n423 0.110872
R6341 VGND.n2494 VGND.n2493 0.110872
R6342 VGND.n432 VGND.n431 0.110872
R6343 VGND.n2468 VGND.n2467 0.110872
R6344 VGND.n440 VGND.n439 0.110872
R6345 VGND.n2442 VGND.n2441 0.110872
R6346 VGND.n448 VGND.n447 0.110872
R6347 VGND.n2416 VGND.n2415 0.110872
R6348 VGND.n456 VGND.n455 0.110872
R6349 VGND.n2390 VGND.n2389 0.110872
R6350 VGND.n464 VGND.n463 0.110872
R6351 VGND.n2364 VGND.n2363 0.110872
R6352 VGND.n1988 VGND.n1987 0.110872
R6353 VGND.n1982 VGND.n1981 0.110872
R6354 VGND.n1977 VGND.n1976 0.110872
R6355 VGND.n608 VGND.n607 0.110872
R6356 VGND.n1966 VGND.n1965 0.110872
R6357 VGND.n611 VGND.n610 0.110872
R6358 VGND.n1955 VGND.n1954 0.110872
R6359 VGND.n614 VGND.n613 0.110872
R6360 VGND.n1944 VGND.n1943 0.110872
R6361 VGND.n617 VGND.n616 0.110872
R6362 VGND.n1933 VGND.n1932 0.110872
R6363 VGND.n620 VGND.n619 0.110872
R6364 VGND.n1922 VGND.n1921 0.110872
R6365 VGND.n623 VGND.n622 0.110872
R6366 VGND.n1911 VGND.n1910 0.110872
R6367 VGND.n1995 VGND.n1994 0.110872
R6368 VGND.n2001 VGND.n2000 0.110872
R6369 VGND.n2006 VGND.n2005 0.110872
R6370 VGND.n2011 VGND.n2010 0.110872
R6371 VGND.n2016 VGND.n2015 0.110872
R6372 VGND.n2021 VGND.n2020 0.110872
R6373 VGND.n2026 VGND.n2025 0.110872
R6374 VGND.n2031 VGND.n2030 0.110872
R6375 VGND.n2036 VGND.n2035 0.110872
R6376 VGND.n2041 VGND.n2040 0.110872
R6377 VGND.n2046 VGND.n2045 0.110872
R6378 VGND.n2051 VGND.n2050 0.110872
R6379 VGND.n2056 VGND.n2055 0.110872
R6380 VGND.n594 VGND.n593 0.110872
R6381 VGND.n597 VGND.n596 0.110872
R6382 VGND.n2841 VGND.n2840 0.110872
R6383 VGND.n2835 VGND.n2834 0.110872
R6384 VGND.n2125 VGND.n2124 0.110872
R6385 VGND.n585 VGND.n584 0.110872
R6386 VGND.n2120 VGND.n2119 0.110872
R6387 VGND.n2115 VGND.n2114 0.110872
R6388 VGND.n2110 VGND.n2109 0.110872
R6389 VGND.n2105 VGND.n2104 0.110872
R6390 VGND.n2100 VGND.n2099 0.110872
R6391 VGND.n2095 VGND.n2094 0.110872
R6392 VGND.n2090 VGND.n2089 0.110872
R6393 VGND.n2085 VGND.n2084 0.110872
R6394 VGND.n2080 VGND.n2079 0.110872
R6395 VGND.n2075 VGND.n2074 0.110872
R6396 VGND.n2070 VGND.n2069 0.110872
R6397 VGND.n1828 VGND.n1827 0.110872
R6398 VGND.n1822 VGND.n1821 0.110872
R6399 VGND.n1817 VGND.n1816 0.110872
R6400 VGND.n1741 VGND.n1740 0.110872
R6401 VGND.n1806 VGND.n1805 0.110872
R6402 VGND.n1744 VGND.n1743 0.110872
R6403 VGND.n1795 VGND.n1794 0.110872
R6404 VGND.n1747 VGND.n1746 0.110872
R6405 VGND.n1784 VGND.n1783 0.110872
R6406 VGND.n1750 VGND.n1749 0.110872
R6407 VGND.n1773 VGND.n1772 0.110872
R6408 VGND.n1753 VGND.n1752 0.110872
R6409 VGND.n1762 VGND.n1761 0.110872
R6410 VGND.n1757 VGND.n1756 0.110872
R6411 VGND.n2177 VGND.n2176 0.110872
R6412 VGND.n1835 VGND.n1834 0.110872
R6413 VGND.n1841 VGND.n1840 0.110872
R6414 VGND.n1846 VGND.n1845 0.110872
R6415 VGND.n1673 VGND.n1672 0.110872
R6416 VGND.n1730 VGND.n1729 0.110872
R6417 VGND.n1725 VGND.n1724 0.110872
R6418 VGND.n1720 VGND.n1719 0.110872
R6419 VGND.n1715 VGND.n1714 0.110872
R6420 VGND.n1710 VGND.n1709 0.110872
R6421 VGND.n1705 VGND.n1704 0.110872
R6422 VGND.n1700 VGND.n1699 0.110872
R6423 VGND.n1695 VGND.n1694 0.110872
R6424 VGND.n1690 VGND.n1689 0.110872
R6425 VGND.n1676 VGND.n1675 0.110872
R6426 VGND.n1679 VGND.n1678 0.110872
R6427 VGND.n2866 VGND.n2865 0.110872
R6428 VGND.n2860 VGND.n2859 0.110872
R6429 VGND.n725 VGND.n724 0.110872
R6430 VGND.n667 VGND.n666 0.110872
R6431 VGND.n720 VGND.n719 0.110872
R6432 VGND.n715 VGND.n714 0.110872
R6433 VGND.n710 VGND.n709 0.110872
R6434 VGND.n705 VGND.n704 0.110872
R6435 VGND.n700 VGND.n699 0.110872
R6436 VGND.n695 VGND.n694 0.110872
R6437 VGND.n690 VGND.n689 0.110872
R6438 VGND.n685 VGND.n684 0.110872
R6439 VGND.n680 VGND.n679 0.110872
R6440 VGND.n675 VGND.n674 0.110872
R6441 VGND.n670 VGND.n669 0.110872
R6442 VGND.n1657 VGND.n1656 0.110872
R6443 VGND.n1662 VGND.n1661 0.110872
R6444 VGND.n735 VGND.n734 0.110872
R6445 VGND.n854 VGND.n853 0.110872
R6446 VGND.n820 VGND.n819 0.110872
R6447 VGND.n849 VGND.n848 0.110872
R6448 VGND.n844 VGND.n843 0.110872
R6449 VGND.n839 VGND.n838 0.110872
R6450 VGND.n834 VGND.n833 0.110872
R6451 VGND.n829 VGND.n828 0.110872
R6452 VGND.n824 VGND.n823 0.110872
R6453 VGND.n811 VGND.n810 0.110872
R6454 VGND.n870 VGND.n869 0.110872
R6455 VGND.n875 VGND.n874 0.110872
R6456 VGND.n1353 VGND.n1352 0.110872
R6457 VGND.n1649 VGND.n1648 0.110872
R6458 VGND.n1643 VGND.n1642 0.110872
R6459 VGND.n1638 VGND.n1637 0.110872
R6460 VGND.n1633 VGND.n1632 0.110872
R6461 VGND.n1553 VGND.n1552 0.110872
R6462 VGND.n761 VGND.n760 0.110872
R6463 VGND.n1548 VGND.n1547 0.110872
R6464 VGND.n1543 VGND.n1542 0.110872
R6465 VGND.n769 VGND.n768 0.110872
R6466 VGND.n1517 VGND.n1516 0.110872
R6467 VGND.n777 VGND.n776 0.110872
R6468 VGND.n1491 VGND.n1490 0.110872
R6469 VGND.n805 VGND.n804 0.110872
R6470 VGND.n1396 VGND.n1395 0.110872
R6471 VGND.n1391 VGND.n1390 0.110872
R6472 VGND.n2891 VGND.n2890 0.110872
R6473 VGND.n2885 VGND.n2884 0.110872
R6474 VGND.n1572 VGND.n1571 0.110872
R6475 VGND.n1577 VGND.n1576 0.110872
R6476 VGND.n1582 VGND.n1581 0.110872
R6477 VGND.n756 VGND.n755 0.110872
R6478 VGND.n1567 VGND.n1566 0.110872
R6479 VGND.n765 VGND.n764 0.110872
R6480 VGND.n1530 VGND.n1529 0.110872
R6481 VGND.n773 VGND.n772 0.110872
R6482 VGND.n1504 VGND.n1503 0.110872
R6483 VGND.n781 VGND.n780 0.110872
R6484 VGND.n1478 VGND.n1477 0.110872
R6485 VGND.n795 VGND.n794 0.110872
R6486 VGND.n1411 VGND.n1410 0.110872
R6487 VGND.n1609 VGND.n1608 0.110872
R6488 VGND.n1614 VGND.n1613 0.110872
R6489 VGND.n750 VGND.n749 0.110872
R6490 VGND.n1601 VGND.n1600 0.110872
R6491 VGND.n1596 VGND.n1595 0.110872
R6492 VGND.n1459 VGND.n1458 0.110872
R6493 VGND.n791 VGND.n790 0.110872
R6494 VGND.n1454 VGND.n1453 0.110872
R6495 VGND.n1449 VGND.n1448 0.110872
R6496 VGND.n1444 VGND.n1443 0.110872
R6497 VGND.n1439 VGND.n1438 0.110872
R6498 VGND.n1434 VGND.n1433 0.110872
R6499 VGND.n1429 VGND.n1428 0.110872
R6500 VGND.n1424 VGND.n1423 0.110872
R6501 VGND.n885 VGND.n884 0.110872
R6502 VGND.n2911 VGND.n2910 0.110872
R6503 VGND.n2905 VGND.n2904 0.110872
R6504 VGND.n1049 VGND.n1048 0.110872
R6505 VGND.n1058 VGND.n1057 0.110872
R6506 VGND.n1053 VGND.n1052 0.110872
R6507 VGND.n1044 VGND.n1043 0.110872
R6508 VGND.n1070 VGND.n1069 0.110872
R6509 VGND.n1075 VGND.n1074 0.110872
R6510 VGND.n1080 VGND.n1079 0.110872
R6511 VGND.n1085 VGND.n1084 0.110872
R6512 VGND.n1090 VGND.n1089 0.110872
R6513 VGND.n1095 VGND.n1094 0.110872
R6514 VGND.n1029 VGND.n1028 0.110872
R6515 VGND.n1037 VGND.n1036 0.110872
R6516 VGND.n1032 VGND.n1031 0.110872
R6517 VGND.n1169 VGND.n1168 0.110872
R6518 VGND.n1173 VGND.n1172 0.110872
R6519 VGND.n1179 VGND.n1178 0.110872
R6520 VGND.n1186 VGND.n1185 0.110872
R6521 VGND.n1009 VGND.n1008 0.110872
R6522 VGND.n1205 VGND.n1204 0.110872
R6523 VGND.n1211 VGND.n1210 0.110872
R6524 VGND.n1218 VGND.n1217 0.110872
R6525 VGND.n1222 VGND.n1001 0.110872
R6526 VGND.n1244 VGND.n1243 0.110872
R6527 VGND.n1227 VGND.n1225 0.110872
R6528 VGND.n1237 VGND.n1236 0.110872
R6529 VGND.n1232 VGND.n1231 0.110872
R6530 VGND.n1275 VGND.n1274 0.110872
R6531 VGND.n1281 VGND.n1280 0.110872
R6532 VGND.n928 VGND.n927 0.110872
R6533 VGND.n987 VGND.n986 0.110872
R6534 VGND.n982 VGND.n981 0.110872
R6535 VGND.n977 VGND.n976 0.110872
R6536 VGND.n972 VGND.n971 0.110872
R6537 VGND.n967 VGND.n966 0.110872
R6538 VGND.n962 VGND.n961 0.110872
R6539 VGND.n957 VGND.n956 0.110872
R6540 VGND.n952 VGND.n951 0.110872
R6541 VGND.n947 VGND.n946 0.110872
R6542 VGND.n942 VGND.n941 0.110872
R6543 VGND.n937 VGND.n936 0.110872
R6544 VGND.n932 VGND.n931 0.110872
R6545 VGND.n895 VGND.n894 0.110872
R6546 VGND.n1333 VGND.n1332 0.110872
R6547 VGND.n1130 VGND 0.0981562
R6548 VGND.n2214 VGND 0.0981562
R6549 VGND.n1362 VGND 0.0981562
R6550 VGND.n19 VGND 0.0968542
R6551 VGND.n2952 VGND 0.0968542
R6552 VGND.n45 VGND 0.0968542
R6553 VGND VGND.n91 0.0968542
R6554 VGND VGND.n130 0.0968542
R6555 VGND VGND.n499 0.0968542
R6556 VGND VGND.n2280 0.0968542
R6557 VGND VGND.n535 0.0968542
R6558 VGND VGND.n2207 0.0968542
R6559 VGND.n2224 VGND 0.0968542
R6560 VGND.n2982 VGND 0.0968542
R6561 VGND.n2562 VGND 0.088625
R6562 VGND.n2633 VGND 0.0790114
R6563 VGND.n2695 VGND 0.0790114
R6564 VGND.n2690 VGND 0.0790114
R6565 VGND VGND.n2689 0.0790114
R6566 VGND.n2684 VGND 0.0790114
R6567 VGND VGND.n2683 0.0790114
R6568 VGND.n2678 VGND 0.0790114
R6569 VGND VGND.n2677 0.0790114
R6570 VGND.n2709 VGND 0.0790114
R6571 VGND.n2723 VGND 0.0790114
R6572 VGND.n2742 VGND 0.0790114
R6573 VGND.n2761 VGND 0.0790114
R6574 VGND.n2781 VGND 0.0790114
R6575 VGND VGND.n2780 0.0790114
R6576 VGND VGND.n284 0.0790114
R6577 VGND.n2940 VGND 0.0790114
R6578 VGND.n2635 VGND 0.0790114
R6579 VGND.n2693 VGND 0.0790114
R6580 VGND VGND.n2692 0.0790114
R6581 VGND.n2687 VGND 0.0790114
R6582 VGND VGND.n2686 0.0790114
R6583 VGND.n2681 VGND 0.0790114
R6584 VGND VGND.n2680 0.0790114
R6585 VGND.n2675 VGND 0.0790114
R6586 VGND.n2711 VGND 0.0790114
R6587 VGND.n2721 VGND 0.0790114
R6588 VGND.n2744 VGND 0.0790114
R6589 VGND.n2759 VGND 0.0790114
R6590 VGND.n2783 VGND 0.0790114
R6591 VGND.n2784 VGND 0.0790114
R6592 VGND.n2794 VGND 0.0790114
R6593 VGND.n2937 VGND 0.0790114
R6594 VGND VGND.n2559 0.0790114
R6595 VGND VGND.n2558 0.0790114
R6596 VGND VGND.n2557 0.0790114
R6597 VGND VGND.n2556 0.0790114
R6598 VGND VGND.n2555 0.0790114
R6599 VGND VGND.n2554 0.0790114
R6600 VGND VGND.n2553 0.0790114
R6601 VGND VGND.n2552 0.0790114
R6602 VGND VGND.n2551 0.0790114
R6603 VGND VGND.n2550 0.0790114
R6604 VGND VGND.n2549 0.0790114
R6605 VGND VGND.n2548 0.0790114
R6606 VGND VGND.n2547 0.0790114
R6607 VGND.n2798 VGND 0.0790114
R6608 VGND VGND.n2797 0.0790114
R6609 VGND.n2533 VGND 0.0790114
R6610 VGND.n2357 VGND 0.0790114
R6611 VGND.n2373 VGND 0.0790114
R6612 VGND.n2383 VGND 0.0790114
R6613 VGND.n2399 VGND 0.0790114
R6614 VGND.n2409 VGND 0.0790114
R6615 VGND.n2425 VGND 0.0790114
R6616 VGND.n2435 VGND 0.0790114
R6617 VGND.n2451 VGND 0.0790114
R6618 VGND.n2461 VGND 0.0790114
R6619 VGND.n2477 VGND 0.0790114
R6620 VGND.n2487 VGND 0.0790114
R6621 VGND.n2508 VGND 0.0790114
R6622 VGND.n2802 VGND 0.0790114
R6623 VGND VGND.n2801 0.0790114
R6624 VGND.n419 VGND 0.0790114
R6625 VGND.n2530 VGND 0.0790114
R6626 VGND.n2360 VGND 0.0790114
R6627 VGND.n2370 VGND 0.0790114
R6628 VGND.n2386 VGND 0.0790114
R6629 VGND.n2396 VGND 0.0790114
R6630 VGND.n2412 VGND 0.0790114
R6631 VGND.n2422 VGND 0.0790114
R6632 VGND.n2438 VGND 0.0790114
R6633 VGND.n2448 VGND 0.0790114
R6634 VGND.n2464 VGND 0.0790114
R6635 VGND.n2474 VGND 0.0790114
R6636 VGND.n2490 VGND 0.0790114
R6637 VGND.n2505 VGND 0.0790114
R6638 VGND.n2805 VGND 0.0790114
R6639 VGND.n2806 VGND 0.0790114
R6640 VGND.n2819 VGND 0.0790114
R6641 VGND VGND.n2818 0.0790114
R6642 VGND.n1907 VGND 0.0790114
R6643 VGND.n1917 VGND 0.0790114
R6644 VGND.n1918 VGND 0.0790114
R6645 VGND.n1928 VGND 0.0790114
R6646 VGND.n1929 VGND 0.0790114
R6647 VGND.n1939 VGND 0.0790114
R6648 VGND.n1940 VGND 0.0790114
R6649 VGND.n1950 VGND 0.0790114
R6650 VGND.n1951 VGND 0.0790114
R6651 VGND.n1961 VGND 0.0790114
R6652 VGND.n1962 VGND 0.0790114
R6653 VGND.n1972 VGND 0.0790114
R6654 VGND.n1973 VGND 0.0790114
R6655 VGND.n2823 VGND 0.0790114
R6656 VGND VGND.n2822 0.0790114
R6657 VGND.n1990 VGND 0.0790114
R6658 VGND.n2063 VGND 0.0790114
R6659 VGND VGND.n2062 0.0790114
R6660 VGND.n2167 VGND 0.0790114
R6661 VGND VGND.n2166 0.0790114
R6662 VGND.n2159 VGND 0.0790114
R6663 VGND VGND.n2158 0.0790114
R6664 VGND.n2151 VGND 0.0790114
R6665 VGND VGND.n2150 0.0790114
R6666 VGND.n2143 VGND 0.0790114
R6667 VGND VGND.n2142 0.0790114
R6668 VGND.n2135 VGND 0.0790114
R6669 VGND VGND.n2134 0.0790114
R6670 VGND.n2827 VGND 0.0790114
R6671 VGND VGND.n2826 0.0790114
R6672 VGND.n1998 VGND 0.0790114
R6673 VGND VGND.n1997 0.0790114
R6674 VGND.n2066 VGND 0.0790114
R6675 VGND.n2171 VGND 0.0790114
R6676 VGND VGND.n2170 0.0790114
R6677 VGND.n2163 VGND 0.0790114
R6678 VGND VGND.n2162 0.0790114
R6679 VGND.n2155 VGND 0.0790114
R6680 VGND VGND.n2154 0.0790114
R6681 VGND.n2147 VGND 0.0790114
R6682 VGND VGND.n2146 0.0790114
R6683 VGND.n2139 VGND 0.0790114
R6684 VGND VGND.n2138 0.0790114
R6685 VGND.n2131 VGND 0.0790114
R6686 VGND.n2830 VGND 0.0790114
R6687 VGND.n2831 VGND 0.0790114
R6688 VGND.n2844 VGND 0.0790114
R6689 VGND VGND.n2843 0.0790114
R6690 VGND VGND.n1901 0.0790114
R6691 VGND.n2174 VGND 0.0790114
R6692 VGND.n1758 VGND 0.0790114
R6693 VGND.n1768 VGND 0.0790114
R6694 VGND.n1769 VGND 0.0790114
R6695 VGND.n1779 VGND 0.0790114
R6696 VGND.n1780 VGND 0.0790114
R6697 VGND.n1790 VGND 0.0790114
R6698 VGND.n1791 VGND 0.0790114
R6699 VGND.n1801 VGND 0.0790114
R6700 VGND.n1802 VGND 0.0790114
R6701 VGND.n1812 VGND 0.0790114
R6702 VGND.n1813 VGND 0.0790114
R6703 VGND.n2848 VGND 0.0790114
R6704 VGND VGND.n2847 0.0790114
R6705 VGND.n1830 VGND 0.0790114
R6706 VGND VGND.n1899 0.0790114
R6707 VGND.n1685 VGND 0.0790114
R6708 VGND.n1686 VGND 0.0790114
R6709 VGND.n1884 VGND 0.0790114
R6710 VGND VGND.n1883 0.0790114
R6711 VGND.n1876 VGND 0.0790114
R6712 VGND VGND.n1875 0.0790114
R6713 VGND.n1868 VGND 0.0790114
R6714 VGND VGND.n1867 0.0790114
R6715 VGND.n1860 VGND 0.0790114
R6716 VGND VGND.n1859 0.0790114
R6717 VGND.n1852 VGND 0.0790114
R6718 VGND.n2852 VGND 0.0790114
R6719 VGND VGND.n2851 0.0790114
R6720 VGND.n1838 VGND 0.0790114
R6721 VGND VGND.n1837 0.0790114
R6722 VGND.n1896 VGND 0.0790114
R6723 VGND VGND.n1895 0.0790114
R6724 VGND.n1888 VGND 0.0790114
R6725 VGND VGND.n1887 0.0790114
R6726 VGND.n1880 VGND 0.0790114
R6727 VGND VGND.n1879 0.0790114
R6728 VGND.n1872 VGND 0.0790114
R6729 VGND VGND.n1871 0.0790114
R6730 VGND.n1864 VGND 0.0790114
R6731 VGND VGND.n1863 0.0790114
R6732 VGND.n1856 VGND 0.0790114
R6733 VGND VGND.n1855 0.0790114
R6734 VGND.n2855 VGND 0.0790114
R6735 VGND.n2856 VGND 0.0790114
R6736 VGND.n2869 VGND 0.0790114
R6737 VGND VGND.n2868 0.0790114
R6738 VGND.n1349 VGND 0.0790114
R6739 VGND.n1892 VGND 0.0790114
R6740 VGND VGND.n1891 0.0790114
R6741 VGND.n867 VGND 0.0790114
R6742 VGND VGND.n866 0.0790114
R6743 VGND VGND.n865 0.0790114
R6744 VGND VGND.n864 0.0790114
R6745 VGND VGND.n863 0.0790114
R6746 VGND VGND.n862 0.0790114
R6747 VGND VGND.n861 0.0790114
R6748 VGND VGND.n860 0.0790114
R6749 VGND.n1669 VGND 0.0790114
R6750 VGND VGND.n1668 0.0790114
R6751 VGND.n2873 VGND 0.0790114
R6752 VGND VGND.n2872 0.0790114
R6753 VGND.n1654 VGND 0.0790114
R6754 VGND.n1404 VGND 0.0790114
R6755 VGND VGND.n1403 0.0790114
R6756 VGND VGND.n1402 0.0790114
R6757 VGND.n1487 VGND 0.0790114
R6758 VGND.n1497 VGND 0.0790114
R6759 VGND.n1513 VGND 0.0790114
R6760 VGND.n1523 VGND 0.0790114
R6761 VGND.n1539 VGND 0.0790114
R6762 VGND.n1560 VGND 0.0790114
R6763 VGND VGND.n1559 0.0790114
R6764 VGND.n1628 VGND 0.0790114
R6765 VGND.n1629 VGND 0.0790114
R6766 VGND.n2877 VGND 0.0790114
R6767 VGND VGND.n2876 0.0790114
R6768 VGND.n740 VGND 0.0790114
R6769 VGND.n1651 VGND 0.0790114
R6770 VGND.n1407 VGND 0.0790114
R6771 VGND.n1417 VGND 0.0790114
R6772 VGND.n1474 VGND 0.0790114
R6773 VGND.n1484 VGND 0.0790114
R6774 VGND.n1500 VGND 0.0790114
R6775 VGND.n1510 VGND 0.0790114
R6776 VGND.n1526 VGND 0.0790114
R6777 VGND.n1536 VGND 0.0790114
R6778 VGND.n1563 VGND 0.0790114
R6779 VGND.n1588 VGND 0.0790114
R6780 VGND.n1625 VGND 0.0790114
R6781 VGND VGND.n1624 0.0790114
R6782 VGND.n2880 VGND 0.0790114
R6783 VGND.n2881 VGND 0.0790114
R6784 VGND.n2894 VGND 0.0790114
R6785 VGND VGND.n2893 0.0790114
R6786 VGND VGND.n1344 0.0790114
R6787 VGND.n1420 VGND 0.0790114
R6788 VGND.n1471 VGND 0.0790114
R6789 VGND VGND.n1470 0.0790114
R6790 VGND VGND.n1469 0.0790114
R6791 VGND VGND.n1468 0.0790114
R6792 VGND VGND.n1467 0.0790114
R6793 VGND VGND.n1466 0.0790114
R6794 VGND VGND.n1465 0.0790114
R6795 VGND.n1591 VGND 0.0790114
R6796 VGND.n1592 VGND 0.0790114
R6797 VGND.n1621 VGND 0.0790114
R6798 VGND VGND.n1620 0.0790114
R6799 VGND.n2898 VGND 0.0790114
R6800 VGND VGND.n2897 0.0790114
R6801 VGND.n1606 VGND 0.0790114
R6802 VGND.n1103 VGND 0.0790114
R6803 VGND VGND.n1102 0.0790114
R6804 VGND VGND.n1101 0.0790114
R6805 VGND.n1321 VGND 0.0790114
R6806 VGND VGND.n1320 0.0790114
R6807 VGND.n1313 VGND 0.0790114
R6808 VGND VGND.n1312 0.0790114
R6809 VGND.n1305 VGND 0.0790114
R6810 VGND VGND.n1304 0.0790114
R6811 VGND.n1067 VGND 0.0790114
R6812 VGND VGND.n1066 0.0790114
R6813 VGND VGND.n1065 0.0790114
R6814 VGND VGND.n1064 0.0790114
R6815 VGND.n2901 VGND 0.0790114
R6816 VGND.n233 VGND 0.0790114
R6817 VGND.n2913 VGND 0.0790114
R6818 VGND.n1163 VGND 0.0790114
R6819 VGND.n1328 VGND 0.0790114
R6820 VGND VGND.n1327 0.0790114
R6821 VGND.n898 VGND 0.0790114
R6822 VGND.n901 VGND 0.0790114
R6823 VGND.n904 VGND 0.0790114
R6824 VGND.n907 VGND 0.0790114
R6825 VGND.n910 VGND 0.0790114
R6826 VGND.n913 VGND 0.0790114
R6827 VGND.n1298 VGND 0.0790114
R6828 VGND VGND.n1297 0.0790114
R6829 VGND.n1292 VGND 0.0790114
R6830 VGND VGND.n1291 0.0790114
R6831 VGND.n1270 VGND 0.0790114
R6832 VGND.n1285 VGND 0.0790114
R6833 VGND VGND.n1284 0.0790114
R6834 VGND.n1161 VGND 0.0790114
R6835 VGND.n1330 VGND 0.0790114
R6836 VGND.n1325 VGND 0.0790114
R6837 VGND VGND.n1324 0.0790114
R6838 VGND.n1317 VGND 0.0790114
R6839 VGND VGND.n1316 0.0790114
R6840 VGND.n1309 VGND 0.0790114
R6841 VGND VGND.n1308 0.0790114
R6842 VGND.n1301 VGND 0.0790114
R6843 VGND VGND.n1300 0.0790114
R6844 VGND.n1295 VGND 0.0790114
R6845 VGND VGND.n1294 0.0790114
R6846 VGND.n1289 VGND 0.0790114
R6847 VGND VGND.n1288 0.0790114
R6848 VGND VGND.n1287 0.0790114
R6849 VGND.n2916 VGND 0.0790114
R6850 VGND.n2699 VGND.n2698 0.0656596
R6851 VGND.n357 VGND.n355 0.0656596
R6852 VGND.n364 VGND.n362 0.0656596
R6853 VGND.n368 VGND.n367 0.0656596
R6854 VGND.n375 VGND.n373 0.0656596
R6855 VGND.n379 VGND.n378 0.0656596
R6856 VGND.n386 VGND.n384 0.0656596
R6857 VGND.n387 VGND.n325 0.0656596
R6858 VGND.n326 VGND.n314 0.0656596
R6859 VGND.n2726 VGND.n309 0.0656596
R6860 VGND.n312 VGND.n311 0.0656596
R6861 VGND.n2735 VGND.n2734 0.0656596
R6862 VGND.n2730 VGND.n293 0.0656596
R6863 VGND.n296 VGND.n294 0.0656596
R6864 VGND.n2773 VGND.n203 0.0656596
R6865 VGND.n2606 VGND 0.063
R6866 VGND.n2603 VGND 0.063
R6867 VGND.n2600 VGND 0.063
R6868 VGND.n2597 VGND 0.063
R6869 VGND.n2594 VGND 0.063
R6870 VGND.n2591 VGND 0.063
R6871 VGND.n2588 VGND 0.063
R6872 VGND.n2585 VGND 0.063
R6873 VGND.n2582 VGND 0.063
R6874 VGND.n2579 VGND 0.063
R6875 VGND.n2576 VGND 0.063
R6876 VGND.n2573 VGND 0.063
R6877 VGND.n2570 VGND 0.063
R6878 VGND.n2567 VGND 0.063
R6879 VGND.n2564 VGND 0.063
R6880 VGND VGND.n31 0.0603958
R6881 VGND.n3009 VGND 0.0603958
R6882 VGND VGND.n3008 0.0603958
R6883 VGND.n192 VGND 0.0603958
R6884 VGND VGND.n191 0.0603958
R6885 VGND VGND.n2964 0.0603958
R6886 VGND.n2965 VGND 0.0603958
R6887 VGND VGND.n57 0.0603958
R6888 VGND.n64 VGND 0.0603958
R6889 VGND VGND.n63 0.0603958
R6890 VGND.n118 VGND 0.0603958
R6891 VGND.n119 VGND 0.0603958
R6892 VGND.n132 VGND 0.0603958
R6893 VGND VGND.n131 0.0603958
R6894 VGND.n127 VGND 0.0603958
R6895 VGND.n163 VGND 0.0603958
R6896 VGND VGND.n162 0.0603958
R6897 VGND.n1152 VGND 0.0603958
R6898 VGND.n1129 VGND 0.0603958
R6899 VGND VGND.n1128 0.0603958
R6900 VGND.n1125 VGND 0.0603958
R6901 VGND.n501 VGND 0.0603958
R6902 VGND VGND.n500 0.0603958
R6903 VGND.n483 VGND 0.0603958
R6904 VGND.n2282 VGND 0.0603958
R6905 VGND VGND.n2281 0.0603958
R6906 VGND.n2264 VGND 0.0603958
R6907 VGND.n537 VGND 0.0603958
R6908 VGND VGND.n536 0.0603958
R6909 VGND.n519 VGND 0.0603958
R6910 VGND.n2209 VGND 0.0603958
R6911 VGND VGND.n2208 0.0603958
R6912 VGND.n2201 VGND 0.0603958
R6913 VGND.n2198 VGND 0.0603958
R6914 VGND.n2193 VGND 0.0603958
R6915 VGND VGND.n2225 0.0603958
R6916 VGND.n2246 VGND 0.0603958
R6917 VGND VGND.n2245 0.0603958
R6918 VGND VGND.n1363 0.0603958
R6919 VGND.n1384 VGND 0.0603958
R6920 VGND VGND.n1383 0.0603958
R6921 VGND VGND.n2994 0.0603958
R6922 VGND.n2995 VGND 0.0603958
R6923 VGND.n2996 VGND 0.0603958
R6924 VGND.n2698 VGND 0.0574853
R6925 VGND.n357 VGND 0.0574853
R6926 VGND.n364 VGND 0.0574853
R6927 VGND.n367 VGND 0.0574853
R6928 VGND.n375 VGND 0.0574853
R6929 VGND.n378 VGND 0.0574853
R6930 VGND.n386 VGND 0.0574853
R6931 VGND.n325 VGND 0.0574853
R6932 VGND.n314 VGND 0.0574853
R6933 VGND.n309 VGND 0.0574853
R6934 VGND.n311 VGND 0.0574853
R6935 VGND.n2734 VGND 0.0574853
R6936 VGND.n293 VGND 0.0574853
R6937 VGND.n296 VGND 0.0574853
R6938 VGND.n203 VGND 0.0574853
R6939 VGND.n1021 VGND 0.0489375
R6940 VGND.n994 VGND 0.0489375
R6941 VGND.n2630 VGND 0.0489375
R6942 VGND.n204 VGND 0.0489375
R6943 VGND.n334 VGND 0.0489375
R6944 VGND.n2626 VGND 0.0489375
R6945 VGND.n2623 VGND 0.0489375
R6946 VGND.n2620 VGND 0.0489375
R6947 VGND.n2617 VGND 0.0489375
R6948 VGND.n2614 VGND 0.0489375
R6949 VGND.n2611 VGND 0.0489375
R6950 VGND.n322 VGND 0.0489375
R6951 VGND.n315 VGND 0.0489375
R6952 VGND.n306 VGND 0.0489375
R6953 VGND.n299 VGND 0.0489375
R6954 VGND.n2765 VGND 0.0489375
R6955 VGND.n290 VGND 0.0489375
R6956 VGND.n297 VGND 0.0489375
R6957 VGND.n1018 VGND 0.0489375
R6958 VGND.n1015 VGND 0.0489375
R6959 VGND.n1180 VGND 0.0489375
R6960 VGND.n1006 VGND 0.0489375
R6961 VGND.n1004 VGND 0.0489375
R6962 VGND.n1195 VGND 0.0489375
R6963 VGND.n1212 VGND 0.0489375
R6964 VGND.n1000 VGND 0.0489375
R6965 VGND.n1253 VGND 0.0489375
R6966 VGND.n1256 VGND 0.0489375
R6967 VGND.n1259 VGND 0.0489375
R6968 VGND.n1262 VGND 0.0489375
R6969 VGND.n998 VGND 0.0489375
R6970 VGND.n1265 VGND 0.0489375
R6971 VGND VGND.n330 0.037734
R6972 VGND.n286 VGND 0.037734
R6973 VGND.n2787 VGND 0.037734
R6974 VGND.n2752 VGND 0.037734
R6975 VGND.n303 VGND 0.037734
R6976 VGND.n2747 VGND 0.037734
R6977 VGND.n319 VGND 0.037734
R6978 VGND.n2714 VGND 0.037734
R6979 VGND.n393 VGND 0.037734
R6980 VGND.n2668 VGND 0.037734
R6981 VGND.n2663 VGND 0.037734
R6982 VGND.n2658 VGND 0.037734
R6983 VGND.n2653 VGND 0.037734
R6984 VGND.n2648 VGND 0.037734
R6985 VGND.n2643 VGND 0.037734
R6986 VGND.n2638 VGND 0.037734
R6987 VGND VGND.n396 0.037734
R6988 VGND.n2535 VGND 0.037734
R6989 VGND.n2540 VGND 0.037734
R6990 VGND.n414 VGND 0.037734
R6991 VGND.n2287 VGND 0.037734
R6992 VGND.n2292 VGND 0.037734
R6993 VGND.n2297 VGND 0.037734
R6994 VGND.n2302 VGND 0.037734
R6995 VGND.n2307 VGND 0.037734
R6996 VGND.n2312 VGND 0.037734
R6997 VGND.n2317 VGND 0.037734
R6998 VGND.n2322 VGND 0.037734
R6999 VGND.n2327 VGND 0.037734
R7000 VGND.n2332 VGND 0.037734
R7001 VGND.n2337 VGND 0.037734
R7002 VGND.n2342 VGND 0.037734
R7003 VGND VGND.n400 0.037734
R7004 VGND VGND.n2528 0.037734
R7005 VGND.n2521 VGND 0.037734
R7006 VGND.n2516 VGND 0.037734
R7007 VGND.n2511 VGND 0.037734
R7008 VGND.n427 VGND 0.037734
R7009 VGND.n2480 VGND 0.037734
R7010 VGND.n435 VGND 0.037734
R7011 VGND.n2454 VGND 0.037734
R7012 VGND.n443 VGND 0.037734
R7013 VGND.n2428 VGND 0.037734
R7014 VGND.n451 VGND 0.037734
R7015 VGND.n2402 VGND 0.037734
R7016 VGND.n459 VGND 0.037734
R7017 VGND.n2376 VGND 0.037734
R7018 VGND.n471 VGND 0.037734
R7019 VGND VGND.n469 0.037734
R7020 VGND VGND.n2816 0.037734
R7021 VGND.n2809 VGND 0.037734
R7022 VGND.n2498 VGND 0.037734
R7023 VGND.n423 VGND 0.037734
R7024 VGND.n2493 VGND 0.037734
R7025 VGND.n431 VGND 0.037734
R7026 VGND.n2467 VGND 0.037734
R7027 VGND.n439 VGND 0.037734
R7028 VGND.n2441 VGND 0.037734
R7029 VGND.n447 VGND 0.037734
R7030 VGND.n2415 VGND 0.037734
R7031 VGND.n455 VGND 0.037734
R7032 VGND.n2389 VGND 0.037734
R7033 VGND.n463 VGND 0.037734
R7034 VGND.n2363 VGND 0.037734
R7035 VGND VGND.n466 0.037734
R7036 VGND VGND.n1988 0.037734
R7037 VGND.n1981 VGND 0.037734
R7038 VGND.n1976 VGND 0.037734
R7039 VGND.n607 VGND 0.037734
R7040 VGND.n1965 VGND 0.037734
R7041 VGND.n610 VGND 0.037734
R7042 VGND.n1954 VGND 0.037734
R7043 VGND.n613 VGND 0.037734
R7044 VGND.n1943 VGND 0.037734
R7045 VGND.n616 VGND 0.037734
R7046 VGND.n1932 VGND 0.037734
R7047 VGND.n619 VGND 0.037734
R7048 VGND.n1921 VGND 0.037734
R7049 VGND.n622 VGND 0.037734
R7050 VGND.n1910 VGND 0.037734
R7051 VGND VGND.n625 0.037734
R7052 VGND VGND.n1995 0.037734
R7053 VGND.n2000 VGND 0.037734
R7054 VGND.n2005 VGND 0.037734
R7055 VGND.n2010 VGND 0.037734
R7056 VGND.n2015 VGND 0.037734
R7057 VGND.n2020 VGND 0.037734
R7058 VGND.n2025 VGND 0.037734
R7059 VGND.n2030 VGND 0.037734
R7060 VGND.n2035 VGND 0.037734
R7061 VGND.n2040 VGND 0.037734
R7062 VGND.n2045 VGND 0.037734
R7063 VGND.n2050 VGND 0.037734
R7064 VGND.n2055 VGND 0.037734
R7065 VGND.n593 VGND 0.037734
R7066 VGND.n596 VGND 0.037734
R7067 VGND VGND.n590 0.037734
R7068 VGND VGND.n2841 0.037734
R7069 VGND.n2834 VGND 0.037734
R7070 VGND.n2124 VGND 0.037734
R7071 VGND.n584 VGND 0.037734
R7072 VGND.n2119 VGND 0.037734
R7073 VGND.n2114 VGND 0.037734
R7074 VGND.n2109 VGND 0.037734
R7075 VGND.n2104 VGND 0.037734
R7076 VGND.n2099 VGND 0.037734
R7077 VGND.n2094 VGND 0.037734
R7078 VGND.n2089 VGND 0.037734
R7079 VGND.n2084 VGND 0.037734
R7080 VGND.n2079 VGND 0.037734
R7081 VGND.n2074 VGND 0.037734
R7082 VGND.n2069 VGND 0.037734
R7083 VGND VGND.n587 0.037734
R7084 VGND VGND.n1828 0.037734
R7085 VGND.n1821 VGND 0.037734
R7086 VGND.n1816 VGND 0.037734
R7087 VGND.n1740 VGND 0.037734
R7088 VGND.n1805 VGND 0.037734
R7089 VGND.n1743 VGND 0.037734
R7090 VGND.n1794 VGND 0.037734
R7091 VGND.n1746 VGND 0.037734
R7092 VGND.n1783 VGND 0.037734
R7093 VGND.n1749 VGND 0.037734
R7094 VGND.n1772 VGND 0.037734
R7095 VGND.n1752 VGND 0.037734
R7096 VGND.n1761 VGND 0.037734
R7097 VGND VGND.n1757 0.037734
R7098 VGND.n2176 VGND 0.037734
R7099 VGND VGND.n547 0.037734
R7100 VGND VGND.n1835 0.037734
R7101 VGND.n1840 VGND 0.037734
R7102 VGND.n1845 VGND 0.037734
R7103 VGND.n1672 VGND 0.037734
R7104 VGND.n1729 VGND 0.037734
R7105 VGND.n1724 VGND 0.037734
R7106 VGND.n1719 VGND 0.037734
R7107 VGND.n1714 VGND 0.037734
R7108 VGND.n1709 VGND 0.037734
R7109 VGND.n1704 VGND 0.037734
R7110 VGND.n1699 VGND 0.037734
R7111 VGND.n1694 VGND 0.037734
R7112 VGND.n1689 VGND 0.037734
R7113 VGND.n1675 VGND 0.037734
R7114 VGND.n1678 VGND 0.037734
R7115 VGND VGND.n628 0.037734
R7116 VGND VGND.n2866 0.037734
R7117 VGND.n2859 VGND 0.037734
R7118 VGND.n724 VGND 0.037734
R7119 VGND.n666 VGND 0.037734
R7120 VGND.n719 VGND 0.037734
R7121 VGND.n714 VGND 0.037734
R7122 VGND.n709 VGND 0.037734
R7123 VGND.n704 VGND 0.037734
R7124 VGND.n699 VGND 0.037734
R7125 VGND.n694 VGND 0.037734
R7126 VGND.n689 VGND 0.037734
R7127 VGND.n684 VGND 0.037734
R7128 VGND.n679 VGND 0.037734
R7129 VGND.n674 VGND 0.037734
R7130 VGND.n669 VGND 0.037734
R7131 VGND VGND.n632 0.037734
R7132 VGND.n1656 VGND 0.037734
R7133 VGND.n1661 VGND 0.037734
R7134 VGND.n734 VGND 0.037734
R7135 VGND.n853 VGND 0.037734
R7136 VGND.n819 VGND 0.037734
R7137 VGND.n848 VGND 0.037734
R7138 VGND.n843 VGND 0.037734
R7139 VGND.n838 VGND 0.037734
R7140 VGND.n833 VGND 0.037734
R7141 VGND.n828 VGND 0.037734
R7142 VGND.n823 VGND 0.037734
R7143 VGND VGND.n811 0.037734
R7144 VGND.n869 VGND 0.037734
R7145 VGND.n874 VGND 0.037734
R7146 VGND.n1352 VGND 0.037734
R7147 VGND VGND.n879 0.037734
R7148 VGND VGND.n1649 0.037734
R7149 VGND.n1642 VGND 0.037734
R7150 VGND.n1637 VGND 0.037734
R7151 VGND.n1632 VGND 0.037734
R7152 VGND.n1552 VGND 0.037734
R7153 VGND.n760 VGND 0.037734
R7154 VGND.n1547 VGND 0.037734
R7155 VGND.n1542 VGND 0.037734
R7156 VGND.n768 VGND 0.037734
R7157 VGND.n1516 VGND 0.037734
R7158 VGND.n776 VGND 0.037734
R7159 VGND.n1490 VGND 0.037734
R7160 VGND.n804 VGND 0.037734
R7161 VGND.n1395 VGND 0.037734
R7162 VGND.n1390 VGND 0.037734
R7163 VGND VGND.n800 0.037734
R7164 VGND VGND.n2891 0.037734
R7165 VGND.n2884 VGND 0.037734
R7166 VGND.n1571 VGND 0.037734
R7167 VGND.n1576 VGND 0.037734
R7168 VGND.n1581 VGND 0.037734
R7169 VGND.n755 VGND 0.037734
R7170 VGND.n1566 VGND 0.037734
R7171 VGND.n764 VGND 0.037734
R7172 VGND.n1529 VGND 0.037734
R7173 VGND.n772 VGND 0.037734
R7174 VGND.n1503 VGND 0.037734
R7175 VGND.n780 VGND 0.037734
R7176 VGND.n1477 VGND 0.037734
R7177 VGND.n794 VGND 0.037734
R7178 VGND.n1410 VGND 0.037734
R7179 VGND VGND.n797 0.037734
R7180 VGND.n1608 VGND 0.037734
R7181 VGND.n1613 VGND 0.037734
R7182 VGND.n749 VGND 0.037734
R7183 VGND.n1600 VGND 0.037734
R7184 VGND.n1595 VGND 0.037734
R7185 VGND.n1458 VGND 0.037734
R7186 VGND.n790 VGND 0.037734
R7187 VGND.n1453 VGND 0.037734
R7188 VGND.n1448 VGND 0.037734
R7189 VGND.n1443 VGND 0.037734
R7190 VGND.n1438 VGND 0.037734
R7191 VGND.n1433 VGND 0.037734
R7192 VGND.n1428 VGND 0.037734
R7193 VGND.n1423 VGND 0.037734
R7194 VGND.n884 VGND 0.037734
R7195 VGND VGND.n882 0.037734
R7196 VGND VGND.n2911 0.037734
R7197 VGND.n2904 VGND 0.037734
R7198 VGND.n1048 VGND 0.037734
R7199 VGND.n1057 VGND 0.037734
R7200 VGND.n1052 VGND 0.037734
R7201 VGND VGND.n1044 0.037734
R7202 VGND.n1069 VGND 0.037734
R7203 VGND.n1074 VGND 0.037734
R7204 VGND.n1079 VGND 0.037734
R7205 VGND.n1084 VGND 0.037734
R7206 VGND.n1089 VGND 0.037734
R7207 VGND.n1094 VGND 0.037734
R7208 VGND.n1028 VGND 0.037734
R7209 VGND.n1036 VGND 0.037734
R7210 VGND.n1031 VGND 0.037734
R7211 VGND VGND.n1024 0.037734
R7212 VGND VGND.n1014 0.037734
R7213 VGND VGND.n1169 0.037734
R7214 VGND.n1172 VGND 0.037734
R7215 VGND VGND.n1179 0.037734
R7216 VGND.n1185 VGND 0.037734
R7217 VGND.n1008 VGND 0.037734
R7218 VGND.n1204 VGND 0.037734
R7219 VGND VGND.n1211 0.037734
R7220 VGND.n1217 VGND 0.037734
R7221 VGND VGND.n1222 0.037734
R7222 VGND.n1243 VGND 0.037734
R7223 VGND VGND.n1227 0.037734
R7224 VGND.n1236 VGND 0.037734
R7225 VGND.n1231 VGND 0.037734
R7226 VGND.n1274 VGND 0.037734
R7227 VGND VGND.n1281 0.037734
R7228 VGND.n927 VGND 0.037734
R7229 VGND.n986 VGND 0.037734
R7230 VGND.n981 VGND 0.037734
R7231 VGND.n976 VGND 0.037734
R7232 VGND.n971 VGND 0.037734
R7233 VGND.n966 VGND 0.037734
R7234 VGND.n961 VGND 0.037734
R7235 VGND.n956 VGND 0.037734
R7236 VGND.n951 VGND 0.037734
R7237 VGND.n946 VGND 0.037734
R7238 VGND.n941 VGND 0.037734
R7239 VGND.n936 VGND 0.037734
R7240 VGND.n931 VGND 0.037734
R7241 VGND VGND.n895 0.037734
R7242 VGND.n1332 VGND 0.037734
R7243 VGND VGND.n887 0.037734
R7244 VGND.n1156 VGND 0.0343542
R7245 VGND.n1128 VGND 0.0343542
R7246 VGND.n501 VGND 0.0343542
R7247 VGND.n2282 VGND 0.0343542
R7248 VGND.n537 VGND 0.0343542
R7249 VGND.n2209 VGND 0.0343542
R7250 VGND.n2246 VGND 0.0343542
R7251 VGND.n1384 VGND 0.0343542
R7252 VGND.n3009 VGND 0.0330521
R7253 VGND.n192 VGND 0.0330521
R7254 VGND.n2965 VGND 0.0330521
R7255 VGND.n64 VGND 0.0330521
R7256 VGND VGND.n118 0.0330521
R7257 VGND.n132 VGND 0.0330521
R7258 VGND.n163 VGND 0.0330521
R7259 VGND VGND.n2995 0.0330521
R7260 VGND.n33 VGND 0.024
R7261 VGND.n1 VGND 0.024
R7262 VGND.n119 VGND 0.0239375
R7263 VGND.n131 VGND 0.0239375
R7264 VGND.n500 VGND 0.0239375
R7265 VGND.n2281 VGND 0.0239375
R7266 VGND.n536 VGND 0.0239375
R7267 VGND.n3003 VGND 0.0226354
R7268 VGND VGND.n124 0.0226354
R7269 VGND.n1133 VGND 0.0226354
R7270 VGND VGND.n2256 0.0226354
R7271 VGND.n2217 VGND 0.0226354
R7272 VGND.n2208 VGND 0.0226354
R7273 VGND.n2220 VGND 0.0226354
R7274 VGND VGND.n3000 0.0226354
R7275 VGND VGND.n189 0.0213333
R7276 VGND.n191 VGND 0.0213333
R7277 VGND.n58 VGND 0.0213333
R7278 VGND.n113 VGND 0.0213333
R7279 VGND VGND.n90 0.0213333
R7280 VGND VGND.n158 0.0213333
R7281 VGND.n162 VGND 0.0213333
R7282 VGND VGND.n511 0.0213333
R7283 VGND.n2213 VGND 0.0213333
R7284 VGND.n1358 VGND 0.0213333
R7285 VGND VGND.n3024 0.0193356
R7286 VGND.n33 VGND 0.0161667
R7287 VGND.n331 VGND 0.00980851
R7288 VGND.n2936 VGND 0.00980851
R7289 VGND.n2793 VGND 0.00980851
R7290 VGND.n2785 VGND 0.00980851
R7291 VGND VGND.n288 0.00980851
R7292 VGND.n2758 VGND 0.00980851
R7293 VGND.n2745 VGND 0.00980851
R7294 VGND.n2720 VGND 0.00980851
R7295 VGND.n2712 VGND 0.00980851
R7296 VGND.n2674 VGND 0.00980851
R7297 VGND VGND.n350 0.00980851
R7298 VGND VGND.n349 0.00980851
R7299 VGND VGND.n344 0.00980851
R7300 VGND VGND.n343 0.00980851
R7301 VGND VGND.n338 0.00980851
R7302 VGND VGND.n337 0.00980851
R7303 VGND.n2636 VGND 0.00980851
R7304 VGND VGND.n2534 0.00980851
R7305 VGND VGND.n283 0.00980851
R7306 VGND VGND.n282 0.00980851
R7307 VGND.n2546 VGND 0.00980851
R7308 VGND VGND.n412 0.00980851
R7309 VGND VGND.n411 0.00980851
R7310 VGND VGND.n410 0.00980851
R7311 VGND VGND.n409 0.00980851
R7312 VGND VGND.n408 0.00980851
R7313 VGND VGND.n407 0.00980851
R7314 VGND VGND.n406 0.00980851
R7315 VGND VGND.n405 0.00980851
R7316 VGND VGND.n404 0.00980851
R7317 VGND VGND.n403 0.00980851
R7318 VGND VGND.n402 0.00980851
R7319 VGND.n401 VGND 0.00980851
R7320 VGND.n2529 VGND 0.00980851
R7321 VGND VGND.n420 0.00980851
R7322 VGND VGND.n280 0.00980851
R7323 VGND VGND.n279 0.00980851
R7324 VGND.n2509 VGND 0.00980851
R7325 VGND.n2486 VGND 0.00980851
R7326 VGND.n2478 VGND 0.00980851
R7327 VGND.n2460 VGND 0.00980851
R7328 VGND.n2452 VGND 0.00980851
R7329 VGND.n2434 VGND 0.00980851
R7330 VGND.n2426 VGND 0.00980851
R7331 VGND.n2408 VGND 0.00980851
R7332 VGND.n2400 VGND 0.00980851
R7333 VGND.n2382 VGND 0.00980851
R7334 VGND.n2374 VGND 0.00980851
R7335 VGND.n2356 VGND 0.00980851
R7336 VGND.n2817 VGND 0.00980851
R7337 VGND VGND.n273 0.00980851
R7338 VGND.n2807 VGND 0.00980851
R7339 VGND VGND.n277 0.00980851
R7340 VGND.n2504 VGND 0.00980851
R7341 VGND.n2491 VGND 0.00980851
R7342 VGND.n2473 VGND 0.00980851
R7343 VGND.n2465 VGND 0.00980851
R7344 VGND.n2447 VGND 0.00980851
R7345 VGND.n2439 VGND 0.00980851
R7346 VGND.n2421 VGND 0.00980851
R7347 VGND.n2413 VGND 0.00980851
R7348 VGND.n2395 VGND 0.00980851
R7349 VGND.n2387 VGND 0.00980851
R7350 VGND.n2369 VGND 0.00980851
R7351 VGND.n2361 VGND 0.00980851
R7352 VGND.n1989 VGND 0.00980851
R7353 VGND VGND.n271 0.00980851
R7354 VGND VGND.n270 0.00980851
R7355 VGND.n1974 VGND 0.00980851
R7356 VGND.n1971 VGND 0.00980851
R7357 VGND.n1963 VGND 0.00980851
R7358 VGND.n1960 VGND 0.00980851
R7359 VGND.n1952 VGND 0.00980851
R7360 VGND.n1949 VGND 0.00980851
R7361 VGND.n1941 VGND 0.00980851
R7362 VGND.n1938 VGND 0.00980851
R7363 VGND.n1930 VGND 0.00980851
R7364 VGND.n1927 VGND 0.00980851
R7365 VGND.n1919 VGND 0.00980851
R7366 VGND.n1916 VGND 0.00980851
R7367 VGND.n1908 VGND 0.00980851
R7368 VGND.n1996 VGND 0.00980851
R7369 VGND VGND.n1999 0.00980851
R7370 VGND VGND.n268 0.00980851
R7371 VGND VGND.n267 0.00980851
R7372 VGND VGND.n581 0.00980851
R7373 VGND VGND.n580 0.00980851
R7374 VGND VGND.n575 0.00980851
R7375 VGND VGND.n574 0.00980851
R7376 VGND VGND.n569 0.00980851
R7377 VGND VGND.n568 0.00980851
R7378 VGND VGND.n563 0.00980851
R7379 VGND VGND.n562 0.00980851
R7380 VGND VGND.n557 0.00980851
R7381 VGND VGND.n556 0.00980851
R7382 VGND.n2061 VGND 0.00980851
R7383 VGND.n591 VGND 0.00980851
R7384 VGND.n2842 VGND 0.00980851
R7385 VGND VGND.n261 0.00980851
R7386 VGND.n2832 VGND 0.00980851
R7387 VGND VGND.n265 0.00980851
R7388 VGND.n2130 VGND 0.00980851
R7389 VGND VGND.n578 0.00980851
R7390 VGND VGND.n577 0.00980851
R7391 VGND VGND.n572 0.00980851
R7392 VGND VGND.n571 0.00980851
R7393 VGND VGND.n566 0.00980851
R7394 VGND VGND.n565 0.00980851
R7395 VGND VGND.n560 0.00980851
R7396 VGND VGND.n559 0.00980851
R7397 VGND VGND.n554 0.00980851
R7398 VGND VGND.n553 0.00980851
R7399 VGND.n2067 VGND 0.00980851
R7400 VGND.n1829 VGND 0.00980851
R7401 VGND VGND.n259 0.00980851
R7402 VGND VGND.n258 0.00980851
R7403 VGND.n1814 VGND 0.00980851
R7404 VGND.n1811 VGND 0.00980851
R7405 VGND.n1803 VGND 0.00980851
R7406 VGND.n1800 VGND 0.00980851
R7407 VGND.n1792 VGND 0.00980851
R7408 VGND.n1789 VGND 0.00980851
R7409 VGND.n1781 VGND 0.00980851
R7410 VGND.n1778 VGND 0.00980851
R7411 VGND.n1770 VGND 0.00980851
R7412 VGND.n1767 VGND 0.00980851
R7413 VGND.n1759 VGND 0.00980851
R7414 VGND VGND.n2175 0.00980851
R7415 VGND.n548 VGND 0.00980851
R7416 VGND.n1836 VGND 0.00980851
R7417 VGND VGND.n1839 0.00980851
R7418 VGND VGND.n256 0.00980851
R7419 VGND VGND.n255 0.00980851
R7420 VGND.n1851 VGND 0.00980851
R7421 VGND VGND.n662 0.00980851
R7422 VGND VGND.n661 0.00980851
R7423 VGND VGND.n656 0.00980851
R7424 VGND VGND.n655 0.00980851
R7425 VGND VGND.n650 0.00980851
R7426 VGND VGND.n649 0.00980851
R7427 VGND VGND.n644 0.00980851
R7428 VGND VGND.n643 0.00980851
R7429 VGND.n1687 VGND 0.00980851
R7430 VGND.n1684 VGND 0.00980851
R7431 VGND.n629 VGND 0.00980851
R7432 VGND.n2867 VGND 0.00980851
R7433 VGND VGND.n249 0.00980851
R7434 VGND.n2857 VGND 0.00980851
R7435 VGND VGND.n253 0.00980851
R7436 VGND.n730 VGND 0.00980851
R7437 VGND VGND.n664 0.00980851
R7438 VGND VGND.n659 0.00980851
R7439 VGND VGND.n658 0.00980851
R7440 VGND VGND.n653 0.00980851
R7441 VGND VGND.n652 0.00980851
R7442 VGND VGND.n647 0.00980851
R7443 VGND VGND.n646 0.00980851
R7444 VGND VGND.n641 0.00980851
R7445 VGND VGND.n640 0.00980851
R7446 VGND VGND.n634 0.00980851
R7447 VGND.n633 VGND 0.00980851
R7448 VGND VGND.n1655 0.00980851
R7449 VGND VGND.n247 0.00980851
R7450 VGND VGND.n246 0.00980851
R7451 VGND.n1667 VGND 0.00980851
R7452 VGND VGND.n732 0.00980851
R7453 VGND.n859 VGND 0.00980851
R7454 VGND VGND.n817 0.00980851
R7455 VGND VGND.n816 0.00980851
R7456 VGND VGND.n815 0.00980851
R7457 VGND VGND.n814 0.00980851
R7458 VGND VGND.n813 0.00980851
R7459 VGND.n812 VGND 0.00980851
R7460 VGND VGND.n868 0.00980851
R7461 VGND VGND.n637 0.00980851
R7462 VGND VGND.n636 0.00980851
R7463 VGND.n1350 VGND 0.00980851
R7464 VGND.n1650 VGND 0.00980851
R7465 VGND VGND.n741 0.00980851
R7466 VGND VGND.n244 0.00980851
R7467 VGND VGND.n243 0.00980851
R7468 VGND.n1630 VGND 0.00980851
R7469 VGND VGND.n742 0.00980851
R7470 VGND.n1558 VGND 0.00980851
R7471 VGND VGND.n758 0.00980851
R7472 VGND.n1540 VGND 0.00980851
R7473 VGND.n1522 VGND 0.00980851
R7474 VGND.n1514 VGND 0.00980851
R7475 VGND.n1496 VGND 0.00980851
R7476 VGND.n1488 VGND 0.00980851
R7477 VGND.n1401 VGND 0.00980851
R7478 VGND VGND.n802 0.00980851
R7479 VGND.n801 VGND 0.00980851
R7480 VGND.n2892 VGND 0.00980851
R7481 VGND VGND.n236 0.00980851
R7482 VGND.n2882 VGND 0.00980851
R7483 VGND VGND.n240 0.00980851
R7484 VGND VGND.n745 0.00980851
R7485 VGND VGND.n744 0.00980851
R7486 VGND.n1587 VGND 0.00980851
R7487 VGND.n1564 VGND 0.00980851
R7488 VGND.n1535 VGND 0.00980851
R7489 VGND.n1527 VGND 0.00980851
R7490 VGND.n1509 VGND 0.00980851
R7491 VGND.n1501 VGND 0.00980851
R7492 VGND.n1483 VGND 0.00980851
R7493 VGND.n1475 VGND 0.00980851
R7494 VGND.n1416 VGND 0.00980851
R7495 VGND.n1408 VGND 0.00980851
R7496 VGND VGND.n1607 0.00980851
R7497 VGND VGND.n232 0.00980851
R7498 VGND VGND.n231 0.00980851
R7499 VGND.n1619 VGND 0.00980851
R7500 VGND VGND.n747 0.00980851
R7501 VGND.n1593 VGND 0.00980851
R7502 VGND VGND.n751 0.00980851
R7503 VGND.n1464 VGND 0.00980851
R7504 VGND VGND.n788 0.00980851
R7505 VGND VGND.n787 0.00980851
R7506 VGND VGND.n786 0.00980851
R7507 VGND VGND.n785 0.00980851
R7508 VGND VGND.n784 0.00980851
R7509 VGND VGND.n783 0.00980851
R7510 VGND.n1421 VGND 0.00980851
R7511 VGND.n1343 VGND 0.00980851
R7512 VGND.n2912 VGND 0.00980851
R7513 VGND VGND.n228 0.00980851
R7514 VGND.n2902 VGND 0.00980851
R7515 VGND.n1063 VGND 0.00980851
R7516 VGND VGND.n1046 0.00980851
R7517 VGND.n1045 VGND 0.00980851
R7518 VGND VGND.n1068 0.00980851
R7519 VGND VGND.n912 0.00980851
R7520 VGND VGND.n911 0.00980851
R7521 VGND VGND.n906 0.00980851
R7522 VGND VGND.n905 0.00980851
R7523 VGND VGND.n900 0.00980851
R7524 VGND VGND.n899 0.00980851
R7525 VGND.n1100 VGND 0.00980851
R7526 VGND VGND.n1026 0.00980851
R7527 VGND.n1025 VGND 0.00980851
R7528 VGND.n1165 VGND 0.00980851
R7529 VGND.n1170 VGND 0.00980851
R7530 VGND VGND.n1011 0.00980851
R7531 VGND.n1183 VGND 0.00980851
R7532 VGND.n1191 VGND 0.00980851
R7533 VGND.n1202 VGND 0.00980851
R7534 VGND VGND.n1003 0.00980851
R7535 VGND.n1215 VGND 0.00980851
R7536 VGND.n1249 VGND 0.00980851
R7537 VGND.n1223 VGND 0.00980851
R7538 VGND VGND.n1242 0.00980851
R7539 VGND.n1228 VGND 0.00980851
R7540 VGND VGND.n1235 0.00980851
R7541 VGND.n1272 VGND 0.00980851
R7542 VGND VGND.n997 0.00980851
R7543 VGND.n1282 VGND 0.00980851
R7544 VGND.n2917 VGND 0.00980851
R7545 VGND.n992 VGND 0.00980851
R7546 VGND VGND.n925 0.00980851
R7547 VGND VGND.n924 0.00980851
R7548 VGND VGND.n920 0.00980851
R7549 VGND VGND.n919 0.00980851
R7550 VGND VGND.n915 0.00980851
R7551 VGND VGND.n914 0.00980851
R7552 VGND VGND.n909 0.00980851
R7553 VGND VGND.n908 0.00980851
R7554 VGND VGND.n903 0.00980851
R7555 VGND VGND.n902 0.00980851
R7556 VGND VGND.n897 0.00980851
R7557 VGND.n896 VGND 0.00980851
R7558 VGND VGND.n1331 0.00980851
R7559 VGND.n888 VGND 0.00980851
R7560 VGND.n2698 VGND.n2697 0.00182979
R7561 VGND.n358 VGND.n357 0.00182979
R7562 VGND.n365 VGND.n364 0.00182979
R7563 VGND.n367 VGND.n354 0.00182979
R7564 VGND.n376 VGND.n375 0.00182979
R7565 VGND.n378 VGND.n353 0.00182979
R7566 VGND.n389 VGND.n386 0.00182979
R7567 VGND.n2707 VGND.n325 0.00182979
R7568 VGND.n2725 VGND.n314 0.00182979
R7569 VGND.n2740 VGND.n309 0.00182979
R7570 VGND.n311 VGND.n300 0.00182979
R7571 VGND.n2734 VGND.n2733 0.00182979
R7572 VGND.n2778 VGND.n293 0.00182979
R7573 VGND.n2772 VGND.n296 0.00182979
R7574 VGND.n2942 VGND.n203 0.00182979
R7575 XThR.Tn[2].n2 XThR.Tn[2].n1 332.332
R7576 XThR.Tn[2].n2 XThR.Tn[2].n0 296.493
R7577 XThR.Tn[2] XThR.Tn[2].n82 161.363
R7578 XThR.Tn[2] XThR.Tn[2].n77 161.363
R7579 XThR.Tn[2] XThR.Tn[2].n72 161.363
R7580 XThR.Tn[2] XThR.Tn[2].n67 161.363
R7581 XThR.Tn[2] XThR.Tn[2].n62 161.363
R7582 XThR.Tn[2] XThR.Tn[2].n57 161.363
R7583 XThR.Tn[2] XThR.Tn[2].n52 161.363
R7584 XThR.Tn[2] XThR.Tn[2].n47 161.363
R7585 XThR.Tn[2] XThR.Tn[2].n42 161.363
R7586 XThR.Tn[2] XThR.Tn[2].n37 161.363
R7587 XThR.Tn[2] XThR.Tn[2].n32 161.363
R7588 XThR.Tn[2] XThR.Tn[2].n27 161.363
R7589 XThR.Tn[2] XThR.Tn[2].n22 161.363
R7590 XThR.Tn[2] XThR.Tn[2].n17 161.363
R7591 XThR.Tn[2] XThR.Tn[2].n12 161.363
R7592 XThR.Tn[2] XThR.Tn[2].n10 161.363
R7593 XThR.Tn[2].n84 XThR.Tn[2].n83 161.3
R7594 XThR.Tn[2].n79 XThR.Tn[2].n78 161.3
R7595 XThR.Tn[2].n74 XThR.Tn[2].n73 161.3
R7596 XThR.Tn[2].n69 XThR.Tn[2].n68 161.3
R7597 XThR.Tn[2].n64 XThR.Tn[2].n63 161.3
R7598 XThR.Tn[2].n59 XThR.Tn[2].n58 161.3
R7599 XThR.Tn[2].n54 XThR.Tn[2].n53 161.3
R7600 XThR.Tn[2].n49 XThR.Tn[2].n48 161.3
R7601 XThR.Tn[2].n44 XThR.Tn[2].n43 161.3
R7602 XThR.Tn[2].n39 XThR.Tn[2].n38 161.3
R7603 XThR.Tn[2].n34 XThR.Tn[2].n33 161.3
R7604 XThR.Tn[2].n29 XThR.Tn[2].n28 161.3
R7605 XThR.Tn[2].n24 XThR.Tn[2].n23 161.3
R7606 XThR.Tn[2].n19 XThR.Tn[2].n18 161.3
R7607 XThR.Tn[2].n14 XThR.Tn[2].n13 161.3
R7608 XThR.Tn[2].n82 XThR.Tn[2].t65 161.106
R7609 XThR.Tn[2].n77 XThR.Tn[2].t72 161.106
R7610 XThR.Tn[2].n72 XThR.Tn[2].t51 161.106
R7611 XThR.Tn[2].n67 XThR.Tn[2].t36 161.106
R7612 XThR.Tn[2].n62 XThR.Tn[2].t64 161.106
R7613 XThR.Tn[2].n57 XThR.Tn[2].t26 161.106
R7614 XThR.Tn[2].n52 XThR.Tn[2].t69 161.106
R7615 XThR.Tn[2].n47 XThR.Tn[2].t49 161.106
R7616 XThR.Tn[2].n42 XThR.Tn[2].t35 161.106
R7617 XThR.Tn[2].n37 XThR.Tn[2].t41 161.106
R7618 XThR.Tn[2].n32 XThR.Tn[2].t25 161.106
R7619 XThR.Tn[2].n27 XThR.Tn[2].t50 161.106
R7620 XThR.Tn[2].n22 XThR.Tn[2].t23 161.106
R7621 XThR.Tn[2].n17 XThR.Tn[2].t67 161.106
R7622 XThR.Tn[2].n12 XThR.Tn[2].t31 161.106
R7623 XThR.Tn[2].n10 XThR.Tn[2].t14 161.106
R7624 XThR.Tn[2].n83 XThR.Tn[2].t38 159.978
R7625 XThR.Tn[2].n78 XThR.Tn[2].t46 159.978
R7626 XThR.Tn[2].n73 XThR.Tn[2].t29 159.978
R7627 XThR.Tn[2].n68 XThR.Tn[2].t13 159.978
R7628 XThR.Tn[2].n63 XThR.Tn[2].t37 159.978
R7629 XThR.Tn[2].n58 XThR.Tn[2].t63 159.978
R7630 XThR.Tn[2].n53 XThR.Tn[2].t45 159.978
R7631 XThR.Tn[2].n48 XThR.Tn[2].t27 159.978
R7632 XThR.Tn[2].n43 XThR.Tn[2].t12 159.978
R7633 XThR.Tn[2].n38 XThR.Tn[2].t20 159.978
R7634 XThR.Tn[2].n33 XThR.Tn[2].t62 159.978
R7635 XThR.Tn[2].n28 XThR.Tn[2].t28 159.978
R7636 XThR.Tn[2].n23 XThR.Tn[2].t60 159.978
R7637 XThR.Tn[2].n18 XThR.Tn[2].t43 159.978
R7638 XThR.Tn[2].n13 XThR.Tn[2].t66 159.978
R7639 XThR.Tn[2].n82 XThR.Tn[2].t53 145.038
R7640 XThR.Tn[2].n77 XThR.Tn[2].t19 145.038
R7641 XThR.Tn[2].n72 XThR.Tn[2].t59 145.038
R7642 XThR.Tn[2].n67 XThR.Tn[2].t42 145.038
R7643 XThR.Tn[2].n62 XThR.Tn[2].t73 145.038
R7644 XThR.Tn[2].n57 XThR.Tn[2].t52 145.038
R7645 XThR.Tn[2].n52 XThR.Tn[2].t61 145.038
R7646 XThR.Tn[2].n47 XThR.Tn[2].t44 145.038
R7647 XThR.Tn[2].n42 XThR.Tn[2].t39 145.038
R7648 XThR.Tn[2].n37 XThR.Tn[2].t70 145.038
R7649 XThR.Tn[2].n32 XThR.Tn[2].t34 145.038
R7650 XThR.Tn[2].n27 XThR.Tn[2].t58 145.038
R7651 XThR.Tn[2].n22 XThR.Tn[2].t32 145.038
R7652 XThR.Tn[2].n17 XThR.Tn[2].t15 145.038
R7653 XThR.Tn[2].n12 XThR.Tn[2].t40 145.038
R7654 XThR.Tn[2].n10 XThR.Tn[2].t21 145.038
R7655 XThR.Tn[2].n83 XThR.Tn[2].t71 143.911
R7656 XThR.Tn[2].n78 XThR.Tn[2].t33 143.911
R7657 XThR.Tn[2].n73 XThR.Tn[2].t17 143.911
R7658 XThR.Tn[2].n68 XThR.Tn[2].t56 143.911
R7659 XThR.Tn[2].n63 XThR.Tn[2].t24 143.911
R7660 XThR.Tn[2].n58 XThR.Tn[2].t68 143.911
R7661 XThR.Tn[2].n53 XThR.Tn[2].t18 143.911
R7662 XThR.Tn[2].n48 XThR.Tn[2].t57 143.911
R7663 XThR.Tn[2].n43 XThR.Tn[2].t54 143.911
R7664 XThR.Tn[2].n38 XThR.Tn[2].t22 143.911
R7665 XThR.Tn[2].n33 XThR.Tn[2].t48 143.911
R7666 XThR.Tn[2].n28 XThR.Tn[2].t16 143.911
R7667 XThR.Tn[2].n23 XThR.Tn[2].t47 143.911
R7668 XThR.Tn[2].n18 XThR.Tn[2].t30 143.911
R7669 XThR.Tn[2].n13 XThR.Tn[2].t55 143.911
R7670 XThR.Tn[2].n7 XThR.Tn[2].n6 135.249
R7671 XThR.Tn[2].n9 XThR.Tn[2].n3 98.982
R7672 XThR.Tn[2].n8 XThR.Tn[2].n4 98.982
R7673 XThR.Tn[2].n7 XThR.Tn[2].n5 98.982
R7674 XThR.Tn[2].n9 XThR.Tn[2].n8 36.2672
R7675 XThR.Tn[2].n8 XThR.Tn[2].n7 36.2672
R7676 XThR.Tn[2].n88 XThR.Tn[2].n9 32.6405
R7677 XThR.Tn[2].n1 XThR.Tn[2].t10 26.5955
R7678 XThR.Tn[2].n1 XThR.Tn[2].t9 26.5955
R7679 XThR.Tn[2].n0 XThR.Tn[2].t11 26.5955
R7680 XThR.Tn[2].n0 XThR.Tn[2].t8 26.5955
R7681 XThR.Tn[2].n3 XThR.Tn[2].t6 24.9236
R7682 XThR.Tn[2].n3 XThR.Tn[2].t7 24.9236
R7683 XThR.Tn[2].n4 XThR.Tn[2].t5 24.9236
R7684 XThR.Tn[2].n4 XThR.Tn[2].t4 24.9236
R7685 XThR.Tn[2].n5 XThR.Tn[2].t2 24.9236
R7686 XThR.Tn[2].n5 XThR.Tn[2].t3 24.9236
R7687 XThR.Tn[2].n6 XThR.Tn[2].t0 24.9236
R7688 XThR.Tn[2].n6 XThR.Tn[2].t1 24.9236
R7689 XThR.Tn[2] XThR.Tn[2].n2 23.3605
R7690 XThR.Tn[2] XThR.Tn[2].n88 6.7205
R7691 XThR.Tn[2].n88 XThR.Tn[2] 6.30883
R7692 XThR.Tn[2] XThR.Tn[2].n11 5.34038
R7693 XThR.Tn[2].n16 XThR.Tn[2].n15 4.5005
R7694 XThR.Tn[2].n21 XThR.Tn[2].n20 4.5005
R7695 XThR.Tn[2].n26 XThR.Tn[2].n25 4.5005
R7696 XThR.Tn[2].n31 XThR.Tn[2].n30 4.5005
R7697 XThR.Tn[2].n36 XThR.Tn[2].n35 4.5005
R7698 XThR.Tn[2].n41 XThR.Tn[2].n40 4.5005
R7699 XThR.Tn[2].n46 XThR.Tn[2].n45 4.5005
R7700 XThR.Tn[2].n51 XThR.Tn[2].n50 4.5005
R7701 XThR.Tn[2].n56 XThR.Tn[2].n55 4.5005
R7702 XThR.Tn[2].n61 XThR.Tn[2].n60 4.5005
R7703 XThR.Tn[2].n66 XThR.Tn[2].n65 4.5005
R7704 XThR.Tn[2].n71 XThR.Tn[2].n70 4.5005
R7705 XThR.Tn[2].n76 XThR.Tn[2].n75 4.5005
R7706 XThR.Tn[2].n81 XThR.Tn[2].n80 4.5005
R7707 XThR.Tn[2].n86 XThR.Tn[2].n85 4.5005
R7708 XThR.Tn[2].n87 XThR.Tn[2] 3.70586
R7709 XThR.Tn[2].n16 XThR.Tn[2] 2.52282
R7710 XThR.Tn[2].n21 XThR.Tn[2] 2.52282
R7711 XThR.Tn[2].n26 XThR.Tn[2] 2.52282
R7712 XThR.Tn[2].n31 XThR.Tn[2] 2.52282
R7713 XThR.Tn[2].n36 XThR.Tn[2] 2.52282
R7714 XThR.Tn[2].n41 XThR.Tn[2] 2.52282
R7715 XThR.Tn[2].n46 XThR.Tn[2] 2.52282
R7716 XThR.Tn[2].n51 XThR.Tn[2] 2.52282
R7717 XThR.Tn[2].n56 XThR.Tn[2] 2.52282
R7718 XThR.Tn[2].n61 XThR.Tn[2] 2.52282
R7719 XThR.Tn[2].n66 XThR.Tn[2] 2.52282
R7720 XThR.Tn[2].n71 XThR.Tn[2] 2.52282
R7721 XThR.Tn[2].n76 XThR.Tn[2] 2.52282
R7722 XThR.Tn[2].n81 XThR.Tn[2] 2.52282
R7723 XThR.Tn[2].n86 XThR.Tn[2] 2.52282
R7724 XThR.Tn[2].n84 XThR.Tn[2] 1.08677
R7725 XThR.Tn[2].n79 XThR.Tn[2] 1.08677
R7726 XThR.Tn[2].n74 XThR.Tn[2] 1.08677
R7727 XThR.Tn[2].n69 XThR.Tn[2] 1.08677
R7728 XThR.Tn[2].n64 XThR.Tn[2] 1.08677
R7729 XThR.Tn[2].n59 XThR.Tn[2] 1.08677
R7730 XThR.Tn[2].n54 XThR.Tn[2] 1.08677
R7731 XThR.Tn[2].n49 XThR.Tn[2] 1.08677
R7732 XThR.Tn[2].n44 XThR.Tn[2] 1.08677
R7733 XThR.Tn[2].n39 XThR.Tn[2] 1.08677
R7734 XThR.Tn[2].n34 XThR.Tn[2] 1.08677
R7735 XThR.Tn[2].n29 XThR.Tn[2] 1.08677
R7736 XThR.Tn[2].n24 XThR.Tn[2] 1.08677
R7737 XThR.Tn[2].n19 XThR.Tn[2] 1.08677
R7738 XThR.Tn[2].n14 XThR.Tn[2] 1.08677
R7739 XThR.Tn[2] XThR.Tn[2].n16 0.839786
R7740 XThR.Tn[2] XThR.Tn[2].n21 0.839786
R7741 XThR.Tn[2] XThR.Tn[2].n26 0.839786
R7742 XThR.Tn[2] XThR.Tn[2].n31 0.839786
R7743 XThR.Tn[2] XThR.Tn[2].n36 0.839786
R7744 XThR.Tn[2] XThR.Tn[2].n41 0.839786
R7745 XThR.Tn[2] XThR.Tn[2].n46 0.839786
R7746 XThR.Tn[2] XThR.Tn[2].n51 0.839786
R7747 XThR.Tn[2] XThR.Tn[2].n56 0.839786
R7748 XThR.Tn[2] XThR.Tn[2].n61 0.839786
R7749 XThR.Tn[2] XThR.Tn[2].n66 0.839786
R7750 XThR.Tn[2] XThR.Tn[2].n71 0.839786
R7751 XThR.Tn[2] XThR.Tn[2].n76 0.839786
R7752 XThR.Tn[2] XThR.Tn[2].n81 0.839786
R7753 XThR.Tn[2] XThR.Tn[2].n86 0.839786
R7754 XThR.Tn[2].n11 XThR.Tn[2] 0.499542
R7755 XThR.Tn[2].n85 XThR.Tn[2] 0.063
R7756 XThR.Tn[2].n80 XThR.Tn[2] 0.063
R7757 XThR.Tn[2].n75 XThR.Tn[2] 0.063
R7758 XThR.Tn[2].n70 XThR.Tn[2] 0.063
R7759 XThR.Tn[2].n65 XThR.Tn[2] 0.063
R7760 XThR.Tn[2].n60 XThR.Tn[2] 0.063
R7761 XThR.Tn[2].n55 XThR.Tn[2] 0.063
R7762 XThR.Tn[2].n50 XThR.Tn[2] 0.063
R7763 XThR.Tn[2].n45 XThR.Tn[2] 0.063
R7764 XThR.Tn[2].n40 XThR.Tn[2] 0.063
R7765 XThR.Tn[2].n35 XThR.Tn[2] 0.063
R7766 XThR.Tn[2].n30 XThR.Tn[2] 0.063
R7767 XThR.Tn[2].n25 XThR.Tn[2] 0.063
R7768 XThR.Tn[2].n20 XThR.Tn[2] 0.063
R7769 XThR.Tn[2].n15 XThR.Tn[2] 0.063
R7770 XThR.Tn[2].n87 XThR.Tn[2] 0.0540714
R7771 XThR.Tn[2] XThR.Tn[2].n87 0.038
R7772 XThR.Tn[2].n11 XThR.Tn[2] 0.0143889
R7773 XThR.Tn[2].n85 XThR.Tn[2].n84 0.00771154
R7774 XThR.Tn[2].n80 XThR.Tn[2].n79 0.00771154
R7775 XThR.Tn[2].n75 XThR.Tn[2].n74 0.00771154
R7776 XThR.Tn[2].n70 XThR.Tn[2].n69 0.00771154
R7777 XThR.Tn[2].n65 XThR.Tn[2].n64 0.00771154
R7778 XThR.Tn[2].n60 XThR.Tn[2].n59 0.00771154
R7779 XThR.Tn[2].n55 XThR.Tn[2].n54 0.00771154
R7780 XThR.Tn[2].n50 XThR.Tn[2].n49 0.00771154
R7781 XThR.Tn[2].n45 XThR.Tn[2].n44 0.00771154
R7782 XThR.Tn[2].n40 XThR.Tn[2].n39 0.00771154
R7783 XThR.Tn[2].n35 XThR.Tn[2].n34 0.00771154
R7784 XThR.Tn[2].n30 XThR.Tn[2].n29 0.00771154
R7785 XThR.Tn[2].n25 XThR.Tn[2].n24 0.00771154
R7786 XThR.Tn[2].n20 XThR.Tn[2].n19 0.00771154
R7787 XThR.Tn[2].n15 XThR.Tn[2].n14 0.00771154
R7788 VPWR.n2837 VPWR.n2823 2618.82
R7789 VPWR.n2835 VPWR.n2829 2618.82
R7790 VPWR.n2853 VPWR.n2823 1916.47
R7791 VPWR.n2828 VPWR.n2827 1916.47
R7792 VPWR.n2827 VPWR.n2821 1916.47
R7793 VPWR.n2829 VPWR.n2822 1916.47
R7794 VPWR.n2852 VPWR.n2824 1912.94
R7795 VPWR.n2849 VPWR.n2843 1560
R7796 VPWR.n2850 VPWR.n2824 1408.24
R7797 VPWR.n2853 VPWR.n2852 1210.59
R7798 VPWR.n2851 VPWR.n2821 1210.59
R7799 VPWR.n2380 VPWR.t148 1005.7
R7800 VPWR.t366 VPWR.n485 1005.7
R7801 VPWR.t215 VPWR.n2210 1005.7
R7802 VPWR.n639 VPWR.t323 1005.7
R7803 VPWR.n2184 VPWR.t49 1005.7
R7804 VPWR.t156 VPWR.n677 1005.7
R7805 VPWR.t116 VPWR.n2014 1005.7
R7806 VPWR.n831 VPWR.t221 1005.7
R7807 VPWR.n1988 VPWR.t44 1005.7
R7808 VPWR.t228 VPWR.n869 1005.7
R7809 VPWR.n447 VPWR.t36 1005.7
R7810 VPWR.t336 VPWR.n1818 1005.7
R7811 VPWR.t315 VPWR.n2406 1005.7
R7812 VPWR.n1023 VPWR.t188 1005.7
R7813 VPWR.t358 VPWR.n293 1005.7
R7814 VPWR.n1792 VPWR.t299 1005.7
R7815 VPWR.n2591 VPWR.t250 1005.7
R7816 VPWR.n1062 VPWR.t134 1005.7
R7817 VPWR.t1191 VPWR.n2309 983.14
R7818 VPWR.n2310 VPWR.t689 983.14
R7819 VPWR.t1492 VPWR.n2319 983.14
R7820 VPWR.n2320 VPWR.t1508 983.14
R7821 VPWR.t1595 VPWR.n2329 983.14
R7822 VPWR.n2330 VPWR.t959 983.14
R7823 VPWR.t1579 VPWR.n2339 983.14
R7824 VPWR.n2340 VPWR.t900 983.14
R7825 VPWR.t1684 VPWR.n2349 983.14
R7826 VPWR.n2350 VPWR.t745 983.14
R7827 VPWR.t1605 VPWR.n2359 983.14
R7828 VPWR.n2360 VPWR.t1573 983.14
R7829 VPWR.t1077 VPWR.n2369 983.14
R7830 VPWR.n2370 VPWR.t412 983.14
R7831 VPWR.t1846 VPWR.n2379 983.14
R7832 VPWR.n542 VPWR.t1201 983.14
R7833 VPWR.n541 VPWR.t1674 983.14
R7834 VPWR.n537 VPWR.t1470 983.14
R7835 VPWR.n533 VPWR.t390 983.14
R7836 VPWR.n529 VPWR.t1335 983.14
R7837 VPWR.n525 VPWR.t1145 983.14
R7838 VPWR.n521 VPWR.t800 983.14
R7839 VPWR.n517 VPWR.t831 983.14
R7840 VPWR.n513 VPWR.t839 983.14
R7841 VPWR.n509 VPWR.t518 983.14
R7842 VPWR.n505 VPWR.t1310 983.14
R7843 VPWR.n501 VPWR.t1258 983.14
R7844 VPWR.n497 VPWR.t1306 983.14
R7845 VPWR.n493 VPWR.t1358 983.14
R7846 VPWR.n489 VPWR.t598 983.14
R7847 VPWR.n2281 VPWR.t852 983.14
R7848 VPWR.n2280 VPWR.t1709 983.14
R7849 VPWR.n2271 VPWR.t1446 983.14
R7850 VPWR.n2270 VPWR.t1274 983.14
R7851 VPWR.n2261 VPWR.t1695 983.14
R7852 VPWR.n2260 VPWR.t911 983.14
R7853 VPWR.n2251 VPWR.t482 983.14
R7854 VPWR.n2250 VPWR.t886 983.14
R7855 VPWR.n2241 VPWR.t884 983.14
R7856 VPWR.n2240 VPWR.t723 983.14
R7857 VPWR.n2231 VPWR.t1174 983.14
R7858 VPWR.n2230 VPWR.t1828 983.14
R7859 VPWR.n2221 VPWR.t1916 983.14
R7860 VPWR.n2220 VPWR.t564 983.14
R7861 VPWR.n2211 VPWR.t780 983.14
R7862 VPWR.t1018 VPWR.n582 983.14
R7863 VPWR.t471 VPWR.n586 983.14
R7864 VPWR.t1460 VPWR.n590 983.14
R7865 VPWR.t396 VPWR.n594 983.14
R7866 VPWR.t1545 VPWR.n598 983.14
R7867 VPWR.t1155 VPWR.n602 983.14
R7868 VPWR.t810 VPWR.n606 983.14
R7869 VPWR.t932 VPWR.n610 983.14
R7870 VPWR.t945 VPWR.n614 983.14
R7871 VPWR.t1234 VPWR.n618 983.14
R7872 VPWR.t1320 VPWR.n622 983.14
R7873 VPWR.t1248 VPWR.n626 983.14
R7874 VPWR.t1715 VPWR.n630 983.14
R7875 VPWR.t735 VPWR.n634 983.14
R7876 VPWR.t604 VPWR.n638 983.14
R7877 VPWR.t824 VPWR.n2113 983.14
R7878 VPWR.n2114 VPWR.t1551 983.14
R7879 VPWR.t1482 VPWR.n2123 983.14
R7880 VPWR.n2124 VPWR.t998 983.14
R7881 VPWR.t1329 VPWR.n2133 983.14
R7882 VPWR.n2134 VPWR.t620 983.14
R7883 VPWR.t1589 VPWR.n2143 983.14
R7884 VPWR.n2144 VPWR.t871 983.14
R7885 VPWR.t544 VPWR.n2153 983.14
R7886 VPWR.n2154 VPWR.t506 983.14
R7887 VPWR.t1664 VPWR.n2163 983.14
R7888 VPWR.n2164 VPWR.t1282 983.14
R7889 VPWR.t1296 VPWR.n2173 983.14
R7890 VPWR.n2174 VPWR.t1496 983.14
R7891 VPWR.t522 VPWR.n2183 983.14
R7892 VPWR.n734 VPWR.t1189 983.14
R7893 VPWR.n733 VPWR.t687 983.14
R7894 VPWR.n729 VPWR.t1494 983.14
R7895 VPWR.n725 VPWR.t1506 983.14
R7896 VPWR.n721 VPWR.t1593 983.14
R7897 VPWR.n717 VPWR.t957 983.14
R7898 VPWR.n713 VPWR.t1577 983.14
R7899 VPWR.n709 VPWR.t898 983.14
R7900 VPWR.n705 VPWR.t1682 983.14
R7901 VPWR.n701 VPWR.t743 983.14
R7902 VPWR.n697 VPWR.t1619 983.14
R7903 VPWR.n693 VPWR.t1571 983.14
R7904 VPWR.n689 VPWR.t1075 983.14
R7905 VPWR.n685 VPWR.t410 983.14
R7906 VPWR.n681 VPWR.t1844 983.14
R7907 VPWR.n2085 VPWR.t1012 983.14
R7908 VPWR.n2084 VPWR.t1028 983.14
R7909 VPWR.n2075 VPWR.t1488 983.14
R7910 VPWR.n2074 VPWR.t1510 983.14
R7911 VPWR.n2065 VPWR.t1625 983.14
R7912 VPWR.n2064 VPWR.t654 983.14
R7913 VPWR.n2055 VPWR.t1585 983.14
R7914 VPWR.n2054 VPWR.t664 983.14
R7915 VPWR.n2045 VPWR.t1034 983.14
R7916 VPWR.n2044 VPWR.t751 983.14
R7917 VPWR.n2035 VPWR.t878 983.14
R7918 VPWR.n2034 VPWR.t1567 983.14
R7919 VPWR.n2025 VPWR.t1079 983.14
R7920 VPWR.n2024 VPWR.t418 983.14
R7921 VPWR.n2015 VPWR.t1848 983.14
R7922 VPWR.t433 VPWR.n774 983.14
R7923 VPWR.t1707 VPWR.n778 983.14
R7924 VPWR.t1448 VPWR.n782 983.14
R7925 VPWR.t1270 VPWR.n786 983.14
R7926 VPWR.t1693 VPWR.n790 983.14
R7927 VPWR.t909 VPWR.n794 983.14
R7928 VPWR.t480 VPWR.n798 983.14
R7929 VPWR.t648 VPWR.n802 983.14
R7930 VPWR.t882 VPWR.n806 983.14
R7931 VPWR.t721 VPWR.n810 983.14
R7932 VPWR.t1172 VPWR.n814 983.14
R7933 VPWR.t536 VPWR.n818 983.14
R7934 VPWR.t1912 VPWR.n822 983.14
R7935 VPWR.t562 VPWR.n826 983.14
R7936 VPWR.t776 VPWR.n830 983.14
R7937 VPWR.t826 VPWR.n1917 983.14
R7938 VPWR.n1918 VPWR.t1553 983.14
R7939 VPWR.t1480 VPWR.n1927 983.14
R7940 VPWR.n1928 VPWR.t1390 983.14
R7941 VPWR.t1331 VPWR.n1937 983.14
R7942 VPWR.n1938 VPWR.t622 983.14
R7943 VPWR.t790 VPWR.n1947 983.14
R7944 VPWR.n1948 VPWR.t873 983.14
R7945 VPWR.t546 VPWR.n1957 983.14
R7946 VPWR.n1958 VPWR.t508 983.14
R7947 VPWR.t1666 VPWR.n1967 983.14
R7948 VPWR.n1968 VPWR.t1284 983.14
R7949 VPWR.t1298 VPWR.n1977 983.14
R7950 VPWR.n1978 VPWR.t1498 983.14
R7951 VPWR.t524 VPWR.n1987 983.14
R7952 VPWR.n926 VPWR.t431 983.14
R7953 VPWR.n925 VPWR.t1705 983.14
R7954 VPWR.n921 VPWR.t1450 983.14
R7955 VPWR.n917 VPWR.t1268 983.14
R7956 VPWR.n913 VPWR.t1672 983.14
R7957 VPWR.n909 VPWR.t907 983.14
R7958 VPWR.n905 VPWR.t478 983.14
R7959 VPWR.n901 VPWR.t644 983.14
R7960 VPWR.n897 VPWR.t880 983.14
R7961 VPWR.n893 VPWR.t719 983.14
R7962 VPWR.n889 VPWR.t1170 983.14
R7963 VPWR.n885 VPWR.t534 983.14
R7964 VPWR.n881 VPWR.t1908 983.14
R7965 VPWR.n877 VPWR.t560 983.14
R7966 VPWR.n873 VPWR.t774 983.14
R7967 VPWR.t828 VPWR.n390 983.14
R7968 VPWR.t1555 VPWR.n394 983.14
R7969 VPWR.t1478 VPWR.n398 983.14
R7970 VPWR.t1394 VPWR.n402 983.14
R7971 VPWR.t1333 VPWR.n406 983.14
R7972 VPWR.t624 VPWR.n410 983.14
R7973 VPWR.t792 VPWR.n414 983.14
R7974 VPWR.t658 VPWR.n418 983.14
R7975 VPWR.t548 VPWR.n422 983.14
R7976 VPWR.t510 VPWR.n426 983.14
R7977 VPWR.t1668 VPWR.n430 983.14
R7978 VPWR.t1286 VPWR.n434 983.14
R7979 VPWR.t1300 VPWR.n438 983.14
R7980 VPWR.t1500 VPWR.n442 983.14
R7981 VPWR.t528 VPWR.n446 983.14
R7982 VPWR.n1889 VPWR.t1016 983.14
R7983 VPWR.n1888 VPWR.t1680 983.14
R7984 VPWR.n1879 VPWR.t1462 983.14
R7985 VPWR.n1878 VPWR.t394 983.14
R7986 VPWR.n1869 VPWR.t1541 983.14
R7987 VPWR.n1868 VPWR.t1151 983.14
R7988 VPWR.n1859 VPWR.t806 983.14
R7989 VPWR.n1858 VPWR.t930 983.14
R7990 VPWR.n1849 VPWR.t941 983.14
R7991 VPWR.n1848 VPWR.t1232 983.14
R7992 VPWR.n1839 VPWR.t1316 983.14
R7993 VPWR.n1838 VPWR.t1246 983.14
R7994 VPWR.n1829 VPWR.t1713 983.14
R7995 VPWR.n1828 VPWR.t733 983.14
R7996 VPWR.n1819 VPWR.t602 983.14
R7997 VPWR.n2477 VPWR.t1020 983.14
R7998 VPWR.n2476 VPWR.t473 983.14
R7999 VPWR.n2467 VPWR.t1458 983.14
R8000 VPWR.n2466 VPWR.t1514 983.14
R8001 VPWR.n2457 VPWR.t1547 983.14
R8002 VPWR.n2456 VPWR.t1134 983.14
R8003 VPWR.n2447 VPWR.t812 983.14
R8004 VPWR.n2446 VPWR.t934 983.14
R8005 VPWR.n2437 VPWR.t947 983.14
R8006 VPWR.n2436 VPWR.t1236 983.14
R8007 VPWR.n2427 VPWR.t1322 983.14
R8008 VPWR.n2426 VPWR.t1250 983.14
R8009 VPWR.n2417 VPWR.t1717 983.14
R8010 VPWR.n2416 VPWR.t737 983.14
R8011 VPWR.n2407 VPWR.t608 983.14
R8012 VPWR.t854 VPWR.n966 983.14
R8013 VPWR.t1900 VPWR.n970 983.14
R8014 VPWR.t1440 VPWR.n974 983.14
R8015 VPWR.t1280 VPWR.n978 983.14
R8016 VPWR.t1701 VPWR.n982 983.14
R8017 VPWR.t917 VPWR.n986 983.14
R8018 VPWR.t488 VPWR.n990 983.14
R8019 VPWR.t890 VPWR.n994 983.14
R8020 VPWR.t1183 VPWR.n998 983.14
R8021 VPWR.t725 VPWR.n1002 983.14
R8022 VPWR.t1613 VPWR.n1006 983.14
R8023 VPWR.t1830 VPWR.n1010 983.14
R8024 VPWR.t1920 VPWR.n1014 983.14
R8025 VPWR.t402 VPWR.n1018 983.14
R8026 VPWR.t786 VPWR.n1022 983.14
R8027 VPWR.n350 VPWR.t1203 983.14
R8028 VPWR.n349 VPWR.t1676 983.14
R8029 VPWR.n345 VPWR.t1466 983.14
R8030 VPWR.n341 VPWR.t392 983.14
R8031 VPWR.n337 VPWR.t1337 983.14
R8032 VPWR.n333 VPWR.t1147 983.14
R8033 VPWR.n329 VPWR.t802 983.14
R8034 VPWR.n325 VPWR.t835 983.14
R8035 VPWR.n321 VPWR.t841 983.14
R8036 VPWR.n317 VPWR.t1230 983.14
R8037 VPWR.n313 VPWR.t1312 983.14
R8038 VPWR.n309 VPWR.t1260 983.14
R8039 VPWR.n305 VPWR.t1711 983.14
R8040 VPWR.n301 VPWR.t1360 983.14
R8041 VPWR.n297 VPWR.t600 983.14
R8042 VPWR.t269 VPWR.n1468 983.14
R8043 VPWR.t371 VPWR.n1475 983.14
R8044 VPWR.t142 VPWR.n1481 983.14
R8045 VPWR.t244 VPWR.n1492 983.14
R8046 VPWR.n1493 VPWR.t266 983.14
R8047 VPWR.t17 VPWR.n1506 983.14
R8048 VPWR.n1507 VPWR.t139 983.14
R8049 VPWR.t280 VPWR.n1520 983.14
R8050 VPWR.n1521 VPWR.t296 983.14
R8051 VPWR.n1536 VPWR.t39 983.14
R8052 VPWR.n1535 VPWR.t169 983.14
R8053 VPWR.n1761 VPWR.t210 983.14
R8054 VPWR.n1760 VPWR.t33 983.14
R8055 VPWR.n1749 VPWR.t83 983.14
R8056 VPWR.t191 VPWR.n1791 983.14
R8057 VPWR.t197 VPWR.n2506 983.14
R8058 VPWR.n2507 VPWR.t309 983.14
R8059 VPWR.t74 VPWR.n2518 983.14
R8060 VPWR.n2519 VPWR.t185 983.14
R8061 VPWR.t194 VPWR.n2530 983.14
R8062 VPWR.n2531 VPWR.t350 983.14
R8063 VPWR.t71 VPWR.n2542 983.14
R8064 VPWR.n2543 VPWR.t231 983.14
R8065 VPWR.t247 VPWR.n2554 983.14
R8066 VPWR.n2555 VPWR.t377 983.14
R8067 VPWR.t121 VPWR.n2566 983.14
R8068 VPWR.n2567 VPWR.t151 983.14
R8069 VPWR.t1 VPWR.n2578 983.14
R8070 VPWR.n2579 VPWR.t20 983.14
R8071 VPWR.t145 VPWR.n2590 983.14
R8072 VPWR.n1594 VPWR.t80 983.14
R8073 VPWR.n1593 VPWR.t182 983.14
R8074 VPWR.t347 VPWR.n1182 983.14
R8075 VPWR.t65 VPWR.n1185 983.14
R8076 VPWR.n1220 VPWR.t77 983.14
R8077 VPWR.n1219 VPWR.t236 983.14
R8078 VPWR.n1216 VPWR.t344 983.14
R8079 VPWR.n1213 VPWR.t105 983.14
R8080 VPWR.n1205 VPWR.t131 983.14
R8081 VPWR.n1202 VPWR.t258 983.14
R8082 VPWR.n1199 VPWR.t4 983.14
R8083 VPWR.n1191 VPWR.t25 983.14
R8084 VPWR.n1188 VPWR.t263 983.14
R8085 VPWR.n1740 VPWR.t291 983.14
R8086 VPWR.n1739 VPWR.t10 983.14
R8087 VPWR.n1308 VPWR.t423 877.144
R8088 VPWR.n2723 VPWR.t1792 877.144
R8089 VPWR.n2843 VPWR.n2822 857.648
R8090 VPWR.n1122 VPWR.t313 738.074
R8091 VPWR.n99 VPWR.t53 738.074
R8092 VPWR.n290 VPWR.t1118 738.074
R8093 VPWR.n68 VPWR.t122 738.074
R8094 VPWR.n346 VPWR.t1204 738.074
R8095 VPWR.n98 VPWR.t198 738.074
R8096 VPWR.n963 VPWR.t1104 738.074
R8097 VPWR.n356 VPWR.t1112 738.074
R8098 VPWR.n357 VPWR.t1021 738.074
R8099 VPWR.n318 VPWR.t836 738.074
R8100 VPWR.n75 VPWR.t232 738.074
R8101 VPWR.n971 VPWR.t1901 738.074
R8102 VPWR.n369 VPWR.t813 738.074
R8103 VPWR.n322 VPWR.t803 738.074
R8104 VPWR.n80 VPWR.t72 738.074
R8105 VPWR.n932 VPWR.t1116 738.074
R8106 VPWR.n933 VPWR.t1017 738.074
R8107 VPWR.n936 VPWR.t1681 738.074
R8108 VPWR.n387 VPWR.t1122 738.074
R8109 VPWR.n391 VPWR.t829 738.074
R8110 VPWR.n395 VPWR.t1556 738.074
R8111 VPWR.n365 VPWR.t1548 738.074
R8112 VPWR.n330 VPWR.t1338 738.074
R8113 VPWR.n86 VPWR.t195 738.074
R8114 VPWR.n937 VPWR.t1463 738.074
R8115 VPWR.n403 VPWR.t1395 738.074
R8116 VPWR.n364 VPWR.t1515 738.074
R8117 VPWR.n334 VPWR.t393 738.074
R8118 VPWR.n87 VPWR.t186 738.074
R8119 VPWR.n481 VPWR.t1131 738.074
R8120 VPWR.n480 VPWR.t1192 738.074
R8121 VPWR.n477 VPWR.t690 738.074
R8122 VPWR.n476 VPWR.t1493 738.074
R8123 VPWR.n472 VPWR.t1596 738.074
R8124 VPWR.n469 VPWR.t960 738.074
R8125 VPWR.n468 VPWR.t1580 738.074
R8126 VPWR.n465 VPWR.t901 738.074
R8127 VPWR.n464 VPWR.t1685 738.074
R8128 VPWR.n461 VPWR.t746 738.074
R8129 VPWR.n460 VPWR.t1606 738.074
R8130 VPWR.n457 VPWR.t1574 738.074
R8131 VPWR.n456 VPWR.t1078 738.074
R8132 VPWR.n453 VPWR.t413 738.074
R8133 VPWR.n452 VPWR.t1847 738.074
R8134 VPWR.n473 VPWR.t1509 738.074
R8135 VPWR.n482 VPWR.t1120 738.074
R8136 VPWR.n538 VPWR.t1202 738.074
R8137 VPWR.n534 VPWR.t1675 738.074
R8138 VPWR.n530 VPWR.t1471 738.074
R8139 VPWR.n522 VPWR.t1336 738.074
R8140 VPWR.n518 VPWR.t1146 738.074
R8141 VPWR.n514 VPWR.t801 738.074
R8142 VPWR.n510 VPWR.t832 738.074
R8143 VPWR.n506 VPWR.t840 738.074
R8144 VPWR.n502 VPWR.t519 738.074
R8145 VPWR.n498 VPWR.t1311 738.074
R8146 VPWR.n494 VPWR.t1259 738.074
R8147 VPWR.n490 VPWR.t1307 738.074
R8148 VPWR.n486 VPWR.t1359 738.074
R8149 VPWR.n483 VPWR.t599 738.074
R8150 VPWR.n526 VPWR.t391 738.074
R8151 VPWR.n548 VPWR.t1106 738.074
R8152 VPWR.n549 VPWR.t853 738.074
R8153 VPWR.n552 VPWR.t1710 738.074
R8154 VPWR.n553 VPWR.t1447 738.074
R8155 VPWR.n557 VPWR.t1696 738.074
R8156 VPWR.n560 VPWR.t912 738.074
R8157 VPWR.n561 VPWR.t483 738.074
R8158 VPWR.n564 VPWR.t887 738.074
R8159 VPWR.n565 VPWR.t885 738.074
R8160 VPWR.n568 VPWR.t724 738.074
R8161 VPWR.n569 VPWR.t1175 738.074
R8162 VPWR.n572 VPWR.t1829 738.074
R8163 VPWR.n573 VPWR.t1917 738.074
R8164 VPWR.n576 VPWR.t565 738.074
R8165 VPWR.n577 VPWR.t781 738.074
R8166 VPWR.n556 VPWR.t1275 738.074
R8167 VPWR.n579 VPWR.t1114 738.074
R8168 VPWR.n583 VPWR.t1019 738.074
R8169 VPWR.n587 VPWR.t472 738.074
R8170 VPWR.n591 VPWR.t1461 738.074
R8171 VPWR.n599 VPWR.t1546 738.074
R8172 VPWR.n603 VPWR.t1156 738.074
R8173 VPWR.n607 VPWR.t811 738.074
R8174 VPWR.n611 VPWR.t933 738.074
R8175 VPWR.n615 VPWR.t946 738.074
R8176 VPWR.n619 VPWR.t1235 738.074
R8177 VPWR.n623 VPWR.t1321 738.074
R8178 VPWR.n627 VPWR.t1249 738.074
R8179 VPWR.n631 VPWR.t1716 738.074
R8180 VPWR.n635 VPWR.t736 738.074
R8181 VPWR.n578 VPWR.t605 738.074
R8182 VPWR.n595 VPWR.t397 738.074
R8183 VPWR.n673 VPWR.t1126 738.074
R8184 VPWR.n672 VPWR.t825 738.074
R8185 VPWR.n669 VPWR.t1552 738.074
R8186 VPWR.n668 VPWR.t1483 738.074
R8187 VPWR.n664 VPWR.t1330 738.074
R8188 VPWR.n661 VPWR.t621 738.074
R8189 VPWR.n660 VPWR.t1590 738.074
R8190 VPWR.n657 VPWR.t872 738.074
R8191 VPWR.n656 VPWR.t545 738.074
R8192 VPWR.n653 VPWR.t507 738.074
R8193 VPWR.n652 VPWR.t1665 738.074
R8194 VPWR.n649 VPWR.t1283 738.074
R8195 VPWR.n648 VPWR.t1297 738.074
R8196 VPWR.n645 VPWR.t1497 738.074
R8197 VPWR.n644 VPWR.t523 738.074
R8198 VPWR.n665 VPWR.t999 738.074
R8199 VPWR.n674 VPWR.t1133 738.074
R8200 VPWR.n730 VPWR.t1190 738.074
R8201 VPWR.n726 VPWR.t688 738.074
R8202 VPWR.n722 VPWR.t1495 738.074
R8203 VPWR.n714 VPWR.t1594 738.074
R8204 VPWR.n710 VPWR.t958 738.074
R8205 VPWR.n706 VPWR.t1578 738.074
R8206 VPWR.n702 VPWR.t899 738.074
R8207 VPWR.n698 VPWR.t1683 738.074
R8208 VPWR.n694 VPWR.t744 738.074
R8209 VPWR.n690 VPWR.t1620 738.074
R8210 VPWR.n686 VPWR.t1572 738.074
R8211 VPWR.n682 VPWR.t1076 738.074
R8212 VPWR.n678 VPWR.t411 738.074
R8213 VPWR.n675 VPWR.t1845 738.074
R8214 VPWR.n718 VPWR.t1507 738.074
R8215 VPWR.n740 VPWR.t1129 738.074
R8216 VPWR.n741 VPWR.t1013 738.074
R8217 VPWR.n744 VPWR.t1029 738.074
R8218 VPWR.n745 VPWR.t1489 738.074
R8219 VPWR.n749 VPWR.t1626 738.074
R8220 VPWR.n752 VPWR.t655 738.074
R8221 VPWR.n753 VPWR.t1586 738.074
R8222 VPWR.n756 VPWR.t665 738.074
R8223 VPWR.n757 VPWR.t1035 738.074
R8224 VPWR.n760 VPWR.t752 738.074
R8225 VPWR.n761 VPWR.t879 738.074
R8226 VPWR.n764 VPWR.t1568 738.074
R8227 VPWR.n765 VPWR.t1080 738.074
R8228 VPWR.n768 VPWR.t419 738.074
R8229 VPWR.n769 VPWR.t1849 738.074
R8230 VPWR.n748 VPWR.t1511 738.074
R8231 VPWR.n771 VPWR.t1108 738.074
R8232 VPWR.n775 VPWR.t434 738.074
R8233 VPWR.n779 VPWR.t1708 738.074
R8234 VPWR.n783 VPWR.t1449 738.074
R8235 VPWR.n791 VPWR.t1694 738.074
R8236 VPWR.n795 VPWR.t910 738.074
R8237 VPWR.n799 VPWR.t481 738.074
R8238 VPWR.n803 VPWR.t649 738.074
R8239 VPWR.n807 VPWR.t883 738.074
R8240 VPWR.n811 VPWR.t722 738.074
R8241 VPWR.n815 VPWR.t1173 738.074
R8242 VPWR.n819 VPWR.t537 738.074
R8243 VPWR.n823 VPWR.t1913 738.074
R8244 VPWR.n827 VPWR.t563 738.074
R8245 VPWR.n770 VPWR.t777 738.074
R8246 VPWR.n787 VPWR.t1271 738.074
R8247 VPWR.n865 VPWR.t1124 738.074
R8248 VPWR.n864 VPWR.t827 738.074
R8249 VPWR.n861 VPWR.t1554 738.074
R8250 VPWR.n860 VPWR.t1481 738.074
R8251 VPWR.n856 VPWR.t1332 738.074
R8252 VPWR.n853 VPWR.t623 738.074
R8253 VPWR.n852 VPWR.t791 738.074
R8254 VPWR.n849 VPWR.t874 738.074
R8255 VPWR.n848 VPWR.t547 738.074
R8256 VPWR.n845 VPWR.t509 738.074
R8257 VPWR.n844 VPWR.t1667 738.074
R8258 VPWR.n841 VPWR.t1285 738.074
R8259 VPWR.n840 VPWR.t1299 738.074
R8260 VPWR.n837 VPWR.t1499 738.074
R8261 VPWR.n836 VPWR.t525 738.074
R8262 VPWR.n857 VPWR.t1391 738.074
R8263 VPWR.n866 VPWR.t1110 738.074
R8264 VPWR.n922 VPWR.t432 738.074
R8265 VPWR.n918 VPWR.t1706 738.074
R8266 VPWR.n914 VPWR.t1451 738.074
R8267 VPWR.n906 VPWR.t1673 738.074
R8268 VPWR.n902 VPWR.t908 738.074
R8269 VPWR.n898 VPWR.t479 738.074
R8270 VPWR.n894 VPWR.t645 738.074
R8271 VPWR.n890 VPWR.t881 738.074
R8272 VPWR.n886 VPWR.t720 738.074
R8273 VPWR.n882 VPWR.t1171 738.074
R8274 VPWR.n878 VPWR.t535 738.074
R8275 VPWR.n874 VPWR.t1909 738.074
R8276 VPWR.n870 VPWR.t561 738.074
R8277 VPWR.n867 VPWR.t775 738.074
R8278 VPWR.n910 VPWR.t1269 738.074
R8279 VPWR.n940 VPWR.t395 738.074
R8280 VPWR.n979 VPWR.t1281 738.074
R8281 VPWR.n1179 VPWR.t66 738.074
R8282 VPWR.n399 VPWR.t1479 738.074
R8283 VPWR.n361 VPWR.t1459 738.074
R8284 VPWR.n338 VPWR.t1467 738.074
R8285 VPWR.n92 VPWR.t75 738.074
R8286 VPWR.n975 VPWR.t1441 738.074
R8287 VPWR.n1183 VPWR.t348 738.074
R8288 VPWR.n941 VPWR.t1542 738.074
R8289 VPWR.n983 VPWR.t1702 738.074
R8290 VPWR.n1217 VPWR.t78 738.074
R8291 VPWR.n407 VPWR.t1334 738.074
R8292 VPWR.n415 VPWR.t793 738.074
R8293 VPWR.n419 VPWR.t659 738.074
R8294 VPWR.n423 VPWR.t549 738.074
R8295 VPWR.n427 VPWR.t511 738.074
R8296 VPWR.n431 VPWR.t1669 738.074
R8297 VPWR.n435 VPWR.t1287 738.074
R8298 VPWR.n439 VPWR.t1301 738.074
R8299 VPWR.n443 VPWR.t1501 738.074
R8300 VPWR.n386 VPWR.t529 738.074
R8301 VPWR.n411 VPWR.t625 738.074
R8302 VPWR.n368 VPWR.t1135 738.074
R8303 VPWR.n326 VPWR.t1148 738.074
R8304 VPWR.n81 VPWR.t351 738.074
R8305 VPWR.n987 VPWR.t918 738.074
R8306 VPWR.n1214 VPWR.t237 738.074
R8307 VPWR.n944 VPWR.t1152 738.074
R8308 VPWR.n948 VPWR.t931 738.074
R8309 VPWR.n949 VPWR.t942 738.074
R8310 VPWR.n952 VPWR.t1233 738.074
R8311 VPWR.n953 VPWR.t1317 738.074
R8312 VPWR.n956 VPWR.t1247 738.074
R8313 VPWR.n957 VPWR.t1714 738.074
R8314 VPWR.n960 VPWR.t734 738.074
R8315 VPWR.n961 VPWR.t603 738.074
R8316 VPWR.n945 VPWR.t807 738.074
R8317 VPWR.n991 VPWR.t489 738.074
R8318 VPWR.n1206 VPWR.t345 738.074
R8319 VPWR.n360 VPWR.t474 738.074
R8320 VPWR.n342 VPWR.t1677 738.074
R8321 VPWR.n93 VPWR.t310 738.074
R8322 VPWR.n1180 VPWR.t183 738.074
R8323 VPWR.n995 VPWR.t891 738.074
R8324 VPWR.n1203 VPWR.t106 738.074
R8325 VPWR.n372 VPWR.t935 738.074
R8326 VPWR.n376 VPWR.t1237 738.074
R8327 VPWR.n377 VPWR.t1323 738.074
R8328 VPWR.n380 VPWR.t1251 738.074
R8329 VPWR.n381 VPWR.t1718 738.074
R8330 VPWR.n384 VPWR.t738 738.074
R8331 VPWR.n385 VPWR.t609 738.074
R8332 VPWR.n373 VPWR.t948 738.074
R8333 VPWR.n314 VPWR.t842 738.074
R8334 VPWR.n74 VPWR.t248 738.074
R8335 VPWR.n1200 VPWR.t132 738.074
R8336 VPWR.n999 VPWR.t1184 738.074
R8337 VPWR.n1003 VPWR.t726 738.074
R8338 VPWR.n1007 VPWR.t1614 738.074
R8339 VPWR.n1011 VPWR.t1831 738.074
R8340 VPWR.n1015 VPWR.t1921 738.074
R8341 VPWR.n1019 VPWR.t403 738.074
R8342 VPWR.n962 VPWR.t787 738.074
R8343 VPWR.n967 VPWR.t855 738.074
R8344 VPWR.n1123 VPWR.t81 738.074
R8345 VPWR.n310 VPWR.t1231 738.074
R8346 VPWR.n69 VPWR.t378 738.074
R8347 VPWR.n1192 VPWR.t259 738.074
R8348 VPWR.n1189 VPWR.t5 738.074
R8349 VPWR.n306 VPWR.t1313 738.074
R8350 VPWR.n302 VPWR.t1261 738.074
R8351 VPWR.n294 VPWR.t1361 738.074
R8352 VPWR.n291 VPWR.t601 738.074
R8353 VPWR.n298 VPWR.t1712 738.074
R8354 VPWR.n1058 VPWR.t264 738.074
R8355 VPWR.n1186 VPWR.t26 738.074
R8356 VPWR.n63 VPWR.t152 738.074
R8357 VPWR.n62 VPWR.t2 738.074
R8358 VPWR.n57 VPWR.t21 738.074
R8359 VPWR.n56 VPWR.t146 738.074
R8360 VPWR.n1059 VPWR.t292 738.074
R8361 VPWR.n1061 VPWR.t11 738.074
R8362 VPWR.n2856 VPWR.n2821 702.354
R8363 VPWR.n2856 VPWR.n2822 702.354
R8364 VPWR.n2854 VPWR.n2853 702.354
R8365 VPWR.n2854 VPWR.n2821 702.354
R8366 VPWR.n2837 VPWR.n2828 702.354
R8367 VPWR.n2850 VPWR.n2849 702.354
R8368 VPWR.n2835 VPWR.n2828 702.354
R8369 VPWR.n2815 VPWR.t1042 651.634
R8370 VPWR.n2831 VPWR.t1127 651.505
R8371 VPWR.n2825 VPWR.t571 651.505
R8372 VPWR.n2862 VPWR.t1404 651.431
R8373 VPWR.n1061 VPWR.t135 646.071
R8374 VPWR.n1122 VPWR.t31 646.071
R8375 VPWR.n1059 VPWR.t284 646.071
R8376 VPWR.n56 VPWR.t251 646.071
R8377 VPWR.n62 VPWR.t375 646.071
R8378 VPWR.n99 VPWR.t160 646.071
R8379 VPWR.n1053 VPWR.t1074 646.071
R8380 VPWR.n1231 VPWR.t430 646.071
R8381 VPWR.n298 VPWR.t742 646.071
R8382 VPWR.n290 VPWR.t1025 646.071
R8383 VPWR.n306 VPWR.t1255 646.071
R8384 VPWR.n68 VPWR.t114 646.071
R8385 VPWR.n1153 VPWR.t1346 646.071
R8386 VPWR.n346 VPWR.t470 646.071
R8387 VPWR.n98 VPWR.t289 646.071
R8388 VPWR.n967 VPWR.t1905 646.071
R8389 VPWR.n963 VPWR.t1194 646.071
R8390 VPWR.n999 VPWR.t748 646.071
R8391 VPWR.n373 VPWR.t1871 646.071
R8392 VPWR.n356 VPWR.t1200 646.071
R8393 VPWR.n357 VPWR.t1562 646.071
R8394 VPWR.n372 VPWR.t555 646.071
R8395 VPWR.n318 VPWR.t944 646.071
R8396 VPWR.n75 VPWR.t219 646.071
R8397 VPWR.n971 VPWR.t1477 646.071
R8398 VPWR.n369 VPWR.t895 646.071
R8399 VPWR.n322 VPWR.t651 646.071
R8400 VPWR.n80 VPWR.t91 646.071
R8401 VPWR.n945 VPWR.t889 646.071
R8402 VPWR.n932 VPWR.t1196 646.071
R8403 VPWR.n933 VPWR.t476 646.071
R8404 VPWR.n936 VPWR.t1439 646.071
R8405 VPWR.n944 VPWR.t815 646.071
R8406 VPWR.n411 VPWR.t799 646.071
R8407 VPWR.n387 VPWR.t974 646.071
R8408 VPWR.n391 VPWR.t838 646.071
R8409 VPWR.n395 VPWR.t1453 646.071
R8410 VPWR.n407 VPWR.t631 646.071
R8411 VPWR.n365 VPWR.t1141 646.071
R8412 VPWR.n330 VPWR.t1154 646.071
R8413 VPWR.n86 VPWR.t332 646.071
R8414 VPWR.n937 VPWR.t1273 646.071
R8415 VPWR.n403 VPWR.t1640 646.071
R8416 VPWR.n364 VPWR.t589 646.071
R8417 VPWR.n334 VPWR.t1544 646.071
R8418 VPWR.n87 VPWR.t177 646.071
R8419 VPWR.n473 VPWR.t1624 646.071
R8420 VPWR.n481 VPWR.t1015 646.071
R8421 VPWR.n480 VPWR.t1027 646.071
R8422 VPWR.n477 VPWR.t1473 646.071
R8423 VPWR.n476 VPWR.t1397 646.071
R8424 VPWR.n472 VPWR.t653 646.071
R8425 VPWR.n469 VPWR.t1584 646.071
R8426 VPWR.n468 VPWR.t663 646.071
R8427 VPWR.n465 VPWR.t1033 646.071
R8428 VPWR.n464 VPWR.t754 646.071
R8429 VPWR.n461 VPWR.t1610 646.071
R8430 VPWR.n460 VPWR.t1570 646.071
R8431 VPWR.n457 VPWR.t1305 646.071
R8432 VPWR.n456 VPWR.t1880 646.071
R8433 VPWR.n453 VPWR.t531 646.071
R8434 VPWR.n452 VPWR.t149 646.071
R8435 VPWR.n526 VPWR.t1540 646.071
R8436 VPWR.n482 VPWR.t1023 646.071
R8437 VPWR.n538 VPWR.t1679 646.071
R8438 VPWR.n534 VPWR.t1445 646.071
R8439 VPWR.n530 VPWR.t1265 646.071
R8440 VPWR.n522 VPWR.t1150 646.071
R8441 VPWR.n518 VPWR.t805 646.071
R8442 VPWR.n514 VPWR.t647 646.071
R8443 VPWR.n510 VPWR.t844 646.071
R8444 VPWR.n506 VPWR.t1239 646.071
R8445 VPWR.n502 VPWR.t1315 646.071
R8446 VPWR.n498 VPWR.t1253 646.071
R8447 VPWR.n494 VPWR.t1911 646.071
R8448 VPWR.n490 VPWR.t740 646.071
R8449 VPWR.n486 VPWR.t771 646.071
R8450 VPWR.n483 VPWR.t367 646.071
R8451 VPWR.n556 VPWR.t1704 646.071
R8452 VPWR.n548 VPWR.t861 646.071
R8453 VPWR.n549 VPWR.t1903 646.071
R8454 VPWR.n552 VPWR.t1485 646.071
R8455 VPWR.n553 VPWR.t995 646.071
R8456 VPWR.n557 VPWR.t954 646.071
R8457 VPWR.n560 VPWR.t491 646.071
R8458 VPWR.n561 VPWR.t868 646.071
R8459 VPWR.n564 VPWR.t1186 646.071
R8460 VPWR.n565 VPWR.t732 646.071
R8461 VPWR.n568 VPWR.t1616 646.071
R8462 VPWR.n569 VPWR.t1837 646.071
R8463 VPWR.n572 VPWR.t1086 646.071
R8464 VPWR.n573 VPWR.t409 646.071
R8465 VPWR.n576 VPWR.t505 646.071
R8466 VPWR.n577 VPWR.t216 646.071
R8467 VPWR.n595 VPWR.t587 646.071
R8468 VPWR.n579 VPWR.t1198 646.071
R8469 VPWR.n583 VPWR.t1598 646.071
R8470 VPWR.n587 VPWR.t1437 646.071
R8471 VPWR.n591 VPWR.t1277 646.071
R8472 VPWR.n599 VPWR.t1139 646.071
R8473 VPWR.n603 VPWR.t817 646.071
R8474 VPWR.n607 VPWR.t893 646.071
R8475 VPWR.n611 VPWR.t952 646.071
R8476 VPWR.n615 VPWR.t1245 646.071
R8477 VPWR.n619 VPWR.t1342 646.071
R8478 VPWR.n623 VPWR.t1839 646.071
R8479 VPWR.n627 VPWR.t1923 646.071
R8480 VPWR.n631 VPWR.t760 646.071
R8481 VPWR.n635 VPWR.t783 646.071
R8482 VPWR.n578 VPWR.t324 646.071
R8483 VPWR.n665 VPWR.t1636 646.071
R8484 VPWR.n673 VPWR.t970 646.071
R8485 VPWR.n672 VPWR.t1558 646.071
R8486 VPWR.n669 VPWR.t1457 646.071
R8487 VPWR.n668 VPWR.t399 646.071
R8488 VPWR.n664 VPWR.t627 646.071
R8489 VPWR.n661 VPWR.t795 646.071
R8490 VPWR.n660 VPWR.t937 646.071
R8491 VPWR.n657 VPWR.t551 646.071
R8492 VPWR.n656 VPWR.t513 646.071
R8493 VPWR.n653 VPWR.t923 646.071
R8494 VPWR.n652 VPWR.t1353 646.071
R8495 VPWR.n649 VPWR.t1720 646.071
R8496 VPWR.n648 VPWR.t1503 646.071
R8497 VPWR.n645 VPWR.t607 646.071
R8498 VPWR.n644 VPWR.t50 646.071
R8499 VPWR.n718 VPWR.t1622 646.071
R8500 VPWR.n674 VPWR.t1011 646.071
R8501 VPWR.n730 VPWR.t692 646.071
R8502 VPWR.n726 VPWR.t1475 646.071
R8503 VPWR.n722 VPWR.t1393 646.071
R8504 VPWR.n714 VPWR.t962 646.071
R8505 VPWR.n710 VPWR.t1582 646.071
R8506 VPWR.n706 VPWR.t661 646.071
R8507 VPWR.n702 VPWR.t1687 646.071
R8508 VPWR.n698 VPWR.t750 646.071
R8509 VPWR.n694 VPWR.t1608 646.071
R8510 VPWR.n690 VPWR.t1566 646.071
R8511 VPWR.n686 VPWR.t1303 646.071
R8512 VPWR.n682 VPWR.t417 646.071
R8513 VPWR.n678 VPWR.t527 646.071
R8514 VPWR.n675 VPWR.t157 646.071
R8515 VPWR.n748 VPWR.t1628 646.071
R8516 VPWR.n740 VPWR.t823 646.071
R8517 VPWR.n741 VPWR.t1031 646.071
R8518 VPWR.n744 VPWR.t1465 646.071
R8519 VPWR.n745 VPWR.t389 646.071
R8520 VPWR.n749 VPWR.t657 646.071
R8521 VPWR.n752 VPWR.t1588 646.071
R8522 VPWR.n753 VPWR.t834 646.071
R8523 VPWR.n756 VPWR.t1037 646.071
R8524 VPWR.n757 VPWR.t756 646.071
R8525 VPWR.n760 VPWR.t1663 646.071
R8526 VPWR.n761 VPWR.t1533 646.071
R8527 VPWR.n764 VPWR.t1309 646.071
R8528 VPWR.n765 VPWR.t1882 646.071
R8529 VPWR.n768 VPWR.t533 646.071
R8530 VPWR.n769 VPWR.t117 646.071
R8531 VPWR.n787 VPWR.t1700 646.071
R8532 VPWR.n771 VPWR.t859 646.071
R8533 VPWR.n775 VPWR.t1899 646.071
R8534 VPWR.n779 VPWR.t1469 646.071
R8535 VPWR.n783 VPWR.t993 646.071
R8536 VPWR.n791 VPWR.t916 646.071
R8537 VPWR.n795 VPWR.t487 646.071
R8538 VPWR.n799 VPWR.t669 646.071
R8539 VPWR.n803 VPWR.t1182 646.071
R8540 VPWR.n807 VPWR.t730 646.071
R8541 VPWR.n811 VPWR.t1612 646.071
R8542 VPWR.n815 VPWR.t1835 646.071
R8543 VPWR.n819 VPWR.t1084 646.071
R8544 VPWR.n823 VPWR.t407 646.071
R8545 VPWR.n827 VPWR.t1853 646.071
R8546 VPWR.n770 VPWR.t222 646.071
R8547 VPWR.n857 VPWR.t1638 646.071
R8548 VPWR.n865 VPWR.t972 646.071
R8549 VPWR.n864 VPWR.t1560 646.071
R8550 VPWR.n861 VPWR.t1455 646.071
R8551 VPWR.n860 VPWR.t1517 646.071
R8552 VPWR.n856 VPWR.t629 646.071
R8553 VPWR.n853 VPWR.t797 646.071
R8554 VPWR.n852 VPWR.t939 646.071
R8555 VPWR.n849 VPWR.t553 646.071
R8556 VPWR.n848 VPWR.t515 646.071
R8557 VPWR.n845 VPWR.t925 646.071
R8558 VPWR.n844 VPWR.t1355 646.071
R8559 VPWR.n841 VPWR.t1722 646.071
R8560 VPWR.n840 VPWR.t1371 646.071
R8561 VPWR.n837 VPWR.t611 646.071
R8562 VPWR.n836 VPWR.t45 646.071
R8563 VPWR.n910 VPWR.t1698 646.071
R8564 VPWR.n866 VPWR.t857 646.071
R8565 VPWR.n922 VPWR.t1897 646.071
R8566 VPWR.n918 VPWR.t1487 646.071
R8567 VPWR.n914 VPWR.t1513 646.071
R8568 VPWR.n906 VPWR.t914 646.071
R8569 VPWR.n902 VPWR.t485 646.071
R8570 VPWR.n898 VPWR.t667 646.071
R8571 VPWR.n894 VPWR.t1180 646.071
R8572 VPWR.n890 VPWR.t728 646.071
R8573 VPWR.n886 VPWR.t1177 646.071
R8574 VPWR.n882 VPWR.t1833 646.071
R8575 VPWR.n878 VPWR.t1082 646.071
R8576 VPWR.n874 VPWR.t405 646.071
R8577 VPWR.n870 VPWR.t1851 646.071
R8578 VPWR.n867 VPWR.t229 646.071
R8579 VPWR.n940 VPWR.t1550 646.071
R8580 VPWR.n979 VPWR.t1592 646.071
R8581 VPWR.n1227 VPWR.t591 646.071
R8582 VPWR.n1179 VPWR.t61 646.071
R8583 VPWR.n399 VPWR.t1519 646.071
R8584 VPWR.n361 VPWR.t1279 646.071
R8585 VPWR.n338 VPWR.t1267 646.071
R8586 VPWR.n92 VPWR.t69 646.071
R8587 VPWR.n975 VPWR.t997 646.071
R8588 VPWR.n1485 VPWR.t1505 646.071
R8589 VPWR.n1183 VPWR.t340 646.071
R8590 VPWR.n941 VPWR.t1137 646.071
R8591 VPWR.n983 VPWR.t956 646.071
R8592 VPWR.n1173 VPWR.t1143 646.071
R8593 VPWR.n1217 VPWR.t208 646.071
R8594 VPWR.n415 VPWR.t401 646.071
R8595 VPWR.n419 VPWR.t700 646.071
R8596 VPWR.n423 VPWR.t517 646.071
R8597 VPWR.n427 VPWR.t927 646.071
R8598 VPWR.n431 VPWR.t1357 646.071
R8599 VPWR.n435 VPWR.t1724 646.071
R8600 VPWR.n439 VPWR.t1373 646.071
R8601 VPWR.n443 VPWR.t613 646.071
R8602 VPWR.n386 VPWR.t37 646.071
R8603 VPWR.n368 VPWR.t819 646.071
R8604 VPWR.n326 VPWR.t809 646.071
R8605 VPWR.n81 VPWR.t56 646.071
R8606 VPWR.n987 VPWR.t493 646.071
R8607 VPWR.n1169 VPWR.t821 646.071
R8608 VPWR.n1214 VPWR.t319 646.071
R8609 VPWR.n948 VPWR.t950 646.071
R8610 VPWR.n949 VPWR.t1243 646.071
R8611 VPWR.n952 VPWR.t1340 646.071
R8612 VPWR.n953 VPWR.t1257 646.071
R8613 VPWR.n956 VPWR.t1919 646.071
R8614 VPWR.n957 VPWR.t758 646.071
R8615 VPWR.n960 VPWR.t779 646.071
R8616 VPWR.n961 VPWR.t337 646.071
R8617 VPWR.n991 VPWR.t870 646.071
R8618 VPWR.n1163 VPWR.t897 646.071
R8619 VPWR.n1206 VPWR.t356 646.071
R8620 VPWR.n360 VPWR.t1435 646.071
R8621 VPWR.n342 VPWR.t1443 646.071
R8622 VPWR.n93 VPWR.t307 646.071
R8623 VPWR.n1479 VPWR.t1491 646.071
R8624 VPWR.n1180 VPWR.t180 646.071
R8625 VPWR.n995 VPWR.t1188 646.071
R8626 VPWR.n1159 VPWR.t557 646.071
R8627 VPWR.n1203 VPWR.t101 646.071
R8628 VPWR.n376 VPWR.t1344 646.071
R8629 VPWR.n377 VPWR.t1841 646.071
R8630 VPWR.n380 VPWR.t1925 646.071
R8631 VPWR.n381 VPWR.t762 646.071
R8632 VPWR.n384 VPWR.t785 646.071
R8633 VPWR.n385 VPWR.t316 646.071
R8634 VPWR.n314 VPWR.t1241 646.071
R8635 VPWR.n74 VPWR.t329 646.071
R8636 VPWR.n1149 VPWR.t1873 646.071
R8637 VPWR.n1200 VPWR.t205 646.071
R8638 VPWR.n1003 VPWR.t1618 646.071
R8639 VPWR.n1007 VPWR.t1576 646.071
R8640 VPWR.n1011 VPWR.t1295 646.071
R8641 VPWR.n1015 VPWR.t415 646.071
R8642 VPWR.n1019 VPWR.t521 646.071
R8643 VPWR.n962 VPWR.t189 646.071
R8644 VPWR.n1472 VPWR.t1564 646.071
R8645 VPWR.n1123 VPWR.t167 646.071
R8646 VPWR.n310 VPWR.t1319 646.071
R8647 VPWR.n69 VPWR.t96 646.071
R8648 VPWR.n1192 VPWR.t364 646.071
R8649 VPWR.n1049 VPWR.t1843 646.071
R8650 VPWR.n1189 VPWR.t383 646.071
R8651 VPWR.n302 VPWR.t1915 646.071
R8652 VPWR.n294 VPWR.t773 646.071
R8653 VPWR.n291 VPWR.t359 646.071
R8654 VPWR.n1058 VPWR.t256 646.071
R8655 VPWR.n1748 VPWR.t686 646.071
R8656 VPWR.n1036 VPWR.t789 646.071
R8657 VPWR.n1032 VPWR.t300 646.071
R8658 VPWR.n1186 VPWR.t127 646.071
R8659 VPWR.n63 VPWR.t242 646.071
R8660 VPWR.n57 VPWR.t8 646.071
R8661 VPWR.n1230 VPWR.t109 642.13
R8662 VPWR.n1152 VPWR.t40 642.13
R8663 VPWR.n1226 VPWR.t245 642.13
R8664 VPWR.n1484 VPWR.t143 642.13
R8665 VPWR.n1172 VPWR.t267 642.13
R8666 VPWR.n1168 VPWR.t18 642.13
R8667 VPWR.n1162 VPWR.t140 642.13
R8668 VPWR.n1478 VPWR.t372 642.13
R8669 VPWR.n1158 VPWR.t281 642.13
R8670 VPWR.n1148 VPWR.t297 642.13
R8671 VPWR.n1471 VPWR.t270 642.13
R8672 VPWR.n1048 VPWR.t170 642.13
R8673 VPWR.n1747 VPWR.t34 642.13
R8674 VPWR.n1035 VPWR.t84 642.13
R8675 VPWR.n1031 VPWR.t192 642.13
R8676 VPWR.n1052 VPWR.t211 642.13
R8677 VPWR.n2309 VPWR.t1014 629.652
R8678 VPWR.n2310 VPWR.t1026 629.652
R8679 VPWR.n2319 VPWR.t1472 629.652
R8680 VPWR.n2320 VPWR.t1396 629.652
R8681 VPWR.n2329 VPWR.t1623 629.652
R8682 VPWR.n2330 VPWR.t652 629.652
R8683 VPWR.n2339 VPWR.t1583 629.652
R8684 VPWR.n2340 VPWR.t662 629.652
R8685 VPWR.n2349 VPWR.t1032 629.652
R8686 VPWR.n2350 VPWR.t753 629.652
R8687 VPWR.n2359 VPWR.t1609 629.652
R8688 VPWR.n2360 VPWR.t1569 629.652
R8689 VPWR.n2369 VPWR.t1304 629.652
R8690 VPWR.n2370 VPWR.t1879 629.652
R8691 VPWR.n2379 VPWR.t530 629.652
R8692 VPWR.n542 VPWR.t1022 629.652
R8693 VPWR.t1678 VPWR.n541 629.652
R8694 VPWR.t1444 VPWR.n537 629.652
R8695 VPWR.t1264 VPWR.n533 629.652
R8696 VPWR.t1539 VPWR.n529 629.652
R8697 VPWR.t1149 VPWR.n525 629.652
R8698 VPWR.t804 VPWR.n521 629.652
R8699 VPWR.t646 VPWR.n517 629.652
R8700 VPWR.t843 VPWR.n513 629.652
R8701 VPWR.t1238 VPWR.n509 629.652
R8702 VPWR.t1314 VPWR.n505 629.652
R8703 VPWR.t1252 VPWR.n501 629.652
R8704 VPWR.t1910 VPWR.n497 629.652
R8705 VPWR.t739 VPWR.n493 629.652
R8706 VPWR.t770 VPWR.n489 629.652
R8707 VPWR.n2281 VPWR.t860 629.652
R8708 VPWR.t1902 VPWR.n2280 629.652
R8709 VPWR.n2271 VPWR.t1484 629.652
R8710 VPWR.t994 VPWR.n2270 629.652
R8711 VPWR.n2261 VPWR.t1703 629.652
R8712 VPWR.t953 VPWR.n2260 629.652
R8713 VPWR.n2251 VPWR.t490 629.652
R8714 VPWR.t867 VPWR.n2250 629.652
R8715 VPWR.n2241 VPWR.t1185 629.652
R8716 VPWR.t731 VPWR.n2240 629.652
R8717 VPWR.n2231 VPWR.t1615 629.652
R8718 VPWR.t1836 VPWR.n2230 629.652
R8719 VPWR.n2221 VPWR.t1085 629.652
R8720 VPWR.t408 VPWR.n2220 629.652
R8721 VPWR.n2211 VPWR.t504 629.652
R8722 VPWR.n582 VPWR.t1197 629.652
R8723 VPWR.n586 VPWR.t1597 629.652
R8724 VPWR.n590 VPWR.t1436 629.652
R8725 VPWR.n594 VPWR.t1276 629.652
R8726 VPWR.n598 VPWR.t586 629.652
R8727 VPWR.n602 VPWR.t1138 629.652
R8728 VPWR.n606 VPWR.t816 629.652
R8729 VPWR.n610 VPWR.t892 629.652
R8730 VPWR.n614 VPWR.t951 629.652
R8731 VPWR.n618 VPWR.t1244 629.652
R8732 VPWR.n622 VPWR.t1341 629.652
R8733 VPWR.n626 VPWR.t1838 629.652
R8734 VPWR.n630 VPWR.t1922 629.652
R8735 VPWR.n634 VPWR.t759 629.652
R8736 VPWR.n638 VPWR.t782 629.652
R8737 VPWR.n2113 VPWR.t969 629.652
R8738 VPWR.n2114 VPWR.t1557 629.652
R8739 VPWR.n2123 VPWR.t1456 629.652
R8740 VPWR.n2124 VPWR.t398 629.652
R8741 VPWR.n2133 VPWR.t1635 629.652
R8742 VPWR.n2134 VPWR.t626 629.652
R8743 VPWR.n2143 VPWR.t794 629.652
R8744 VPWR.n2144 VPWR.t936 629.652
R8745 VPWR.n2153 VPWR.t550 629.652
R8746 VPWR.n2154 VPWR.t512 629.652
R8747 VPWR.n2163 VPWR.t922 629.652
R8748 VPWR.n2164 VPWR.t1352 629.652
R8749 VPWR.n2173 VPWR.t1719 629.652
R8750 VPWR.n2174 VPWR.t1502 629.652
R8751 VPWR.n2183 VPWR.t606 629.652
R8752 VPWR.n734 VPWR.t1010 629.652
R8753 VPWR.t691 VPWR.n733 629.652
R8754 VPWR.t1474 VPWR.n729 629.652
R8755 VPWR.t1392 VPWR.n725 629.652
R8756 VPWR.t1621 VPWR.n721 629.652
R8757 VPWR.t961 VPWR.n717 629.652
R8758 VPWR.t1581 VPWR.n713 629.652
R8759 VPWR.t660 VPWR.n709 629.652
R8760 VPWR.t1686 VPWR.n705 629.652
R8761 VPWR.t749 VPWR.n701 629.652
R8762 VPWR.t1607 VPWR.n697 629.652
R8763 VPWR.t1565 VPWR.n693 629.652
R8764 VPWR.t1302 VPWR.n689 629.652
R8765 VPWR.t416 VPWR.n685 629.652
R8766 VPWR.t526 VPWR.n681 629.652
R8767 VPWR.n2085 VPWR.t822 629.652
R8768 VPWR.t1030 VPWR.n2084 629.652
R8769 VPWR.n2075 VPWR.t1464 629.652
R8770 VPWR.t388 VPWR.n2074 629.652
R8771 VPWR.n2065 VPWR.t1627 629.652
R8772 VPWR.t656 VPWR.n2064 629.652
R8773 VPWR.n2055 VPWR.t1587 629.652
R8774 VPWR.t833 VPWR.n2054 629.652
R8775 VPWR.n2045 VPWR.t1036 629.652
R8776 VPWR.t755 VPWR.n2044 629.652
R8777 VPWR.n2035 VPWR.t1662 629.652
R8778 VPWR.t1532 VPWR.n2034 629.652
R8779 VPWR.n2025 VPWR.t1308 629.652
R8780 VPWR.t1881 VPWR.n2024 629.652
R8781 VPWR.n2015 VPWR.t532 629.652
R8782 VPWR.n774 VPWR.t858 629.652
R8783 VPWR.n778 VPWR.t1898 629.652
R8784 VPWR.n782 VPWR.t1468 629.652
R8785 VPWR.n786 VPWR.t992 629.652
R8786 VPWR.n790 VPWR.t1699 629.652
R8787 VPWR.n794 VPWR.t915 629.652
R8788 VPWR.n798 VPWR.t486 629.652
R8789 VPWR.n802 VPWR.t668 629.652
R8790 VPWR.n806 VPWR.t1181 629.652
R8791 VPWR.n810 VPWR.t729 629.652
R8792 VPWR.n814 VPWR.t1611 629.652
R8793 VPWR.n818 VPWR.t1834 629.652
R8794 VPWR.n822 VPWR.t1083 629.652
R8795 VPWR.n826 VPWR.t406 629.652
R8796 VPWR.n830 VPWR.t1852 629.652
R8797 VPWR.n1917 VPWR.t971 629.652
R8798 VPWR.n1918 VPWR.t1559 629.652
R8799 VPWR.n1927 VPWR.t1454 629.652
R8800 VPWR.n1928 VPWR.t1516 629.652
R8801 VPWR.n1937 VPWR.t1637 629.652
R8802 VPWR.n1938 VPWR.t628 629.652
R8803 VPWR.n1947 VPWR.t796 629.652
R8804 VPWR.n1948 VPWR.t938 629.652
R8805 VPWR.n1957 VPWR.t552 629.652
R8806 VPWR.n1958 VPWR.t514 629.652
R8807 VPWR.n1967 VPWR.t924 629.652
R8808 VPWR.n1968 VPWR.t1354 629.652
R8809 VPWR.n1977 VPWR.t1721 629.652
R8810 VPWR.n1978 VPWR.t1370 629.652
R8811 VPWR.n1987 VPWR.t610 629.652
R8812 VPWR.n926 VPWR.t856 629.652
R8813 VPWR.t1896 VPWR.n925 629.652
R8814 VPWR.t1486 VPWR.n921 629.652
R8815 VPWR.t1512 VPWR.n917 629.652
R8816 VPWR.t1697 VPWR.n913 629.652
R8817 VPWR.t913 VPWR.n909 629.652
R8818 VPWR.t484 VPWR.n905 629.652
R8819 VPWR.t666 VPWR.n901 629.652
R8820 VPWR.t1179 VPWR.n897 629.652
R8821 VPWR.t727 VPWR.n893 629.652
R8822 VPWR.t1176 VPWR.n889 629.652
R8823 VPWR.t1832 VPWR.n885 629.652
R8824 VPWR.t1081 VPWR.n881 629.652
R8825 VPWR.t404 VPWR.n877 629.652
R8826 VPWR.t1850 VPWR.n873 629.652
R8827 VPWR.n390 VPWR.t973 629.652
R8828 VPWR.n394 VPWR.t837 629.652
R8829 VPWR.n398 VPWR.t1452 629.652
R8830 VPWR.n402 VPWR.t1518 629.652
R8831 VPWR.n406 VPWR.t1639 629.652
R8832 VPWR.n410 VPWR.t630 629.652
R8833 VPWR.n414 VPWR.t798 629.652
R8834 VPWR.n418 VPWR.t400 629.652
R8835 VPWR.n422 VPWR.t699 629.652
R8836 VPWR.n426 VPWR.t516 629.652
R8837 VPWR.n430 VPWR.t926 629.652
R8838 VPWR.n434 VPWR.t1356 629.652
R8839 VPWR.n438 VPWR.t1723 629.652
R8840 VPWR.n442 VPWR.t1372 629.652
R8841 VPWR.n446 VPWR.t612 629.652
R8842 VPWR.n1889 VPWR.t1195 629.652
R8843 VPWR.t475 VPWR.n1888 629.652
R8844 VPWR.n1879 VPWR.t1438 629.652
R8845 VPWR.t1272 VPWR.n1878 629.652
R8846 VPWR.n1869 VPWR.t1549 629.652
R8847 VPWR.t1136 VPWR.n1868 629.652
R8848 VPWR.n1859 VPWR.t814 629.652
R8849 VPWR.t888 VPWR.n1858 629.652
R8850 VPWR.n1849 VPWR.t949 629.652
R8851 VPWR.t1242 VPWR.n1848 629.652
R8852 VPWR.n1839 VPWR.t1339 629.652
R8853 VPWR.t1256 VPWR.n1838 629.652
R8854 VPWR.n1829 VPWR.t1918 629.652
R8855 VPWR.t757 VPWR.n1828 629.652
R8856 VPWR.n1819 VPWR.t778 629.652
R8857 VPWR.n2477 VPWR.t1199 629.652
R8858 VPWR.t1561 VPWR.n2476 629.652
R8859 VPWR.n2467 VPWR.t1434 629.652
R8860 VPWR.t1278 VPWR.n2466 629.652
R8861 VPWR.n2457 VPWR.t588 629.652
R8862 VPWR.t1140 VPWR.n2456 629.652
R8863 VPWR.n2447 VPWR.t818 629.652
R8864 VPWR.t894 VPWR.n2446 629.652
R8865 VPWR.n2437 VPWR.t554 629.652
R8866 VPWR.t1870 VPWR.n2436 629.652
R8867 VPWR.n2427 VPWR.t1343 629.652
R8868 VPWR.t1840 VPWR.n2426 629.652
R8869 VPWR.n2417 VPWR.t1924 629.652
R8870 VPWR.t761 VPWR.n2416 629.652
R8871 VPWR.n2407 VPWR.t784 629.652
R8872 VPWR.n966 VPWR.t1193 629.652
R8873 VPWR.n970 VPWR.t1904 629.652
R8874 VPWR.n974 VPWR.t1476 629.652
R8875 VPWR.n978 VPWR.t996 629.652
R8876 VPWR.n982 VPWR.t1591 629.652
R8877 VPWR.n986 VPWR.t955 629.652
R8878 VPWR.n990 VPWR.t492 629.652
R8879 VPWR.n994 VPWR.t869 629.652
R8880 VPWR.n998 VPWR.t1187 629.652
R8881 VPWR.n1002 VPWR.t747 629.652
R8882 VPWR.n1006 VPWR.t1617 629.652
R8883 VPWR.n1010 VPWR.t1575 629.652
R8884 VPWR.n1014 VPWR.t1294 629.652
R8885 VPWR.n1018 VPWR.t414 629.652
R8886 VPWR.n1022 VPWR.t520 629.652
R8887 VPWR.n350 VPWR.t1024 629.652
R8888 VPWR.t469 VPWR.n349 629.652
R8889 VPWR.t1442 VPWR.n345 629.652
R8890 VPWR.t1266 VPWR.n341 629.652
R8891 VPWR.t1543 VPWR.n337 629.652
R8892 VPWR.t1153 VPWR.n333 629.652
R8893 VPWR.t808 VPWR.n329 629.652
R8894 VPWR.t650 VPWR.n325 629.652
R8895 VPWR.t943 VPWR.n321 629.652
R8896 VPWR.t1240 VPWR.n317 629.652
R8897 VPWR.t1318 VPWR.n313 629.652
R8898 VPWR.t1254 VPWR.n309 629.652
R8899 VPWR.t1914 VPWR.n305 629.652
R8900 VPWR.t741 VPWR.n301 629.652
R8901 VPWR.t772 VPWR.n297 629.652
R8902 VPWR.n1468 VPWR.t429 629.652
R8903 VPWR.n1475 VPWR.t1563 629.652
R8904 VPWR.n1481 VPWR.t1490 629.652
R8905 VPWR.n1492 VPWR.t1504 629.652
R8906 VPWR.n1493 VPWR.t590 629.652
R8907 VPWR.n1506 VPWR.t1142 629.652
R8908 VPWR.n1507 VPWR.t820 629.652
R8909 VPWR.n1520 VPWR.t896 629.652
R8910 VPWR.n1521 VPWR.t556 629.652
R8911 VPWR.n1536 VPWR.t1872 629.652
R8912 VPWR.t1345 VPWR.n1535 629.652
R8913 VPWR.n1761 VPWR.t1842 629.652
R8914 VPWR.t1073 VPWR.n1760 629.652
R8915 VPWR.n1749 VPWR.t685 629.652
R8916 VPWR.n1791 VPWR.t788 629.652
R8917 VPWR.n2506 VPWR.t159 629.652
R8918 VPWR.n2507 VPWR.t288 629.652
R8919 VPWR.n2518 VPWR.t306 629.652
R8920 VPWR.n2519 VPWR.t68 629.652
R8921 VPWR.n2530 VPWR.t176 629.652
R8922 VPWR.n2531 VPWR.t331 629.652
R8923 VPWR.n2542 VPWR.t55 629.652
R8924 VPWR.n2543 VPWR.t90 629.652
R8925 VPWR.n2554 VPWR.t218 629.652
R8926 VPWR.n2555 VPWR.t328 629.652
R8927 VPWR.n2566 VPWR.t95 629.652
R8928 VPWR.n2567 VPWR.t113 629.652
R8929 VPWR.n2578 VPWR.t241 629.652
R8930 VPWR.n2579 VPWR.t374 629.652
R8931 VPWR.n2590 VPWR.t7 629.652
R8932 VPWR.n1594 VPWR.t30 629.652
R8933 VPWR.t166 VPWR.n1593 629.652
R8934 VPWR.n1182 VPWR.t179 629.652
R8935 VPWR.n1185 VPWR.t339 629.652
R8936 VPWR.n1220 VPWR.t60 629.652
R8937 VPWR.t207 VPWR.n1219 629.652
R8938 VPWR.t318 VPWR.n1216 629.652
R8939 VPWR.t355 VPWR.n1213 629.652
R8940 VPWR.t100 VPWR.n1205 629.652
R8941 VPWR.t204 VPWR.n1202 629.652
R8942 VPWR.t363 VPWR.n1199 629.652
R8943 VPWR.t382 VPWR.n1191 629.652
R8944 VPWR.t126 VPWR.n1188 629.652
R8945 VPWR.n1740 VPWR.t255 629.652
R8946 VPWR.t283 VPWR.n1739 629.652
R8947 VPWR.n2836 VPWR.t570 531.804
R8948 VPWR.n2855 VPWR.t570 531.804
R8949 VPWR.n2851 VPWR.n2850 504.707
R8950 VPWR.t1014 VPWR.t769 486.048
R8951 VPWR.t1026 VPWR.t1731 486.048
R8952 VPWR.t1327 VPWR.t1472 486.048
R8953 VPWR.t1396 VPWR.t1326 486.048
R8954 VPWR.t768 VPWR.t1623 486.048
R8955 VPWR.t652 VPWR.t1163 486.048
R8956 VPWR.t1162 VPWR.t1583 486.048
R8957 VPWR.t662 VPWR.t767 486.048
R8958 VPWR.t1733 VPWR.t1032 486.048
R8959 VPWR.t753 VPWR.t1164 486.048
R8960 VPWR.t1325 VPWR.t1609 486.048
R8961 VPWR.t1569 VPWR.t1324 486.048
R8962 VPWR.t1161 VPWR.t1304 486.048
R8963 VPWR.t1879 VPWR.t1160 486.048
R8964 VPWR.t1328 VPWR.t530 486.048
R8965 VPWR.t148 VPWR.t1732 486.048
R8966 VPWR.t1022 VPWR.t1867 486.048
R8967 VPWR.t977 VPWR.t1678 486.048
R8968 VPWR.t1377 VPWR.t1444 486.048
R8969 VPWR.t1376 VPWR.t1264 486.048
R8970 VPWR.t1866 VPWR.t1539 486.048
R8971 VPWR.t1660 VPWR.t1149 486.048
R8972 VPWR.t1659 VPWR.t804 486.048
R8973 VPWR.t1865 VPWR.t646 486.048
R8974 VPWR.t979 VPWR.t843 486.048
R8975 VPWR.t1661 VPWR.t1238 486.048
R8976 VPWR.t1375 VPWR.t1314 486.048
R8977 VPWR.t1868 VPWR.t1252 486.048
R8978 VPWR.t1658 VPWR.t1910 486.048
R8979 VPWR.t1657 VPWR.t739 486.048
R8980 VPWR.t1378 VPWR.t770 486.048
R8981 VPWR.t978 VPWR.t366 486.048
R8982 VPWR.t860 VPWR.t1263 486.048
R8983 VPWR.t1053 VPWR.t1902 486.048
R8984 VPWR.t1484 VPWR.t1644 486.048
R8985 VPWR.t1643 VPWR.t994 486.048
R8986 VPWR.t1703 VPWR.t1262 486.048
R8987 VPWR.t1051 VPWR.t953 486.048
R8988 VPWR.t490 VPWR.t1050 486.048
R8989 VPWR.t1056 VPWR.t867 486.048
R8990 VPWR.t1185 VPWR.t1055 486.048
R8991 VPWR.t1052 VPWR.t731 486.048
R8992 VPWR.t1615 VPWR.t1642 486.048
R8993 VPWR.t1641 VPWR.t1836 486.048
R8994 VPWR.t1085 VPWR.t1049 486.048
R8995 VPWR.t1646 VPWR.t408 486.048
R8996 VPWR.t504 VPWR.t1645 486.048
R8997 VPWR.t1054 VPWR.t215 486.048
R8998 VPWR.t1197 VPWR.t1428 486.048
R8999 VPWR.t1597 VPWR.t1423 486.048
R9000 VPWR.t1436 VPWR.t698 486.048
R9001 VPWR.t1276 VPWR.t697 486.048
R9002 VPWR.t586 VPWR.t1427 486.048
R9003 VPWR.t1138 VPWR.t1878 486.048
R9004 VPWR.t816 VPWR.t1877 486.048
R9005 VPWR.t892 VPWR.t1426 486.048
R9006 VPWR.t951 VPWR.t1425 486.048
R9007 VPWR.t1244 VPWR.t1422 486.048
R9008 VPWR.t1341 VPWR.t696 486.048
R9009 VPWR.t1838 VPWR.t695 486.048
R9010 VPWR.t1922 VPWR.t1876 486.048
R9011 VPWR.t759 VPWR.t1875 486.048
R9012 VPWR.t782 VPWR.t1874 486.048
R9013 VPWR.t323 VPWR.t1424 486.048
R9014 VPWR.t969 VPWR.t1061 486.048
R9015 VPWR.t1557 VPWR.t982 486.048
R9016 VPWR.t1158 VPWR.t1456 486.048
R9017 VPWR.t398 VPWR.t1157 486.048
R9018 VPWR.t877 VPWR.t1635 486.048
R9019 VPWR.t626 VPWR.t1691 486.048
R9020 VPWR.t1690 VPWR.t794 486.048
R9021 VPWR.t936 VPWR.t876 486.048
R9022 VPWR.t875 VPWR.t550 486.048
R9023 VPWR.t512 VPWR.t1692 486.048
R9024 VPWR.t1063 VPWR.t922 486.048
R9025 VPWR.t1352 VPWR.t1062 486.048
R9026 VPWR.t1689 VPWR.t1719 486.048
R9027 VPWR.t1502 VPWR.t1688 486.048
R9028 VPWR.t1159 VPWR.t606 486.048
R9029 VPWR.t49 VPWR.t983 486.048
R9030 VPWR.t1010 VPWR.t633 486.048
R9031 VPWR.t1821 VPWR.t691 486.048
R9032 VPWR.t1350 VPWR.t1474 486.048
R9033 VPWR.t1349 VPWR.t1392 486.048
R9034 VPWR.t632 VPWR.t1621 486.048
R9035 VPWR.t1067 VPWR.t961 486.048
R9036 VPWR.t1066 VPWR.t1581 486.048
R9037 VPWR.t1144 VPWR.t660 486.048
R9038 VPWR.t1823 VPWR.t1686 486.048
R9039 VPWR.t1068 VPWR.t749 486.048
R9040 VPWR.t1348 VPWR.t1607 486.048
R9041 VPWR.t634 VPWR.t1565 486.048
R9042 VPWR.t1065 VPWR.t1302 486.048
R9043 VPWR.t1064 VPWR.t416 486.048
R9044 VPWR.t1351 VPWR.t526 486.048
R9045 VPWR.t1822 VPWR.t156 486.048
R9046 VPWR.t822 VPWR.t1629 486.048
R9047 VPWR.t1604 VPWR.t1030 486.048
R9048 VPWR.t1464 VPWR.t1633 486.048
R9049 VPWR.t1632 VPWR.t388 486.048
R9050 VPWR.t1627 VPWR.t468 486.048
R9051 VPWR.t1602 VPWR.t656 486.048
R9052 VPWR.t1587 VPWR.t1601 486.048
R9053 VPWR.t467 VPWR.t833 486.048
R9054 VPWR.t1036 VPWR.t466 486.048
R9055 VPWR.t1603 VPWR.t755 486.048
R9056 VPWR.t1662 VPWR.t1631 486.048
R9057 VPWR.t1630 VPWR.t1532 486.048
R9058 VPWR.t1308 VPWR.t1600 486.048
R9059 VPWR.t1599 VPWR.t1881 486.048
R9060 VPWR.t532 VPWR.t1634 486.048
R9061 VPWR.t465 VPWR.t116 486.048
R9062 VPWR.t858 VPWR.t707 486.048
R9063 VPWR.t1898 VPWR.t702 486.048
R9064 VPWR.t1468 VPWR.t1004 486.048
R9065 VPWR.t992 VPWR.t1003 486.048
R9066 VPWR.t1699 VPWR.t706 486.048
R9067 VPWR.t915 VPWR.t1009 486.048
R9068 VPWR.t486 VPWR.t1008 486.048
R9069 VPWR.t668 VPWR.t705 486.048
R9070 VPWR.t1181 VPWR.t704 486.048
R9071 VPWR.t729 VPWR.t701 486.048
R9072 VPWR.t1611 VPWR.t1002 486.048
R9073 VPWR.t1834 VPWR.t1001 486.048
R9074 VPWR.t1083 VPWR.t1007 486.048
R9075 VPWR.t406 VPWR.t1006 486.048
R9076 VPWR.t1852 VPWR.t1005 486.048
R9077 VPWR.t221 VPWR.t703 486.048
R9078 VPWR.t971 VPWR.t713 486.048
R9079 VPWR.t1559 VPWR.t1824 486.048
R9080 VPWR.t717 VPWR.t1454 486.048
R9081 VPWR.t1516 VPWR.t716 486.048
R9082 VPWR.t712 VPWR.t1637 486.048
R9083 VPWR.t628 VPWR.t1530 486.048
R9084 VPWR.t1529 VPWR.t796 486.048
R9085 VPWR.t938 VPWR.t1827 486.048
R9086 VPWR.t1826 VPWR.t552 486.048
R9087 VPWR.t514 VPWR.t1531 486.048
R9088 VPWR.t715 VPWR.t924 486.048
R9089 VPWR.t1354 VPWR.t714 486.048
R9090 VPWR.t1528 VPWR.t1721 486.048
R9091 VPWR.t1370 VPWR.t1527 486.048
R9092 VPWR.t718 VPWR.t610 486.048
R9093 VPWR.t44 VPWR.t1825 486.048
R9094 VPWR.t856 VPWR.t968 486.048
R9095 VPWR.t963 VPWR.t1896 486.048
R9096 VPWR.t845 VPWR.t1486 486.048
R9097 VPWR.t1861 VPWR.t1512 486.048
R9098 VPWR.t967 VPWR.t1697 486.048
R9099 VPWR.t850 VPWR.t913 486.048
R9100 VPWR.t849 VPWR.t484 486.048
R9101 VPWR.t966 VPWR.t666 486.048
R9102 VPWR.t965 VPWR.t1179 486.048
R9103 VPWR.t851 VPWR.t727 486.048
R9104 VPWR.t1860 VPWR.t1176 486.048
R9105 VPWR.t1859 VPWR.t1832 486.048
R9106 VPWR.t848 VPWR.t1081 486.048
R9107 VPWR.t847 VPWR.t404 486.048
R9108 VPWR.t846 VPWR.t1850 486.048
R9109 VPWR.t964 VPWR.t228 486.048
R9110 VPWR.t973 VPWR.t1433 486.048
R9111 VPWR.t837 VPWR.t1347 486.048
R9112 VPWR.t1452 VPWR.t1650 486.048
R9113 VPWR.t1518 VPWR.t1649 486.048
R9114 VPWR.t1639 VPWR.t1432 486.048
R9115 VPWR.t630 VPWR.t1655 486.048
R9116 VPWR.t798 VPWR.t1654 486.048
R9117 VPWR.t400 VPWR.t1431 486.048
R9118 VPWR.t699 VPWR.t1430 486.048
R9119 VPWR.t516 VPWR.t1656 486.048
R9120 VPWR.t926 VPWR.t1648 486.048
R9121 VPWR.t1356 VPWR.t1647 486.048
R9122 VPWR.t1723 VPWR.t1653 486.048
R9123 VPWR.t1372 VPWR.t1652 486.048
R9124 VPWR.t612 VPWR.t1651 486.048
R9125 VPWR.t36 VPWR.t1429 486.048
R9126 VPWR.t1195 VPWR.t539 486.048
R9127 VPWR.t1855 VPWR.t475 486.048
R9128 VPWR.t1438 VPWR.t543 486.048
R9129 VPWR.t542 VPWR.t1272 486.048
R9130 VPWR.t1549 VPWR.t538 486.048
R9131 VPWR.t906 VPWR.t1136 486.048
R9132 VPWR.t814 VPWR.t905 486.048
R9133 VPWR.t1858 VPWR.t888 486.048
R9134 VPWR.t949 VPWR.t1857 486.048
R9135 VPWR.t1854 VPWR.t1242 486.048
R9136 VPWR.t1339 VPWR.t541 486.048
R9137 VPWR.t540 VPWR.t1256 486.048
R9138 VPWR.t1918 VPWR.t904 486.048
R9139 VPWR.t903 VPWR.t757 486.048
R9140 VPWR.t778 VPWR.t902 486.048
R9141 VPWR.t1856 VPWR.t336 486.048
R9142 VPWR.t1199 VPWR.t1169 486.048
R9143 VPWR.t1221 VPWR.t1561 486.048
R9144 VPWR.t1434 VPWR.t763 486.048
R9145 VPWR.t921 VPWR.t1278 486.048
R9146 VPWR.t588 VPWR.t1168 486.048
R9147 VPWR.t1219 VPWR.t1140 486.048
R9148 VPWR.t818 VPWR.t1218 486.048
R9149 VPWR.t1167 VPWR.t894 486.048
R9150 VPWR.t554 VPWR.t1166 486.048
R9151 VPWR.t1220 VPWR.t1870 486.048
R9152 VPWR.t1343 VPWR.t920 486.048
R9153 VPWR.t919 VPWR.t1840 486.048
R9154 VPWR.t1924 VPWR.t766 486.048
R9155 VPWR.t765 VPWR.t761 486.048
R9156 VPWR.t784 VPWR.t764 486.048
R9157 VPWR.t1165 VPWR.t315 486.048
R9158 VPWR.t1193 VPWR.t1038 486.048
R9159 VPWR.t1904 VPWR.t1383 486.048
R9160 VPWR.t1476 VPWR.t1044 486.048
R9161 VPWR.t996 VPWR.t1043 486.048
R9162 VPWR.t1591 VPWR.t940 486.048
R9163 VPWR.t955 VPWR.t1381 486.048
R9164 VPWR.t492 VPWR.t1380 486.048
R9165 VPWR.t869 VPWR.t594 486.048
R9166 VPWR.t1187 VPWR.t593 486.048
R9167 VPWR.t747 VPWR.t1382 486.048
R9168 VPWR.t1617 VPWR.t1040 486.048
R9169 VPWR.t1575 VPWR.t1039 486.048
R9170 VPWR.t1294 VPWR.t1379 486.048
R9171 VPWR.t414 VPWR.t1046 486.048
R9172 VPWR.t520 VPWR.t1045 486.048
R9173 VPWR.t188 VPWR.t592 486.048
R9174 VPWR.t1024 VPWR.t1389 486.048
R9175 VPWR.t1384 VPWR.t469 486.048
R9176 VPWR.t1886 VPWR.t1442 486.048
R9177 VPWR.t1885 VPWR.t1266 486.048
R9178 VPWR.t1388 VPWR.t1543 486.048
R9179 VPWR.t990 VPWR.t1153 486.048
R9180 VPWR.t989 VPWR.t808 486.048
R9181 VPWR.t1387 VPWR.t650 486.048
R9182 VPWR.t1386 VPWR.t943 486.048
R9183 VPWR.t991 VPWR.t1240 486.048
R9184 VPWR.t1884 VPWR.t1318 486.048
R9185 VPWR.t1883 VPWR.t1254 486.048
R9186 VPWR.t988 VPWR.t1914 486.048
R9187 VPWR.t987 VPWR.t741 486.048
R9188 VPWR.t1887 VPWR.t772 486.048
R9189 VPWR.t1385 VPWR.t358 486.048
R9190 VPWR.t429 VPWR.t93 486.048
R9191 VPWR.t1563 VPWR.t224 486.048
R9192 VPWR.t1490 VPWR.t353 486.048
R9193 VPWR.t1504 VPWR.t15 486.048
R9194 VPWR.t590 VPWR.t119 486.048
R9195 VPWR.t274 VPWR.t1142 486.048
R9196 VPWR.t820 VPWR.t276 486.048
R9197 VPWR.t124 VPWR.t896 486.048
R9198 VPWR.t556 VPWR.t154 486.048
R9199 VPWR.t272 VPWR.t1872 486.048
R9200 VPWR.t23 VPWR.t1345 486.048
R9201 VPWR.t42 VPWR.t1842 486.048
R9202 VPWR.t286 VPWR.t1073 486.048
R9203 VPWR.t685 VPWR.t304 486.048
R9204 VPWR.t342 VPWR.t788 486.048
R9205 VPWR.t299 VPWR.t174 486.048
R9206 VPWR.t159 VPWR.t28 486.048
R9207 VPWR.t288 VPWR.t164 486.048
R9208 VPWR.t294 VPWR.t306 486.048
R9209 VPWR.t68 VPWR.t334 486.048
R9210 VPWR.t58 VPWR.t176 486.048
R9211 VPWR.t331 VPWR.t202 486.048
R9212 VPWR.t226 VPWR.t55 486.048
R9213 VPWR.t90 VPWR.t63 486.048
R9214 VPWR.t98 VPWR.t218 486.048
R9215 VPWR.t328 VPWR.t200 486.048
R9216 VPWR.t361 VPWR.t95 486.048
R9217 VPWR.t113 VPWR.t380 486.048
R9218 VPWR.t234 VPWR.t241 486.048
R9219 VPWR.t374 VPWR.t253 486.048
R9220 VPWR.t278 VPWR.t7 486.048
R9221 VPWR.t250 VPWR.t129 486.048
R9222 VPWR.t30 VPWR.t302 486.048
R9223 VPWR.t47 VPWR.t166 486.048
R9224 VPWR.t179 VPWR.t172 486.048
R9225 VPWR.t339 VPWR.t213 486.048
R9226 VPWR.t60 VPWR.t321 486.048
R9227 VPWR.t88 VPWR.t207 486.048
R9228 VPWR.t103 VPWR.t318 486.048
R9229 VPWR.t326 VPWR.t355 486.048
R9230 VPWR.t369 VPWR.t100 486.048
R9231 VPWR.t86 VPWR.t204 486.048
R9232 VPWR.t239 VPWR.t363 486.048
R9233 VPWR.t261 VPWR.t382 486.048
R9234 VPWR.t111 VPWR.t126 486.048
R9235 VPWR.t137 VPWR.t255 486.048
R9236 VPWR.t162 VPWR.t283 486.048
R9237 VPWR.t134 VPWR.t13 486.048
R9238 VPWR.t769 VPWR.t1130 463.954
R9239 VPWR.t1731 VPWR.t1191 463.954
R9240 VPWR.t689 VPWR.t1327 463.954
R9241 VPWR.t1326 VPWR.t1492 463.954
R9242 VPWR.t1508 VPWR.t768 463.954
R9243 VPWR.t1163 VPWR.t1595 463.954
R9244 VPWR.t959 VPWR.t1162 463.954
R9245 VPWR.t767 VPWR.t1579 463.954
R9246 VPWR.t900 VPWR.t1733 463.954
R9247 VPWR.t1164 VPWR.t1684 463.954
R9248 VPWR.t745 VPWR.t1325 463.954
R9249 VPWR.t1324 VPWR.t1605 463.954
R9250 VPWR.t1573 VPWR.t1161 463.954
R9251 VPWR.t1160 VPWR.t1077 463.954
R9252 VPWR.t412 VPWR.t1328 463.954
R9253 VPWR.t1732 VPWR.t1846 463.954
R9254 VPWR.t1867 VPWR.t1119 463.954
R9255 VPWR.t1201 VPWR.t977 463.954
R9256 VPWR.t1674 VPWR.t1377 463.954
R9257 VPWR.t1470 VPWR.t1376 463.954
R9258 VPWR.t390 VPWR.t1866 463.954
R9259 VPWR.t1335 VPWR.t1660 463.954
R9260 VPWR.t1145 VPWR.t1659 463.954
R9261 VPWR.t800 VPWR.t1865 463.954
R9262 VPWR.t831 VPWR.t979 463.954
R9263 VPWR.t839 VPWR.t1661 463.954
R9264 VPWR.t518 VPWR.t1375 463.954
R9265 VPWR.t1310 VPWR.t1868 463.954
R9266 VPWR.t1258 VPWR.t1658 463.954
R9267 VPWR.t1306 VPWR.t1657 463.954
R9268 VPWR.t1358 VPWR.t1378 463.954
R9269 VPWR.t598 VPWR.t978 463.954
R9270 VPWR.t1263 VPWR.t1105 463.954
R9271 VPWR.t852 VPWR.t1053 463.954
R9272 VPWR.t1644 VPWR.t1709 463.954
R9273 VPWR.t1446 VPWR.t1643 463.954
R9274 VPWR.t1262 VPWR.t1274 463.954
R9275 VPWR.t1695 VPWR.t1051 463.954
R9276 VPWR.t1050 VPWR.t911 463.954
R9277 VPWR.t482 VPWR.t1056 463.954
R9278 VPWR.t1055 VPWR.t886 463.954
R9279 VPWR.t884 VPWR.t1052 463.954
R9280 VPWR.t1642 VPWR.t723 463.954
R9281 VPWR.t1174 VPWR.t1641 463.954
R9282 VPWR.t1049 VPWR.t1828 463.954
R9283 VPWR.t1916 VPWR.t1646 463.954
R9284 VPWR.t1645 VPWR.t564 463.954
R9285 VPWR.t780 VPWR.t1054 463.954
R9286 VPWR.t1428 VPWR.t1113 463.954
R9287 VPWR.t1423 VPWR.t1018 463.954
R9288 VPWR.t698 VPWR.t471 463.954
R9289 VPWR.t697 VPWR.t1460 463.954
R9290 VPWR.t1427 VPWR.t396 463.954
R9291 VPWR.t1878 VPWR.t1545 463.954
R9292 VPWR.t1877 VPWR.t1155 463.954
R9293 VPWR.t1426 VPWR.t810 463.954
R9294 VPWR.t1425 VPWR.t932 463.954
R9295 VPWR.t1422 VPWR.t945 463.954
R9296 VPWR.t696 VPWR.t1234 463.954
R9297 VPWR.t695 VPWR.t1320 463.954
R9298 VPWR.t1876 VPWR.t1248 463.954
R9299 VPWR.t1875 VPWR.t1715 463.954
R9300 VPWR.t1874 VPWR.t735 463.954
R9301 VPWR.t1424 VPWR.t604 463.954
R9302 VPWR.t1061 VPWR.t1125 463.954
R9303 VPWR.t982 VPWR.t824 463.954
R9304 VPWR.t1551 VPWR.t1158 463.954
R9305 VPWR.t1157 VPWR.t1482 463.954
R9306 VPWR.t998 VPWR.t877 463.954
R9307 VPWR.t1691 VPWR.t1329 463.954
R9308 VPWR.t620 VPWR.t1690 463.954
R9309 VPWR.t876 VPWR.t1589 463.954
R9310 VPWR.t871 VPWR.t875 463.954
R9311 VPWR.t1692 VPWR.t544 463.954
R9312 VPWR.t506 VPWR.t1063 463.954
R9313 VPWR.t1062 VPWR.t1664 463.954
R9314 VPWR.t1282 VPWR.t1689 463.954
R9315 VPWR.t1688 VPWR.t1296 463.954
R9316 VPWR.t1496 VPWR.t1159 463.954
R9317 VPWR.t983 VPWR.t522 463.954
R9318 VPWR.t633 VPWR.t1132 463.954
R9319 VPWR.t1189 VPWR.t1821 463.954
R9320 VPWR.t687 VPWR.t1350 463.954
R9321 VPWR.t1494 VPWR.t1349 463.954
R9322 VPWR.t1506 VPWR.t632 463.954
R9323 VPWR.t1593 VPWR.t1067 463.954
R9324 VPWR.t957 VPWR.t1066 463.954
R9325 VPWR.t1577 VPWR.t1144 463.954
R9326 VPWR.t898 VPWR.t1823 463.954
R9327 VPWR.t1682 VPWR.t1068 463.954
R9328 VPWR.t743 VPWR.t1348 463.954
R9329 VPWR.t1619 VPWR.t634 463.954
R9330 VPWR.t1571 VPWR.t1065 463.954
R9331 VPWR.t1075 VPWR.t1064 463.954
R9332 VPWR.t410 VPWR.t1351 463.954
R9333 VPWR.t1844 VPWR.t1822 463.954
R9334 VPWR.t1629 VPWR.t1128 463.954
R9335 VPWR.t1012 VPWR.t1604 463.954
R9336 VPWR.t1633 VPWR.t1028 463.954
R9337 VPWR.t1488 VPWR.t1632 463.954
R9338 VPWR.t468 VPWR.t1510 463.954
R9339 VPWR.t1625 VPWR.t1602 463.954
R9340 VPWR.t1601 VPWR.t654 463.954
R9341 VPWR.t1585 VPWR.t467 463.954
R9342 VPWR.t466 VPWR.t664 463.954
R9343 VPWR.t1034 VPWR.t1603 463.954
R9344 VPWR.t1631 VPWR.t751 463.954
R9345 VPWR.t878 VPWR.t1630 463.954
R9346 VPWR.t1600 VPWR.t1567 463.954
R9347 VPWR.t1079 VPWR.t1599 463.954
R9348 VPWR.t1634 VPWR.t418 463.954
R9349 VPWR.t1848 VPWR.t465 463.954
R9350 VPWR.t707 VPWR.t1107 463.954
R9351 VPWR.t702 VPWR.t433 463.954
R9352 VPWR.t1004 VPWR.t1707 463.954
R9353 VPWR.t1003 VPWR.t1448 463.954
R9354 VPWR.t706 VPWR.t1270 463.954
R9355 VPWR.t1009 VPWR.t1693 463.954
R9356 VPWR.t1008 VPWR.t909 463.954
R9357 VPWR.t705 VPWR.t480 463.954
R9358 VPWR.t704 VPWR.t648 463.954
R9359 VPWR.t701 VPWR.t882 463.954
R9360 VPWR.t1002 VPWR.t721 463.954
R9361 VPWR.t1001 VPWR.t1172 463.954
R9362 VPWR.t1007 VPWR.t536 463.954
R9363 VPWR.t1006 VPWR.t1912 463.954
R9364 VPWR.t1005 VPWR.t562 463.954
R9365 VPWR.t703 VPWR.t776 463.954
R9366 VPWR.t713 VPWR.t1123 463.954
R9367 VPWR.t1824 VPWR.t826 463.954
R9368 VPWR.t1553 VPWR.t717 463.954
R9369 VPWR.t716 VPWR.t1480 463.954
R9370 VPWR.t1390 VPWR.t712 463.954
R9371 VPWR.t1530 VPWR.t1331 463.954
R9372 VPWR.t622 VPWR.t1529 463.954
R9373 VPWR.t1827 VPWR.t790 463.954
R9374 VPWR.t873 VPWR.t1826 463.954
R9375 VPWR.t1531 VPWR.t546 463.954
R9376 VPWR.t508 VPWR.t715 463.954
R9377 VPWR.t714 VPWR.t1666 463.954
R9378 VPWR.t1284 VPWR.t1528 463.954
R9379 VPWR.t1527 VPWR.t1298 463.954
R9380 VPWR.t1498 VPWR.t718 463.954
R9381 VPWR.t1825 VPWR.t524 463.954
R9382 VPWR.t968 VPWR.t1109 463.954
R9383 VPWR.t431 VPWR.t963 463.954
R9384 VPWR.t1705 VPWR.t845 463.954
R9385 VPWR.t1450 VPWR.t1861 463.954
R9386 VPWR.t1268 VPWR.t967 463.954
R9387 VPWR.t1672 VPWR.t850 463.954
R9388 VPWR.t907 VPWR.t849 463.954
R9389 VPWR.t478 VPWR.t966 463.954
R9390 VPWR.t644 VPWR.t965 463.954
R9391 VPWR.t880 VPWR.t851 463.954
R9392 VPWR.t719 VPWR.t1860 463.954
R9393 VPWR.t1170 VPWR.t1859 463.954
R9394 VPWR.t534 VPWR.t848 463.954
R9395 VPWR.t1908 VPWR.t847 463.954
R9396 VPWR.t560 VPWR.t846 463.954
R9397 VPWR.t774 VPWR.t964 463.954
R9398 VPWR.t1433 VPWR.t1121 463.954
R9399 VPWR.t1347 VPWR.t828 463.954
R9400 VPWR.t1650 VPWR.t1555 463.954
R9401 VPWR.t1649 VPWR.t1478 463.954
R9402 VPWR.t1432 VPWR.t1394 463.954
R9403 VPWR.t1655 VPWR.t1333 463.954
R9404 VPWR.t1654 VPWR.t624 463.954
R9405 VPWR.t1431 VPWR.t792 463.954
R9406 VPWR.t1430 VPWR.t658 463.954
R9407 VPWR.t1656 VPWR.t548 463.954
R9408 VPWR.t1648 VPWR.t510 463.954
R9409 VPWR.t1647 VPWR.t1668 463.954
R9410 VPWR.t1653 VPWR.t1286 463.954
R9411 VPWR.t1652 VPWR.t1300 463.954
R9412 VPWR.t1651 VPWR.t1500 463.954
R9413 VPWR.t1429 VPWR.t528 463.954
R9414 VPWR.t539 VPWR.t1115 463.954
R9415 VPWR.t1016 VPWR.t1855 463.954
R9416 VPWR.t543 VPWR.t1680 463.954
R9417 VPWR.t1462 VPWR.t542 463.954
R9418 VPWR.t538 VPWR.t394 463.954
R9419 VPWR.t1541 VPWR.t906 463.954
R9420 VPWR.t905 VPWR.t1151 463.954
R9421 VPWR.t806 VPWR.t1858 463.954
R9422 VPWR.t1857 VPWR.t930 463.954
R9423 VPWR.t941 VPWR.t1854 463.954
R9424 VPWR.t541 VPWR.t1232 463.954
R9425 VPWR.t1316 VPWR.t540 463.954
R9426 VPWR.t904 VPWR.t1246 463.954
R9427 VPWR.t1713 VPWR.t903 463.954
R9428 VPWR.t902 VPWR.t733 463.954
R9429 VPWR.t602 VPWR.t1856 463.954
R9430 VPWR.t1169 VPWR.t1111 463.954
R9431 VPWR.t1020 VPWR.t1221 463.954
R9432 VPWR.t763 VPWR.t473 463.954
R9433 VPWR.t1458 VPWR.t921 463.954
R9434 VPWR.t1168 VPWR.t1514 463.954
R9435 VPWR.t1547 VPWR.t1219 463.954
R9436 VPWR.t1218 VPWR.t1134 463.954
R9437 VPWR.t812 VPWR.t1167 463.954
R9438 VPWR.t1166 VPWR.t934 463.954
R9439 VPWR.t947 VPWR.t1220 463.954
R9440 VPWR.t920 VPWR.t1236 463.954
R9441 VPWR.t1322 VPWR.t919 463.954
R9442 VPWR.t766 VPWR.t1250 463.954
R9443 VPWR.t1717 VPWR.t765 463.954
R9444 VPWR.t764 VPWR.t737 463.954
R9445 VPWR.t608 VPWR.t1165 463.954
R9446 VPWR.t1038 VPWR.t1103 463.954
R9447 VPWR.t1383 VPWR.t854 463.954
R9448 VPWR.t1044 VPWR.t1900 463.954
R9449 VPWR.t1043 VPWR.t1440 463.954
R9450 VPWR.t940 VPWR.t1280 463.954
R9451 VPWR.t1381 VPWR.t1701 463.954
R9452 VPWR.t1380 VPWR.t917 463.954
R9453 VPWR.t594 VPWR.t488 463.954
R9454 VPWR.t593 VPWR.t890 463.954
R9455 VPWR.t1382 VPWR.t1183 463.954
R9456 VPWR.t1040 VPWR.t725 463.954
R9457 VPWR.t1039 VPWR.t1613 463.954
R9458 VPWR.t1379 VPWR.t1830 463.954
R9459 VPWR.t1046 VPWR.t1920 463.954
R9460 VPWR.t1045 VPWR.t402 463.954
R9461 VPWR.t592 VPWR.t786 463.954
R9462 VPWR.t1389 VPWR.t1117 463.954
R9463 VPWR.t1203 VPWR.t1384 463.954
R9464 VPWR.t1676 VPWR.t1886 463.954
R9465 VPWR.t1466 VPWR.t1885 463.954
R9466 VPWR.t392 VPWR.t1388 463.954
R9467 VPWR.t1337 VPWR.t990 463.954
R9468 VPWR.t1147 VPWR.t989 463.954
R9469 VPWR.t802 VPWR.t1387 463.954
R9470 VPWR.t835 VPWR.t1386 463.954
R9471 VPWR.t841 VPWR.t991 463.954
R9472 VPWR.t1230 VPWR.t1884 463.954
R9473 VPWR.t1312 VPWR.t1883 463.954
R9474 VPWR.t1260 VPWR.t988 463.954
R9475 VPWR.t1711 VPWR.t987 463.954
R9476 VPWR.t1360 VPWR.t1887 463.954
R9477 VPWR.t600 VPWR.t1385 463.954
R9478 VPWR.t93 VPWR.t108 463.954
R9479 VPWR.t224 VPWR.t269 463.954
R9480 VPWR.t353 VPWR.t371 463.954
R9481 VPWR.t15 VPWR.t142 463.954
R9482 VPWR.t119 VPWR.t244 463.954
R9483 VPWR.t266 VPWR.t274 463.954
R9484 VPWR.t276 VPWR.t17 463.954
R9485 VPWR.t139 VPWR.t124 463.954
R9486 VPWR.t154 VPWR.t280 463.954
R9487 VPWR.t296 VPWR.t272 463.954
R9488 VPWR.t39 VPWR.t23 463.954
R9489 VPWR.t169 VPWR.t42 463.954
R9490 VPWR.t210 VPWR.t286 463.954
R9491 VPWR.t304 VPWR.t33 463.954
R9492 VPWR.t83 VPWR.t342 463.954
R9493 VPWR.t174 VPWR.t191 463.954
R9494 VPWR.t28 VPWR.t52 463.954
R9495 VPWR.t164 VPWR.t197 463.954
R9496 VPWR.t309 VPWR.t294 463.954
R9497 VPWR.t334 VPWR.t74 463.954
R9498 VPWR.t185 VPWR.t58 463.954
R9499 VPWR.t202 VPWR.t194 463.954
R9500 VPWR.t350 VPWR.t226 463.954
R9501 VPWR.t63 VPWR.t71 463.954
R9502 VPWR.t231 VPWR.t98 463.954
R9503 VPWR.t200 VPWR.t247 463.954
R9504 VPWR.t377 VPWR.t361 463.954
R9505 VPWR.t380 VPWR.t121 463.954
R9506 VPWR.t151 VPWR.t234 463.954
R9507 VPWR.t253 VPWR.t1 463.954
R9508 VPWR.t20 VPWR.t278 463.954
R9509 VPWR.t129 VPWR.t145 463.954
R9510 VPWR.t302 VPWR.t312 463.954
R9511 VPWR.t80 VPWR.t47 463.954
R9512 VPWR.t172 VPWR.t182 463.954
R9513 VPWR.t213 VPWR.t347 463.954
R9514 VPWR.t321 VPWR.t65 463.954
R9515 VPWR.t77 VPWR.t88 463.954
R9516 VPWR.t236 VPWR.t103 463.954
R9517 VPWR.t344 VPWR.t326 463.954
R9518 VPWR.t105 VPWR.t369 463.954
R9519 VPWR.t131 VPWR.t86 463.954
R9520 VPWR.t258 VPWR.t239 463.954
R9521 VPWR.t4 VPWR.t261 463.954
R9522 VPWR.t25 VPWR.t111 463.954
R9523 VPWR.t263 VPWR.t137 463.954
R9524 VPWR.t291 VPWR.t162 463.954
R9525 VPWR.t13 VPWR.t10 463.954
R9526 VPWR.n2626 VPWR.t1089 428.822
R9527 VPWR.n1595 VPWR.n1594 376.045
R9528 VPWR.n2506 VPWR.n2505 376.045
R9529 VPWR.n1468 VPWR.n1467 376.045
R9530 VPWR.n351 VPWR.n350 376.045
R9531 VPWR.n2568 VPWR.n2567 376.045
R9532 VPWR.n1535 VPWR.n1534 376.045
R9533 VPWR.n349 VPWR.n348 376.045
R9534 VPWR.n2508 VPWR.n2507 376.045
R9535 VPWR.n966 VPWR.n965 376.045
R9536 VPWR.n2478 VPWR.n2477 376.045
R9537 VPWR.n2476 VPWR.n2475 376.045
R9538 VPWR.n321 VPWR.n320 376.045
R9539 VPWR.n2554 VPWR.n2553 376.045
R9540 VPWR.n974 VPWR.n973 376.045
R9541 VPWR.n2446 VPWR.n2445 376.045
R9542 VPWR.n325 VPWR.n324 376.045
R9543 VPWR.n2544 VPWR.n2543 376.045
R9544 VPWR.n1890 VPWR.n1889 376.045
R9545 VPWR.n1888 VPWR.n1887 376.045
R9546 VPWR.n1880 VPWR.n1879 376.045
R9547 VPWR.n390 VPWR.n389 376.045
R9548 VPWR.n394 VPWR.n393 376.045
R9549 VPWR.n398 VPWR.n397 376.045
R9550 VPWR.n2456 VPWR.n2455 376.045
R9551 VPWR.n333 VPWR.n332 376.045
R9552 VPWR.n2532 VPWR.n2531 376.045
R9553 VPWR.n1878 VPWR.n1877 376.045
R9554 VPWR.n406 VPWR.n405 376.045
R9555 VPWR.n2458 VPWR.n2457 376.045
R9556 VPWR.n337 VPWR.n336 376.045
R9557 VPWR.n2530 VPWR.n2529 376.045
R9558 VPWR.n2309 VPWR.n2308 376.045
R9559 VPWR.n2311 VPWR.n2310 376.045
R9560 VPWR.n2319 VPWR.n2318 376.045
R9561 VPWR.n2321 VPWR.n2320 376.045
R9562 VPWR.n2331 VPWR.n2330 376.045
R9563 VPWR.n2339 VPWR.n2338 376.045
R9564 VPWR.n2341 VPWR.n2340 376.045
R9565 VPWR.n2349 VPWR.n2348 376.045
R9566 VPWR.n2351 VPWR.n2350 376.045
R9567 VPWR.n2359 VPWR.n2358 376.045
R9568 VPWR.n2361 VPWR.n2360 376.045
R9569 VPWR.n2369 VPWR.n2368 376.045
R9570 VPWR.n2371 VPWR.n2370 376.045
R9571 VPWR.n2379 VPWR.n2378 376.045
R9572 VPWR.n2329 VPWR.n2328 376.045
R9573 VPWR.n543 VPWR.n542 376.045
R9574 VPWR.n541 VPWR.n540 376.045
R9575 VPWR.n537 VPWR.n536 376.045
R9576 VPWR.n533 VPWR.n532 376.045
R9577 VPWR.n525 VPWR.n524 376.045
R9578 VPWR.n521 VPWR.n520 376.045
R9579 VPWR.n517 VPWR.n516 376.045
R9580 VPWR.n513 VPWR.n512 376.045
R9581 VPWR.n509 VPWR.n508 376.045
R9582 VPWR.n505 VPWR.n504 376.045
R9583 VPWR.n501 VPWR.n500 376.045
R9584 VPWR.n497 VPWR.n496 376.045
R9585 VPWR.n493 VPWR.n492 376.045
R9586 VPWR.n489 VPWR.n488 376.045
R9587 VPWR.n529 VPWR.n528 376.045
R9588 VPWR.n2282 VPWR.n2281 376.045
R9589 VPWR.n2280 VPWR.n2279 376.045
R9590 VPWR.n2272 VPWR.n2271 376.045
R9591 VPWR.n2270 VPWR.n2269 376.045
R9592 VPWR.n2260 VPWR.n2259 376.045
R9593 VPWR.n2252 VPWR.n2251 376.045
R9594 VPWR.n2250 VPWR.n2249 376.045
R9595 VPWR.n2242 VPWR.n2241 376.045
R9596 VPWR.n2240 VPWR.n2239 376.045
R9597 VPWR.n2232 VPWR.n2231 376.045
R9598 VPWR.n2230 VPWR.n2229 376.045
R9599 VPWR.n2222 VPWR.n2221 376.045
R9600 VPWR.n2220 VPWR.n2219 376.045
R9601 VPWR.n2212 VPWR.n2211 376.045
R9602 VPWR.n2262 VPWR.n2261 376.045
R9603 VPWR.n582 VPWR.n581 376.045
R9604 VPWR.n586 VPWR.n585 376.045
R9605 VPWR.n590 VPWR.n589 376.045
R9606 VPWR.n594 VPWR.n593 376.045
R9607 VPWR.n602 VPWR.n601 376.045
R9608 VPWR.n606 VPWR.n605 376.045
R9609 VPWR.n610 VPWR.n609 376.045
R9610 VPWR.n614 VPWR.n613 376.045
R9611 VPWR.n618 VPWR.n617 376.045
R9612 VPWR.n622 VPWR.n621 376.045
R9613 VPWR.n626 VPWR.n625 376.045
R9614 VPWR.n630 VPWR.n629 376.045
R9615 VPWR.n634 VPWR.n633 376.045
R9616 VPWR.n638 VPWR.n637 376.045
R9617 VPWR.n598 VPWR.n597 376.045
R9618 VPWR.n2113 VPWR.n2112 376.045
R9619 VPWR.n2115 VPWR.n2114 376.045
R9620 VPWR.n2123 VPWR.n2122 376.045
R9621 VPWR.n2125 VPWR.n2124 376.045
R9622 VPWR.n2135 VPWR.n2134 376.045
R9623 VPWR.n2143 VPWR.n2142 376.045
R9624 VPWR.n2145 VPWR.n2144 376.045
R9625 VPWR.n2153 VPWR.n2152 376.045
R9626 VPWR.n2155 VPWR.n2154 376.045
R9627 VPWR.n2163 VPWR.n2162 376.045
R9628 VPWR.n2165 VPWR.n2164 376.045
R9629 VPWR.n2173 VPWR.n2172 376.045
R9630 VPWR.n2175 VPWR.n2174 376.045
R9631 VPWR.n2183 VPWR.n2182 376.045
R9632 VPWR.n2133 VPWR.n2132 376.045
R9633 VPWR.n735 VPWR.n734 376.045
R9634 VPWR.n733 VPWR.n732 376.045
R9635 VPWR.n729 VPWR.n728 376.045
R9636 VPWR.n725 VPWR.n724 376.045
R9637 VPWR.n717 VPWR.n716 376.045
R9638 VPWR.n713 VPWR.n712 376.045
R9639 VPWR.n709 VPWR.n708 376.045
R9640 VPWR.n705 VPWR.n704 376.045
R9641 VPWR.n701 VPWR.n700 376.045
R9642 VPWR.n697 VPWR.n696 376.045
R9643 VPWR.n693 VPWR.n692 376.045
R9644 VPWR.n689 VPWR.n688 376.045
R9645 VPWR.n685 VPWR.n684 376.045
R9646 VPWR.n681 VPWR.n680 376.045
R9647 VPWR.n721 VPWR.n720 376.045
R9648 VPWR.n2086 VPWR.n2085 376.045
R9649 VPWR.n2084 VPWR.n2083 376.045
R9650 VPWR.n2076 VPWR.n2075 376.045
R9651 VPWR.n2074 VPWR.n2073 376.045
R9652 VPWR.n2064 VPWR.n2063 376.045
R9653 VPWR.n2056 VPWR.n2055 376.045
R9654 VPWR.n2054 VPWR.n2053 376.045
R9655 VPWR.n2046 VPWR.n2045 376.045
R9656 VPWR.n2044 VPWR.n2043 376.045
R9657 VPWR.n2036 VPWR.n2035 376.045
R9658 VPWR.n2034 VPWR.n2033 376.045
R9659 VPWR.n2026 VPWR.n2025 376.045
R9660 VPWR.n2024 VPWR.n2023 376.045
R9661 VPWR.n2016 VPWR.n2015 376.045
R9662 VPWR.n2066 VPWR.n2065 376.045
R9663 VPWR.n774 VPWR.n773 376.045
R9664 VPWR.n778 VPWR.n777 376.045
R9665 VPWR.n782 VPWR.n781 376.045
R9666 VPWR.n786 VPWR.n785 376.045
R9667 VPWR.n794 VPWR.n793 376.045
R9668 VPWR.n798 VPWR.n797 376.045
R9669 VPWR.n802 VPWR.n801 376.045
R9670 VPWR.n806 VPWR.n805 376.045
R9671 VPWR.n810 VPWR.n809 376.045
R9672 VPWR.n814 VPWR.n813 376.045
R9673 VPWR.n818 VPWR.n817 376.045
R9674 VPWR.n822 VPWR.n821 376.045
R9675 VPWR.n826 VPWR.n825 376.045
R9676 VPWR.n830 VPWR.n829 376.045
R9677 VPWR.n790 VPWR.n789 376.045
R9678 VPWR.n1917 VPWR.n1916 376.045
R9679 VPWR.n1919 VPWR.n1918 376.045
R9680 VPWR.n1927 VPWR.n1926 376.045
R9681 VPWR.n1929 VPWR.n1928 376.045
R9682 VPWR.n1939 VPWR.n1938 376.045
R9683 VPWR.n1947 VPWR.n1946 376.045
R9684 VPWR.n1949 VPWR.n1948 376.045
R9685 VPWR.n1957 VPWR.n1956 376.045
R9686 VPWR.n1959 VPWR.n1958 376.045
R9687 VPWR.n1967 VPWR.n1966 376.045
R9688 VPWR.n1969 VPWR.n1968 376.045
R9689 VPWR.n1977 VPWR.n1976 376.045
R9690 VPWR.n1979 VPWR.n1978 376.045
R9691 VPWR.n1987 VPWR.n1986 376.045
R9692 VPWR.n1937 VPWR.n1936 376.045
R9693 VPWR.n927 VPWR.n926 376.045
R9694 VPWR.n925 VPWR.n924 376.045
R9695 VPWR.n921 VPWR.n920 376.045
R9696 VPWR.n917 VPWR.n916 376.045
R9697 VPWR.n909 VPWR.n908 376.045
R9698 VPWR.n905 VPWR.n904 376.045
R9699 VPWR.n901 VPWR.n900 376.045
R9700 VPWR.n897 VPWR.n896 376.045
R9701 VPWR.n893 VPWR.n892 376.045
R9702 VPWR.n889 VPWR.n888 376.045
R9703 VPWR.n885 VPWR.n884 376.045
R9704 VPWR.n881 VPWR.n880 376.045
R9705 VPWR.n877 VPWR.n876 376.045
R9706 VPWR.n873 VPWR.n872 376.045
R9707 VPWR.n913 VPWR.n912 376.045
R9708 VPWR.n1870 VPWR.n1869 376.045
R9709 VPWR.n982 VPWR.n981 376.045
R9710 VPWR.n1494 VPWR.n1493 376.045
R9711 VPWR.n1221 VPWR.n1220 376.045
R9712 VPWR.n402 VPWR.n401 376.045
R9713 VPWR.n2466 VPWR.n2465 376.045
R9714 VPWR.n341 VPWR.n340 376.045
R9715 VPWR.n2520 VPWR.n2519 376.045
R9716 VPWR.n978 VPWR.n977 376.045
R9717 VPWR.n1492 VPWR.n1491 376.045
R9718 VPWR.n1185 VPWR.n1184 376.045
R9719 VPWR.n1868 VPWR.n1867 376.045
R9720 VPWR.n986 VPWR.n985 376.045
R9721 VPWR.n1506 VPWR.n1505 376.045
R9722 VPWR.n1219 VPWR.n1218 376.045
R9723 VPWR.n410 VPWR.n409 376.045
R9724 VPWR.n418 VPWR.n417 376.045
R9725 VPWR.n422 VPWR.n421 376.045
R9726 VPWR.n426 VPWR.n425 376.045
R9727 VPWR.n430 VPWR.n429 376.045
R9728 VPWR.n434 VPWR.n433 376.045
R9729 VPWR.n438 VPWR.n437 376.045
R9730 VPWR.n442 VPWR.n441 376.045
R9731 VPWR.n446 VPWR.n445 376.045
R9732 VPWR.n414 VPWR.n413 376.045
R9733 VPWR.n2448 VPWR.n2447 376.045
R9734 VPWR.n329 VPWR.n328 376.045
R9735 VPWR.n2542 VPWR.n2541 376.045
R9736 VPWR.n990 VPWR.n989 376.045
R9737 VPWR.n1508 VPWR.n1507 376.045
R9738 VPWR.n1216 VPWR.n1215 376.045
R9739 VPWR.n1860 VPWR.n1859 376.045
R9740 VPWR.n1850 VPWR.n1849 376.045
R9741 VPWR.n1848 VPWR.n1847 376.045
R9742 VPWR.n1840 VPWR.n1839 376.045
R9743 VPWR.n1838 VPWR.n1837 376.045
R9744 VPWR.n1830 VPWR.n1829 376.045
R9745 VPWR.n1828 VPWR.n1827 376.045
R9746 VPWR.n1820 VPWR.n1819 376.045
R9747 VPWR.n1858 VPWR.n1857 376.045
R9748 VPWR.n994 VPWR.n993 376.045
R9749 VPWR.n1520 VPWR.n1519 376.045
R9750 VPWR.n1213 VPWR.n1212 376.045
R9751 VPWR.n2468 VPWR.n2467 376.045
R9752 VPWR.n345 VPWR.n344 376.045
R9753 VPWR.n2518 VPWR.n2517 376.045
R9754 VPWR.n1481 VPWR.n1480 376.045
R9755 VPWR.n1182 VPWR.n1181 376.045
R9756 VPWR.n998 VPWR.n997 376.045
R9757 VPWR.n1522 VPWR.n1521 376.045
R9758 VPWR.n1205 VPWR.n1204 376.045
R9759 VPWR.n2438 VPWR.n2437 376.045
R9760 VPWR.n2428 VPWR.n2427 376.045
R9761 VPWR.n2426 VPWR.n2425 376.045
R9762 VPWR.n2418 VPWR.n2417 376.045
R9763 VPWR.n2416 VPWR.n2415 376.045
R9764 VPWR.n2408 VPWR.n2407 376.045
R9765 VPWR.n2436 VPWR.n2435 376.045
R9766 VPWR.n317 VPWR.n316 376.045
R9767 VPWR.n2556 VPWR.n2555 376.045
R9768 VPWR.n1537 VPWR.n1536 376.045
R9769 VPWR.n1202 VPWR.n1201 376.045
R9770 VPWR.n1002 VPWR.n1001 376.045
R9771 VPWR.n1006 VPWR.n1005 376.045
R9772 VPWR.n1010 VPWR.n1009 376.045
R9773 VPWR.n1014 VPWR.n1013 376.045
R9774 VPWR.n1018 VPWR.n1017 376.045
R9775 VPWR.n1022 VPWR.n1021 376.045
R9776 VPWR.n970 VPWR.n969 376.045
R9777 VPWR.n1475 VPWR.n1474 376.045
R9778 VPWR.n1593 VPWR.n1592 376.045
R9779 VPWR.n313 VPWR.n312 376.045
R9780 VPWR.n2566 VPWR.n2565 376.045
R9781 VPWR.n1199 VPWR.n1198 376.045
R9782 VPWR.n1762 VPWR.n1761 376.045
R9783 VPWR.n1191 VPWR.n1190 376.045
R9784 VPWR.n309 VPWR.n308 376.045
R9785 VPWR.n305 VPWR.n304 376.045
R9786 VPWR.n297 VPWR.n296 376.045
R9787 VPWR.n301 VPWR.n300 376.045
R9788 VPWR.n1741 VPWR.n1740 376.045
R9789 VPWR.n1750 VPWR.n1749 376.045
R9790 VPWR.n1791 VPWR.n1790 376.045
R9791 VPWR.n1760 VPWR.n1759 376.045
R9792 VPWR.n1188 VPWR.n1187 376.045
R9793 VPWR.n2578 VPWR.n2577 376.045
R9794 VPWR.n2580 VPWR.n2579 376.045
R9795 VPWR.n2590 VPWR.n2589 376.045
R9796 VPWR.n1739 VPWR.n1738 376.045
R9797 VPWR.n1339 VPWR.t1743 342.841
R9798 VPWR.n1378 VPWR.t497 342.841
R9799 VPWR.n1415 VPWR.t1211 342.841
R9800 VPWR.n2693 VPWR.t477 342.841
R9801 VPWR.n2656 VPWR.t676 342.841
R9802 VPWR.n2599 VPWR.t1364 342.841
R9803 VPWR.n1339 VPWR.t1740 342.839
R9804 VPWR.n1378 VPWR.t1288 342.839
R9805 VPWR.n1415 VPWR.t1407 342.839
R9806 VPWR.n2693 VPWR.t456 342.839
R9807 VPWR.n2656 VPWR.t1863 342.839
R9808 VPWR.n2599 VPWR.t1090 342.839
R9809 VPWR.n2842 VPWR.n2824 339.212
R9810 VPWR.n1306 VPWR.t619 338.488
R9811 VPWR.n2729 VPWR.t1893 338.488
R9812 VPWR.n1315 VPWR.n1314 327.377
R9813 VPWR.n1308 VPWR.n1307 327.377
R9814 VPWR.n1322 VPWR.n1321 327.377
R9815 VPWR.n1352 VPWR.n1350 327.377
R9816 VPWR.n1345 VPWR.n1343 327.377
R9817 VPWR.n1360 VPWR.n1358 327.377
R9818 VPWR.n1391 VPWR.n1389 327.377
R9819 VPWR.n1384 VPWR.n1382 327.377
R9820 VPWR.n1399 VPWR.n1397 327.377
R9821 VPWR.n1428 VPWR.n1426 327.377
R9822 VPWR.n1421 VPWR.n1419 327.377
R9823 VPWR.n1436 VPWR.n1434 327.377
R9824 VPWR.n1324 VPWR.n1323 327.375
R9825 VPWR.n1352 VPWR.n1351 327.375
R9826 VPWR.n1345 VPWR.n1344 327.375
R9827 VPWR.n1360 VPWR.n1359 327.375
R9828 VPWR.n1391 VPWR.n1390 327.375
R9829 VPWR.n1384 VPWR.n1383 327.375
R9830 VPWR.n1399 VPWR.n1398 327.375
R9831 VPWR.n1428 VPWR.n1427 327.375
R9832 VPWR.n1421 VPWR.n1420 327.375
R9833 VPWR.n1436 VPWR.n1435 327.375
R9834 VPWR.n1 VPWR 325.546
R9835 VPWR.n2667 VPWR.t455 322.262
R9836 VPWR.n2630 VPWR.t675 322.262
R9837 VPWR.n2805 VPWR.n2804 321.642
R9838 VPWR.n2722 VPWR.n2712 320.976
R9839 VPWR.n2716 VPWR.n2715 320.976
R9840 VPWR.n2710 VPWR.n2709 320.976
R9841 VPWR.n2680 VPWR.n2679 320.976
R9842 VPWR.n2686 VPWR.n2675 320.976
R9843 VPWR.n2672 VPWR.n2671 320.976
R9844 VPWR.n2643 VPWR.n2642 320.976
R9845 VPWR.n2649 VPWR.n2638 320.976
R9846 VPWR.n2635 VPWR.n2634 320.976
R9847 VPWR.n2610 VPWR.n2606 320.976
R9848 VPWR.n2614 VPWR.n2613 320.976
R9849 VPWR.n2620 VPWR.n2602 320.976
R9850 VPWR.n2727 VPWR.n2708 320.976
R9851 VPWR.n2680 VPWR.n2678 320.976
R9852 VPWR.n2686 VPWR.n2674 320.976
R9853 VPWR.n2672 VPWR.n2670 320.976
R9854 VPWR.n2643 VPWR.n2641 320.976
R9855 VPWR.n2649 VPWR.n2637 320.976
R9856 VPWR.n2635 VPWR.n2633 320.976
R9857 VPWR.n2610 VPWR.n2605 320.976
R9858 VPWR.n2614 VPWR.n2612 320.976
R9859 VPWR.n2620 VPWR.n2601 320.976
R9860 VPWR.n2801 VPWR 319.627
R9861 VPWR.n6 VPWR.n5 316.245
R9862 VPWR.n1241 VPWR.n1239 316.245
R9863 VPWR.n1264 VPWR.n1262 316.245
R9864 VPWR.n1288 VPWR.n1286 316.245
R9865 VPWR.n2784 VPWR.n2783 316.245
R9866 VPWR.n2764 VPWR.n2763 316.245
R9867 VPWR.n2745 VPWR.n2744 316.245
R9868 VPWR.n1241 VPWR.n1240 316.245
R9869 VPWR.n1264 VPWR.n1263 316.245
R9870 VPWR.n1288 VPWR.n1287 316.245
R9871 VPWR.n2784 VPWR.n2782 316.245
R9872 VPWR.n2764 VPWR.n2762 316.245
R9873 VPWR.n2745 VPWR.n2743 316.245
R9874 VPWR.n2630 VPWR.t975 313.87
R9875 VPWR.n10 VPWR.n4 310.502
R9876 VPWR.n1246 VPWR.n1238 310.502
R9877 VPWR.n1269 VPWR.n1261 310.502
R9878 VPWR.n1293 VPWR.n1285 310.502
R9879 VPWR.n2803 VPWR.n2802 310.502
R9880 VPWR.n2788 VPWR.n2787 310.502
R9881 VPWR.n2768 VPWR.n2767 310.502
R9882 VPWR.n2749 VPWR.n2748 310.502
R9883 VPWR.n1246 VPWR.n1245 310.5
R9884 VPWR.n1269 VPWR.n1268 310.5
R9885 VPWR.n1293 VPWR.n1292 310.5
R9886 VPWR.n2788 VPWR.n2786 310.5
R9887 VPWR.n2768 VPWR.n2766 310.5
R9888 VPWR.n2749 VPWR.n2747 310.5
R9889 VPWR.n2834 VPWR.n2833 279.341
R9890 VPWR.n2839 VPWR.n2838 279.341
R9891 VPWR.n1412 VPWR.t1071 255.905
R9892 VPWR.n2663 VPWR.t1869 255.905
R9893 VPWR.n1275 VPWR.t1217 255.904
R9894 VPWR.n1412 VPWR.t1072 255.904
R9895 VPWR.n2774 VPWR.t1749 255.904
R9896 VPWR.n2663 VPWR.t976 255.904
R9897 VPWR.n1303 VPWR.t1730 254.019
R9898 VPWR.n2735 VPWR.t1293 254.019
R9899 VPWR.n1335 VPWR.t1728 252.948
R9900 VPWR.n2737 VPWR.t1291 252.948
R9901 VPWR.n1373 VPWR.t984 250.722
R9902 VPWR.n2700 VPWR.t597 250.722
R9903 VPWR.n1310 VPWR.t1224 249.901
R9904 VPWR.n1346 VPWR.t1524 249.901
R9905 VPWR.n1385 VPWR.t708 249.901
R9906 VPWR.n1422 VPWR.t1526 249.901
R9907 VPWR.n2714 VPWR.t1804 249.901
R9908 VPWR.n2677 VPWR.t1801 249.901
R9909 VPWR.n2640 VPWR.t1815 249.901
R9910 VPWR.n2607 VPWR.t1769 249.901
R9911 VPWR.n1346 VPWR.t641 249.901
R9912 VPWR.n1385 VPWR.t1521 249.901
R9913 VPWR.n1422 VPWR.t866 249.901
R9914 VPWR.n2677 VPWR.t1814 249.901
R9915 VPWR.n2640 VPWR.t1767 249.901
R9916 VPWR.n2607 VPWR.t1790 249.901
R9917 VPWR.n1253 VPWR.t583 249.363
R9918 VPWR.n1338 VPWR.t1374 249.363
R9919 VPWR.n2811 VPWR.t385 249.363
R9920 VPWR.n2795 VPWR.t1534 249.363
R9921 VPWR.n2698 VPWR.t929 249.363
R9922 VPWR.n17 VPWR.t1415 249.362
R9923 VPWR.n1253 VPWR.t567 249.362
R9924 VPWR.n2795 VPWR.t448 249.362
R9925 VPWR.t1213 VPWR.t1414 248.599
R9926 VPWR.t616 VPWR.t435 248.599
R9927 VPWR.t435 VPWR.t439 248.599
R9928 VPWR.t439 VPWR.t443 248.599
R9929 VPWR.t443 VPWR.t420 248.599
R9930 VPWR.t420 VPWR.t424 248.599
R9931 VPWR.t424 VPWR.t1523 248.599
R9932 VPWR.t1523 VPWR.t1417 248.599
R9933 VPWR.t635 VPWR.t638 248.599
R9934 VPWR.t638 VPWR.t1223 248.599
R9935 VPWR.t1817 VPWR.t1793 248.599
R9936 VPWR.t1781 VPWR.t1817 248.599
R9937 VPWR.t1755 VPWR.t1781 248.599
R9938 VPWR.t1890 VPWR.t1755 248.599
R9939 VPWR.t683 VPWR.t1890 248.599
R9940 VPWR.t693 VPWR.t683 248.599
R9941 VPWR.t558 VPWR.t693 248.599
R9942 VPWR.t1750 VPWR.t384 248.599
R9943 VPWR.t1761 VPWR.t1803 248.599
R9944 VPWR.t1809 VPWR.t1761 248.599
R9945 VPWR.n15 VPWR.t1214 247.394
R9946 VPWR.n1251 VPWR.t1216 247.394
R9947 VPWR.n2809 VPWR.t1751 247.394
R9948 VPWR.n2793 VPWR.t1745 247.394
R9949 VPWR.n1251 VPWR.t1215 247.394
R9950 VPWR.n2793 VPWR.t1747 247.394
R9951 VPWR.n1304 VPWR.t1227 244.737
R9952 VPWR.n2730 VPWR.t1819 244.737
R9953 VPWR.n1374 VPWR.t569 243.886
R9954 VPWR.n2701 VPWR.t1402 243.886
R9955 VPWR.n1277 VPWR.t1413 243.512
R9956 VPWR.n1300 VPWR.t585 243.512
R9957 VPWR.n1303 VPWR.t1070 243.512
R9958 VPWR.n2776 VPWR.t387 243.512
R9959 VPWR.n2756 VPWR.t1535 243.512
R9960 VPWR.n2735 VPWR.t1671 243.512
R9961 VPWR.n1300 VPWR.t568 243.512
R9962 VPWR.n2756 VPWR.t446 243.512
R9963 VPWR.n1329 VPWR.t1729 238.339
R9964 VPWR.n2705 VPWR.t1292 238.339
R9965 VPWR.n2855 VPWR.t1041 237.99
R9966 VPWR.n2667 VPWR.t928 234.982
R9967 VPWR.t1420 VPWR.t635 228.101
R9968 VPWR.t1787 VPWR.t1809 228.101
R9969 VPWR.n2801 VPWR 224.923
R9970 VPWR.n1 VPWR 219.004
R9971 VPWR.n1444 VPWR.n1443 214.613
R9972 VPWR.n1444 VPWR.n1442 214.613
R9973 VPWR.n1236 VPWR.n1235 214.326
R9974 VPWR.n1259 VPWR.n1258 214.326
R9975 VPWR.n1283 VPWR.n1282 214.326
R9976 VPWR.n1368 VPWR.n1367 214.326
R9977 VPWR.n1407 VPWR.n1406 214.326
R9978 VPWR.n1236 VPWR.n1234 214.326
R9979 VPWR.n1259 VPWR.n1257 214.326
R9980 VPWR.n1283 VPWR.n1281 214.326
R9981 VPWR.n1368 VPWR.n1366 214.326
R9982 VPWR.n1407 VPWR.n1405 214.326
R9983 VPWR.n2 VPWR.n1 213.119
R9984 VPWR.n2808 VPWR.n2801 213.119
R9985 VPWR VPWR.t1213 207.166
R9986 VPWR.n2840 VPWR.n2839 204.424
R9987 VPWR.n2830 VPWR.n2817 204.424
R9988 VPWR.n2833 VPWR.n2820 204.424
R9989 VPWR.n2844 VPWR.n2841 204.048
R9990 VPWR VPWR.t558 201.246
R9991 VPWR.t1223 VPWR 189.409
R9992 VPWR.n2741 VPWR 184.63
R9993 VPWR.n1329 VPWR 182.952
R9994 VPWR.n2760 VPWR 182.952
R9995 VPWR.n2780 VPWR 181.273
R9996 VPWR.t975 VPWR 177.916
R9997 VPWR.n2848 VPWR.n2847 166.4
R9998 VPWR.n1770 VPWR.n1768 161.365
R9999 VPWR.n1041 VPWR.n1039 161.365
R10000 VPWR.n1545 VPWR.n1543 161.365
R10001 VPWR.n1550 VPWR.n1548 161.365
R10002 VPWR.n1555 VPWR.n1553 161.365
R10003 VPWR.n1560 VPWR.n1558 161.365
R10004 VPWR.n1565 VPWR.n1563 161.365
R10005 VPWR.n1570 VPWR.n1568 161.365
R10006 VPWR.n1575 VPWR.n1573 161.365
R10007 VPWR.n1580 VPWR.n1578 161.365
R10008 VPWR.n1135 VPWR.n1133 161.365
R10009 VPWR.n1460 VPWR.n1458 161.365
R10010 VPWR.n1455 VPWR.n1453 161.365
R10011 VPWR.n1775 VPWR.n1773 161.365
R10012 VPWR.n1783 VPWR.n1781 161.365
R10013 VPWR.n1779 VPWR.n1777 161.365
R10014 VPWR VPWR.n53 161.363
R10015 VPWR VPWR.n51 161.363
R10016 VPWR VPWR.n49 161.363
R10017 VPWR VPWR.n47 161.363
R10018 VPWR VPWR.n45 161.363
R10019 VPWR VPWR.n43 161.363
R10020 VPWR VPWR.n41 161.363
R10021 VPWR VPWR.n39 161.363
R10022 VPWR VPWR.n37 161.363
R10023 VPWR VPWR.n35 161.363
R10024 VPWR VPWR.n33 161.363
R10025 VPWR VPWR.n31 161.363
R10026 VPWR VPWR.n29 161.363
R10027 VPWR VPWR.n27 161.363
R10028 VPWR VPWR.n25 161.363
R10029 VPWR VPWR.n23 161.363
R10030 VPWR.n1115 VPWR.n1114 161.303
R10031 VPWR.n107 VPWR.n106 161.303
R10032 VPWR.n1120 VPWR.n1119 161.3
R10033 VPWR.n1599 VPWR.n1598 161.3
R10034 VPWR.n1602 VPWR.n1601 161.3
R10035 VPWR.n1111 VPWR.n1110 161.3
R10036 VPWR.n1126 VPWR.n1125 161.3
R10037 VPWR.n1107 VPWR.n1106 161.3
R10038 VPWR.n1612 VPWR.n1611 161.3
R10039 VPWR.n1615 VPWR.n1614 161.3
R10040 VPWR.n1618 VPWR.n1617 161.3
R10041 VPWR.n1623 VPWR.n1622 161.3
R10042 VPWR.n1626 VPWR.n1625 161.3
R10043 VPWR.n1629 VPWR.n1628 161.3
R10044 VPWR.n1101 VPWR.n1100 161.3
R10045 VPWR.n1177 VPWR.n1176 161.3
R10046 VPWR.n1097 VPWR.n1096 161.3
R10047 VPWR.n1639 VPWR.n1638 161.3
R10048 VPWR.n1642 VPWR.n1641 161.3
R10049 VPWR.n1645 VPWR.n1644 161.3
R10050 VPWR.n1650 VPWR.n1649 161.3
R10051 VPWR.n1653 VPWR.n1652 161.3
R10052 VPWR.n1656 VPWR.n1655 161.3
R10053 VPWR.n1091 VPWR.n1090 161.3
R10054 VPWR.n1209 VPWR.n1208 161.3
R10055 VPWR.n1087 VPWR.n1086 161.3
R10056 VPWR.n1666 VPWR.n1665 161.3
R10057 VPWR.n1669 VPWR.n1668 161.3
R10058 VPWR.n1672 VPWR.n1671 161.3
R10059 VPWR.n1677 VPWR.n1676 161.3
R10060 VPWR.n1680 VPWR.n1679 161.3
R10061 VPWR.n1683 VPWR.n1682 161.3
R10062 VPWR.n1081 VPWR.n1080 161.3
R10063 VPWR.n1195 VPWR.n1194 161.3
R10064 VPWR.n1077 VPWR.n1076 161.3
R10065 VPWR.n1693 VPWR.n1692 161.3
R10066 VPWR.n1696 VPWR.n1695 161.3
R10067 VPWR.n1699 VPWR.n1698 161.3
R10068 VPWR.n1704 VPWR.n1703 161.3
R10069 VPWR.n1707 VPWR.n1706 161.3
R10070 VPWR.n1710 VPWR.n1709 161.3
R10071 VPWR.n1070 VPWR.n1069 161.3
R10072 VPWR.n1719 VPWR.n1718 161.3
R10073 VPWR.n1722 VPWR.n1721 161.3
R10074 VPWR.n1717 VPWR.n1716 161.3
R10075 VPWR.n1734 VPWR.n1733 161.3
R10076 VPWR.n1117 VPWR.n1116 161.3
R10077 VPWR.n1731 VPWR.n1730 161.3
R10078 VPWR.n1065 VPWR.n1064 161.3
R10079 VPWR.n126 VPWR.n125 161.3
R10080 VPWR.n117 VPWR.n116 161.3
R10081 VPWR.n120 VPWR.n119 161.3
R10082 VPWR.n115 VPWR.n114 161.3
R10083 VPWR.n138 VPWR.n137 161.3
R10084 VPWR.n128 VPWR.n127 161.3
R10085 VPWR.n109 VPWR.n108 161.3
R10086 VPWR.n105 VPWR.n104 161.3
R10087 VPWR.n288 VPWR.n287 161.3
R10088 VPWR.n285 VPWR.n284 161.3
R10089 VPWR.n101 VPWR.n100 161.3
R10090 VPWR.n272 VPWR.n271 161.3
R10091 VPWR.n275 VPWR.n274 161.3
R10092 VPWR.n270 VPWR.n269 161.3
R10093 VPWR.n260 VPWR.n259 161.3
R10094 VPWR.n263 VPWR.n262 161.3
R10095 VPWR.n258 VPWR.n257 161.3
R10096 VPWR.n248 VPWR.n247 161.3
R10097 VPWR.n251 VPWR.n250 161.3
R10098 VPWR.n246 VPWR.n245 161.3
R10099 VPWR.n236 VPWR.n235 161.3
R10100 VPWR.n239 VPWR.n238 161.3
R10101 VPWR.n234 VPWR.n233 161.3
R10102 VPWR.n224 VPWR.n223 161.3
R10103 VPWR.n227 VPWR.n226 161.3
R10104 VPWR.n222 VPWR.n221 161.3
R10105 VPWR.n212 VPWR.n211 161.3
R10106 VPWR.n215 VPWR.n214 161.3
R10107 VPWR.n210 VPWR.n209 161.3
R10108 VPWR.n200 VPWR.n199 161.3
R10109 VPWR.n203 VPWR.n202 161.3
R10110 VPWR.n198 VPWR.n197 161.3
R10111 VPWR.n188 VPWR.n187 161.3
R10112 VPWR.n191 VPWR.n190 161.3
R10113 VPWR.n186 VPWR.n185 161.3
R10114 VPWR.n176 VPWR.n175 161.3
R10115 VPWR.n179 VPWR.n178 161.3
R10116 VPWR.n174 VPWR.n173 161.3
R10117 VPWR.n164 VPWR.n163 161.3
R10118 VPWR.n167 VPWR.n166 161.3
R10119 VPWR.n162 VPWR.n161 161.3
R10120 VPWR.n152 VPWR.n151 161.3
R10121 VPWR.n155 VPWR.n154 161.3
R10122 VPWR.n150 VPWR.n149 161.3
R10123 VPWR.n140 VPWR.n139 161.3
R10124 VPWR.n143 VPWR.n142 161.3
R10125 VPWR.n131 VPWR.n130 161.3
R10126 VPWR.n1601 VPWR.t46 161.202
R10127 VPWR.n1106 VPWR.t171 161.202
R10128 VPWR.n1617 VPWR.t212 161.202
R10129 VPWR.n1628 VPWR.t320 161.202
R10130 VPWR.n1096 VPWR.t87 161.202
R10131 VPWR.n1644 VPWR.t102 161.202
R10132 VPWR.n1655 VPWR.t325 161.202
R10133 VPWR.n1086 VPWR.t368 161.202
R10134 VPWR.n1671 VPWR.t85 161.202
R10135 VPWR.n1682 VPWR.t238 161.202
R10136 VPWR.n1076 VPWR.t260 161.202
R10137 VPWR.n1698 VPWR.t110 161.202
R10138 VPWR.n1709 VPWR.t136 161.202
R10139 VPWR.n1721 VPWR.t161 161.202
R10140 VPWR.n1116 VPWR.t301 161.202
R10141 VPWR.n1730 VPWR.t12 161.202
R10142 VPWR.n119 VPWR.t128 161.202
R10143 VPWR.n108 VPWR.t27 161.202
R10144 VPWR.n284 VPWR.t163 161.202
R10145 VPWR.n274 VPWR.t293 161.202
R10146 VPWR.n262 VPWR.t333 161.202
R10147 VPWR.n250 VPWR.t57 161.202
R10148 VPWR.n238 VPWR.t201 161.202
R10149 VPWR.n226 VPWR.t225 161.202
R10150 VPWR.n214 VPWR.t62 161.202
R10151 VPWR.n202 VPWR.t97 161.202
R10152 VPWR.n190 VPWR.t199 161.202
R10153 VPWR.n178 VPWR.t360 161.202
R10154 VPWR.n166 VPWR.t379 161.202
R10155 VPWR.n154 VPWR.t233 161.202
R10156 VPWR.n1768 VPWR.t285 161.202
R10157 VPWR.n1039 VPWR.t41 161.202
R10158 VPWR.n1543 VPWR.t22 161.202
R10159 VPWR.n1548 VPWR.t271 161.202
R10160 VPWR.n1553 VPWR.t153 161.202
R10161 VPWR.n1558 VPWR.t123 161.202
R10162 VPWR.n1563 VPWR.t275 161.202
R10163 VPWR.n1568 VPWR.t273 161.202
R10164 VPWR.n1573 VPWR.t118 161.202
R10165 VPWR.n1578 VPWR.t14 161.202
R10166 VPWR.n1133 VPWR.t352 161.202
R10167 VPWR.n1458 VPWR.t223 161.202
R10168 VPWR.n1453 VPWR.t92 161.202
R10169 VPWR.n1773 VPWR.t303 161.202
R10170 VPWR.n1781 VPWR.t341 161.202
R10171 VPWR.n1777 VPWR.t173 161.202
R10172 VPWR.n142 VPWR.t252 161.202
R10173 VPWR.n130 VPWR.t277 161.202
R10174 VPWR.n1119 VPWR.t29 161.106
R10175 VPWR.n1110 VPWR.t165 161.106
R10176 VPWR.n1611 VPWR.t178 161.106
R10177 VPWR.n1622 VPWR.t338 161.106
R10178 VPWR.n1100 VPWR.t59 161.106
R10179 VPWR.n1638 VPWR.t206 161.106
R10180 VPWR.n1649 VPWR.t317 161.106
R10181 VPWR.n1090 VPWR.t354 161.106
R10182 VPWR.n1665 VPWR.t99 161.106
R10183 VPWR.n1676 VPWR.t203 161.106
R10184 VPWR.n1080 VPWR.t362 161.106
R10185 VPWR.n1692 VPWR.t381 161.106
R10186 VPWR.n1703 VPWR.t125 161.106
R10187 VPWR.n1069 VPWR.t254 161.106
R10188 VPWR.n1716 VPWR.t282 161.106
R10189 VPWR.n1064 VPWR.t133 161.106
R10190 VPWR.n125 VPWR.t6 161.106
R10191 VPWR.n114 VPWR.t249 161.106
R10192 VPWR.n137 VPWR.t373 161.106
R10193 VPWR.n104 VPWR.t158 161.106
R10194 VPWR.n100 VPWR.t287 161.106
R10195 VPWR.n269 VPWR.t305 161.106
R10196 VPWR.n257 VPWR.t67 161.106
R10197 VPWR.n245 VPWR.t175 161.106
R10198 VPWR.n233 VPWR.t330 161.106
R10199 VPWR.n221 VPWR.t54 161.106
R10200 VPWR.n209 VPWR.t89 161.106
R10201 VPWR.n197 VPWR.t217 161.106
R10202 VPWR.n185 VPWR.t327 161.106
R10203 VPWR.n173 VPWR.t94 161.106
R10204 VPWR.n161 VPWR.t112 161.106
R10205 VPWR.n149 VPWR.t240 161.106
R10206 VPWR.n53 VPWR.t357 161.106
R10207 VPWR.n51 VPWR.t314 161.106
R10208 VPWR.n49 VPWR.t35 161.106
R10209 VPWR.n47 VPWR.t147 161.106
R10210 VPWR.n45 VPWR.t365 161.106
R10211 VPWR.n43 VPWR.t214 161.106
R10212 VPWR.n41 VPWR.t322 161.106
R10213 VPWR.n39 VPWR.t48 161.106
R10214 VPWR.n37 VPWR.t155 161.106
R10215 VPWR.n35 VPWR.t115 161.106
R10216 VPWR.n33 VPWR.t220 161.106
R10217 VPWR.n31 VPWR.t43 161.106
R10218 VPWR.n29 VPWR.t227 161.106
R10219 VPWR.n27 VPWR.t335 161.106
R10220 VPWR.n25 VPWR.t187 161.106
R10221 VPWR.n23 VPWR.t298 161.106
R10222 VPWR.n1598 VPWR.t79 159.978
R10223 VPWR.n1125 VPWR.t181 159.978
R10224 VPWR.n1614 VPWR.t346 159.978
R10225 VPWR.n1625 VPWR.t64 159.978
R10226 VPWR.n1176 VPWR.t76 159.978
R10227 VPWR.n1641 VPWR.t235 159.978
R10228 VPWR.n1652 VPWR.t343 159.978
R10229 VPWR.n1208 VPWR.t104 159.978
R10230 VPWR.n1668 VPWR.t130 159.978
R10231 VPWR.n1679 VPWR.t257 159.978
R10232 VPWR.n1194 VPWR.t3 159.978
R10233 VPWR.n1695 VPWR.t24 159.978
R10234 VPWR.n1706 VPWR.t262 159.978
R10235 VPWR.n1718 VPWR.t290 159.978
R10236 VPWR.n1733 VPWR.t9 159.978
R10237 VPWR.n1114 VPWR.t311 159.978
R10238 VPWR.n116 VPWR.t144 159.978
R10239 VPWR.n127 VPWR.t19 159.978
R10240 VPWR.n106 VPWR.t51 159.978
R10241 VPWR.n287 VPWR.t196 159.978
R10242 VPWR.n271 VPWR.t308 159.978
R10243 VPWR.n259 VPWR.t73 159.978
R10244 VPWR.n247 VPWR.t184 159.978
R10245 VPWR.n235 VPWR.t193 159.978
R10246 VPWR.n223 VPWR.t349 159.978
R10247 VPWR.n211 VPWR.t70 159.978
R10248 VPWR.n199 VPWR.t230 159.978
R10249 VPWR.n187 VPWR.t246 159.978
R10250 VPWR.n175 VPWR.t376 159.978
R10251 VPWR.n163 VPWR.t120 159.978
R10252 VPWR.n151 VPWR.t150 159.978
R10253 VPWR.n1228 VPWR.t107 159.978
R10254 VPWR.n1150 VPWR.t38 159.978
R10255 VPWR.n1224 VPWR.t243 159.978
R10256 VPWR.n1482 VPWR.t141 159.978
R10257 VPWR.n1170 VPWR.t265 159.978
R10258 VPWR.n1166 VPWR.t16 159.978
R10259 VPWR.n1160 VPWR.t138 159.978
R10260 VPWR.n1476 VPWR.t370 159.978
R10261 VPWR.n1156 VPWR.t279 159.978
R10262 VPWR.n1146 VPWR.t295 159.978
R10263 VPWR.n1469 VPWR.t268 159.978
R10264 VPWR.n1046 VPWR.t168 159.978
R10265 VPWR.n1745 VPWR.t32 159.978
R10266 VPWR.n1033 VPWR.t82 159.978
R10267 VPWR.n1029 VPWR.t190 159.978
R10268 VPWR.n1050 VPWR.t209 159.978
R10269 VPWR.n139 VPWR.t0 159.978
R10270 VPWR.n1229 VPWR.n1228 152
R10271 VPWR.n1151 VPWR.n1150 152
R10272 VPWR.n1225 VPWR.n1224 152
R10273 VPWR.n1483 VPWR.n1482 152
R10274 VPWR.n1171 VPWR.n1170 152
R10275 VPWR.n1167 VPWR.n1166 152
R10276 VPWR.n1161 VPWR.n1160 152
R10277 VPWR.n1477 VPWR.n1476 152
R10278 VPWR.n1157 VPWR.n1156 152
R10279 VPWR.n1147 VPWR.n1146 152
R10280 VPWR.n1470 VPWR.n1469 152
R10281 VPWR.n1047 VPWR.n1046 152
R10282 VPWR.n1746 VPWR.n1745 152
R10283 VPWR.n1034 VPWR.n1033 152
R10284 VPWR.n1030 VPWR.n1029 152
R10285 VPWR.n1051 VPWR.n1050 152
R10286 VPWR.n2845 VPWR.n2844 150.213
R10287 VPWR.n1601 VPWR.t2063 145.137
R10288 VPWR.n1106 VPWR.t2014 145.137
R10289 VPWR.n1617 VPWR.t2000 145.137
R10290 VPWR.n1628 VPWR.t1962 145.137
R10291 VPWR.n1096 VPWR.t2049 145.137
R10292 VPWR.n1644 VPWR.t2042 145.137
R10293 VPWR.n1655 VPWR.t1959 145.137
R10294 VPWR.n1086 VPWR.t1945 145.137
R10295 VPWR.n1671 VPWR.t2050 145.137
R10296 VPWR.n1682 VPWR.t1993 145.137
R10297 VPWR.n1076 VPWR.t1988 145.137
R10298 VPWR.n1698 VPWR.t2040 145.137
R10299 VPWR.n1709 VPWR.t2033 145.137
R10300 VPWR.n1721 VPWR.t2019 145.137
R10301 VPWR.n1116 VPWR.t1969 145.137
R10302 VPWR.n1730 VPWR.t1937 145.137
R10303 VPWR.n119 VPWR.t2048 145.137
R10304 VPWR.n108 VPWR.t1934 145.137
R10305 VPWR.n284 VPWR.t2030 145.137
R10306 VPWR.n274 VPWR.t1983 145.137
R10307 VPWR.n262 VPWR.t1971 145.137
R10308 VPWR.n250 VPWR.t1930 145.137
R10309 VPWR.n238 VPWR.t2016 145.137
R10310 VPWR.n226 VPWR.t2008 145.137
R10311 VPWR.n214 VPWR.t1928 145.137
R10312 VPWR.n202 VPWR.t2057 145.137
R10313 VPWR.n190 VPWR.t2017 145.137
R10314 VPWR.n178 VPWR.t1961 145.137
R10315 VPWR.n166 VPWR.t1952 145.137
R10316 VPWR.n154 VPWR.t2007 145.137
R10317 VPWR.n1768 VPWR.t1976 145.137
R10318 VPWR.n1039 VPWR.t2065 145.137
R10319 VPWR.n1543 VPWR.t1929 145.137
R10320 VPWR.n1548 VPWR.t1986 145.137
R10321 VPWR.n1553 VPWR.t2025 145.137
R10322 VPWR.n1558 VPWR.t2037 145.137
R10323 VPWR.n1563 VPWR.t1979 145.137
R10324 VPWR.n1568 VPWR.t1985 145.137
R10325 VPWR.n1573 VPWR.t2039 145.137
R10326 VPWR.n1578 VPWR.t1936 145.137
R10327 VPWR.n1133 VPWR.t1950 145.137
R10328 VPWR.n1458 VPWR.t1996 145.137
R10329 VPWR.n1453 VPWR.t2045 145.137
R10330 VPWR.n1773 VPWR.t1968 145.137
R10331 VPWR.n1781 VPWR.t1953 145.137
R10332 VPWR.n1777 VPWR.t2013 145.137
R10333 VPWR.n142 VPWR.t1999 145.137
R10334 VPWR.n130 VPWR.t1990 145.137
R10335 VPWR.n1119 VPWR.t2067 145.038
R10336 VPWR.n1110 VPWR.t2018 145.038
R10337 VPWR.n1611 VPWR.t2010 145.038
R10338 VPWR.n1622 VPWR.t1955 145.038
R10339 VPWR.n1100 VPWR.t2059 145.038
R10340 VPWR.n1638 VPWR.t2002 145.038
R10341 VPWR.n1649 VPWR.t1964 145.038
R10342 VPWR.n1090 VPWR.t1949 145.038
R10343 VPWR.n1665 VPWR.t2043 145.038
R10344 VPWR.n1676 VPWR.t2003 145.038
R10345 VPWR.n1080 VPWR.t1947 145.038
R10346 VPWR.n1692 VPWR.t1939 145.038
R10347 VPWR.n1703 VPWR.t2036 145.038
R10348 VPWR.n1069 VPWR.t1989 145.038
R10349 VPWR.n1716 VPWR.t1977 145.038
R10350 VPWR.n1064 VPWR.t2034 145.038
R10351 VPWR.n125 VPWR.t1940 145.038
R10352 VPWR.n114 VPWR.t2001 145.038
R10353 VPWR.n137 VPWR.t1954 145.038
R10354 VPWR.n104 VPWR.t2032 145.038
R10355 VPWR.n100 VPWR.t1987 145.038
R10356 VPWR.n269 VPWR.t1980 145.038
R10357 VPWR.n257 VPWR.t2068 145.038
R10358 VPWR.n245 VPWR.t2027 145.038
R10359 VPWR.n233 VPWR.t1972 145.038
R10360 VPWR.n221 VPWR.t1931 145.038
R10361 VPWR.n209 VPWR.t2060 145.038
R10362 VPWR.n197 VPWR.t2009 145.038
R10363 VPWR.n185 VPWR.t1973 145.038
R10364 VPWR.n173 VPWR.t2058 145.038
R10365 VPWR.n161 VPWR.t2052 145.038
R10366 VPWR.n149 VPWR.t2004 145.038
R10367 VPWR.n53 VPWR.t2053 145.038
R10368 VPWR.n51 VPWR.t1963 145.038
R10369 VPWR.n49 VPWR.t2066 145.038
R10370 VPWR.n47 VPWR.t2026 145.038
R10371 VPWR.n45 VPWR.t1946 145.038
R10372 VPWR.n43 VPWR.t2051 145.038
R10373 VPWR.n41 VPWR.t2069 145.038
R10374 VPWR.n39 VPWR.t2028 145.038
R10375 VPWR.n37 VPWR.t2022 145.038
R10376 VPWR.n35 VPWR.t1943 145.038
R10377 VPWR.n33 VPWR.t1997 145.038
R10378 VPWR.n31 VPWR.t2064 145.038
R10379 VPWR.n29 VPWR.t1995 145.038
R10380 VPWR.n27 VPWR.t1956 145.038
R10381 VPWR.n25 VPWR.t2021 145.038
R10382 VPWR.n23 VPWR.t1970 145.038
R10383 VPWR.n1598 VPWR.t1966 143.911
R10384 VPWR.n1125 VPWR.t2062 143.911
R10385 VPWR.n1614 VPWR.t2047 143.911
R10386 VPWR.n1625 VPWR.t1965 143.911
R10387 VPWR.n1176 VPWR.t1958 143.911
R10388 VPWR.n1641 VPWR.t1944 143.911
R10389 VPWR.n1652 VPWR.t2005 143.911
R10390 VPWR.n1208 VPWR.t1992 143.911
R10391 VPWR.n1668 VPWR.t1941 143.911
R10392 VPWR.n1679 VPWR.t2038 143.911
R10393 VPWR.n1194 VPWR.t2031 143.911
R10394 VPWR.n1695 VPWR.t1978 143.911
R10395 VPWR.n1706 VPWR.t1935 143.911
R10396 VPWR.n1718 VPWR.t2024 143.911
R10397 VPWR.n1733 VPWR.t1984 143.911
R10398 VPWR.n1114 VPWR.t2012 143.911
R10399 VPWR.n116 VPWR.t1951 143.911
R10400 VPWR.n127 VPWR.t1991 143.911
R10401 VPWR.n106 VPWR.t1981 143.911
R10402 VPWR.n287 VPWR.t1933 143.911
R10403 VPWR.n271 VPWR.t2029 143.911
R10404 VPWR.n259 VPWR.t2015 143.911
R10405 VPWR.n247 VPWR.t1932 143.911
R10406 VPWR.n235 VPWR.t1926 143.911
R10407 VPWR.n223 VPWR.t2056 143.911
R10408 VPWR.n211 VPWR.t1974 143.911
R10409 VPWR.n199 VPWR.t1960 143.911
R10410 VPWR.n187 VPWR.t2054 143.911
R10411 VPWR.n175 VPWR.t2006 143.911
R10412 VPWR.n163 VPWR.t1998 143.911
R10413 VPWR.n151 VPWR.t1942 143.911
R10414 VPWR.n1228 VPWR.t1948 143.911
R10415 VPWR.n1150 VPWR.t1975 143.911
R10416 VPWR.n1224 VPWR.t2041 143.911
R10417 VPWR.n1482 VPWR.t1982 143.911
R10418 VPWR.n1170 VPWR.t2035 143.911
R10419 VPWR.n1166 VPWR.t2023 143.911
R10420 VPWR.n1160 VPWR.t1938 143.911
R10421 VPWR.n1476 VPWR.t1994 143.911
R10422 VPWR.n1156 VPWR.t1927 143.911
R10423 VPWR.n1146 VPWR.t2020 143.911
R10424 VPWR.n1469 VPWR.t2044 143.911
R10425 VPWR.n1046 VPWR.t1967 143.911
R10426 VPWR.n1745 VPWR.t2011 143.911
R10427 VPWR.n1033 VPWR.t1957 143.911
R10428 VPWR.n1029 VPWR.t2061 143.911
R10429 VPWR.n1050 VPWR.t2055 143.911
R10430 VPWR.n139 VPWR.t2046 143.911
R10431 VPWR.t441 VPWR.t1420 140.989
R10432 VPWR.t1772 VPWR.t1759 140.989
R10433 VPWR.t1799 VPWR.t1772 140.989
R10434 VPWR.t1775 VPWR.t1799 140.989
R10435 VPWR.t463 VPWR.t1775 140.989
R10436 VPWR.t457 VPWR.t463 140.989
R10437 VPWR.t449 VPWR.t457 140.989
R10438 VPWR.t451 VPWR.t449 140.989
R10439 VPWR.t1744 VPWR.t447 140.989
R10440 VPWR.t1811 VPWR.t1778 140.989
R10441 VPWR.t1765 VPWR.t1811 140.989
R10442 VPWR.t1812 VPWR.t1765 140.989
R10443 VPWR.t572 VPWR.t1812 140.989
R10444 VPWR.t680 VPWR.t572 140.989
R10445 VPWR.t673 VPWR.t680 140.989
R10446 VPWR.t677 VPWR.t673 140.989
R10447 VPWR.t1756 VPWR.t1797 140.989
R10448 VPWR.t1786 VPWR.t1756 140.989
R10449 VPWR.t1760 VPWR.t1786 140.989
R10450 VPWR.t1097 VPWR.t1760 140.989
R10451 VPWR.t1091 VPWR.t1097 140.989
R10452 VPWR.t1099 VPWR.t1091 140.989
R10453 VPWR.t1101 VPWR.t1099 140.989
R10454 VPWR.t1888 VPWR.t1787 140.989
R10455 VPWR.t1757 VPWR.t1800 140.989
R10456 VPWR.t1807 VPWR.t1757 140.989
R10457 VPWR.t1784 VPWR.t1807 140.989
R10458 VPWR.t459 VPWR.t1784 140.989
R10459 VPWR.t453 VPWR.t459 140.989
R10460 VPWR.t461 VPWR.t453 140.989
R10461 VPWR.t455 VPWR.t461 140.989
R10462 VPWR.t1779 VPWR.t1766 140.989
R10463 VPWR.t1753 VPWR.t1779 140.989
R10464 VPWR.t1805 VPWR.t1753 140.989
R10465 VPWR.t576 VPWR.t1805 140.989
R10466 VPWR.t671 VPWR.t576 140.989
R10467 VPWR.t574 VPWR.t671 140.989
R10468 VPWR.t675 VPWR.t574 140.989
R10469 VPWR.t1776 VPWR.t1768 140.989
R10470 VPWR.t1782 VPWR.t1776 140.989
R10471 VPWR.t1770 VPWR.t1782 140.989
R10472 VPWR.t1093 VPWR.t1770 140.989
R10473 VPWR.t1087 VPWR.t1093 140.989
R10474 VPWR.t1095 VPWR.t1087 140.989
R10475 VPWR.t1089 VPWR.t1095 140.989
R10476 VPWR VPWR.n1442 133.312
R10477 VPWR.n2841 VPWR.n2840 129.13
R10478 VPWR.n2858 VPWR.n2819 129.13
R10479 VPWR.n2780 VPWR 127.562
R10480 VPWR.n2760 VPWR 127.562
R10481 VPWR.n2741 VPWR 127.562
R10482 VPWR VPWR.t1818 125.883
R10483 VPWR.n2705 VPWR 125.883
R10484 VPWR.t1746 VPWR.t445 120.849
R10485 VPWR.t1069 VPWR.t1727 117.492
R10486 VPWR.t1670 VPWR.t1290 117.492
R10487 VPWR.t1401 VPWR 115.814
R10488 VPWR VPWR.t451 114.135
R10489 VPWR VPWR.t677 114.135
R10490 VPWR VPWR.t1101 114.135
R10491 VPWR.n2859 VPWR.n2817 111.059
R10492 VPWR.t1536 VPWR 107.421
R10493 VPWR.n1330 VPWR.n1329 106.561
R10494 VPWR.n2781 VPWR.n2780 106.561
R10495 VPWR.n2761 VPWR.n2760 106.561
R10496 VPWR.n2742 VPWR.n2741 106.561
R10497 VPWR.n2706 VPWR.n2705 106.561
R10498 VPWR.n2668 VPWR.n2667 106.561
R10499 VPWR.n2631 VPWR.n2630 106.561
R10500 VPWR VPWR.t1750 106.543
R10501 VPWR VPWR.n1234 104.8
R10502 VPWR VPWR.n1257 104.8
R10503 VPWR VPWR.n1281 104.8
R10504 VPWR VPWR.n1366 104.8
R10505 VPWR VPWR.n1405 104.8
R10506 VPWR.n1443 VPWR 100.883
R10507 VPWR VPWR.t616 100.624
R10508 VPWR.t1403 VPWR.t1041 97.9386
R10509 VPWR.n2859 VPWR.n2858 93.3652
R10510 VPWR.n1231 VPWR.n1230 91.8492
R10511 VPWR.n1153 VPWR.n1152 91.8492
R10512 VPWR.n1227 VPWR.n1226 91.8492
R10513 VPWR.n1485 VPWR.n1484 91.8492
R10514 VPWR.n1173 VPWR.n1172 91.8492
R10515 VPWR.n1169 VPWR.n1168 91.8492
R10516 VPWR.n1163 VPWR.n1162 91.8492
R10517 VPWR.n1479 VPWR.n1478 91.8492
R10518 VPWR.n1159 VPWR.n1158 91.8492
R10519 VPWR.n1149 VPWR.n1148 91.8492
R10520 VPWR.n1472 VPWR.n1471 91.8492
R10521 VPWR.n1049 VPWR.n1048 91.8492
R10522 VPWR.n1748 VPWR.n1747 91.8492
R10523 VPWR.n1036 VPWR.n1035 91.8492
R10524 VPWR.n1032 VPWR.n1031 91.8492
R10525 VPWR.n1053 VPWR.n1052 91.8492
R10526 VPWR.n2847 VPWR.n2820 91.4829
R10527 VPWR.t1403 VPWR.n2842 90.0872
R10528 VPWR.t1803 VPWR 88.7855
R10529 VPWR.n1235 VPWR 79.407
R10530 VPWR.n1258 VPWR 79.407
R10531 VPWR.n1282 VPWR 79.407
R10532 VPWR.n1367 VPWR 79.407
R10533 VPWR.n1406 VPWR 79.407
R10534 VPWR.t928 VPWR.t596 78.8874
R10535 VPWR.n2840 VPWR.n2818 74.9181
R10536 VPWR.n2858 VPWR.n2818 74.9181
R10537 VPWR.n2858 VPWR.n2857 74.9181
R10538 VPWR.n2857 VPWR.n2820 74.9181
R10539 VPWR.t1226 VPWR.t618 70.4952
R10540 VPWR.t618 VPWR.t1228 70.4952
R10541 VPWR.t1228 VPWR.t437 70.4952
R10542 VPWR.t437 VPWR.t863 70.4952
R10543 VPWR.t863 VPWR.t614 70.4952
R10544 VPWR.t614 VPWR.t422 70.4952
R10545 VPWR.t422 VPWR.t441 70.4952
R10546 VPWR.t1791 VPWR.t1888 70.4952
R10547 VPWR.t1894 VPWR.t1791 70.4952
R10548 VPWR.t1763 VPWR.t1894 70.4952
R10549 VPWR.t578 VPWR.t1763 70.4952
R10550 VPWR.t1795 VPWR.t578 70.4952
R10551 VPWR.t1892 VPWR.t1795 70.4952
R10552 VPWR.t1818 VPWR.t1892 70.4952
R10553 VPWR VPWR.t1226 68.8168
R10554 VPWR.t1752 VPWR.t1748 68.8168
R10555 VPWR.t596 VPWR.t1401 62.103
R10556 VPWR VPWR.t1744 60.4245
R10557 VPWR.n2849 VPWR.n2842 59.762
R10558 VPWR.n2845 VPWR.n2819 53.8358
R10559 VPWR.t1748 VPWR.t386 52.0323
R10560 VPWR.t1047 VPWR 50.3539
R10561 VPWR VPWR.t1752 50.3539
R10562 VPWR VPWR.t1746 50.3539
R10563 VPWR.t1800 VPWR 50.3539
R10564 VPWR.t1766 VPWR 50.3539
R10565 VPWR.t1768 VPWR 50.3539
R10566 VPWR.n2854 VPWR.n2818 46.2505
R10567 VPWR.n2855 VPWR.n2854 46.2505
R10568 VPWR.n2835 VPWR.n2834 46.2505
R10569 VPWR.n2836 VPWR.n2835 46.2505
R10570 VPWR.n2838 VPWR.n2837 46.2505
R10571 VPWR.n2837 VPWR.n2836 46.2505
R10572 VPWR.n2844 VPWR.n2824 46.2505
R10573 VPWR.n2857 VPWR.n2856 46.2505
R10574 VPWR.n2856 VPWR.n2855 46.2505
R10575 VPWR.n2849 VPWR.n2848 46.2505
R10576 VPWR.n2846 VPWR.n2845 45.9299
R10577 VPWR.n2832 VPWR.n2830 44.8005
R10578 VPWR.n2830 VPWR.n2826 44.8005
R10579 VPWR.n2847 VPWR.n2843 37.0005
R10580 VPWR.n2843 VPWR.t1041 37.0005
R10581 VPWR.n1230 VPWR.n1229 34.7473
R10582 VPWR.n1152 VPWR.n1151 34.7473
R10583 VPWR.n1226 VPWR.n1225 34.7473
R10584 VPWR.n1484 VPWR.n1483 34.7473
R10585 VPWR.n1172 VPWR.n1171 34.7473
R10586 VPWR.n1168 VPWR.n1167 34.7473
R10587 VPWR.n1162 VPWR.n1161 34.7473
R10588 VPWR.n1478 VPWR.n1477 34.7473
R10589 VPWR.n1158 VPWR.n1157 34.7473
R10590 VPWR.n1148 VPWR.n1147 34.7473
R10591 VPWR.n1471 VPWR.n1470 34.7473
R10592 VPWR.n1048 VPWR.n1047 34.7473
R10593 VPWR.n1747 VPWR.n1746 34.7473
R10594 VPWR.n1035 VPWR.n1034 34.7473
R10595 VPWR.n1031 VPWR.n1030 34.7473
R10596 VPWR.n1052 VPWR.n1051 34.7473
R10597 VPWR.n1299 VPWR.n1298 34.6358
R10598 VPWR.n1357 VPWR.n1341 34.6358
R10599 VPWR.n1362 VPWR.n1361 34.6358
R10600 VPWR.n1396 VPWR.n1380 34.6358
R10601 VPWR.n1401 VPWR.n1400 34.6358
R10602 VPWR.n1411 VPWR.n1377 34.6358
R10603 VPWR.n1433 VPWR.n1417 34.6358
R10604 VPWR.n1438 VPWR.n1437 34.6358
R10605 VPWR.n2755 VPWR.n2754 34.6358
R10606 VPWR.n2721 VPWR.n2713 34.6358
R10607 VPWR.n2728 VPWR.n2727 34.6358
R10608 VPWR.n2685 VPWR.n2676 34.6358
R10609 VPWR.n2688 VPWR.n2687 34.6358
R10610 VPWR.n2692 VPWR.n2691 34.6358
R10611 VPWR.n2648 VPWR.n2639 34.6358
R10612 VPWR.n2651 VPWR.n2650 34.6358
R10613 VPWR.n2655 VPWR.n2654 34.6358
R10614 VPWR.n2662 VPWR.n2661 34.6358
R10615 VPWR.n2615 VPWR.n2611 34.6358
R10616 VPWR.n2619 VPWR.n2603 34.6358
R10617 VPWR.n2622 VPWR.n2621 34.6358
R10618 VPWR.n1316 VPWR.n1315 32.0005
R10619 VPWR.n1353 VPWR.n1352 32.0005
R10620 VPWR.n1392 VPWR.n1391 32.0005
R10621 VPWR.n1429 VPWR.n1428 32.0005
R10622 VPWR.n2717 VPWR.n2716 30.8711
R10623 VPWR.n2681 VPWR.n2680 30.8711
R10624 VPWR.n2644 VPWR.n2643 30.8711
R10625 VPWR.n2610 VPWR.n2609 30.8711
R10626 VPWR.n2834 VPWR.n2832 30.1181
R10627 VPWR.n2838 VPWR.n2826 30.1181
R10628 VPWR.n2848 VPWR.n2846 28.9887
R10629 VPWR.n1325 VPWR.n1324 28.2358
R10630 VPWR.n5 VPWR.t440 26.5955
R10631 VPWR.n5 VPWR.t444 26.5955
R10632 VPWR.n4 VPWR.t617 26.5955
R10633 VPWR.n4 VPWR.t436 26.5955
R10634 VPWR.n1240 VPWR.t1738 26.5955
R10635 VPWR.n1240 VPWR.t1737 26.5955
R10636 VPWR.n1239 VPWR.t1742 26.5955
R10637 VPWR.n1239 VPWR.t581 26.5955
R10638 VPWR.n1245 VPWR.t1734 26.5955
R10639 VPWR.n1245 VPWR.t1739 26.5955
R10640 VPWR.n1238 VPWR.t1057 26.5955
R10641 VPWR.n1238 VPWR.t1060 26.5955
R10642 VPWR.n1263 VPWR.t980 26.5955
R10643 VPWR.n1263 VPWR.t981 26.5955
R10644 VPWR.n1262 VPWR.t498 26.5955
R10645 VPWR.n1262 VPWR.t495 26.5955
R10646 VPWR.n1268 VPWR.t1538 26.5955
R10647 VPWR.n1268 VPWR.t1289 26.5955
R10648 VPWR.n1261 VPWR.t501 26.5955
R10649 VPWR.n1261 VPWR.t499 26.5955
R10650 VPWR.n1287 VPWR.t1405 26.5955
R10651 VPWR.n1287 VPWR.t1412 26.5955
R10652 VPWR.n1286 VPWR.t1209 26.5955
R10653 VPWR.n1286 VPWR.t1208 26.5955
R10654 VPWR.n1292 VPWR.t1409 26.5955
R10655 VPWR.n1292 VPWR.t1406 26.5955
R10656 VPWR.n1285 VPWR.t1212 26.5955
R10657 VPWR.n1285 VPWR.t1210 26.5955
R10658 VPWR.n1314 VPWR.t636 26.5955
R10659 VPWR.n1314 VPWR.t639 26.5955
R10660 VPWR.n1307 VPWR.t442 26.5955
R10661 VPWR.n1307 VPWR.t1421 26.5955
R10662 VPWR.n1321 VPWR.t438 26.5955
R10663 VPWR.n1321 VPWR.t615 26.5955
R10664 VPWR.n1323 VPWR.t1229 26.5955
R10665 VPWR.n1323 VPWR.t864 26.5955
R10666 VPWR.n1351 VPWR.t1416 26.5955
R10667 VPWR.n1351 VPWR.t1419 26.5955
R10668 VPWR.n1350 VPWR.t1398 26.5955
R10669 VPWR.n1350 VPWR.t426 26.5955
R10670 VPWR.n1344 VPWR.t1741 26.5955
R10671 VPWR.n1344 VPWR.t1522 26.5955
R10672 VPWR.n1343 VPWR.t1058 26.5955
R10673 VPWR.n1343 VPWR.t710 26.5955
R10674 VPWR.n1359 VPWR.t1736 26.5955
R10675 VPWR.n1359 VPWR.t1735 26.5955
R10676 VPWR.n1358 VPWR.t582 26.5955
R10677 VPWR.n1358 VPWR.t1059 26.5955
R10678 VPWR.n1390 VPWR.t709 26.5955
R10679 VPWR.n1390 VPWR.t1400 26.5955
R10680 VPWR.n1389 VPWR.t1418 26.5955
R10681 VPWR.n1389 VPWR.t862 26.5955
R10682 VPWR.n1383 VPWR.t1726 26.5955
R10683 VPWR.n1383 VPWR.t643 26.5955
R10684 VPWR.n1382 VPWR.t502 26.5955
R10685 VPWR.n1382 VPWR.t1525 26.5955
R10686 VPWR.n1398 VPWR.t1725 26.5955
R10687 VPWR.n1398 VPWR.t1537 26.5955
R10688 VPWR.n1397 VPWR.t503 26.5955
R10689 VPWR.n1397 VPWR.t500 26.5955
R10690 VPWR.n1427 VPWR.t1225 26.5955
R10691 VPWR.n1427 VPWR.t1520 26.5955
R10692 VPWR.n1426 VPWR.t1399 26.5955
R10693 VPWR.n1426 VPWR.t428 26.5955
R10694 VPWR.n1420 VPWR.t1408 26.5955
R10695 VPWR.n1420 VPWR.t1222 26.5955
R10696 VPWR.n1419 VPWR.t1206 26.5955
R10697 VPWR.n1419 VPWR.t711 26.5955
R10698 VPWR.n1435 VPWR.t1411 26.5955
R10699 VPWR.n1435 VPWR.t1410 26.5955
R10700 VPWR.n1434 VPWR.t1207 26.5955
R10701 VPWR.n1434 VPWR.t1205 26.5955
R10702 VPWR.n2802 VPWR.t694 26.5955
R10703 VPWR.n2802 VPWR.t559 26.5955
R10704 VPWR.n2804 VPWR.t1891 26.5955
R10705 VPWR.n2804 VPWR.t684 26.5955
R10706 VPWR.n2782 VPWR.t464 26.5955
R10707 VPWR.n2782 VPWR.t458 26.5955
R10708 VPWR.n2783 VPWR.t985 26.5955
R10709 VPWR.n2783 VPWR.t1048 26.5955
R10710 VPWR.n2786 VPWR.t450 26.5955
R10711 VPWR.n2786 VPWR.t452 26.5955
R10712 VPWR.n2787 VPWR.t986 26.5955
R10713 VPWR.n2787 VPWR.t830 26.5955
R10714 VPWR.n2762 VPWR.t573 26.5955
R10715 VPWR.n2762 VPWR.t1862 26.5955
R10716 VPWR.n2763 VPWR.t670 26.5955
R10717 VPWR.n2763 VPWR.t681 26.5955
R10718 VPWR.n2766 VPWR.t1907 26.5955
R10719 VPWR.n2766 VPWR.t1906 26.5955
R10720 VPWR.n2767 VPWR.t674 26.5955
R10721 VPWR.n2767 VPWR.t678 26.5955
R10722 VPWR.n2743 VPWR.t1098 26.5955
R10723 VPWR.n2743 VPWR.t1092 26.5955
R10724 VPWR.n2744 VPWR.t1366 26.5955
R10725 VPWR.n2744 VPWR.t1365 26.5955
R10726 VPWR.n2747 VPWR.t1100 26.5955
R10727 VPWR.n2747 VPWR.t1102 26.5955
R10728 VPWR.n2748 VPWR.t1368 26.5955
R10729 VPWR.n2748 VPWR.t1362 26.5955
R10730 VPWR.n2708 VPWR.t1764 26.5955
R10731 VPWR.n2708 VPWR.t1796 26.5955
R10732 VPWR.n2712 VPWR.t1788 26.5955
R10733 VPWR.n2712 VPWR.t1889 26.5955
R10734 VPWR.n2715 VPWR.t1762 26.5955
R10735 VPWR.n2715 VPWR.t1810 26.5955
R10736 VPWR.n2709 VPWR.t1895 26.5955
R10737 VPWR.n2709 VPWR.t579 26.5955
R10738 VPWR.n2679 VPWR.t1758 26.5955
R10739 VPWR.n2679 VPWR.t1808 26.5955
R10740 VPWR.n2678 VPWR.t1774 26.5955
R10741 VPWR.n2678 VPWR.t1820 26.5955
R10742 VPWR.n2675 VPWR.t1785 26.5955
R10743 VPWR.n2675 VPWR.t1000 26.5955
R10744 VPWR.n2674 VPWR.t1802 26.5955
R10745 VPWR.n2674 VPWR.t460 26.5955
R10746 VPWR.n2671 VPWR.t1178 26.5955
R10747 VPWR.n2671 VPWR.t595 26.5955
R10748 VPWR.n2670 VPWR.t454 26.5955
R10749 VPWR.n2670 VPWR.t462 26.5955
R10750 VPWR.n2642 VPWR.t1780 26.5955
R10751 VPWR.n2642 VPWR.t1754 26.5955
R10752 VPWR.n2641 VPWR.t1798 26.5955
R10753 VPWR.n2641 VPWR.t1773 26.5955
R10754 VPWR.n2638 VPWR.t1806 26.5955
R10755 VPWR.n2638 VPWR.t679 26.5955
R10756 VPWR.n2637 VPWR.t1816 26.5955
R10757 VPWR.n2637 VPWR.t577 26.5955
R10758 VPWR.n2634 VPWR.t672 26.5955
R10759 VPWR.n2634 VPWR.t682 26.5955
R10760 VPWR.n2633 VPWR.t1864 26.5955
R10761 VPWR.n2633 VPWR.t575 26.5955
R10762 VPWR.n2606 VPWR.t1777 26.5955
R10763 VPWR.n2606 VPWR.t1783 26.5955
R10764 VPWR.n2605 VPWR.t1813 26.5955
R10765 VPWR.n2605 VPWR.t1794 26.5955
R10766 VPWR.n2613 VPWR.t1789 26.5955
R10767 VPWR.n2613 VPWR.t1367 26.5955
R10768 VPWR.n2612 VPWR.t1771 26.5955
R10769 VPWR.n2612 VPWR.t1094 26.5955
R10770 VPWR.n2602 VPWR.t1369 26.5955
R10771 VPWR.n2602 VPWR.t1363 26.5955
R10772 VPWR.n2601 VPWR.t1088 26.5955
R10773 VPWR.n2601 VPWR.t1096 26.5955
R10774 VPWR.n17 VPWR.n16 25.977
R10775 VPWR.n1253 VPWR.n1252 25.977
R10776 VPWR.n1313 VPWR.n1310 25.977
R10777 VPWR.n1349 VPWR.n1346 25.977
R10778 VPWR.n1372 VPWR.n1338 25.977
R10779 VPWR.n1388 VPWR.n1385 25.977
R10780 VPWR.n1425 VPWR.n1422 25.977
R10781 VPWR.n2811 VPWR.n2810 25.977
R10782 VPWR.n2795 VPWR.n2794 25.977
R10783 VPWR.n2717 VPWR.n2714 25.977
R10784 VPWR.n2681 VPWR.n2677 25.977
R10785 VPWR.n2699 VPWR.n2698 25.977
R10786 VPWR.n2644 VPWR.n2640 25.977
R10787 VPWR.n2609 VPWR.n2607 25.977
R10788 VPWR.n1335 VPWR.n1334 25.224
R10789 VPWR.n2737 VPWR.n2736 25.224
R10790 VPWR.n2722 VPWR.n2721 24.8476
R10791 VPWR.n2686 VPWR.n2685 24.8476
R10792 VPWR.n2649 VPWR.n2648 24.8476
R10793 VPWR.n2615 VPWR.n2614 24.8476
R10794 VPWR.n16 VPWR.n15 24.4711
R10795 VPWR.n1252 VPWR.n1251 24.4711
R10796 VPWR.n1315 VPWR.n1313 24.4711
R10797 VPWR.n1352 VPWR.n1349 24.4711
R10798 VPWR.n1391 VPWR.n1388 24.4711
R10799 VPWR.n1428 VPWR.n1425 24.4711
R10800 VPWR.n2810 VPWR.n2809 24.4711
R10801 VPWR.n2794 VPWR.n2793 24.4711
R10802 VPWR.n11 VPWR.n2 23.7181
R10803 VPWR.n1247 VPWR.n1236 23.7181
R10804 VPWR.n1270 VPWR.n1259 23.7181
R10805 VPWR.n1274 VPWR.n1259 23.7181
R10806 VPWR.n1294 VPWR.n1283 23.7181
R10807 VPWR.n1298 VPWR.n1283 23.7181
R10808 VPWR.n1330 VPWR.n1328 23.7181
R10809 VPWR.n1368 VPWR.n1365 23.7181
R10810 VPWR.n1407 VPWR.n1404 23.7181
R10811 VPWR.n1407 VPWR.n1377 23.7181
R10812 VPWR.n1444 VPWR.n1441 23.7181
R10813 VPWR.n2808 VPWR.n2807 23.7181
R10814 VPWR.n2789 VPWR.n2781 23.7181
R10815 VPWR.n2769 VPWR.n2761 23.7181
R10816 VPWR.n2773 VPWR.n2761 23.7181
R10817 VPWR.n2750 VPWR.n2742 23.7181
R10818 VPWR.n2754 VPWR.n2742 23.7181
R10819 VPWR.n2731 VPWR.n2706 23.7181
R10820 VPWR.n2694 VPWR.n2668 23.7181
R10821 VPWR.n2657 VPWR.n2631 23.7181
R10822 VPWR.n2661 VPWR.n2631 23.7181
R10823 VPWR.n2626 VPWR.n2625 23.7181
R10824 VPWR.t1729 VPWR.t1069 23.4987
R10825 VPWR.t1292 VPWR.t1670 23.4987
R10826 VPWR.n2852 VPWR.n2841 23.1255
R10827 VPWR.n2852 VPWR.t1403 23.1255
R10828 VPWR.n2851 VPWR.n2819 23.1255
R10829 VPWR.t1403 VPWR.n2851 23.1255
R10830 VPWR.n11 VPWR.n10 22.9652
R10831 VPWR.n1247 VPWR.n1246 22.9652
R10832 VPWR.n1270 VPWR.n1269 22.9652
R10833 VPWR.n1294 VPWR.n1293 22.9652
R10834 VPWR.n2807 VPWR.n2803 22.9652
R10835 VPWR.n2789 VPWR.n2788 22.9652
R10836 VPWR.n2769 VPWR.n2768 22.9652
R10837 VPWR.n2750 VPWR.n2749 22.9652
R10838 VPWR.n1320 VPWR.n1308 22.2123
R10839 VPWR.n2724 VPWR.n2723 22.2123
R10840 VPWR.n10 VPWR.n3 21.4593
R10841 VPWR.n1246 VPWR.n1237 21.4593
R10842 VPWR.n1269 VPWR.n1260 21.4593
R10843 VPWR.n1293 VPWR.n1284 21.4593
R10844 VPWR.n1442 VPWR.t427 20.5957
R10845 VPWR.n1443 VPWR.t865 20.5957
R10846 VPWR.n1277 VPWR.n1276 19.9534
R10847 VPWR.n1300 VPWR.n1299 19.9534
R10848 VPWR.n1334 VPWR.n1303 19.9534
R10849 VPWR.n2776 VPWR.n2775 19.9534
R10850 VPWR.n2756 VPWR.n2755 19.9534
R10851 VPWR.n2736 VPWR.n2735 19.9534
R10852 VPWR.n2724 VPWR.n2710 18.824
R10853 VPWR.n2688 VPWR.n2672 18.824
R10854 VPWR.n2651 VPWR.n2635 18.824
R10855 VPWR.n2620 VPWR.n2619 18.824
R10856 VPWR.n1316 VPWR.n1308 18.4476
R10857 VPWR.n1353 VPWR.n1345 18.4476
R10858 VPWR.n1373 VPWR.n1372 18.4476
R10859 VPWR.n1392 VPWR.n1384 18.4476
R10860 VPWR.n1429 VPWR.n1421 18.4476
R10861 VPWR.n2700 VPWR.n2699 18.4476
R10862 VPWR.n1413 VPWR.n1412 17.5829
R10863 VPWR.n2664 VPWR.n2663 17.5829
R10864 VPWR.n6 VPWR.n3 16.9417
R10865 VPWR.n1241 VPWR.n1237 16.9417
R10866 VPWR.n1264 VPWR.n1260 16.9417
R10867 VPWR.n1288 VPWR.n1284 16.9417
R10868 VPWR.n2730 VPWR.n2729 16.5652
R10869 VPWR.n1306 VPWR.n1304 16.1887
R10870 VPWR.n1374 VPWR.n1373 16.1887
R10871 VPWR.n2701 VPWR.n2700 16.1887
R10872 VPWR.n1235 VPWR.t566 16.0935
R10873 VPWR.n1258 VPWR.t637 16.0935
R10874 VPWR.n1282 VPWR.t421 16.0935
R10875 VPWR.n1367 VPWR.t640 16.0935
R10876 VPWR.n1406 VPWR.t642 16.0935
R10877 VPWR.n1234 VPWR.t580 16.0935
R10878 VPWR.n1257 VPWR.t494 16.0935
R10879 VPWR.n1281 VPWR.t584 16.0935
R10880 VPWR.n1366 VPWR.t425 16.0935
R10881 VPWR.n1405 VPWR.t496 16.0935
R10882 VPWR.n1325 VPWR.n1306 15.8123
R10883 VPWR.n2727 VPWR.n2710 15.8123
R10884 VPWR.n2729 VPWR.n2728 15.8123
R10885 VPWR.n2691 VPWR.n2672 15.8123
R10886 VPWR.n2654 VPWR.n2635 15.8123
R10887 VPWR.n2621 VPWR.n2620 15.8123
R10888 VPWR.n1330 VPWR.n1303 13.5534
R10889 VPWR.n2735 VPWR.n2706 13.5534
R10890 VPWR.n2839 VPWR.n2823 13.2148
R10891 VPWR.n2823 VPWR.t570 13.2148
R10892 VPWR.n2827 VPWR.n2817 13.2148
R10893 VPWR.n2827 VPWR.t570 13.2148
R10894 VPWR.n2833 VPWR.n2829 13.2148
R10895 VPWR.n2829 VPWR.t570 13.2148
R10896 VPWR.n15 VPWR.n2 12.8005
R10897 VPWR.n1251 VPWR.n1236 12.8005
R10898 VPWR.n1368 VPWR.n1338 12.8005
R10899 VPWR.n2809 VPWR.n2808 12.8005
R10900 VPWR.n2793 VPWR.n2781 12.8005
R10901 VPWR.n2698 VPWR.n2668 12.8005
R10902 VPWR.n1322 VPWR.n1320 12.424
R10903 VPWR.n1360 VPWR.n1357 12.424
R10904 VPWR.n1399 VPWR.n1396 12.424
R10905 VPWR.n1436 VPWR.n1433 12.424
R10906 VPWR.n1276 VPWR.n1275 10.5417
R10907 VPWR.n1412 VPWR.n1411 10.5417
R10908 VPWR.n2775 VPWR.n2774 10.5417
R10909 VPWR.n2663 VPWR.n2662 10.5417
R10910 VPWR.n2687 VPWR.n2686 9.78874
R10911 VPWR.n2650 VPWR.n2649 9.78874
R10912 VPWR.n2614 VPWR.n2603 9.78874
R10913 VPWR.n1361 VPWR.n1360 9.41227
R10914 VPWR.n1365 VPWR.n1339 9.41227
R10915 VPWR.n1400 VPWR.n1399 9.41227
R10916 VPWR.n1404 VPWR.n1378 9.41227
R10917 VPWR.n1437 VPWR.n1436 9.41227
R10918 VPWR.n1441 VPWR.n1415 9.41227
R10919 VPWR.n2694 VPWR.n2693 9.41227
R10920 VPWR.n2657 VPWR.n2656 9.41227
R10921 VPWR.n2625 VPWR.n2599 9.41227
R10922 VPWR.n1229 VPWR 9.37021
R10923 VPWR.n1151 VPWR 9.37021
R10924 VPWR.n1225 VPWR 9.37021
R10925 VPWR.n1483 VPWR 9.37021
R10926 VPWR.n1171 VPWR 9.37021
R10927 VPWR.n1167 VPWR 9.37021
R10928 VPWR.n1161 VPWR 9.37021
R10929 VPWR.n1477 VPWR 9.37021
R10930 VPWR.n1157 VPWR 9.37021
R10931 VPWR.n1147 VPWR 9.37021
R10932 VPWR.n1470 VPWR 9.37021
R10933 VPWR.n1047 VPWR 9.37021
R10934 VPWR.n1746 VPWR 9.37021
R10935 VPWR.n1034 VPWR 9.37021
R10936 VPWR.n1030 VPWR 9.37021
R10937 VPWR.n1051 VPWR 9.37021
R10938 VPWR.n1467 VPWR.n1466 9.33404
R10939 VPWR.n352 VPWR.n351 9.33404
R10940 VPWR.n1534 VPWR.n1533 9.33404
R10941 VPWR.n348 VPWR.n347 9.33404
R10942 VPWR.n965 VPWR.n964 9.33404
R10943 VPWR.n2479 VPWR.n2478 9.33404
R10944 VPWR.n2475 VPWR.n2474 9.33404
R10945 VPWR.n320 VPWR.n319 9.33404
R10946 VPWR.n973 VPWR.n972 9.33404
R10947 VPWR.n2445 VPWR.n2444 9.33404
R10948 VPWR.n324 VPWR.n323 9.33404
R10949 VPWR.n1891 VPWR.n1890 9.33404
R10950 VPWR.n1887 VPWR.n1886 9.33404
R10951 VPWR.n1881 VPWR.n1880 9.33404
R10952 VPWR.n389 VPWR.n388 9.33404
R10953 VPWR.n393 VPWR.n392 9.33404
R10954 VPWR.n397 VPWR.n396 9.33404
R10955 VPWR.n2455 VPWR.n2454 9.33404
R10956 VPWR.n332 VPWR.n331 9.33404
R10957 VPWR.n1877 VPWR.n1876 9.33404
R10958 VPWR.n405 VPWR.n404 9.33404
R10959 VPWR.n2459 VPWR.n2458 9.33404
R10960 VPWR.n336 VPWR.n335 9.33404
R10961 VPWR.n2308 VPWR.n2307 9.33404
R10962 VPWR.n2312 VPWR.n2311 9.33404
R10963 VPWR.n2318 VPWR.n2317 9.33404
R10964 VPWR.n2322 VPWR.n2321 9.33404
R10965 VPWR.n2332 VPWR.n2331 9.33404
R10966 VPWR.n2338 VPWR.n2337 9.33404
R10967 VPWR.n2342 VPWR.n2341 9.33404
R10968 VPWR.n2348 VPWR.n2347 9.33404
R10969 VPWR.n2352 VPWR.n2351 9.33404
R10970 VPWR.n2358 VPWR.n2357 9.33404
R10971 VPWR.n2362 VPWR.n2361 9.33404
R10972 VPWR.n2368 VPWR.n2367 9.33404
R10973 VPWR.n2372 VPWR.n2371 9.33404
R10974 VPWR.n2378 VPWR.n2377 9.33404
R10975 VPWR.n2381 VPWR.n2380 9.33404
R10976 VPWR.n2328 VPWR.n2327 9.33404
R10977 VPWR.n544 VPWR.n543 9.33404
R10978 VPWR.n540 VPWR.n539 9.33404
R10979 VPWR.n536 VPWR.n535 9.33404
R10980 VPWR.n532 VPWR.n531 9.33404
R10981 VPWR.n524 VPWR.n523 9.33404
R10982 VPWR.n520 VPWR.n519 9.33404
R10983 VPWR.n516 VPWR.n515 9.33404
R10984 VPWR.n512 VPWR.n511 9.33404
R10985 VPWR.n508 VPWR.n507 9.33404
R10986 VPWR.n504 VPWR.n503 9.33404
R10987 VPWR.n500 VPWR.n499 9.33404
R10988 VPWR.n496 VPWR.n495 9.33404
R10989 VPWR.n492 VPWR.n491 9.33404
R10990 VPWR.n488 VPWR.n487 9.33404
R10991 VPWR.n485 VPWR.n484 9.33404
R10992 VPWR.n528 VPWR.n527 9.33404
R10993 VPWR.n2283 VPWR.n2282 9.33404
R10994 VPWR.n2279 VPWR.n2278 9.33404
R10995 VPWR.n2273 VPWR.n2272 9.33404
R10996 VPWR.n2269 VPWR.n2268 9.33404
R10997 VPWR.n2259 VPWR.n2258 9.33404
R10998 VPWR.n2253 VPWR.n2252 9.33404
R10999 VPWR.n2249 VPWR.n2248 9.33404
R11000 VPWR.n2243 VPWR.n2242 9.33404
R11001 VPWR.n2239 VPWR.n2238 9.33404
R11002 VPWR.n2233 VPWR.n2232 9.33404
R11003 VPWR.n2229 VPWR.n2228 9.33404
R11004 VPWR.n2223 VPWR.n2222 9.33404
R11005 VPWR.n2219 VPWR.n2218 9.33404
R11006 VPWR.n2213 VPWR.n2212 9.33404
R11007 VPWR.n2210 VPWR.n2209 9.33404
R11008 VPWR.n2263 VPWR.n2262 9.33404
R11009 VPWR.n581 VPWR.n580 9.33404
R11010 VPWR.n585 VPWR.n584 9.33404
R11011 VPWR.n589 VPWR.n588 9.33404
R11012 VPWR.n593 VPWR.n592 9.33404
R11013 VPWR.n601 VPWR.n600 9.33404
R11014 VPWR.n605 VPWR.n604 9.33404
R11015 VPWR.n609 VPWR.n608 9.33404
R11016 VPWR.n613 VPWR.n612 9.33404
R11017 VPWR.n617 VPWR.n616 9.33404
R11018 VPWR.n621 VPWR.n620 9.33404
R11019 VPWR.n625 VPWR.n624 9.33404
R11020 VPWR.n629 VPWR.n628 9.33404
R11021 VPWR.n633 VPWR.n632 9.33404
R11022 VPWR.n637 VPWR.n636 9.33404
R11023 VPWR.n640 VPWR.n639 9.33404
R11024 VPWR.n597 VPWR.n596 9.33404
R11025 VPWR.n2112 VPWR.n2111 9.33404
R11026 VPWR.n2116 VPWR.n2115 9.33404
R11027 VPWR.n2122 VPWR.n2121 9.33404
R11028 VPWR.n2126 VPWR.n2125 9.33404
R11029 VPWR.n2136 VPWR.n2135 9.33404
R11030 VPWR.n2142 VPWR.n2141 9.33404
R11031 VPWR.n2146 VPWR.n2145 9.33404
R11032 VPWR.n2152 VPWR.n2151 9.33404
R11033 VPWR.n2156 VPWR.n2155 9.33404
R11034 VPWR.n2162 VPWR.n2161 9.33404
R11035 VPWR.n2166 VPWR.n2165 9.33404
R11036 VPWR.n2172 VPWR.n2171 9.33404
R11037 VPWR.n2176 VPWR.n2175 9.33404
R11038 VPWR.n2182 VPWR.n2181 9.33404
R11039 VPWR.n2185 VPWR.n2184 9.33404
R11040 VPWR.n2132 VPWR.n2131 9.33404
R11041 VPWR.n736 VPWR.n735 9.33404
R11042 VPWR.n732 VPWR.n731 9.33404
R11043 VPWR.n728 VPWR.n727 9.33404
R11044 VPWR.n724 VPWR.n723 9.33404
R11045 VPWR.n716 VPWR.n715 9.33404
R11046 VPWR.n712 VPWR.n711 9.33404
R11047 VPWR.n708 VPWR.n707 9.33404
R11048 VPWR.n704 VPWR.n703 9.33404
R11049 VPWR.n700 VPWR.n699 9.33404
R11050 VPWR.n696 VPWR.n695 9.33404
R11051 VPWR.n692 VPWR.n691 9.33404
R11052 VPWR.n688 VPWR.n687 9.33404
R11053 VPWR.n684 VPWR.n683 9.33404
R11054 VPWR.n680 VPWR.n679 9.33404
R11055 VPWR.n677 VPWR.n676 9.33404
R11056 VPWR.n720 VPWR.n719 9.33404
R11057 VPWR.n2087 VPWR.n2086 9.33404
R11058 VPWR.n2083 VPWR.n2082 9.33404
R11059 VPWR.n2077 VPWR.n2076 9.33404
R11060 VPWR.n2073 VPWR.n2072 9.33404
R11061 VPWR.n2063 VPWR.n2062 9.33404
R11062 VPWR.n2057 VPWR.n2056 9.33404
R11063 VPWR.n2053 VPWR.n2052 9.33404
R11064 VPWR.n2047 VPWR.n2046 9.33404
R11065 VPWR.n2043 VPWR.n2042 9.33404
R11066 VPWR.n2037 VPWR.n2036 9.33404
R11067 VPWR.n2033 VPWR.n2032 9.33404
R11068 VPWR.n2027 VPWR.n2026 9.33404
R11069 VPWR.n2023 VPWR.n2022 9.33404
R11070 VPWR.n2017 VPWR.n2016 9.33404
R11071 VPWR.n2014 VPWR.n2013 9.33404
R11072 VPWR.n2067 VPWR.n2066 9.33404
R11073 VPWR.n773 VPWR.n772 9.33404
R11074 VPWR.n777 VPWR.n776 9.33404
R11075 VPWR.n781 VPWR.n780 9.33404
R11076 VPWR.n785 VPWR.n784 9.33404
R11077 VPWR.n793 VPWR.n792 9.33404
R11078 VPWR.n797 VPWR.n796 9.33404
R11079 VPWR.n801 VPWR.n800 9.33404
R11080 VPWR.n805 VPWR.n804 9.33404
R11081 VPWR.n809 VPWR.n808 9.33404
R11082 VPWR.n813 VPWR.n812 9.33404
R11083 VPWR.n817 VPWR.n816 9.33404
R11084 VPWR.n821 VPWR.n820 9.33404
R11085 VPWR.n825 VPWR.n824 9.33404
R11086 VPWR.n829 VPWR.n828 9.33404
R11087 VPWR.n832 VPWR.n831 9.33404
R11088 VPWR.n789 VPWR.n788 9.33404
R11089 VPWR.n1916 VPWR.n1915 9.33404
R11090 VPWR.n1920 VPWR.n1919 9.33404
R11091 VPWR.n1926 VPWR.n1925 9.33404
R11092 VPWR.n1930 VPWR.n1929 9.33404
R11093 VPWR.n1940 VPWR.n1939 9.33404
R11094 VPWR.n1946 VPWR.n1945 9.33404
R11095 VPWR.n1950 VPWR.n1949 9.33404
R11096 VPWR.n1956 VPWR.n1955 9.33404
R11097 VPWR.n1960 VPWR.n1959 9.33404
R11098 VPWR.n1966 VPWR.n1965 9.33404
R11099 VPWR.n1970 VPWR.n1969 9.33404
R11100 VPWR.n1976 VPWR.n1975 9.33404
R11101 VPWR.n1980 VPWR.n1979 9.33404
R11102 VPWR.n1986 VPWR.n1985 9.33404
R11103 VPWR.n1989 VPWR.n1988 9.33404
R11104 VPWR.n1936 VPWR.n1935 9.33404
R11105 VPWR.n928 VPWR.n927 9.33404
R11106 VPWR.n924 VPWR.n923 9.33404
R11107 VPWR.n920 VPWR.n919 9.33404
R11108 VPWR.n916 VPWR.n915 9.33404
R11109 VPWR.n908 VPWR.n907 9.33404
R11110 VPWR.n904 VPWR.n903 9.33404
R11111 VPWR.n900 VPWR.n899 9.33404
R11112 VPWR.n896 VPWR.n895 9.33404
R11113 VPWR.n892 VPWR.n891 9.33404
R11114 VPWR.n888 VPWR.n887 9.33404
R11115 VPWR.n884 VPWR.n883 9.33404
R11116 VPWR.n880 VPWR.n879 9.33404
R11117 VPWR.n876 VPWR.n875 9.33404
R11118 VPWR.n872 VPWR.n871 9.33404
R11119 VPWR.n869 VPWR.n868 9.33404
R11120 VPWR.n912 VPWR.n911 9.33404
R11121 VPWR.n1871 VPWR.n1870 9.33404
R11122 VPWR.n981 VPWR.n980 9.33404
R11123 VPWR.n1495 VPWR.n1494 9.33404
R11124 VPWR.n401 VPWR.n400 9.33404
R11125 VPWR.n2465 VPWR.n2464 9.33404
R11126 VPWR.n340 VPWR.n339 9.33404
R11127 VPWR.n977 VPWR.n976 9.33404
R11128 VPWR.n1491 VPWR.n1490 9.33404
R11129 VPWR.n1867 VPWR.n1866 9.33404
R11130 VPWR.n985 VPWR.n984 9.33404
R11131 VPWR.n1505 VPWR.n1504 9.33404
R11132 VPWR.n409 VPWR.n408 9.33404
R11133 VPWR.n417 VPWR.n416 9.33404
R11134 VPWR.n421 VPWR.n420 9.33404
R11135 VPWR.n425 VPWR.n424 9.33404
R11136 VPWR.n429 VPWR.n428 9.33404
R11137 VPWR.n433 VPWR.n432 9.33404
R11138 VPWR.n437 VPWR.n436 9.33404
R11139 VPWR.n441 VPWR.n440 9.33404
R11140 VPWR.n445 VPWR.n444 9.33404
R11141 VPWR.n448 VPWR.n447 9.33404
R11142 VPWR.n413 VPWR.n412 9.33404
R11143 VPWR.n2449 VPWR.n2448 9.33404
R11144 VPWR.n328 VPWR.n327 9.33404
R11145 VPWR.n989 VPWR.n988 9.33404
R11146 VPWR.n1509 VPWR.n1508 9.33404
R11147 VPWR.n1861 VPWR.n1860 9.33404
R11148 VPWR.n1851 VPWR.n1850 9.33404
R11149 VPWR.n1847 VPWR.n1846 9.33404
R11150 VPWR.n1841 VPWR.n1840 9.33404
R11151 VPWR.n1837 VPWR.n1836 9.33404
R11152 VPWR.n1831 VPWR.n1830 9.33404
R11153 VPWR.n1827 VPWR.n1826 9.33404
R11154 VPWR.n1821 VPWR.n1820 9.33404
R11155 VPWR.n1818 VPWR.n1817 9.33404
R11156 VPWR.n1857 VPWR.n1856 9.33404
R11157 VPWR.n993 VPWR.n992 9.33404
R11158 VPWR.n1519 VPWR.n1518 9.33404
R11159 VPWR.n2469 VPWR.n2468 9.33404
R11160 VPWR.n344 VPWR.n343 9.33404
R11161 VPWR.n1480 VPWR.n1130 9.33404
R11162 VPWR.n997 VPWR.n996 9.33404
R11163 VPWR.n1523 VPWR.n1522 9.33404
R11164 VPWR.n2439 VPWR.n2438 9.33404
R11165 VPWR.n2429 VPWR.n2428 9.33404
R11166 VPWR.n2425 VPWR.n2424 9.33404
R11167 VPWR.n2419 VPWR.n2418 9.33404
R11168 VPWR.n2415 VPWR.n2414 9.33404
R11169 VPWR.n2409 VPWR.n2408 9.33404
R11170 VPWR.n2406 VPWR.n2405 9.33404
R11171 VPWR.n2435 VPWR.n2434 9.33404
R11172 VPWR.n316 VPWR.n315 9.33404
R11173 VPWR.n1538 VPWR.n1537 9.33404
R11174 VPWR.n1001 VPWR.n1000 9.33404
R11175 VPWR.n1005 VPWR.n1004 9.33404
R11176 VPWR.n1009 VPWR.n1008 9.33404
R11177 VPWR.n1013 VPWR.n1012 9.33404
R11178 VPWR.n1017 VPWR.n1016 9.33404
R11179 VPWR.n1021 VPWR.n1020 9.33404
R11180 VPWR.n1024 VPWR.n1023 9.33404
R11181 VPWR.n969 VPWR.n968 9.33404
R11182 VPWR.n1474 VPWR.n1473 9.33404
R11183 VPWR.n312 VPWR.n311 9.33404
R11184 VPWR.n1763 VPWR.n1762 9.33404
R11185 VPWR.n308 VPWR.n307 9.33404
R11186 VPWR.n304 VPWR.n303 9.33404
R11187 VPWR.n296 VPWR.n295 9.33404
R11188 VPWR.n293 VPWR.n292 9.33404
R11189 VPWR.n300 VPWR.n299 9.33404
R11190 VPWR.n1751 VPWR.n1750 9.33404
R11191 VPWR.n1790 VPWR.n1789 9.33404
R11192 VPWR.n1793 VPWR.n1792 9.33404
R11193 VPWR.n1759 VPWR.n1758 9.33404
R11194 VPWR.n2714 VPWR 9.32394
R11195 VPWR.n2677 VPWR 9.32394
R11196 VPWR.n2640 VPWR 9.32394
R11197 VPWR VPWR.n2607 9.32394
R11198 VPWR.n18 VPWR.n17 9.3005
R11199 VPWR.n15 VPWR.n14 9.3005
R11200 VPWR.n13 VPWR.n2 9.3005
R11201 VPWR.n10 VPWR.n9 9.3005
R11202 VPWR.n8 VPWR.n3 9.3005
R11203 VPWR.n12 VPWR.n11 9.3005
R11204 VPWR.n16 VPWR.n0 9.3005
R11205 VPWR.n1254 VPWR.n1253 9.3005
R11206 VPWR.n1251 VPWR.n1250 9.3005
R11207 VPWR.n1249 VPWR.n1236 9.3005
R11208 VPWR.n1246 VPWR.n1244 9.3005
R11209 VPWR.n1243 VPWR.n1237 9.3005
R11210 VPWR.n1248 VPWR.n1247 9.3005
R11211 VPWR.n1252 VPWR.n1233 9.3005
R11212 VPWR.n1278 VPWR.n1277 9.3005
R11213 VPWR.n1272 VPWR.n1259 9.3005
R11214 VPWR.n1269 VPWR.n1267 9.3005
R11215 VPWR.n1266 VPWR.n1260 9.3005
R11216 VPWR.n1271 VPWR.n1270 9.3005
R11217 VPWR.n1274 VPWR.n1273 9.3005
R11218 VPWR.n1276 VPWR.n1256 9.3005
R11219 VPWR.n1301 VPWR.n1300 9.3005
R11220 VPWR.n1296 VPWR.n1283 9.3005
R11221 VPWR.n1293 VPWR.n1291 9.3005
R11222 VPWR.n1290 VPWR.n1284 9.3005
R11223 VPWR.n1295 VPWR.n1294 9.3005
R11224 VPWR.n1298 VPWR.n1297 9.3005
R11225 VPWR.n1299 VPWR.n1280 9.3005
R11226 VPWR.n1332 VPWR.n1303 9.3005
R11227 VPWR.n1331 VPWR.n1330 9.3005
R11228 VPWR.n1311 VPWR.n1310 9.3005
R11229 VPWR.n1313 VPWR.n1312 9.3005
R11230 VPWR.n1315 VPWR.n1309 9.3005
R11231 VPWR.n1317 VPWR.n1316 9.3005
R11232 VPWR.n1318 VPWR.n1308 9.3005
R11233 VPWR.n1320 VPWR.n1319 9.3005
R11234 VPWR.n1324 VPWR.n1305 9.3005
R11235 VPWR.n1326 VPWR.n1325 9.3005
R11236 VPWR.n1328 VPWR.n1327 9.3005
R11237 VPWR.n1334 VPWR.n1333 9.3005
R11238 VPWR.n1336 VPWR.n1335 9.3005
R11239 VPWR.n1375 VPWR.n1374 9.3005
R11240 VPWR.n1370 VPWR.n1338 9.3005
R11241 VPWR.n1369 VPWR.n1368 9.3005
R11242 VPWR.n1347 VPWR.n1346 9.3005
R11243 VPWR.n1349 VPWR.n1348 9.3005
R11244 VPWR.n1352 VPWR.n1342 9.3005
R11245 VPWR.n1354 VPWR.n1353 9.3005
R11246 VPWR.n1355 VPWR.n1341 9.3005
R11247 VPWR.n1357 VPWR.n1356 9.3005
R11248 VPWR.n1361 VPWR.n1340 9.3005
R11249 VPWR.n1363 VPWR.n1362 9.3005
R11250 VPWR.n1365 VPWR.n1364 9.3005
R11251 VPWR.n1372 VPWR.n1371 9.3005
R11252 VPWR.n1408 VPWR.n1407 9.3005
R11253 VPWR.n1386 VPWR.n1385 9.3005
R11254 VPWR.n1388 VPWR.n1387 9.3005
R11255 VPWR.n1391 VPWR.n1381 9.3005
R11256 VPWR.n1393 VPWR.n1392 9.3005
R11257 VPWR.n1394 VPWR.n1380 9.3005
R11258 VPWR.n1396 VPWR.n1395 9.3005
R11259 VPWR.n1400 VPWR.n1379 9.3005
R11260 VPWR.n1402 VPWR.n1401 9.3005
R11261 VPWR.n1404 VPWR.n1403 9.3005
R11262 VPWR.n1409 VPWR.n1377 9.3005
R11263 VPWR.n1411 VPWR.n1410 9.3005
R11264 VPWR.n1445 VPWR.n1444 9.3005
R11265 VPWR.n1423 VPWR.n1422 9.3005
R11266 VPWR.n1425 VPWR.n1424 9.3005
R11267 VPWR.n1428 VPWR.n1418 9.3005
R11268 VPWR.n1430 VPWR.n1429 9.3005
R11269 VPWR.n1431 VPWR.n1417 9.3005
R11270 VPWR.n1433 VPWR.n1432 9.3005
R11271 VPWR.n1437 VPWR.n1416 9.3005
R11272 VPWR.n1439 VPWR.n1438 9.3005
R11273 VPWR.n1441 VPWR.n1440 9.3005
R11274 VPWR.n2807 VPWR.n2806 9.3005
R11275 VPWR.n2808 VPWR.n2800 9.3005
R11276 VPWR.n2809 VPWR.n2799 9.3005
R11277 VPWR.n2810 VPWR.n2798 9.3005
R11278 VPWR.n2812 VPWR.n2811 9.3005
R11279 VPWR.n2796 VPWR.n2795 9.3005
R11280 VPWR.n2790 VPWR.n2789 9.3005
R11281 VPWR.n2791 VPWR.n2781 9.3005
R11282 VPWR.n2793 VPWR.n2792 9.3005
R11283 VPWR.n2794 VPWR.n2779 9.3005
R11284 VPWR.n2777 VPWR.n2776 9.3005
R11285 VPWR.n2775 VPWR.n2759 9.3005
R11286 VPWR.n2770 VPWR.n2769 9.3005
R11287 VPWR.n2771 VPWR.n2761 9.3005
R11288 VPWR.n2773 VPWR.n2772 9.3005
R11289 VPWR.n2757 VPWR.n2756 9.3005
R11290 VPWR.n2751 VPWR.n2750 9.3005
R11291 VPWR.n2752 VPWR.n2742 9.3005
R11292 VPWR.n2754 VPWR.n2753 9.3005
R11293 VPWR.n2755 VPWR.n2740 9.3005
R11294 VPWR.n2738 VPWR.n2737 9.3005
R11295 VPWR.n2718 VPWR.n2717 9.3005
R11296 VPWR.n2719 VPWR.n2713 9.3005
R11297 VPWR.n2721 VPWR.n2720 9.3005
R11298 VPWR.n2723 VPWR.n2711 9.3005
R11299 VPWR.n2725 VPWR.n2724 9.3005
R11300 VPWR.n2727 VPWR.n2726 9.3005
R11301 VPWR.n2728 VPWR.n2707 9.3005
R11302 VPWR.n2732 VPWR.n2731 9.3005
R11303 VPWR.n2733 VPWR.n2706 9.3005
R11304 VPWR.n2735 VPWR.n2734 9.3005
R11305 VPWR.n2736 VPWR.n2704 9.3005
R11306 VPWR.n2702 VPWR.n2701 9.3005
R11307 VPWR.n2682 VPWR.n2681 9.3005
R11308 VPWR.n2683 VPWR.n2676 9.3005
R11309 VPWR.n2685 VPWR.n2684 9.3005
R11310 VPWR.n2687 VPWR.n2673 9.3005
R11311 VPWR.n2689 VPWR.n2688 9.3005
R11312 VPWR.n2691 VPWR.n2690 9.3005
R11313 VPWR.n2692 VPWR.n2669 9.3005
R11314 VPWR.n2695 VPWR.n2694 9.3005
R11315 VPWR.n2696 VPWR.n2668 9.3005
R11316 VPWR.n2698 VPWR.n2697 9.3005
R11317 VPWR.n2699 VPWR.n2666 9.3005
R11318 VPWR.n2645 VPWR.n2644 9.3005
R11319 VPWR.n2646 VPWR.n2639 9.3005
R11320 VPWR.n2648 VPWR.n2647 9.3005
R11321 VPWR.n2650 VPWR.n2636 9.3005
R11322 VPWR.n2652 VPWR.n2651 9.3005
R11323 VPWR.n2654 VPWR.n2653 9.3005
R11324 VPWR.n2655 VPWR.n2632 9.3005
R11325 VPWR.n2658 VPWR.n2657 9.3005
R11326 VPWR.n2659 VPWR.n2631 9.3005
R11327 VPWR.n2661 VPWR.n2660 9.3005
R11328 VPWR.n2662 VPWR.n2629 9.3005
R11329 VPWR.n2627 VPWR.n2626 9.3005
R11330 VPWR.n2609 VPWR.n2608 9.3005
R11331 VPWR.n2611 VPWR.n2604 9.3005
R11332 VPWR.n2616 VPWR.n2615 9.3005
R11333 VPWR.n2617 VPWR.n2603 9.3005
R11334 VPWR.n2619 VPWR.n2618 9.3005
R11335 VPWR.n2621 VPWR.n2600 9.3005
R11336 VPWR.n2623 VPWR.n2622 9.3005
R11337 VPWR.n2625 VPWR.n2624 9.3005
R11338 VPWR.n2505 VPWR.n2504 9.3005
R11339 VPWR.n2569 VPWR.n2568 9.3005
R11340 VPWR.n2509 VPWR.n2508 9.3005
R11341 VPWR.n2553 VPWR.n2552 9.3005
R11342 VPWR.n2545 VPWR.n2544 9.3005
R11343 VPWR.n2533 VPWR.n2532 9.3005
R11344 VPWR.n2529 VPWR.n2528 9.3005
R11345 VPWR.n1222 VPWR.n1221 9.3005
R11346 VPWR.n2521 VPWR.n2520 9.3005
R11347 VPWR.n1184 VPWR.n1102 9.3005
R11348 VPWR.n1218 VPWR.n1094 9.3005
R11349 VPWR.n2541 VPWR.n2540 9.3005
R11350 VPWR.n1215 VPWR.n1092 9.3005
R11351 VPWR.n1212 VPWR.n1211 9.3005
R11352 VPWR.n2517 VPWR.n2516 9.3005
R11353 VPWR.n1181 VPWR.n1104 9.3005
R11354 VPWR.n1204 VPWR.n1084 9.3005
R11355 VPWR.n2557 VPWR.n2556 9.3005
R11356 VPWR.n1201 VPWR.n1082 9.3005
R11357 VPWR.n1592 VPWR.n1591 9.3005
R11358 VPWR.n2565 VPWR.n2564 9.3005
R11359 VPWR.n1198 VPWR.n1197 9.3005
R11360 VPWR.n1190 VPWR.n1074 9.3005
R11361 VPWR.n1742 VPWR.n1741 9.3005
R11362 VPWR.n1187 VPWR.n1071 9.3005
R11363 VPWR.n2577 VPWR.n2576 9.3005
R11364 VPWR.n2581 VPWR.n2580 9.3005
R11365 VPWR.n2592 VPWR.n2591 9.3005
R11366 VPWR.n2589 VPWR.n2588 9.3005
R11367 VPWR.n1738 VPWR.n1737 9.3005
R11368 VPWR.n1063 VPWR.n1062 9.3005
R11369 VPWR.n1596 VPWR.n1595 9.3005
R11370 VPWR.n1275 VPWR.n1274 8.28285
R11371 VPWR.n2774 VPWR.n2773 8.28285
R11372 VPWR.n1607 VPWR.n1109 8.25914
R11373 VPWR.n1728 VPWR.n1727 8.25914
R11374 VPWR.n281 VPWR.n113 8.25914
R11375 VPWR.n136 VPWR.n124 8.25914
R11376 VPWR.n1780 VPWR.n1779 7.91351
R11377 VPWR.n1771 VPWR.n1770 7.9105
R11378 VPWR.n1042 VPWR.n1041 7.9105
R11379 VPWR.n1546 VPWR.n1545 7.9105
R11380 VPWR.n1551 VPWR.n1550 7.9105
R11381 VPWR.n1556 VPWR.n1555 7.9105
R11382 VPWR.n1561 VPWR.n1560 7.9105
R11383 VPWR.n1566 VPWR.n1565 7.9105
R11384 VPWR.n1571 VPWR.n1570 7.9105
R11385 VPWR.n1576 VPWR.n1575 7.9105
R11386 VPWR.n1581 VPWR.n1580 7.9105
R11387 VPWR.n1136 VPWR.n1135 7.9105
R11388 VPWR.n1461 VPWR.n1460 7.9105
R11389 VPWR.n1456 VPWR.n1455 7.9105
R11390 VPWR.n1776 VPWR.n1775 7.9105
R11391 VPWR.n1784 VPWR.n1783 7.9105
R11392 VPWR.n282 VPWR.n281 7.9105
R11393 VPWR.n280 VPWR.n279 7.9105
R11394 VPWR.n268 VPWR.n267 7.9105
R11395 VPWR.n256 VPWR.n255 7.9105
R11396 VPWR.n244 VPWR.n243 7.9105
R11397 VPWR.n232 VPWR.n231 7.9105
R11398 VPWR.n220 VPWR.n219 7.9105
R11399 VPWR.n208 VPWR.n207 7.9105
R11400 VPWR.n196 VPWR.n195 7.9105
R11401 VPWR.n184 VPWR.n183 7.9105
R11402 VPWR.n172 VPWR.n171 7.9105
R11403 VPWR.n160 VPWR.n159 7.9105
R11404 VPWR.n148 VPWR.n147 7.9105
R11405 VPWR.n136 VPWR.n135 7.9105
R11406 VPWR.n1727 VPWR.n1726 7.9105
R11407 VPWR.n1715 VPWR.n1714 7.9105
R11408 VPWR.n1701 VPWR.n1068 7.9105
R11409 VPWR.n1690 VPWR.n1689 7.9105
R11410 VPWR.n1688 VPWR.n1687 7.9105
R11411 VPWR.n1674 VPWR.n1079 7.9105
R11412 VPWR.n1663 VPWR.n1662 7.9105
R11413 VPWR.n1661 VPWR.n1660 7.9105
R11414 VPWR.n1647 VPWR.n1089 7.9105
R11415 VPWR.n1636 VPWR.n1635 7.9105
R11416 VPWR.n1634 VPWR.n1633 7.9105
R11417 VPWR.n1620 VPWR.n1099 7.9105
R11418 VPWR.n1609 VPWR.n1608 7.9105
R11419 VPWR.n1607 VPWR.n1606 7.9105
R11420 VPWR.n26 VPWR.n24 7.8627
R11421 VPWR.n7 VPWR.n6 7.56315
R11422 VPWR.n1242 VPWR.n1241 7.56315
R11423 VPWR.n1265 VPWR.n1264 7.56315
R11424 VPWR.n1289 VPWR.n1288 7.56315
R11425 VPWR.n2805 VPWR.n2803 6.4511
R11426 VPWR.n2788 VPWR.n2785 6.4511
R11427 VPWR.n2768 VPWR.n2765 6.4511
R11428 VPWR.n2749 VPWR.n2746 6.4511
R11429 VPWR.n1362 VPWR.n1339 6.4005
R11430 VPWR.n1401 VPWR.n1378 6.4005
R11431 VPWR.n1438 VPWR.n1415 6.4005
R11432 VPWR.n2723 VPWR.n2722 6.4005
R11433 VPWR.n2693 VPWR.n2692 6.4005
R11434 VPWR.n2656 VPWR.n2655 6.4005
R11435 VPWR.n2622 VPWR.n2599 6.4005
R11436 VPWR.n1595 VPWR.n1122 6.04494
R11437 VPWR.n2505 VPWR.n99 6.04494
R11438 VPWR.n1467 VPWR.n1231 6.04494
R11439 VPWR.n351 VPWR.n290 6.04494
R11440 VPWR.n2568 VPWR.n68 6.04494
R11441 VPWR.n1534 VPWR.n1153 6.04494
R11442 VPWR.n348 VPWR.n346 6.04494
R11443 VPWR.n2508 VPWR.n98 6.04494
R11444 VPWR.n965 VPWR.n963 6.04494
R11445 VPWR.n2478 VPWR.n356 6.04494
R11446 VPWR.n2475 VPWR.n357 6.04494
R11447 VPWR.n320 VPWR.n318 6.04494
R11448 VPWR.n2553 VPWR.n75 6.04494
R11449 VPWR.n973 VPWR.n971 6.04494
R11450 VPWR.n2445 VPWR.n369 6.04494
R11451 VPWR.n324 VPWR.n322 6.04494
R11452 VPWR.n2544 VPWR.n80 6.04494
R11453 VPWR.n1890 VPWR.n932 6.04494
R11454 VPWR.n1887 VPWR.n933 6.04494
R11455 VPWR.n1880 VPWR.n936 6.04494
R11456 VPWR.n389 VPWR.n387 6.04494
R11457 VPWR.n393 VPWR.n391 6.04494
R11458 VPWR.n397 VPWR.n395 6.04494
R11459 VPWR.n2455 VPWR.n365 6.04494
R11460 VPWR.n332 VPWR.n330 6.04494
R11461 VPWR.n2532 VPWR.n86 6.04494
R11462 VPWR.n1877 VPWR.n937 6.04494
R11463 VPWR.n405 VPWR.n403 6.04494
R11464 VPWR.n2458 VPWR.n364 6.04494
R11465 VPWR.n336 VPWR.n334 6.04494
R11466 VPWR.n2529 VPWR.n87 6.04494
R11467 VPWR.n2308 VPWR.n481 6.04494
R11468 VPWR.n2311 VPWR.n480 6.04494
R11469 VPWR.n2318 VPWR.n477 6.04494
R11470 VPWR.n2321 VPWR.n476 6.04494
R11471 VPWR.n2331 VPWR.n472 6.04494
R11472 VPWR.n2338 VPWR.n469 6.04494
R11473 VPWR.n2341 VPWR.n468 6.04494
R11474 VPWR.n2348 VPWR.n465 6.04494
R11475 VPWR.n2351 VPWR.n464 6.04494
R11476 VPWR.n2358 VPWR.n461 6.04494
R11477 VPWR.n2361 VPWR.n460 6.04494
R11478 VPWR.n2368 VPWR.n457 6.04494
R11479 VPWR.n2371 VPWR.n456 6.04494
R11480 VPWR.n2378 VPWR.n453 6.04494
R11481 VPWR.n2380 VPWR.n452 6.04494
R11482 VPWR.n2328 VPWR.n473 6.04494
R11483 VPWR.n543 VPWR.n482 6.04494
R11484 VPWR.n540 VPWR.n538 6.04494
R11485 VPWR.n536 VPWR.n534 6.04494
R11486 VPWR.n532 VPWR.n530 6.04494
R11487 VPWR.n524 VPWR.n522 6.04494
R11488 VPWR.n520 VPWR.n518 6.04494
R11489 VPWR.n516 VPWR.n514 6.04494
R11490 VPWR.n512 VPWR.n510 6.04494
R11491 VPWR.n508 VPWR.n506 6.04494
R11492 VPWR.n504 VPWR.n502 6.04494
R11493 VPWR.n500 VPWR.n498 6.04494
R11494 VPWR.n496 VPWR.n494 6.04494
R11495 VPWR.n492 VPWR.n490 6.04494
R11496 VPWR.n488 VPWR.n486 6.04494
R11497 VPWR.n485 VPWR.n483 6.04494
R11498 VPWR.n528 VPWR.n526 6.04494
R11499 VPWR.n2282 VPWR.n548 6.04494
R11500 VPWR.n2279 VPWR.n549 6.04494
R11501 VPWR.n2272 VPWR.n552 6.04494
R11502 VPWR.n2269 VPWR.n553 6.04494
R11503 VPWR.n2259 VPWR.n557 6.04494
R11504 VPWR.n2252 VPWR.n560 6.04494
R11505 VPWR.n2249 VPWR.n561 6.04494
R11506 VPWR.n2242 VPWR.n564 6.04494
R11507 VPWR.n2239 VPWR.n565 6.04494
R11508 VPWR.n2232 VPWR.n568 6.04494
R11509 VPWR.n2229 VPWR.n569 6.04494
R11510 VPWR.n2222 VPWR.n572 6.04494
R11511 VPWR.n2219 VPWR.n573 6.04494
R11512 VPWR.n2212 VPWR.n576 6.04494
R11513 VPWR.n2210 VPWR.n577 6.04494
R11514 VPWR.n2262 VPWR.n556 6.04494
R11515 VPWR.n581 VPWR.n579 6.04494
R11516 VPWR.n585 VPWR.n583 6.04494
R11517 VPWR.n589 VPWR.n587 6.04494
R11518 VPWR.n593 VPWR.n591 6.04494
R11519 VPWR.n601 VPWR.n599 6.04494
R11520 VPWR.n605 VPWR.n603 6.04494
R11521 VPWR.n609 VPWR.n607 6.04494
R11522 VPWR.n613 VPWR.n611 6.04494
R11523 VPWR.n617 VPWR.n615 6.04494
R11524 VPWR.n621 VPWR.n619 6.04494
R11525 VPWR.n625 VPWR.n623 6.04494
R11526 VPWR.n629 VPWR.n627 6.04494
R11527 VPWR.n633 VPWR.n631 6.04494
R11528 VPWR.n637 VPWR.n635 6.04494
R11529 VPWR.n639 VPWR.n578 6.04494
R11530 VPWR.n597 VPWR.n595 6.04494
R11531 VPWR.n2112 VPWR.n673 6.04494
R11532 VPWR.n2115 VPWR.n672 6.04494
R11533 VPWR.n2122 VPWR.n669 6.04494
R11534 VPWR.n2125 VPWR.n668 6.04494
R11535 VPWR.n2135 VPWR.n664 6.04494
R11536 VPWR.n2142 VPWR.n661 6.04494
R11537 VPWR.n2145 VPWR.n660 6.04494
R11538 VPWR.n2152 VPWR.n657 6.04494
R11539 VPWR.n2155 VPWR.n656 6.04494
R11540 VPWR.n2162 VPWR.n653 6.04494
R11541 VPWR.n2165 VPWR.n652 6.04494
R11542 VPWR.n2172 VPWR.n649 6.04494
R11543 VPWR.n2175 VPWR.n648 6.04494
R11544 VPWR.n2182 VPWR.n645 6.04494
R11545 VPWR.n2184 VPWR.n644 6.04494
R11546 VPWR.n2132 VPWR.n665 6.04494
R11547 VPWR.n735 VPWR.n674 6.04494
R11548 VPWR.n732 VPWR.n730 6.04494
R11549 VPWR.n728 VPWR.n726 6.04494
R11550 VPWR.n724 VPWR.n722 6.04494
R11551 VPWR.n716 VPWR.n714 6.04494
R11552 VPWR.n712 VPWR.n710 6.04494
R11553 VPWR.n708 VPWR.n706 6.04494
R11554 VPWR.n704 VPWR.n702 6.04494
R11555 VPWR.n700 VPWR.n698 6.04494
R11556 VPWR.n696 VPWR.n694 6.04494
R11557 VPWR.n692 VPWR.n690 6.04494
R11558 VPWR.n688 VPWR.n686 6.04494
R11559 VPWR.n684 VPWR.n682 6.04494
R11560 VPWR.n680 VPWR.n678 6.04494
R11561 VPWR.n677 VPWR.n675 6.04494
R11562 VPWR.n720 VPWR.n718 6.04494
R11563 VPWR.n2086 VPWR.n740 6.04494
R11564 VPWR.n2083 VPWR.n741 6.04494
R11565 VPWR.n2076 VPWR.n744 6.04494
R11566 VPWR.n2073 VPWR.n745 6.04494
R11567 VPWR.n2063 VPWR.n749 6.04494
R11568 VPWR.n2056 VPWR.n752 6.04494
R11569 VPWR.n2053 VPWR.n753 6.04494
R11570 VPWR.n2046 VPWR.n756 6.04494
R11571 VPWR.n2043 VPWR.n757 6.04494
R11572 VPWR.n2036 VPWR.n760 6.04494
R11573 VPWR.n2033 VPWR.n761 6.04494
R11574 VPWR.n2026 VPWR.n764 6.04494
R11575 VPWR.n2023 VPWR.n765 6.04494
R11576 VPWR.n2016 VPWR.n768 6.04494
R11577 VPWR.n2014 VPWR.n769 6.04494
R11578 VPWR.n2066 VPWR.n748 6.04494
R11579 VPWR.n773 VPWR.n771 6.04494
R11580 VPWR.n777 VPWR.n775 6.04494
R11581 VPWR.n781 VPWR.n779 6.04494
R11582 VPWR.n785 VPWR.n783 6.04494
R11583 VPWR.n793 VPWR.n791 6.04494
R11584 VPWR.n797 VPWR.n795 6.04494
R11585 VPWR.n801 VPWR.n799 6.04494
R11586 VPWR.n805 VPWR.n803 6.04494
R11587 VPWR.n809 VPWR.n807 6.04494
R11588 VPWR.n813 VPWR.n811 6.04494
R11589 VPWR.n817 VPWR.n815 6.04494
R11590 VPWR.n821 VPWR.n819 6.04494
R11591 VPWR.n825 VPWR.n823 6.04494
R11592 VPWR.n829 VPWR.n827 6.04494
R11593 VPWR.n831 VPWR.n770 6.04494
R11594 VPWR.n789 VPWR.n787 6.04494
R11595 VPWR.n1916 VPWR.n865 6.04494
R11596 VPWR.n1919 VPWR.n864 6.04494
R11597 VPWR.n1926 VPWR.n861 6.04494
R11598 VPWR.n1929 VPWR.n860 6.04494
R11599 VPWR.n1939 VPWR.n856 6.04494
R11600 VPWR.n1946 VPWR.n853 6.04494
R11601 VPWR.n1949 VPWR.n852 6.04494
R11602 VPWR.n1956 VPWR.n849 6.04494
R11603 VPWR.n1959 VPWR.n848 6.04494
R11604 VPWR.n1966 VPWR.n845 6.04494
R11605 VPWR.n1969 VPWR.n844 6.04494
R11606 VPWR.n1976 VPWR.n841 6.04494
R11607 VPWR.n1979 VPWR.n840 6.04494
R11608 VPWR.n1986 VPWR.n837 6.04494
R11609 VPWR.n1988 VPWR.n836 6.04494
R11610 VPWR.n1936 VPWR.n857 6.04494
R11611 VPWR.n927 VPWR.n866 6.04494
R11612 VPWR.n924 VPWR.n922 6.04494
R11613 VPWR.n920 VPWR.n918 6.04494
R11614 VPWR.n916 VPWR.n914 6.04494
R11615 VPWR.n908 VPWR.n906 6.04494
R11616 VPWR.n904 VPWR.n902 6.04494
R11617 VPWR.n900 VPWR.n898 6.04494
R11618 VPWR.n896 VPWR.n894 6.04494
R11619 VPWR.n892 VPWR.n890 6.04494
R11620 VPWR.n888 VPWR.n886 6.04494
R11621 VPWR.n884 VPWR.n882 6.04494
R11622 VPWR.n880 VPWR.n878 6.04494
R11623 VPWR.n876 VPWR.n874 6.04494
R11624 VPWR.n872 VPWR.n870 6.04494
R11625 VPWR.n869 VPWR.n867 6.04494
R11626 VPWR.n912 VPWR.n910 6.04494
R11627 VPWR.n1870 VPWR.n940 6.04494
R11628 VPWR.n981 VPWR.n979 6.04494
R11629 VPWR.n1494 VPWR.n1227 6.04494
R11630 VPWR.n1221 VPWR.n1179 6.04494
R11631 VPWR.n401 VPWR.n399 6.04494
R11632 VPWR.n2465 VPWR.n361 6.04494
R11633 VPWR.n340 VPWR.n338 6.04494
R11634 VPWR.n2520 VPWR.n92 6.04494
R11635 VPWR.n977 VPWR.n975 6.04494
R11636 VPWR.n1491 VPWR.n1485 6.04494
R11637 VPWR.n1184 VPWR.n1183 6.04494
R11638 VPWR.n1867 VPWR.n941 6.04494
R11639 VPWR.n985 VPWR.n983 6.04494
R11640 VPWR.n1505 VPWR.n1173 6.04494
R11641 VPWR.n1218 VPWR.n1217 6.04494
R11642 VPWR.n409 VPWR.n407 6.04494
R11643 VPWR.n417 VPWR.n415 6.04494
R11644 VPWR.n421 VPWR.n419 6.04494
R11645 VPWR.n425 VPWR.n423 6.04494
R11646 VPWR.n429 VPWR.n427 6.04494
R11647 VPWR.n433 VPWR.n431 6.04494
R11648 VPWR.n437 VPWR.n435 6.04494
R11649 VPWR.n441 VPWR.n439 6.04494
R11650 VPWR.n445 VPWR.n443 6.04494
R11651 VPWR.n447 VPWR.n386 6.04494
R11652 VPWR.n413 VPWR.n411 6.04494
R11653 VPWR.n2448 VPWR.n368 6.04494
R11654 VPWR.n328 VPWR.n326 6.04494
R11655 VPWR.n2541 VPWR.n81 6.04494
R11656 VPWR.n989 VPWR.n987 6.04494
R11657 VPWR.n1508 VPWR.n1169 6.04494
R11658 VPWR.n1215 VPWR.n1214 6.04494
R11659 VPWR.n1860 VPWR.n944 6.04494
R11660 VPWR.n1850 VPWR.n948 6.04494
R11661 VPWR.n1847 VPWR.n949 6.04494
R11662 VPWR.n1840 VPWR.n952 6.04494
R11663 VPWR.n1837 VPWR.n953 6.04494
R11664 VPWR.n1830 VPWR.n956 6.04494
R11665 VPWR.n1827 VPWR.n957 6.04494
R11666 VPWR.n1820 VPWR.n960 6.04494
R11667 VPWR.n1818 VPWR.n961 6.04494
R11668 VPWR.n1857 VPWR.n945 6.04494
R11669 VPWR.n993 VPWR.n991 6.04494
R11670 VPWR.n1519 VPWR.n1163 6.04494
R11671 VPWR.n1212 VPWR.n1206 6.04494
R11672 VPWR.n2468 VPWR.n360 6.04494
R11673 VPWR.n344 VPWR.n342 6.04494
R11674 VPWR.n2517 VPWR.n93 6.04494
R11675 VPWR.n1480 VPWR.n1479 6.04494
R11676 VPWR.n1181 VPWR.n1180 6.04494
R11677 VPWR.n997 VPWR.n995 6.04494
R11678 VPWR.n1522 VPWR.n1159 6.04494
R11679 VPWR.n1204 VPWR.n1203 6.04494
R11680 VPWR.n2438 VPWR.n372 6.04494
R11681 VPWR.n2428 VPWR.n376 6.04494
R11682 VPWR.n2425 VPWR.n377 6.04494
R11683 VPWR.n2418 VPWR.n380 6.04494
R11684 VPWR.n2415 VPWR.n381 6.04494
R11685 VPWR.n2408 VPWR.n384 6.04494
R11686 VPWR.n2406 VPWR.n385 6.04494
R11687 VPWR.n2435 VPWR.n373 6.04494
R11688 VPWR.n316 VPWR.n314 6.04494
R11689 VPWR.n2556 VPWR.n74 6.04494
R11690 VPWR.n1537 VPWR.n1149 6.04494
R11691 VPWR.n1201 VPWR.n1200 6.04494
R11692 VPWR.n1001 VPWR.n999 6.04494
R11693 VPWR.n1005 VPWR.n1003 6.04494
R11694 VPWR.n1009 VPWR.n1007 6.04494
R11695 VPWR.n1013 VPWR.n1011 6.04494
R11696 VPWR.n1017 VPWR.n1015 6.04494
R11697 VPWR.n1021 VPWR.n1019 6.04494
R11698 VPWR.n1023 VPWR.n962 6.04494
R11699 VPWR.n969 VPWR.n967 6.04494
R11700 VPWR.n1474 VPWR.n1472 6.04494
R11701 VPWR.n1592 VPWR.n1123 6.04494
R11702 VPWR.n312 VPWR.n310 6.04494
R11703 VPWR.n2565 VPWR.n69 6.04494
R11704 VPWR.n1198 VPWR.n1192 6.04494
R11705 VPWR.n1762 VPWR.n1049 6.04494
R11706 VPWR.n1190 VPWR.n1189 6.04494
R11707 VPWR.n308 VPWR.n306 6.04494
R11708 VPWR.n304 VPWR.n302 6.04494
R11709 VPWR.n296 VPWR.n294 6.04494
R11710 VPWR.n293 VPWR.n291 6.04494
R11711 VPWR.n300 VPWR.n298 6.04494
R11712 VPWR.n1741 VPWR.n1058 6.04494
R11713 VPWR.n1750 VPWR.n1748 6.04494
R11714 VPWR.n1790 VPWR.n1036 6.04494
R11715 VPWR.n1792 VPWR.n1032 6.04494
R11716 VPWR.n1759 VPWR.n1053 6.04494
R11717 VPWR.n1187 VPWR.n1186 6.04494
R11718 VPWR.n2577 VPWR.n63 6.04494
R11719 VPWR.n2580 VPWR.n62 6.04494
R11720 VPWR.n2589 VPWR.n57 6.04494
R11721 VPWR.n2591 VPWR.n56 6.04494
R11722 VPWR.n1738 VPWR.n1059 6.04494
R11723 VPWR.n1062 VPWR.n1061 6.04494
R11724 VPWR.n2785 VPWR.n2784 5.39628
R11725 VPWR.n2765 VPWR.n2764 5.39628
R11726 VPWR.n2746 VPWR.n2745 5.39628
R11727 VPWR.n54 VPWR 4.72593
R11728 VPWR.n52 VPWR 4.72593
R11729 VPWR.n50 VPWR 4.72593
R11730 VPWR.n48 VPWR 4.72593
R11731 VPWR.n46 VPWR 4.72593
R11732 VPWR.n44 VPWR 4.72593
R11733 VPWR.n42 VPWR 4.72593
R11734 VPWR.n40 VPWR 4.72593
R11735 VPWR.n38 VPWR 4.72593
R11736 VPWR.n36 VPWR 4.72593
R11737 VPWR.n34 VPWR 4.72593
R11738 VPWR.n32 VPWR 4.72593
R11739 VPWR.n30 VPWR 4.72593
R11740 VPWR.n28 VPWR 4.72593
R11741 VPWR.n26 VPWR 4.72593
R11742 VPWR.n1446 VPWR.n1445 4.55954
R11743 VPWR.n2571 VPWR.n2570 4.5005
R11744 VPWR.n2511 VPWR.n2510 4.5005
R11745 VPWR.n2551 VPWR.n2550 4.5005
R11746 VPWR.n319 VPWR.n77 4.5005
R11747 VPWR.n2547 VPWR.n2546 4.5005
R11748 VPWR.n323 VPWR.n78 4.5005
R11749 VPWR.n2535 VPWR.n2534 4.5005
R11750 VPWR.n331 VPWR.n84 4.5005
R11751 VPWR.n2454 VPWR.n2453 4.5005
R11752 VPWR.n2527 VPWR.n2526 4.5005
R11753 VPWR.n335 VPWR.n89 4.5005
R11754 VPWR.n2460 VPWR.n2459 4.5005
R11755 VPWR.n1498 VPWR.n1223 4.5005
R11756 VPWR.n1497 VPWR.n1495 4.5005
R11757 VPWR.n980 VPWR.n939 4.5005
R11758 VPWR.n1872 VPWR.n1871 4.5005
R11759 VPWR.n911 VPWR.n858 4.5005
R11760 VPWR.n1935 VPWR.n1934 4.5005
R11761 VPWR.n788 VPWR.n747 4.5005
R11762 VPWR.n2068 VPWR.n2067 4.5005
R11763 VPWR.n719 VPWR.n666 4.5005
R11764 VPWR.n2131 VPWR.n2130 4.5005
R11765 VPWR.n596 VPWR.n555 4.5005
R11766 VPWR.n2264 VPWR.n2263 4.5005
R11767 VPWR.n527 VPWR.n474 4.5005
R11768 VPWR.n2327 VPWR.n2326 4.5005
R11769 VPWR.n404 VPWR.n363 4.5005
R11770 VPWR.n2523 VPWR.n2522 4.5005
R11771 VPWR.n339 VPWR.n90 4.5005
R11772 VPWR.n2464 VPWR.n2463 4.5005
R11773 VPWR.n400 VPWR.n362 4.5005
R11774 VPWR.n2323 VPWR.n2322 4.5005
R11775 VPWR.n531 VPWR.n475 4.5005
R11776 VPWR.n2268 VPWR.n2267 4.5005
R11777 VPWR.n592 VPWR.n554 4.5005
R11778 VPWR.n2127 VPWR.n2126 4.5005
R11779 VPWR.n723 VPWR.n667 4.5005
R11780 VPWR.n2072 VPWR.n2071 4.5005
R11781 VPWR.n784 VPWR.n746 4.5005
R11782 VPWR.n1931 VPWR.n1930 4.5005
R11783 VPWR.n915 VPWR.n859 4.5005
R11784 VPWR.n1488 VPWR.n1486 4.5005
R11785 VPWR.n1490 VPWR.n1489 4.5005
R11786 VPWR.n976 VPWR.n938 4.5005
R11787 VPWR.n1876 VPWR.n1875 4.5005
R11788 VPWR.n1501 VPWR.n1174 4.5005
R11789 VPWR.n1504 VPWR.n1503 4.5005
R11790 VPWR.n984 VPWR.n942 4.5005
R11791 VPWR.n1866 VPWR.n1865 4.5005
R11792 VPWR.n907 VPWR.n855 4.5005
R11793 VPWR.n1941 VPWR.n1940 4.5005
R11794 VPWR.n792 VPWR.n750 4.5005
R11795 VPWR.n2062 VPWR.n2061 4.5005
R11796 VPWR.n715 VPWR.n663 4.5005
R11797 VPWR.n2137 VPWR.n2136 4.5005
R11798 VPWR.n600 VPWR.n558 4.5005
R11799 VPWR.n2258 VPWR.n2257 4.5005
R11800 VPWR.n523 VPWR.n471 4.5005
R11801 VPWR.n2333 VPWR.n2332 4.5005
R11802 VPWR.n408 VPWR.n366 4.5005
R11803 VPWR.n2539 VPWR.n2538 4.5005
R11804 VPWR.n327 VPWR.n83 4.5005
R11805 VPWR.n2450 VPWR.n2449 4.5005
R11806 VPWR.n412 VPWR.n367 4.5005
R11807 VPWR.n2337 VPWR.n2336 4.5005
R11808 VPWR.n519 VPWR.n470 4.5005
R11809 VPWR.n2254 VPWR.n2253 4.5005
R11810 VPWR.n604 VPWR.n559 4.5005
R11811 VPWR.n2141 VPWR.n2140 4.5005
R11812 VPWR.n711 VPWR.n662 4.5005
R11813 VPWR.n2058 VPWR.n2057 4.5005
R11814 VPWR.n796 VPWR.n751 4.5005
R11815 VPWR.n1945 VPWR.n1944 4.5005
R11816 VPWR.n903 VPWR.n854 4.5005
R11817 VPWR.n1512 VPWR.n1165 4.5005
R11818 VPWR.n1511 VPWR.n1509 4.5005
R11819 VPWR.n988 VPWR.n943 4.5005
R11820 VPWR.n1862 VPWR.n1861 4.5005
R11821 VPWR.n1515 VPWR.n1164 4.5005
R11822 VPWR.n1518 VPWR.n1517 4.5005
R11823 VPWR.n992 VPWR.n946 4.5005
R11824 VPWR.n1856 VPWR.n1855 4.5005
R11825 VPWR.n899 VPWR.n851 4.5005
R11826 VPWR.n1951 VPWR.n1950 4.5005
R11827 VPWR.n800 VPWR.n754 4.5005
R11828 VPWR.n2052 VPWR.n2051 4.5005
R11829 VPWR.n707 VPWR.n659 4.5005
R11830 VPWR.n2147 VPWR.n2146 4.5005
R11831 VPWR.n608 VPWR.n562 4.5005
R11832 VPWR.n2248 VPWR.n2247 4.5005
R11833 VPWR.n515 VPWR.n467 4.5005
R11834 VPWR.n2343 VPWR.n2342 4.5005
R11835 VPWR.n416 VPWR.n370 4.5005
R11836 VPWR.n2444 VPWR.n2443 4.5005
R11837 VPWR.n2515 VPWR.n2514 4.5005
R11838 VPWR.n343 VPWR.n95 4.5005
R11839 VPWR.n2470 VPWR.n2469 4.5005
R11840 VPWR.n396 VPWR.n359 4.5005
R11841 VPWR.n2317 VPWR.n2316 4.5005
R11842 VPWR.n535 VPWR.n478 4.5005
R11843 VPWR.n2274 VPWR.n2273 4.5005
R11844 VPWR.n588 VPWR.n551 4.5005
R11845 VPWR.n2121 VPWR.n2120 4.5005
R11846 VPWR.n727 VPWR.n670 4.5005
R11847 VPWR.n2078 VPWR.n2077 4.5005
R11848 VPWR.n780 VPWR.n743 4.5005
R11849 VPWR.n1925 VPWR.n1924 4.5005
R11850 VPWR.n919 VPWR.n862 4.5005
R11851 VPWR.n1882 VPWR.n1881 4.5005
R11852 VPWR.n1586 VPWR.n1129 4.5005
R11853 VPWR.n1585 VPWR.n1130 4.5005
R11854 VPWR.n972 VPWR.n935 4.5005
R11855 VPWR.n1526 VPWR.n1155 4.5005
R11856 VPWR.n1525 VPWR.n1523 4.5005
R11857 VPWR.n996 VPWR.n947 4.5005
R11858 VPWR.n1852 VPWR.n1851 4.5005
R11859 VPWR.n895 VPWR.n850 4.5005
R11860 VPWR.n1955 VPWR.n1954 4.5005
R11861 VPWR.n804 VPWR.n755 4.5005
R11862 VPWR.n2048 VPWR.n2047 4.5005
R11863 VPWR.n703 VPWR.n658 4.5005
R11864 VPWR.n2151 VPWR.n2150 4.5005
R11865 VPWR.n612 VPWR.n563 4.5005
R11866 VPWR.n2244 VPWR.n2243 4.5005
R11867 VPWR.n511 VPWR.n466 4.5005
R11868 VPWR.n2347 VPWR.n2346 4.5005
R11869 VPWR.n420 VPWR.n371 4.5005
R11870 VPWR.n2440 VPWR.n2439 4.5005
R11871 VPWR.n2559 VPWR.n2558 4.5005
R11872 VPWR.n315 VPWR.n72 4.5005
R11873 VPWR.n2434 VPWR.n2433 4.5005
R11874 VPWR.n424 VPWR.n374 4.5005
R11875 VPWR.n2353 VPWR.n2352 4.5005
R11876 VPWR.n507 VPWR.n463 4.5005
R11877 VPWR.n2238 VPWR.n2237 4.5005
R11878 VPWR.n616 VPWR.n566 4.5005
R11879 VPWR.n2157 VPWR.n2156 4.5005
R11880 VPWR.n699 VPWR.n655 4.5005
R11881 VPWR.n2042 VPWR.n2041 4.5005
R11882 VPWR.n808 VPWR.n758 4.5005
R11883 VPWR.n1961 VPWR.n1960 4.5005
R11884 VPWR.n891 VPWR.n847 4.5005
R11885 VPWR.n1846 VPWR.n1845 4.5005
R11886 VPWR.n1145 VPWR.n1144 4.5005
R11887 VPWR.n1539 VPWR.n1538 4.5005
R11888 VPWR.n1000 VPWR.n950 4.5005
R11889 VPWR.n1590 VPWR.n1589 4.5005
R11890 VPWR.n1473 VPWR.n1128 4.5005
R11891 VPWR.n968 VPWR.n934 4.5005
R11892 VPWR.n1886 VPWR.n1885 4.5005
R11893 VPWR.n923 VPWR.n863 4.5005
R11894 VPWR.n1921 VPWR.n1920 4.5005
R11895 VPWR.n776 VPWR.n742 4.5005
R11896 VPWR.n2082 VPWR.n2081 4.5005
R11897 VPWR.n731 VPWR.n671 4.5005
R11898 VPWR.n2117 VPWR.n2116 4.5005
R11899 VPWR.n584 VPWR.n550 4.5005
R11900 VPWR.n2278 VPWR.n2277 4.5005
R11901 VPWR.n539 VPWR.n479 4.5005
R11902 VPWR.n2313 VPWR.n2312 4.5005
R11903 VPWR.n392 VPWR.n358 4.5005
R11904 VPWR.n2474 VPWR.n2473 4.5005
R11905 VPWR.n347 VPWR.n96 4.5005
R11906 VPWR.n2563 VPWR.n2562 4.5005
R11907 VPWR.n311 VPWR.n71 4.5005
R11908 VPWR.n2430 VPWR.n2429 4.5005
R11909 VPWR.n428 VPWR.n375 4.5005
R11910 VPWR.n2357 VPWR.n2356 4.5005
R11911 VPWR.n503 VPWR.n462 4.5005
R11912 VPWR.n2234 VPWR.n2233 4.5005
R11913 VPWR.n620 VPWR.n567 4.5005
R11914 VPWR.n2161 VPWR.n2160 4.5005
R11915 VPWR.n695 VPWR.n654 4.5005
R11916 VPWR.n2038 VPWR.n2037 4.5005
R11917 VPWR.n812 VPWR.n759 4.5005
R11918 VPWR.n1965 VPWR.n1964 4.5005
R11919 VPWR.n887 VPWR.n846 4.5005
R11920 VPWR.n1842 VPWR.n1841 4.5005
R11921 VPWR.n1004 VPWR.n951 4.5005
R11922 VPWR.n1531 VPWR.n1154 4.5005
R11923 VPWR.n1533 VPWR.n1532 4.5005
R11924 VPWR.n1073 VPWR.n1045 4.5005
R11925 VPWR.n1764 VPWR.n1763 4.5005
R11926 VPWR.n1008 VPWR.n954 4.5005
R11927 VPWR.n1836 VPWR.n1835 4.5005
R11928 VPWR.n883 VPWR.n843 4.5005
R11929 VPWR.n1971 VPWR.n1970 4.5005
R11930 VPWR.n816 VPWR.n762 4.5005
R11931 VPWR.n2032 VPWR.n2031 4.5005
R11932 VPWR.n691 VPWR.n651 4.5005
R11933 VPWR.n2167 VPWR.n2166 4.5005
R11934 VPWR.n624 VPWR.n570 4.5005
R11935 VPWR.n2228 VPWR.n2227 4.5005
R11936 VPWR.n499 VPWR.n459 4.5005
R11937 VPWR.n2363 VPWR.n2362 4.5005
R11938 VPWR.n432 VPWR.n378 4.5005
R11939 VPWR.n2424 VPWR.n2423 4.5005
R11940 VPWR.n307 VPWR.n66 4.5005
R11941 VPWR.n299 VPWR.n60 4.5005
R11942 VPWR.n2414 VPWR.n2413 4.5005
R11943 VPWR.n440 VPWR.n382 4.5005
R11944 VPWR.n2373 VPWR.n2372 4.5005
R11945 VPWR.n491 VPWR.n455 4.5005
R11946 VPWR.n2218 VPWR.n2217 4.5005
R11947 VPWR.n632 VPWR.n574 4.5005
R11948 VPWR.n2177 VPWR.n2176 4.5005
R11949 VPWR.n683 VPWR.n647 4.5005
R11950 VPWR.n2022 VPWR.n2021 4.5005
R11951 VPWR.n824 VPWR.n766 4.5005
R11952 VPWR.n1981 VPWR.n1980 4.5005
R11953 VPWR.n875 VPWR.n839 4.5005
R11954 VPWR.n1826 VPWR.n1825 4.5005
R11955 VPWR.n1016 VPWR.n958 4.5005
R11956 VPWR.n1753 VPWR.n1743 4.5005
R11957 VPWR.n1752 VPWR.n1751 4.5005
R11958 VPWR.n1756 VPWR.n1054 4.5005
R11959 VPWR.n1758 VPWR.n1757 4.5005
R11960 VPWR.n1012 VPWR.n955 4.5005
R11961 VPWR.n1832 VPWR.n1831 4.5005
R11962 VPWR.n879 VPWR.n842 4.5005
R11963 VPWR.n1975 VPWR.n1974 4.5005
R11964 VPWR.n820 VPWR.n763 4.5005
R11965 VPWR.n2028 VPWR.n2027 4.5005
R11966 VPWR.n687 VPWR.n650 4.5005
R11967 VPWR.n2171 VPWR.n2170 4.5005
R11968 VPWR.n628 VPWR.n571 4.5005
R11969 VPWR.n2224 VPWR.n2223 4.5005
R11970 VPWR.n495 VPWR.n458 4.5005
R11971 VPWR.n2367 VPWR.n2366 4.5005
R11972 VPWR.n436 VPWR.n379 4.5005
R11973 VPWR.n2420 VPWR.n2419 4.5005
R11974 VPWR.n303 VPWR.n65 4.5005
R11975 VPWR.n2575 VPWR.n2574 4.5005
R11976 VPWR.n2583 VPWR.n2582 4.5005
R11977 VPWR.n2587 VPWR.n2586 4.5005
R11978 VPWR.n295 VPWR.n59 4.5005
R11979 VPWR.n2410 VPWR.n2409 4.5005
R11980 VPWR.n444 VPWR.n383 4.5005
R11981 VPWR.n2377 VPWR.n2376 4.5005
R11982 VPWR.n487 VPWR.n454 4.5005
R11983 VPWR.n2214 VPWR.n2213 4.5005
R11984 VPWR.n636 VPWR.n575 4.5005
R11985 VPWR.n2181 VPWR.n2180 4.5005
R11986 VPWR.n679 VPWR.n646 4.5005
R11987 VPWR.n2018 VPWR.n2017 4.5005
R11988 VPWR.n828 VPWR.n767 4.5005
R11989 VPWR.n1985 VPWR.n1984 4.5005
R11990 VPWR.n871 VPWR.n838 4.5005
R11991 VPWR.n1822 VPWR.n1821 4.5005
R11992 VPWR.n1020 VPWR.n959 4.5005
R11993 VPWR.n1789 VPWR.n1788 4.5005
R11994 VPWR.n1736 VPWR.n1037 4.5005
R11995 VPWR.n1232 VPWR.n1121 4.5005
R11996 VPWR.n1466 VPWR.n1465 4.5005
R11997 VPWR.n964 VPWR.n931 4.5005
R11998 VPWR.n1892 VPWR.n1891 4.5005
R11999 VPWR.n929 VPWR.n928 4.5005
R12000 VPWR.n1915 VPWR.n1914 4.5005
R12001 VPWR.n772 VPWR.n739 4.5005
R12002 VPWR.n2088 VPWR.n2087 4.5005
R12003 VPWR.n737 VPWR.n736 4.5005
R12004 VPWR.n2111 VPWR.n2110 4.5005
R12005 VPWR.n580 VPWR.n547 4.5005
R12006 VPWR.n2284 VPWR.n2283 4.5005
R12007 VPWR.n545 VPWR.n544 4.5005
R12008 VPWR.n2307 VPWR.n2306 4.5005
R12009 VPWR.n388 VPWR.n355 4.5005
R12010 VPWR.n2480 VPWR.n2479 4.5005
R12011 VPWR.n353 VPWR.n352 4.5005
R12012 VPWR.n2503 VPWR.n2502 4.5005
R12013 VPWR.n2594 VPWR.n2593 4.5005
R12014 VPWR.n292 VPWR.n22 4.5005
R12015 VPWR.n2405 VPWR.n2404 4.5005
R12016 VPWR.n449 VPWR.n448 4.5005
R12017 VPWR.n2382 VPWR.n2381 4.5005
R12018 VPWR.n484 VPWR.n451 4.5005
R12019 VPWR.n2209 VPWR.n2208 4.5005
R12020 VPWR.n641 VPWR.n640 4.5005
R12021 VPWR.n2186 VPWR.n2185 4.5005
R12022 VPWR.n676 VPWR.n643 4.5005
R12023 VPWR.n2013 VPWR.n2012 4.5005
R12024 VPWR.n833 VPWR.n832 4.5005
R12025 VPWR.n1990 VPWR.n1989 4.5005
R12026 VPWR.n868 VPWR.n835 4.5005
R12027 VPWR.n1817 VPWR.n1816 4.5005
R12028 VPWR.n1025 VPWR.n1024 4.5005
R12029 VPWR.n1794 VPWR.n1793 4.5005
R12030 VPWR.n1060 VPWR.n1028 4.5005
R12031 VPWR.n2628 VPWR 4.49965
R12032 VPWR.n19 VPWR.n18 4.20017
R12033 VPWR.n1255 VPWR.n1254 4.20017
R12034 VPWR.n1279 VPWR.n1278 4.20017
R12035 VPWR.n1302 VPWR.n1301 4.20017
R12036 VPWR.n1337 VPWR.n1336 4.20017
R12037 VPWR.n1376 VPWR.n1375 4.20017
R12038 VPWR.n1414 VPWR.n1413 4.20017
R12039 VPWR.n2813 VPWR 4.14027
R12040 VPWR.n2797 VPWR 4.14027
R12041 VPWR.n2778 VPWR 4.14027
R12042 VPWR.n2758 VPWR 4.14027
R12043 VPWR.n2739 VPWR 4.14027
R12044 VPWR.n2703 VPWR 4.14027
R12045 VPWR.n2665 VPWR 4.14027
R12046 VPWR.n55 VPWR.n54 4.0005
R12047 VPWR.n2716 VPWR.n2713 3.76521
R12048 VPWR.n2680 VPWR.n2676 3.76521
R12049 VPWR.n2643 VPWR.n2639 3.76521
R12050 VPWR.n2611 VPWR.n2610 3.76521
R12051 VPWR.n1906 VPWR.n858 3.4105
R12052 VPWR.n1934 VPWR.n1933 3.4105
R12053 VPWR.n1997 VPWR.n747 3.4105
R12054 VPWR.n2069 VPWR.n2068 3.4105
R12055 VPWR.n2102 VPWR.n666 3.4105
R12056 VPWR.n2130 VPWR.n2129 3.4105
R12057 VPWR.n2193 VPWR.n555 3.4105
R12058 VPWR.n2265 VPWR.n2264 3.4105
R12059 VPWR.n2298 VPWR.n474 3.4105
R12060 VPWR.n2326 VPWR.n2325 3.4105
R12061 VPWR.n2389 VPWR.n363 3.4105
R12062 VPWR.n2388 VPWR.n362 3.4105
R12063 VPWR.n2324 VPWR.n2323 3.4105
R12064 VPWR.n2299 VPWR.n475 3.4105
R12065 VPWR.n2267 VPWR.n2266 3.4105
R12066 VPWR.n2192 VPWR.n554 3.4105
R12067 VPWR.n2128 VPWR.n2127 3.4105
R12068 VPWR.n2103 VPWR.n667 3.4105
R12069 VPWR.n2071 VPWR.n2070 3.4105
R12070 VPWR.n1996 VPWR.n746 3.4105
R12071 VPWR.n1932 VPWR.n1931 3.4105
R12072 VPWR.n1907 VPWR.n859 3.4105
R12073 VPWR.n1875 VPWR.n1874 3.4105
R12074 VPWR.n1873 VPWR.n1872 3.4105
R12075 VPWR.n1865 VPWR.n1864 3.4105
R12076 VPWR.n1905 VPWR.n855 3.4105
R12077 VPWR.n1942 VPWR.n1941 3.4105
R12078 VPWR.n1998 VPWR.n750 3.4105
R12079 VPWR.n2061 VPWR.n2060 3.4105
R12080 VPWR.n2101 VPWR.n663 3.4105
R12081 VPWR.n2138 VPWR.n2137 3.4105
R12082 VPWR.n2194 VPWR.n558 3.4105
R12083 VPWR.n2257 VPWR.n2256 3.4105
R12084 VPWR.n2297 VPWR.n471 3.4105
R12085 VPWR.n2334 VPWR.n2333 3.4105
R12086 VPWR.n2390 VPWR.n366 3.4105
R12087 VPWR.n2391 VPWR.n367 3.4105
R12088 VPWR.n2336 VPWR.n2335 3.4105
R12089 VPWR.n2296 VPWR.n470 3.4105
R12090 VPWR.n2255 VPWR.n2254 3.4105
R12091 VPWR.n2195 VPWR.n559 3.4105
R12092 VPWR.n2140 VPWR.n2139 3.4105
R12093 VPWR.n2100 VPWR.n662 3.4105
R12094 VPWR.n2059 VPWR.n2058 3.4105
R12095 VPWR.n1999 VPWR.n751 3.4105
R12096 VPWR.n1944 VPWR.n1943 3.4105
R12097 VPWR.n1904 VPWR.n854 3.4105
R12098 VPWR.n1863 VPWR.n1862 3.4105
R12099 VPWR.n1855 VPWR.n1854 3.4105
R12100 VPWR.n1903 VPWR.n851 3.4105
R12101 VPWR.n1952 VPWR.n1951 3.4105
R12102 VPWR.n2000 VPWR.n754 3.4105
R12103 VPWR.n2051 VPWR.n2050 3.4105
R12104 VPWR.n2099 VPWR.n659 3.4105
R12105 VPWR.n2148 VPWR.n2147 3.4105
R12106 VPWR.n2196 VPWR.n562 3.4105
R12107 VPWR.n2247 VPWR.n2246 3.4105
R12108 VPWR.n2295 VPWR.n467 3.4105
R12109 VPWR.n2344 VPWR.n2343 3.4105
R12110 VPWR.n2392 VPWR.n370 3.4105
R12111 VPWR.n2443 VPWR.n2442 3.4105
R12112 VPWR.n2451 VPWR.n2450 3.4105
R12113 VPWR.n2453 VPWR.n2452 3.4105
R12114 VPWR.n2461 VPWR.n2460 3.4105
R12115 VPWR.n2463 VPWR.n2462 3.4105
R12116 VPWR.n2471 VPWR.n2470 3.4105
R12117 VPWR.n2387 VPWR.n359 3.4105
R12118 VPWR.n2316 VPWR.n2315 3.4105
R12119 VPWR.n2300 VPWR.n478 3.4105
R12120 VPWR.n2275 VPWR.n2274 3.4105
R12121 VPWR.n2191 VPWR.n551 3.4105
R12122 VPWR.n2120 VPWR.n2119 3.4105
R12123 VPWR.n2104 VPWR.n670 3.4105
R12124 VPWR.n2079 VPWR.n2078 3.4105
R12125 VPWR.n1995 VPWR.n743 3.4105
R12126 VPWR.n1924 VPWR.n1923 3.4105
R12127 VPWR.n1908 VPWR.n862 3.4105
R12128 VPWR.n1883 VPWR.n1882 3.4105
R12129 VPWR.n1799 VPWR.n935 3.4105
R12130 VPWR.n1800 VPWR.n938 3.4105
R12131 VPWR.n1801 VPWR.n939 3.4105
R12132 VPWR.n1802 VPWR.n942 3.4105
R12133 VPWR.n1803 VPWR.n943 3.4105
R12134 VPWR.n1804 VPWR.n946 3.4105
R12135 VPWR.n1805 VPWR.n947 3.4105
R12136 VPWR.n1853 VPWR.n1852 3.4105
R12137 VPWR.n1902 VPWR.n850 3.4105
R12138 VPWR.n1954 VPWR.n1953 3.4105
R12139 VPWR.n2001 VPWR.n755 3.4105
R12140 VPWR.n2049 VPWR.n2048 3.4105
R12141 VPWR.n2098 VPWR.n658 3.4105
R12142 VPWR.n2150 VPWR.n2149 3.4105
R12143 VPWR.n2197 VPWR.n563 3.4105
R12144 VPWR.n2245 VPWR.n2244 3.4105
R12145 VPWR.n2294 VPWR.n466 3.4105
R12146 VPWR.n2346 VPWR.n2345 3.4105
R12147 VPWR.n2393 VPWR.n371 3.4105
R12148 VPWR.n2441 VPWR.n2440 3.4105
R12149 VPWR.n2433 VPWR.n2432 3.4105
R12150 VPWR.n2394 VPWR.n374 3.4105
R12151 VPWR.n2354 VPWR.n2353 3.4105
R12152 VPWR.n2293 VPWR.n463 3.4105
R12153 VPWR.n2237 VPWR.n2236 3.4105
R12154 VPWR.n2198 VPWR.n566 3.4105
R12155 VPWR.n2158 VPWR.n2157 3.4105
R12156 VPWR.n2097 VPWR.n655 3.4105
R12157 VPWR.n2041 VPWR.n2040 3.4105
R12158 VPWR.n2002 VPWR.n758 3.4105
R12159 VPWR.n1962 VPWR.n1961 3.4105
R12160 VPWR.n1901 VPWR.n847 3.4105
R12161 VPWR.n1845 VPWR.n1844 3.4105
R12162 VPWR.n1806 VPWR.n950 3.4105
R12163 VPWR.n1798 VPWR.n934 3.4105
R12164 VPWR.n1885 VPWR.n1884 3.4105
R12165 VPWR.n1909 VPWR.n863 3.4105
R12166 VPWR.n1922 VPWR.n1921 3.4105
R12167 VPWR.n1994 VPWR.n742 3.4105
R12168 VPWR.n2081 VPWR.n2080 3.4105
R12169 VPWR.n2105 VPWR.n671 3.4105
R12170 VPWR.n2118 VPWR.n2117 3.4105
R12171 VPWR.n2190 VPWR.n550 3.4105
R12172 VPWR.n2277 VPWR.n2276 3.4105
R12173 VPWR.n2301 VPWR.n479 3.4105
R12174 VPWR.n2314 VPWR.n2313 3.4105
R12175 VPWR.n2386 VPWR.n358 3.4105
R12176 VPWR.n2473 VPWR.n2472 3.4105
R12177 VPWR.n2497 VPWR.n96 3.4105
R12178 VPWR.n2496 VPWR.n95 3.4105
R12179 VPWR.n2495 VPWR.n90 3.4105
R12180 VPWR.n2494 VPWR.n89 3.4105
R12181 VPWR.n2493 VPWR.n84 3.4105
R12182 VPWR.n2492 VPWR.n83 3.4105
R12183 VPWR.n2491 VPWR.n78 3.4105
R12184 VPWR.n2490 VPWR.n77 3.4105
R12185 VPWR.n2489 VPWR.n72 3.4105
R12186 VPWR.n2488 VPWR.n71 3.4105
R12187 VPWR.n2431 VPWR.n2430 3.4105
R12188 VPWR.n2395 VPWR.n375 3.4105
R12189 VPWR.n2356 VPWR.n2355 3.4105
R12190 VPWR.n2292 VPWR.n462 3.4105
R12191 VPWR.n2235 VPWR.n2234 3.4105
R12192 VPWR.n2199 VPWR.n567 3.4105
R12193 VPWR.n2160 VPWR.n2159 3.4105
R12194 VPWR.n2096 VPWR.n654 3.4105
R12195 VPWR.n2039 VPWR.n2038 3.4105
R12196 VPWR.n2003 VPWR.n759 3.4105
R12197 VPWR.n1964 VPWR.n1963 3.4105
R12198 VPWR.n1900 VPWR.n846 3.4105
R12199 VPWR.n1843 VPWR.n1842 3.4105
R12200 VPWR.n1807 VPWR.n951 3.4105
R12201 VPWR.n1532 VPWR.n1143 3.4105
R12202 VPWR.n1540 VPWR.n1539 3.4105
R12203 VPWR.n1525 VPWR.n1524 3.4105
R12204 VPWR.n1517 VPWR.n1516 3.4105
R12205 VPWR.n1511 VPWR.n1510 3.4105
R12206 VPWR.n1503 VPWR.n1502 3.4105
R12207 VPWR.n1497 VPWR.n1496 3.4105
R12208 VPWR.n1489 VPWR.n1132 3.4105
R12209 VPWR.n1585 VPWR.n1584 3.4105
R12210 VPWR.n1452 VPWR.n1128 3.4105
R12211 VPWR.n1765 VPWR.n1764 3.4105
R12212 VPWR.n1808 VPWR.n954 3.4105
R12213 VPWR.n1835 VPWR.n1834 3.4105
R12214 VPWR.n1899 VPWR.n843 3.4105
R12215 VPWR.n1972 VPWR.n1971 3.4105
R12216 VPWR.n2004 VPWR.n762 3.4105
R12217 VPWR.n2031 VPWR.n2030 3.4105
R12218 VPWR.n2095 VPWR.n651 3.4105
R12219 VPWR.n2168 VPWR.n2167 3.4105
R12220 VPWR.n2200 VPWR.n570 3.4105
R12221 VPWR.n2227 VPWR.n2226 3.4105
R12222 VPWR.n2291 VPWR.n459 3.4105
R12223 VPWR.n2364 VPWR.n2363 3.4105
R12224 VPWR.n2396 VPWR.n378 3.4105
R12225 VPWR.n2423 VPWR.n2422 3.4105
R12226 VPWR.n2487 VPWR.n66 3.4105
R12227 VPWR.n2485 VPWR.n60 3.4105
R12228 VPWR.n2413 VPWR.n2412 3.4105
R12229 VPWR.n2398 VPWR.n382 3.4105
R12230 VPWR.n2374 VPWR.n2373 3.4105
R12231 VPWR.n2289 VPWR.n455 3.4105
R12232 VPWR.n2217 VPWR.n2216 3.4105
R12233 VPWR.n2202 VPWR.n574 3.4105
R12234 VPWR.n2178 VPWR.n2177 3.4105
R12235 VPWR.n2093 VPWR.n647 3.4105
R12236 VPWR.n2021 VPWR.n2020 3.4105
R12237 VPWR.n2006 VPWR.n766 3.4105
R12238 VPWR.n1982 VPWR.n1981 3.4105
R12239 VPWR.n1897 VPWR.n839 3.4105
R12240 VPWR.n1825 VPWR.n1824 3.4105
R12241 VPWR.n1810 VPWR.n958 3.4105
R12242 VPWR.n1752 VPWR.n1744 3.4105
R12243 VPWR.n1757 VPWR.n1043 3.4105
R12244 VPWR.n1809 VPWR.n955 3.4105
R12245 VPWR.n1833 VPWR.n1832 3.4105
R12246 VPWR.n1898 VPWR.n842 3.4105
R12247 VPWR.n1974 VPWR.n1973 3.4105
R12248 VPWR.n2005 VPWR.n763 3.4105
R12249 VPWR.n2029 VPWR.n2028 3.4105
R12250 VPWR.n2094 VPWR.n650 3.4105
R12251 VPWR.n2170 VPWR.n2169 3.4105
R12252 VPWR.n2201 VPWR.n571 3.4105
R12253 VPWR.n2225 VPWR.n2224 3.4105
R12254 VPWR.n2290 VPWR.n458 3.4105
R12255 VPWR.n2366 VPWR.n2365 3.4105
R12256 VPWR.n2397 VPWR.n379 3.4105
R12257 VPWR.n2421 VPWR.n2420 3.4105
R12258 VPWR.n2486 VPWR.n65 3.4105
R12259 VPWR.n2484 VPWR.n59 3.4105
R12260 VPWR.n2411 VPWR.n2410 3.4105
R12261 VPWR.n2399 VPWR.n383 3.4105
R12262 VPWR.n2376 VPWR.n2375 3.4105
R12263 VPWR.n2288 VPWR.n454 3.4105
R12264 VPWR.n2215 VPWR.n2214 3.4105
R12265 VPWR.n2203 VPWR.n575 3.4105
R12266 VPWR.n2180 VPWR.n2179 3.4105
R12267 VPWR.n2092 VPWR.n646 3.4105
R12268 VPWR.n2019 VPWR.n2018 3.4105
R12269 VPWR.n2007 VPWR.n767 3.4105
R12270 VPWR.n1984 VPWR.n1983 3.4105
R12271 VPWR.n1896 VPWR.n838 3.4105
R12272 VPWR.n1823 VPWR.n1822 3.4105
R12273 VPWR.n1811 VPWR.n959 3.4105
R12274 VPWR.n1788 VPWR.n1787 3.4105
R12275 VPWR.n1465 VPWR.n1464 3.4105
R12276 VPWR.n1797 VPWR.n931 3.4105
R12277 VPWR.n1893 VPWR.n1892 3.4105
R12278 VPWR.n1910 VPWR.n929 3.4105
R12279 VPWR.n1914 VPWR.n1913 3.4105
R12280 VPWR.n1993 VPWR.n739 3.4105
R12281 VPWR.n2089 VPWR.n2088 3.4105
R12282 VPWR.n2106 VPWR.n737 3.4105
R12283 VPWR.n2110 VPWR.n2109 3.4105
R12284 VPWR.n2189 VPWR.n547 3.4105
R12285 VPWR.n2285 VPWR.n2284 3.4105
R12286 VPWR.n2302 VPWR.n545 3.4105
R12287 VPWR.n2306 VPWR.n2305 3.4105
R12288 VPWR.n2385 VPWR.n355 3.4105
R12289 VPWR.n2481 VPWR.n2480 3.4105
R12290 VPWR.n2498 VPWR.n353 3.4105
R12291 VPWR.n2502 VPWR.n2501 3.4105
R12292 VPWR.n2512 VPWR.n2511 3.4105
R12293 VPWR.n2514 VPWR.n2513 3.4105
R12294 VPWR.n2524 VPWR.n2523 3.4105
R12295 VPWR.n2526 VPWR.n2525 3.4105
R12296 VPWR.n2536 VPWR.n2535 3.4105
R12297 VPWR.n2538 VPWR.n2537 3.4105
R12298 VPWR.n2548 VPWR.n2547 3.4105
R12299 VPWR.n2550 VPWR.n2549 3.4105
R12300 VPWR.n2560 VPWR.n2559 3.4105
R12301 VPWR.n2562 VPWR.n2561 3.4105
R12302 VPWR.n2572 VPWR.n2571 3.4105
R12303 VPWR.n2574 VPWR.n2573 3.4105
R12304 VPWR.n2584 VPWR.n2583 3.4105
R12305 VPWR.n2586 VPWR.n2585 3.4105
R12306 VPWR.n2595 VPWR.n2594 3.4105
R12307 VPWR.n2483 VPWR.n22 3.4105
R12308 VPWR.n2404 VPWR.n2403 3.4105
R12309 VPWR.n2400 VPWR.n449 3.4105
R12310 VPWR.n2383 VPWR.n2382 3.4105
R12311 VPWR.n2287 VPWR.n451 3.4105
R12312 VPWR.n2208 VPWR.n2207 3.4105
R12313 VPWR.n2204 VPWR.n641 3.4105
R12314 VPWR.n2187 VPWR.n2186 3.4105
R12315 VPWR.n2091 VPWR.n643 3.4105
R12316 VPWR.n2012 VPWR.n2011 3.4105
R12317 VPWR.n2008 VPWR.n833 3.4105
R12318 VPWR.n1991 VPWR.n1990 3.4105
R12319 VPWR.n1895 VPWR.n835 3.4105
R12320 VPWR.n1816 VPWR.n1815 3.4105
R12321 VPWR.n1812 VPWR.n1025 3.4105
R12322 VPWR.n1795 VPWR.n1794 3.4105
R12323 VPWR.n1055 VPWR.n1028 3.4105
R12324 VPWR.n1056 VPWR.n1037 3.4105
R12325 VPWR.n1754 VPWR.n1753 3.4105
R12326 VPWR.n1756 VPWR.n1755 3.4105
R12327 VPWR.n1529 VPWR.n1045 3.4105
R12328 VPWR.n1531 VPWR.n1530 3.4105
R12329 VPWR.n1528 VPWR.n1145 3.4105
R12330 VPWR.n1527 VPWR.n1526 3.4105
R12331 VPWR.n1515 VPWR.n1514 3.4105
R12332 VPWR.n1513 VPWR.n1512 3.4105
R12333 VPWR.n1501 VPWR.n1500 3.4105
R12334 VPWR.n1499 VPWR.n1498 3.4105
R12335 VPWR.n1488 VPWR.n1487 3.4105
R12336 VPWR.n1587 VPWR.n1586 3.4105
R12337 VPWR.n1589 VPWR.n1588 3.4105
R12338 VPWR.n1448 VPWR.n1232 3.4105
R12339 VPWR.n1345 VPWR.n1341 3.38874
R12340 VPWR.n1384 VPWR.n1380 3.38874
R12341 VPWR.n1421 VPWR.n1417 3.38874
R12342 VPWR.n28 VPWR.n26 3.36211
R12343 VPWR.n30 VPWR.n28 3.36211
R12344 VPWR.n32 VPWR.n30 3.36211
R12345 VPWR.n34 VPWR.n32 3.36211
R12346 VPWR.n36 VPWR.n34 3.36211
R12347 VPWR.n38 VPWR.n36 3.36211
R12348 VPWR.n40 VPWR.n38 3.36211
R12349 VPWR.n42 VPWR.n40 3.36211
R12350 VPWR.n44 VPWR.n42 3.36211
R12351 VPWR.n46 VPWR.n44 3.36211
R12352 VPWR.n48 VPWR.n46 3.36211
R12353 VPWR.n50 VPWR.n48 3.36211
R12354 VPWR.n52 VPWR.n50 3.36211
R12355 VPWR.n54 VPWR.n52 3.36211
R12356 VPWR.t1727 VPWR.t1047 3.35739
R12357 VPWR.t1290 VPWR.t1536 3.35739
R12358 VPWR.n2571 VPWR.n66 3.28012
R12359 VPWR.n2511 VPWR.n96 3.28012
R12360 VPWR.n2550 VPWR.n77 3.28012
R12361 VPWR.n2440 VPWR.n77 3.28012
R12362 VPWR.n2547 VPWR.n78 3.28012
R12363 VPWR.n2443 VPWR.n78 3.28012
R12364 VPWR.n2535 VPWR.n84 3.28012
R12365 VPWR.n2453 VPWR.n84 3.28012
R12366 VPWR.n2453 VPWR.n366 3.28012
R12367 VPWR.n2526 VPWR.n89 3.28012
R12368 VPWR.n2460 VPWR.n89 3.28012
R12369 VPWR.n2460 VPWR.n363 3.28012
R12370 VPWR.n1498 VPWR.n1497 3.28012
R12371 VPWR.n1497 VPWR.n939 3.28012
R12372 VPWR.n1872 VPWR.n939 3.28012
R12373 VPWR.n1872 VPWR.n858 3.28012
R12374 VPWR.n1934 VPWR.n858 3.28012
R12375 VPWR.n1934 VPWR.n747 3.28012
R12376 VPWR.n2068 VPWR.n747 3.28012
R12377 VPWR.n2068 VPWR.n666 3.28012
R12378 VPWR.n2130 VPWR.n666 3.28012
R12379 VPWR.n2130 VPWR.n555 3.28012
R12380 VPWR.n2264 VPWR.n555 3.28012
R12381 VPWR.n2264 VPWR.n474 3.28012
R12382 VPWR.n2326 VPWR.n474 3.28012
R12383 VPWR.n2326 VPWR.n363 3.28012
R12384 VPWR.n2523 VPWR.n90 3.28012
R12385 VPWR.n2463 VPWR.n90 3.28012
R12386 VPWR.n2463 VPWR.n362 3.28012
R12387 VPWR.n2323 VPWR.n362 3.28012
R12388 VPWR.n2323 VPWR.n475 3.28012
R12389 VPWR.n2267 VPWR.n475 3.28012
R12390 VPWR.n2267 VPWR.n554 3.28012
R12391 VPWR.n2127 VPWR.n554 3.28012
R12392 VPWR.n2127 VPWR.n667 3.28012
R12393 VPWR.n2071 VPWR.n667 3.28012
R12394 VPWR.n2071 VPWR.n746 3.28012
R12395 VPWR.n1931 VPWR.n746 3.28012
R12396 VPWR.n1931 VPWR.n859 3.28012
R12397 VPWR.n1875 VPWR.n859 3.28012
R12398 VPWR.n1489 VPWR.n1488 3.28012
R12399 VPWR.n1489 VPWR.n938 3.28012
R12400 VPWR.n1875 VPWR.n938 3.28012
R12401 VPWR.n1503 VPWR.n1501 3.28012
R12402 VPWR.n1503 VPWR.n942 3.28012
R12403 VPWR.n1865 VPWR.n942 3.28012
R12404 VPWR.n1865 VPWR.n855 3.28012
R12405 VPWR.n1941 VPWR.n855 3.28012
R12406 VPWR.n1941 VPWR.n750 3.28012
R12407 VPWR.n2061 VPWR.n750 3.28012
R12408 VPWR.n2061 VPWR.n663 3.28012
R12409 VPWR.n2137 VPWR.n663 3.28012
R12410 VPWR.n2137 VPWR.n558 3.28012
R12411 VPWR.n2257 VPWR.n558 3.28012
R12412 VPWR.n2257 VPWR.n471 3.28012
R12413 VPWR.n2333 VPWR.n471 3.28012
R12414 VPWR.n2333 VPWR.n366 3.28012
R12415 VPWR.n2538 VPWR.n83 3.28012
R12416 VPWR.n2450 VPWR.n83 3.28012
R12417 VPWR.n2450 VPWR.n367 3.28012
R12418 VPWR.n2336 VPWR.n367 3.28012
R12419 VPWR.n2336 VPWR.n470 3.28012
R12420 VPWR.n2254 VPWR.n470 3.28012
R12421 VPWR.n2254 VPWR.n559 3.28012
R12422 VPWR.n2140 VPWR.n559 3.28012
R12423 VPWR.n2140 VPWR.n662 3.28012
R12424 VPWR.n2058 VPWR.n662 3.28012
R12425 VPWR.n2058 VPWR.n751 3.28012
R12426 VPWR.n1944 VPWR.n751 3.28012
R12427 VPWR.n1944 VPWR.n854 3.28012
R12428 VPWR.n1862 VPWR.n854 3.28012
R12429 VPWR.n1512 VPWR.n1511 3.28012
R12430 VPWR.n1511 VPWR.n943 3.28012
R12431 VPWR.n1862 VPWR.n943 3.28012
R12432 VPWR.n1517 VPWR.n1515 3.28012
R12433 VPWR.n1517 VPWR.n946 3.28012
R12434 VPWR.n1855 VPWR.n946 3.28012
R12435 VPWR.n1855 VPWR.n851 3.28012
R12436 VPWR.n1951 VPWR.n851 3.28012
R12437 VPWR.n1951 VPWR.n754 3.28012
R12438 VPWR.n2051 VPWR.n754 3.28012
R12439 VPWR.n2051 VPWR.n659 3.28012
R12440 VPWR.n2147 VPWR.n659 3.28012
R12441 VPWR.n2147 VPWR.n562 3.28012
R12442 VPWR.n2247 VPWR.n562 3.28012
R12443 VPWR.n2247 VPWR.n467 3.28012
R12444 VPWR.n2343 VPWR.n467 3.28012
R12445 VPWR.n2343 VPWR.n370 3.28012
R12446 VPWR.n2443 VPWR.n370 3.28012
R12447 VPWR.n2514 VPWR.n95 3.28012
R12448 VPWR.n2470 VPWR.n95 3.28012
R12449 VPWR.n2470 VPWR.n359 3.28012
R12450 VPWR.n2316 VPWR.n359 3.28012
R12451 VPWR.n2316 VPWR.n478 3.28012
R12452 VPWR.n2274 VPWR.n478 3.28012
R12453 VPWR.n2274 VPWR.n551 3.28012
R12454 VPWR.n2120 VPWR.n551 3.28012
R12455 VPWR.n2120 VPWR.n670 3.28012
R12456 VPWR.n2078 VPWR.n670 3.28012
R12457 VPWR.n2078 VPWR.n743 3.28012
R12458 VPWR.n1924 VPWR.n743 3.28012
R12459 VPWR.n1924 VPWR.n862 3.28012
R12460 VPWR.n1882 VPWR.n862 3.28012
R12461 VPWR.n1882 VPWR.n935 3.28012
R12462 VPWR.n1586 VPWR.n1585 3.28012
R12463 VPWR.n1585 VPWR.n935 3.28012
R12464 VPWR.n1526 VPWR.n1525 3.28012
R12465 VPWR.n1525 VPWR.n947 3.28012
R12466 VPWR.n1852 VPWR.n947 3.28012
R12467 VPWR.n1852 VPWR.n850 3.28012
R12468 VPWR.n1954 VPWR.n850 3.28012
R12469 VPWR.n1954 VPWR.n755 3.28012
R12470 VPWR.n2048 VPWR.n755 3.28012
R12471 VPWR.n2048 VPWR.n658 3.28012
R12472 VPWR.n2150 VPWR.n658 3.28012
R12473 VPWR.n2150 VPWR.n563 3.28012
R12474 VPWR.n2244 VPWR.n563 3.28012
R12475 VPWR.n2244 VPWR.n466 3.28012
R12476 VPWR.n2346 VPWR.n466 3.28012
R12477 VPWR.n2346 VPWR.n371 3.28012
R12478 VPWR.n2440 VPWR.n371 3.28012
R12479 VPWR.n2559 VPWR.n72 3.28012
R12480 VPWR.n2433 VPWR.n72 3.28012
R12481 VPWR.n2433 VPWR.n374 3.28012
R12482 VPWR.n2353 VPWR.n374 3.28012
R12483 VPWR.n2353 VPWR.n463 3.28012
R12484 VPWR.n2237 VPWR.n463 3.28012
R12485 VPWR.n2237 VPWR.n566 3.28012
R12486 VPWR.n2157 VPWR.n566 3.28012
R12487 VPWR.n2157 VPWR.n655 3.28012
R12488 VPWR.n2041 VPWR.n655 3.28012
R12489 VPWR.n2041 VPWR.n758 3.28012
R12490 VPWR.n1961 VPWR.n758 3.28012
R12491 VPWR.n1961 VPWR.n847 3.28012
R12492 VPWR.n1845 VPWR.n847 3.28012
R12493 VPWR.n1845 VPWR.n950 3.28012
R12494 VPWR.n1539 VPWR.n1145 3.28012
R12495 VPWR.n1539 VPWR.n950 3.28012
R12496 VPWR.n1589 VPWR.n1128 3.28012
R12497 VPWR.n1128 VPWR.n934 3.28012
R12498 VPWR.n1885 VPWR.n934 3.28012
R12499 VPWR.n1885 VPWR.n863 3.28012
R12500 VPWR.n1921 VPWR.n863 3.28012
R12501 VPWR.n1921 VPWR.n742 3.28012
R12502 VPWR.n2081 VPWR.n742 3.28012
R12503 VPWR.n2081 VPWR.n671 3.28012
R12504 VPWR.n2117 VPWR.n671 3.28012
R12505 VPWR.n2117 VPWR.n550 3.28012
R12506 VPWR.n2277 VPWR.n550 3.28012
R12507 VPWR.n2277 VPWR.n479 3.28012
R12508 VPWR.n2313 VPWR.n479 3.28012
R12509 VPWR.n2313 VPWR.n358 3.28012
R12510 VPWR.n2473 VPWR.n358 3.28012
R12511 VPWR.n2473 VPWR.n96 3.28012
R12512 VPWR.n2562 VPWR.n71 3.28012
R12513 VPWR.n2430 VPWR.n71 3.28012
R12514 VPWR.n2430 VPWR.n375 3.28012
R12515 VPWR.n2356 VPWR.n375 3.28012
R12516 VPWR.n2356 VPWR.n462 3.28012
R12517 VPWR.n2234 VPWR.n462 3.28012
R12518 VPWR.n2234 VPWR.n567 3.28012
R12519 VPWR.n2160 VPWR.n567 3.28012
R12520 VPWR.n2160 VPWR.n654 3.28012
R12521 VPWR.n2038 VPWR.n654 3.28012
R12522 VPWR.n2038 VPWR.n759 3.28012
R12523 VPWR.n1964 VPWR.n759 3.28012
R12524 VPWR.n1964 VPWR.n846 3.28012
R12525 VPWR.n1842 VPWR.n846 3.28012
R12526 VPWR.n1842 VPWR.n951 3.28012
R12527 VPWR.n1532 VPWR.n951 3.28012
R12528 VPWR.n1532 VPWR.n1531 3.28012
R12529 VPWR.n1764 VPWR.n1045 3.28012
R12530 VPWR.n1764 VPWR.n954 3.28012
R12531 VPWR.n1835 VPWR.n954 3.28012
R12532 VPWR.n1835 VPWR.n843 3.28012
R12533 VPWR.n1971 VPWR.n843 3.28012
R12534 VPWR.n1971 VPWR.n762 3.28012
R12535 VPWR.n2031 VPWR.n762 3.28012
R12536 VPWR.n2031 VPWR.n651 3.28012
R12537 VPWR.n2167 VPWR.n651 3.28012
R12538 VPWR.n2167 VPWR.n570 3.28012
R12539 VPWR.n2227 VPWR.n570 3.28012
R12540 VPWR.n2227 VPWR.n459 3.28012
R12541 VPWR.n2363 VPWR.n459 3.28012
R12542 VPWR.n2363 VPWR.n378 3.28012
R12543 VPWR.n2423 VPWR.n378 3.28012
R12544 VPWR.n2423 VPWR.n66 3.28012
R12545 VPWR.n2583 VPWR.n60 3.28012
R12546 VPWR.n2413 VPWR.n60 3.28012
R12547 VPWR.n2413 VPWR.n382 3.28012
R12548 VPWR.n2373 VPWR.n382 3.28012
R12549 VPWR.n2373 VPWR.n455 3.28012
R12550 VPWR.n2217 VPWR.n455 3.28012
R12551 VPWR.n2217 VPWR.n574 3.28012
R12552 VPWR.n2177 VPWR.n574 3.28012
R12553 VPWR.n2177 VPWR.n647 3.28012
R12554 VPWR.n2021 VPWR.n647 3.28012
R12555 VPWR.n2021 VPWR.n766 3.28012
R12556 VPWR.n1981 VPWR.n766 3.28012
R12557 VPWR.n1981 VPWR.n839 3.28012
R12558 VPWR.n1825 VPWR.n839 3.28012
R12559 VPWR.n1825 VPWR.n958 3.28012
R12560 VPWR.n1752 VPWR.n958 3.28012
R12561 VPWR.n1753 VPWR.n1752 3.28012
R12562 VPWR.n1757 VPWR.n1756 3.28012
R12563 VPWR.n1757 VPWR.n955 3.28012
R12564 VPWR.n1832 VPWR.n955 3.28012
R12565 VPWR.n1832 VPWR.n842 3.28012
R12566 VPWR.n1974 VPWR.n842 3.28012
R12567 VPWR.n1974 VPWR.n763 3.28012
R12568 VPWR.n2028 VPWR.n763 3.28012
R12569 VPWR.n2028 VPWR.n650 3.28012
R12570 VPWR.n2170 VPWR.n650 3.28012
R12571 VPWR.n2170 VPWR.n571 3.28012
R12572 VPWR.n2224 VPWR.n571 3.28012
R12573 VPWR.n2224 VPWR.n458 3.28012
R12574 VPWR.n2366 VPWR.n458 3.28012
R12575 VPWR.n2366 VPWR.n379 3.28012
R12576 VPWR.n2420 VPWR.n379 3.28012
R12577 VPWR.n2420 VPWR.n65 3.28012
R12578 VPWR.n2574 VPWR.n65 3.28012
R12579 VPWR.n2586 VPWR.n59 3.28012
R12580 VPWR.n2410 VPWR.n59 3.28012
R12581 VPWR.n2410 VPWR.n383 3.28012
R12582 VPWR.n2376 VPWR.n383 3.28012
R12583 VPWR.n2376 VPWR.n454 3.28012
R12584 VPWR.n2214 VPWR.n454 3.28012
R12585 VPWR.n2214 VPWR.n575 3.28012
R12586 VPWR.n2180 VPWR.n575 3.28012
R12587 VPWR.n2180 VPWR.n646 3.28012
R12588 VPWR.n2018 VPWR.n646 3.28012
R12589 VPWR.n2018 VPWR.n767 3.28012
R12590 VPWR.n1984 VPWR.n767 3.28012
R12591 VPWR.n1984 VPWR.n838 3.28012
R12592 VPWR.n1822 VPWR.n838 3.28012
R12593 VPWR.n1822 VPWR.n959 3.28012
R12594 VPWR.n1788 VPWR.n959 3.28012
R12595 VPWR.n1788 VPWR.n1037 3.28012
R12596 VPWR.n1465 VPWR.n1232 3.28012
R12597 VPWR.n1465 VPWR.n931 3.28012
R12598 VPWR.n1892 VPWR.n931 3.28012
R12599 VPWR.n1892 VPWR.n929 3.28012
R12600 VPWR.n1914 VPWR.n929 3.28012
R12601 VPWR.n1914 VPWR.n739 3.28012
R12602 VPWR.n2088 VPWR.n739 3.28012
R12603 VPWR.n2088 VPWR.n737 3.28012
R12604 VPWR.n2110 VPWR.n737 3.28012
R12605 VPWR.n2110 VPWR.n547 3.28012
R12606 VPWR.n2284 VPWR.n547 3.28012
R12607 VPWR.n2284 VPWR.n545 3.28012
R12608 VPWR.n2306 VPWR.n545 3.28012
R12609 VPWR.n2306 VPWR.n355 3.28012
R12610 VPWR.n2480 VPWR.n355 3.28012
R12611 VPWR.n2480 VPWR.n353 3.28012
R12612 VPWR.n2502 VPWR.n353 3.28012
R12613 VPWR.n2404 VPWR.n22 3.28012
R12614 VPWR.n2404 VPWR.n449 3.28012
R12615 VPWR.n2382 VPWR.n449 3.28012
R12616 VPWR.n2382 VPWR.n451 3.28012
R12617 VPWR.n2208 VPWR.n451 3.28012
R12618 VPWR.n2208 VPWR.n641 3.28012
R12619 VPWR.n2186 VPWR.n641 3.28012
R12620 VPWR.n2186 VPWR.n643 3.28012
R12621 VPWR.n2012 VPWR.n643 3.28012
R12622 VPWR.n2012 VPWR.n833 3.28012
R12623 VPWR.n1990 VPWR.n833 3.28012
R12624 VPWR.n1990 VPWR.n835 3.28012
R12625 VPWR.n1816 VPWR.n835 3.28012
R12626 VPWR.n1816 VPWR.n1025 3.28012
R12627 VPWR.n1794 VPWR.n1025 3.28012
R12628 VPWR.n1794 VPWR.n1028 3.28012
R12629 VPWR.n2594 VPWR.n22 3.26393
R12630 VPWR.n2863 VPWR 3.18182
R12631 VPWR.n2832 VPWR.n2831 3.1005
R12632 VPWR.n2826 VPWR.n2825 3.1005
R12633 VPWR.n2846 VPWR.n2815 3.1005
R12634 VPWR.n1324 VPWR.n1322 3.01226
R12635 VPWR.n1328 VPWR.n1304 2.63579
R12636 VPWR.n2731 VPWR.n2730 2.25932
R12637 VPWR.n1447 VPWR.n1446 2.06026
R12638 VPWR.n1447 VPWR.n1026 1.78803
R12639 VPWR.n2384 VPWR.n2383 1.32852
R12640 VPWR.n2287 VPWR.n450 1.32852
R12641 VPWR.n2207 VPWR.n2206 1.32852
R12642 VPWR.n2205 VPWR.n2204 1.32852
R12643 VPWR.n2188 VPWR.n2187 1.32852
R12644 VPWR.n2091 VPWR.n642 1.32852
R12645 VPWR.n2011 VPWR.n2010 1.32852
R12646 VPWR.n2009 VPWR.n2008 1.32852
R12647 VPWR.n1992 VPWR.n1991 1.32852
R12648 VPWR.n1895 VPWR.n834 1.32852
R12649 VPWR.n2401 VPWR.n2400 1.32852
R12650 VPWR.n1815 VPWR.n1814 1.32852
R12651 VPWR.n2403 VPWR.n2402 1.32852
R12652 VPWR.n1813 VPWR.n1812 1.32852
R12653 VPWR.n2483 VPWR.n21 1.32852
R12654 VPWR.n1796 VPWR.n1795 1.32852
R12655 VPWR.n2596 VPWR.n2595 1.32852
R12656 VPWR.n1055 VPWR.n1026 1.32852
R12657 VPWR.n2482 VPWR 1.25994
R12658 VPWR VPWR.n354 1.25994
R12659 VPWR VPWR.n2304 1.25994
R12660 VPWR.n2303 VPWR 1.25994
R12661 VPWR.n2286 VPWR 1.25994
R12662 VPWR VPWR.n546 1.25994
R12663 VPWR VPWR.n2108 1.25994
R12664 VPWR.n2107 VPWR 1.25994
R12665 VPWR.n2090 VPWR 1.25994
R12666 VPWR VPWR.n738 1.25994
R12667 VPWR VPWR.n1912 1.25994
R12668 VPWR.n1911 VPWR 1.25994
R12669 VPWR.n1894 VPWR 1.25994
R12670 VPWR VPWR.n930 1.25994
R12671 VPWR.n2499 VPWR 1.25994
R12672 VPWR VPWR.n1450 1.25994
R12673 VPWR VPWR.n2500 1.25994
R12674 VPWR.n1449 VPWR 1.25994
R12675 VPWR.n2597 VPWR.n2596 1.144
R12676 VPWR.n2861 VPWR.n2860 0.936724
R12677 VPWR.n2592 VPWR 0.925943
R12678 VPWR VPWR.n1063 0.925943
R12679 VPWR.n2860 VPWR.n2816 0.925245
R12680 VPWR.n2569 VPWR.n67 0.904391
R12681 VPWR.n2509 VPWR.n97 0.904391
R12682 VPWR.n2552 VPWR.n76 0.904391
R12683 VPWR.n2545 VPWR.n79 0.904391
R12684 VPWR.n2533 VPWR.n85 0.904391
R12685 VPWR.n2528 VPWR.n88 0.904391
R12686 VPWR.n1222 VPWR.n1178 0.904391
R12687 VPWR.n2521 VPWR.n91 0.904391
R12688 VPWR.n1624 VPWR.n1102 0.904391
R12689 VPWR.n1640 VPWR.n1094 0.904391
R12690 VPWR.n2540 VPWR.n82 0.904391
R12691 VPWR.n1651 VPWR.n1092 0.904391
R12692 VPWR.n1211 VPWR.n1210 0.904391
R12693 VPWR.n2516 VPWR.n94 0.904391
R12694 VPWR.n1613 VPWR.n1104 0.904391
R12695 VPWR.n1667 VPWR.n1084 0.904391
R12696 VPWR.n2557 VPWR.n73 0.904391
R12697 VPWR.n1678 VPWR.n1082 0.904391
R12698 VPWR.n1591 VPWR.n1127 0.904391
R12699 VPWR.n2564 VPWR.n70 0.904391
R12700 VPWR.n1197 VPWR.n1196 0.904391
R12701 VPWR.n1694 VPWR.n1074 0.904391
R12702 VPWR.n1742 VPWR.n1057 0.904391
R12703 VPWR.n1705 VPWR.n1071 0.904391
R12704 VPWR.n2581 VPWR.n61 0.904391
R12705 VPWR.n2588 VPWR.n58 0.904391
R12706 VPWR.n1737 VPWR.n1735 0.904391
R12707 VPWR.n1597 VPWR.n1596 0.904391
R12708 VPWR.n2504 VPWR.n289 0.904391
R12709 VPWR.n2576 VPWR.n64 0.904391
R12710 VPWR VPWR.n2863 0.812229
R12711 VPWR.n140 VPWR.n64 0.675548
R12712 VPWR.n152 VPWR.n67 0.675548
R12713 VPWR.n164 VPWR.n70 0.675548
R12714 VPWR.n176 VPWR.n73 0.675548
R12715 VPWR.n188 VPWR.n76 0.675548
R12716 VPWR.n200 VPWR.n79 0.675548
R12717 VPWR.n212 VPWR.n82 0.675548
R12718 VPWR.n224 VPWR.n85 0.675548
R12719 VPWR.n236 VPWR.n88 0.675548
R12720 VPWR.n248 VPWR.n91 0.675548
R12721 VPWR.n260 VPWR.n94 0.675548
R12722 VPWR.n272 VPWR.n97 0.675548
R12723 VPWR.n289 VPWR.n288 0.675548
R12724 VPWR.n128 VPWR.n61 0.675548
R12725 VPWR.n117 VPWR.n58 0.675548
R12726 VPWR.n1735 VPWR.n1734 0.675548
R12727 VPWR.n1719 VPWR.n1057 0.675548
R12728 VPWR.n1707 VPWR.n1705 0.675548
R12729 VPWR.n1696 VPWR.n1694 0.675548
R12730 VPWR.n1196 VPWR.n1195 0.675548
R12731 VPWR.n1680 VPWR.n1678 0.675548
R12732 VPWR.n1669 VPWR.n1667 0.675548
R12733 VPWR.n1210 VPWR.n1209 0.675548
R12734 VPWR.n1653 VPWR.n1651 0.675548
R12735 VPWR.n1642 VPWR.n1640 0.675548
R12736 VPWR.n1178 VPWR.n1177 0.675548
R12737 VPWR.n1626 VPWR.n1624 0.675548
R12738 VPWR.n1615 VPWR.n1613 0.675548
R12739 VPWR.n1127 VPWR.n1126 0.675548
R12740 VPWR.n1599 VPWR.n1597 0.675548
R12741 VPWR.n2806 VPWR.n2805 0.672385
R12742 VPWR.n2790 VPWR.n2785 0.672385
R12743 VPWR.n2770 VPWR.n2765 0.672385
R12744 VPWR.n2751 VPWR.n2746 0.672385
R12745 VPWR.n7 VPWR 0.63497
R12746 VPWR.n1242 VPWR 0.63497
R12747 VPWR.n1265 VPWR 0.63497
R12748 VPWR.n1289 VPWR 0.63497
R12749 VPWR.n24 VPWR 0.499542
R12750 VPWR.n2814 VPWR.n2813 0.442692
R12751 VPWR.n1120 VPWR.n1118 0.404056
R12752 VPWR.n144 VPWR.n138 0.404056
R12753 VPWR.n156 VPWR.n150 0.404056
R12754 VPWR.n168 VPWR.n162 0.404056
R12755 VPWR.n180 VPWR.n174 0.404056
R12756 VPWR.n192 VPWR.n186 0.404056
R12757 VPWR.n204 VPWR.n198 0.404056
R12758 VPWR.n216 VPWR.n210 0.404056
R12759 VPWR.n228 VPWR.n222 0.404056
R12760 VPWR.n240 VPWR.n234 0.404056
R12761 VPWR.n252 VPWR.n246 0.404056
R12762 VPWR.n264 VPWR.n258 0.404056
R12763 VPWR.n276 VPWR.n270 0.404056
R12764 VPWR.n283 VPWR.n101 0.404056
R12765 VPWR.n110 VPWR.n105 0.404056
R12766 VPWR.n132 VPWR.n126 0.404056
R12767 VPWR.n121 VPWR.n115 0.404056
R12768 VPWR.n1729 VPWR.n1065 0.404056
R12769 VPWR.n1723 VPWR.n1717 0.404056
R12770 VPWR.n1711 VPWR.n1070 0.404056
R12771 VPWR.n1704 VPWR.n1702 0.404056
R12772 VPWR.n1693 VPWR.n1691 0.404056
R12773 VPWR.n1684 VPWR.n1081 0.404056
R12774 VPWR.n1677 VPWR.n1675 0.404056
R12775 VPWR.n1666 VPWR.n1664 0.404056
R12776 VPWR.n1657 VPWR.n1091 0.404056
R12777 VPWR.n1650 VPWR.n1648 0.404056
R12778 VPWR.n1639 VPWR.n1637 0.404056
R12779 VPWR.n1630 VPWR.n1101 0.404056
R12780 VPWR.n1623 VPWR.n1621 0.404056
R12781 VPWR.n1612 VPWR.n1610 0.404056
R12782 VPWR.n1603 VPWR.n1111 0.404056
R12783 VPWR.n2860 VPWR.n2859 0.388
R12784 VPWR.n1608 VPWR.n1607 0.349144
R12785 VPWR.n1608 VPWR.n1099 0.349144
R12786 VPWR.n1634 VPWR.n1099 0.349144
R12787 VPWR.n1635 VPWR.n1634 0.349144
R12788 VPWR.n1635 VPWR.n1089 0.349144
R12789 VPWR.n1661 VPWR.n1089 0.349144
R12790 VPWR.n1662 VPWR.n1661 0.349144
R12791 VPWR.n1662 VPWR.n1079 0.349144
R12792 VPWR.n1688 VPWR.n1079 0.349144
R12793 VPWR.n1689 VPWR.n1688 0.349144
R12794 VPWR.n1689 VPWR.n1068 0.349144
R12795 VPWR.n1715 VPWR.n1068 0.349144
R12796 VPWR.n1727 VPWR.n1715 0.349144
R12797 VPWR.n281 VPWR.n280 0.349144
R12798 VPWR.n280 VPWR.n268 0.349144
R12799 VPWR.n268 VPWR.n256 0.349144
R12800 VPWR.n256 VPWR.n244 0.349144
R12801 VPWR.n244 VPWR.n232 0.349144
R12802 VPWR.n232 VPWR.n220 0.349144
R12803 VPWR.n220 VPWR.n208 0.349144
R12804 VPWR.n208 VPWR.n196 0.349144
R12805 VPWR.n196 VPWR.n184 0.349144
R12806 VPWR.n184 VPWR.n172 0.349144
R12807 VPWR.n172 VPWR.n160 0.349144
R12808 VPWR.n160 VPWR.n148 0.349144
R12809 VPWR.n148 VPWR.n136 0.349144
R12810 VPWR.n1462 VPWR.n1456 0.346131
R12811 VPWR.n1461 VPWR.n1457 0.346131
R12812 VPWR.n1582 VPWR.n1136 0.346131
R12813 VPWR.n1581 VPWR.n1577 0.346131
R12814 VPWR.n1576 VPWR.n1572 0.346131
R12815 VPWR.n1571 VPWR.n1567 0.346131
R12816 VPWR.n1566 VPWR.n1562 0.346131
R12817 VPWR.n1561 VPWR.n1557 0.346131
R12818 VPWR.n1556 VPWR.n1552 0.346131
R12819 VPWR.n1551 VPWR.n1547 0.346131
R12820 VPWR.n1546 VPWR.n1542 0.346131
R12821 VPWR.n1767 VPWR.n1042 0.346131
R12822 VPWR.n1784 VPWR.n1780 0.346131
R12823 VPWR.n1785 VPWR.n1776 0.346131
R12824 VPWR.n1772 VPWR.n1771 0.346131
R12825 VPWR.n2862 VPWR.n2861 0.304571
R12826 VPWR.n2594 VPWR.n55 0.300179
R12827 VPWR.n1118 VPWR.n1113 0.286958
R12828 VPWR.n145 VPWR.n144 0.286958
R12829 VPWR.n157 VPWR.n156 0.286958
R12830 VPWR.n169 VPWR.n168 0.286958
R12831 VPWR.n181 VPWR.n180 0.286958
R12832 VPWR.n193 VPWR.n192 0.286958
R12833 VPWR.n205 VPWR.n204 0.286958
R12834 VPWR.n217 VPWR.n216 0.286958
R12835 VPWR.n229 VPWR.n228 0.286958
R12836 VPWR.n241 VPWR.n240 0.286958
R12837 VPWR.n253 VPWR.n252 0.286958
R12838 VPWR.n265 VPWR.n264 0.286958
R12839 VPWR.n277 VPWR.n276 0.286958
R12840 VPWR.n283 VPWR.n102 0.286958
R12841 VPWR.n111 VPWR.n110 0.286958
R12842 VPWR.n133 VPWR.n132 0.286958
R12843 VPWR.n122 VPWR.n121 0.286958
R12844 VPWR.n1729 VPWR.n1066 0.286958
R12845 VPWR.n1724 VPWR.n1723 0.286958
R12846 VPWR.n1712 VPWR.n1711 0.286958
R12847 VPWR.n1702 VPWR.n1072 0.286958
R12848 VPWR.n1691 VPWR.n1075 0.286958
R12849 VPWR.n1685 VPWR.n1684 0.286958
R12850 VPWR.n1675 VPWR.n1083 0.286958
R12851 VPWR.n1664 VPWR.n1085 0.286958
R12852 VPWR.n1658 VPWR.n1657 0.286958
R12853 VPWR.n1648 VPWR.n1093 0.286958
R12854 VPWR.n1637 VPWR.n1095 0.286958
R12855 VPWR.n1631 VPWR.n1630 0.286958
R12856 VPWR.n1621 VPWR.n1103 0.286958
R12857 VPWR.n1610 VPWR.n1105 0.286958
R12858 VPWR.n1604 VPWR.n1603 0.286958
R12859 VPWR.n55 VPWR 0.2505
R12860 VPWR VPWR.n2481 0.249238
R12861 VPWR.n2472 VPWR 0.249238
R12862 VPWR VPWR.n2471 0.249238
R12863 VPWR.n2385 VPWR 0.249238
R12864 VPWR.n2386 VPWR 0.249238
R12865 VPWR.n2387 VPWR 0.249238
R12866 VPWR.n2388 VPWR 0.249238
R12867 VPWR.n2305 VPWR 0.249238
R12868 VPWR.n2314 VPWR 0.249238
R12869 VPWR.n2315 VPWR 0.249238
R12870 VPWR.n2324 VPWR 0.249238
R12871 VPWR.n2325 VPWR 0.249238
R12872 VPWR.n2383 VPWR 0.249238
R12873 VPWR.n2375 VPWR 0.249238
R12874 VPWR.n2374 VPWR 0.249238
R12875 VPWR.n2365 VPWR 0.249238
R12876 VPWR.n2364 VPWR 0.249238
R12877 VPWR.n2355 VPWR 0.249238
R12878 VPWR.n2354 VPWR 0.249238
R12879 VPWR.n2345 VPWR 0.249238
R12880 VPWR.n2344 VPWR 0.249238
R12881 VPWR.n2335 VPWR 0.249238
R12882 VPWR.n2334 VPWR 0.249238
R12883 VPWR VPWR.n2302 0.249238
R12884 VPWR VPWR.n2301 0.249238
R12885 VPWR VPWR.n2300 0.249238
R12886 VPWR VPWR.n2299 0.249238
R12887 VPWR VPWR.n2298 0.249238
R12888 VPWR VPWR.n2287 0.249238
R12889 VPWR VPWR.n2288 0.249238
R12890 VPWR VPWR.n2289 0.249238
R12891 VPWR VPWR.n2290 0.249238
R12892 VPWR VPWR.n2291 0.249238
R12893 VPWR VPWR.n2292 0.249238
R12894 VPWR VPWR.n2293 0.249238
R12895 VPWR VPWR.n2294 0.249238
R12896 VPWR VPWR.n2295 0.249238
R12897 VPWR VPWR.n2296 0.249238
R12898 VPWR VPWR.n2297 0.249238
R12899 VPWR VPWR.n2285 0.249238
R12900 VPWR.n2276 VPWR 0.249238
R12901 VPWR VPWR.n2275 0.249238
R12902 VPWR.n2266 VPWR 0.249238
R12903 VPWR VPWR.n2265 0.249238
R12904 VPWR.n2207 VPWR 0.249238
R12905 VPWR VPWR.n2215 0.249238
R12906 VPWR.n2216 VPWR 0.249238
R12907 VPWR VPWR.n2225 0.249238
R12908 VPWR.n2226 VPWR 0.249238
R12909 VPWR VPWR.n2235 0.249238
R12910 VPWR.n2236 VPWR 0.249238
R12911 VPWR VPWR.n2245 0.249238
R12912 VPWR.n2246 VPWR 0.249238
R12913 VPWR VPWR.n2255 0.249238
R12914 VPWR.n2256 VPWR 0.249238
R12915 VPWR.n2189 VPWR 0.249238
R12916 VPWR.n2190 VPWR 0.249238
R12917 VPWR.n2191 VPWR 0.249238
R12918 VPWR.n2192 VPWR 0.249238
R12919 VPWR.n2193 VPWR 0.249238
R12920 VPWR.n2204 VPWR 0.249238
R12921 VPWR.n2203 VPWR 0.249238
R12922 VPWR.n2202 VPWR 0.249238
R12923 VPWR.n2201 VPWR 0.249238
R12924 VPWR.n2200 VPWR 0.249238
R12925 VPWR.n2199 VPWR 0.249238
R12926 VPWR.n2198 VPWR 0.249238
R12927 VPWR.n2197 VPWR 0.249238
R12928 VPWR.n2196 VPWR 0.249238
R12929 VPWR.n2195 VPWR 0.249238
R12930 VPWR.n2194 VPWR 0.249238
R12931 VPWR.n2109 VPWR 0.249238
R12932 VPWR.n2118 VPWR 0.249238
R12933 VPWR.n2119 VPWR 0.249238
R12934 VPWR.n2128 VPWR 0.249238
R12935 VPWR.n2129 VPWR 0.249238
R12936 VPWR.n2187 VPWR 0.249238
R12937 VPWR.n2179 VPWR 0.249238
R12938 VPWR.n2178 VPWR 0.249238
R12939 VPWR.n2169 VPWR 0.249238
R12940 VPWR.n2168 VPWR 0.249238
R12941 VPWR.n2159 VPWR 0.249238
R12942 VPWR.n2158 VPWR 0.249238
R12943 VPWR.n2149 VPWR 0.249238
R12944 VPWR.n2148 VPWR 0.249238
R12945 VPWR.n2139 VPWR 0.249238
R12946 VPWR.n2138 VPWR 0.249238
R12947 VPWR VPWR.n2106 0.249238
R12948 VPWR VPWR.n2105 0.249238
R12949 VPWR VPWR.n2104 0.249238
R12950 VPWR VPWR.n2103 0.249238
R12951 VPWR VPWR.n2102 0.249238
R12952 VPWR VPWR.n2091 0.249238
R12953 VPWR VPWR.n2092 0.249238
R12954 VPWR VPWR.n2093 0.249238
R12955 VPWR VPWR.n2094 0.249238
R12956 VPWR VPWR.n2095 0.249238
R12957 VPWR VPWR.n2096 0.249238
R12958 VPWR VPWR.n2097 0.249238
R12959 VPWR VPWR.n2098 0.249238
R12960 VPWR VPWR.n2099 0.249238
R12961 VPWR VPWR.n2100 0.249238
R12962 VPWR VPWR.n2101 0.249238
R12963 VPWR VPWR.n2089 0.249238
R12964 VPWR.n2080 VPWR 0.249238
R12965 VPWR VPWR.n2079 0.249238
R12966 VPWR.n2070 VPWR 0.249238
R12967 VPWR VPWR.n2069 0.249238
R12968 VPWR.n2011 VPWR 0.249238
R12969 VPWR VPWR.n2019 0.249238
R12970 VPWR.n2020 VPWR 0.249238
R12971 VPWR VPWR.n2029 0.249238
R12972 VPWR.n2030 VPWR 0.249238
R12973 VPWR VPWR.n2039 0.249238
R12974 VPWR.n2040 VPWR 0.249238
R12975 VPWR VPWR.n2049 0.249238
R12976 VPWR.n2050 VPWR 0.249238
R12977 VPWR VPWR.n2059 0.249238
R12978 VPWR.n2060 VPWR 0.249238
R12979 VPWR.n1993 VPWR 0.249238
R12980 VPWR.n1994 VPWR 0.249238
R12981 VPWR.n1995 VPWR 0.249238
R12982 VPWR.n1996 VPWR 0.249238
R12983 VPWR.n1997 VPWR 0.249238
R12984 VPWR.n2008 VPWR 0.249238
R12985 VPWR.n2007 VPWR 0.249238
R12986 VPWR.n2006 VPWR 0.249238
R12987 VPWR.n2005 VPWR 0.249238
R12988 VPWR.n2004 VPWR 0.249238
R12989 VPWR.n2003 VPWR 0.249238
R12990 VPWR.n2002 VPWR 0.249238
R12991 VPWR.n2001 VPWR 0.249238
R12992 VPWR.n2000 VPWR 0.249238
R12993 VPWR.n1999 VPWR 0.249238
R12994 VPWR.n1998 VPWR 0.249238
R12995 VPWR.n1913 VPWR 0.249238
R12996 VPWR.n1922 VPWR 0.249238
R12997 VPWR.n1923 VPWR 0.249238
R12998 VPWR.n1932 VPWR 0.249238
R12999 VPWR.n1933 VPWR 0.249238
R13000 VPWR.n1991 VPWR 0.249238
R13001 VPWR.n1983 VPWR 0.249238
R13002 VPWR.n1982 VPWR 0.249238
R13003 VPWR.n1973 VPWR 0.249238
R13004 VPWR.n1972 VPWR 0.249238
R13005 VPWR.n1963 VPWR 0.249238
R13006 VPWR.n1962 VPWR 0.249238
R13007 VPWR.n1953 VPWR 0.249238
R13008 VPWR.n1952 VPWR 0.249238
R13009 VPWR.n1943 VPWR 0.249238
R13010 VPWR.n1942 VPWR 0.249238
R13011 VPWR VPWR.n1910 0.249238
R13012 VPWR VPWR.n1909 0.249238
R13013 VPWR VPWR.n1908 0.249238
R13014 VPWR VPWR.n1907 0.249238
R13015 VPWR VPWR.n1906 0.249238
R13016 VPWR VPWR.n1895 0.249238
R13017 VPWR VPWR.n1896 0.249238
R13018 VPWR VPWR.n1897 0.249238
R13019 VPWR VPWR.n1898 0.249238
R13020 VPWR VPWR.n1899 0.249238
R13021 VPWR VPWR.n1900 0.249238
R13022 VPWR VPWR.n1901 0.249238
R13023 VPWR VPWR.n1902 0.249238
R13024 VPWR VPWR.n1903 0.249238
R13025 VPWR VPWR.n1904 0.249238
R13026 VPWR VPWR.n1905 0.249238
R13027 VPWR.n2400 VPWR 0.249238
R13028 VPWR.n2399 VPWR 0.249238
R13029 VPWR.n2398 VPWR 0.249238
R13030 VPWR.n2397 VPWR 0.249238
R13031 VPWR.n2396 VPWR 0.249238
R13032 VPWR.n2395 VPWR 0.249238
R13033 VPWR.n2394 VPWR 0.249238
R13034 VPWR.n2393 VPWR 0.249238
R13035 VPWR.n2392 VPWR 0.249238
R13036 VPWR.n2391 VPWR 0.249238
R13037 VPWR.n2390 VPWR 0.249238
R13038 VPWR.n2389 VPWR 0.249238
R13039 VPWR VPWR.n1893 0.249238
R13040 VPWR.n1884 VPWR 0.249238
R13041 VPWR VPWR.n1883 0.249238
R13042 VPWR.n1874 VPWR 0.249238
R13043 VPWR VPWR.n1873 0.249238
R13044 VPWR.n1864 VPWR 0.249238
R13045 VPWR.n1815 VPWR 0.249238
R13046 VPWR VPWR.n1823 0.249238
R13047 VPWR.n1824 VPWR 0.249238
R13048 VPWR VPWR.n1833 0.249238
R13049 VPWR.n1834 VPWR 0.249238
R13050 VPWR VPWR.n1843 0.249238
R13051 VPWR.n1844 VPWR 0.249238
R13052 VPWR VPWR.n1853 0.249238
R13053 VPWR.n1854 VPWR 0.249238
R13054 VPWR VPWR.n1863 0.249238
R13055 VPWR.n2403 VPWR 0.249238
R13056 VPWR VPWR.n2411 0.249238
R13057 VPWR.n2412 VPWR 0.249238
R13058 VPWR VPWR.n2421 0.249238
R13059 VPWR.n2422 VPWR 0.249238
R13060 VPWR VPWR.n2431 0.249238
R13061 VPWR.n2432 VPWR 0.249238
R13062 VPWR VPWR.n2441 0.249238
R13063 VPWR.n2442 VPWR 0.249238
R13064 VPWR VPWR.n2451 0.249238
R13065 VPWR.n2452 VPWR 0.249238
R13066 VPWR VPWR.n2461 0.249238
R13067 VPWR.n2462 VPWR 0.249238
R13068 VPWR.n1797 VPWR 0.249238
R13069 VPWR.n1798 VPWR 0.249238
R13070 VPWR.n1799 VPWR 0.249238
R13071 VPWR.n1800 VPWR 0.249238
R13072 VPWR.n1801 VPWR 0.249238
R13073 VPWR.n1802 VPWR 0.249238
R13074 VPWR.n1803 VPWR 0.249238
R13075 VPWR.n1804 VPWR 0.249238
R13076 VPWR.n1805 VPWR 0.249238
R13077 VPWR.n1812 VPWR 0.249238
R13078 VPWR.n1811 VPWR 0.249238
R13079 VPWR.n1810 VPWR 0.249238
R13080 VPWR.n1809 VPWR 0.249238
R13081 VPWR.n1808 VPWR 0.249238
R13082 VPWR.n1807 VPWR 0.249238
R13083 VPWR.n1806 VPWR 0.249238
R13084 VPWR VPWR.n2498 0.249238
R13085 VPWR VPWR.n2497 0.249238
R13086 VPWR VPWR.n2496 0.249238
R13087 VPWR VPWR.n2495 0.249238
R13088 VPWR VPWR.n2494 0.249238
R13089 VPWR VPWR.n2493 0.249238
R13090 VPWR VPWR.n2492 0.249238
R13091 VPWR VPWR.n2491 0.249238
R13092 VPWR VPWR.n2490 0.249238
R13093 VPWR VPWR.n2489 0.249238
R13094 VPWR VPWR.n2488 0.249238
R13095 VPWR VPWR.n2483 0.249238
R13096 VPWR VPWR.n2484 0.249238
R13097 VPWR VPWR.n2485 0.249238
R13098 VPWR VPWR.n2486 0.249238
R13099 VPWR VPWR.n2487 0.249238
R13100 VPWR.n2501 VPWR 0.249238
R13101 VPWR.n2512 VPWR 0.249238
R13102 VPWR.n2513 VPWR 0.249238
R13103 VPWR.n2524 VPWR 0.249238
R13104 VPWR.n2525 VPWR 0.249238
R13105 VPWR.n2536 VPWR 0.249238
R13106 VPWR.n2537 VPWR 0.249238
R13107 VPWR.n2548 VPWR 0.249238
R13108 VPWR.n2549 VPWR 0.249238
R13109 VPWR.n2560 VPWR 0.249238
R13110 VPWR.n2561 VPWR 0.249238
R13111 VPWR.n2572 VPWR 0.249238
R13112 VPWR.n2573 VPWR 0.249238
R13113 VPWR.n2584 VPWR 0.249238
R13114 VPWR.n2585 VPWR 0.249238
R13115 VPWR.n2595 VPWR 0.249238
R13116 VPWR VPWR.n1055 0.249238
R13117 VPWR VPWR.n1056 0.249238
R13118 VPWR VPWR.n1754 0.249238
R13119 VPWR.n1755 VPWR 0.249238
R13120 VPWR VPWR.n1529 0.249238
R13121 VPWR.n1530 VPWR 0.249238
R13122 VPWR.n1528 VPWR 0.249238
R13123 VPWR.n1527 VPWR 0.249238
R13124 VPWR.n1514 VPWR 0.249238
R13125 VPWR.n1513 VPWR 0.249238
R13126 VPWR.n1500 VPWR 0.249238
R13127 VPWR.n1499 VPWR 0.249238
R13128 VPWR.n1487 VPWR 0.249238
R13129 VPWR VPWR.n1587 0.249238
R13130 VPWR.n1588 VPWR 0.249238
R13131 VPWR VPWR.n1448 0.249238
R13132 VPWR.n2861 VPWR.n2815 0.245065
R13133 VPWR.n2813 VPWR.n2797 0.213567
R13134 VPWR.n2797 VPWR.n2778 0.213567
R13135 VPWR.n2778 VPWR.n2758 0.213567
R13136 VPWR.n2758 VPWR.n2739 0.213567
R13137 VPWR.n2739 VPWR.n2703 0.213567
R13138 VPWR.n2703 VPWR.n2665 0.213567
R13139 VPWR.n2665 VPWR.n2628 0.213567
R13140 VPWR.n1446 VPWR.n1414 0.213567
R13141 VPWR.n1414 VPWR.n1376 0.213567
R13142 VPWR.n1376 VPWR.n1337 0.213567
R13143 VPWR.n1337 VPWR.n1302 0.213567
R13144 VPWR.n1302 VPWR.n1279 0.213567
R13145 VPWR.n1279 VPWR.n1255 0.213567
R13146 VPWR.n1255 VPWR.n19 0.213567
R13147 VPWR VPWR.n2862 0.204304
R13148 VPWR.n1449 VPWR.n1447 0.179202
R13149 VPWR.n1450 VPWR.n1449 0.154425
R13150 VPWR.n1450 VPWR.n930 0.154425
R13151 VPWR.n1894 VPWR.n930 0.154425
R13152 VPWR.n1911 VPWR.n1894 0.154425
R13153 VPWR.n1912 VPWR.n1911 0.154425
R13154 VPWR.n1912 VPWR.n738 0.154425
R13155 VPWR.n2090 VPWR.n738 0.154425
R13156 VPWR.n2107 VPWR.n2090 0.154425
R13157 VPWR.n2108 VPWR.n2107 0.154425
R13158 VPWR.n2108 VPWR.n546 0.154425
R13159 VPWR.n2286 VPWR.n546 0.154425
R13160 VPWR.n2303 VPWR.n2286 0.154425
R13161 VPWR.n2304 VPWR.n2303 0.154425
R13162 VPWR.n2304 VPWR.n354 0.154425
R13163 VPWR.n2482 VPWR.n354 0.154425
R13164 VPWR.n2499 VPWR.n2482 0.154425
R13165 VPWR.n2500 VPWR.n2499 0.154425
R13166 VPWR.n1796 VPWR.n1026 0.154425
R13167 VPWR.n1813 VPWR.n1796 0.154425
R13168 VPWR.n1814 VPWR.n1813 0.154425
R13169 VPWR.n1814 VPWR.n834 0.154425
R13170 VPWR.n1992 VPWR.n834 0.154425
R13171 VPWR.n2009 VPWR.n1992 0.154425
R13172 VPWR.n2010 VPWR.n2009 0.154425
R13173 VPWR.n2010 VPWR.n642 0.154425
R13174 VPWR.n2188 VPWR.n642 0.154425
R13175 VPWR.n2205 VPWR.n2188 0.154425
R13176 VPWR.n2206 VPWR.n2205 0.154425
R13177 VPWR.n2206 VPWR.n450 0.154425
R13178 VPWR.n2384 VPWR.n450 0.154425
R13179 VPWR.n2401 VPWR.n2384 0.154425
R13180 VPWR.n2402 VPWR.n2401 0.154425
R13181 VPWR.n2402 VPWR.n21 0.154425
R13182 VPWR.n2596 VPWR.n21 0.154425
R13183 VPWR.n8 VPWR.n7 0.147771
R13184 VPWR.n1243 VPWR.n1242 0.147771
R13185 VPWR.n1266 VPWR.n1265 0.147771
R13186 VPWR.n1290 VPWR.n1289 0.147771
R13187 VPWR.n1113 VPWR 0.135917
R13188 VPWR.n145 VPWR 0.135917
R13189 VPWR.n157 VPWR 0.135917
R13190 VPWR.n169 VPWR 0.135917
R13191 VPWR.n181 VPWR 0.135917
R13192 VPWR.n193 VPWR 0.135917
R13193 VPWR.n205 VPWR 0.135917
R13194 VPWR.n217 VPWR 0.135917
R13195 VPWR.n229 VPWR 0.135917
R13196 VPWR.n241 VPWR 0.135917
R13197 VPWR.n253 VPWR 0.135917
R13198 VPWR.n265 VPWR 0.135917
R13199 VPWR.n277 VPWR 0.135917
R13200 VPWR.n102 VPWR 0.135917
R13201 VPWR.n111 VPWR 0.135917
R13202 VPWR.n133 VPWR 0.135917
R13203 VPWR.n122 VPWR 0.135917
R13204 VPWR.n1066 VPWR 0.135917
R13205 VPWR.n1724 VPWR 0.135917
R13206 VPWR.n1712 VPWR 0.135917
R13207 VPWR.n1072 VPWR 0.135917
R13208 VPWR.n1075 VPWR 0.135917
R13209 VPWR.n1685 VPWR 0.135917
R13210 VPWR.n1083 VPWR 0.135917
R13211 VPWR.n1085 VPWR 0.135917
R13212 VPWR.n1658 VPWR 0.135917
R13213 VPWR.n1093 VPWR 0.135917
R13214 VPWR.n1095 VPWR 0.135917
R13215 VPWR.n1631 VPWR 0.135917
R13216 VPWR.n1103 VPWR 0.135917
R13217 VPWR.n1105 VPWR 0.135917
R13218 VPWR.n1604 VPWR 0.135917
R13219 VPWR.n2863 VPWR.n2814 0.127988
R13220 VPWR.n2825 VPWR.n2816 0.1255
R13221 VPWR.n2831 VPWR.n2816 0.1255
R13222 VPWR.n18 VPWR.n0 0.120292
R13223 VPWR.n14 VPWR.n0 0.120292
R13224 VPWR.n9 VPWR.n8 0.120292
R13225 VPWR.n1254 VPWR.n1233 0.120292
R13226 VPWR.n1250 VPWR.n1233 0.120292
R13227 VPWR.n1244 VPWR.n1243 0.120292
R13228 VPWR.n1278 VPWR.n1256 0.120292
R13229 VPWR.n1273 VPWR.n1256 0.120292
R13230 VPWR.n1267 VPWR.n1266 0.120292
R13231 VPWR.n1301 VPWR.n1280 0.120292
R13232 VPWR.n1297 VPWR.n1280 0.120292
R13233 VPWR.n1291 VPWR.n1290 0.120292
R13234 VPWR.n1333 VPWR.n1332 0.120292
R13235 VPWR.n1326 VPWR.n1305 0.120292
R13236 VPWR.n1319 VPWR.n1305 0.120292
R13237 VPWR.n1319 VPWR.n1318 0.120292
R13238 VPWR.n1317 VPWR.n1309 0.120292
R13239 VPWR.n1312 VPWR.n1309 0.120292
R13240 VPWR.n1312 VPWR.n1311 0.120292
R13241 VPWR.n1371 VPWR.n1370 0.120292
R13242 VPWR.n1364 VPWR.n1363 0.120292
R13243 VPWR.n1363 VPWR.n1340 0.120292
R13244 VPWR.n1356 VPWR.n1340 0.120292
R13245 VPWR.n1356 VPWR.n1355 0.120292
R13246 VPWR.n1355 VPWR.n1354 0.120292
R13247 VPWR.n1354 VPWR.n1342 0.120292
R13248 VPWR.n1348 VPWR.n1342 0.120292
R13249 VPWR.n1348 VPWR.n1347 0.120292
R13250 VPWR.n1410 VPWR.n1409 0.120292
R13251 VPWR.n1403 VPWR.n1402 0.120292
R13252 VPWR.n1402 VPWR.n1379 0.120292
R13253 VPWR.n1395 VPWR.n1379 0.120292
R13254 VPWR.n1395 VPWR.n1394 0.120292
R13255 VPWR.n1394 VPWR.n1393 0.120292
R13256 VPWR.n1393 VPWR.n1381 0.120292
R13257 VPWR.n1387 VPWR.n1381 0.120292
R13258 VPWR.n1387 VPWR.n1386 0.120292
R13259 VPWR.n1440 VPWR.n1439 0.120292
R13260 VPWR.n1439 VPWR.n1416 0.120292
R13261 VPWR.n1432 VPWR.n1416 0.120292
R13262 VPWR.n1432 VPWR.n1431 0.120292
R13263 VPWR.n1431 VPWR.n1430 0.120292
R13264 VPWR.n1430 VPWR.n1418 0.120292
R13265 VPWR.n1424 VPWR.n1418 0.120292
R13266 VPWR.n1424 VPWR.n1423 0.120292
R13267 VPWR.n2812 VPWR.n2798 0.120292
R13268 VPWR.n2796 VPWR.n2779 0.120292
R13269 VPWR.n2777 VPWR.n2759 0.120292
R13270 VPWR.n2757 VPWR.n2740 0.120292
R13271 VPWR.n2719 VPWR.n2718 0.120292
R13272 VPWR.n2720 VPWR.n2719 0.120292
R13273 VPWR.n2720 VPWR.n2711 0.120292
R13274 VPWR.n2725 VPWR.n2711 0.120292
R13275 VPWR.n2726 VPWR.n2725 0.120292
R13276 VPWR.n2726 VPWR.n2707 0.120292
R13277 VPWR.n2732 VPWR.n2707 0.120292
R13278 VPWR.n2734 VPWR.n2704 0.120292
R13279 VPWR.n2738 VPWR.n2704 0.120292
R13280 VPWR.n2683 VPWR.n2682 0.120292
R13281 VPWR.n2684 VPWR.n2683 0.120292
R13282 VPWR.n2684 VPWR.n2673 0.120292
R13283 VPWR.n2689 VPWR.n2673 0.120292
R13284 VPWR.n2690 VPWR.n2689 0.120292
R13285 VPWR.n2690 VPWR.n2669 0.120292
R13286 VPWR.n2695 VPWR.n2669 0.120292
R13287 VPWR.n2697 VPWR.n2666 0.120292
R13288 VPWR.n2702 VPWR.n2666 0.120292
R13289 VPWR.n2646 VPWR.n2645 0.120292
R13290 VPWR.n2647 VPWR.n2646 0.120292
R13291 VPWR.n2647 VPWR.n2636 0.120292
R13292 VPWR.n2652 VPWR.n2636 0.120292
R13293 VPWR.n2653 VPWR.n2652 0.120292
R13294 VPWR.n2653 VPWR.n2632 0.120292
R13295 VPWR.n2658 VPWR.n2632 0.120292
R13296 VPWR.n2660 VPWR.n2629 0.120292
R13297 VPWR.n2664 VPWR.n2629 0.120292
R13298 VPWR.n2608 VPWR.n2604 0.120292
R13299 VPWR.n2616 VPWR.n2604 0.120292
R13300 VPWR.n2617 VPWR.n2616 0.120292
R13301 VPWR.n2618 VPWR.n2617 0.120292
R13302 VPWR.n2618 VPWR.n2600 0.120292
R13303 VPWR.n2623 VPWR.n2600 0.120292
R13304 VPWR.n2624 VPWR.n2623 0.120292
R13305 VPWR.n1605 VPWR 0.118556
R13306 VPWR.n1108 VPWR 0.118556
R13307 VPWR.n1619 VPWR 0.118556
R13308 VPWR.n1632 VPWR 0.118556
R13309 VPWR.n1098 VPWR 0.118556
R13310 VPWR.n1646 VPWR 0.118556
R13311 VPWR.n1659 VPWR 0.118556
R13312 VPWR.n1088 VPWR 0.118556
R13313 VPWR.n1673 VPWR 0.118556
R13314 VPWR.n1686 VPWR 0.118556
R13315 VPWR.n1078 VPWR 0.118556
R13316 VPWR.n1700 VPWR 0.118556
R13317 VPWR.n1713 VPWR 0.118556
R13318 VPWR.n1725 VPWR 0.118556
R13319 VPWR VPWR.n1112 0.118556
R13320 VPWR.n1067 VPWR 0.118556
R13321 VPWR.n123 VPWR 0.118556
R13322 VPWR.n112 VPWR 0.118556
R13323 VPWR.n103 VPWR 0.118556
R13324 VPWR.n278 VPWR 0.118556
R13325 VPWR.n266 VPWR 0.118556
R13326 VPWR.n254 VPWR 0.118556
R13327 VPWR.n242 VPWR 0.118556
R13328 VPWR.n230 VPWR 0.118556
R13329 VPWR.n218 VPWR 0.118556
R13330 VPWR.n206 VPWR 0.118556
R13331 VPWR.n194 VPWR 0.118556
R13332 VPWR.n182 VPWR 0.118556
R13333 VPWR.n170 VPWR 0.118556
R13334 VPWR.n158 VPWR 0.118556
R13335 VPWR.n146 VPWR 0.118556
R13336 VPWR.n134 VPWR 0.118556
R13337 VPWR.n1765 VPWR.n1044 0.108238
R13338 VPWR.n1541 VPWR.n1143 0.108238
R13339 VPWR.n1540 VPWR.n1142 0.108238
R13340 VPWR.n1524 VPWR.n1141 0.108238
R13341 VPWR.n1516 VPWR.n1140 0.108238
R13342 VPWR.n1510 VPWR.n1139 0.108238
R13343 VPWR.n1502 VPWR.n1138 0.108238
R13344 VPWR.n1496 VPWR.n1137 0.108238
R13345 VPWR.n1583 VPWR.n1132 0.108238
R13346 VPWR.n1584 VPWR.n1131 0.108238
R13347 VPWR.n1463 VPWR.n1452 0.108238
R13348 VPWR.n1464 VPWR.n1451 0.108238
R13349 VPWR.n1795 VPWR.n1027 0.108238
R13350 VPWR.n1766 VPWR.n1043 0.108238
R13351 VPWR.n1744 VPWR.n1038 0.108238
R13352 VPWR.n1787 VPWR.n1786 0.108238
R13353 VPWR.n2481 VPWR 0.100405
R13354 VPWR.n2472 VPWR 0.100405
R13355 VPWR VPWR.n2385 0.100405
R13356 VPWR VPWR.n2386 0.100405
R13357 VPWR VPWR.n2387 0.100405
R13358 VPWR.n2305 VPWR 0.100405
R13359 VPWR VPWR.n2314 0.100405
R13360 VPWR.n2315 VPWR 0.100405
R13361 VPWR VPWR.n2324 0.100405
R13362 VPWR.n2375 VPWR 0.100405
R13363 VPWR VPWR.n2374 0.100405
R13364 VPWR.n2365 VPWR 0.100405
R13365 VPWR VPWR.n2364 0.100405
R13366 VPWR.n2355 VPWR 0.100405
R13367 VPWR VPWR.n2354 0.100405
R13368 VPWR.n2345 VPWR 0.100405
R13369 VPWR VPWR.n2344 0.100405
R13370 VPWR.n2335 VPWR 0.100405
R13371 VPWR VPWR.n2334 0.100405
R13372 VPWR.n2325 VPWR 0.100405
R13373 VPWR.n2302 VPWR 0.100405
R13374 VPWR.n2301 VPWR 0.100405
R13375 VPWR.n2300 VPWR 0.100405
R13376 VPWR.n2299 VPWR 0.100405
R13377 VPWR.n2288 VPWR 0.100405
R13378 VPWR.n2289 VPWR 0.100405
R13379 VPWR.n2290 VPWR 0.100405
R13380 VPWR.n2291 VPWR 0.100405
R13381 VPWR.n2292 VPWR 0.100405
R13382 VPWR.n2293 VPWR 0.100405
R13383 VPWR.n2294 VPWR 0.100405
R13384 VPWR.n2295 VPWR 0.100405
R13385 VPWR.n2296 VPWR 0.100405
R13386 VPWR.n2297 VPWR 0.100405
R13387 VPWR.n2298 VPWR 0.100405
R13388 VPWR.n2285 VPWR 0.100405
R13389 VPWR.n2276 VPWR 0.100405
R13390 VPWR.n2275 VPWR 0.100405
R13391 VPWR.n2266 VPWR 0.100405
R13392 VPWR.n2215 VPWR 0.100405
R13393 VPWR.n2216 VPWR 0.100405
R13394 VPWR.n2225 VPWR 0.100405
R13395 VPWR.n2226 VPWR 0.100405
R13396 VPWR.n2235 VPWR 0.100405
R13397 VPWR.n2236 VPWR 0.100405
R13398 VPWR.n2245 VPWR 0.100405
R13399 VPWR.n2246 VPWR 0.100405
R13400 VPWR.n2255 VPWR 0.100405
R13401 VPWR.n2256 VPWR 0.100405
R13402 VPWR.n2265 VPWR 0.100405
R13403 VPWR VPWR.n2189 0.100405
R13404 VPWR VPWR.n2190 0.100405
R13405 VPWR VPWR.n2191 0.100405
R13406 VPWR VPWR.n2192 0.100405
R13407 VPWR VPWR.n2203 0.100405
R13408 VPWR VPWR.n2202 0.100405
R13409 VPWR VPWR.n2201 0.100405
R13410 VPWR VPWR.n2200 0.100405
R13411 VPWR VPWR.n2199 0.100405
R13412 VPWR VPWR.n2198 0.100405
R13413 VPWR VPWR.n2197 0.100405
R13414 VPWR VPWR.n2196 0.100405
R13415 VPWR VPWR.n2195 0.100405
R13416 VPWR VPWR.n2194 0.100405
R13417 VPWR VPWR.n2193 0.100405
R13418 VPWR.n2109 VPWR 0.100405
R13419 VPWR VPWR.n2118 0.100405
R13420 VPWR.n2119 VPWR 0.100405
R13421 VPWR VPWR.n2128 0.100405
R13422 VPWR.n2179 VPWR 0.100405
R13423 VPWR VPWR.n2178 0.100405
R13424 VPWR.n2169 VPWR 0.100405
R13425 VPWR VPWR.n2168 0.100405
R13426 VPWR.n2159 VPWR 0.100405
R13427 VPWR VPWR.n2158 0.100405
R13428 VPWR.n2149 VPWR 0.100405
R13429 VPWR VPWR.n2148 0.100405
R13430 VPWR.n2139 VPWR 0.100405
R13431 VPWR VPWR.n2138 0.100405
R13432 VPWR.n2129 VPWR 0.100405
R13433 VPWR.n2106 VPWR 0.100405
R13434 VPWR.n2105 VPWR 0.100405
R13435 VPWR.n2104 VPWR 0.100405
R13436 VPWR.n2103 VPWR 0.100405
R13437 VPWR.n2092 VPWR 0.100405
R13438 VPWR.n2093 VPWR 0.100405
R13439 VPWR.n2094 VPWR 0.100405
R13440 VPWR.n2095 VPWR 0.100405
R13441 VPWR.n2096 VPWR 0.100405
R13442 VPWR.n2097 VPWR 0.100405
R13443 VPWR.n2098 VPWR 0.100405
R13444 VPWR.n2099 VPWR 0.100405
R13445 VPWR.n2100 VPWR 0.100405
R13446 VPWR.n2101 VPWR 0.100405
R13447 VPWR.n2102 VPWR 0.100405
R13448 VPWR.n2089 VPWR 0.100405
R13449 VPWR.n2080 VPWR 0.100405
R13450 VPWR.n2079 VPWR 0.100405
R13451 VPWR.n2070 VPWR 0.100405
R13452 VPWR.n2019 VPWR 0.100405
R13453 VPWR.n2020 VPWR 0.100405
R13454 VPWR.n2029 VPWR 0.100405
R13455 VPWR.n2030 VPWR 0.100405
R13456 VPWR.n2039 VPWR 0.100405
R13457 VPWR.n2040 VPWR 0.100405
R13458 VPWR.n2049 VPWR 0.100405
R13459 VPWR.n2050 VPWR 0.100405
R13460 VPWR.n2059 VPWR 0.100405
R13461 VPWR.n2060 VPWR 0.100405
R13462 VPWR.n2069 VPWR 0.100405
R13463 VPWR VPWR.n1993 0.100405
R13464 VPWR VPWR.n1994 0.100405
R13465 VPWR VPWR.n1995 0.100405
R13466 VPWR VPWR.n1996 0.100405
R13467 VPWR VPWR.n2007 0.100405
R13468 VPWR VPWR.n2006 0.100405
R13469 VPWR VPWR.n2005 0.100405
R13470 VPWR VPWR.n2004 0.100405
R13471 VPWR VPWR.n2003 0.100405
R13472 VPWR VPWR.n2002 0.100405
R13473 VPWR VPWR.n2001 0.100405
R13474 VPWR VPWR.n2000 0.100405
R13475 VPWR VPWR.n1999 0.100405
R13476 VPWR VPWR.n1998 0.100405
R13477 VPWR VPWR.n1997 0.100405
R13478 VPWR.n1913 VPWR 0.100405
R13479 VPWR VPWR.n1922 0.100405
R13480 VPWR.n1923 VPWR 0.100405
R13481 VPWR VPWR.n1932 0.100405
R13482 VPWR.n1983 VPWR 0.100405
R13483 VPWR VPWR.n1982 0.100405
R13484 VPWR.n1973 VPWR 0.100405
R13485 VPWR VPWR.n1972 0.100405
R13486 VPWR.n1963 VPWR 0.100405
R13487 VPWR VPWR.n1962 0.100405
R13488 VPWR.n1953 VPWR 0.100405
R13489 VPWR VPWR.n1952 0.100405
R13490 VPWR.n1943 VPWR 0.100405
R13491 VPWR VPWR.n1942 0.100405
R13492 VPWR.n1933 VPWR 0.100405
R13493 VPWR.n1910 VPWR 0.100405
R13494 VPWR.n1909 VPWR 0.100405
R13495 VPWR.n1908 VPWR 0.100405
R13496 VPWR.n1907 VPWR 0.100405
R13497 VPWR.n1896 VPWR 0.100405
R13498 VPWR.n1897 VPWR 0.100405
R13499 VPWR.n1898 VPWR 0.100405
R13500 VPWR.n1899 VPWR 0.100405
R13501 VPWR.n1900 VPWR 0.100405
R13502 VPWR.n1901 VPWR 0.100405
R13503 VPWR.n1902 VPWR 0.100405
R13504 VPWR.n1903 VPWR 0.100405
R13505 VPWR.n1904 VPWR 0.100405
R13506 VPWR.n1905 VPWR 0.100405
R13507 VPWR.n1906 VPWR 0.100405
R13508 VPWR VPWR.n2399 0.100405
R13509 VPWR VPWR.n2398 0.100405
R13510 VPWR VPWR.n2397 0.100405
R13511 VPWR VPWR.n2396 0.100405
R13512 VPWR VPWR.n2395 0.100405
R13513 VPWR VPWR.n2394 0.100405
R13514 VPWR VPWR.n2393 0.100405
R13515 VPWR VPWR.n2392 0.100405
R13516 VPWR VPWR.n2391 0.100405
R13517 VPWR VPWR.n2390 0.100405
R13518 VPWR VPWR.n2389 0.100405
R13519 VPWR VPWR.n2388 0.100405
R13520 VPWR.n1893 VPWR 0.100405
R13521 VPWR.n1884 VPWR 0.100405
R13522 VPWR.n1883 VPWR 0.100405
R13523 VPWR.n1874 VPWR 0.100405
R13524 VPWR.n1873 VPWR 0.100405
R13525 VPWR.n1823 VPWR 0.100405
R13526 VPWR.n1824 VPWR 0.100405
R13527 VPWR.n1833 VPWR 0.100405
R13528 VPWR.n1834 VPWR 0.100405
R13529 VPWR.n1843 VPWR 0.100405
R13530 VPWR.n1844 VPWR 0.100405
R13531 VPWR.n1853 VPWR 0.100405
R13532 VPWR.n1854 VPWR 0.100405
R13533 VPWR.n1863 VPWR 0.100405
R13534 VPWR.n1864 VPWR 0.100405
R13535 VPWR.n2411 VPWR 0.100405
R13536 VPWR.n2412 VPWR 0.100405
R13537 VPWR.n2421 VPWR 0.100405
R13538 VPWR.n2422 VPWR 0.100405
R13539 VPWR.n2431 VPWR 0.100405
R13540 VPWR.n2432 VPWR 0.100405
R13541 VPWR.n2441 VPWR 0.100405
R13542 VPWR.n2442 VPWR 0.100405
R13543 VPWR.n2451 VPWR 0.100405
R13544 VPWR.n2452 VPWR 0.100405
R13545 VPWR.n2461 VPWR 0.100405
R13546 VPWR.n2462 VPWR 0.100405
R13547 VPWR.n2471 VPWR 0.100405
R13548 VPWR VPWR.n1797 0.100405
R13549 VPWR VPWR.n1798 0.100405
R13550 VPWR VPWR.n1799 0.100405
R13551 VPWR VPWR.n1800 0.100405
R13552 VPWR VPWR.n1801 0.100405
R13553 VPWR VPWR.n1802 0.100405
R13554 VPWR VPWR.n1803 0.100405
R13555 VPWR VPWR.n1804 0.100405
R13556 VPWR VPWR.n1811 0.100405
R13557 VPWR VPWR.n1810 0.100405
R13558 VPWR VPWR.n1809 0.100405
R13559 VPWR VPWR.n1808 0.100405
R13560 VPWR VPWR.n1807 0.100405
R13561 VPWR VPWR.n1806 0.100405
R13562 VPWR VPWR.n1805 0.100405
R13563 VPWR.n2498 VPWR 0.100405
R13564 VPWR.n2497 VPWR 0.100405
R13565 VPWR.n2496 VPWR 0.100405
R13566 VPWR.n2495 VPWR 0.100405
R13567 VPWR.n2494 VPWR 0.100405
R13568 VPWR.n2493 VPWR 0.100405
R13569 VPWR.n2492 VPWR 0.100405
R13570 VPWR.n2491 VPWR 0.100405
R13571 VPWR.n2490 VPWR 0.100405
R13572 VPWR.n2489 VPWR 0.100405
R13573 VPWR.n2484 VPWR 0.100405
R13574 VPWR.n2485 VPWR 0.100405
R13575 VPWR.n2486 VPWR 0.100405
R13576 VPWR.n2487 VPWR 0.100405
R13577 VPWR.n2488 VPWR 0.100405
R13578 VPWR.n1143 VPWR 0.100405
R13579 VPWR VPWR.n1540 0.100405
R13580 VPWR.n1524 VPWR 0.100405
R13581 VPWR.n1516 VPWR 0.100405
R13582 VPWR.n1510 VPWR 0.100405
R13583 VPWR.n1502 VPWR 0.100405
R13584 VPWR.n1496 VPWR 0.100405
R13585 VPWR VPWR.n1132 0.100405
R13586 VPWR.n1584 VPWR 0.100405
R13587 VPWR.n1452 VPWR 0.100405
R13588 VPWR.n1464 VPWR 0.100405
R13589 VPWR.n1043 VPWR 0.100405
R13590 VPWR.n1744 VPWR 0.100405
R13591 VPWR.n1787 VPWR 0.100405
R13592 VPWR VPWR.n1765 0.100405
R13593 VPWR.n2501 VPWR 0.100405
R13594 VPWR VPWR.n2512 0.100405
R13595 VPWR.n2513 VPWR 0.100405
R13596 VPWR VPWR.n2524 0.100405
R13597 VPWR.n2525 VPWR 0.100405
R13598 VPWR VPWR.n2536 0.100405
R13599 VPWR.n2537 VPWR 0.100405
R13600 VPWR VPWR.n2548 0.100405
R13601 VPWR.n2549 VPWR 0.100405
R13602 VPWR VPWR.n2560 0.100405
R13603 VPWR.n2561 VPWR 0.100405
R13604 VPWR VPWR.n2572 0.100405
R13605 VPWR.n2573 VPWR 0.100405
R13606 VPWR VPWR.n2584 0.100405
R13607 VPWR.n2585 VPWR 0.100405
R13608 VPWR.n1056 VPWR 0.100405
R13609 VPWR.n1754 VPWR 0.100405
R13610 VPWR.n1755 VPWR 0.100405
R13611 VPWR.n1529 VPWR 0.100405
R13612 VPWR.n1530 VPWR 0.100405
R13613 VPWR VPWR.n1528 0.100405
R13614 VPWR VPWR.n1527 0.100405
R13615 VPWR.n1514 VPWR 0.100405
R13616 VPWR VPWR.n1513 0.100405
R13617 VPWR.n1500 VPWR 0.100405
R13618 VPWR VPWR.n1499 0.100405
R13619 VPWR.n1487 VPWR 0.100405
R13620 VPWR.n1587 VPWR 0.100405
R13621 VPWR.n1588 VPWR 0.100405
R13622 VPWR.n1448 VPWR 0.100405
R13623 VPWR VPWR.n2798 0.0994583
R13624 VPWR VPWR.n2779 0.0994583
R13625 VPWR VPWR.n1326 0.0981562
R13626 VPWR.n1371 VPWR 0.0981562
R13627 VPWR.n1410 VPWR 0.0981562
R13628 VPWR.n9 VPWR 0.0968542
R13629 VPWR.n1244 VPWR 0.0968542
R13630 VPWR.n1267 VPWR 0.0968542
R13631 VPWR.n1291 VPWR 0.0968542
R13632 VPWR.n1333 VPWR 0.0968542
R13633 VPWR VPWR.n2759 0.0968542
R13634 VPWR VPWR.n2740 0.0968542
R13635 VPWR.n2718 VPWR 0.0968542
R13636 VPWR.n2682 VPWR 0.0968542
R13637 VPWR.n2645 VPWR 0.0968542
R13638 VPWR.n2608 VPWR 0.0968542
R13639 VPWR VPWR.n1044 0.0945
R13640 VPWR.n1541 VPWR 0.0945
R13641 VPWR VPWR.n1142 0.0945
R13642 VPWR VPWR.n1141 0.0945
R13643 VPWR VPWR.n1140 0.0945
R13644 VPWR VPWR.n1139 0.0945
R13645 VPWR VPWR.n1138 0.0945
R13646 VPWR.n1137 VPWR 0.0945
R13647 VPWR VPWR.n1583 0.0945
R13648 VPWR VPWR.n1131 0.0945
R13649 VPWR VPWR.n1463 0.0945
R13650 VPWR.n1451 VPWR 0.0945
R13651 VPWR VPWR.n1038 0.0945
R13652 VPWR.n1786 VPWR 0.0945
R13653 VPWR VPWR.n1027 0.0945
R13654 VPWR.n1766 VPWR 0.0945
R13655 VPWR.n1117 VPWR 0.093504
R13656 VPWR.n109 VPWR 0.093504
R13657 VPWR.n143 VPWR 0.093504
R13658 VPWR.n155 VPWR 0.093504
R13659 VPWR.n167 VPWR 0.093504
R13660 VPWR.n179 VPWR 0.093504
R13661 VPWR.n191 VPWR 0.093504
R13662 VPWR.n203 VPWR 0.093504
R13663 VPWR.n215 VPWR 0.093504
R13664 VPWR.n227 VPWR 0.093504
R13665 VPWR.n239 VPWR 0.093504
R13666 VPWR.n251 VPWR 0.093504
R13667 VPWR.n263 VPWR 0.093504
R13668 VPWR.n275 VPWR 0.093504
R13669 VPWR VPWR.n285 0.093504
R13670 VPWR.n131 VPWR 0.093504
R13671 VPWR.n120 VPWR 0.093504
R13672 VPWR VPWR.n1731 0.093504
R13673 VPWR.n1722 VPWR 0.093504
R13674 VPWR.n1710 VPWR 0.093504
R13675 VPWR.n1699 VPWR 0.093504
R13676 VPWR VPWR.n1077 0.093504
R13677 VPWR.n1683 VPWR 0.093504
R13678 VPWR.n1672 VPWR 0.093504
R13679 VPWR VPWR.n1087 0.093504
R13680 VPWR.n1656 VPWR 0.093504
R13681 VPWR.n1645 VPWR 0.093504
R13682 VPWR VPWR.n1097 0.093504
R13683 VPWR.n1629 VPWR 0.093504
R13684 VPWR.n1618 VPWR 0.093504
R13685 VPWR VPWR.n1107 0.093504
R13686 VPWR.n1602 VPWR 0.093504
R13687 VPWR.n2598 VPWR 0.0849042
R13688 VPWR.n1112 VPWR.n1109 0.0845517
R13689 VPWR.n147 VPWR.n146 0.0845517
R13690 VPWR.n159 VPWR.n158 0.0845517
R13691 VPWR.n171 VPWR.n170 0.0845517
R13692 VPWR.n183 VPWR.n182 0.0845517
R13693 VPWR.n195 VPWR.n194 0.0845517
R13694 VPWR.n207 VPWR.n206 0.0845517
R13695 VPWR.n219 VPWR.n218 0.0845517
R13696 VPWR.n231 VPWR.n230 0.0845517
R13697 VPWR.n243 VPWR.n242 0.0845517
R13698 VPWR.n255 VPWR.n254 0.0845517
R13699 VPWR.n267 VPWR.n266 0.0845517
R13700 VPWR.n279 VPWR.n278 0.0845517
R13701 VPWR.n282 VPWR.n103 0.0845517
R13702 VPWR.n113 VPWR.n112 0.0845517
R13703 VPWR.n135 VPWR.n134 0.0845517
R13704 VPWR.n124 VPWR.n123 0.0845517
R13705 VPWR.n1728 VPWR.n1067 0.0845517
R13706 VPWR.n1726 VPWR.n1725 0.0845517
R13707 VPWR.n1714 VPWR.n1713 0.0845517
R13708 VPWR.n1701 VPWR.n1700 0.0845517
R13709 VPWR.n1690 VPWR.n1078 0.0845517
R13710 VPWR.n1687 VPWR.n1686 0.0845517
R13711 VPWR.n1674 VPWR.n1673 0.0845517
R13712 VPWR.n1663 VPWR.n1088 0.0845517
R13713 VPWR.n1660 VPWR.n1659 0.0845517
R13714 VPWR.n1647 VPWR.n1646 0.0845517
R13715 VPWR.n1636 VPWR.n1098 0.0845517
R13716 VPWR.n1633 VPWR.n1632 0.0845517
R13717 VPWR.n1620 VPWR.n1619 0.0845517
R13718 VPWR.n1609 VPWR.n1108 0.0845517
R13719 VPWR.n1606 VPWR.n1605 0.0845517
R13720 VPWR.n1456 VPWR.n1451 0.0740128
R13721 VPWR.n1542 VPWR.n1044 0.071
R13722 VPWR.n1547 VPWR.n1541 0.071
R13723 VPWR.n1552 VPWR.n1142 0.071
R13724 VPWR.n1557 VPWR.n1141 0.071
R13725 VPWR.n1562 VPWR.n1140 0.071
R13726 VPWR.n1567 VPWR.n1139 0.071
R13727 VPWR.n1572 VPWR.n1138 0.071
R13728 VPWR.n1577 VPWR.n1137 0.071
R13729 VPWR.n1583 VPWR.n1582 0.071
R13730 VPWR.n1457 VPWR.n1131 0.071
R13731 VPWR.n1463 VPWR.n1462 0.071
R13732 VPWR.n1772 VPWR.n1038 0.071
R13733 VPWR.n1786 VPWR.n1785 0.071
R13734 VPWR.n1780 VPWR.n1027 0.071
R13735 VPWR.n1767 VPWR.n1766 0.071
R13736 VPWR VPWR.n1115 0.0678077
R13737 VPWR VPWR.n107 0.0678077
R13738 VPWR VPWR.n141 0.0678077
R13739 VPWR VPWR.n153 0.0678077
R13740 VPWR VPWR.n165 0.0678077
R13741 VPWR VPWR.n177 0.0678077
R13742 VPWR VPWR.n189 0.0678077
R13743 VPWR VPWR.n201 0.0678077
R13744 VPWR VPWR.n213 0.0678077
R13745 VPWR VPWR.n225 0.0678077
R13746 VPWR VPWR.n237 0.0678077
R13747 VPWR VPWR.n249 0.0678077
R13748 VPWR VPWR.n261 0.0678077
R13749 VPWR VPWR.n273 0.0678077
R13750 VPWR.n286 VPWR 0.0678077
R13751 VPWR VPWR.n129 0.0678077
R13752 VPWR VPWR.n118 0.0678077
R13753 VPWR.n1732 VPWR 0.0678077
R13754 VPWR VPWR.n1720 0.0678077
R13755 VPWR VPWR.n1708 0.0678077
R13756 VPWR VPWR.n1697 0.0678077
R13757 VPWR.n1193 VPWR 0.0678077
R13758 VPWR VPWR.n1681 0.0678077
R13759 VPWR VPWR.n1670 0.0678077
R13760 VPWR.n1207 VPWR 0.0678077
R13761 VPWR VPWR.n1654 0.0678077
R13762 VPWR VPWR.n1643 0.0678077
R13763 VPWR.n1175 VPWR 0.0678077
R13764 VPWR VPWR.n1627 0.0678077
R13765 VPWR VPWR.n1616 0.0678077
R13766 VPWR.n1124 VPWR 0.0678077
R13767 VPWR VPWR.n1600 0.0678077
R13768 VPWR.n150 VPWR 0.063
R13769 VPWR.n162 VPWR 0.063
R13770 VPWR.n174 VPWR 0.063
R13771 VPWR.n186 VPWR 0.063
R13772 VPWR.n198 VPWR 0.063
R13773 VPWR.n210 VPWR 0.063
R13774 VPWR.n222 VPWR 0.063
R13775 VPWR.n234 VPWR 0.063
R13776 VPWR.n246 VPWR 0.063
R13777 VPWR.n258 VPWR 0.063
R13778 VPWR.n270 VPWR 0.063
R13779 VPWR.n101 VPWR 0.063
R13780 VPWR.n105 VPWR 0.063
R13781 VPWR.n138 VPWR 0.063
R13782 VPWR.n115 VPWR 0.063
R13783 VPWR.n126 VPWR 0.063
R13784 VPWR.n1065 VPWR 0.063
R13785 VPWR.n1717 VPWR 0.063
R13786 VPWR.n1070 VPWR 0.063
R13787 VPWR VPWR.n1704 0.063
R13788 VPWR VPWR.n1693 0.063
R13789 VPWR VPWR.n1081 0.063
R13790 VPWR VPWR.n1677 0.063
R13791 VPWR VPWR.n1666 0.063
R13792 VPWR VPWR.n1091 0.063
R13793 VPWR VPWR.n1650 0.063
R13794 VPWR VPWR.n1639 0.063
R13795 VPWR VPWR.n1101 0.063
R13796 VPWR VPWR.n1623 0.063
R13797 VPWR VPWR.n1612 0.063
R13798 VPWR VPWR.n1111 0.063
R13799 VPWR VPWR.n1120 0.063
R13800 VPWR.n1115 VPWR 0.0608448
R13801 VPWR.n107 VPWR 0.0608448
R13802 VPWR.n141 VPWR 0.0608448
R13803 VPWR.n153 VPWR 0.0608448
R13804 VPWR.n165 VPWR 0.0608448
R13805 VPWR.n177 VPWR 0.0608448
R13806 VPWR.n189 VPWR 0.0608448
R13807 VPWR.n201 VPWR 0.0608448
R13808 VPWR.n213 VPWR 0.0608448
R13809 VPWR.n225 VPWR 0.0608448
R13810 VPWR.n237 VPWR 0.0608448
R13811 VPWR.n249 VPWR 0.0608448
R13812 VPWR.n261 VPWR 0.0608448
R13813 VPWR.n273 VPWR 0.0608448
R13814 VPWR.n286 VPWR 0.0608448
R13815 VPWR.n129 VPWR 0.0608448
R13816 VPWR.n118 VPWR 0.0608448
R13817 VPWR.n1732 VPWR 0.0608448
R13818 VPWR.n1720 VPWR 0.0608448
R13819 VPWR.n1708 VPWR 0.0608448
R13820 VPWR.n1697 VPWR 0.0608448
R13821 VPWR.n1193 VPWR 0.0608448
R13822 VPWR.n1681 VPWR 0.0608448
R13823 VPWR.n1670 VPWR 0.0608448
R13824 VPWR.n1207 VPWR 0.0608448
R13825 VPWR.n1654 VPWR 0.0608448
R13826 VPWR.n1643 VPWR 0.0608448
R13827 VPWR.n1175 VPWR 0.0608448
R13828 VPWR.n1627 VPWR 0.0608448
R13829 VPWR.n1616 VPWR 0.0608448
R13830 VPWR.n1124 VPWR 0.0608448
R13831 VPWR.n1600 VPWR 0.0608448
R13832 VPWR VPWR.n13 0.0603958
R13833 VPWR VPWR.n12 0.0603958
R13834 VPWR VPWR.n1249 0.0603958
R13835 VPWR VPWR.n1248 0.0603958
R13836 VPWR VPWR.n1272 0.0603958
R13837 VPWR VPWR.n1271 0.0603958
R13838 VPWR VPWR.n1296 0.0603958
R13839 VPWR VPWR.n1295 0.0603958
R13840 VPWR.n1332 VPWR 0.0603958
R13841 VPWR VPWR.n1331 0.0603958
R13842 VPWR.n1327 VPWR 0.0603958
R13843 VPWR.n1318 VPWR 0.0603958
R13844 VPWR VPWR.n1317 0.0603958
R13845 VPWR.n1370 VPWR 0.0603958
R13846 VPWR VPWR.n1369 0.0603958
R13847 VPWR.n1364 VPWR 0.0603958
R13848 VPWR.n1409 VPWR 0.0603958
R13849 VPWR VPWR.n1408 0.0603958
R13850 VPWR.n1403 VPWR 0.0603958
R13851 VPWR.n1440 VPWR 0.0603958
R13852 VPWR VPWR.n2800 0.0603958
R13853 VPWR VPWR.n2799 0.0603958
R13854 VPWR VPWR.n2812 0.0603958
R13855 VPWR.n2791 VPWR 0.0603958
R13856 VPWR.n2792 VPWR 0.0603958
R13857 VPWR VPWR.n2796 0.0603958
R13858 VPWR.n2771 VPWR 0.0603958
R13859 VPWR.n2772 VPWR 0.0603958
R13860 VPWR VPWR.n2777 0.0603958
R13861 VPWR.n2752 VPWR 0.0603958
R13862 VPWR.n2753 VPWR 0.0603958
R13863 VPWR VPWR.n2757 0.0603958
R13864 VPWR.n2733 VPWR 0.0603958
R13865 VPWR.n2734 VPWR 0.0603958
R13866 VPWR VPWR.n2695 0.0603958
R13867 VPWR.n2696 VPWR 0.0603958
R13868 VPWR.n2697 VPWR 0.0603958
R13869 VPWR VPWR.n2658 0.0603958
R13870 VPWR.n2659 VPWR 0.0603958
R13871 VPWR.n2660 VPWR 0.0603958
R13872 VPWR.n2624 VPWR 0.0603958
R13873 VPWR.n2627 VPWR 0.0603958
R13874 VPWR.n1770 VPWR.n1769 0.0599512
R13875 VPWR.n1041 VPWR.n1040 0.0599512
R13876 VPWR.n1545 VPWR.n1544 0.0599512
R13877 VPWR.n1550 VPWR.n1549 0.0599512
R13878 VPWR.n1555 VPWR.n1554 0.0599512
R13879 VPWR.n1560 VPWR.n1559 0.0599512
R13880 VPWR.n1565 VPWR.n1564 0.0599512
R13881 VPWR.n1570 VPWR.n1569 0.0599512
R13882 VPWR.n1575 VPWR.n1574 0.0599512
R13883 VPWR.n1580 VPWR.n1579 0.0599512
R13884 VPWR.n1135 VPWR.n1134 0.0599512
R13885 VPWR.n1460 VPWR.n1459 0.0599512
R13886 VPWR.n1455 VPWR.n1454 0.0599512
R13887 VPWR.n1775 VPWR.n1774 0.0599512
R13888 VPWR.n1783 VPWR.n1782 0.0599512
R13889 VPWR.n1779 VPWR.n1778 0.0599512
R13890 VPWR.n1118 VPWR.n1117 0.0565345
R13891 VPWR.n1112 VPWR 0.0565345
R13892 VPWR.n144 VPWR.n143 0.0565345
R13893 VPWR.n146 VPWR 0.0565345
R13894 VPWR.n156 VPWR.n155 0.0565345
R13895 VPWR.n158 VPWR 0.0565345
R13896 VPWR.n168 VPWR.n167 0.0565345
R13897 VPWR.n170 VPWR 0.0565345
R13898 VPWR.n180 VPWR.n179 0.0565345
R13899 VPWR.n182 VPWR 0.0565345
R13900 VPWR.n192 VPWR.n191 0.0565345
R13901 VPWR.n194 VPWR 0.0565345
R13902 VPWR.n204 VPWR.n203 0.0565345
R13903 VPWR.n206 VPWR 0.0565345
R13904 VPWR.n216 VPWR.n215 0.0565345
R13905 VPWR.n218 VPWR 0.0565345
R13906 VPWR.n228 VPWR.n227 0.0565345
R13907 VPWR.n230 VPWR 0.0565345
R13908 VPWR.n240 VPWR.n239 0.0565345
R13909 VPWR.n242 VPWR 0.0565345
R13910 VPWR.n252 VPWR.n251 0.0565345
R13911 VPWR.n254 VPWR 0.0565345
R13912 VPWR.n264 VPWR.n263 0.0565345
R13913 VPWR.n266 VPWR 0.0565345
R13914 VPWR.n276 VPWR.n275 0.0565345
R13915 VPWR.n278 VPWR 0.0565345
R13916 VPWR.n285 VPWR.n283 0.0565345
R13917 VPWR.n103 VPWR 0.0565345
R13918 VPWR.n110 VPWR.n109 0.0565345
R13919 VPWR.n112 VPWR 0.0565345
R13920 VPWR.n132 VPWR.n131 0.0565345
R13921 VPWR.n134 VPWR 0.0565345
R13922 VPWR.n121 VPWR.n120 0.0565345
R13923 VPWR.n123 VPWR 0.0565345
R13924 VPWR.n1731 VPWR.n1729 0.0565345
R13925 VPWR.n1067 VPWR 0.0565345
R13926 VPWR.n1723 VPWR.n1722 0.0565345
R13927 VPWR.n1725 VPWR 0.0565345
R13928 VPWR.n1711 VPWR.n1710 0.0565345
R13929 VPWR.n1713 VPWR 0.0565345
R13930 VPWR.n1702 VPWR.n1699 0.0565345
R13931 VPWR.n1700 VPWR 0.0565345
R13932 VPWR.n1691 VPWR.n1077 0.0565345
R13933 VPWR.n1078 VPWR 0.0565345
R13934 VPWR.n1684 VPWR.n1683 0.0565345
R13935 VPWR.n1686 VPWR 0.0565345
R13936 VPWR.n1675 VPWR.n1672 0.0565345
R13937 VPWR.n1673 VPWR 0.0565345
R13938 VPWR.n1664 VPWR.n1087 0.0565345
R13939 VPWR.n1088 VPWR 0.0565345
R13940 VPWR.n1657 VPWR.n1656 0.0565345
R13941 VPWR.n1659 VPWR 0.0565345
R13942 VPWR.n1648 VPWR.n1645 0.0565345
R13943 VPWR.n1646 VPWR 0.0565345
R13944 VPWR.n1637 VPWR.n1097 0.0565345
R13945 VPWR.n1098 VPWR 0.0565345
R13946 VPWR.n1630 VPWR.n1629 0.0565345
R13947 VPWR.n1632 VPWR 0.0565345
R13948 VPWR.n1621 VPWR.n1618 0.0565345
R13949 VPWR.n1619 VPWR 0.0565345
R13950 VPWR.n1610 VPWR.n1107 0.0565345
R13951 VPWR.n1108 VPWR 0.0565345
R13952 VPWR.n1603 VPWR.n1602 0.0565345
R13953 VPWR.n1605 VPWR 0.0565345
R13954 VPWR.n1769 VPWR 0.0469286
R13955 VPWR.n1040 VPWR 0.0469286
R13956 VPWR.n1544 VPWR 0.0469286
R13957 VPWR.n1549 VPWR 0.0469286
R13958 VPWR.n1554 VPWR 0.0469286
R13959 VPWR.n1559 VPWR 0.0469286
R13960 VPWR.n1564 VPWR 0.0469286
R13961 VPWR.n1569 VPWR 0.0469286
R13962 VPWR.n1574 VPWR 0.0469286
R13963 VPWR.n1579 VPWR 0.0469286
R13964 VPWR.n1134 VPWR 0.0469286
R13965 VPWR.n1459 VPWR 0.0469286
R13966 VPWR.n1454 VPWR 0.0469286
R13967 VPWR.n1774 VPWR 0.0469286
R13968 VPWR.n1782 VPWR 0.0469286
R13969 VPWR.n1778 VPWR 0.0469286
R13970 VPWR.n1769 VPWR 0.0401341
R13971 VPWR.n1040 VPWR 0.0401341
R13972 VPWR.n1544 VPWR 0.0401341
R13973 VPWR.n1549 VPWR 0.0401341
R13974 VPWR.n1554 VPWR 0.0401341
R13975 VPWR.n1559 VPWR 0.0401341
R13976 VPWR.n1564 VPWR 0.0401341
R13977 VPWR.n1569 VPWR 0.0401341
R13978 VPWR.n1574 VPWR 0.0401341
R13979 VPWR.n1579 VPWR 0.0401341
R13980 VPWR.n1134 VPWR 0.0401341
R13981 VPWR.n1459 VPWR 0.0401341
R13982 VPWR.n1454 VPWR 0.0401341
R13983 VPWR.n1774 VPWR 0.0401341
R13984 VPWR.n1782 VPWR 0.0401341
R13985 VPWR.n1778 VPWR 0.0401341
R13986 VPWR.n13 VPWR 0.0382604
R13987 VPWR.n1249 VPWR 0.0382604
R13988 VPWR.n1272 VPWR 0.0382604
R13989 VPWR.n1296 VPWR 0.0382604
R13990 VPWR.n1331 VPWR 0.0382604
R13991 VPWR.n1369 VPWR 0.0382604
R13992 VPWR.n1408 VPWR 0.0382604
R13993 VPWR.n1445 VPWR 0.0382604
R13994 VPWR.n20 VPWR 0.0375125
R13995 VPWR.n20 VPWR 0.0373589
R13996 VPWR.n1118 VPWR.n1109 0.0349828
R13997 VPWR.n147 VPWR.n144 0.0349828
R13998 VPWR.n159 VPWR.n156 0.0349828
R13999 VPWR.n171 VPWR.n168 0.0349828
R14000 VPWR.n183 VPWR.n180 0.0349828
R14001 VPWR.n195 VPWR.n192 0.0349828
R14002 VPWR.n207 VPWR.n204 0.0349828
R14003 VPWR.n219 VPWR.n216 0.0349828
R14004 VPWR.n231 VPWR.n228 0.0349828
R14005 VPWR.n243 VPWR.n240 0.0349828
R14006 VPWR.n255 VPWR.n252 0.0349828
R14007 VPWR.n267 VPWR.n264 0.0349828
R14008 VPWR.n279 VPWR.n276 0.0349828
R14009 VPWR.n283 VPWR.n282 0.0349828
R14010 VPWR.n113 VPWR.n110 0.0349828
R14011 VPWR.n135 VPWR.n132 0.0349828
R14012 VPWR.n124 VPWR.n121 0.0349828
R14013 VPWR.n1729 VPWR.n1728 0.0349828
R14014 VPWR.n1726 VPWR.n1723 0.0349828
R14015 VPWR.n1714 VPWR.n1711 0.0349828
R14016 VPWR.n1702 VPWR.n1701 0.0349828
R14017 VPWR.n1691 VPWR.n1690 0.0349828
R14018 VPWR.n1687 VPWR.n1684 0.0349828
R14019 VPWR.n1675 VPWR.n1674 0.0349828
R14020 VPWR.n1664 VPWR.n1663 0.0349828
R14021 VPWR.n1660 VPWR.n1657 0.0349828
R14022 VPWR.n1648 VPWR.n1647 0.0349828
R14023 VPWR.n1637 VPWR.n1636 0.0349828
R14024 VPWR.n1633 VPWR.n1630 0.0349828
R14025 VPWR.n1621 VPWR.n1620 0.0349828
R14026 VPWR.n1610 VPWR.n1609 0.0349828
R14027 VPWR.n1606 VPWR.n1603 0.0349828
R14028 VPWR.n2504 VPWR.n2503 0.0340366
R14029 VPWR.n2570 VPWR.n2569 0.0340366
R14030 VPWR.n2510 VPWR.n2509 0.0340366
R14031 VPWR.n2552 VPWR.n2551 0.0340366
R14032 VPWR.n2546 VPWR.n2545 0.0340366
R14033 VPWR.n2534 VPWR.n2533 0.0340366
R14034 VPWR.n2528 VPWR.n2527 0.0340366
R14035 VPWR.n1223 VPWR.n1222 0.0340366
R14036 VPWR.n2522 VPWR.n2521 0.0340366
R14037 VPWR.n1486 VPWR.n1102 0.0340366
R14038 VPWR.n1174 VPWR.n1094 0.0340366
R14039 VPWR.n2540 VPWR.n2539 0.0340366
R14040 VPWR.n1165 VPWR.n1092 0.0340366
R14041 VPWR.n1211 VPWR.n1164 0.0340366
R14042 VPWR.n2516 VPWR.n2515 0.0340366
R14043 VPWR.n1129 VPWR.n1104 0.0340366
R14044 VPWR.n1155 VPWR.n1084 0.0340366
R14045 VPWR.n2558 VPWR.n2557 0.0340366
R14046 VPWR.n1144 VPWR.n1082 0.0340366
R14047 VPWR.n1591 VPWR.n1590 0.0340366
R14048 VPWR.n2564 VPWR.n2563 0.0340366
R14049 VPWR.n1197 VPWR.n1154 0.0340366
R14050 VPWR.n1074 VPWR.n1073 0.0340366
R14051 VPWR.n1743 VPWR.n1742 0.0340366
R14052 VPWR.n1071 VPWR.n1054 0.0340366
R14053 VPWR.n2576 VPWR.n2575 0.0340366
R14054 VPWR.n2582 VPWR.n2581 0.0340366
R14055 VPWR.n2593 VPWR.n2592 0.0340366
R14056 VPWR.n2588 VPWR.n2587 0.0340366
R14057 VPWR.n1737 VPWR.n1736 0.0340366
R14058 VPWR.n1063 VPWR.n1060 0.0340366
R14059 VPWR.n1596 VPWR.n1121 0.0340366
R14060 VPWR.n2628 VPWR.n2598 0.0320292
R14061 VPWR.n2800 VPWR 0.03175
R14062 VPWR VPWR.n2791 0.03175
R14063 VPWR VPWR.n2771 0.03175
R14064 VPWR VPWR.n2752 0.03175
R14065 VPWR VPWR.n2733 0.03175
R14066 VPWR VPWR.n2696 0.03175
R14067 VPWR VPWR.n2659 0.03175
R14068 VPWR VPWR.n2627 0.03175
R14069 VPWR.n2598 VPWR.n2597 0.0240975
R14070 VPWR.n2597 VPWR.n20 0.0240975
R14071 VPWR.n2814 VPWR 0.024
R14072 VPWR.n14 VPWR 0.0239375
R14073 VPWR.n12 VPWR 0.0239375
R14074 VPWR.n1250 VPWR 0.0239375
R14075 VPWR.n1248 VPWR 0.0239375
R14076 VPWR.n1271 VPWR 0.0239375
R14077 VPWR.n1295 VPWR 0.0239375
R14078 VPWR.n2753 VPWR 0.0239375
R14079 VPWR.n2503 VPWR 0.0233659
R14080 VPWR.n1466 VPWR 0.0233659
R14081 VPWR.n352 VPWR 0.0233659
R14082 VPWR.n2570 VPWR 0.0233659
R14083 VPWR.n1533 VPWR 0.0233659
R14084 VPWR.n347 VPWR 0.0233659
R14085 VPWR.n2510 VPWR 0.0233659
R14086 VPWR.n964 VPWR 0.0233659
R14087 VPWR.n2479 VPWR 0.0233659
R14088 VPWR.n2474 VPWR 0.0233659
R14089 VPWR.n319 VPWR 0.0233659
R14090 VPWR.n2551 VPWR 0.0233659
R14091 VPWR.n972 VPWR 0.0233659
R14092 VPWR.n2444 VPWR 0.0233659
R14093 VPWR.n323 VPWR 0.0233659
R14094 VPWR.n2546 VPWR 0.0233659
R14095 VPWR.n1891 VPWR 0.0233659
R14096 VPWR.n1886 VPWR 0.0233659
R14097 VPWR.n1881 VPWR 0.0233659
R14098 VPWR.n388 VPWR 0.0233659
R14099 VPWR.n392 VPWR 0.0233659
R14100 VPWR.n396 VPWR 0.0233659
R14101 VPWR.n2454 VPWR 0.0233659
R14102 VPWR.n331 VPWR 0.0233659
R14103 VPWR.n2534 VPWR 0.0233659
R14104 VPWR.n1876 VPWR 0.0233659
R14105 VPWR.n404 VPWR 0.0233659
R14106 VPWR.n2459 VPWR 0.0233659
R14107 VPWR.n335 VPWR 0.0233659
R14108 VPWR.n2527 VPWR 0.0233659
R14109 VPWR.n2307 VPWR 0.0233659
R14110 VPWR.n2312 VPWR 0.0233659
R14111 VPWR.n2317 VPWR 0.0233659
R14112 VPWR.n2322 VPWR 0.0233659
R14113 VPWR.n2332 VPWR 0.0233659
R14114 VPWR.n2337 VPWR 0.0233659
R14115 VPWR.n2342 VPWR 0.0233659
R14116 VPWR.n2347 VPWR 0.0233659
R14117 VPWR.n2352 VPWR 0.0233659
R14118 VPWR.n2357 VPWR 0.0233659
R14119 VPWR.n2362 VPWR 0.0233659
R14120 VPWR.n2367 VPWR 0.0233659
R14121 VPWR.n2372 VPWR 0.0233659
R14122 VPWR.n2377 VPWR 0.0233659
R14123 VPWR.n2381 VPWR 0.0233659
R14124 VPWR.n2327 VPWR 0.0233659
R14125 VPWR.n544 VPWR 0.0233659
R14126 VPWR.n539 VPWR 0.0233659
R14127 VPWR.n535 VPWR 0.0233659
R14128 VPWR.n531 VPWR 0.0233659
R14129 VPWR.n523 VPWR 0.0233659
R14130 VPWR.n519 VPWR 0.0233659
R14131 VPWR.n515 VPWR 0.0233659
R14132 VPWR.n511 VPWR 0.0233659
R14133 VPWR.n507 VPWR 0.0233659
R14134 VPWR.n503 VPWR 0.0233659
R14135 VPWR.n499 VPWR 0.0233659
R14136 VPWR.n495 VPWR 0.0233659
R14137 VPWR.n491 VPWR 0.0233659
R14138 VPWR.n487 VPWR 0.0233659
R14139 VPWR.n484 VPWR 0.0233659
R14140 VPWR.n527 VPWR 0.0233659
R14141 VPWR.n2283 VPWR 0.0233659
R14142 VPWR.n2278 VPWR 0.0233659
R14143 VPWR.n2273 VPWR 0.0233659
R14144 VPWR.n2268 VPWR 0.0233659
R14145 VPWR.n2258 VPWR 0.0233659
R14146 VPWR.n2253 VPWR 0.0233659
R14147 VPWR.n2248 VPWR 0.0233659
R14148 VPWR.n2243 VPWR 0.0233659
R14149 VPWR.n2238 VPWR 0.0233659
R14150 VPWR.n2233 VPWR 0.0233659
R14151 VPWR.n2228 VPWR 0.0233659
R14152 VPWR.n2223 VPWR 0.0233659
R14153 VPWR.n2218 VPWR 0.0233659
R14154 VPWR.n2213 VPWR 0.0233659
R14155 VPWR.n2209 VPWR 0.0233659
R14156 VPWR.n2263 VPWR 0.0233659
R14157 VPWR.n580 VPWR 0.0233659
R14158 VPWR.n584 VPWR 0.0233659
R14159 VPWR.n588 VPWR 0.0233659
R14160 VPWR.n592 VPWR 0.0233659
R14161 VPWR.n600 VPWR 0.0233659
R14162 VPWR.n604 VPWR 0.0233659
R14163 VPWR.n608 VPWR 0.0233659
R14164 VPWR.n612 VPWR 0.0233659
R14165 VPWR.n616 VPWR 0.0233659
R14166 VPWR.n620 VPWR 0.0233659
R14167 VPWR.n624 VPWR 0.0233659
R14168 VPWR.n628 VPWR 0.0233659
R14169 VPWR.n632 VPWR 0.0233659
R14170 VPWR.n636 VPWR 0.0233659
R14171 VPWR.n640 VPWR 0.0233659
R14172 VPWR.n596 VPWR 0.0233659
R14173 VPWR.n2111 VPWR 0.0233659
R14174 VPWR.n2116 VPWR 0.0233659
R14175 VPWR.n2121 VPWR 0.0233659
R14176 VPWR.n2126 VPWR 0.0233659
R14177 VPWR.n2136 VPWR 0.0233659
R14178 VPWR.n2141 VPWR 0.0233659
R14179 VPWR.n2146 VPWR 0.0233659
R14180 VPWR.n2151 VPWR 0.0233659
R14181 VPWR.n2156 VPWR 0.0233659
R14182 VPWR.n2161 VPWR 0.0233659
R14183 VPWR.n2166 VPWR 0.0233659
R14184 VPWR.n2171 VPWR 0.0233659
R14185 VPWR.n2176 VPWR 0.0233659
R14186 VPWR.n2181 VPWR 0.0233659
R14187 VPWR.n2185 VPWR 0.0233659
R14188 VPWR.n2131 VPWR 0.0233659
R14189 VPWR.n736 VPWR 0.0233659
R14190 VPWR.n731 VPWR 0.0233659
R14191 VPWR.n727 VPWR 0.0233659
R14192 VPWR.n723 VPWR 0.0233659
R14193 VPWR.n715 VPWR 0.0233659
R14194 VPWR.n711 VPWR 0.0233659
R14195 VPWR.n707 VPWR 0.0233659
R14196 VPWR.n703 VPWR 0.0233659
R14197 VPWR.n699 VPWR 0.0233659
R14198 VPWR.n695 VPWR 0.0233659
R14199 VPWR.n691 VPWR 0.0233659
R14200 VPWR.n687 VPWR 0.0233659
R14201 VPWR.n683 VPWR 0.0233659
R14202 VPWR.n679 VPWR 0.0233659
R14203 VPWR.n676 VPWR 0.0233659
R14204 VPWR.n719 VPWR 0.0233659
R14205 VPWR.n2087 VPWR 0.0233659
R14206 VPWR.n2082 VPWR 0.0233659
R14207 VPWR.n2077 VPWR 0.0233659
R14208 VPWR.n2072 VPWR 0.0233659
R14209 VPWR.n2062 VPWR 0.0233659
R14210 VPWR.n2057 VPWR 0.0233659
R14211 VPWR.n2052 VPWR 0.0233659
R14212 VPWR.n2047 VPWR 0.0233659
R14213 VPWR.n2042 VPWR 0.0233659
R14214 VPWR.n2037 VPWR 0.0233659
R14215 VPWR.n2032 VPWR 0.0233659
R14216 VPWR.n2027 VPWR 0.0233659
R14217 VPWR.n2022 VPWR 0.0233659
R14218 VPWR.n2017 VPWR 0.0233659
R14219 VPWR.n2013 VPWR 0.0233659
R14220 VPWR.n2067 VPWR 0.0233659
R14221 VPWR.n772 VPWR 0.0233659
R14222 VPWR.n776 VPWR 0.0233659
R14223 VPWR.n780 VPWR 0.0233659
R14224 VPWR.n784 VPWR 0.0233659
R14225 VPWR.n792 VPWR 0.0233659
R14226 VPWR.n796 VPWR 0.0233659
R14227 VPWR.n800 VPWR 0.0233659
R14228 VPWR.n804 VPWR 0.0233659
R14229 VPWR.n808 VPWR 0.0233659
R14230 VPWR.n812 VPWR 0.0233659
R14231 VPWR.n816 VPWR 0.0233659
R14232 VPWR.n820 VPWR 0.0233659
R14233 VPWR.n824 VPWR 0.0233659
R14234 VPWR.n828 VPWR 0.0233659
R14235 VPWR.n832 VPWR 0.0233659
R14236 VPWR.n788 VPWR 0.0233659
R14237 VPWR.n1915 VPWR 0.0233659
R14238 VPWR.n1920 VPWR 0.0233659
R14239 VPWR.n1925 VPWR 0.0233659
R14240 VPWR.n1930 VPWR 0.0233659
R14241 VPWR.n1940 VPWR 0.0233659
R14242 VPWR.n1945 VPWR 0.0233659
R14243 VPWR.n1950 VPWR 0.0233659
R14244 VPWR.n1955 VPWR 0.0233659
R14245 VPWR.n1960 VPWR 0.0233659
R14246 VPWR.n1965 VPWR 0.0233659
R14247 VPWR.n1970 VPWR 0.0233659
R14248 VPWR.n1975 VPWR 0.0233659
R14249 VPWR.n1980 VPWR 0.0233659
R14250 VPWR.n1985 VPWR 0.0233659
R14251 VPWR.n1989 VPWR 0.0233659
R14252 VPWR.n1935 VPWR 0.0233659
R14253 VPWR.n928 VPWR 0.0233659
R14254 VPWR.n923 VPWR 0.0233659
R14255 VPWR.n919 VPWR 0.0233659
R14256 VPWR.n915 VPWR 0.0233659
R14257 VPWR.n907 VPWR 0.0233659
R14258 VPWR.n903 VPWR 0.0233659
R14259 VPWR.n899 VPWR 0.0233659
R14260 VPWR.n895 VPWR 0.0233659
R14261 VPWR.n891 VPWR 0.0233659
R14262 VPWR.n887 VPWR 0.0233659
R14263 VPWR.n883 VPWR 0.0233659
R14264 VPWR.n879 VPWR 0.0233659
R14265 VPWR.n875 VPWR 0.0233659
R14266 VPWR.n871 VPWR 0.0233659
R14267 VPWR.n868 VPWR 0.0233659
R14268 VPWR.n911 VPWR 0.0233659
R14269 VPWR.n1871 VPWR 0.0233659
R14270 VPWR.n980 VPWR 0.0233659
R14271 VPWR.n1495 VPWR 0.0233659
R14272 VPWR.n1223 VPWR 0.0233659
R14273 VPWR.n400 VPWR 0.0233659
R14274 VPWR.n2464 VPWR 0.0233659
R14275 VPWR.n339 VPWR 0.0233659
R14276 VPWR.n2522 VPWR 0.0233659
R14277 VPWR.n976 VPWR 0.0233659
R14278 VPWR.n1490 VPWR 0.0233659
R14279 VPWR.n1486 VPWR 0.0233659
R14280 VPWR.n1866 VPWR 0.0233659
R14281 VPWR.n984 VPWR 0.0233659
R14282 VPWR.n1504 VPWR 0.0233659
R14283 VPWR.n1174 VPWR 0.0233659
R14284 VPWR.n408 VPWR 0.0233659
R14285 VPWR.n416 VPWR 0.0233659
R14286 VPWR.n420 VPWR 0.0233659
R14287 VPWR.n424 VPWR 0.0233659
R14288 VPWR.n428 VPWR 0.0233659
R14289 VPWR.n432 VPWR 0.0233659
R14290 VPWR.n436 VPWR 0.0233659
R14291 VPWR.n440 VPWR 0.0233659
R14292 VPWR.n444 VPWR 0.0233659
R14293 VPWR.n448 VPWR 0.0233659
R14294 VPWR.n412 VPWR 0.0233659
R14295 VPWR.n2449 VPWR 0.0233659
R14296 VPWR.n327 VPWR 0.0233659
R14297 VPWR.n2539 VPWR 0.0233659
R14298 VPWR.n988 VPWR 0.0233659
R14299 VPWR.n1509 VPWR 0.0233659
R14300 VPWR.n1165 VPWR 0.0233659
R14301 VPWR.n1861 VPWR 0.0233659
R14302 VPWR.n1851 VPWR 0.0233659
R14303 VPWR.n1846 VPWR 0.0233659
R14304 VPWR.n1841 VPWR 0.0233659
R14305 VPWR.n1836 VPWR 0.0233659
R14306 VPWR.n1831 VPWR 0.0233659
R14307 VPWR.n1826 VPWR 0.0233659
R14308 VPWR.n1821 VPWR 0.0233659
R14309 VPWR.n1817 VPWR 0.0233659
R14310 VPWR.n1856 VPWR 0.0233659
R14311 VPWR.n992 VPWR 0.0233659
R14312 VPWR.n1518 VPWR 0.0233659
R14313 VPWR.n1164 VPWR 0.0233659
R14314 VPWR.n2469 VPWR 0.0233659
R14315 VPWR.n343 VPWR 0.0233659
R14316 VPWR.n2515 VPWR 0.0233659
R14317 VPWR.n1130 VPWR 0.0233659
R14318 VPWR.n1129 VPWR 0.0233659
R14319 VPWR.n996 VPWR 0.0233659
R14320 VPWR.n1523 VPWR 0.0233659
R14321 VPWR.n1155 VPWR 0.0233659
R14322 VPWR.n2439 VPWR 0.0233659
R14323 VPWR.n2429 VPWR 0.0233659
R14324 VPWR.n2424 VPWR 0.0233659
R14325 VPWR.n2419 VPWR 0.0233659
R14326 VPWR.n2414 VPWR 0.0233659
R14327 VPWR.n2409 VPWR 0.0233659
R14328 VPWR.n2405 VPWR 0.0233659
R14329 VPWR.n2434 VPWR 0.0233659
R14330 VPWR.n315 VPWR 0.0233659
R14331 VPWR.n2558 VPWR 0.0233659
R14332 VPWR.n1538 VPWR 0.0233659
R14333 VPWR.n1144 VPWR 0.0233659
R14334 VPWR.n1000 VPWR 0.0233659
R14335 VPWR.n1004 VPWR 0.0233659
R14336 VPWR.n1008 VPWR 0.0233659
R14337 VPWR.n1012 VPWR 0.0233659
R14338 VPWR.n1016 VPWR 0.0233659
R14339 VPWR.n1020 VPWR 0.0233659
R14340 VPWR.n1024 VPWR 0.0233659
R14341 VPWR.n968 VPWR 0.0233659
R14342 VPWR.n1473 VPWR 0.0233659
R14343 VPWR.n1590 VPWR 0.0233659
R14344 VPWR.n311 VPWR 0.0233659
R14345 VPWR.n2563 VPWR 0.0233659
R14346 VPWR.n1154 VPWR 0.0233659
R14347 VPWR.n1763 VPWR 0.0233659
R14348 VPWR.n1073 VPWR 0.0233659
R14349 VPWR.n307 VPWR 0.0233659
R14350 VPWR.n303 VPWR 0.0233659
R14351 VPWR.n295 VPWR 0.0233659
R14352 VPWR.n292 VPWR 0.0233659
R14353 VPWR.n299 VPWR 0.0233659
R14354 VPWR.n1743 VPWR 0.0233659
R14355 VPWR.n1751 VPWR 0.0233659
R14356 VPWR.n1789 VPWR 0.0233659
R14357 VPWR.n1793 VPWR 0.0233659
R14358 VPWR.n1758 VPWR 0.0233659
R14359 VPWR.n1054 VPWR 0.0233659
R14360 VPWR.n2575 VPWR 0.0233659
R14361 VPWR.n2582 VPWR 0.0233659
R14362 VPWR.n2593 VPWR 0.0233659
R14363 VPWR.n2587 VPWR 0.0233659
R14364 VPWR.n1736 VPWR 0.0233659
R14365 VPWR.n1060 VPWR 0.0233659
R14366 VPWR.n1121 VPWR 0.0233659
R14367 VPWR.n1336 VPWR 0.0226354
R14368 VPWR.n1327 VPWR 0.0226354
R14369 VPWR.n1413 VPWR 0.0226354
R14370 VPWR.n2772 VPWR 0.0226354
R14371 VPWR VPWR.n2732 0.0226354
R14372 VPWR VPWR.n2702 0.0226354
R14373 VPWR VPWR.n2664 0.0226354
R14374 VPWR VPWR.n64 0.0220517
R14375 VPWR VPWR.n67 0.0220517
R14376 VPWR VPWR.n70 0.0220517
R14377 VPWR VPWR.n73 0.0220517
R14378 VPWR VPWR.n76 0.0220517
R14379 VPWR VPWR.n79 0.0220517
R14380 VPWR VPWR.n82 0.0220517
R14381 VPWR VPWR.n85 0.0220517
R14382 VPWR VPWR.n88 0.0220517
R14383 VPWR VPWR.n91 0.0220517
R14384 VPWR VPWR.n94 0.0220517
R14385 VPWR VPWR.n97 0.0220517
R14386 VPWR.n289 VPWR 0.0220517
R14387 VPWR VPWR.n61 0.0220517
R14388 VPWR VPWR.n58 0.0220517
R14389 VPWR.n1735 VPWR 0.0220517
R14390 VPWR VPWR.n1057 0.0220517
R14391 VPWR.n1705 VPWR 0.0220517
R14392 VPWR.n1694 VPWR 0.0220517
R14393 VPWR.n1196 VPWR 0.0220517
R14394 VPWR.n1678 VPWR 0.0220517
R14395 VPWR.n1667 VPWR 0.0220517
R14396 VPWR.n1210 VPWR 0.0220517
R14397 VPWR.n1651 VPWR 0.0220517
R14398 VPWR.n1640 VPWR 0.0220517
R14399 VPWR.n1178 VPWR 0.0220517
R14400 VPWR.n1624 VPWR 0.0220517
R14401 VPWR.n1613 VPWR 0.0220517
R14402 VPWR.n1127 VPWR 0.0220517
R14403 VPWR.n1597 VPWR 0.0220517
R14404 VPWR.n1273 VPWR 0.0213333
R14405 VPWR.n1297 VPWR 0.0213333
R14406 VPWR.n1311 VPWR 0.0213333
R14407 VPWR.n1375 VPWR 0.0213333
R14408 VPWR.n1347 VPWR 0.0213333
R14409 VPWR.n1386 VPWR 0.0213333
R14410 VPWR.n1423 VPWR 0.0213333
R14411 VPWR.n2806 VPWR 0.0213333
R14412 VPWR.n2799 VPWR 0.0213333
R14413 VPWR VPWR.n2790 0.0213333
R14414 VPWR.n2792 VPWR 0.0213333
R14415 VPWR VPWR.n2770 0.0213333
R14416 VPWR VPWR.n2751 0.0213333
R14417 VPWR VPWR.n2738 0.0213333
R14418 VPWR.n2500 VPWR 0.0196917
R14419 VPWR.n24 VPWR 0.0143889
R14420 VPWR VPWR.n19 0.0099
R14421 VPWR VPWR.n1604 0.00397222
R14422 VPWR VPWR.n1105 0.00397222
R14423 VPWR VPWR.n1103 0.00397222
R14424 VPWR VPWR.n1631 0.00397222
R14425 VPWR VPWR.n1095 0.00397222
R14426 VPWR VPWR.n1093 0.00397222
R14427 VPWR VPWR.n1658 0.00397222
R14428 VPWR VPWR.n1085 0.00397222
R14429 VPWR VPWR.n1083 0.00397222
R14430 VPWR VPWR.n1685 0.00397222
R14431 VPWR VPWR.n1075 0.00397222
R14432 VPWR VPWR.n1072 0.00397222
R14433 VPWR VPWR.n1712 0.00397222
R14434 VPWR VPWR.n1724 0.00397222
R14435 VPWR.n1113 VPWR 0.00397222
R14436 VPWR VPWR.n1066 0.00397222
R14437 VPWR VPWR.n122 0.00397222
R14438 VPWR VPWR.n111 0.00397222
R14439 VPWR VPWR.n102 0.00397222
R14440 VPWR VPWR.n277 0.00397222
R14441 VPWR VPWR.n265 0.00397222
R14442 VPWR VPWR.n253 0.00397222
R14443 VPWR VPWR.n241 0.00397222
R14444 VPWR VPWR.n229 0.00397222
R14445 VPWR VPWR.n217 0.00397222
R14446 VPWR VPWR.n205 0.00397222
R14447 VPWR VPWR.n193 0.00397222
R14448 VPWR VPWR.n181 0.00397222
R14449 VPWR VPWR.n169 0.00397222
R14450 VPWR VPWR.n157 0.00397222
R14451 VPWR VPWR.n145 0.00397222
R14452 VPWR VPWR.n133 0.00397222
R14453 VPWR.n1462 VPWR.n1461 0.00351282
R14454 VPWR.n1457 VPWR.n1136 0.00351282
R14455 VPWR.n1582 VPWR.n1581 0.00351282
R14456 VPWR.n1577 VPWR.n1576 0.00351282
R14457 VPWR.n1572 VPWR.n1571 0.00351282
R14458 VPWR.n1567 VPWR.n1566 0.00351282
R14459 VPWR.n1562 VPWR.n1561 0.00351282
R14460 VPWR.n1557 VPWR.n1556 0.00351282
R14461 VPWR.n1552 VPWR.n1551 0.00351282
R14462 VPWR.n1547 VPWR.n1546 0.00351282
R14463 VPWR.n1542 VPWR.n1042 0.00351282
R14464 VPWR.n1785 VPWR.n1784 0.00351282
R14465 VPWR.n1776 VPWR.n1772 0.00351282
R14466 VPWR.n1771 VPWR.n1767 0.00351282
R14467 VPWR.n141 VPWR.n140 0.00265517
R14468 VPWR.n153 VPWR.n152 0.00265517
R14469 VPWR.n165 VPWR.n164 0.00265517
R14470 VPWR.n177 VPWR.n176 0.00265517
R14471 VPWR.n189 VPWR.n188 0.00265517
R14472 VPWR.n201 VPWR.n200 0.00265517
R14473 VPWR.n213 VPWR.n212 0.00265517
R14474 VPWR.n225 VPWR.n224 0.00265517
R14475 VPWR.n237 VPWR.n236 0.00265517
R14476 VPWR.n249 VPWR.n248 0.00265517
R14477 VPWR.n261 VPWR.n260 0.00265517
R14478 VPWR.n273 VPWR.n272 0.00265517
R14479 VPWR.n288 VPWR.n286 0.00265517
R14480 VPWR.n129 VPWR.n128 0.00265517
R14481 VPWR.n118 VPWR.n117 0.00265517
R14482 VPWR.n1734 VPWR.n1732 0.00265517
R14483 VPWR.n1720 VPWR.n1719 0.00265517
R14484 VPWR.n1708 VPWR.n1707 0.00265517
R14485 VPWR.n1697 VPWR.n1696 0.00265517
R14486 VPWR.n1195 VPWR.n1193 0.00265517
R14487 VPWR.n1681 VPWR.n1680 0.00265517
R14488 VPWR.n1670 VPWR.n1669 0.00265517
R14489 VPWR.n1209 VPWR.n1207 0.00265517
R14490 VPWR.n1654 VPWR.n1653 0.00265517
R14491 VPWR.n1643 VPWR.n1642 0.00265517
R14492 VPWR.n1177 VPWR.n1175 0.00265517
R14493 VPWR.n1627 VPWR.n1626 0.00265517
R14494 VPWR.n1616 VPWR.n1615 0.00265517
R14495 VPWR.n1126 VPWR.n1124 0.00265517
R14496 VPWR.n1600 VPWR.n1599 0.00265517
R14497 Iout.n1020 Iout.t64 239.927
R14498 Iout.n509 Iout.t33 239.927
R14499 Iout.n513 Iout.t9 239.927
R14500 Iout.n507 Iout.t86 239.927
R14501 Iout.n504 Iout.t39 239.927
R14502 Iout.n500 Iout.t249 239.927
R14503 Iout.n192 Iout.t234 239.927
R14504 Iout.n195 Iout.t133 239.927
R14505 Iout.n199 Iout.t20 239.927
R14506 Iout.n202 Iout.t35 239.927
R14507 Iout.n206 Iout.t61 239.927
R14508 Iout.n210 Iout.t205 239.927
R14509 Iout.n214 Iout.t62 239.927
R14510 Iout.n218 Iout.t160 239.927
R14511 Iout.n222 Iout.t139 239.927
R14512 Iout.n226 Iout.t75 239.927
R14513 Iout.n232 Iout.t117 239.927
R14514 Iout.n235 Iout.t72 239.927
R14515 Iout.n238 Iout.t3 239.927
R14516 Iout.n241 Iout.t118 239.927
R14517 Iout.n244 Iout.t216 239.927
R14518 Iout.n247 Iout.t42 239.927
R14519 Iout.n250 Iout.t178 239.927
R14520 Iout.n255 Iout.t110 239.927
R14521 Iout.n252 Iout.t121 239.927
R14522 Iout.n489 Iout.t124 239.927
R14523 Iout.n494 Iout.t93 239.927
R14524 Iout.n491 Iout.t203 239.927
R14525 Iout.n519 Iout.t95 239.927
R14526 Iout.n149 Iout.t153 239.927
R14527 Iout.n146 Iout.t145 239.927
R14528 Iout.n1010 Iout.t200 239.927
R14529 Iout.n1007 Iout.t63 239.927
R14530 Iout.n140 Iout.t135 239.927
R14531 Iout.n143 Iout.t91 239.927
R14532 Iout.n525 Iout.t214 239.927
R14533 Iout.n480 Iout.t143 239.927
R14534 Iout.n483 Iout.t26 239.927
R14535 Iout.n478 Iout.t168 239.927
R14536 Iout.n259 Iout.t13 239.927
R14537 Iout.n186 Iout.t182 239.927
R14538 Iout.n271 Iout.t243 239.927
R14539 Iout.n180 Iout.t245 239.927
R14540 Iout.n283 Iout.t114 239.927
R14541 Iout.n174 Iout.t76 239.927
R14542 Iout.n168 Iout.t80 239.927
R14543 Iout.n301 Iout.t2 239.927
R14544 Iout.n289 Iout.t226 239.927
R14545 Iout.n177 Iout.t255 239.927
R14546 Iout.n277 Iout.t179 239.927
R14547 Iout.n183 Iout.t5 239.927
R14548 Iout.n265 Iout.t210 239.927
R14549 Iout.n189 Iout.t248 239.927
R14550 Iout.n472 Iout.t19 239.927
R14551 Iout.n469 Iout.t74 239.927
R14552 Iout.n156 Iout.t108 239.927
R14553 Iout.n531 Iout.t125 239.927
R14554 Iout.n534 Iout.t69 239.927
R14555 Iout.n536 Iout.t58 239.927
R14556 Iout.n133 Iout.t220 239.927
R14557 Iout.n136 Iout.t55 239.927
R14558 Iout.n542 Iout.t16 239.927
R14559 Iout.n460 Iout.t136 239.927
R14560 Iout.n463 Iout.t173 239.927
R14561 Iout.n458 Iout.t73 239.927
R14562 Iout.n305 Iout.t183 239.927
R14563 Iout.n308 Iout.t194 239.927
R14564 Iout.n311 Iout.t18 239.927
R14565 Iout.n314 Iout.t165 239.927
R14566 Iout.n317 Iout.t191 239.927
R14567 Iout.n320 Iout.t176 239.927
R14568 Iout.n392 Iout.t30 239.927
R14569 Iout.n378 Iout.t237 239.927
R14570 Iout.n376 Iout.t25 239.927
R14571 Iout.n394 Iout.t7 239.927
R14572 Iout.n408 Iout.t14 239.927
R14573 Iout.n410 Iout.t154 239.927
R14574 Iout.n424 Iout.t185 239.927
R14575 Iout.n426 Iout.t207 239.927
R14576 Iout.n447 Iout.t190 239.927
R14577 Iout.n452 Iout.t152 239.927
R14578 Iout.n449 Iout.t45 239.927
R14579 Iout.n548 Iout.t89 239.927
R14580 Iout.n130 Iout.t232 239.927
R14581 Iout.n559 Iout.t49 239.927
R14582 Iout.n557 Iout.t166 239.927
R14583 Iout.n554 Iout.t184 239.927
R14584 Iout.n434 Iout.t112 239.927
R14585 Iout.n438 Iout.t247 239.927
R14586 Iout.n441 Iout.t126 239.927
R14587 Iout.n432 Iout.t15 239.927
R14588 Iout.n418 Iout.t111 239.927
R14589 Iout.n416 Iout.t206 239.927
R14590 Iout.n402 Iout.t6 239.927
R14591 Iout.n357 Iout.t204 239.927
R14592 Iout.n360 Iout.t212 239.927
R14593 Iout.n363 Iout.t102 239.927
R14594 Iout.n366 Iout.t81 239.927
R14595 Iout.n354 Iout.t222 239.927
R14596 Iout.n351 Iout.t96 239.927
R14597 Iout.n348 Iout.t107 239.927
R14598 Iout.n345 Iout.t40 239.927
R14599 Iout.n342 Iout.t115 239.927
R14600 Iout.n339 Iout.t28 239.927
R14601 Iout.n336 Iout.t83 239.927
R14602 Iout.n333 Iout.t180 239.927
R14603 Iout.n117 Iout.t34 239.927
R14604 Iout.n582 Iout.t169 239.927
R14605 Iout.n111 Iout.t84 239.927
R14606 Iout.n594 Iout.t219 239.927
R14607 Iout.n105 Iout.t138 239.927
R14608 Iout.n606 Iout.t99 239.927
R14609 Iout.n99 Iout.t48 239.927
R14610 Iout.n618 Iout.t177 239.927
R14611 Iout.n624 Iout.t17 239.927
R14612 Iout.n90 Iout.t52 239.927
R14613 Iout.n636 Iout.t29 239.927
R14614 Iout.n81 Iout.t187 239.927
R14615 Iout.n648 Iout.t164 239.927
R14616 Iout.n96 Iout.t238 239.927
R14617 Iout.n612 Iout.t11 239.927
R14618 Iout.n102 Iout.t188 239.927
R14619 Iout.n600 Iout.t32 239.927
R14620 Iout.n108 Iout.t239 239.927
R14621 Iout.n588 Iout.t66 239.927
R14622 Iout.n687 Iout.t151 239.927
R14623 Iout.n684 Iout.t225 239.927
R14624 Iout.n681 Iout.t85 239.927
R14625 Iout.n678 Iout.t156 239.927
R14626 Iout.n675 Iout.t56 239.927
R14627 Iout.n672 Iout.t224 239.927
R14628 Iout.n747 Iout.t130 239.927
R14629 Iout.n50 Iout.t218 239.927
R14630 Iout.n759 Iout.t106 239.927
R14631 Iout.n44 Iout.t67 239.927
R14632 Iout.n771 Iout.t41 239.927
R14633 Iout.n42 Iout.t244 239.927
R14634 Iout.n56 Iout.t159 239.927
R14635 Iout.n735 Iout.t202 239.927
R14636 Iout.n62 Iout.t198 239.927
R14637 Iout.n723 Iout.t242 239.927
R14638 Iout.n717 Iout.t46 239.927
R14639 Iout.n65 Iout.t65 239.927
R14640 Iout.n729 Iout.t231 239.927
R14641 Iout.n59 Iout.t170 239.927
R14642 Iout.n805 Iout.t122 239.927
R14643 Iout.n808 Iout.t189 239.927
R14644 Iout.n811 Iout.t228 239.927
R14645 Iout.n814 Iout.t47 239.927
R14646 Iout.n817 Iout.t92 239.927
R14647 Iout.n820 Iout.t252 239.927
R14648 Iout.n823 Iout.t233 239.927
R14649 Iout.n802 Iout.t230 239.927
R14650 Iout.n799 Iout.t131 239.927
R14651 Iout.n890 Iout.t94 239.927
R14652 Iout.n888 Iout.t60 239.927
R14653 Iout.n881 Iout.t82 239.927
R14654 Iout.n869 Iout.t253 239.927
R14655 Iout.n867 Iout.t146 239.927
R14656 Iout.n855 Iout.t43 239.927
R14657 Iout.n853 Iout.t87 239.927
R14658 Iout.n841 Iout.t158 239.927
R14659 Iout.n839 Iout.t254 239.927
R14660 Iout.n827 Iout.t163 239.927
R14661 Iout.n883 Iout.t68 239.927
R14662 Iout.n895 Iout.t150 239.927
R14663 Iout.n897 Iout.t246 239.927
R14664 Iout.n909 Iout.t120 239.927
R14665 Iout.n911 Iout.t251 239.927
R14666 Iout.n923 Iout.t0 239.927
R14667 Iout.n926 Iout.t90 239.927
R14668 Iout.n22 Iout.t57 239.927
R14669 Iout.n876 Iout.t175 239.927
R14670 Iout.n874 Iout.t241 239.927
R14671 Iout.n862 Iout.t119 239.927
R14672 Iout.n860 Iout.t149 239.927
R14673 Iout.n848 Iout.t217 239.927
R14674 Iout.n846 Iout.t70 239.927
R14675 Iout.n834 Iout.t141 239.927
R14676 Iout.n832 Iout.t116 239.927
R14677 Iout.n902 Iout.t38 239.927
R14678 Iout.n904 Iout.t127 239.927
R14679 Iout.n916 Iout.t215 239.927
R14680 Iout.n918 Iout.t209 239.927
R14681 Iout.n931 Iout.t4 239.927
R14682 Iout.n934 Iout.t1 239.927
R14683 Iout.n796 Iout.t174 239.927
R14684 Iout.n793 Iout.t22 239.927
R14685 Iout.n790 Iout.t27 239.927
R14686 Iout.n787 Iout.t197 239.927
R14687 Iout.n784 Iout.t147 239.927
R14688 Iout.n781 Iout.t53 239.927
R14689 Iout.n938 Iout.t221 239.927
R14690 Iout.n741 Iout.t137 239.927
R14691 Iout.n53 Iout.t123 239.927
R14692 Iout.n753 Iout.t88 239.927
R14693 Iout.n47 Iout.t199 239.927
R14694 Iout.n765 Iout.t100 239.927
R14695 Iout.n38 Iout.t103 239.927
R14696 Iout.n777 Iout.t51 239.927
R14697 Iout.n71 Iout.t211 239.927
R14698 Iout.n705 Iout.t23 239.927
R14699 Iout.n77 Iout.t132 239.927
R14700 Iout.n944 Iout.t155 239.927
R14701 Iout.n19 Iout.t50 239.927
R14702 Iout.n68 Iout.t37 239.927
R14703 Iout.n711 Iout.t98 239.927
R14704 Iout.n74 Iout.t105 239.927
R14705 Iout.n699 Iout.t101 239.927
R14706 Iout.n950 Iout.t196 239.927
R14707 Iout.n953 Iout.t227 239.927
R14708 Iout.n669 Iout.t104 239.927
R14709 Iout.n666 Iout.t71 239.927
R14710 Iout.n663 Iout.t12 239.927
R14711 Iout.n660 Iout.t109 239.927
R14712 Iout.n657 Iout.t208 239.927
R14713 Iout.n654 Iout.t235 239.927
R14714 Iout.n690 Iout.t229 239.927
R14715 Iout.n695 Iout.t59 239.927
R14716 Iout.n692 Iout.t193 239.927
R14717 Iout.n957 Iout.t36 239.927
R14718 Iout.n114 Iout.t161 239.927
R14719 Iout.n576 Iout.t167 239.927
R14720 Iout.n573 Iout.t162 239.927
R14721 Iout.n963 Iout.t142 239.927
R14722 Iout.n14 Iout.t157 239.927
R14723 Iout.n93 Iout.t79 239.927
R14724 Iout.n630 Iout.t129 239.927
R14725 Iout.n87 Iout.t192 239.927
R14726 Iout.n642 Iout.t144 239.927
R14727 Iout.n85 Iout.t77 239.927
R14728 Iout.n563 Iout.t44 239.927
R14729 Iout.n969 Iout.t10 239.927
R14730 Iout.n972 Iout.t172 239.927
R14731 Iout.n569 Iout.t24 239.927
R14732 Iout.n123 Iout.t148 239.927
R14733 Iout.n120 Iout.t240 239.927
R14734 Iout.n976 Iout.t201 239.927
R14735 Iout.n400 Iout.t140 239.927
R14736 Iout.n386 Iout.t113 239.927
R14737 Iout.n384 Iout.t97 239.927
R14738 Iout.n370 Iout.t223 239.927
R14739 Iout.n982 Iout.t195 239.927
R14740 Iout.n9 Iout.t31 239.927
R14741 Iout.n127 Iout.t78 239.927
R14742 Iout.n988 Iout.t250 239.927
R14743 Iout.n991 Iout.t8 239.927
R14744 Iout.n323 Iout.t186 239.927
R14745 Iout.n326 Iout.t171 239.927
R14746 Iout.n329 Iout.t128 239.927
R14747 Iout.n995 Iout.t236 239.927
R14748 Iout.n1001 Iout.t213 239.927
R14749 Iout.n4 Iout.t21 239.927
R14750 Iout.n295 Iout.t181 239.927
R14751 Iout.n172 Iout.t134 239.927
R14752 Iout.n1014 Iout.t54 239.927
R14753 Iout.n1021 Iout.n1020 7.9105
R14754 Iout.n510 Iout.n509 7.9105
R14755 Iout.n514 Iout.n513 7.9105
R14756 Iout.n508 Iout.n507 7.9105
R14757 Iout.n505 Iout.n504 7.9105
R14758 Iout.n501 Iout.n500 7.9105
R14759 Iout.n193 Iout.n192 7.9105
R14760 Iout.n196 Iout.n195 7.9105
R14761 Iout.n200 Iout.n199 7.9105
R14762 Iout.n203 Iout.n202 7.9105
R14763 Iout.n207 Iout.n206 7.9105
R14764 Iout.n211 Iout.n210 7.9105
R14765 Iout.n215 Iout.n214 7.9105
R14766 Iout.n219 Iout.n218 7.9105
R14767 Iout.n223 Iout.n222 7.9105
R14768 Iout.n227 Iout.n226 7.9105
R14769 Iout.n233 Iout.n232 7.9105
R14770 Iout.n236 Iout.n235 7.9105
R14771 Iout.n239 Iout.n238 7.9105
R14772 Iout.n242 Iout.n241 7.9105
R14773 Iout.n245 Iout.n244 7.9105
R14774 Iout.n248 Iout.n247 7.9105
R14775 Iout.n251 Iout.n250 7.9105
R14776 Iout.n256 Iout.n255 7.9105
R14777 Iout.n253 Iout.n252 7.9105
R14778 Iout.n490 Iout.n489 7.9105
R14779 Iout.n495 Iout.n494 7.9105
R14780 Iout.n492 Iout.n491 7.9105
R14781 Iout.n520 Iout.n519 7.9105
R14782 Iout.n150 Iout.n149 7.9105
R14783 Iout.n147 Iout.n146 7.9105
R14784 Iout.n1011 Iout.n1010 7.9105
R14785 Iout.n1008 Iout.n1007 7.9105
R14786 Iout.n141 Iout.n140 7.9105
R14787 Iout.n144 Iout.n143 7.9105
R14788 Iout.n526 Iout.n525 7.9105
R14789 Iout.n481 Iout.n480 7.9105
R14790 Iout.n484 Iout.n483 7.9105
R14791 Iout.n479 Iout.n478 7.9105
R14792 Iout.n260 Iout.n259 7.9105
R14793 Iout.n187 Iout.n186 7.9105
R14794 Iout.n272 Iout.n271 7.9105
R14795 Iout.n181 Iout.n180 7.9105
R14796 Iout.n284 Iout.n283 7.9105
R14797 Iout.n175 Iout.n174 7.9105
R14798 Iout.n169 Iout.n168 7.9105
R14799 Iout.n302 Iout.n301 7.9105
R14800 Iout.n290 Iout.n289 7.9105
R14801 Iout.n178 Iout.n177 7.9105
R14802 Iout.n278 Iout.n277 7.9105
R14803 Iout.n184 Iout.n183 7.9105
R14804 Iout.n266 Iout.n265 7.9105
R14805 Iout.n190 Iout.n189 7.9105
R14806 Iout.n473 Iout.n472 7.9105
R14807 Iout.n470 Iout.n469 7.9105
R14808 Iout.n157 Iout.n156 7.9105
R14809 Iout.n532 Iout.n531 7.9105
R14810 Iout.n535 Iout.n534 7.9105
R14811 Iout.n537 Iout.n536 7.9105
R14812 Iout.n134 Iout.n133 7.9105
R14813 Iout.n137 Iout.n136 7.9105
R14814 Iout.n543 Iout.n542 7.9105
R14815 Iout.n461 Iout.n460 7.9105
R14816 Iout.n464 Iout.n463 7.9105
R14817 Iout.n459 Iout.n458 7.9105
R14818 Iout.n306 Iout.n305 7.9105
R14819 Iout.n309 Iout.n308 7.9105
R14820 Iout.n312 Iout.n311 7.9105
R14821 Iout.n315 Iout.n314 7.9105
R14822 Iout.n318 Iout.n317 7.9105
R14823 Iout.n321 Iout.n320 7.9105
R14824 Iout.n393 Iout.n392 7.9105
R14825 Iout.n379 Iout.n378 7.9105
R14826 Iout.n377 Iout.n376 7.9105
R14827 Iout.n395 Iout.n394 7.9105
R14828 Iout.n409 Iout.n408 7.9105
R14829 Iout.n411 Iout.n410 7.9105
R14830 Iout.n425 Iout.n424 7.9105
R14831 Iout.n427 Iout.n426 7.9105
R14832 Iout.n448 Iout.n447 7.9105
R14833 Iout.n453 Iout.n452 7.9105
R14834 Iout.n450 Iout.n449 7.9105
R14835 Iout.n549 Iout.n548 7.9105
R14836 Iout.n131 Iout.n130 7.9105
R14837 Iout.n560 Iout.n559 7.9105
R14838 Iout.n558 Iout.n557 7.9105
R14839 Iout.n555 Iout.n554 7.9105
R14840 Iout.n435 Iout.n434 7.9105
R14841 Iout.n439 Iout.n438 7.9105
R14842 Iout.n442 Iout.n441 7.9105
R14843 Iout.n433 Iout.n432 7.9105
R14844 Iout.n419 Iout.n418 7.9105
R14845 Iout.n417 Iout.n416 7.9105
R14846 Iout.n403 Iout.n402 7.9105
R14847 Iout.n358 Iout.n357 7.9105
R14848 Iout.n361 Iout.n360 7.9105
R14849 Iout.n364 Iout.n363 7.9105
R14850 Iout.n367 Iout.n366 7.9105
R14851 Iout.n355 Iout.n354 7.9105
R14852 Iout.n352 Iout.n351 7.9105
R14853 Iout.n349 Iout.n348 7.9105
R14854 Iout.n346 Iout.n345 7.9105
R14855 Iout.n343 Iout.n342 7.9105
R14856 Iout.n340 Iout.n339 7.9105
R14857 Iout.n337 Iout.n336 7.9105
R14858 Iout.n334 Iout.n333 7.9105
R14859 Iout.n118 Iout.n117 7.9105
R14860 Iout.n583 Iout.n582 7.9105
R14861 Iout.n112 Iout.n111 7.9105
R14862 Iout.n595 Iout.n594 7.9105
R14863 Iout.n106 Iout.n105 7.9105
R14864 Iout.n607 Iout.n606 7.9105
R14865 Iout.n100 Iout.n99 7.9105
R14866 Iout.n619 Iout.n618 7.9105
R14867 Iout.n625 Iout.n624 7.9105
R14868 Iout.n91 Iout.n90 7.9105
R14869 Iout.n637 Iout.n636 7.9105
R14870 Iout.n82 Iout.n81 7.9105
R14871 Iout.n649 Iout.n648 7.9105
R14872 Iout.n97 Iout.n96 7.9105
R14873 Iout.n613 Iout.n612 7.9105
R14874 Iout.n103 Iout.n102 7.9105
R14875 Iout.n601 Iout.n600 7.9105
R14876 Iout.n109 Iout.n108 7.9105
R14877 Iout.n589 Iout.n588 7.9105
R14878 Iout.n688 Iout.n687 7.9105
R14879 Iout.n685 Iout.n684 7.9105
R14880 Iout.n682 Iout.n681 7.9105
R14881 Iout.n679 Iout.n678 7.9105
R14882 Iout.n676 Iout.n675 7.9105
R14883 Iout.n673 Iout.n672 7.9105
R14884 Iout.n748 Iout.n747 7.9105
R14885 Iout.n51 Iout.n50 7.9105
R14886 Iout.n760 Iout.n759 7.9105
R14887 Iout.n45 Iout.n44 7.9105
R14888 Iout.n772 Iout.n771 7.9105
R14889 Iout.n43 Iout.n42 7.9105
R14890 Iout.n57 Iout.n56 7.9105
R14891 Iout.n736 Iout.n735 7.9105
R14892 Iout.n63 Iout.n62 7.9105
R14893 Iout.n724 Iout.n723 7.9105
R14894 Iout.n718 Iout.n717 7.9105
R14895 Iout.n66 Iout.n65 7.9105
R14896 Iout.n730 Iout.n729 7.9105
R14897 Iout.n60 Iout.n59 7.9105
R14898 Iout.n806 Iout.n805 7.9105
R14899 Iout.n809 Iout.n808 7.9105
R14900 Iout.n812 Iout.n811 7.9105
R14901 Iout.n815 Iout.n814 7.9105
R14902 Iout.n818 Iout.n817 7.9105
R14903 Iout.n821 Iout.n820 7.9105
R14904 Iout.n824 Iout.n823 7.9105
R14905 Iout.n803 Iout.n802 7.9105
R14906 Iout.n800 Iout.n799 7.9105
R14907 Iout.n891 Iout.n890 7.9105
R14908 Iout.n889 Iout.n888 7.9105
R14909 Iout.n882 Iout.n881 7.9105
R14910 Iout.n870 Iout.n869 7.9105
R14911 Iout.n868 Iout.n867 7.9105
R14912 Iout.n856 Iout.n855 7.9105
R14913 Iout.n854 Iout.n853 7.9105
R14914 Iout.n842 Iout.n841 7.9105
R14915 Iout.n840 Iout.n839 7.9105
R14916 Iout.n828 Iout.n827 7.9105
R14917 Iout.n884 Iout.n883 7.9105
R14918 Iout.n896 Iout.n895 7.9105
R14919 Iout.n898 Iout.n897 7.9105
R14920 Iout.n910 Iout.n909 7.9105
R14921 Iout.n912 Iout.n911 7.9105
R14922 Iout.n924 Iout.n923 7.9105
R14923 Iout.n927 Iout.n926 7.9105
R14924 Iout.n23 Iout.n22 7.9105
R14925 Iout.n877 Iout.n876 7.9105
R14926 Iout.n875 Iout.n874 7.9105
R14927 Iout.n863 Iout.n862 7.9105
R14928 Iout.n861 Iout.n860 7.9105
R14929 Iout.n849 Iout.n848 7.9105
R14930 Iout.n847 Iout.n846 7.9105
R14931 Iout.n835 Iout.n834 7.9105
R14932 Iout.n833 Iout.n832 7.9105
R14933 Iout.n903 Iout.n902 7.9105
R14934 Iout.n905 Iout.n904 7.9105
R14935 Iout.n917 Iout.n916 7.9105
R14936 Iout.n919 Iout.n918 7.9105
R14937 Iout.n932 Iout.n931 7.9105
R14938 Iout.n935 Iout.n934 7.9105
R14939 Iout.n797 Iout.n796 7.9105
R14940 Iout.n794 Iout.n793 7.9105
R14941 Iout.n791 Iout.n790 7.9105
R14942 Iout.n788 Iout.n787 7.9105
R14943 Iout.n785 Iout.n784 7.9105
R14944 Iout.n782 Iout.n781 7.9105
R14945 Iout.n939 Iout.n938 7.9105
R14946 Iout.n742 Iout.n741 7.9105
R14947 Iout.n54 Iout.n53 7.9105
R14948 Iout.n754 Iout.n753 7.9105
R14949 Iout.n48 Iout.n47 7.9105
R14950 Iout.n766 Iout.n765 7.9105
R14951 Iout.n39 Iout.n38 7.9105
R14952 Iout.n778 Iout.n777 7.9105
R14953 Iout.n72 Iout.n71 7.9105
R14954 Iout.n706 Iout.n705 7.9105
R14955 Iout.n78 Iout.n77 7.9105
R14956 Iout.n945 Iout.n944 7.9105
R14957 Iout.n20 Iout.n19 7.9105
R14958 Iout.n69 Iout.n68 7.9105
R14959 Iout.n712 Iout.n711 7.9105
R14960 Iout.n75 Iout.n74 7.9105
R14961 Iout.n700 Iout.n699 7.9105
R14962 Iout.n951 Iout.n950 7.9105
R14963 Iout.n954 Iout.n953 7.9105
R14964 Iout.n670 Iout.n669 7.9105
R14965 Iout.n667 Iout.n666 7.9105
R14966 Iout.n664 Iout.n663 7.9105
R14967 Iout.n661 Iout.n660 7.9105
R14968 Iout.n658 Iout.n657 7.9105
R14969 Iout.n655 Iout.n654 7.9105
R14970 Iout.n691 Iout.n690 7.9105
R14971 Iout.n696 Iout.n695 7.9105
R14972 Iout.n693 Iout.n692 7.9105
R14973 Iout.n958 Iout.n957 7.9105
R14974 Iout.n115 Iout.n114 7.9105
R14975 Iout.n577 Iout.n576 7.9105
R14976 Iout.n574 Iout.n573 7.9105
R14977 Iout.n964 Iout.n963 7.9105
R14978 Iout.n15 Iout.n14 7.9105
R14979 Iout.n94 Iout.n93 7.9105
R14980 Iout.n631 Iout.n630 7.9105
R14981 Iout.n88 Iout.n87 7.9105
R14982 Iout.n643 Iout.n642 7.9105
R14983 Iout.n86 Iout.n85 7.9105
R14984 Iout.n564 Iout.n563 7.9105
R14985 Iout.n970 Iout.n969 7.9105
R14986 Iout.n973 Iout.n972 7.9105
R14987 Iout.n570 Iout.n569 7.9105
R14988 Iout.n124 Iout.n123 7.9105
R14989 Iout.n121 Iout.n120 7.9105
R14990 Iout.n977 Iout.n976 7.9105
R14991 Iout.n401 Iout.n400 7.9105
R14992 Iout.n387 Iout.n386 7.9105
R14993 Iout.n385 Iout.n384 7.9105
R14994 Iout.n371 Iout.n370 7.9105
R14995 Iout.n983 Iout.n982 7.9105
R14996 Iout.n10 Iout.n9 7.9105
R14997 Iout.n128 Iout.n127 7.9105
R14998 Iout.n989 Iout.n988 7.9105
R14999 Iout.n992 Iout.n991 7.9105
R15000 Iout.n324 Iout.n323 7.9105
R15001 Iout.n327 Iout.n326 7.9105
R15002 Iout.n330 Iout.n329 7.9105
R15003 Iout.n996 Iout.n995 7.9105
R15004 Iout.n1002 Iout.n1001 7.9105
R15005 Iout.n5 Iout.n4 7.9105
R15006 Iout.n296 Iout.n295 7.9105
R15007 Iout.n173 Iout.n172 7.9105
R15008 Iout.n1015 Iout.n1014 7.9105
R15009 Iout.n886 Iout.n885 3.86101
R15010 Iout.n880 Iout.n879 3.86101
R15011 Iout.n894 Iout.n893 3.86101
R15012 Iout.n872 Iout.n871 3.86101
R15013 Iout.n900 Iout.n899 3.86101
R15014 Iout.n866 Iout.n865 3.86101
R15015 Iout.n908 Iout.n907 3.86101
R15016 Iout.n858 Iout.n857 3.86101
R15017 Iout.n914 Iout.n913 3.86101
R15018 Iout.n852 Iout.n851 3.86101
R15019 Iout.n922 Iout.n921 3.86101
R15020 Iout.n844 Iout.n843 3.86101
R15021 Iout.n929 Iout.n928 3.86101
R15022 Iout.n838 Iout.n837 3.86101
R15023 Iout.n925 Iout.n21 3.86101
R15024 Iout.n830 Iout.n829 3.86101
R15025 Iout.n879 Iout.n878 3.4105
R15026 Iout.n887 Iout.n886 3.4105
R15027 Iout.n893 Iout.n892 3.4105
R15028 Iout.n798 Iout.n28 3.4105
R15029 Iout.n801 Iout.n29 3.4105
R15030 Iout.n804 Iout.n30 3.4105
R15031 Iout.n807 Iout.n31 3.4105
R15032 Iout.n873 Iout.n872 3.4105
R15033 Iout.n744 Iout.n743 3.4105
R15034 Iout.n740 Iout.n739 3.4105
R15035 Iout.n732 Iout.n731 3.4105
R15036 Iout.n728 Iout.n727 3.4105
R15037 Iout.n720 Iout.n719 3.4105
R15038 Iout.n795 Iout.n27 3.4105
R15039 Iout.n901 Iout.n900 3.4105
R15040 Iout.n722 Iout.n721 3.4105
R15041 Iout.n726 Iout.n725 3.4105
R15042 Iout.n734 Iout.n733 3.4105
R15043 Iout.n738 Iout.n737 3.4105
R15044 Iout.n746 Iout.n745 3.4105
R15045 Iout.n750 Iout.n749 3.4105
R15046 Iout.n752 Iout.n751 3.4105
R15047 Iout.n810 Iout.n32 3.4105
R15048 Iout.n865 Iout.n864 3.4105
R15049 Iout.n668 Iout.n55 3.4105
R15050 Iout.n671 Iout.n58 3.4105
R15051 Iout.n674 Iout.n61 3.4105
R15052 Iout.n677 Iout.n64 3.4105
R15053 Iout.n680 Iout.n67 3.4105
R15054 Iout.n683 Iout.n70 3.4105
R15055 Iout.n686 Iout.n73 3.4105
R15056 Iout.n714 Iout.n713 3.4105
R15057 Iout.n716 Iout.n715 3.4105
R15058 Iout.n792 Iout.n26 3.4105
R15059 Iout.n907 Iout.n906 3.4105
R15060 Iout.n587 Iout.n586 3.4105
R15061 Iout.n591 Iout.n590 3.4105
R15062 Iout.n599 Iout.n598 3.4105
R15063 Iout.n603 Iout.n602 3.4105
R15064 Iout.n611 Iout.n610 3.4105
R15065 Iout.n615 Iout.n614 3.4105
R15066 Iout.n623 Iout.n622 3.4105
R15067 Iout.n627 Iout.n626 3.4105
R15068 Iout.n665 Iout.n52 3.4105
R15069 Iout.n758 Iout.n757 3.4105
R15070 Iout.n756 Iout.n755 3.4105
R15071 Iout.n813 Iout.n33 3.4105
R15072 Iout.n859 Iout.n858 3.4105
R15073 Iout.n629 Iout.n628 3.4105
R15074 Iout.n621 Iout.n620 3.4105
R15075 Iout.n617 Iout.n616 3.4105
R15076 Iout.n609 Iout.n608 3.4105
R15077 Iout.n605 Iout.n604 3.4105
R15078 Iout.n597 Iout.n596 3.4105
R15079 Iout.n593 Iout.n592 3.4105
R15080 Iout.n585 Iout.n584 3.4105
R15081 Iout.n581 Iout.n580 3.4105
R15082 Iout.n579 Iout.n578 3.4105
R15083 Iout.n689 Iout.n76 3.4105
R15084 Iout.n710 Iout.n709 3.4105
R15085 Iout.n708 Iout.n707 3.4105
R15086 Iout.n789 Iout.n25 3.4105
R15087 Iout.n915 Iout.n914 3.4105
R15088 Iout.n572 Iout.n571 3.4105
R15089 Iout.n335 Iout.n116 3.4105
R15090 Iout.n338 Iout.n113 3.4105
R15091 Iout.n341 Iout.n110 3.4105
R15092 Iout.n344 Iout.n107 3.4105
R15093 Iout.n347 Iout.n104 3.4105
R15094 Iout.n350 Iout.n101 3.4105
R15095 Iout.n353 Iout.n98 3.4105
R15096 Iout.n356 Iout.n95 3.4105
R15097 Iout.n359 Iout.n92 3.4105
R15098 Iout.n633 Iout.n632 3.4105
R15099 Iout.n635 Iout.n634 3.4105
R15100 Iout.n662 Iout.n49 3.4105
R15101 Iout.n762 Iout.n761 3.4105
R15102 Iout.n764 Iout.n763 3.4105
R15103 Iout.n816 Iout.n34 3.4105
R15104 Iout.n851 Iout.n850 3.4105
R15105 Iout.n399 Iout.n398 3.4105
R15106 Iout.n405 Iout.n404 3.4105
R15107 Iout.n415 Iout.n414 3.4105
R15108 Iout.n421 Iout.n420 3.4105
R15109 Iout.n431 Iout.n430 3.4105
R15110 Iout.n444 Iout.n443 3.4105
R15111 Iout.n440 Iout.n159 3.4105
R15112 Iout.n437 Iout.n436 3.4105
R15113 Iout.n553 Iout.n552 3.4105
R15114 Iout.n556 Iout.n119 3.4105
R15115 Iout.n562 Iout.n561 3.4105
R15116 Iout.n568 Iout.n567 3.4105
R15117 Iout.n566 Iout.n565 3.4105
R15118 Iout.n575 Iout.n79 3.4105
R15119 Iout.n698 Iout.n697 3.4105
R15120 Iout.n702 Iout.n701 3.4105
R15121 Iout.n704 Iout.n703 3.4105
R15122 Iout.n786 Iout.n24 3.4105
R15123 Iout.n921 Iout.n920 3.4105
R15124 Iout.n129 Iout.n125 3.4105
R15125 Iout.n547 Iout.n546 3.4105
R15126 Iout.n551 Iout.n550 3.4105
R15127 Iout.n451 Iout.n158 3.4105
R15128 Iout.n455 Iout.n454 3.4105
R15129 Iout.n446 Iout.n445 3.4105
R15130 Iout.n429 Iout.n428 3.4105
R15131 Iout.n423 Iout.n422 3.4105
R15132 Iout.n413 Iout.n412 3.4105
R15133 Iout.n407 Iout.n406 3.4105
R15134 Iout.n397 Iout.n396 3.4105
R15135 Iout.n391 Iout.n390 3.4105
R15136 Iout.n389 Iout.n388 3.4105
R15137 Iout.n362 Iout.n89 3.4105
R15138 Iout.n641 Iout.n640 3.4105
R15139 Iout.n639 Iout.n638 3.4105
R15140 Iout.n659 Iout.n46 3.4105
R15141 Iout.n770 Iout.n769 3.4105
R15142 Iout.n768 Iout.n767 3.4105
R15143 Iout.n819 Iout.n35 3.4105
R15144 Iout.n845 Iout.n844 3.4105
R15145 Iout.n325 Iout.n165 3.4105
R15146 Iout.n322 Iout.n164 3.4105
R15147 Iout.n319 Iout.n163 3.4105
R15148 Iout.n316 Iout.n162 3.4105
R15149 Iout.n313 Iout.n161 3.4105
R15150 Iout.n310 Iout.n160 3.4105
R15151 Iout.n307 Iout.n155 3.4105
R15152 Iout.n457 Iout.n456 3.4105
R15153 Iout.n466 Iout.n465 3.4105
R15154 Iout.n462 Iout.n126 3.4105
R15155 Iout.n545 Iout.n544 3.4105
R15156 Iout.n541 Iout.n540 3.4105
R15157 Iout.n135 Iout.n3 3.4105
R15158 Iout.n987 Iout.n986 3.4105
R15159 Iout.n985 Iout.n984 3.4105
R15160 Iout.n122 Iout.n8 3.4105
R15161 Iout.n968 Iout.n967 3.4105
R15162 Iout.n966 Iout.n965 3.4105
R15163 Iout.n694 Iout.n13 3.4105
R15164 Iout.n949 Iout.n948 3.4105
R15165 Iout.n947 Iout.n946 3.4105
R15166 Iout.n783 Iout.n18 3.4105
R15167 Iout.n930 Iout.n929 3.4105
R15168 Iout.n1004 Iout.n1003 3.4105
R15169 Iout.n539 Iout.n538 3.4105
R15170 Iout.n533 Iout.n132 3.4105
R15171 Iout.n530 Iout.n529 3.4105
R15172 Iout.n468 Iout.n467 3.4105
R15173 Iout.n471 Iout.n153 3.4105
R15174 Iout.n475 Iout.n474 3.4105
R15175 Iout.n264 Iout.n263 3.4105
R15176 Iout.n268 Iout.n267 3.4105
R15177 Iout.n276 Iout.n275 3.4105
R15178 Iout.n280 Iout.n279 3.4105
R15179 Iout.n288 Iout.n287 3.4105
R15180 Iout.n292 Iout.n291 3.4105
R15181 Iout.n300 Iout.n299 3.4105
R15182 Iout.n328 Iout.n166 3.4105
R15183 Iout.n381 Iout.n380 3.4105
R15184 Iout.n383 Iout.n382 3.4105
R15185 Iout.n365 Iout.n83 3.4105
R15186 Iout.n645 Iout.n644 3.4105
R15187 Iout.n647 Iout.n646 3.4105
R15188 Iout.n656 Iout.n40 3.4105
R15189 Iout.n774 Iout.n773 3.4105
R15190 Iout.n776 Iout.n775 3.4105
R15191 Iout.n822 Iout.n36 3.4105
R15192 Iout.n837 Iout.n836 3.4105
R15193 Iout.n298 Iout.n297 3.4105
R15194 Iout.n294 Iout.n293 3.4105
R15195 Iout.n286 Iout.n285 3.4105
R15196 Iout.n282 Iout.n281 3.4105
R15197 Iout.n274 Iout.n273 3.4105
R15198 Iout.n270 Iout.n269 3.4105
R15199 Iout.n262 Iout.n261 3.4105
R15200 Iout.n477 Iout.n476 3.4105
R15201 Iout.n486 Iout.n485 3.4105
R15202 Iout.n482 Iout.n151 3.4105
R15203 Iout.n528 Iout.n527 3.4105
R15204 Iout.n524 Iout.n523 3.4105
R15205 Iout.n142 Iout.n138 3.4105
R15206 Iout.n1006 Iout.n1005 3.4105
R15207 Iout.n1009 Iout.n0 3.4105
R15208 Iout.n1000 Iout.n999 3.4105
R15209 Iout.n998 Iout.n997 3.4105
R15210 Iout.n990 Iout.n6 3.4105
R15211 Iout.n981 Iout.n980 3.4105
R15212 Iout.n979 Iout.n978 3.4105
R15213 Iout.n971 Iout.n11 3.4105
R15214 Iout.n962 Iout.n961 3.4105
R15215 Iout.n960 Iout.n959 3.4105
R15216 Iout.n952 Iout.n16 3.4105
R15217 Iout.n943 Iout.n942 3.4105
R15218 Iout.n941 Iout.n940 3.4105
R15219 Iout.n933 Iout.n21 3.4105
R15220 Iout.n1017 Iout.n1016 3.4105
R15221 Iout.n148 Iout.n2 3.4105
R15222 Iout.n518 Iout.n517 3.4105
R15223 Iout.n522 Iout.n521 3.4105
R15224 Iout.n493 Iout.n139 3.4105
R15225 Iout.n497 Iout.n496 3.4105
R15226 Iout.n488 Iout.n487 3.4105
R15227 Iout.n254 Iout.n154 3.4105
R15228 Iout.n258 Iout.n257 3.4105
R15229 Iout.n249 Iout.n188 3.4105
R15230 Iout.n246 Iout.n185 3.4105
R15231 Iout.n243 Iout.n182 3.4105
R15232 Iout.n240 Iout.n179 3.4105
R15233 Iout.n237 Iout.n176 3.4105
R15234 Iout.n234 Iout.n170 3.4105
R15235 Iout.n231 Iout.n230 3.4105
R15236 Iout.n171 Iout.n167 3.4105
R15237 Iout.n304 Iout.n303 3.4105
R15238 Iout.n332 Iout.n331 3.4105
R15239 Iout.n375 Iout.n374 3.4105
R15240 Iout.n373 Iout.n372 3.4105
R15241 Iout.n369 Iout.n368 3.4105
R15242 Iout.n84 Iout.n80 3.4105
R15243 Iout.n651 Iout.n650 3.4105
R15244 Iout.n653 Iout.n652 3.4105
R15245 Iout.n41 Iout.n37 3.4105
R15246 Iout.n780 Iout.n779 3.4105
R15247 Iout.n826 Iout.n825 3.4105
R15248 Iout.n831 Iout.n830 3.4105
R15249 Iout.n229 Iout.n228 3.4105
R15250 Iout.n225 Iout.n224 3.4105
R15251 Iout.n221 Iout.n220 3.4105
R15252 Iout.n217 Iout.n216 3.4105
R15253 Iout.n213 Iout.n212 3.4105
R15254 Iout.n209 Iout.n208 3.4105
R15255 Iout.n205 Iout.n204 3.4105
R15256 Iout.n201 Iout.n191 3.4105
R15257 Iout.n198 Iout.n197 3.4105
R15258 Iout.n194 Iout.n152 3.4105
R15259 Iout.n499 Iout.n498 3.4105
R15260 Iout.n503 Iout.n502 3.4105
R15261 Iout.n506 Iout.n145 3.4105
R15262 Iout.n516 Iout.n515 3.4105
R15263 Iout.n512 Iout.n511 3.4105
R15264 Iout.n1019 Iout.n1018 3.4105
R15265 Iout.n936 Iout.n23 1.43848
R15266 Iout.n936 Iout.n935 1.34612
R15267 Iout.n939 Iout.n937 1.34612
R15268 Iout.n20 Iout.n17 1.34612
R15269 Iout.n955 Iout.n954 1.34612
R15270 Iout.n958 Iout.n956 1.34612
R15271 Iout.n15 Iout.n12 1.34612
R15272 Iout.n974 Iout.n973 1.34612
R15273 Iout.n977 Iout.n975 1.34612
R15274 Iout.n10 Iout.n7 1.34612
R15275 Iout.n993 Iout.n992 1.34612
R15276 Iout.n996 Iout.n994 1.34612
R15277 Iout.n5 Iout.n1 1.34612
R15278 Iout.n1012 Iout.n1011 1.34612
R15279 Iout.n1015 Iout.n1013 1.34612
R15280 Iout.n1022 Iout.n1021 1.34612
R15281 Iout.n197 Iout.n154 0.451012
R15282 Iout.n476 Iout.n154 0.451012
R15283 Iout.n476 Iout.n475 0.451012
R15284 Iout.n475 Iout.n155 0.451012
R15285 Iout.n445 Iout.n155 0.451012
R15286 Iout.n445 Iout.n444 0.451012
R15287 Iout.n444 Iout.n107 0.451012
R15288 Iout.n604 Iout.n107 0.451012
R15289 Iout.n604 Iout.n603 0.451012
R15290 Iout.n603 Iout.n64 0.451012
R15291 Iout.n733 Iout.n64 0.451012
R15292 Iout.n733 Iout.n732 0.451012
R15293 Iout.n732 Iout.n29 0.451012
R15294 Iout.n886 Iout.n29 0.451012
R15295 Iout.n258 Iout.n191 0.451012
R15296 Iout.n262 Iout.n258 0.451012
R15297 Iout.n263 Iout.n262 0.451012
R15298 Iout.n263 Iout.n160 0.451012
R15299 Iout.n429 Iout.n160 0.451012
R15300 Iout.n430 Iout.n429 0.451012
R15301 Iout.n430 Iout.n104 0.451012
R15302 Iout.n609 Iout.n104 0.451012
R15303 Iout.n610 Iout.n609 0.451012
R15304 Iout.n610 Iout.n61 0.451012
R15305 Iout.n738 Iout.n61 0.451012
R15306 Iout.n739 Iout.n738 0.451012
R15307 Iout.n739 Iout.n30 0.451012
R15308 Iout.n879 Iout.n30 0.451012
R15309 Iout.n487 Iout.n152 0.451012
R15310 Iout.n487 Iout.n486 0.451012
R15311 Iout.n486 Iout.n153 0.451012
R15312 Iout.n456 Iout.n153 0.451012
R15313 Iout.n456 Iout.n455 0.451012
R15314 Iout.n455 Iout.n159 0.451012
R15315 Iout.n159 Iout.n110 0.451012
R15316 Iout.n597 Iout.n110 0.451012
R15317 Iout.n598 Iout.n597 0.451012
R15318 Iout.n598 Iout.n67 0.451012
R15319 Iout.n726 Iout.n67 0.451012
R15320 Iout.n727 Iout.n726 0.451012
R15321 Iout.n727 Iout.n28 0.451012
R15322 Iout.n893 Iout.n28 0.451012
R15323 Iout.n204 Iout.n188 0.451012
R15324 Iout.n269 Iout.n188 0.451012
R15325 Iout.n269 Iout.n268 0.451012
R15326 Iout.n268 Iout.n161 0.451012
R15327 Iout.n422 Iout.n161 0.451012
R15328 Iout.n422 Iout.n421 0.451012
R15329 Iout.n421 Iout.n101 0.451012
R15330 Iout.n616 Iout.n101 0.451012
R15331 Iout.n616 Iout.n615 0.451012
R15332 Iout.n615 Iout.n58 0.451012
R15333 Iout.n745 Iout.n58 0.451012
R15334 Iout.n745 Iout.n744 0.451012
R15335 Iout.n744 Iout.n31 0.451012
R15336 Iout.n872 Iout.n31 0.451012
R15337 Iout.n498 Iout.n497 0.451012
R15338 Iout.n497 Iout.n151 0.451012
R15339 Iout.n467 Iout.n151 0.451012
R15340 Iout.n467 Iout.n466 0.451012
R15341 Iout.n466 Iout.n158 0.451012
R15342 Iout.n436 Iout.n158 0.451012
R15343 Iout.n436 Iout.n113 0.451012
R15344 Iout.n592 Iout.n113 0.451012
R15345 Iout.n592 Iout.n591 0.451012
R15346 Iout.n591 Iout.n70 0.451012
R15347 Iout.n721 Iout.n70 0.451012
R15348 Iout.n721 Iout.n720 0.451012
R15349 Iout.n720 Iout.n27 0.451012
R15350 Iout.n900 Iout.n27 0.451012
R15351 Iout.n208 Iout.n185 0.451012
R15352 Iout.n274 Iout.n185 0.451012
R15353 Iout.n275 Iout.n274 0.451012
R15354 Iout.n275 Iout.n162 0.451012
R15355 Iout.n413 Iout.n162 0.451012
R15356 Iout.n414 Iout.n413 0.451012
R15357 Iout.n414 Iout.n98 0.451012
R15358 Iout.n621 Iout.n98 0.451012
R15359 Iout.n622 Iout.n621 0.451012
R15360 Iout.n622 Iout.n55 0.451012
R15361 Iout.n750 Iout.n55 0.451012
R15362 Iout.n751 Iout.n750 0.451012
R15363 Iout.n751 Iout.n32 0.451012
R15364 Iout.n865 Iout.n32 0.451012
R15365 Iout.n502 Iout.n139 0.451012
R15366 Iout.n528 Iout.n139 0.451012
R15367 Iout.n529 Iout.n528 0.451012
R15368 Iout.n529 Iout.n126 0.451012
R15369 Iout.n551 Iout.n126 0.451012
R15370 Iout.n552 Iout.n551 0.451012
R15371 Iout.n552 Iout.n116 0.451012
R15372 Iout.n585 Iout.n116 0.451012
R15373 Iout.n586 Iout.n585 0.451012
R15374 Iout.n586 Iout.n73 0.451012
R15375 Iout.n714 Iout.n73 0.451012
R15376 Iout.n715 Iout.n714 0.451012
R15377 Iout.n715 Iout.n26 0.451012
R15378 Iout.n907 Iout.n26 0.451012
R15379 Iout.n212 Iout.n182 0.451012
R15380 Iout.n281 Iout.n182 0.451012
R15381 Iout.n281 Iout.n280 0.451012
R15382 Iout.n280 Iout.n163 0.451012
R15383 Iout.n406 Iout.n163 0.451012
R15384 Iout.n406 Iout.n405 0.451012
R15385 Iout.n405 Iout.n95 0.451012
R15386 Iout.n628 Iout.n95 0.451012
R15387 Iout.n628 Iout.n627 0.451012
R15388 Iout.n627 Iout.n52 0.451012
R15389 Iout.n757 Iout.n52 0.451012
R15390 Iout.n757 Iout.n756 0.451012
R15391 Iout.n756 Iout.n33 0.451012
R15392 Iout.n858 Iout.n33 0.451012
R15393 Iout.n522 Iout.n145 0.451012
R15394 Iout.n523 Iout.n522 0.451012
R15395 Iout.n523 Iout.n132 0.451012
R15396 Iout.n545 Iout.n132 0.451012
R15397 Iout.n546 Iout.n545 0.451012
R15398 Iout.n546 Iout.n119 0.451012
R15399 Iout.n572 Iout.n119 0.451012
R15400 Iout.n580 Iout.n572 0.451012
R15401 Iout.n580 Iout.n579 0.451012
R15402 Iout.n579 Iout.n76 0.451012
R15403 Iout.n709 Iout.n76 0.451012
R15404 Iout.n709 Iout.n708 0.451012
R15405 Iout.n708 Iout.n25 0.451012
R15406 Iout.n914 Iout.n25 0.451012
R15407 Iout.n216 Iout.n179 0.451012
R15408 Iout.n286 Iout.n179 0.451012
R15409 Iout.n287 Iout.n286 0.451012
R15410 Iout.n287 Iout.n164 0.451012
R15411 Iout.n397 Iout.n164 0.451012
R15412 Iout.n398 Iout.n397 0.451012
R15413 Iout.n398 Iout.n92 0.451012
R15414 Iout.n633 Iout.n92 0.451012
R15415 Iout.n634 Iout.n633 0.451012
R15416 Iout.n634 Iout.n49 0.451012
R15417 Iout.n762 Iout.n49 0.451012
R15418 Iout.n763 Iout.n762 0.451012
R15419 Iout.n763 Iout.n34 0.451012
R15420 Iout.n851 Iout.n34 0.451012
R15421 Iout.n517 Iout.n516 0.451012
R15422 Iout.n517 Iout.n138 0.451012
R15423 Iout.n539 Iout.n138 0.451012
R15424 Iout.n540 Iout.n539 0.451012
R15425 Iout.n540 Iout.n125 0.451012
R15426 Iout.n562 Iout.n125 0.451012
R15427 Iout.n567 Iout.n562 0.451012
R15428 Iout.n567 Iout.n566 0.451012
R15429 Iout.n566 Iout.n79 0.451012
R15430 Iout.n698 Iout.n79 0.451012
R15431 Iout.n702 Iout.n698 0.451012
R15432 Iout.n703 Iout.n702 0.451012
R15433 Iout.n703 Iout.n24 0.451012
R15434 Iout.n921 Iout.n24 0.451012
R15435 Iout.n220 Iout.n176 0.451012
R15436 Iout.n293 Iout.n176 0.451012
R15437 Iout.n293 Iout.n292 0.451012
R15438 Iout.n292 Iout.n165 0.451012
R15439 Iout.n390 Iout.n165 0.451012
R15440 Iout.n390 Iout.n389 0.451012
R15441 Iout.n389 Iout.n89 0.451012
R15442 Iout.n640 Iout.n89 0.451012
R15443 Iout.n640 Iout.n639 0.451012
R15444 Iout.n639 Iout.n46 0.451012
R15445 Iout.n769 Iout.n46 0.451012
R15446 Iout.n769 Iout.n768 0.451012
R15447 Iout.n768 Iout.n35 0.451012
R15448 Iout.n844 Iout.n35 0.451012
R15449 Iout.n511 Iout.n2 0.451012
R15450 Iout.n1005 Iout.n2 0.451012
R15451 Iout.n1005 Iout.n1004 0.451012
R15452 Iout.n1004 Iout.n3 0.451012
R15453 Iout.n986 Iout.n3 0.451012
R15454 Iout.n986 Iout.n985 0.451012
R15455 Iout.n985 Iout.n8 0.451012
R15456 Iout.n967 Iout.n8 0.451012
R15457 Iout.n967 Iout.n966 0.451012
R15458 Iout.n966 Iout.n13 0.451012
R15459 Iout.n948 Iout.n13 0.451012
R15460 Iout.n948 Iout.n947 0.451012
R15461 Iout.n947 Iout.n18 0.451012
R15462 Iout.n929 Iout.n18 0.451012
R15463 Iout.n224 Iout.n170 0.451012
R15464 Iout.n298 Iout.n170 0.451012
R15465 Iout.n299 Iout.n298 0.451012
R15466 Iout.n299 Iout.n166 0.451012
R15467 Iout.n381 Iout.n166 0.451012
R15468 Iout.n382 Iout.n381 0.451012
R15469 Iout.n382 Iout.n83 0.451012
R15470 Iout.n645 Iout.n83 0.451012
R15471 Iout.n646 Iout.n645 0.451012
R15472 Iout.n646 Iout.n40 0.451012
R15473 Iout.n774 Iout.n40 0.451012
R15474 Iout.n775 Iout.n774 0.451012
R15475 Iout.n775 Iout.n36 0.451012
R15476 Iout.n837 Iout.n36 0.451012
R15477 Iout.n1018 Iout.n1017 0.451012
R15478 Iout.n1017 Iout.n0 0.451012
R15479 Iout.n999 Iout.n0 0.451012
R15480 Iout.n999 Iout.n998 0.451012
R15481 Iout.n998 Iout.n6 0.451012
R15482 Iout.n980 Iout.n6 0.451012
R15483 Iout.n980 Iout.n979 0.451012
R15484 Iout.n979 Iout.n11 0.451012
R15485 Iout.n961 Iout.n11 0.451012
R15486 Iout.n961 Iout.n960 0.451012
R15487 Iout.n960 Iout.n16 0.451012
R15488 Iout.n942 Iout.n16 0.451012
R15489 Iout.n942 Iout.n941 0.451012
R15490 Iout.n941 Iout.n21 0.451012
R15491 Iout.n230 Iout.n229 0.451012
R15492 Iout.n230 Iout.n167 0.451012
R15493 Iout.n304 Iout.n167 0.451012
R15494 Iout.n332 Iout.n304 0.451012
R15495 Iout.n374 Iout.n332 0.451012
R15496 Iout.n374 Iout.n373 0.451012
R15497 Iout.n373 Iout.n369 0.451012
R15498 Iout.n369 Iout.n80 0.451012
R15499 Iout.n651 Iout.n80 0.451012
R15500 Iout.n652 Iout.n651 0.451012
R15501 Iout.n652 Iout.n37 0.451012
R15502 Iout.n780 Iout.n37 0.451012
R15503 Iout.n826 Iout.n780 0.451012
R15504 Iout.n830 Iout.n826 0.451012
R15505 Iout.n231 Iout 0.2919
R15506 Iout.n303 Iout 0.2919
R15507 Iout Iout.n300 0.2919
R15508 Iout.n375 Iout 0.2919
R15509 Iout.n380 Iout 0.2919
R15510 Iout.n391 Iout 0.2919
R15511 Iout.n368 Iout 0.2919
R15512 Iout Iout.n365 0.2919
R15513 Iout Iout.n362 0.2919
R15514 Iout Iout.n359 0.2919
R15515 Iout.n650 Iout 0.2919
R15516 Iout Iout.n647 0.2919
R15517 Iout.n638 Iout 0.2919
R15518 Iout Iout.n635 0.2919
R15519 Iout.n626 Iout 0.2919
R15520 Iout.n41 Iout 0.2919
R15521 Iout.n773 Iout 0.2919
R15522 Iout Iout.n770 0.2919
R15523 Iout.n761 Iout 0.2919
R15524 Iout Iout.n758 0.2919
R15525 Iout.n749 Iout 0.2919
R15526 Iout.n825 Iout 0.2919
R15527 Iout Iout.n822 0.2919
R15528 Iout Iout.n819 0.2919
R15529 Iout Iout.n816 0.2919
R15530 Iout Iout.n813 0.2919
R15531 Iout Iout.n810 0.2919
R15532 Iout Iout.n807 0.2919
R15533 Iout.n829 Iout 0.2919
R15534 Iout.n838 Iout 0.2919
R15535 Iout.n843 Iout 0.2919
R15536 Iout.n852 Iout 0.2919
R15537 Iout.n857 Iout 0.2919
R15538 Iout.n866 Iout 0.2919
R15539 Iout.n871 Iout 0.2919
R15540 Iout.n880 Iout 0.2919
R15541 Iout Iout.n925 0.2919
R15542 Iout.n928 Iout 0.2919
R15543 Iout.n922 Iout 0.2919
R15544 Iout.n913 Iout 0.2919
R15545 Iout.n908 Iout 0.2919
R15546 Iout.n899 Iout 0.2919
R15547 Iout.n894 Iout 0.2919
R15548 Iout.n885 Iout 0.2919
R15549 Iout.n831 Iout 0.2919
R15550 Iout.n836 Iout 0.2919
R15551 Iout.n845 Iout 0.2919
R15552 Iout.n850 Iout 0.2919
R15553 Iout.n859 Iout 0.2919
R15554 Iout.n864 Iout 0.2919
R15555 Iout.n873 Iout 0.2919
R15556 Iout.n878 Iout 0.2919
R15557 Iout.n887 Iout 0.2919
R15558 Iout.n892 Iout 0.2919
R15559 Iout.n933 Iout 0.2919
R15560 Iout.n930 Iout 0.2919
R15561 Iout.n920 Iout 0.2919
R15562 Iout.n915 Iout 0.2919
R15563 Iout.n906 Iout 0.2919
R15564 Iout.n901 Iout 0.2919
R15565 Iout.n940 Iout 0.2919
R15566 Iout Iout.n783 0.2919
R15567 Iout Iout.n786 0.2919
R15568 Iout Iout.n789 0.2919
R15569 Iout Iout.n792 0.2919
R15570 Iout Iout.n795 0.2919
R15571 Iout Iout.n798 0.2919
R15572 Iout Iout.n801 0.2919
R15573 Iout Iout.n804 0.2919
R15574 Iout.n779 Iout 0.2919
R15575 Iout Iout.n776 0.2919
R15576 Iout.n767 Iout 0.2919
R15577 Iout Iout.n764 0.2919
R15578 Iout.n755 Iout 0.2919
R15579 Iout Iout.n752 0.2919
R15580 Iout.n743 Iout 0.2919
R15581 Iout Iout.n740 0.2919
R15582 Iout.n731 Iout 0.2919
R15583 Iout Iout.n728 0.2919
R15584 Iout.n719 Iout 0.2919
R15585 Iout Iout.n943 0.2919
R15586 Iout.n946 Iout 0.2919
R15587 Iout Iout.n704 0.2919
R15588 Iout.n707 Iout 0.2919
R15589 Iout Iout.n716 0.2919
R15590 Iout.n952 Iout 0.2919
R15591 Iout.n949 Iout 0.2919
R15592 Iout.n701 Iout 0.2919
R15593 Iout Iout.n710 0.2919
R15594 Iout.n713 Iout 0.2919
R15595 Iout Iout.n722 0.2919
R15596 Iout.n725 Iout 0.2919
R15597 Iout Iout.n734 0.2919
R15598 Iout.n737 Iout 0.2919
R15599 Iout Iout.n746 0.2919
R15600 Iout.n653 Iout 0.2919
R15601 Iout.n656 Iout 0.2919
R15602 Iout.n659 Iout 0.2919
R15603 Iout.n662 Iout 0.2919
R15604 Iout.n665 Iout 0.2919
R15605 Iout.n668 Iout 0.2919
R15606 Iout.n671 Iout 0.2919
R15607 Iout.n674 Iout 0.2919
R15608 Iout.n677 Iout 0.2919
R15609 Iout.n680 Iout 0.2919
R15610 Iout.n683 Iout 0.2919
R15611 Iout.n686 Iout 0.2919
R15612 Iout.n959 Iout 0.2919
R15613 Iout Iout.n694 0.2919
R15614 Iout.n697 Iout 0.2919
R15615 Iout.n689 Iout 0.2919
R15616 Iout Iout.n962 0.2919
R15617 Iout.n965 Iout 0.2919
R15618 Iout Iout.n575 0.2919
R15619 Iout.n578 Iout 0.2919
R15620 Iout Iout.n587 0.2919
R15621 Iout.n590 Iout 0.2919
R15622 Iout Iout.n599 0.2919
R15623 Iout.n602 Iout 0.2919
R15624 Iout Iout.n611 0.2919
R15625 Iout.n614 Iout 0.2919
R15626 Iout Iout.n623 0.2919
R15627 Iout.n84 Iout 0.2919
R15628 Iout.n644 Iout 0.2919
R15629 Iout Iout.n641 0.2919
R15630 Iout.n632 Iout 0.2919
R15631 Iout Iout.n629 0.2919
R15632 Iout.n620 Iout 0.2919
R15633 Iout Iout.n617 0.2919
R15634 Iout.n608 Iout 0.2919
R15635 Iout Iout.n605 0.2919
R15636 Iout.n596 Iout 0.2919
R15637 Iout Iout.n593 0.2919
R15638 Iout.n584 Iout 0.2919
R15639 Iout Iout.n581 0.2919
R15640 Iout.n971 Iout 0.2919
R15641 Iout.n968 Iout 0.2919
R15642 Iout.n565 Iout 0.2919
R15643 Iout.n978 Iout 0.2919
R15644 Iout Iout.n122 0.2919
R15645 Iout Iout.n568 0.2919
R15646 Iout.n571 Iout 0.2919
R15647 Iout Iout.n335 0.2919
R15648 Iout Iout.n338 0.2919
R15649 Iout Iout.n341 0.2919
R15650 Iout Iout.n344 0.2919
R15651 Iout Iout.n347 0.2919
R15652 Iout Iout.n350 0.2919
R15653 Iout Iout.n353 0.2919
R15654 Iout Iout.n356 0.2919
R15655 Iout.n372 Iout 0.2919
R15656 Iout.n383 Iout 0.2919
R15657 Iout.n388 Iout 0.2919
R15658 Iout.n399 Iout 0.2919
R15659 Iout.n404 Iout 0.2919
R15660 Iout.n415 Iout 0.2919
R15661 Iout.n420 Iout 0.2919
R15662 Iout.n431 Iout 0.2919
R15663 Iout.n443 Iout 0.2919
R15664 Iout Iout.n440 0.2919
R15665 Iout Iout.n437 0.2919
R15666 Iout.n553 Iout 0.2919
R15667 Iout.n556 Iout 0.2919
R15668 Iout.n561 Iout 0.2919
R15669 Iout Iout.n981 0.2919
R15670 Iout.n984 Iout 0.2919
R15671 Iout.n990 Iout 0.2919
R15672 Iout.n987 Iout 0.2919
R15673 Iout Iout.n129 0.2919
R15674 Iout Iout.n547 0.2919
R15675 Iout.n550 Iout 0.2919
R15676 Iout Iout.n451 0.2919
R15677 Iout.n454 Iout 0.2919
R15678 Iout.n446 Iout 0.2919
R15679 Iout.n428 Iout 0.2919
R15680 Iout.n423 Iout 0.2919
R15681 Iout.n412 Iout 0.2919
R15682 Iout.n407 Iout 0.2919
R15683 Iout.n396 Iout 0.2919
R15684 Iout.n331 Iout 0.2919
R15685 Iout Iout.n328 0.2919
R15686 Iout Iout.n325 0.2919
R15687 Iout Iout.n322 0.2919
R15688 Iout Iout.n319 0.2919
R15689 Iout Iout.n316 0.2919
R15690 Iout Iout.n313 0.2919
R15691 Iout Iout.n310 0.2919
R15692 Iout Iout.n307 0.2919
R15693 Iout.n457 Iout 0.2919
R15694 Iout.n465 Iout 0.2919
R15695 Iout Iout.n462 0.2919
R15696 Iout.n544 Iout 0.2919
R15697 Iout Iout.n541 0.2919
R15698 Iout Iout.n135 0.2919
R15699 Iout.n997 Iout 0.2919
R15700 Iout Iout.n1000 0.2919
R15701 Iout.n1003 Iout 0.2919
R15702 Iout.n538 Iout 0.2919
R15703 Iout.n533 Iout 0.2919
R15704 Iout.n530 Iout 0.2919
R15705 Iout Iout.n468 0.2919
R15706 Iout Iout.n471 0.2919
R15707 Iout.n474 Iout 0.2919
R15708 Iout Iout.n264 0.2919
R15709 Iout.n267 Iout 0.2919
R15710 Iout Iout.n276 0.2919
R15711 Iout.n279 Iout 0.2919
R15712 Iout Iout.n288 0.2919
R15713 Iout.n291 Iout 0.2919
R15714 Iout.n171 Iout 0.2919
R15715 Iout.n297 Iout 0.2919
R15716 Iout Iout.n294 0.2919
R15717 Iout.n285 Iout 0.2919
R15718 Iout Iout.n282 0.2919
R15719 Iout.n273 Iout 0.2919
R15720 Iout Iout.n270 0.2919
R15721 Iout.n261 Iout 0.2919
R15722 Iout.n477 Iout 0.2919
R15723 Iout.n485 Iout 0.2919
R15724 Iout Iout.n482 0.2919
R15725 Iout.n527 Iout 0.2919
R15726 Iout Iout.n524 0.2919
R15727 Iout Iout.n142 0.2919
R15728 Iout.n1006 Iout 0.2919
R15729 Iout.n1009 Iout 0.2919
R15730 Iout.n1016 Iout 0.2919
R15731 Iout Iout.n148 0.2919
R15732 Iout Iout.n518 0.2919
R15733 Iout.n521 Iout 0.2919
R15734 Iout Iout.n493 0.2919
R15735 Iout.n496 Iout 0.2919
R15736 Iout.n488 Iout 0.2919
R15737 Iout Iout.n254 0.2919
R15738 Iout.n257 Iout 0.2919
R15739 Iout.n249 Iout 0.2919
R15740 Iout.n246 Iout 0.2919
R15741 Iout.n243 Iout 0.2919
R15742 Iout.n240 Iout 0.2919
R15743 Iout.n237 Iout 0.2919
R15744 Iout.n234 Iout 0.2919
R15745 Iout.n228 Iout 0.2919
R15746 Iout Iout.n225 0.2919
R15747 Iout Iout.n221 0.2919
R15748 Iout Iout.n217 0.2919
R15749 Iout Iout.n213 0.2919
R15750 Iout Iout.n209 0.2919
R15751 Iout Iout.n205 0.2919
R15752 Iout Iout.n201 0.2919
R15753 Iout Iout.n198 0.2919
R15754 Iout Iout.n194 0.2919
R15755 Iout.n499 Iout 0.2919
R15756 Iout.n503 Iout 0.2919
R15757 Iout.n506 Iout 0.2919
R15758 Iout.n515 Iout 0.2919
R15759 Iout Iout.n512 0.2919
R15760 Iout.n1019 Iout 0.2919
R15761 Iout.n1013 Iout.n1012 0.092855
R15762 Iout.n1012 Iout.n1 0.092855
R15763 Iout.n994 Iout.n1 0.092855
R15764 Iout.n994 Iout.n993 0.092855
R15765 Iout.n993 Iout.n7 0.092855
R15766 Iout.n975 Iout.n7 0.092855
R15767 Iout.n975 Iout.n974 0.092855
R15768 Iout.n974 Iout.n12 0.092855
R15769 Iout.n956 Iout.n12 0.092855
R15770 Iout.n956 Iout.n955 0.092855
R15771 Iout.n955 Iout.n17 0.092855
R15772 Iout.n937 Iout.n17 0.092855
R15773 Iout.n937 Iout.n936 0.092855
R15774 Iout.n197 Iout 0.0818902
R15775 Iout.n191 Iout 0.0818902
R15776 Iout.n152 Iout 0.0818902
R15777 Iout.n204 Iout 0.0818902
R15778 Iout.n498 Iout 0.0818902
R15779 Iout.n208 Iout 0.0818902
R15780 Iout.n502 Iout 0.0818902
R15781 Iout.n212 Iout 0.0818902
R15782 Iout.n145 Iout 0.0818902
R15783 Iout.n216 Iout 0.0818902
R15784 Iout.n516 Iout 0.0818902
R15785 Iout.n220 Iout 0.0818902
R15786 Iout.n511 Iout 0.0818902
R15787 Iout.n224 Iout 0.0818902
R15788 Iout.n1018 Iout 0.0818902
R15789 Iout.n229 Iout 0.0818902
R15790 Iout.n1013 Iout 0.072645
R15791 Iout.n302 Iout 0.0532071
R15792 Iout Iout.n377 0.0532071
R15793 Iout.n379 Iout 0.0532071
R15794 Iout.n367 Iout 0.0532071
R15795 Iout.n364 Iout 0.0532071
R15796 Iout.n361 Iout 0.0532071
R15797 Iout.n649 Iout 0.0532071
R15798 Iout Iout.n82 0.0532071
R15799 Iout.n637 Iout 0.0532071
R15800 Iout Iout.n91 0.0532071
R15801 Iout Iout.n43 0.0532071
R15802 Iout.n772 Iout 0.0532071
R15803 Iout Iout.n45 0.0532071
R15804 Iout.n760 Iout 0.0532071
R15805 Iout Iout.n51 0.0532071
R15806 Iout.n824 Iout 0.0532071
R15807 Iout.n821 Iout 0.0532071
R15808 Iout.n818 Iout 0.0532071
R15809 Iout.n815 Iout 0.0532071
R15810 Iout.n812 Iout 0.0532071
R15811 Iout.n809 Iout 0.0532071
R15812 Iout.n828 Iout 0.0532071
R15813 Iout Iout.n840 0.0532071
R15814 Iout.n842 Iout 0.0532071
R15815 Iout Iout.n854 0.0532071
R15816 Iout.n856 Iout 0.0532071
R15817 Iout Iout.n868 0.0532071
R15818 Iout.n870 Iout 0.0532071
R15819 Iout.n927 Iout 0.0532071
R15820 Iout Iout.n924 0.0532071
R15821 Iout.n912 Iout 0.0532071
R15822 Iout Iout.n910 0.0532071
R15823 Iout.n898 Iout 0.0532071
R15824 Iout Iout.n896 0.0532071
R15825 Iout.n884 Iout 0.0532071
R15826 Iout Iout.n882 0.0532071
R15827 Iout Iout.n833 0.0532071
R15828 Iout.n835 Iout 0.0532071
R15829 Iout Iout.n847 0.0532071
R15830 Iout.n849 Iout 0.0532071
R15831 Iout Iout.n861 0.0532071
R15832 Iout.n863 Iout 0.0532071
R15833 Iout Iout.n875 0.0532071
R15834 Iout.n877 Iout 0.0532071
R15835 Iout Iout.n889 0.0532071
R15836 Iout Iout.n932 0.0532071
R15837 Iout.n919 Iout 0.0532071
R15838 Iout Iout.n917 0.0532071
R15839 Iout.n905 Iout 0.0532071
R15840 Iout Iout.n903 0.0532071
R15841 Iout.n891 Iout 0.0532071
R15842 Iout.n782 Iout 0.0532071
R15843 Iout.n785 Iout 0.0532071
R15844 Iout.n788 Iout 0.0532071
R15845 Iout.n791 Iout 0.0532071
R15846 Iout.n794 Iout 0.0532071
R15847 Iout.n797 Iout 0.0532071
R15848 Iout.n800 Iout 0.0532071
R15849 Iout.n803 Iout 0.0532071
R15850 Iout.n806 Iout 0.0532071
R15851 Iout.n778 Iout 0.0532071
R15852 Iout Iout.n39 0.0532071
R15853 Iout.n766 Iout 0.0532071
R15854 Iout Iout.n48 0.0532071
R15855 Iout.n754 Iout 0.0532071
R15856 Iout Iout.n54 0.0532071
R15857 Iout.n742 Iout 0.0532071
R15858 Iout Iout.n60 0.0532071
R15859 Iout.n730 Iout 0.0532071
R15860 Iout Iout.n66 0.0532071
R15861 Iout.n945 Iout 0.0532071
R15862 Iout.n78 Iout 0.0532071
R15863 Iout.n706 Iout 0.0532071
R15864 Iout Iout.n72 0.0532071
R15865 Iout.n718 Iout 0.0532071
R15866 Iout Iout.n951 0.0532071
R15867 Iout.n700 Iout 0.0532071
R15868 Iout Iout.n75 0.0532071
R15869 Iout.n712 Iout 0.0532071
R15870 Iout Iout.n69 0.0532071
R15871 Iout.n724 Iout 0.0532071
R15872 Iout Iout.n63 0.0532071
R15873 Iout.n736 Iout 0.0532071
R15874 Iout Iout.n57 0.0532071
R15875 Iout.n748 Iout 0.0532071
R15876 Iout Iout.n655 0.0532071
R15877 Iout Iout.n658 0.0532071
R15878 Iout Iout.n661 0.0532071
R15879 Iout Iout.n664 0.0532071
R15880 Iout Iout.n667 0.0532071
R15881 Iout Iout.n670 0.0532071
R15882 Iout Iout.n673 0.0532071
R15883 Iout Iout.n676 0.0532071
R15884 Iout Iout.n679 0.0532071
R15885 Iout Iout.n682 0.0532071
R15886 Iout Iout.n685 0.0532071
R15887 Iout.n693 Iout 0.0532071
R15888 Iout.n696 Iout 0.0532071
R15889 Iout Iout.n691 0.0532071
R15890 Iout Iout.n688 0.0532071
R15891 Iout.n964 Iout 0.0532071
R15892 Iout.n574 Iout 0.0532071
R15893 Iout.n577 Iout 0.0532071
R15894 Iout Iout.n115 0.0532071
R15895 Iout.n589 Iout 0.0532071
R15896 Iout Iout.n109 0.0532071
R15897 Iout.n601 Iout 0.0532071
R15898 Iout Iout.n103 0.0532071
R15899 Iout.n613 Iout 0.0532071
R15900 Iout Iout.n97 0.0532071
R15901 Iout.n625 Iout 0.0532071
R15902 Iout Iout.n86 0.0532071
R15903 Iout.n643 Iout 0.0532071
R15904 Iout Iout.n88 0.0532071
R15905 Iout.n631 Iout 0.0532071
R15906 Iout Iout.n94 0.0532071
R15907 Iout.n619 Iout 0.0532071
R15908 Iout Iout.n100 0.0532071
R15909 Iout.n607 Iout 0.0532071
R15910 Iout Iout.n106 0.0532071
R15911 Iout.n595 Iout 0.0532071
R15912 Iout Iout.n112 0.0532071
R15913 Iout.n583 Iout 0.0532071
R15914 Iout Iout.n970 0.0532071
R15915 Iout.n564 Iout 0.0532071
R15916 Iout Iout.n118 0.0532071
R15917 Iout.n121 Iout 0.0532071
R15918 Iout.n124 Iout 0.0532071
R15919 Iout.n570 Iout 0.0532071
R15920 Iout.n334 Iout 0.0532071
R15921 Iout.n337 Iout 0.0532071
R15922 Iout.n340 Iout 0.0532071
R15923 Iout.n343 Iout 0.0532071
R15924 Iout.n346 Iout 0.0532071
R15925 Iout.n349 Iout 0.0532071
R15926 Iout.n352 Iout 0.0532071
R15927 Iout.n355 Iout 0.0532071
R15928 Iout.n358 Iout 0.0532071
R15929 Iout.n371 Iout 0.0532071
R15930 Iout Iout.n385 0.0532071
R15931 Iout.n387 Iout 0.0532071
R15932 Iout Iout.n401 0.0532071
R15933 Iout.n403 Iout 0.0532071
R15934 Iout Iout.n417 0.0532071
R15935 Iout.n419 Iout 0.0532071
R15936 Iout Iout.n433 0.0532071
R15937 Iout.n442 Iout 0.0532071
R15938 Iout.n439 Iout 0.0532071
R15939 Iout.n435 Iout 0.0532071
R15940 Iout Iout.n555 0.0532071
R15941 Iout Iout.n558 0.0532071
R15942 Iout.n983 Iout 0.0532071
R15943 Iout.n560 Iout 0.0532071
R15944 Iout Iout.n989 0.0532071
R15945 Iout.n128 Iout 0.0532071
R15946 Iout.n131 Iout 0.0532071
R15947 Iout.n549 Iout 0.0532071
R15948 Iout.n450 Iout 0.0532071
R15949 Iout.n453 Iout 0.0532071
R15950 Iout Iout.n448 0.0532071
R15951 Iout.n427 Iout 0.0532071
R15952 Iout Iout.n425 0.0532071
R15953 Iout.n411 Iout 0.0532071
R15954 Iout Iout.n409 0.0532071
R15955 Iout.n395 Iout 0.0532071
R15956 Iout Iout.n393 0.0532071
R15957 Iout.n330 Iout 0.0532071
R15958 Iout.n327 Iout 0.0532071
R15959 Iout.n324 Iout 0.0532071
R15960 Iout.n321 Iout 0.0532071
R15961 Iout.n318 Iout 0.0532071
R15962 Iout.n315 Iout 0.0532071
R15963 Iout.n312 Iout 0.0532071
R15964 Iout.n309 Iout 0.0532071
R15965 Iout.n306 Iout 0.0532071
R15966 Iout Iout.n459 0.0532071
R15967 Iout.n464 Iout 0.0532071
R15968 Iout.n461 Iout 0.0532071
R15969 Iout.n543 Iout 0.0532071
R15970 Iout.n137 Iout 0.0532071
R15971 Iout.n134 Iout 0.0532071
R15972 Iout.n1002 Iout 0.0532071
R15973 Iout.n537 Iout 0.0532071
R15974 Iout Iout.n535 0.0532071
R15975 Iout Iout.n532 0.0532071
R15976 Iout.n157 Iout 0.0532071
R15977 Iout.n470 Iout 0.0532071
R15978 Iout.n473 Iout 0.0532071
R15979 Iout.n190 Iout 0.0532071
R15980 Iout.n266 Iout 0.0532071
R15981 Iout Iout.n184 0.0532071
R15982 Iout.n278 Iout 0.0532071
R15983 Iout Iout.n178 0.0532071
R15984 Iout.n290 Iout 0.0532071
R15985 Iout Iout.n169 0.0532071
R15986 Iout Iout.n173 0.0532071
R15987 Iout.n296 Iout 0.0532071
R15988 Iout Iout.n175 0.0532071
R15989 Iout.n284 Iout 0.0532071
R15990 Iout Iout.n181 0.0532071
R15991 Iout.n272 Iout 0.0532071
R15992 Iout Iout.n187 0.0532071
R15993 Iout.n260 Iout 0.0532071
R15994 Iout Iout.n479 0.0532071
R15995 Iout.n484 Iout 0.0532071
R15996 Iout.n481 Iout 0.0532071
R15997 Iout.n526 Iout 0.0532071
R15998 Iout.n144 Iout 0.0532071
R15999 Iout.n141 Iout 0.0532071
R16000 Iout Iout.n1008 0.0532071
R16001 Iout.n147 Iout 0.0532071
R16002 Iout.n150 Iout 0.0532071
R16003 Iout.n520 Iout 0.0532071
R16004 Iout.n492 Iout 0.0532071
R16005 Iout.n495 Iout 0.0532071
R16006 Iout Iout.n490 0.0532071
R16007 Iout.n253 Iout 0.0532071
R16008 Iout.n256 Iout 0.0532071
R16009 Iout Iout.n251 0.0532071
R16010 Iout Iout.n248 0.0532071
R16011 Iout Iout.n245 0.0532071
R16012 Iout Iout.n242 0.0532071
R16013 Iout Iout.n239 0.0532071
R16014 Iout Iout.n236 0.0532071
R16015 Iout Iout.n233 0.0532071
R16016 Iout.n227 Iout 0.0532071
R16017 Iout.n223 Iout 0.0532071
R16018 Iout.n219 Iout 0.0532071
R16019 Iout.n215 Iout 0.0532071
R16020 Iout.n211 Iout 0.0532071
R16021 Iout.n207 Iout 0.0532071
R16022 Iout.n203 Iout 0.0532071
R16023 Iout.n200 Iout 0.0532071
R16024 Iout.n196 Iout 0.0532071
R16025 Iout.n193 Iout 0.0532071
R16026 Iout Iout.n501 0.0532071
R16027 Iout Iout.n505 0.0532071
R16028 Iout Iout.n508 0.0532071
R16029 Iout.n514 Iout 0.0532071
R16030 Iout.n510 Iout 0.0532071
R16031 Iout.n1020 Iout 0.03925
R16032 Iout.n509 Iout 0.03925
R16033 Iout.n513 Iout 0.03925
R16034 Iout.n507 Iout 0.03925
R16035 Iout.n504 Iout 0.03925
R16036 Iout.n500 Iout 0.03925
R16037 Iout.n192 Iout 0.03925
R16038 Iout.n195 Iout 0.03925
R16039 Iout.n199 Iout 0.03925
R16040 Iout.n202 Iout 0.03925
R16041 Iout.n206 Iout 0.03925
R16042 Iout.n210 Iout 0.03925
R16043 Iout.n214 Iout 0.03925
R16044 Iout.n218 Iout 0.03925
R16045 Iout.n222 Iout 0.03925
R16046 Iout.n226 Iout 0.03925
R16047 Iout.n232 Iout 0.03925
R16048 Iout.n235 Iout 0.03925
R16049 Iout.n238 Iout 0.03925
R16050 Iout.n241 Iout 0.03925
R16051 Iout.n244 Iout 0.03925
R16052 Iout.n247 Iout 0.03925
R16053 Iout.n250 Iout 0.03925
R16054 Iout.n255 Iout 0.03925
R16055 Iout.n252 Iout 0.03925
R16056 Iout.n489 Iout 0.03925
R16057 Iout.n494 Iout 0.03925
R16058 Iout.n491 Iout 0.03925
R16059 Iout.n519 Iout 0.03925
R16060 Iout.n149 Iout 0.03925
R16061 Iout.n146 Iout 0.03925
R16062 Iout.n1010 Iout 0.03925
R16063 Iout.n1007 Iout 0.03925
R16064 Iout.n140 Iout 0.03925
R16065 Iout.n143 Iout 0.03925
R16066 Iout.n525 Iout 0.03925
R16067 Iout.n480 Iout 0.03925
R16068 Iout.n483 Iout 0.03925
R16069 Iout.n478 Iout 0.03925
R16070 Iout.n259 Iout 0.03925
R16071 Iout.n186 Iout 0.03925
R16072 Iout.n271 Iout 0.03925
R16073 Iout.n180 Iout 0.03925
R16074 Iout.n283 Iout 0.03925
R16075 Iout.n174 Iout 0.03925
R16076 Iout.n168 Iout 0.03925
R16077 Iout.n301 Iout 0.03925
R16078 Iout.n289 Iout 0.03925
R16079 Iout.n177 Iout 0.03925
R16080 Iout.n277 Iout 0.03925
R16081 Iout.n183 Iout 0.03925
R16082 Iout.n265 Iout 0.03925
R16083 Iout.n189 Iout 0.03925
R16084 Iout.n472 Iout 0.03925
R16085 Iout.n469 Iout 0.03925
R16086 Iout.n156 Iout 0.03925
R16087 Iout.n531 Iout 0.03925
R16088 Iout.n534 Iout 0.03925
R16089 Iout.n536 Iout 0.03925
R16090 Iout.n133 Iout 0.03925
R16091 Iout.n136 Iout 0.03925
R16092 Iout.n542 Iout 0.03925
R16093 Iout.n460 Iout 0.03925
R16094 Iout.n463 Iout 0.03925
R16095 Iout.n458 Iout 0.03925
R16096 Iout.n305 Iout 0.03925
R16097 Iout.n308 Iout 0.03925
R16098 Iout.n311 Iout 0.03925
R16099 Iout.n314 Iout 0.03925
R16100 Iout.n317 Iout 0.03925
R16101 Iout.n320 Iout 0.03925
R16102 Iout.n392 Iout 0.03925
R16103 Iout.n378 Iout 0.03925
R16104 Iout.n376 Iout 0.03925
R16105 Iout.n394 Iout 0.03925
R16106 Iout.n408 Iout 0.03925
R16107 Iout.n410 Iout 0.03925
R16108 Iout.n424 Iout 0.03925
R16109 Iout.n426 Iout 0.03925
R16110 Iout.n447 Iout 0.03925
R16111 Iout.n452 Iout 0.03925
R16112 Iout.n449 Iout 0.03925
R16113 Iout.n548 Iout 0.03925
R16114 Iout.n130 Iout 0.03925
R16115 Iout.n559 Iout 0.03925
R16116 Iout.n557 Iout 0.03925
R16117 Iout.n554 Iout 0.03925
R16118 Iout.n434 Iout 0.03925
R16119 Iout.n438 Iout 0.03925
R16120 Iout.n441 Iout 0.03925
R16121 Iout.n432 Iout 0.03925
R16122 Iout.n418 Iout 0.03925
R16123 Iout.n416 Iout 0.03925
R16124 Iout.n402 Iout 0.03925
R16125 Iout.n357 Iout 0.03925
R16126 Iout.n360 Iout 0.03925
R16127 Iout.n363 Iout 0.03925
R16128 Iout.n366 Iout 0.03925
R16129 Iout.n354 Iout 0.03925
R16130 Iout.n351 Iout 0.03925
R16131 Iout.n348 Iout 0.03925
R16132 Iout.n345 Iout 0.03925
R16133 Iout.n342 Iout 0.03925
R16134 Iout.n339 Iout 0.03925
R16135 Iout.n336 Iout 0.03925
R16136 Iout.n333 Iout 0.03925
R16137 Iout.n117 Iout 0.03925
R16138 Iout.n582 Iout 0.03925
R16139 Iout.n111 Iout 0.03925
R16140 Iout.n594 Iout 0.03925
R16141 Iout.n105 Iout 0.03925
R16142 Iout.n606 Iout 0.03925
R16143 Iout.n99 Iout 0.03925
R16144 Iout.n618 Iout 0.03925
R16145 Iout.n624 Iout 0.03925
R16146 Iout.n90 Iout 0.03925
R16147 Iout.n636 Iout 0.03925
R16148 Iout.n81 Iout 0.03925
R16149 Iout.n648 Iout 0.03925
R16150 Iout.n96 Iout 0.03925
R16151 Iout.n612 Iout 0.03925
R16152 Iout.n102 Iout 0.03925
R16153 Iout.n600 Iout 0.03925
R16154 Iout.n108 Iout 0.03925
R16155 Iout.n588 Iout 0.03925
R16156 Iout.n687 Iout 0.03925
R16157 Iout.n684 Iout 0.03925
R16158 Iout.n681 Iout 0.03925
R16159 Iout.n678 Iout 0.03925
R16160 Iout.n675 Iout 0.03925
R16161 Iout.n672 Iout 0.03925
R16162 Iout.n747 Iout 0.03925
R16163 Iout.n50 Iout 0.03925
R16164 Iout.n759 Iout 0.03925
R16165 Iout.n44 Iout 0.03925
R16166 Iout.n771 Iout 0.03925
R16167 Iout.n42 Iout 0.03925
R16168 Iout.n56 Iout 0.03925
R16169 Iout.n735 Iout 0.03925
R16170 Iout.n62 Iout 0.03925
R16171 Iout.n723 Iout 0.03925
R16172 Iout.n717 Iout 0.03925
R16173 Iout.n65 Iout 0.03925
R16174 Iout.n729 Iout 0.03925
R16175 Iout.n59 Iout 0.03925
R16176 Iout.n805 Iout 0.03925
R16177 Iout.n808 Iout 0.03925
R16178 Iout.n811 Iout 0.03925
R16179 Iout.n814 Iout 0.03925
R16180 Iout.n817 Iout 0.03925
R16181 Iout.n820 Iout 0.03925
R16182 Iout.n823 Iout 0.03925
R16183 Iout.n802 Iout 0.03925
R16184 Iout.n799 Iout 0.03925
R16185 Iout.n890 Iout 0.03925
R16186 Iout.n888 Iout 0.03925
R16187 Iout.n881 Iout 0.03925
R16188 Iout.n869 Iout 0.03925
R16189 Iout.n867 Iout 0.03925
R16190 Iout.n855 Iout 0.03925
R16191 Iout.n853 Iout 0.03925
R16192 Iout.n841 Iout 0.03925
R16193 Iout.n839 Iout 0.03925
R16194 Iout.n827 Iout 0.03925
R16195 Iout.n883 Iout 0.03925
R16196 Iout.n895 Iout 0.03925
R16197 Iout.n897 Iout 0.03925
R16198 Iout.n909 Iout 0.03925
R16199 Iout.n911 Iout 0.03925
R16200 Iout.n923 Iout 0.03925
R16201 Iout.n926 Iout 0.03925
R16202 Iout.n22 Iout 0.03925
R16203 Iout.n876 Iout 0.03925
R16204 Iout.n874 Iout 0.03925
R16205 Iout.n862 Iout 0.03925
R16206 Iout.n860 Iout 0.03925
R16207 Iout.n848 Iout 0.03925
R16208 Iout.n846 Iout 0.03925
R16209 Iout.n834 Iout 0.03925
R16210 Iout.n832 Iout 0.03925
R16211 Iout.n902 Iout 0.03925
R16212 Iout.n904 Iout 0.03925
R16213 Iout.n916 Iout 0.03925
R16214 Iout.n918 Iout 0.03925
R16215 Iout.n931 Iout 0.03925
R16216 Iout.n934 Iout 0.03925
R16217 Iout.n796 Iout 0.03925
R16218 Iout.n793 Iout 0.03925
R16219 Iout.n790 Iout 0.03925
R16220 Iout.n787 Iout 0.03925
R16221 Iout.n784 Iout 0.03925
R16222 Iout.n781 Iout 0.03925
R16223 Iout.n938 Iout 0.03925
R16224 Iout.n741 Iout 0.03925
R16225 Iout.n53 Iout 0.03925
R16226 Iout.n753 Iout 0.03925
R16227 Iout.n47 Iout 0.03925
R16228 Iout.n765 Iout 0.03925
R16229 Iout.n38 Iout 0.03925
R16230 Iout.n777 Iout 0.03925
R16231 Iout.n71 Iout 0.03925
R16232 Iout.n705 Iout 0.03925
R16233 Iout.n77 Iout 0.03925
R16234 Iout.n944 Iout 0.03925
R16235 Iout.n19 Iout 0.03925
R16236 Iout.n68 Iout 0.03925
R16237 Iout.n711 Iout 0.03925
R16238 Iout.n74 Iout 0.03925
R16239 Iout.n699 Iout 0.03925
R16240 Iout.n950 Iout 0.03925
R16241 Iout.n953 Iout 0.03925
R16242 Iout.n669 Iout 0.03925
R16243 Iout.n666 Iout 0.03925
R16244 Iout.n663 Iout 0.03925
R16245 Iout.n660 Iout 0.03925
R16246 Iout.n657 Iout 0.03925
R16247 Iout.n654 Iout 0.03925
R16248 Iout.n690 Iout 0.03925
R16249 Iout.n695 Iout 0.03925
R16250 Iout.n692 Iout 0.03925
R16251 Iout.n957 Iout 0.03925
R16252 Iout.n114 Iout 0.03925
R16253 Iout.n576 Iout 0.03925
R16254 Iout.n573 Iout 0.03925
R16255 Iout.n963 Iout 0.03925
R16256 Iout.n14 Iout 0.03925
R16257 Iout.n93 Iout 0.03925
R16258 Iout.n630 Iout 0.03925
R16259 Iout.n87 Iout 0.03925
R16260 Iout.n642 Iout 0.03925
R16261 Iout.n85 Iout 0.03925
R16262 Iout.n563 Iout 0.03925
R16263 Iout.n969 Iout 0.03925
R16264 Iout.n972 Iout 0.03925
R16265 Iout.n569 Iout 0.03925
R16266 Iout.n123 Iout 0.03925
R16267 Iout.n120 Iout 0.03925
R16268 Iout.n976 Iout 0.03925
R16269 Iout.n400 Iout 0.03925
R16270 Iout.n386 Iout 0.03925
R16271 Iout.n384 Iout 0.03925
R16272 Iout.n370 Iout 0.03925
R16273 Iout.n982 Iout 0.03925
R16274 Iout.n9 Iout 0.03925
R16275 Iout.n127 Iout 0.03925
R16276 Iout.n988 Iout 0.03925
R16277 Iout.n991 Iout 0.03925
R16278 Iout.n323 Iout 0.03925
R16279 Iout.n326 Iout 0.03925
R16280 Iout.n329 Iout 0.03925
R16281 Iout.n995 Iout 0.03925
R16282 Iout.n1001 Iout 0.03925
R16283 Iout.n4 Iout 0.03925
R16284 Iout.n295 Iout 0.03925
R16285 Iout.n172 Iout 0.03925
R16286 Iout.n1014 Iout 0.03925
R16287 Iout.n1022 Iout 0.02071
R16288 Iout Iout.n1022 0.00379
R16289 Iout.n303 Iout.n302 0.00105952
R16290 Iout.n377 Iout.n375 0.00105952
R16291 Iout.n380 Iout.n379 0.00105952
R16292 Iout.n368 Iout.n367 0.00105952
R16293 Iout.n365 Iout.n364 0.00105952
R16294 Iout.n362 Iout.n361 0.00105952
R16295 Iout.n650 Iout.n649 0.00105952
R16296 Iout.n647 Iout.n82 0.00105952
R16297 Iout.n638 Iout.n637 0.00105952
R16298 Iout.n635 Iout.n91 0.00105952
R16299 Iout.n43 Iout.n41 0.00105952
R16300 Iout.n773 Iout.n772 0.00105952
R16301 Iout.n770 Iout.n45 0.00105952
R16302 Iout.n761 Iout.n760 0.00105952
R16303 Iout.n758 Iout.n51 0.00105952
R16304 Iout.n825 Iout.n824 0.00105952
R16305 Iout.n822 Iout.n821 0.00105952
R16306 Iout.n819 Iout.n818 0.00105952
R16307 Iout.n816 Iout.n815 0.00105952
R16308 Iout.n813 Iout.n812 0.00105952
R16309 Iout.n810 Iout.n809 0.00105952
R16310 Iout.n829 Iout.n828 0.00105952
R16311 Iout.n840 Iout.n838 0.00105952
R16312 Iout.n843 Iout.n842 0.00105952
R16313 Iout.n854 Iout.n852 0.00105952
R16314 Iout.n857 Iout.n856 0.00105952
R16315 Iout.n868 Iout.n866 0.00105952
R16316 Iout.n871 Iout.n870 0.00105952
R16317 Iout.n925 Iout.n23 0.00105952
R16318 Iout.n928 Iout.n927 0.00105952
R16319 Iout.n924 Iout.n922 0.00105952
R16320 Iout.n913 Iout.n912 0.00105952
R16321 Iout.n910 Iout.n908 0.00105952
R16322 Iout.n899 Iout.n898 0.00105952
R16323 Iout.n896 Iout.n894 0.00105952
R16324 Iout.n885 Iout.n884 0.00105952
R16325 Iout.n882 Iout.n880 0.00105952
R16326 Iout.n833 Iout.n831 0.00105952
R16327 Iout.n836 Iout.n835 0.00105952
R16328 Iout.n847 Iout.n845 0.00105952
R16329 Iout.n850 Iout.n849 0.00105952
R16330 Iout.n861 Iout.n859 0.00105952
R16331 Iout.n864 Iout.n863 0.00105952
R16332 Iout.n875 Iout.n873 0.00105952
R16333 Iout.n878 Iout.n877 0.00105952
R16334 Iout.n889 Iout.n887 0.00105952
R16335 Iout.n935 Iout.n933 0.00105952
R16336 Iout.n932 Iout.n930 0.00105952
R16337 Iout.n920 Iout.n919 0.00105952
R16338 Iout.n917 Iout.n915 0.00105952
R16339 Iout.n906 Iout.n905 0.00105952
R16340 Iout.n903 Iout.n901 0.00105952
R16341 Iout.n892 Iout.n891 0.00105952
R16342 Iout.n940 Iout.n939 0.00105952
R16343 Iout.n783 Iout.n782 0.00105952
R16344 Iout.n786 Iout.n785 0.00105952
R16345 Iout.n789 Iout.n788 0.00105952
R16346 Iout.n792 Iout.n791 0.00105952
R16347 Iout.n795 Iout.n794 0.00105952
R16348 Iout.n798 Iout.n797 0.00105952
R16349 Iout.n801 Iout.n800 0.00105952
R16350 Iout.n804 Iout.n803 0.00105952
R16351 Iout.n807 Iout.n806 0.00105952
R16352 Iout.n779 Iout.n778 0.00105952
R16353 Iout.n776 Iout.n39 0.00105952
R16354 Iout.n767 Iout.n766 0.00105952
R16355 Iout.n764 Iout.n48 0.00105952
R16356 Iout.n755 Iout.n754 0.00105952
R16357 Iout.n752 Iout.n54 0.00105952
R16358 Iout.n743 Iout.n742 0.00105952
R16359 Iout.n740 Iout.n60 0.00105952
R16360 Iout.n731 Iout.n730 0.00105952
R16361 Iout.n728 Iout.n66 0.00105952
R16362 Iout.n943 Iout.n20 0.00105952
R16363 Iout.n946 Iout.n945 0.00105952
R16364 Iout.n704 Iout.n78 0.00105952
R16365 Iout.n707 Iout.n706 0.00105952
R16366 Iout.n716 Iout.n72 0.00105952
R16367 Iout.n719 Iout.n718 0.00105952
R16368 Iout.n954 Iout.n952 0.00105952
R16369 Iout.n951 Iout.n949 0.00105952
R16370 Iout.n701 Iout.n700 0.00105952
R16371 Iout.n710 Iout.n75 0.00105952
R16372 Iout.n713 Iout.n712 0.00105952
R16373 Iout.n722 Iout.n69 0.00105952
R16374 Iout.n725 Iout.n724 0.00105952
R16375 Iout.n734 Iout.n63 0.00105952
R16376 Iout.n737 Iout.n736 0.00105952
R16377 Iout.n746 Iout.n57 0.00105952
R16378 Iout.n749 Iout.n748 0.00105952
R16379 Iout.n655 Iout.n653 0.00105952
R16380 Iout.n658 Iout.n656 0.00105952
R16381 Iout.n661 Iout.n659 0.00105952
R16382 Iout.n664 Iout.n662 0.00105952
R16383 Iout.n667 Iout.n665 0.00105952
R16384 Iout.n670 Iout.n668 0.00105952
R16385 Iout.n673 Iout.n671 0.00105952
R16386 Iout.n676 Iout.n674 0.00105952
R16387 Iout.n679 Iout.n677 0.00105952
R16388 Iout.n682 Iout.n680 0.00105952
R16389 Iout.n685 Iout.n683 0.00105952
R16390 Iout.n959 Iout.n958 0.00105952
R16391 Iout.n694 Iout.n693 0.00105952
R16392 Iout.n697 Iout.n696 0.00105952
R16393 Iout.n691 Iout.n689 0.00105952
R16394 Iout.n688 Iout.n686 0.00105952
R16395 Iout.n962 Iout.n15 0.00105952
R16396 Iout.n965 Iout.n964 0.00105952
R16397 Iout.n575 Iout.n574 0.00105952
R16398 Iout.n578 Iout.n577 0.00105952
R16399 Iout.n587 Iout.n115 0.00105952
R16400 Iout.n590 Iout.n589 0.00105952
R16401 Iout.n599 Iout.n109 0.00105952
R16402 Iout.n602 Iout.n601 0.00105952
R16403 Iout.n611 Iout.n103 0.00105952
R16404 Iout.n614 Iout.n613 0.00105952
R16405 Iout.n623 Iout.n97 0.00105952
R16406 Iout.n626 Iout.n625 0.00105952
R16407 Iout.n86 Iout.n84 0.00105952
R16408 Iout.n644 Iout.n643 0.00105952
R16409 Iout.n641 Iout.n88 0.00105952
R16410 Iout.n632 Iout.n631 0.00105952
R16411 Iout.n629 Iout.n94 0.00105952
R16412 Iout.n620 Iout.n619 0.00105952
R16413 Iout.n617 Iout.n100 0.00105952
R16414 Iout.n608 Iout.n607 0.00105952
R16415 Iout.n605 Iout.n106 0.00105952
R16416 Iout.n596 Iout.n595 0.00105952
R16417 Iout.n593 Iout.n112 0.00105952
R16418 Iout.n584 Iout.n583 0.00105952
R16419 Iout.n973 Iout.n971 0.00105952
R16420 Iout.n970 Iout.n968 0.00105952
R16421 Iout.n565 Iout.n564 0.00105952
R16422 Iout.n581 Iout.n118 0.00105952
R16423 Iout.n978 Iout.n977 0.00105952
R16424 Iout.n122 Iout.n121 0.00105952
R16425 Iout.n568 Iout.n124 0.00105952
R16426 Iout.n571 Iout.n570 0.00105952
R16427 Iout.n335 Iout.n334 0.00105952
R16428 Iout.n338 Iout.n337 0.00105952
R16429 Iout.n341 Iout.n340 0.00105952
R16430 Iout.n344 Iout.n343 0.00105952
R16431 Iout.n347 Iout.n346 0.00105952
R16432 Iout.n350 Iout.n349 0.00105952
R16433 Iout.n353 Iout.n352 0.00105952
R16434 Iout.n356 Iout.n355 0.00105952
R16435 Iout.n359 Iout.n358 0.00105952
R16436 Iout.n372 Iout.n371 0.00105952
R16437 Iout.n385 Iout.n383 0.00105952
R16438 Iout.n388 Iout.n387 0.00105952
R16439 Iout.n401 Iout.n399 0.00105952
R16440 Iout.n404 Iout.n403 0.00105952
R16441 Iout.n417 Iout.n415 0.00105952
R16442 Iout.n420 Iout.n419 0.00105952
R16443 Iout.n433 Iout.n431 0.00105952
R16444 Iout.n443 Iout.n442 0.00105952
R16445 Iout.n440 Iout.n439 0.00105952
R16446 Iout.n437 Iout.n435 0.00105952
R16447 Iout.n555 Iout.n553 0.00105952
R16448 Iout.n558 Iout.n556 0.00105952
R16449 Iout.n981 Iout.n10 0.00105952
R16450 Iout.n984 Iout.n983 0.00105952
R16451 Iout.n561 Iout.n560 0.00105952
R16452 Iout.n992 Iout.n990 0.00105952
R16453 Iout.n989 Iout.n987 0.00105952
R16454 Iout.n129 Iout.n128 0.00105952
R16455 Iout.n547 Iout.n131 0.00105952
R16456 Iout.n550 Iout.n549 0.00105952
R16457 Iout.n451 Iout.n450 0.00105952
R16458 Iout.n454 Iout.n453 0.00105952
R16459 Iout.n448 Iout.n446 0.00105952
R16460 Iout.n428 Iout.n427 0.00105952
R16461 Iout.n425 Iout.n423 0.00105952
R16462 Iout.n412 Iout.n411 0.00105952
R16463 Iout.n409 Iout.n407 0.00105952
R16464 Iout.n396 Iout.n395 0.00105952
R16465 Iout.n393 Iout.n391 0.00105952
R16466 Iout.n331 Iout.n330 0.00105952
R16467 Iout.n328 Iout.n327 0.00105952
R16468 Iout.n325 Iout.n324 0.00105952
R16469 Iout.n322 Iout.n321 0.00105952
R16470 Iout.n319 Iout.n318 0.00105952
R16471 Iout.n316 Iout.n315 0.00105952
R16472 Iout.n313 Iout.n312 0.00105952
R16473 Iout.n310 Iout.n309 0.00105952
R16474 Iout.n307 Iout.n306 0.00105952
R16475 Iout.n459 Iout.n457 0.00105952
R16476 Iout.n465 Iout.n464 0.00105952
R16477 Iout.n462 Iout.n461 0.00105952
R16478 Iout.n544 Iout.n543 0.00105952
R16479 Iout.n541 Iout.n137 0.00105952
R16480 Iout.n997 Iout.n996 0.00105952
R16481 Iout.n135 Iout.n134 0.00105952
R16482 Iout.n1000 Iout.n5 0.00105952
R16483 Iout.n1003 Iout.n1002 0.00105952
R16484 Iout.n538 Iout.n537 0.00105952
R16485 Iout.n535 Iout.n533 0.00105952
R16486 Iout.n532 Iout.n530 0.00105952
R16487 Iout.n468 Iout.n157 0.00105952
R16488 Iout.n471 Iout.n470 0.00105952
R16489 Iout.n474 Iout.n473 0.00105952
R16490 Iout.n264 Iout.n190 0.00105952
R16491 Iout.n267 Iout.n266 0.00105952
R16492 Iout.n276 Iout.n184 0.00105952
R16493 Iout.n279 Iout.n278 0.00105952
R16494 Iout.n288 Iout.n178 0.00105952
R16495 Iout.n291 Iout.n290 0.00105952
R16496 Iout.n300 Iout.n169 0.00105952
R16497 Iout.n173 Iout.n171 0.00105952
R16498 Iout.n297 Iout.n296 0.00105952
R16499 Iout.n294 Iout.n175 0.00105952
R16500 Iout.n285 Iout.n284 0.00105952
R16501 Iout.n282 Iout.n181 0.00105952
R16502 Iout.n273 Iout.n272 0.00105952
R16503 Iout.n270 Iout.n187 0.00105952
R16504 Iout.n261 Iout.n260 0.00105952
R16505 Iout.n479 Iout.n477 0.00105952
R16506 Iout.n485 Iout.n484 0.00105952
R16507 Iout.n482 Iout.n481 0.00105952
R16508 Iout.n527 Iout.n526 0.00105952
R16509 Iout.n524 Iout.n144 0.00105952
R16510 Iout.n142 Iout.n141 0.00105952
R16511 Iout.n1008 Iout.n1006 0.00105952
R16512 Iout.n1011 Iout.n1009 0.00105952
R16513 Iout.n1016 Iout.n1015 0.00105952
R16514 Iout.n148 Iout.n147 0.00105952
R16515 Iout.n518 Iout.n150 0.00105952
R16516 Iout.n521 Iout.n520 0.00105952
R16517 Iout.n493 Iout.n492 0.00105952
R16518 Iout.n496 Iout.n495 0.00105952
R16519 Iout.n490 Iout.n488 0.00105952
R16520 Iout.n254 Iout.n253 0.00105952
R16521 Iout.n257 Iout.n256 0.00105952
R16522 Iout.n251 Iout.n249 0.00105952
R16523 Iout.n248 Iout.n246 0.00105952
R16524 Iout.n245 Iout.n243 0.00105952
R16525 Iout.n242 Iout.n240 0.00105952
R16526 Iout.n239 Iout.n237 0.00105952
R16527 Iout.n236 Iout.n234 0.00105952
R16528 Iout.n233 Iout.n231 0.00105952
R16529 Iout.n228 Iout.n227 0.00105952
R16530 Iout.n225 Iout.n223 0.00105952
R16531 Iout.n221 Iout.n219 0.00105952
R16532 Iout.n217 Iout.n215 0.00105952
R16533 Iout.n213 Iout.n211 0.00105952
R16534 Iout.n209 Iout.n207 0.00105952
R16535 Iout.n205 Iout.n203 0.00105952
R16536 Iout.n201 Iout.n200 0.00105952
R16537 Iout.n198 Iout.n196 0.00105952
R16538 Iout.n194 Iout.n193 0.00105952
R16539 Iout.n501 Iout.n499 0.00105952
R16540 Iout.n505 Iout.n503 0.00105952
R16541 Iout.n508 Iout.n506 0.00105952
R16542 Iout.n515 Iout.n514 0.00105952
R16543 Iout.n512 Iout.n510 0.00105952
R16544 Iout.n1021 Iout.n1019 0.00105952
R16545 XThC.Tn[10].n71 XThC.Tn[10].n70 256.104
R16546 XThC.Tn[10].n75 XThC.Tn[10].n74 243.679
R16547 XThC.Tn[10].n2 XThC.Tn[10].n0 241.847
R16548 XThC.Tn[10].n75 XThC.Tn[10].n73 205.28
R16549 XThC.Tn[10].n71 XThC.Tn[10].n69 202.095
R16550 XThC.Tn[10].n2 XThC.Tn[10].n1 185
R16551 XThC.Tn[10].n65 XThC.Tn[10].n63 161.365
R16552 XThC.Tn[10].n61 XThC.Tn[10].n59 161.365
R16553 XThC.Tn[10].n57 XThC.Tn[10].n55 161.365
R16554 XThC.Tn[10].n53 XThC.Tn[10].n51 161.365
R16555 XThC.Tn[10].n49 XThC.Tn[10].n47 161.365
R16556 XThC.Tn[10].n45 XThC.Tn[10].n43 161.365
R16557 XThC.Tn[10].n41 XThC.Tn[10].n39 161.365
R16558 XThC.Tn[10].n37 XThC.Tn[10].n35 161.365
R16559 XThC.Tn[10].n33 XThC.Tn[10].n31 161.365
R16560 XThC.Tn[10].n29 XThC.Tn[10].n27 161.365
R16561 XThC.Tn[10].n25 XThC.Tn[10].n23 161.365
R16562 XThC.Tn[10].n21 XThC.Tn[10].n19 161.365
R16563 XThC.Tn[10].n17 XThC.Tn[10].n15 161.365
R16564 XThC.Tn[10].n13 XThC.Tn[10].n11 161.365
R16565 XThC.Tn[10].n9 XThC.Tn[10].n7 161.365
R16566 XThC.Tn[10].n6 XThC.Tn[10].n4 161.365
R16567 XThC.Tn[10].n63 XThC.Tn[10].t42 161.202
R16568 XThC.Tn[10].n59 XThC.Tn[10].t32 161.202
R16569 XThC.Tn[10].n55 XThC.Tn[10].t19 161.202
R16570 XThC.Tn[10].n51 XThC.Tn[10].t16 161.202
R16571 XThC.Tn[10].n47 XThC.Tn[10].t40 161.202
R16572 XThC.Tn[10].n43 XThC.Tn[10].t27 161.202
R16573 XThC.Tn[10].n39 XThC.Tn[10].t26 161.202
R16574 XThC.Tn[10].n35 XThC.Tn[10].t39 161.202
R16575 XThC.Tn[10].n31 XThC.Tn[10].t37 161.202
R16576 XThC.Tn[10].n27 XThC.Tn[10].t28 161.202
R16577 XThC.Tn[10].n23 XThC.Tn[10].t15 161.202
R16578 XThC.Tn[10].n19 XThC.Tn[10].t14 161.202
R16579 XThC.Tn[10].n15 XThC.Tn[10].t25 161.202
R16580 XThC.Tn[10].n11 XThC.Tn[10].t23 161.202
R16581 XThC.Tn[10].n7 XThC.Tn[10].t21 161.202
R16582 XThC.Tn[10].n4 XThC.Tn[10].t36 161.202
R16583 XThC.Tn[10].n63 XThC.Tn[10].t13 145.137
R16584 XThC.Tn[10].n59 XThC.Tn[10].t35 145.137
R16585 XThC.Tn[10].n55 XThC.Tn[10].t22 145.137
R16586 XThC.Tn[10].n51 XThC.Tn[10].t20 145.137
R16587 XThC.Tn[10].n47 XThC.Tn[10].t12 145.137
R16588 XThC.Tn[10].n43 XThC.Tn[10].t33 145.137
R16589 XThC.Tn[10].n39 XThC.Tn[10].t31 145.137
R16590 XThC.Tn[10].n35 XThC.Tn[10].t43 145.137
R16591 XThC.Tn[10].n31 XThC.Tn[10].t41 145.137
R16592 XThC.Tn[10].n27 XThC.Tn[10].t34 145.137
R16593 XThC.Tn[10].n23 XThC.Tn[10].t18 145.137
R16594 XThC.Tn[10].n19 XThC.Tn[10].t17 145.137
R16595 XThC.Tn[10].n15 XThC.Tn[10].t30 145.137
R16596 XThC.Tn[10].n11 XThC.Tn[10].t29 145.137
R16597 XThC.Tn[10].n7 XThC.Tn[10].t24 145.137
R16598 XThC.Tn[10].n4 XThC.Tn[10].t38 145.137
R16599 XThC.Tn[10].n69 XThC.Tn[10].t6 26.5955
R16600 XThC.Tn[10].n69 XThC.Tn[10].t5 26.5955
R16601 XThC.Tn[10].n70 XThC.Tn[10].t10 26.5955
R16602 XThC.Tn[10].n70 XThC.Tn[10].t1 26.5955
R16603 XThC.Tn[10].n73 XThC.Tn[10].t4 26.5955
R16604 XThC.Tn[10].n73 XThC.Tn[10].t8 26.5955
R16605 XThC.Tn[10].n74 XThC.Tn[10].t0 26.5955
R16606 XThC.Tn[10].n74 XThC.Tn[10].t9 26.5955
R16607 XThC.Tn[10].n1 XThC.Tn[10].t11 24.9236
R16608 XThC.Tn[10].n1 XThC.Tn[10].t3 24.9236
R16609 XThC.Tn[10].n0 XThC.Tn[10].t2 24.9236
R16610 XThC.Tn[10].n0 XThC.Tn[10].t7 24.9236
R16611 XThC.Tn[10] XThC.Tn[10].n75 22.9652
R16612 XThC.Tn[10] XThC.Tn[10].n2 22.9615
R16613 XThC.Tn[10].n72 XThC.Tn[10].n71 13.9299
R16614 XThC.Tn[10] XThC.Tn[10].n72 13.9299
R16615 XThC.Tn[10] XThC.Tn[10].n6 8.0245
R16616 XThC.Tn[10].n66 XThC.Tn[10].n65 7.9105
R16617 XThC.Tn[10].n62 XThC.Tn[10].n61 7.9105
R16618 XThC.Tn[10].n58 XThC.Tn[10].n57 7.9105
R16619 XThC.Tn[10].n54 XThC.Tn[10].n53 7.9105
R16620 XThC.Tn[10].n50 XThC.Tn[10].n49 7.9105
R16621 XThC.Tn[10].n46 XThC.Tn[10].n45 7.9105
R16622 XThC.Tn[10].n42 XThC.Tn[10].n41 7.9105
R16623 XThC.Tn[10].n38 XThC.Tn[10].n37 7.9105
R16624 XThC.Tn[10].n34 XThC.Tn[10].n33 7.9105
R16625 XThC.Tn[10].n30 XThC.Tn[10].n29 7.9105
R16626 XThC.Tn[10].n26 XThC.Tn[10].n25 7.9105
R16627 XThC.Tn[10].n22 XThC.Tn[10].n21 7.9105
R16628 XThC.Tn[10].n18 XThC.Tn[10].n17 7.9105
R16629 XThC.Tn[10].n14 XThC.Tn[10].n13 7.9105
R16630 XThC.Tn[10].n10 XThC.Tn[10].n9 7.9105
R16631 XThC.Tn[10].n68 XThC.Tn[10].n67 7.40985
R16632 XThC.Tn[10].n67 XThC.Tn[10] 4.38575
R16633 XThC.Tn[10].n72 XThC.Tn[10].n68 2.99115
R16634 XThC.Tn[10].n72 XThC.Tn[10] 2.87153
R16635 XThC.Tn[10].n3 XThC.Tn[10] 2.688
R16636 XThC.Tn[10].n68 XThC.Tn[10] 2.2734
R16637 XThC.Tn[10].n67 XThC.Tn[10].n3 0.244922
R16638 XThC.Tn[10].n10 XThC.Tn[10] 0.235138
R16639 XThC.Tn[10].n14 XThC.Tn[10] 0.235138
R16640 XThC.Tn[10].n18 XThC.Tn[10] 0.235138
R16641 XThC.Tn[10].n22 XThC.Tn[10] 0.235138
R16642 XThC.Tn[10].n26 XThC.Tn[10] 0.235138
R16643 XThC.Tn[10].n30 XThC.Tn[10] 0.235138
R16644 XThC.Tn[10].n34 XThC.Tn[10] 0.235138
R16645 XThC.Tn[10].n38 XThC.Tn[10] 0.235138
R16646 XThC.Tn[10].n42 XThC.Tn[10] 0.235138
R16647 XThC.Tn[10].n46 XThC.Tn[10] 0.235138
R16648 XThC.Tn[10].n50 XThC.Tn[10] 0.235138
R16649 XThC.Tn[10].n54 XThC.Tn[10] 0.235138
R16650 XThC.Tn[10].n58 XThC.Tn[10] 0.235138
R16651 XThC.Tn[10].n62 XThC.Tn[10] 0.235138
R16652 XThC.Tn[10].n66 XThC.Tn[10] 0.235138
R16653 XThC.Tn[10].n3 XThC.Tn[10] 0.141947
R16654 XThC.Tn[10] XThC.Tn[10].n10 0.114505
R16655 XThC.Tn[10] XThC.Tn[10].n14 0.114505
R16656 XThC.Tn[10] XThC.Tn[10].n18 0.114505
R16657 XThC.Tn[10] XThC.Tn[10].n22 0.114505
R16658 XThC.Tn[10] XThC.Tn[10].n26 0.114505
R16659 XThC.Tn[10] XThC.Tn[10].n30 0.114505
R16660 XThC.Tn[10] XThC.Tn[10].n34 0.114505
R16661 XThC.Tn[10] XThC.Tn[10].n38 0.114505
R16662 XThC.Tn[10] XThC.Tn[10].n42 0.114505
R16663 XThC.Tn[10] XThC.Tn[10].n46 0.114505
R16664 XThC.Tn[10] XThC.Tn[10].n50 0.114505
R16665 XThC.Tn[10] XThC.Tn[10].n54 0.114505
R16666 XThC.Tn[10] XThC.Tn[10].n58 0.114505
R16667 XThC.Tn[10] XThC.Tn[10].n62 0.114505
R16668 XThC.Tn[10] XThC.Tn[10].n66 0.114505
R16669 XThC.Tn[10].n65 XThC.Tn[10].n64 0.0599512
R16670 XThC.Tn[10].n61 XThC.Tn[10].n60 0.0599512
R16671 XThC.Tn[10].n57 XThC.Tn[10].n56 0.0599512
R16672 XThC.Tn[10].n53 XThC.Tn[10].n52 0.0599512
R16673 XThC.Tn[10].n49 XThC.Tn[10].n48 0.0599512
R16674 XThC.Tn[10].n45 XThC.Tn[10].n44 0.0599512
R16675 XThC.Tn[10].n41 XThC.Tn[10].n40 0.0599512
R16676 XThC.Tn[10].n37 XThC.Tn[10].n36 0.0599512
R16677 XThC.Tn[10].n33 XThC.Tn[10].n32 0.0599512
R16678 XThC.Tn[10].n29 XThC.Tn[10].n28 0.0599512
R16679 XThC.Tn[10].n25 XThC.Tn[10].n24 0.0599512
R16680 XThC.Tn[10].n21 XThC.Tn[10].n20 0.0599512
R16681 XThC.Tn[10].n17 XThC.Tn[10].n16 0.0599512
R16682 XThC.Tn[10].n13 XThC.Tn[10].n12 0.0599512
R16683 XThC.Tn[10].n9 XThC.Tn[10].n8 0.0599512
R16684 XThC.Tn[10].n6 XThC.Tn[10].n5 0.0599512
R16685 XThC.Tn[10].n64 XThC.Tn[10] 0.0469286
R16686 XThC.Tn[10].n60 XThC.Tn[10] 0.0469286
R16687 XThC.Tn[10].n56 XThC.Tn[10] 0.0469286
R16688 XThC.Tn[10].n52 XThC.Tn[10] 0.0469286
R16689 XThC.Tn[10].n48 XThC.Tn[10] 0.0469286
R16690 XThC.Tn[10].n44 XThC.Tn[10] 0.0469286
R16691 XThC.Tn[10].n40 XThC.Tn[10] 0.0469286
R16692 XThC.Tn[10].n36 XThC.Tn[10] 0.0469286
R16693 XThC.Tn[10].n32 XThC.Tn[10] 0.0469286
R16694 XThC.Tn[10].n28 XThC.Tn[10] 0.0469286
R16695 XThC.Tn[10].n24 XThC.Tn[10] 0.0469286
R16696 XThC.Tn[10].n20 XThC.Tn[10] 0.0469286
R16697 XThC.Tn[10].n16 XThC.Tn[10] 0.0469286
R16698 XThC.Tn[10].n12 XThC.Tn[10] 0.0469286
R16699 XThC.Tn[10].n8 XThC.Tn[10] 0.0469286
R16700 XThC.Tn[10].n5 XThC.Tn[10] 0.0469286
R16701 XThC.Tn[10].n64 XThC.Tn[10] 0.0401341
R16702 XThC.Tn[10].n60 XThC.Tn[10] 0.0401341
R16703 XThC.Tn[10].n56 XThC.Tn[10] 0.0401341
R16704 XThC.Tn[10].n52 XThC.Tn[10] 0.0401341
R16705 XThC.Tn[10].n48 XThC.Tn[10] 0.0401341
R16706 XThC.Tn[10].n44 XThC.Tn[10] 0.0401341
R16707 XThC.Tn[10].n40 XThC.Tn[10] 0.0401341
R16708 XThC.Tn[10].n36 XThC.Tn[10] 0.0401341
R16709 XThC.Tn[10].n32 XThC.Tn[10] 0.0401341
R16710 XThC.Tn[10].n28 XThC.Tn[10] 0.0401341
R16711 XThC.Tn[10].n24 XThC.Tn[10] 0.0401341
R16712 XThC.Tn[10].n20 XThC.Tn[10] 0.0401341
R16713 XThC.Tn[10].n16 XThC.Tn[10] 0.0401341
R16714 XThC.Tn[10].n12 XThC.Tn[10] 0.0401341
R16715 XThC.Tn[10].n8 XThC.Tn[10] 0.0401341
R16716 XThC.Tn[10].n5 XThC.Tn[10] 0.0401341
R16717 XThR.Tn[6].n2 XThR.Tn[6].n1 332.332
R16718 XThR.Tn[6].n2 XThR.Tn[6].n0 296.493
R16719 XThR.Tn[6] XThR.Tn[6].n82 161.363
R16720 XThR.Tn[6] XThR.Tn[6].n77 161.363
R16721 XThR.Tn[6] XThR.Tn[6].n72 161.363
R16722 XThR.Tn[6] XThR.Tn[6].n67 161.363
R16723 XThR.Tn[6] XThR.Tn[6].n62 161.363
R16724 XThR.Tn[6] XThR.Tn[6].n57 161.363
R16725 XThR.Tn[6] XThR.Tn[6].n52 161.363
R16726 XThR.Tn[6] XThR.Tn[6].n47 161.363
R16727 XThR.Tn[6] XThR.Tn[6].n42 161.363
R16728 XThR.Tn[6] XThR.Tn[6].n37 161.363
R16729 XThR.Tn[6] XThR.Tn[6].n32 161.363
R16730 XThR.Tn[6] XThR.Tn[6].n27 161.363
R16731 XThR.Tn[6] XThR.Tn[6].n22 161.363
R16732 XThR.Tn[6] XThR.Tn[6].n17 161.363
R16733 XThR.Tn[6] XThR.Tn[6].n12 161.363
R16734 XThR.Tn[6] XThR.Tn[6].n10 161.363
R16735 XThR.Tn[6].n84 XThR.Tn[6].n83 161.3
R16736 XThR.Tn[6].n79 XThR.Tn[6].n78 161.3
R16737 XThR.Tn[6].n74 XThR.Tn[6].n73 161.3
R16738 XThR.Tn[6].n69 XThR.Tn[6].n68 161.3
R16739 XThR.Tn[6].n64 XThR.Tn[6].n63 161.3
R16740 XThR.Tn[6].n59 XThR.Tn[6].n58 161.3
R16741 XThR.Tn[6].n54 XThR.Tn[6].n53 161.3
R16742 XThR.Tn[6].n49 XThR.Tn[6].n48 161.3
R16743 XThR.Tn[6].n44 XThR.Tn[6].n43 161.3
R16744 XThR.Tn[6].n39 XThR.Tn[6].n38 161.3
R16745 XThR.Tn[6].n34 XThR.Tn[6].n33 161.3
R16746 XThR.Tn[6].n29 XThR.Tn[6].n28 161.3
R16747 XThR.Tn[6].n24 XThR.Tn[6].n23 161.3
R16748 XThR.Tn[6].n19 XThR.Tn[6].n18 161.3
R16749 XThR.Tn[6].n14 XThR.Tn[6].n13 161.3
R16750 XThR.Tn[6].n82 XThR.Tn[6].t46 161.106
R16751 XThR.Tn[6].n77 XThR.Tn[6].t52 161.106
R16752 XThR.Tn[6].n72 XThR.Tn[6].t32 161.106
R16753 XThR.Tn[6].n67 XThR.Tn[6].t18 161.106
R16754 XThR.Tn[6].n62 XThR.Tn[6].t44 161.106
R16755 XThR.Tn[6].n57 XThR.Tn[6].t69 161.106
R16756 XThR.Tn[6].n52 XThR.Tn[6].t50 161.106
R16757 XThR.Tn[6].n47 XThR.Tn[6].t30 161.106
R16758 XThR.Tn[6].n42 XThR.Tn[6].t17 161.106
R16759 XThR.Tn[6].n37 XThR.Tn[6].t22 161.106
R16760 XThR.Tn[6].n32 XThR.Tn[6].t67 161.106
R16761 XThR.Tn[6].n27 XThR.Tn[6].t31 161.106
R16762 XThR.Tn[6].n22 XThR.Tn[6].t66 161.106
R16763 XThR.Tn[6].n17 XThR.Tn[6].t49 161.106
R16764 XThR.Tn[6].n12 XThR.Tn[6].t72 161.106
R16765 XThR.Tn[6].n10 XThR.Tn[6].t56 161.106
R16766 XThR.Tn[6].n83 XThR.Tn[6].t42 159.978
R16767 XThR.Tn[6].n78 XThR.Tn[6].t48 159.978
R16768 XThR.Tn[6].n73 XThR.Tn[6].t28 159.978
R16769 XThR.Tn[6].n68 XThR.Tn[6].t15 159.978
R16770 XThR.Tn[6].n63 XThR.Tn[6].t39 159.978
R16771 XThR.Tn[6].n58 XThR.Tn[6].t65 159.978
R16772 XThR.Tn[6].n53 XThR.Tn[6].t47 159.978
R16773 XThR.Tn[6].n48 XThR.Tn[6].t25 159.978
R16774 XThR.Tn[6].n43 XThR.Tn[6].t12 159.978
R16775 XThR.Tn[6].n38 XThR.Tn[6].t19 159.978
R16776 XThR.Tn[6].n33 XThR.Tn[6].t64 159.978
R16777 XThR.Tn[6].n28 XThR.Tn[6].t27 159.978
R16778 XThR.Tn[6].n23 XThR.Tn[6].t63 159.978
R16779 XThR.Tn[6].n18 XThR.Tn[6].t45 159.978
R16780 XThR.Tn[6].n13 XThR.Tn[6].t68 159.978
R16781 XThR.Tn[6].n82 XThR.Tn[6].t34 145.038
R16782 XThR.Tn[6].n77 XThR.Tn[6].t58 145.038
R16783 XThR.Tn[6].n72 XThR.Tn[6].t38 145.038
R16784 XThR.Tn[6].n67 XThR.Tn[6].t23 145.038
R16785 XThR.Tn[6].n62 XThR.Tn[6].t53 145.038
R16786 XThR.Tn[6].n57 XThR.Tn[6].t33 145.038
R16787 XThR.Tn[6].n52 XThR.Tn[6].t40 145.038
R16788 XThR.Tn[6].n47 XThR.Tn[6].t24 145.038
R16789 XThR.Tn[6].n42 XThR.Tn[6].t21 145.038
R16790 XThR.Tn[6].n37 XThR.Tn[6].t51 145.038
R16791 XThR.Tn[6].n32 XThR.Tn[6].t13 145.038
R16792 XThR.Tn[6].n27 XThR.Tn[6].t35 145.038
R16793 XThR.Tn[6].n22 XThR.Tn[6].t73 145.038
R16794 XThR.Tn[6].n17 XThR.Tn[6].t57 145.038
R16795 XThR.Tn[6].n12 XThR.Tn[6].t20 145.038
R16796 XThR.Tn[6].n10 XThR.Tn[6].t62 145.038
R16797 XThR.Tn[6].n83 XThR.Tn[6].t55 143.911
R16798 XThR.Tn[6].n78 XThR.Tn[6].t16 143.911
R16799 XThR.Tn[6].n73 XThR.Tn[6].t60 143.911
R16800 XThR.Tn[6].n68 XThR.Tn[6].t41 143.911
R16801 XThR.Tn[6].n63 XThR.Tn[6].t71 143.911
R16802 XThR.Tn[6].n58 XThR.Tn[6].t54 143.911
R16803 XThR.Tn[6].n53 XThR.Tn[6].t61 143.911
R16804 XThR.Tn[6].n48 XThR.Tn[6].t43 143.911
R16805 XThR.Tn[6].n43 XThR.Tn[6].t37 143.911
R16806 XThR.Tn[6].n38 XThR.Tn[6].t70 143.911
R16807 XThR.Tn[6].n33 XThR.Tn[6].t29 143.911
R16808 XThR.Tn[6].n28 XThR.Tn[6].t59 143.911
R16809 XThR.Tn[6].n23 XThR.Tn[6].t26 143.911
R16810 XThR.Tn[6].n18 XThR.Tn[6].t14 143.911
R16811 XThR.Tn[6].n13 XThR.Tn[6].t36 143.911
R16812 XThR.Tn[6].n7 XThR.Tn[6].n5 135.249
R16813 XThR.Tn[6].n9 XThR.Tn[6].n3 98.982
R16814 XThR.Tn[6].n8 XThR.Tn[6].n4 98.982
R16815 XThR.Tn[6].n7 XThR.Tn[6].n6 98.982
R16816 XThR.Tn[6].n9 XThR.Tn[6].n8 36.2672
R16817 XThR.Tn[6].n8 XThR.Tn[6].n7 36.2672
R16818 XThR.Tn[6].n88 XThR.Tn[6].n9 32.6405
R16819 XThR.Tn[6].n1 XThR.Tn[6].t6 26.5955
R16820 XThR.Tn[6].n1 XThR.Tn[6].t5 26.5955
R16821 XThR.Tn[6].n0 XThR.Tn[6].t7 26.5955
R16822 XThR.Tn[6].n0 XThR.Tn[6].t4 26.5955
R16823 XThR.Tn[6].n3 XThR.Tn[6].t8 24.9236
R16824 XThR.Tn[6].n3 XThR.Tn[6].t9 24.9236
R16825 XThR.Tn[6].n4 XThR.Tn[6].t11 24.9236
R16826 XThR.Tn[6].n4 XThR.Tn[6].t10 24.9236
R16827 XThR.Tn[6].n5 XThR.Tn[6].t0 24.9236
R16828 XThR.Tn[6].n5 XThR.Tn[6].t1 24.9236
R16829 XThR.Tn[6].n6 XThR.Tn[6].t3 24.9236
R16830 XThR.Tn[6].n6 XThR.Tn[6].t2 24.9236
R16831 XThR.Tn[6] XThR.Tn[6].n2 23.3605
R16832 XThR.Tn[6] XThR.Tn[6].n88 6.7205
R16833 XThR.Tn[6].n88 XThR.Tn[6] 5.37828
R16834 XThR.Tn[6] XThR.Tn[6].n11 5.34038
R16835 XThR.Tn[6].n16 XThR.Tn[6].n15 4.5005
R16836 XThR.Tn[6].n21 XThR.Tn[6].n20 4.5005
R16837 XThR.Tn[6].n26 XThR.Tn[6].n25 4.5005
R16838 XThR.Tn[6].n31 XThR.Tn[6].n30 4.5005
R16839 XThR.Tn[6].n36 XThR.Tn[6].n35 4.5005
R16840 XThR.Tn[6].n41 XThR.Tn[6].n40 4.5005
R16841 XThR.Tn[6].n46 XThR.Tn[6].n45 4.5005
R16842 XThR.Tn[6].n51 XThR.Tn[6].n50 4.5005
R16843 XThR.Tn[6].n56 XThR.Tn[6].n55 4.5005
R16844 XThR.Tn[6].n61 XThR.Tn[6].n60 4.5005
R16845 XThR.Tn[6].n66 XThR.Tn[6].n65 4.5005
R16846 XThR.Tn[6].n71 XThR.Tn[6].n70 4.5005
R16847 XThR.Tn[6].n76 XThR.Tn[6].n75 4.5005
R16848 XThR.Tn[6].n81 XThR.Tn[6].n80 4.5005
R16849 XThR.Tn[6].n86 XThR.Tn[6].n85 4.5005
R16850 XThR.Tn[6].n87 XThR.Tn[6] 3.70586
R16851 XThR.Tn[6].n16 XThR.Tn[6] 2.52282
R16852 XThR.Tn[6].n21 XThR.Tn[6] 2.52282
R16853 XThR.Tn[6].n26 XThR.Tn[6] 2.52282
R16854 XThR.Tn[6].n31 XThR.Tn[6] 2.52282
R16855 XThR.Tn[6].n36 XThR.Tn[6] 2.52282
R16856 XThR.Tn[6].n41 XThR.Tn[6] 2.52282
R16857 XThR.Tn[6].n46 XThR.Tn[6] 2.52282
R16858 XThR.Tn[6].n51 XThR.Tn[6] 2.52282
R16859 XThR.Tn[6].n56 XThR.Tn[6] 2.52282
R16860 XThR.Tn[6].n61 XThR.Tn[6] 2.52282
R16861 XThR.Tn[6].n66 XThR.Tn[6] 2.52282
R16862 XThR.Tn[6].n71 XThR.Tn[6] 2.52282
R16863 XThR.Tn[6].n76 XThR.Tn[6] 2.52282
R16864 XThR.Tn[6].n81 XThR.Tn[6] 2.52282
R16865 XThR.Tn[6].n86 XThR.Tn[6] 2.52282
R16866 XThR.Tn[6].n84 XThR.Tn[6] 1.08677
R16867 XThR.Tn[6].n79 XThR.Tn[6] 1.08677
R16868 XThR.Tn[6].n74 XThR.Tn[6] 1.08677
R16869 XThR.Tn[6].n69 XThR.Tn[6] 1.08677
R16870 XThR.Tn[6].n64 XThR.Tn[6] 1.08677
R16871 XThR.Tn[6].n59 XThR.Tn[6] 1.08677
R16872 XThR.Tn[6].n54 XThR.Tn[6] 1.08677
R16873 XThR.Tn[6].n49 XThR.Tn[6] 1.08677
R16874 XThR.Tn[6].n44 XThR.Tn[6] 1.08677
R16875 XThR.Tn[6].n39 XThR.Tn[6] 1.08677
R16876 XThR.Tn[6].n34 XThR.Tn[6] 1.08677
R16877 XThR.Tn[6].n29 XThR.Tn[6] 1.08677
R16878 XThR.Tn[6].n24 XThR.Tn[6] 1.08677
R16879 XThR.Tn[6].n19 XThR.Tn[6] 1.08677
R16880 XThR.Tn[6].n14 XThR.Tn[6] 1.08677
R16881 XThR.Tn[6] XThR.Tn[6].n16 0.839786
R16882 XThR.Tn[6] XThR.Tn[6].n21 0.839786
R16883 XThR.Tn[6] XThR.Tn[6].n26 0.839786
R16884 XThR.Tn[6] XThR.Tn[6].n31 0.839786
R16885 XThR.Tn[6] XThR.Tn[6].n36 0.839786
R16886 XThR.Tn[6] XThR.Tn[6].n41 0.839786
R16887 XThR.Tn[6] XThR.Tn[6].n46 0.839786
R16888 XThR.Tn[6] XThR.Tn[6].n51 0.839786
R16889 XThR.Tn[6] XThR.Tn[6].n56 0.839786
R16890 XThR.Tn[6] XThR.Tn[6].n61 0.839786
R16891 XThR.Tn[6] XThR.Tn[6].n66 0.839786
R16892 XThR.Tn[6] XThR.Tn[6].n71 0.839786
R16893 XThR.Tn[6] XThR.Tn[6].n76 0.839786
R16894 XThR.Tn[6] XThR.Tn[6].n81 0.839786
R16895 XThR.Tn[6] XThR.Tn[6].n86 0.839786
R16896 XThR.Tn[6].n11 XThR.Tn[6] 0.499542
R16897 XThR.Tn[6].n85 XThR.Tn[6] 0.063
R16898 XThR.Tn[6].n80 XThR.Tn[6] 0.063
R16899 XThR.Tn[6].n75 XThR.Tn[6] 0.063
R16900 XThR.Tn[6].n70 XThR.Tn[6] 0.063
R16901 XThR.Tn[6].n65 XThR.Tn[6] 0.063
R16902 XThR.Tn[6].n60 XThR.Tn[6] 0.063
R16903 XThR.Tn[6].n55 XThR.Tn[6] 0.063
R16904 XThR.Tn[6].n50 XThR.Tn[6] 0.063
R16905 XThR.Tn[6].n45 XThR.Tn[6] 0.063
R16906 XThR.Tn[6].n40 XThR.Tn[6] 0.063
R16907 XThR.Tn[6].n35 XThR.Tn[6] 0.063
R16908 XThR.Tn[6].n30 XThR.Tn[6] 0.063
R16909 XThR.Tn[6].n25 XThR.Tn[6] 0.063
R16910 XThR.Tn[6].n20 XThR.Tn[6] 0.063
R16911 XThR.Tn[6].n15 XThR.Tn[6] 0.063
R16912 XThR.Tn[6].n87 XThR.Tn[6] 0.0540714
R16913 XThR.Tn[6] XThR.Tn[6].n87 0.038
R16914 XThR.Tn[6].n11 XThR.Tn[6] 0.0143889
R16915 XThR.Tn[6].n85 XThR.Tn[6].n84 0.00771154
R16916 XThR.Tn[6].n80 XThR.Tn[6].n79 0.00771154
R16917 XThR.Tn[6].n75 XThR.Tn[6].n74 0.00771154
R16918 XThR.Tn[6].n70 XThR.Tn[6].n69 0.00771154
R16919 XThR.Tn[6].n65 XThR.Tn[6].n64 0.00771154
R16920 XThR.Tn[6].n60 XThR.Tn[6].n59 0.00771154
R16921 XThR.Tn[6].n55 XThR.Tn[6].n54 0.00771154
R16922 XThR.Tn[6].n50 XThR.Tn[6].n49 0.00771154
R16923 XThR.Tn[6].n45 XThR.Tn[6].n44 0.00771154
R16924 XThR.Tn[6].n40 XThR.Tn[6].n39 0.00771154
R16925 XThR.Tn[6].n35 XThR.Tn[6].n34 0.00771154
R16926 XThR.Tn[6].n30 XThR.Tn[6].n29 0.00771154
R16927 XThR.Tn[6].n25 XThR.Tn[6].n24 0.00771154
R16928 XThR.Tn[6].n20 XThR.Tn[6].n19 0.00771154
R16929 XThR.Tn[6].n15 XThR.Tn[6].n14 0.00771154
R16930 XThR.Tn[14].n87 XThR.Tn[14].n86 256.103
R16931 XThR.Tn[14].n2 XThR.Tn[14].n0 243.68
R16932 XThR.Tn[14].n5 XThR.Tn[14].n3 241.847
R16933 XThR.Tn[14].n2 XThR.Tn[14].n1 205.28
R16934 XThR.Tn[14].n87 XThR.Tn[14].n85 202.094
R16935 XThR.Tn[14].n5 XThR.Tn[14].n4 185
R16936 XThR.Tn[14] XThR.Tn[14].n78 161.363
R16937 XThR.Tn[14] XThR.Tn[14].n73 161.363
R16938 XThR.Tn[14] XThR.Tn[14].n68 161.363
R16939 XThR.Tn[14] XThR.Tn[14].n63 161.363
R16940 XThR.Tn[14] XThR.Tn[14].n58 161.363
R16941 XThR.Tn[14] XThR.Tn[14].n53 161.363
R16942 XThR.Tn[14] XThR.Tn[14].n48 161.363
R16943 XThR.Tn[14] XThR.Tn[14].n43 161.363
R16944 XThR.Tn[14] XThR.Tn[14].n38 161.363
R16945 XThR.Tn[14] XThR.Tn[14].n33 161.363
R16946 XThR.Tn[14] XThR.Tn[14].n28 161.363
R16947 XThR.Tn[14] XThR.Tn[14].n23 161.363
R16948 XThR.Tn[14] XThR.Tn[14].n18 161.363
R16949 XThR.Tn[14] XThR.Tn[14].n13 161.363
R16950 XThR.Tn[14] XThR.Tn[14].n8 161.363
R16951 XThR.Tn[14] XThR.Tn[14].n6 161.363
R16952 XThR.Tn[14].n80 XThR.Tn[14].n79 161.3
R16953 XThR.Tn[14].n75 XThR.Tn[14].n74 161.3
R16954 XThR.Tn[14].n70 XThR.Tn[14].n69 161.3
R16955 XThR.Tn[14].n65 XThR.Tn[14].n64 161.3
R16956 XThR.Tn[14].n60 XThR.Tn[14].n59 161.3
R16957 XThR.Tn[14].n55 XThR.Tn[14].n54 161.3
R16958 XThR.Tn[14].n50 XThR.Tn[14].n49 161.3
R16959 XThR.Tn[14].n45 XThR.Tn[14].n44 161.3
R16960 XThR.Tn[14].n40 XThR.Tn[14].n39 161.3
R16961 XThR.Tn[14].n35 XThR.Tn[14].n34 161.3
R16962 XThR.Tn[14].n30 XThR.Tn[14].n29 161.3
R16963 XThR.Tn[14].n25 XThR.Tn[14].n24 161.3
R16964 XThR.Tn[14].n20 XThR.Tn[14].n19 161.3
R16965 XThR.Tn[14].n15 XThR.Tn[14].n14 161.3
R16966 XThR.Tn[14].n10 XThR.Tn[14].n9 161.3
R16967 XThR.Tn[14].n78 XThR.Tn[14].t51 161.106
R16968 XThR.Tn[14].n73 XThR.Tn[14].t58 161.106
R16969 XThR.Tn[14].n68 XThR.Tn[14].t39 161.106
R16970 XThR.Tn[14].n63 XThR.Tn[14].t22 161.106
R16971 XThR.Tn[14].n58 XThR.Tn[14].t49 161.106
R16972 XThR.Tn[14].n53 XThR.Tn[14].t12 161.106
R16973 XThR.Tn[14].n48 XThR.Tn[14].t56 161.106
R16974 XThR.Tn[14].n43 XThR.Tn[14].t36 161.106
R16975 XThR.Tn[14].n38 XThR.Tn[14].t19 161.106
R16976 XThR.Tn[14].n33 XThR.Tn[14].t25 161.106
R16977 XThR.Tn[14].n28 XThR.Tn[14].t73 161.106
R16978 XThR.Tn[14].n23 XThR.Tn[14].t38 161.106
R16979 XThR.Tn[14].n18 XThR.Tn[14].t72 161.106
R16980 XThR.Tn[14].n13 XThR.Tn[14].t54 161.106
R16981 XThR.Tn[14].n8 XThR.Tn[14].t13 161.106
R16982 XThR.Tn[14].n6 XThR.Tn[14].t62 161.106
R16983 XThR.Tn[14].n79 XThR.Tn[14].t32 159.978
R16984 XThR.Tn[14].n74 XThR.Tn[14].t37 159.978
R16985 XThR.Tn[14].n69 XThR.Tn[14].t20 159.978
R16986 XThR.Tn[14].n64 XThR.Tn[14].t68 159.978
R16987 XThR.Tn[14].n59 XThR.Tn[14].t30 159.978
R16988 XThR.Tn[14].n54 XThR.Tn[14].t55 159.978
R16989 XThR.Tn[14].n49 XThR.Tn[14].t35 159.978
R16990 XThR.Tn[14].n44 XThR.Tn[14].t16 159.978
R16991 XThR.Tn[14].n39 XThR.Tn[14].t66 159.978
R16992 XThR.Tn[14].n34 XThR.Tn[14].t71 159.978
R16993 XThR.Tn[14].n29 XThR.Tn[14].t53 159.978
R16994 XThR.Tn[14].n24 XThR.Tn[14].t18 159.978
R16995 XThR.Tn[14].n19 XThR.Tn[14].t52 159.978
R16996 XThR.Tn[14].n14 XThR.Tn[14].t34 159.978
R16997 XThR.Tn[14].n9 XThR.Tn[14].t60 159.978
R16998 XThR.Tn[14].n78 XThR.Tn[14].t41 145.038
R16999 XThR.Tn[14].n73 XThR.Tn[14].t65 145.038
R17000 XThR.Tn[14].n68 XThR.Tn[14].t45 145.038
R17001 XThR.Tn[14].n63 XThR.Tn[14].t26 145.038
R17002 XThR.Tn[14].n58 XThR.Tn[14].t59 145.038
R17003 XThR.Tn[14].n53 XThR.Tn[14].t40 145.038
R17004 XThR.Tn[14].n48 XThR.Tn[14].t46 145.038
R17005 XThR.Tn[14].n43 XThR.Tn[14].t27 145.038
R17006 XThR.Tn[14].n38 XThR.Tn[14].t23 145.038
R17007 XThR.Tn[14].n33 XThR.Tn[14].t57 145.038
R17008 XThR.Tn[14].n28 XThR.Tn[14].t15 145.038
R17009 XThR.Tn[14].n23 XThR.Tn[14].t44 145.038
R17010 XThR.Tn[14].n18 XThR.Tn[14].t14 145.038
R17011 XThR.Tn[14].n13 XThR.Tn[14].t64 145.038
R17012 XThR.Tn[14].n8 XThR.Tn[14].t24 145.038
R17013 XThR.Tn[14].n6 XThR.Tn[14].t69 145.038
R17014 XThR.Tn[14].n79 XThR.Tn[14].t43 143.911
R17015 XThR.Tn[14].n74 XThR.Tn[14].t70 143.911
R17016 XThR.Tn[14].n69 XThR.Tn[14].t48 143.911
R17017 XThR.Tn[14].n64 XThR.Tn[14].t31 143.911
R17018 XThR.Tn[14].n59 XThR.Tn[14].t63 143.911
R17019 XThR.Tn[14].n54 XThR.Tn[14].t42 143.911
R17020 XThR.Tn[14].n49 XThR.Tn[14].t50 143.911
R17021 XThR.Tn[14].n44 XThR.Tn[14].t33 143.911
R17022 XThR.Tn[14].n39 XThR.Tn[14].t29 143.911
R17023 XThR.Tn[14].n34 XThR.Tn[14].t61 143.911
R17024 XThR.Tn[14].n29 XThR.Tn[14].t21 143.911
R17025 XThR.Tn[14].n24 XThR.Tn[14].t47 143.911
R17026 XThR.Tn[14].n19 XThR.Tn[14].t17 143.911
R17027 XThR.Tn[14].n14 XThR.Tn[14].t67 143.911
R17028 XThR.Tn[14].n9 XThR.Tn[14].t28 143.911
R17029 XThR.Tn[14] XThR.Tn[14].n2 35.7652
R17030 XThR.Tn[14].n86 XThR.Tn[14].t0 26.5955
R17031 XThR.Tn[14].n86 XThR.Tn[14].t1 26.5955
R17032 XThR.Tn[14].n0 XThR.Tn[14].t8 26.5955
R17033 XThR.Tn[14].n0 XThR.Tn[14].t9 26.5955
R17034 XThR.Tn[14].n1 XThR.Tn[14].t10 26.5955
R17035 XThR.Tn[14].n1 XThR.Tn[14].t11 26.5955
R17036 XThR.Tn[14].n85 XThR.Tn[14].t2 26.5955
R17037 XThR.Tn[14].n85 XThR.Tn[14].t3 26.5955
R17038 XThR.Tn[14].n4 XThR.Tn[14].t4 24.9236
R17039 XThR.Tn[14].n4 XThR.Tn[14].t5 24.9236
R17040 XThR.Tn[14].n3 XThR.Tn[14].t6 24.9236
R17041 XThR.Tn[14].n3 XThR.Tn[14].t7 24.9236
R17042 XThR.Tn[14] XThR.Tn[14].n5 18.8943
R17043 XThR.Tn[14].n88 XThR.Tn[14].n87 13.5534
R17044 XThR.Tn[14].n84 XThR.Tn[14] 8.47191
R17045 XThR.Tn[14].n84 XThR.Tn[14] 6.34069
R17046 XThR.Tn[14] XThR.Tn[14].n7 5.34038
R17047 XThR.Tn[14].n12 XThR.Tn[14].n11 4.5005
R17048 XThR.Tn[14].n17 XThR.Tn[14].n16 4.5005
R17049 XThR.Tn[14].n22 XThR.Tn[14].n21 4.5005
R17050 XThR.Tn[14].n27 XThR.Tn[14].n26 4.5005
R17051 XThR.Tn[14].n32 XThR.Tn[14].n31 4.5005
R17052 XThR.Tn[14].n37 XThR.Tn[14].n36 4.5005
R17053 XThR.Tn[14].n42 XThR.Tn[14].n41 4.5005
R17054 XThR.Tn[14].n47 XThR.Tn[14].n46 4.5005
R17055 XThR.Tn[14].n52 XThR.Tn[14].n51 4.5005
R17056 XThR.Tn[14].n57 XThR.Tn[14].n56 4.5005
R17057 XThR.Tn[14].n62 XThR.Tn[14].n61 4.5005
R17058 XThR.Tn[14].n67 XThR.Tn[14].n66 4.5005
R17059 XThR.Tn[14].n72 XThR.Tn[14].n71 4.5005
R17060 XThR.Tn[14].n77 XThR.Tn[14].n76 4.5005
R17061 XThR.Tn[14].n82 XThR.Tn[14].n81 4.5005
R17062 XThR.Tn[14].n83 XThR.Tn[14] 3.70586
R17063 XThR.Tn[14].n12 XThR.Tn[14] 2.52282
R17064 XThR.Tn[14].n17 XThR.Tn[14] 2.52282
R17065 XThR.Tn[14].n22 XThR.Tn[14] 2.52282
R17066 XThR.Tn[14].n27 XThR.Tn[14] 2.52282
R17067 XThR.Tn[14].n32 XThR.Tn[14] 2.52282
R17068 XThR.Tn[14].n37 XThR.Tn[14] 2.52282
R17069 XThR.Tn[14].n42 XThR.Tn[14] 2.52282
R17070 XThR.Tn[14].n47 XThR.Tn[14] 2.52282
R17071 XThR.Tn[14].n52 XThR.Tn[14] 2.52282
R17072 XThR.Tn[14].n57 XThR.Tn[14] 2.52282
R17073 XThR.Tn[14].n62 XThR.Tn[14] 2.52282
R17074 XThR.Tn[14].n67 XThR.Tn[14] 2.52282
R17075 XThR.Tn[14].n72 XThR.Tn[14] 2.52282
R17076 XThR.Tn[14].n77 XThR.Tn[14] 2.52282
R17077 XThR.Tn[14].n82 XThR.Tn[14] 2.52282
R17078 XThR.Tn[14] XThR.Tn[14].n84 1.79489
R17079 XThR.Tn[14] XThR.Tn[14].n88 1.50638
R17080 XThR.Tn[14].n88 XThR.Tn[14] 1.19676
R17081 XThR.Tn[14].n80 XThR.Tn[14] 1.08677
R17082 XThR.Tn[14].n75 XThR.Tn[14] 1.08677
R17083 XThR.Tn[14].n70 XThR.Tn[14] 1.08677
R17084 XThR.Tn[14].n65 XThR.Tn[14] 1.08677
R17085 XThR.Tn[14].n60 XThR.Tn[14] 1.08677
R17086 XThR.Tn[14].n55 XThR.Tn[14] 1.08677
R17087 XThR.Tn[14].n50 XThR.Tn[14] 1.08677
R17088 XThR.Tn[14].n45 XThR.Tn[14] 1.08677
R17089 XThR.Tn[14].n40 XThR.Tn[14] 1.08677
R17090 XThR.Tn[14].n35 XThR.Tn[14] 1.08677
R17091 XThR.Tn[14].n30 XThR.Tn[14] 1.08677
R17092 XThR.Tn[14].n25 XThR.Tn[14] 1.08677
R17093 XThR.Tn[14].n20 XThR.Tn[14] 1.08677
R17094 XThR.Tn[14].n15 XThR.Tn[14] 1.08677
R17095 XThR.Tn[14].n10 XThR.Tn[14] 1.08677
R17096 XThR.Tn[14] XThR.Tn[14].n12 0.839786
R17097 XThR.Tn[14] XThR.Tn[14].n17 0.839786
R17098 XThR.Tn[14] XThR.Tn[14].n22 0.839786
R17099 XThR.Tn[14] XThR.Tn[14].n27 0.839786
R17100 XThR.Tn[14] XThR.Tn[14].n32 0.839786
R17101 XThR.Tn[14] XThR.Tn[14].n37 0.839786
R17102 XThR.Tn[14] XThR.Tn[14].n42 0.839786
R17103 XThR.Tn[14] XThR.Tn[14].n47 0.839786
R17104 XThR.Tn[14] XThR.Tn[14].n52 0.839786
R17105 XThR.Tn[14] XThR.Tn[14].n57 0.839786
R17106 XThR.Tn[14] XThR.Tn[14].n62 0.839786
R17107 XThR.Tn[14] XThR.Tn[14].n67 0.839786
R17108 XThR.Tn[14] XThR.Tn[14].n72 0.839786
R17109 XThR.Tn[14] XThR.Tn[14].n77 0.839786
R17110 XThR.Tn[14] XThR.Tn[14].n82 0.839786
R17111 XThR.Tn[14].n7 XThR.Tn[14] 0.499542
R17112 XThR.Tn[14].n81 XThR.Tn[14] 0.063
R17113 XThR.Tn[14].n76 XThR.Tn[14] 0.063
R17114 XThR.Tn[14].n71 XThR.Tn[14] 0.063
R17115 XThR.Tn[14].n66 XThR.Tn[14] 0.063
R17116 XThR.Tn[14].n61 XThR.Tn[14] 0.063
R17117 XThR.Tn[14].n56 XThR.Tn[14] 0.063
R17118 XThR.Tn[14].n51 XThR.Tn[14] 0.063
R17119 XThR.Tn[14].n46 XThR.Tn[14] 0.063
R17120 XThR.Tn[14].n41 XThR.Tn[14] 0.063
R17121 XThR.Tn[14].n36 XThR.Tn[14] 0.063
R17122 XThR.Tn[14].n31 XThR.Tn[14] 0.063
R17123 XThR.Tn[14].n26 XThR.Tn[14] 0.063
R17124 XThR.Tn[14].n21 XThR.Tn[14] 0.063
R17125 XThR.Tn[14].n16 XThR.Tn[14] 0.063
R17126 XThR.Tn[14].n11 XThR.Tn[14] 0.063
R17127 XThR.Tn[14].n83 XThR.Tn[14] 0.0540714
R17128 XThR.Tn[14] XThR.Tn[14].n83 0.038
R17129 XThR.Tn[14].n7 XThR.Tn[14] 0.0143889
R17130 XThR.Tn[14].n81 XThR.Tn[14].n80 0.00771154
R17131 XThR.Tn[14].n76 XThR.Tn[14].n75 0.00771154
R17132 XThR.Tn[14].n71 XThR.Tn[14].n70 0.00771154
R17133 XThR.Tn[14].n66 XThR.Tn[14].n65 0.00771154
R17134 XThR.Tn[14].n61 XThR.Tn[14].n60 0.00771154
R17135 XThR.Tn[14].n56 XThR.Tn[14].n55 0.00771154
R17136 XThR.Tn[14].n51 XThR.Tn[14].n50 0.00771154
R17137 XThR.Tn[14].n46 XThR.Tn[14].n45 0.00771154
R17138 XThR.Tn[14].n41 XThR.Tn[14].n40 0.00771154
R17139 XThR.Tn[14].n36 XThR.Tn[14].n35 0.00771154
R17140 XThR.Tn[14].n31 XThR.Tn[14].n30 0.00771154
R17141 XThR.Tn[14].n26 XThR.Tn[14].n25 0.00771154
R17142 XThR.Tn[14].n21 XThR.Tn[14].n20 0.00771154
R17143 XThR.Tn[14].n16 XThR.Tn[14].n15 0.00771154
R17144 XThR.Tn[14].n11 XThR.Tn[14].n10 0.00771154
R17145 XThR.Tn[12].n87 XThR.Tn[12].n86 256.103
R17146 XThR.Tn[12].n2 XThR.Tn[12].n0 243.68
R17147 XThR.Tn[12].n5 XThR.Tn[12].n3 241.847
R17148 XThR.Tn[12].n2 XThR.Tn[12].n1 205.28
R17149 XThR.Tn[12].n87 XThR.Tn[12].n85 202.095
R17150 XThR.Tn[12].n5 XThR.Tn[12].n4 185
R17151 XThR.Tn[12] XThR.Tn[12].n78 161.363
R17152 XThR.Tn[12] XThR.Tn[12].n73 161.363
R17153 XThR.Tn[12] XThR.Tn[12].n68 161.363
R17154 XThR.Tn[12] XThR.Tn[12].n63 161.363
R17155 XThR.Tn[12] XThR.Tn[12].n58 161.363
R17156 XThR.Tn[12] XThR.Tn[12].n53 161.363
R17157 XThR.Tn[12] XThR.Tn[12].n48 161.363
R17158 XThR.Tn[12] XThR.Tn[12].n43 161.363
R17159 XThR.Tn[12] XThR.Tn[12].n38 161.363
R17160 XThR.Tn[12] XThR.Tn[12].n33 161.363
R17161 XThR.Tn[12] XThR.Tn[12].n28 161.363
R17162 XThR.Tn[12] XThR.Tn[12].n23 161.363
R17163 XThR.Tn[12] XThR.Tn[12].n18 161.363
R17164 XThR.Tn[12] XThR.Tn[12].n13 161.363
R17165 XThR.Tn[12] XThR.Tn[12].n8 161.363
R17166 XThR.Tn[12] XThR.Tn[12].n6 161.363
R17167 XThR.Tn[12].n80 XThR.Tn[12].n79 161.3
R17168 XThR.Tn[12].n75 XThR.Tn[12].n74 161.3
R17169 XThR.Tn[12].n70 XThR.Tn[12].n69 161.3
R17170 XThR.Tn[12].n65 XThR.Tn[12].n64 161.3
R17171 XThR.Tn[12].n60 XThR.Tn[12].n59 161.3
R17172 XThR.Tn[12].n55 XThR.Tn[12].n54 161.3
R17173 XThR.Tn[12].n50 XThR.Tn[12].n49 161.3
R17174 XThR.Tn[12].n45 XThR.Tn[12].n44 161.3
R17175 XThR.Tn[12].n40 XThR.Tn[12].n39 161.3
R17176 XThR.Tn[12].n35 XThR.Tn[12].n34 161.3
R17177 XThR.Tn[12].n30 XThR.Tn[12].n29 161.3
R17178 XThR.Tn[12].n25 XThR.Tn[12].n24 161.3
R17179 XThR.Tn[12].n20 XThR.Tn[12].n19 161.3
R17180 XThR.Tn[12].n15 XThR.Tn[12].n14 161.3
R17181 XThR.Tn[12].n10 XThR.Tn[12].n9 161.3
R17182 XThR.Tn[12].n78 XThR.Tn[12].t18 161.106
R17183 XThR.Tn[12].n73 XThR.Tn[12].t24 161.106
R17184 XThR.Tn[12].n68 XThR.Tn[12].t67 161.106
R17185 XThR.Tn[12].n63 XThR.Tn[12].t52 161.106
R17186 XThR.Tn[12].n58 XThR.Tn[12].t16 161.106
R17187 XThR.Tn[12].n53 XThR.Tn[12].t40 161.106
R17188 XThR.Tn[12].n48 XThR.Tn[12].t22 161.106
R17189 XThR.Tn[12].n43 XThR.Tn[12].t65 161.106
R17190 XThR.Tn[12].n38 XThR.Tn[12].t51 161.106
R17191 XThR.Tn[12].n33 XThR.Tn[12].t56 161.106
R17192 XThR.Tn[12].n28 XThR.Tn[12].t39 161.106
R17193 XThR.Tn[12].n23 XThR.Tn[12].t66 161.106
R17194 XThR.Tn[12].n18 XThR.Tn[12].t38 161.106
R17195 XThR.Tn[12].n13 XThR.Tn[12].t20 161.106
R17196 XThR.Tn[12].n8 XThR.Tn[12].t43 161.106
R17197 XThR.Tn[12].n6 XThR.Tn[12].t28 161.106
R17198 XThR.Tn[12].n79 XThR.Tn[12].t58 159.978
R17199 XThR.Tn[12].n74 XThR.Tn[12].t62 159.978
R17200 XThR.Tn[12].n69 XThR.Tn[12].t47 159.978
R17201 XThR.Tn[12].n64 XThR.Tn[12].t31 159.978
R17202 XThR.Tn[12].n59 XThR.Tn[12].t55 159.978
R17203 XThR.Tn[12].n54 XThR.Tn[12].t19 159.978
R17204 XThR.Tn[12].n49 XThR.Tn[12].t61 159.978
R17205 XThR.Tn[12].n44 XThR.Tn[12].t44 159.978
R17206 XThR.Tn[12].n39 XThR.Tn[12].t29 159.978
R17207 XThR.Tn[12].n34 XThR.Tn[12].t37 159.978
R17208 XThR.Tn[12].n29 XThR.Tn[12].t17 159.978
R17209 XThR.Tn[12].n24 XThR.Tn[12].t46 159.978
R17210 XThR.Tn[12].n19 XThR.Tn[12].t15 159.978
R17211 XThR.Tn[12].n14 XThR.Tn[12].t60 159.978
R17212 XThR.Tn[12].n9 XThR.Tn[12].t21 159.978
R17213 XThR.Tn[12].n78 XThR.Tn[12].t69 145.038
R17214 XThR.Tn[12].n73 XThR.Tn[12].t32 145.038
R17215 XThR.Tn[12].n68 XThR.Tn[12].t73 145.038
R17216 XThR.Tn[12].n63 XThR.Tn[12].t57 145.038
R17217 XThR.Tn[12].n58 XThR.Tn[12].t25 145.038
R17218 XThR.Tn[12].n53 XThR.Tn[12].t68 145.038
R17219 XThR.Tn[12].n48 XThR.Tn[12].t12 145.038
R17220 XThR.Tn[12].n43 XThR.Tn[12].t59 145.038
R17221 XThR.Tn[12].n38 XThR.Tn[12].t54 145.038
R17222 XThR.Tn[12].n33 XThR.Tn[12].t23 145.038
R17223 XThR.Tn[12].n28 XThR.Tn[12].t48 145.038
R17224 XThR.Tn[12].n23 XThR.Tn[12].t70 145.038
R17225 XThR.Tn[12].n18 XThR.Tn[12].t45 145.038
R17226 XThR.Tn[12].n13 XThR.Tn[12].t30 145.038
R17227 XThR.Tn[12].n8 XThR.Tn[12].t53 145.038
R17228 XThR.Tn[12].n6 XThR.Tn[12].t36 145.038
R17229 XThR.Tn[12].n79 XThR.Tn[12].t27 143.911
R17230 XThR.Tn[12].n74 XThR.Tn[12].t50 143.911
R17231 XThR.Tn[12].n69 XThR.Tn[12].t34 143.911
R17232 XThR.Tn[12].n64 XThR.Tn[12].t13 143.911
R17233 XThR.Tn[12].n59 XThR.Tn[12].t42 143.911
R17234 XThR.Tn[12].n54 XThR.Tn[12].t26 143.911
R17235 XThR.Tn[12].n49 XThR.Tn[12].t35 143.911
R17236 XThR.Tn[12].n44 XThR.Tn[12].t14 143.911
R17237 XThR.Tn[12].n39 XThR.Tn[12].t72 143.911
R17238 XThR.Tn[12].n34 XThR.Tn[12].t41 143.911
R17239 XThR.Tn[12].n29 XThR.Tn[12].t64 143.911
R17240 XThR.Tn[12].n24 XThR.Tn[12].t33 143.911
R17241 XThR.Tn[12].n19 XThR.Tn[12].t63 143.911
R17242 XThR.Tn[12].n14 XThR.Tn[12].t49 143.911
R17243 XThR.Tn[12].n9 XThR.Tn[12].t71 143.911
R17244 XThR.Tn[12] XThR.Tn[12].n2 35.7652
R17245 XThR.Tn[12].n85 XThR.Tn[12].t2 26.5955
R17246 XThR.Tn[12].n85 XThR.Tn[12].t0 26.5955
R17247 XThR.Tn[12].n0 XThR.Tn[12].t11 26.5955
R17248 XThR.Tn[12].n0 XThR.Tn[12].t9 26.5955
R17249 XThR.Tn[12].n1 XThR.Tn[12].t8 26.5955
R17250 XThR.Tn[12].n1 XThR.Tn[12].t10 26.5955
R17251 XThR.Tn[12].n86 XThR.Tn[12].t3 26.5955
R17252 XThR.Tn[12].n86 XThR.Tn[12].t1 26.5955
R17253 XThR.Tn[12].n4 XThR.Tn[12].t6 24.9236
R17254 XThR.Tn[12].n4 XThR.Tn[12].t4 24.9236
R17255 XThR.Tn[12].n3 XThR.Tn[12].t7 24.9236
R17256 XThR.Tn[12].n3 XThR.Tn[12].t5 24.9236
R17257 XThR.Tn[12] XThR.Tn[12].n5 18.8943
R17258 XThR.Tn[12].n88 XThR.Tn[12].n87 13.5534
R17259 XThR.Tn[12].n84 XThR.Tn[12] 8.18715
R17260 XThR.Tn[12].n84 XThR.Tn[12] 6.34069
R17261 XThR.Tn[12] XThR.Tn[12].n7 5.34038
R17262 XThR.Tn[12].n12 XThR.Tn[12].n11 4.5005
R17263 XThR.Tn[12].n17 XThR.Tn[12].n16 4.5005
R17264 XThR.Tn[12].n22 XThR.Tn[12].n21 4.5005
R17265 XThR.Tn[12].n27 XThR.Tn[12].n26 4.5005
R17266 XThR.Tn[12].n32 XThR.Tn[12].n31 4.5005
R17267 XThR.Tn[12].n37 XThR.Tn[12].n36 4.5005
R17268 XThR.Tn[12].n42 XThR.Tn[12].n41 4.5005
R17269 XThR.Tn[12].n47 XThR.Tn[12].n46 4.5005
R17270 XThR.Tn[12].n52 XThR.Tn[12].n51 4.5005
R17271 XThR.Tn[12].n57 XThR.Tn[12].n56 4.5005
R17272 XThR.Tn[12].n62 XThR.Tn[12].n61 4.5005
R17273 XThR.Tn[12].n67 XThR.Tn[12].n66 4.5005
R17274 XThR.Tn[12].n72 XThR.Tn[12].n71 4.5005
R17275 XThR.Tn[12].n77 XThR.Tn[12].n76 4.5005
R17276 XThR.Tn[12].n82 XThR.Tn[12].n81 4.5005
R17277 XThR.Tn[12].n83 XThR.Tn[12] 3.70586
R17278 XThR.Tn[12].n12 XThR.Tn[12] 2.52282
R17279 XThR.Tn[12].n17 XThR.Tn[12] 2.52282
R17280 XThR.Tn[12].n22 XThR.Tn[12] 2.52282
R17281 XThR.Tn[12].n27 XThR.Tn[12] 2.52282
R17282 XThR.Tn[12].n32 XThR.Tn[12] 2.52282
R17283 XThR.Tn[12].n37 XThR.Tn[12] 2.52282
R17284 XThR.Tn[12].n42 XThR.Tn[12] 2.52282
R17285 XThR.Tn[12].n47 XThR.Tn[12] 2.52282
R17286 XThR.Tn[12].n52 XThR.Tn[12] 2.52282
R17287 XThR.Tn[12].n57 XThR.Tn[12] 2.52282
R17288 XThR.Tn[12].n62 XThR.Tn[12] 2.52282
R17289 XThR.Tn[12].n67 XThR.Tn[12] 2.52282
R17290 XThR.Tn[12].n72 XThR.Tn[12] 2.52282
R17291 XThR.Tn[12].n77 XThR.Tn[12] 2.52282
R17292 XThR.Tn[12].n82 XThR.Tn[12] 2.52282
R17293 XThR.Tn[12] XThR.Tn[12].n84 1.79489
R17294 XThR.Tn[12] XThR.Tn[12].n88 1.50638
R17295 XThR.Tn[12].n88 XThR.Tn[12] 1.19676
R17296 XThR.Tn[12].n80 XThR.Tn[12] 1.08677
R17297 XThR.Tn[12].n75 XThR.Tn[12] 1.08677
R17298 XThR.Tn[12].n70 XThR.Tn[12] 1.08677
R17299 XThR.Tn[12].n65 XThR.Tn[12] 1.08677
R17300 XThR.Tn[12].n60 XThR.Tn[12] 1.08677
R17301 XThR.Tn[12].n55 XThR.Tn[12] 1.08677
R17302 XThR.Tn[12].n50 XThR.Tn[12] 1.08677
R17303 XThR.Tn[12].n45 XThR.Tn[12] 1.08677
R17304 XThR.Tn[12].n40 XThR.Tn[12] 1.08677
R17305 XThR.Tn[12].n35 XThR.Tn[12] 1.08677
R17306 XThR.Tn[12].n30 XThR.Tn[12] 1.08677
R17307 XThR.Tn[12].n25 XThR.Tn[12] 1.08677
R17308 XThR.Tn[12].n20 XThR.Tn[12] 1.08677
R17309 XThR.Tn[12].n15 XThR.Tn[12] 1.08677
R17310 XThR.Tn[12].n10 XThR.Tn[12] 1.08677
R17311 XThR.Tn[12] XThR.Tn[12].n12 0.839786
R17312 XThR.Tn[12] XThR.Tn[12].n17 0.839786
R17313 XThR.Tn[12] XThR.Tn[12].n22 0.839786
R17314 XThR.Tn[12] XThR.Tn[12].n27 0.839786
R17315 XThR.Tn[12] XThR.Tn[12].n32 0.839786
R17316 XThR.Tn[12] XThR.Tn[12].n37 0.839786
R17317 XThR.Tn[12] XThR.Tn[12].n42 0.839786
R17318 XThR.Tn[12] XThR.Tn[12].n47 0.839786
R17319 XThR.Tn[12] XThR.Tn[12].n52 0.839786
R17320 XThR.Tn[12] XThR.Tn[12].n57 0.839786
R17321 XThR.Tn[12] XThR.Tn[12].n62 0.839786
R17322 XThR.Tn[12] XThR.Tn[12].n67 0.839786
R17323 XThR.Tn[12] XThR.Tn[12].n72 0.839786
R17324 XThR.Tn[12] XThR.Tn[12].n77 0.839786
R17325 XThR.Tn[12] XThR.Tn[12].n82 0.839786
R17326 XThR.Tn[12].n7 XThR.Tn[12] 0.499542
R17327 XThR.Tn[12].n81 XThR.Tn[12] 0.063
R17328 XThR.Tn[12].n76 XThR.Tn[12] 0.063
R17329 XThR.Tn[12].n71 XThR.Tn[12] 0.063
R17330 XThR.Tn[12].n66 XThR.Tn[12] 0.063
R17331 XThR.Tn[12].n61 XThR.Tn[12] 0.063
R17332 XThR.Tn[12].n56 XThR.Tn[12] 0.063
R17333 XThR.Tn[12].n51 XThR.Tn[12] 0.063
R17334 XThR.Tn[12].n46 XThR.Tn[12] 0.063
R17335 XThR.Tn[12].n41 XThR.Tn[12] 0.063
R17336 XThR.Tn[12].n36 XThR.Tn[12] 0.063
R17337 XThR.Tn[12].n31 XThR.Tn[12] 0.063
R17338 XThR.Tn[12].n26 XThR.Tn[12] 0.063
R17339 XThR.Tn[12].n21 XThR.Tn[12] 0.063
R17340 XThR.Tn[12].n16 XThR.Tn[12] 0.063
R17341 XThR.Tn[12].n11 XThR.Tn[12] 0.063
R17342 XThR.Tn[12].n83 XThR.Tn[12] 0.0540714
R17343 XThR.Tn[12] XThR.Tn[12].n83 0.038
R17344 XThR.Tn[12].n7 XThR.Tn[12] 0.0143889
R17345 XThR.Tn[12].n81 XThR.Tn[12].n80 0.00771154
R17346 XThR.Tn[12].n76 XThR.Tn[12].n75 0.00771154
R17347 XThR.Tn[12].n71 XThR.Tn[12].n70 0.00771154
R17348 XThR.Tn[12].n66 XThR.Tn[12].n65 0.00771154
R17349 XThR.Tn[12].n61 XThR.Tn[12].n60 0.00771154
R17350 XThR.Tn[12].n56 XThR.Tn[12].n55 0.00771154
R17351 XThR.Tn[12].n51 XThR.Tn[12].n50 0.00771154
R17352 XThR.Tn[12].n46 XThR.Tn[12].n45 0.00771154
R17353 XThR.Tn[12].n41 XThR.Tn[12].n40 0.00771154
R17354 XThR.Tn[12].n36 XThR.Tn[12].n35 0.00771154
R17355 XThR.Tn[12].n31 XThR.Tn[12].n30 0.00771154
R17356 XThR.Tn[12].n26 XThR.Tn[12].n25 0.00771154
R17357 XThR.Tn[12].n21 XThR.Tn[12].n20 0.00771154
R17358 XThR.Tn[12].n16 XThR.Tn[12].n15 0.00771154
R17359 XThR.Tn[12].n11 XThR.Tn[12].n10 0.00771154
R17360 XThC.XTBN.Y.n182 XThC.XTBN.Y.t9 212.081
R17361 XThC.XTBN.Y.n181 XThC.XTBN.Y.t75 212.081
R17362 XThC.XTBN.Y.n175 XThC.XTBN.Y.t33 212.081
R17363 XThC.XTBN.Y.n176 XThC.XTBN.Y.t27 212.081
R17364 XThC.XTBN.Y.n87 XThC.XTBN.Y.t25 212.081
R17365 XThC.XTBN.Y.n78 XThC.XTBN.Y.t100 212.081
R17366 XThC.XTBN.Y.n82 XThC.XTBN.Y.t93 212.081
R17367 XThC.XTBN.Y.n80 XThC.XTBN.Y.t90 212.081
R17368 XThC.XTBN.Y.n61 XThC.XTBN.Y.t47 212.081
R17369 XThC.XTBN.Y.n52 XThC.XTBN.Y.t17 212.081
R17370 XThC.XTBN.Y.n56 XThC.XTBN.Y.t116 212.081
R17371 XThC.XTBN.Y.n54 XThC.XTBN.Y.t111 212.081
R17372 XThC.XTBN.Y.n35 XThC.XTBN.Y.t106 212.081
R17373 XThC.XTBN.Y.n26 XThC.XTBN.Y.t70 212.081
R17374 XThC.XTBN.Y.n30 XThC.XTBN.Y.t56 212.081
R17375 XThC.XTBN.Y.n28 XThC.XTBN.Y.t48 212.081
R17376 XThC.XTBN.Y.n10 XThC.XTBN.Y.t50 212.081
R17377 XThC.XTBN.Y.n1 XThC.XTBN.Y.t18 212.081
R17378 XThC.XTBN.Y.n5 XThC.XTBN.Y.t120 212.081
R17379 XThC.XTBN.Y.n3 XThC.XTBN.Y.t114 212.081
R17380 XThC.XTBN.Y.n74 XThC.XTBN.Y.t101 212.081
R17381 XThC.XTBN.Y.n65 XThC.XTBN.Y.t63 212.081
R17382 XThC.XTBN.Y.n69 XThC.XTBN.Y.t52 212.081
R17383 XThC.XTBN.Y.n67 XThC.XTBN.Y.t44 212.081
R17384 XThC.XTBN.Y.n48 XThC.XTBN.Y.t39 212.081
R17385 XThC.XTBN.Y.n39 XThC.XTBN.Y.t122 212.081
R17386 XThC.XTBN.Y.n43 XThC.XTBN.Y.t109 212.081
R17387 XThC.XTBN.Y.n41 XThC.XTBN.Y.t102 212.081
R17388 XThC.XTBN.Y.n22 XThC.XTBN.Y.t79 212.081
R17389 XThC.XTBN.Y.n13 XThC.XTBN.Y.t36 212.081
R17390 XThC.XTBN.Y.n17 XThC.XTBN.Y.t26 212.081
R17391 XThC.XTBN.Y.n15 XThC.XTBN.Y.t21 212.081
R17392 XThC.XTBN.Y.n99 XThC.XTBN.Y.t54 212.081
R17393 XThC.XTBN.Y.n98 XThC.XTBN.Y.t46 212.081
R17394 XThC.XTBN.Y.n93 XThC.XTBN.Y.t12 212.081
R17395 XThC.XTBN.Y.n92 XThC.XTBN.Y.t6 212.081
R17396 XThC.XTBN.Y.n122 XThC.XTBN.Y.t34 212.081
R17397 XThC.XTBN.Y.n121 XThC.XTBN.Y.t30 212.081
R17398 XThC.XTBN.Y.n116 XThC.XTBN.Y.t103 212.081
R17399 XThC.XTBN.Y.n115 XThC.XTBN.Y.t98 212.081
R17400 XThC.XTBN.Y.n146 XThC.XTBN.Y.t91 212.081
R17401 XThC.XTBN.Y.n145 XThC.XTBN.Y.t88 212.081
R17402 XThC.XTBN.Y.n140 XThC.XTBN.Y.t40 212.081
R17403 XThC.XTBN.Y.n139 XThC.XTBN.Y.t37 212.081
R17404 XThC.XTBN.Y.n170 XThC.XTBN.Y.t28 212.081
R17405 XThC.XTBN.Y.n169 XThC.XTBN.Y.t23 212.081
R17406 XThC.XTBN.Y.n164 XThC.XTBN.Y.t97 212.081
R17407 XThC.XTBN.Y.n163 XThC.XTBN.Y.t95 212.081
R17408 XThC.XTBN.Y.n110 XThC.XTBN.Y.t42 212.081
R17409 XThC.XTBN.Y.n109 XThC.XTBN.Y.t38 212.081
R17410 XThC.XTBN.Y.n104 XThC.XTBN.Y.t119 212.081
R17411 XThC.XTBN.Y.n103 XThC.XTBN.Y.t113 212.081
R17412 XThC.XTBN.Y.n134 XThC.XTBN.Y.t99 212.081
R17413 XThC.XTBN.Y.n133 XThC.XTBN.Y.t96 212.081
R17414 XThC.XTBN.Y.n128 XThC.XTBN.Y.t58 212.081
R17415 XThC.XTBN.Y.n127 XThC.XTBN.Y.t51 212.081
R17416 XThC.XTBN.Y.n158 XThC.XTBN.Y.t13 212.081
R17417 XThC.XTBN.Y.n157 XThC.XTBN.Y.t7 212.081
R17418 XThC.XTBN.Y.n152 XThC.XTBN.Y.t86 212.081
R17419 XThC.XTBN.Y.n151 XThC.XTBN.Y.t81 212.081
R17420 XThC.XTBN.Y.n192 XThC.XTBN.Y.n191 208.964
R17421 XThC.XTBN.Y.n176 XThC.XTBN.Y.n0 188.516
R17422 XThC.XTBN.Y.n88 XThC.XTBN.Y.n87 180.482
R17423 XThC.XTBN.Y.n62 XThC.XTBN.Y.n61 180.482
R17424 XThC.XTBN.Y.n36 XThC.XTBN.Y.n35 180.482
R17425 XThC.XTBN.Y.n11 XThC.XTBN.Y.n10 180.482
R17426 XThC.XTBN.Y.n75 XThC.XTBN.Y.n74 180.482
R17427 XThC.XTBN.Y.n49 XThC.XTBN.Y.n48 180.482
R17428 XThC.XTBN.Y.n23 XThC.XTBN.Y.n22 180.482
R17429 XThC.XTBN.Y.n95 XThC.XTBN.Y.n94 173.761
R17430 XThC.XTBN.Y.n118 XThC.XTBN.Y.n117 173.761
R17431 XThC.XTBN.Y.n142 XThC.XTBN.Y.n141 173.761
R17432 XThC.XTBN.Y.n166 XThC.XTBN.Y.n165 173.761
R17433 XThC.XTBN.Y.n106 XThC.XTBN.Y.n105 173.761
R17434 XThC.XTBN.Y.n130 XThC.XTBN.Y.n129 173.761
R17435 XThC.XTBN.Y.n154 XThC.XTBN.Y.n153 173.761
R17436 XThC.XTBN.Y.n81 XThC.XTBN.Y.n79 152
R17437 XThC.XTBN.Y.n84 XThC.XTBN.Y.n83 152
R17438 XThC.XTBN.Y.n86 XThC.XTBN.Y.n85 152
R17439 XThC.XTBN.Y.n55 XThC.XTBN.Y.n53 152
R17440 XThC.XTBN.Y.n58 XThC.XTBN.Y.n57 152
R17441 XThC.XTBN.Y.n60 XThC.XTBN.Y.n59 152
R17442 XThC.XTBN.Y.n29 XThC.XTBN.Y.n27 152
R17443 XThC.XTBN.Y.n32 XThC.XTBN.Y.n31 152
R17444 XThC.XTBN.Y.n34 XThC.XTBN.Y.n33 152
R17445 XThC.XTBN.Y.n4 XThC.XTBN.Y.n2 152
R17446 XThC.XTBN.Y.n7 XThC.XTBN.Y.n6 152
R17447 XThC.XTBN.Y.n9 XThC.XTBN.Y.n8 152
R17448 XThC.XTBN.Y.n68 XThC.XTBN.Y.n66 152
R17449 XThC.XTBN.Y.n71 XThC.XTBN.Y.n70 152
R17450 XThC.XTBN.Y.n73 XThC.XTBN.Y.n72 152
R17451 XThC.XTBN.Y.n42 XThC.XTBN.Y.n40 152
R17452 XThC.XTBN.Y.n45 XThC.XTBN.Y.n44 152
R17453 XThC.XTBN.Y.n47 XThC.XTBN.Y.n46 152
R17454 XThC.XTBN.Y.n16 XThC.XTBN.Y.n14 152
R17455 XThC.XTBN.Y.n19 XThC.XTBN.Y.n18 152
R17456 XThC.XTBN.Y.n21 XThC.XTBN.Y.n20 152
R17457 XThC.XTBN.Y.n95 XThC.XTBN.Y.n91 152
R17458 XThC.XTBN.Y.n97 XThC.XTBN.Y.n96 152
R17459 XThC.XTBN.Y.n101 XThC.XTBN.Y.n100 152
R17460 XThC.XTBN.Y.n118 XThC.XTBN.Y.n114 152
R17461 XThC.XTBN.Y.n120 XThC.XTBN.Y.n119 152
R17462 XThC.XTBN.Y.n124 XThC.XTBN.Y.n123 152
R17463 XThC.XTBN.Y.n142 XThC.XTBN.Y.n138 152
R17464 XThC.XTBN.Y.n144 XThC.XTBN.Y.n143 152
R17465 XThC.XTBN.Y.n148 XThC.XTBN.Y.n147 152
R17466 XThC.XTBN.Y.n166 XThC.XTBN.Y.n162 152
R17467 XThC.XTBN.Y.n168 XThC.XTBN.Y.n167 152
R17468 XThC.XTBN.Y.n172 XThC.XTBN.Y.n171 152
R17469 XThC.XTBN.Y.n106 XThC.XTBN.Y.n102 152
R17470 XThC.XTBN.Y.n108 XThC.XTBN.Y.n107 152
R17471 XThC.XTBN.Y.n112 XThC.XTBN.Y.n111 152
R17472 XThC.XTBN.Y.n130 XThC.XTBN.Y.n126 152
R17473 XThC.XTBN.Y.n132 XThC.XTBN.Y.n131 152
R17474 XThC.XTBN.Y.n136 XThC.XTBN.Y.n135 152
R17475 XThC.XTBN.Y.n154 XThC.XTBN.Y.n150 152
R17476 XThC.XTBN.Y.n156 XThC.XTBN.Y.n155 152
R17477 XThC.XTBN.Y.n160 XThC.XTBN.Y.n159 152
R17478 XThC.XTBN.Y.n178 XThC.XTBN.Y.n177 152
R17479 XThC.XTBN.Y.n180 XThC.XTBN.Y.n179 152
R17480 XThC.XTBN.Y.n184 XThC.XTBN.Y.n183 152
R17481 XThC.XTBN.Y.n182 XThC.XTBN.Y.t14 139.78
R17482 XThC.XTBN.Y.n181 XThC.XTBN.Y.t105 139.78
R17483 XThC.XTBN.Y.n175 XThC.XTBN.Y.t69 139.78
R17484 XThC.XTBN.Y.n176 XThC.XTBN.Y.t61 139.78
R17485 XThC.XTBN.Y.n87 XThC.XTBN.Y.t123 139.78
R17486 XThC.XTBN.Y.n78 XThC.XTBN.Y.t85 139.78
R17487 XThC.XTBN.Y.n82 XThC.XTBN.Y.t74 139.78
R17488 XThC.XTBN.Y.n80 XThC.XTBN.Y.t65 139.78
R17489 XThC.XTBN.Y.n61 XThC.XTBN.Y.t31 139.78
R17490 XThC.XTBN.Y.n52 XThC.XTBN.Y.t104 139.78
R17491 XThC.XTBN.Y.n56 XThC.XTBN.Y.t94 139.78
R17492 XThC.XTBN.Y.n54 XThC.XTBN.Y.t92 139.78
R17493 XThC.XTBN.Y.n35 XThC.XTBN.Y.t89 139.78
R17494 XThC.XTBN.Y.n26 XThC.XTBN.Y.t41 139.78
R17495 XThC.XTBN.Y.n30 XThC.XTBN.Y.t35 139.78
R17496 XThC.XTBN.Y.n28 XThC.XTBN.Y.t32 139.78
R17497 XThC.XTBN.Y.n10 XThC.XTBN.Y.t118 139.78
R17498 XThC.XTBN.Y.n1 XThC.XTBN.Y.t83 139.78
R17499 XThC.XTBN.Y.n5 XThC.XTBN.Y.t71 139.78
R17500 XThC.XTBN.Y.n3 XThC.XTBN.Y.t62 139.78
R17501 XThC.XTBN.Y.n74 XThC.XTBN.Y.t107 139.78
R17502 XThC.XTBN.Y.n65 XThC.XTBN.Y.t72 139.78
R17503 XThC.XTBN.Y.n69 XThC.XTBN.Y.t57 139.78
R17504 XThC.XTBN.Y.n67 XThC.XTBN.Y.t49 139.78
R17505 XThC.XTBN.Y.n48 XThC.XTBN.Y.t43 139.78
R17506 XThC.XTBN.Y.n39 XThC.XTBN.Y.t10 139.78
R17507 XThC.XTBN.Y.n43 XThC.XTBN.Y.t112 139.78
R17508 XThC.XTBN.Y.n41 XThC.XTBN.Y.t108 139.78
R17509 XThC.XTBN.Y.n22 XThC.XTBN.Y.t121 139.78
R17510 XThC.XTBN.Y.n13 XThC.XTBN.Y.t84 139.78
R17511 XThC.XTBN.Y.n17 XThC.XTBN.Y.t73 139.78
R17512 XThC.XTBN.Y.n15 XThC.XTBN.Y.t64 139.78
R17513 XThC.XTBN.Y.n99 XThC.XTBN.Y.t76 139.78
R17514 XThC.XTBN.Y.n98 XThC.XTBN.Y.t67 139.78
R17515 XThC.XTBN.Y.n93 XThC.XTBN.Y.t29 139.78
R17516 XThC.XTBN.Y.n92 XThC.XTBN.Y.t24 139.78
R17517 XThC.XTBN.Y.n122 XThC.XTBN.Y.t15 139.78
R17518 XThC.XTBN.Y.n121 XThC.XTBN.Y.t8 139.78
R17519 XThC.XTBN.Y.n116 XThC.XTBN.Y.t87 139.78
R17520 XThC.XTBN.Y.n115 XThC.XTBN.Y.t82 139.78
R17521 XThC.XTBN.Y.n146 XThC.XTBN.Y.t66 139.78
R17522 XThC.XTBN.Y.n145 XThC.XTBN.Y.t60 139.78
R17523 XThC.XTBN.Y.n140 XThC.XTBN.Y.t22 139.78
R17524 XThC.XTBN.Y.n139 XThC.XTBN.Y.t20 139.78
R17525 XThC.XTBN.Y.n170 XThC.XTBN.Y.t4 139.78
R17526 XThC.XTBN.Y.n169 XThC.XTBN.Y.t117 139.78
R17527 XThC.XTBN.Y.n164 XThC.XTBN.Y.t80 139.78
R17528 XThC.XTBN.Y.n163 XThC.XTBN.Y.t78 139.78
R17529 XThC.XTBN.Y.n110 XThC.XTBN.Y.t59 139.78
R17530 XThC.XTBN.Y.n109 XThC.XTBN.Y.t55 139.78
R17531 XThC.XTBN.Y.n104 XThC.XTBN.Y.t19 139.78
R17532 XThC.XTBN.Y.n103 XThC.XTBN.Y.t16 139.78
R17533 XThC.XTBN.Y.n134 XThC.XTBN.Y.t115 139.78
R17534 XThC.XTBN.Y.n133 XThC.XTBN.Y.t110 139.78
R17535 XThC.XTBN.Y.n128 XThC.XTBN.Y.t77 139.78
R17536 XThC.XTBN.Y.n127 XThC.XTBN.Y.t68 139.78
R17537 XThC.XTBN.Y.n158 XThC.XTBN.Y.t53 139.78
R17538 XThC.XTBN.Y.n157 XThC.XTBN.Y.t45 139.78
R17539 XThC.XTBN.Y.n152 XThC.XTBN.Y.t11 139.78
R17540 XThC.XTBN.Y.n151 XThC.XTBN.Y.t5 139.78
R17541 XThC.XTBN.Y XThC.XTBN.Y.n188 96.8352
R17542 XThC.XTBN.Y.n187 XThC.XTBN.Y.n0 64.6909
R17543 XThC.XTBN.Y.n97 XThC.XTBN.Y.n91 49.6611
R17544 XThC.XTBN.Y.n120 XThC.XTBN.Y.n114 49.6611
R17545 XThC.XTBN.Y.n144 XThC.XTBN.Y.n138 49.6611
R17546 XThC.XTBN.Y.n168 XThC.XTBN.Y.n162 49.6611
R17547 XThC.XTBN.Y.n108 XThC.XTBN.Y.n102 49.6611
R17548 XThC.XTBN.Y.n132 XThC.XTBN.Y.n126 49.6611
R17549 XThC.XTBN.Y.n156 XThC.XTBN.Y.n150 49.6611
R17550 XThC.XTBN.Y.n100 XThC.XTBN.Y.n98 44.549
R17551 XThC.XTBN.Y.n123 XThC.XTBN.Y.n121 44.549
R17552 XThC.XTBN.Y.n147 XThC.XTBN.Y.n145 44.549
R17553 XThC.XTBN.Y.n171 XThC.XTBN.Y.n169 44.549
R17554 XThC.XTBN.Y.n111 XThC.XTBN.Y.n109 44.549
R17555 XThC.XTBN.Y.n135 XThC.XTBN.Y.n133 44.549
R17556 XThC.XTBN.Y.n159 XThC.XTBN.Y.n157 44.549
R17557 XThC.XTBN.Y.n94 XThC.XTBN.Y.n93 43.0884
R17558 XThC.XTBN.Y.n117 XThC.XTBN.Y.n116 43.0884
R17559 XThC.XTBN.Y.n141 XThC.XTBN.Y.n140 43.0884
R17560 XThC.XTBN.Y.n165 XThC.XTBN.Y.n164 43.0884
R17561 XThC.XTBN.Y.n105 XThC.XTBN.Y.n104 43.0884
R17562 XThC.XTBN.Y.n129 XThC.XTBN.Y.n128 43.0884
R17563 XThC.XTBN.Y.n153 XThC.XTBN.Y.n152 43.0884
R17564 XThC.XTBN.Y.n177 XThC.XTBN.Y.n176 30.6732
R17565 XThC.XTBN.Y.n177 XThC.XTBN.Y.n175 30.6732
R17566 XThC.XTBN.Y.n180 XThC.XTBN.Y.n175 30.6732
R17567 XThC.XTBN.Y.n181 XThC.XTBN.Y.n180 30.6732
R17568 XThC.XTBN.Y.n183 XThC.XTBN.Y.n181 30.6732
R17569 XThC.XTBN.Y.n183 XThC.XTBN.Y.n182 30.6732
R17570 XThC.XTBN.Y.n81 XThC.XTBN.Y.n80 30.6732
R17571 XThC.XTBN.Y.n82 XThC.XTBN.Y.n81 30.6732
R17572 XThC.XTBN.Y.n83 XThC.XTBN.Y.n82 30.6732
R17573 XThC.XTBN.Y.n83 XThC.XTBN.Y.n78 30.6732
R17574 XThC.XTBN.Y.n86 XThC.XTBN.Y.n78 30.6732
R17575 XThC.XTBN.Y.n87 XThC.XTBN.Y.n86 30.6732
R17576 XThC.XTBN.Y.n55 XThC.XTBN.Y.n54 30.6732
R17577 XThC.XTBN.Y.n56 XThC.XTBN.Y.n55 30.6732
R17578 XThC.XTBN.Y.n57 XThC.XTBN.Y.n56 30.6732
R17579 XThC.XTBN.Y.n57 XThC.XTBN.Y.n52 30.6732
R17580 XThC.XTBN.Y.n60 XThC.XTBN.Y.n52 30.6732
R17581 XThC.XTBN.Y.n61 XThC.XTBN.Y.n60 30.6732
R17582 XThC.XTBN.Y.n29 XThC.XTBN.Y.n28 30.6732
R17583 XThC.XTBN.Y.n30 XThC.XTBN.Y.n29 30.6732
R17584 XThC.XTBN.Y.n31 XThC.XTBN.Y.n30 30.6732
R17585 XThC.XTBN.Y.n31 XThC.XTBN.Y.n26 30.6732
R17586 XThC.XTBN.Y.n34 XThC.XTBN.Y.n26 30.6732
R17587 XThC.XTBN.Y.n35 XThC.XTBN.Y.n34 30.6732
R17588 XThC.XTBN.Y.n4 XThC.XTBN.Y.n3 30.6732
R17589 XThC.XTBN.Y.n5 XThC.XTBN.Y.n4 30.6732
R17590 XThC.XTBN.Y.n6 XThC.XTBN.Y.n5 30.6732
R17591 XThC.XTBN.Y.n6 XThC.XTBN.Y.n1 30.6732
R17592 XThC.XTBN.Y.n9 XThC.XTBN.Y.n1 30.6732
R17593 XThC.XTBN.Y.n10 XThC.XTBN.Y.n9 30.6732
R17594 XThC.XTBN.Y.n68 XThC.XTBN.Y.n67 30.6732
R17595 XThC.XTBN.Y.n69 XThC.XTBN.Y.n68 30.6732
R17596 XThC.XTBN.Y.n70 XThC.XTBN.Y.n69 30.6732
R17597 XThC.XTBN.Y.n70 XThC.XTBN.Y.n65 30.6732
R17598 XThC.XTBN.Y.n73 XThC.XTBN.Y.n65 30.6732
R17599 XThC.XTBN.Y.n74 XThC.XTBN.Y.n73 30.6732
R17600 XThC.XTBN.Y.n42 XThC.XTBN.Y.n41 30.6732
R17601 XThC.XTBN.Y.n43 XThC.XTBN.Y.n42 30.6732
R17602 XThC.XTBN.Y.n44 XThC.XTBN.Y.n43 30.6732
R17603 XThC.XTBN.Y.n44 XThC.XTBN.Y.n39 30.6732
R17604 XThC.XTBN.Y.n47 XThC.XTBN.Y.n39 30.6732
R17605 XThC.XTBN.Y.n48 XThC.XTBN.Y.n47 30.6732
R17606 XThC.XTBN.Y.n16 XThC.XTBN.Y.n15 30.6732
R17607 XThC.XTBN.Y.n17 XThC.XTBN.Y.n16 30.6732
R17608 XThC.XTBN.Y.n18 XThC.XTBN.Y.n17 30.6732
R17609 XThC.XTBN.Y.n18 XThC.XTBN.Y.n13 30.6732
R17610 XThC.XTBN.Y.n21 XThC.XTBN.Y.n13 30.6732
R17611 XThC.XTBN.Y.n22 XThC.XTBN.Y.n21 30.6732
R17612 XThC.XTBN.Y.n191 XThC.XTBN.Y.t0 26.5955
R17613 XThC.XTBN.Y.n191 XThC.XTBN.Y.t1 26.5955
R17614 XThC.XTBN.Y.n188 XThC.XTBN.Y.t3 24.9236
R17615 XThC.XTBN.Y.n188 XThC.XTBN.Y.t2 24.9236
R17616 XThC.XTBN.Y.n96 XThC.XTBN.Y.n95 21.7605
R17617 XThC.XTBN.Y.n119 XThC.XTBN.Y.n118 21.7605
R17618 XThC.XTBN.Y.n143 XThC.XTBN.Y.n142 21.7605
R17619 XThC.XTBN.Y.n167 XThC.XTBN.Y.n166 21.7605
R17620 XThC.XTBN.Y.n107 XThC.XTBN.Y.n106 21.7605
R17621 XThC.XTBN.Y.n131 XThC.XTBN.Y.n130 21.7605
R17622 XThC.XTBN.Y.n155 XThC.XTBN.Y.n154 21.7605
R17623 XThC.XTBN.Y.n84 XThC.XTBN.Y.n79 21.5045
R17624 XThC.XTBN.Y.n58 XThC.XTBN.Y.n53 21.5045
R17625 XThC.XTBN.Y.n32 XThC.XTBN.Y.n27 21.5045
R17626 XThC.XTBN.Y.n7 XThC.XTBN.Y.n2 21.5045
R17627 XThC.XTBN.Y.n71 XThC.XTBN.Y.n66 21.5045
R17628 XThC.XTBN.Y.n45 XThC.XTBN.Y.n40 21.5045
R17629 XThC.XTBN.Y.n19 XThC.XTBN.Y.n14 21.5045
R17630 XThC.XTBN.Y.n178 XThC.XTBN.Y 21.2485
R17631 XThC.XTBN.Y.n85 XThC.XTBN.Y 19.9685
R17632 XThC.XTBN.Y.n59 XThC.XTBN.Y 19.9685
R17633 XThC.XTBN.Y.n33 XThC.XTBN.Y 19.9685
R17634 XThC.XTBN.Y.n8 XThC.XTBN.Y 19.9685
R17635 XThC.XTBN.Y.n72 XThC.XTBN.Y 19.9685
R17636 XThC.XTBN.Y.n46 XThC.XTBN.Y 19.9685
R17637 XThC.XTBN.Y.n20 XThC.XTBN.Y 19.9685
R17638 XThC.XTBN.Y.n179 XThC.XTBN.Y 19.2005
R17639 XThC.XTBN.Y.n94 XThC.XTBN.Y.n92 18.2581
R17640 XThC.XTBN.Y.n117 XThC.XTBN.Y.n115 18.2581
R17641 XThC.XTBN.Y.n141 XThC.XTBN.Y.n139 18.2581
R17642 XThC.XTBN.Y.n165 XThC.XTBN.Y.n163 18.2581
R17643 XThC.XTBN.Y.n105 XThC.XTBN.Y.n103 18.2581
R17644 XThC.XTBN.Y.n129 XThC.XTBN.Y.n127 18.2581
R17645 XThC.XTBN.Y.n153 XThC.XTBN.Y.n151 18.2581
R17646 XThC.XTBN.Y.n113 XThC.XTBN.Y.n101 17.1655
R17647 XThC.XTBN.Y.n88 XThC.XTBN.Y 17.1525
R17648 XThC.XTBN.Y.n62 XThC.XTBN.Y 17.1525
R17649 XThC.XTBN.Y.n36 XThC.XTBN.Y 17.1525
R17650 XThC.XTBN.Y.n11 XThC.XTBN.Y 17.1525
R17651 XThC.XTBN.Y.n75 XThC.XTBN.Y 17.1525
R17652 XThC.XTBN.Y.n49 XThC.XTBN.Y 17.1525
R17653 XThC.XTBN.Y.n23 XThC.XTBN.Y 17.1525
R17654 XThC.XTBN.Y.n100 XThC.XTBN.Y.n99 16.7975
R17655 XThC.XTBN.Y.n123 XThC.XTBN.Y.n122 16.7975
R17656 XThC.XTBN.Y.n147 XThC.XTBN.Y.n146 16.7975
R17657 XThC.XTBN.Y.n171 XThC.XTBN.Y.n170 16.7975
R17658 XThC.XTBN.Y.n111 XThC.XTBN.Y.n110 16.7975
R17659 XThC.XTBN.Y.n135 XThC.XTBN.Y.n134 16.7975
R17660 XThC.XTBN.Y.n159 XThC.XTBN.Y.n158 16.7975
R17661 XThC.XTBN.Y.n125 XThC.XTBN.Y.n124 16.0405
R17662 XThC.XTBN.Y.n149 XThC.XTBN.Y.n148 16.0405
R17663 XThC.XTBN.Y.n173 XThC.XTBN.Y.n172 16.0405
R17664 XThC.XTBN.Y.n113 XThC.XTBN.Y.n112 16.0405
R17665 XThC.XTBN.Y.n137 XThC.XTBN.Y.n136 16.0405
R17666 XThC.XTBN.Y.n161 XThC.XTBN.Y.n160 16.0405
R17667 XThC.XTBN.Y.n25 XThC.XTBN.Y.n12 15.262
R17668 XThC.XTBN.Y.n101 XThC.XTBN.Y 15.0405
R17669 XThC.XTBN.Y.n124 XThC.XTBN.Y 15.0405
R17670 XThC.XTBN.Y.n148 XThC.XTBN.Y 15.0405
R17671 XThC.XTBN.Y.n172 XThC.XTBN.Y 15.0405
R17672 XThC.XTBN.Y.n112 XThC.XTBN.Y 15.0405
R17673 XThC.XTBN.Y.n136 XThC.XTBN.Y 15.0405
R17674 XThC.XTBN.Y.n160 XThC.XTBN.Y 15.0405
R17675 XThC.XTBN.Y.n90 XThC.XTBN.Y.n89 13.8005
R17676 XThC.XTBN.Y.n64 XThC.XTBN.Y.n63 13.8005
R17677 XThC.XTBN.Y.n38 XThC.XTBN.Y.n37 13.8005
R17678 XThC.XTBN.Y.n77 XThC.XTBN.Y.n76 13.8005
R17679 XThC.XTBN.Y.n51 XThC.XTBN.Y.n50 13.8005
R17680 XThC.XTBN.Y.n25 XThC.XTBN.Y.n24 13.8005
R17681 XThC.XTBN.Y XThC.XTBN.Y.n190 12.5445
R17682 XThC.XTBN.Y XThC.XTBN.Y.n189 11.2645
R17683 XThC.XTBN.Y.n185 XThC.XTBN.Y.n184 9.2165
R17684 XThC.XTBN.Y.n185 XThC.XTBN.Y 7.9365
R17685 XThC.XTBN.Y.n96 XThC.XTBN.Y 6.7205
R17686 XThC.XTBN.Y.n119 XThC.XTBN.Y 6.7205
R17687 XThC.XTBN.Y.n143 XThC.XTBN.Y 6.7205
R17688 XThC.XTBN.Y.n167 XThC.XTBN.Y 6.7205
R17689 XThC.XTBN.Y.n107 XThC.XTBN.Y 6.7205
R17690 XThC.XTBN.Y.n131 XThC.XTBN.Y 6.7205
R17691 XThC.XTBN.Y.n155 XThC.XTBN.Y 6.7205
R17692 XThC.XTBN.Y.n93 XThC.XTBN.Y.n91 6.57323
R17693 XThC.XTBN.Y.n116 XThC.XTBN.Y.n114 6.57323
R17694 XThC.XTBN.Y.n140 XThC.XTBN.Y.n138 6.57323
R17695 XThC.XTBN.Y.n164 XThC.XTBN.Y.n162 6.57323
R17696 XThC.XTBN.Y.n104 XThC.XTBN.Y.n102 6.57323
R17697 XThC.XTBN.Y.n128 XThC.XTBN.Y.n126 6.57323
R17698 XThC.XTBN.Y.n152 XThC.XTBN.Y.n150 6.57323
R17699 XThC.XTBN.Y.n184 XThC.XTBN.Y 6.4005
R17700 XThC.XTBN.Y.n189 XThC.XTBN.Y 6.1445
R17701 XThC.XTBN.Y.n187 XThC.XTBN.Y.n186 5.74665
R17702 XThC.XTBN.Y.n186 XThC.XTBN.Y.n174 5.68319
R17703 XThC.XTBN.Y.n98 XThC.XTBN.Y.n97 5.11262
R17704 XThC.XTBN.Y.n121 XThC.XTBN.Y.n120 5.11262
R17705 XThC.XTBN.Y.n145 XThC.XTBN.Y.n144 5.11262
R17706 XThC.XTBN.Y.n169 XThC.XTBN.Y.n168 5.11262
R17707 XThC.XTBN.Y.n109 XThC.XTBN.Y.n108 5.11262
R17708 XThC.XTBN.Y.n133 XThC.XTBN.Y.n132 5.11262
R17709 XThC.XTBN.Y.n157 XThC.XTBN.Y.n156 5.11262
R17710 XThC.XTBN.Y.n190 XThC.XTBN.Y.n187 5.06717
R17711 XThC.XTBN.Y.n190 XThC.XTBN.Y 4.8645
R17712 XThC.XTBN.Y.n189 XThC.XTBN.Y 4.65505
R17713 XThC.XTBN.Y.n186 XThC.XTBN.Y.n185 4.6505
R17714 XThC.XTBN.Y.n89 XThC.XTBN.Y 4.6085
R17715 XThC.XTBN.Y.n63 XThC.XTBN.Y 4.6085
R17716 XThC.XTBN.Y.n37 XThC.XTBN.Y 4.6085
R17717 XThC.XTBN.Y.n12 XThC.XTBN.Y 4.6085
R17718 XThC.XTBN.Y.n76 XThC.XTBN.Y 4.6085
R17719 XThC.XTBN.Y.n50 XThC.XTBN.Y 4.6085
R17720 XThC.XTBN.Y.n24 XThC.XTBN.Y 4.6085
R17721 XThC.XTBN.Y.n179 XThC.XTBN.Y 4.3525
R17722 XThC.XTBN.Y.n85 XThC.XTBN.Y 3.5845
R17723 XThC.XTBN.Y.n59 XThC.XTBN.Y 3.5845
R17724 XThC.XTBN.Y.n33 XThC.XTBN.Y 3.5845
R17725 XThC.XTBN.Y.n8 XThC.XTBN.Y 3.5845
R17726 XThC.XTBN.Y.n72 XThC.XTBN.Y 3.5845
R17727 XThC.XTBN.Y.n46 XThC.XTBN.Y 3.5845
R17728 XThC.XTBN.Y.n20 XThC.XTBN.Y 3.5845
R17729 XThC.XTBN.Y XThC.XTBN.Y.n0 2.3045
R17730 XThC.XTBN.Y XThC.XTBN.Y.n178 2.3045
R17731 XThC.XTBN.Y.n192 XThC.XTBN.Y 2.0485
R17732 XThC.XTBN.Y.n89 XThC.XTBN.Y.n88 1.7925
R17733 XThC.XTBN.Y.n63 XThC.XTBN.Y.n62 1.7925
R17734 XThC.XTBN.Y.n37 XThC.XTBN.Y.n36 1.7925
R17735 XThC.XTBN.Y.n12 XThC.XTBN.Y.n11 1.7925
R17736 XThC.XTBN.Y.n76 XThC.XTBN.Y.n75 1.7925
R17737 XThC.XTBN.Y.n50 XThC.XTBN.Y.n49 1.7925
R17738 XThC.XTBN.Y.n24 XThC.XTBN.Y.n23 1.7925
R17739 XThC.XTBN.Y.n174 XThC.XTBN.Y.n173 1.59665
R17740 XThC.XTBN.Y XThC.XTBN.Y.n192 1.55202
R17741 XThC.XTBN.Y XThC.XTBN.Y.n84 1.5365
R17742 XThC.XTBN.Y XThC.XTBN.Y.n58 1.5365
R17743 XThC.XTBN.Y XThC.XTBN.Y.n32 1.5365
R17744 XThC.XTBN.Y XThC.XTBN.Y.n7 1.5365
R17745 XThC.XTBN.Y XThC.XTBN.Y.n71 1.5365
R17746 XThC.XTBN.Y XThC.XTBN.Y.n45 1.5365
R17747 XThC.XTBN.Y XThC.XTBN.Y.n19 1.5365
R17748 XThC.XTBN.Y.n149 XThC.XTBN.Y.n137 1.49088
R17749 XThC.XTBN.Y.n125 XThC.XTBN.Y.n113 1.49088
R17750 XThC.XTBN.Y.n173 XThC.XTBN.Y.n161 1.48608
R17751 XThC.XTBN.Y.n51 XThC.XTBN.Y.n38 1.46204
R17752 XThC.XTBN.Y.n77 XThC.XTBN.Y.n64 1.46204
R17753 XThC.XTBN.Y.n38 XThC.XTBN.Y.n25 1.15435
R17754 XThC.XTBN.Y.n64 XThC.XTBN.Y.n51 1.15435
R17755 XThC.XTBN.Y.n90 XThC.XTBN.Y.n77 1.15435
R17756 XThC.XTBN.Y.n174 XThC.XTBN.Y.n90 1.14473
R17757 XThC.XTBN.Y.n161 XThC.XTBN.Y.n149 1.13031
R17758 XThC.XTBN.Y.n137 XThC.XTBN.Y.n125 1.1255
R17759 XThC.XTBN.Y.n79 XThC.XTBN.Y 0.5125
R17760 XThC.XTBN.Y.n53 XThC.XTBN.Y 0.5125
R17761 XThC.XTBN.Y.n27 XThC.XTBN.Y 0.5125
R17762 XThC.XTBN.Y.n2 XThC.XTBN.Y 0.5125
R17763 XThC.XTBN.Y.n66 XThC.XTBN.Y 0.5125
R17764 XThC.XTBN.Y.n40 XThC.XTBN.Y 0.5125
R17765 XThC.XTBN.Y.n14 XThC.XTBN.Y 0.5125
R17766 XThC.Tn[6].n2 XThC.Tn[6].n1 332.332
R17767 XThC.Tn[6].n2 XThC.Tn[6].n0 296.493
R17768 XThC.Tn[6].n71 XThC.Tn[6].n69 161.365
R17769 XThC.Tn[6].n67 XThC.Tn[6].n65 161.365
R17770 XThC.Tn[6].n63 XThC.Tn[6].n61 161.365
R17771 XThC.Tn[6].n59 XThC.Tn[6].n57 161.365
R17772 XThC.Tn[6].n55 XThC.Tn[6].n53 161.365
R17773 XThC.Tn[6].n51 XThC.Tn[6].n49 161.365
R17774 XThC.Tn[6].n47 XThC.Tn[6].n45 161.365
R17775 XThC.Tn[6].n43 XThC.Tn[6].n41 161.365
R17776 XThC.Tn[6].n39 XThC.Tn[6].n37 161.365
R17777 XThC.Tn[6].n35 XThC.Tn[6].n33 161.365
R17778 XThC.Tn[6].n31 XThC.Tn[6].n29 161.365
R17779 XThC.Tn[6].n27 XThC.Tn[6].n25 161.365
R17780 XThC.Tn[6].n23 XThC.Tn[6].n21 161.365
R17781 XThC.Tn[6].n19 XThC.Tn[6].n17 161.365
R17782 XThC.Tn[6].n15 XThC.Tn[6].n13 161.365
R17783 XThC.Tn[6].n12 XThC.Tn[6].n10 161.365
R17784 XThC.Tn[6].n69 XThC.Tn[6].t34 161.202
R17785 XThC.Tn[6].n65 XThC.Tn[6].t24 161.202
R17786 XThC.Tn[6].n61 XThC.Tn[6].t43 161.202
R17787 XThC.Tn[6].n57 XThC.Tn[6].t41 161.202
R17788 XThC.Tn[6].n53 XThC.Tn[6].t32 161.202
R17789 XThC.Tn[6].n49 XThC.Tn[6].t21 161.202
R17790 XThC.Tn[6].n45 XThC.Tn[6].t19 161.202
R17791 XThC.Tn[6].n41 XThC.Tn[6].t31 161.202
R17792 XThC.Tn[6].n37 XThC.Tn[6].t29 161.202
R17793 XThC.Tn[6].n33 XThC.Tn[6].t22 161.202
R17794 XThC.Tn[6].n29 XThC.Tn[6].t38 161.202
R17795 XThC.Tn[6].n25 XThC.Tn[6].t37 161.202
R17796 XThC.Tn[6].n21 XThC.Tn[6].t18 161.202
R17797 XThC.Tn[6].n17 XThC.Tn[6].t17 161.202
R17798 XThC.Tn[6].n13 XThC.Tn[6].t13 161.202
R17799 XThC.Tn[6].n10 XThC.Tn[6].t26 161.202
R17800 XThC.Tn[6].n69 XThC.Tn[6].t30 145.137
R17801 XThC.Tn[6].n65 XThC.Tn[6].t20 145.137
R17802 XThC.Tn[6].n61 XThC.Tn[6].t39 145.137
R17803 XThC.Tn[6].n57 XThC.Tn[6].t36 145.137
R17804 XThC.Tn[6].n53 XThC.Tn[6].t28 145.137
R17805 XThC.Tn[6].n49 XThC.Tn[6].t15 145.137
R17806 XThC.Tn[6].n45 XThC.Tn[6].t14 145.137
R17807 XThC.Tn[6].n41 XThC.Tn[6].t27 145.137
R17808 XThC.Tn[6].n37 XThC.Tn[6].t25 145.137
R17809 XThC.Tn[6].n33 XThC.Tn[6].t16 145.137
R17810 XThC.Tn[6].n29 XThC.Tn[6].t35 145.137
R17811 XThC.Tn[6].n25 XThC.Tn[6].t33 145.137
R17812 XThC.Tn[6].n21 XThC.Tn[6].t12 145.137
R17813 XThC.Tn[6].n17 XThC.Tn[6].t42 145.137
R17814 XThC.Tn[6].n13 XThC.Tn[6].t40 145.137
R17815 XThC.Tn[6].n10 XThC.Tn[6].t23 145.137
R17816 XThC.Tn[6].n5 XThC.Tn[6].n3 135.248
R17817 XThC.Tn[6].n5 XThC.Tn[6].n4 98.982
R17818 XThC.Tn[6].n7 XThC.Tn[6].n6 98.982
R17819 XThC.Tn[6].n9 XThC.Tn[6].n8 98.982
R17820 XThC.Tn[6].n7 XThC.Tn[6].n5 36.2672
R17821 XThC.Tn[6].n9 XThC.Tn[6].n7 36.2672
R17822 XThC.Tn[6].n73 XThC.Tn[6].n9 32.6405
R17823 XThC.Tn[6].n1 XThC.Tn[6].t5 26.5955
R17824 XThC.Tn[6].n1 XThC.Tn[6].t4 26.5955
R17825 XThC.Tn[6].n0 XThC.Tn[6].t7 26.5955
R17826 XThC.Tn[6].n0 XThC.Tn[6].t6 26.5955
R17827 XThC.Tn[6].n3 XThC.Tn[6].t11 24.9236
R17828 XThC.Tn[6].n3 XThC.Tn[6].t10 24.9236
R17829 XThC.Tn[6].n4 XThC.Tn[6].t9 24.9236
R17830 XThC.Tn[6].n4 XThC.Tn[6].t8 24.9236
R17831 XThC.Tn[6].n6 XThC.Tn[6].t2 24.9236
R17832 XThC.Tn[6].n6 XThC.Tn[6].t1 24.9236
R17833 XThC.Tn[6].n8 XThC.Tn[6].t0 24.9236
R17834 XThC.Tn[6].n8 XThC.Tn[6].t3 24.9236
R17835 XThC.Tn[6].n74 XThC.Tn[6].n2 18.5605
R17836 XThC.Tn[6].n74 XThC.Tn[6].n73 11.5205
R17837 XThC.Tn[6] XThC.Tn[6].n12 8.0245
R17838 XThC.Tn[6].n72 XThC.Tn[6].n71 7.9105
R17839 XThC.Tn[6].n68 XThC.Tn[6].n67 7.9105
R17840 XThC.Tn[6].n64 XThC.Tn[6].n63 7.9105
R17841 XThC.Tn[6].n60 XThC.Tn[6].n59 7.9105
R17842 XThC.Tn[6].n56 XThC.Tn[6].n55 7.9105
R17843 XThC.Tn[6].n52 XThC.Tn[6].n51 7.9105
R17844 XThC.Tn[6].n48 XThC.Tn[6].n47 7.9105
R17845 XThC.Tn[6].n44 XThC.Tn[6].n43 7.9105
R17846 XThC.Tn[6].n40 XThC.Tn[6].n39 7.9105
R17847 XThC.Tn[6].n36 XThC.Tn[6].n35 7.9105
R17848 XThC.Tn[6].n32 XThC.Tn[6].n31 7.9105
R17849 XThC.Tn[6].n28 XThC.Tn[6].n27 7.9105
R17850 XThC.Tn[6].n24 XThC.Tn[6].n23 7.9105
R17851 XThC.Tn[6].n20 XThC.Tn[6].n19 7.9105
R17852 XThC.Tn[6].n16 XThC.Tn[6].n15 7.9105
R17853 XThC.Tn[6].n73 XThC.Tn[6] 5.42203
R17854 XThC.Tn[6] XThC.Tn[6].n74 0.6405
R17855 XThC.Tn[6].n16 XThC.Tn[6] 0.235138
R17856 XThC.Tn[6].n20 XThC.Tn[6] 0.235138
R17857 XThC.Tn[6].n24 XThC.Tn[6] 0.235138
R17858 XThC.Tn[6].n28 XThC.Tn[6] 0.235138
R17859 XThC.Tn[6].n32 XThC.Tn[6] 0.235138
R17860 XThC.Tn[6].n36 XThC.Tn[6] 0.235138
R17861 XThC.Tn[6].n40 XThC.Tn[6] 0.235138
R17862 XThC.Tn[6].n44 XThC.Tn[6] 0.235138
R17863 XThC.Tn[6].n48 XThC.Tn[6] 0.235138
R17864 XThC.Tn[6].n52 XThC.Tn[6] 0.235138
R17865 XThC.Tn[6].n56 XThC.Tn[6] 0.235138
R17866 XThC.Tn[6].n60 XThC.Tn[6] 0.235138
R17867 XThC.Tn[6].n64 XThC.Tn[6] 0.235138
R17868 XThC.Tn[6].n68 XThC.Tn[6] 0.235138
R17869 XThC.Tn[6].n72 XThC.Tn[6] 0.235138
R17870 XThC.Tn[6] XThC.Tn[6].n16 0.114505
R17871 XThC.Tn[6] XThC.Tn[6].n20 0.114505
R17872 XThC.Tn[6] XThC.Tn[6].n24 0.114505
R17873 XThC.Tn[6] XThC.Tn[6].n28 0.114505
R17874 XThC.Tn[6] XThC.Tn[6].n32 0.114505
R17875 XThC.Tn[6] XThC.Tn[6].n36 0.114505
R17876 XThC.Tn[6] XThC.Tn[6].n40 0.114505
R17877 XThC.Tn[6] XThC.Tn[6].n44 0.114505
R17878 XThC.Tn[6] XThC.Tn[6].n48 0.114505
R17879 XThC.Tn[6] XThC.Tn[6].n52 0.114505
R17880 XThC.Tn[6] XThC.Tn[6].n56 0.114505
R17881 XThC.Tn[6] XThC.Tn[6].n60 0.114505
R17882 XThC.Tn[6] XThC.Tn[6].n64 0.114505
R17883 XThC.Tn[6] XThC.Tn[6].n68 0.114505
R17884 XThC.Tn[6] XThC.Tn[6].n72 0.114505
R17885 XThC.Tn[6].n71 XThC.Tn[6].n70 0.0599512
R17886 XThC.Tn[6].n67 XThC.Tn[6].n66 0.0599512
R17887 XThC.Tn[6].n63 XThC.Tn[6].n62 0.0599512
R17888 XThC.Tn[6].n59 XThC.Tn[6].n58 0.0599512
R17889 XThC.Tn[6].n55 XThC.Tn[6].n54 0.0599512
R17890 XThC.Tn[6].n51 XThC.Tn[6].n50 0.0599512
R17891 XThC.Tn[6].n47 XThC.Tn[6].n46 0.0599512
R17892 XThC.Tn[6].n43 XThC.Tn[6].n42 0.0599512
R17893 XThC.Tn[6].n39 XThC.Tn[6].n38 0.0599512
R17894 XThC.Tn[6].n35 XThC.Tn[6].n34 0.0599512
R17895 XThC.Tn[6].n31 XThC.Tn[6].n30 0.0599512
R17896 XThC.Tn[6].n27 XThC.Tn[6].n26 0.0599512
R17897 XThC.Tn[6].n23 XThC.Tn[6].n22 0.0599512
R17898 XThC.Tn[6].n19 XThC.Tn[6].n18 0.0599512
R17899 XThC.Tn[6].n15 XThC.Tn[6].n14 0.0599512
R17900 XThC.Tn[6].n12 XThC.Tn[6].n11 0.0599512
R17901 XThC.Tn[6].n70 XThC.Tn[6] 0.0469286
R17902 XThC.Tn[6].n66 XThC.Tn[6] 0.0469286
R17903 XThC.Tn[6].n62 XThC.Tn[6] 0.0469286
R17904 XThC.Tn[6].n58 XThC.Tn[6] 0.0469286
R17905 XThC.Tn[6].n54 XThC.Tn[6] 0.0469286
R17906 XThC.Tn[6].n50 XThC.Tn[6] 0.0469286
R17907 XThC.Tn[6].n46 XThC.Tn[6] 0.0469286
R17908 XThC.Tn[6].n42 XThC.Tn[6] 0.0469286
R17909 XThC.Tn[6].n38 XThC.Tn[6] 0.0469286
R17910 XThC.Tn[6].n34 XThC.Tn[6] 0.0469286
R17911 XThC.Tn[6].n30 XThC.Tn[6] 0.0469286
R17912 XThC.Tn[6].n26 XThC.Tn[6] 0.0469286
R17913 XThC.Tn[6].n22 XThC.Tn[6] 0.0469286
R17914 XThC.Tn[6].n18 XThC.Tn[6] 0.0469286
R17915 XThC.Tn[6].n14 XThC.Tn[6] 0.0469286
R17916 XThC.Tn[6].n11 XThC.Tn[6] 0.0469286
R17917 XThC.Tn[6].n70 XThC.Tn[6] 0.0401341
R17918 XThC.Tn[6].n66 XThC.Tn[6] 0.0401341
R17919 XThC.Tn[6].n62 XThC.Tn[6] 0.0401341
R17920 XThC.Tn[6].n58 XThC.Tn[6] 0.0401341
R17921 XThC.Tn[6].n54 XThC.Tn[6] 0.0401341
R17922 XThC.Tn[6].n50 XThC.Tn[6] 0.0401341
R17923 XThC.Tn[6].n46 XThC.Tn[6] 0.0401341
R17924 XThC.Tn[6].n42 XThC.Tn[6] 0.0401341
R17925 XThC.Tn[6].n38 XThC.Tn[6] 0.0401341
R17926 XThC.Tn[6].n34 XThC.Tn[6] 0.0401341
R17927 XThC.Tn[6].n30 XThC.Tn[6] 0.0401341
R17928 XThC.Tn[6].n26 XThC.Tn[6] 0.0401341
R17929 XThC.Tn[6].n22 XThC.Tn[6] 0.0401341
R17930 XThC.Tn[6].n18 XThC.Tn[6] 0.0401341
R17931 XThC.Tn[6].n14 XThC.Tn[6] 0.0401341
R17932 XThC.Tn[6].n11 XThC.Tn[6] 0.0401341
R17933 XThR.Tn[9].n87 XThR.Tn[9].n86 256.103
R17934 XThR.Tn[9].n2 XThR.Tn[9].n0 243.68
R17935 XThR.Tn[9].n5 XThR.Tn[9].n3 241.847
R17936 XThR.Tn[9].n2 XThR.Tn[9].n1 205.28
R17937 XThR.Tn[9].n87 XThR.Tn[9].n85 202.094
R17938 XThR.Tn[9].n5 XThR.Tn[9].n4 185
R17939 XThR.Tn[9] XThR.Tn[9].n78 161.363
R17940 XThR.Tn[9] XThR.Tn[9].n73 161.363
R17941 XThR.Tn[9] XThR.Tn[9].n68 161.363
R17942 XThR.Tn[9] XThR.Tn[9].n63 161.363
R17943 XThR.Tn[9] XThR.Tn[9].n58 161.363
R17944 XThR.Tn[9] XThR.Tn[9].n53 161.363
R17945 XThR.Tn[9] XThR.Tn[9].n48 161.363
R17946 XThR.Tn[9] XThR.Tn[9].n43 161.363
R17947 XThR.Tn[9] XThR.Tn[9].n38 161.363
R17948 XThR.Tn[9] XThR.Tn[9].n33 161.363
R17949 XThR.Tn[9] XThR.Tn[9].n28 161.363
R17950 XThR.Tn[9] XThR.Tn[9].n23 161.363
R17951 XThR.Tn[9] XThR.Tn[9].n18 161.363
R17952 XThR.Tn[9] XThR.Tn[9].n13 161.363
R17953 XThR.Tn[9] XThR.Tn[9].n8 161.363
R17954 XThR.Tn[9] XThR.Tn[9].n6 161.363
R17955 XThR.Tn[9].n80 XThR.Tn[9].n79 161.3
R17956 XThR.Tn[9].n75 XThR.Tn[9].n74 161.3
R17957 XThR.Tn[9].n70 XThR.Tn[9].n69 161.3
R17958 XThR.Tn[9].n65 XThR.Tn[9].n64 161.3
R17959 XThR.Tn[9].n60 XThR.Tn[9].n59 161.3
R17960 XThR.Tn[9].n55 XThR.Tn[9].n54 161.3
R17961 XThR.Tn[9].n50 XThR.Tn[9].n49 161.3
R17962 XThR.Tn[9].n45 XThR.Tn[9].n44 161.3
R17963 XThR.Tn[9].n40 XThR.Tn[9].n39 161.3
R17964 XThR.Tn[9].n35 XThR.Tn[9].n34 161.3
R17965 XThR.Tn[9].n30 XThR.Tn[9].n29 161.3
R17966 XThR.Tn[9].n25 XThR.Tn[9].n24 161.3
R17967 XThR.Tn[9].n20 XThR.Tn[9].n19 161.3
R17968 XThR.Tn[9].n15 XThR.Tn[9].n14 161.3
R17969 XThR.Tn[9].n10 XThR.Tn[9].n9 161.3
R17970 XThR.Tn[9].n78 XThR.Tn[9].t63 161.106
R17971 XThR.Tn[9].n73 XThR.Tn[9].t69 161.106
R17972 XThR.Tn[9].n68 XThR.Tn[9].t47 161.106
R17973 XThR.Tn[9].n63 XThR.Tn[9].t34 161.106
R17974 XThR.Tn[9].n58 XThR.Tn[9].t62 161.106
R17975 XThR.Tn[9].n53 XThR.Tn[9].t24 161.106
R17976 XThR.Tn[9].n48 XThR.Tn[9].t66 161.106
R17977 XThR.Tn[9].n43 XThR.Tn[9].t45 161.106
R17978 XThR.Tn[9].n38 XThR.Tn[9].t32 161.106
R17979 XThR.Tn[9].n33 XThR.Tn[9].t37 161.106
R17980 XThR.Tn[9].n28 XThR.Tn[9].t23 161.106
R17981 XThR.Tn[9].n23 XThR.Tn[9].t46 161.106
R17982 XThR.Tn[9].n18 XThR.Tn[9].t21 161.106
R17983 XThR.Tn[9].n13 XThR.Tn[9].t64 161.106
R17984 XThR.Tn[9].n8 XThR.Tn[9].t28 161.106
R17985 XThR.Tn[9].n6 XThR.Tn[9].t71 161.106
R17986 XThR.Tn[9].n79 XThR.Tn[9].t54 159.978
R17987 XThR.Tn[9].n74 XThR.Tn[9].t61 159.978
R17988 XThR.Tn[9].n69 XThR.Tn[9].t43 159.978
R17989 XThR.Tn[9].n64 XThR.Tn[9].t27 159.978
R17990 XThR.Tn[9].n59 XThR.Tn[9].t52 159.978
R17991 XThR.Tn[9].n54 XThR.Tn[9].t18 159.978
R17992 XThR.Tn[9].n49 XThR.Tn[9].t60 159.978
R17993 XThR.Tn[9].n44 XThR.Tn[9].t40 159.978
R17994 XThR.Tn[9].n39 XThR.Tn[9].t25 159.978
R17995 XThR.Tn[9].n34 XThR.Tn[9].t33 159.978
R17996 XThR.Tn[9].n29 XThR.Tn[9].t16 159.978
R17997 XThR.Tn[9].n24 XThR.Tn[9].t42 159.978
R17998 XThR.Tn[9].n19 XThR.Tn[9].t15 159.978
R17999 XThR.Tn[9].n14 XThR.Tn[9].t59 159.978
R18000 XThR.Tn[9].n9 XThR.Tn[9].t19 159.978
R18001 XThR.Tn[9].n78 XThR.Tn[9].t49 145.038
R18002 XThR.Tn[9].n73 XThR.Tn[9].t14 145.038
R18003 XThR.Tn[9].n68 XThR.Tn[9].t57 145.038
R18004 XThR.Tn[9].n63 XThR.Tn[9].t38 145.038
R18005 XThR.Tn[9].n58 XThR.Tn[9].t70 145.038
R18006 XThR.Tn[9].n53 XThR.Tn[9].t48 145.038
R18007 XThR.Tn[9].n48 XThR.Tn[9].t58 145.038
R18008 XThR.Tn[9].n43 XThR.Tn[9].t39 145.038
R18009 XThR.Tn[9].n38 XThR.Tn[9].t36 145.038
R18010 XThR.Tn[9].n33 XThR.Tn[9].t67 145.038
R18011 XThR.Tn[9].n28 XThR.Tn[9].t31 145.038
R18012 XThR.Tn[9].n23 XThR.Tn[9].t56 145.038
R18013 XThR.Tn[9].n18 XThR.Tn[9].t29 145.038
R18014 XThR.Tn[9].n13 XThR.Tn[9].t72 145.038
R18015 XThR.Tn[9].n8 XThR.Tn[9].t35 145.038
R18016 XThR.Tn[9].n6 XThR.Tn[9].t17 145.038
R18017 XThR.Tn[9].n79 XThR.Tn[9].t68 143.911
R18018 XThR.Tn[9].n74 XThR.Tn[9].t30 143.911
R18019 XThR.Tn[9].n69 XThR.Tn[9].t12 143.911
R18020 XThR.Tn[9].n64 XThR.Tn[9].t53 143.911
R18021 XThR.Tn[9].n59 XThR.Tn[9].t22 143.911
R18022 XThR.Tn[9].n54 XThR.Tn[9].t65 143.911
R18023 XThR.Tn[9].n49 XThR.Tn[9].t13 143.911
R18024 XThR.Tn[9].n44 XThR.Tn[9].t55 143.911
R18025 XThR.Tn[9].n39 XThR.Tn[9].t51 143.911
R18026 XThR.Tn[9].n34 XThR.Tn[9].t20 143.911
R18027 XThR.Tn[9].n29 XThR.Tn[9].t44 143.911
R18028 XThR.Tn[9].n24 XThR.Tn[9].t73 143.911
R18029 XThR.Tn[9].n19 XThR.Tn[9].t41 143.911
R18030 XThR.Tn[9].n14 XThR.Tn[9].t26 143.911
R18031 XThR.Tn[9].n9 XThR.Tn[9].t50 143.911
R18032 XThR.Tn[9] XThR.Tn[9].n2 35.7652
R18033 XThR.Tn[9].n85 XThR.Tn[9].t2 26.5955
R18034 XThR.Tn[9].n85 XThR.Tn[9].t0 26.5955
R18035 XThR.Tn[9].n0 XThR.Tn[9].t10 26.5955
R18036 XThR.Tn[9].n0 XThR.Tn[9].t8 26.5955
R18037 XThR.Tn[9].n1 XThR.Tn[9].t11 26.5955
R18038 XThR.Tn[9].n1 XThR.Tn[9].t9 26.5955
R18039 XThR.Tn[9].n86 XThR.Tn[9].t3 26.5955
R18040 XThR.Tn[9].n86 XThR.Tn[9].t1 26.5955
R18041 XThR.Tn[9].n4 XThR.Tn[9].t4 24.9236
R18042 XThR.Tn[9].n4 XThR.Tn[9].t6 24.9236
R18043 XThR.Tn[9].n3 XThR.Tn[9].t5 24.9236
R18044 XThR.Tn[9].n3 XThR.Tn[9].t7 24.9236
R18045 XThR.Tn[9] XThR.Tn[9].n5 22.9615
R18046 XThR.Tn[9].n88 XThR.Tn[9].n87 13.5534
R18047 XThR.Tn[9].n84 XThR.Tn[9] 7.97984
R18048 XThR.Tn[9] XThR.Tn[9].n7 5.34038
R18049 XThR.Tn[9].n12 XThR.Tn[9].n11 4.5005
R18050 XThR.Tn[9].n17 XThR.Tn[9].n16 4.5005
R18051 XThR.Tn[9].n22 XThR.Tn[9].n21 4.5005
R18052 XThR.Tn[9].n27 XThR.Tn[9].n26 4.5005
R18053 XThR.Tn[9].n32 XThR.Tn[9].n31 4.5005
R18054 XThR.Tn[9].n37 XThR.Tn[9].n36 4.5005
R18055 XThR.Tn[9].n42 XThR.Tn[9].n41 4.5005
R18056 XThR.Tn[9].n47 XThR.Tn[9].n46 4.5005
R18057 XThR.Tn[9].n52 XThR.Tn[9].n51 4.5005
R18058 XThR.Tn[9].n57 XThR.Tn[9].n56 4.5005
R18059 XThR.Tn[9].n62 XThR.Tn[9].n61 4.5005
R18060 XThR.Tn[9].n67 XThR.Tn[9].n66 4.5005
R18061 XThR.Tn[9].n72 XThR.Tn[9].n71 4.5005
R18062 XThR.Tn[9].n77 XThR.Tn[9].n76 4.5005
R18063 XThR.Tn[9].n82 XThR.Tn[9].n81 4.5005
R18064 XThR.Tn[9].n83 XThR.Tn[9] 3.70586
R18065 XThR.Tn[9].n88 XThR.Tn[9].n84 2.99115
R18066 XThR.Tn[9].n88 XThR.Tn[9] 2.87153
R18067 XThR.Tn[9].n12 XThR.Tn[9] 2.52282
R18068 XThR.Tn[9].n17 XThR.Tn[9] 2.52282
R18069 XThR.Tn[9].n22 XThR.Tn[9] 2.52282
R18070 XThR.Tn[9].n27 XThR.Tn[9] 2.52282
R18071 XThR.Tn[9].n32 XThR.Tn[9] 2.52282
R18072 XThR.Tn[9].n37 XThR.Tn[9] 2.52282
R18073 XThR.Tn[9].n42 XThR.Tn[9] 2.52282
R18074 XThR.Tn[9].n47 XThR.Tn[9] 2.52282
R18075 XThR.Tn[9].n52 XThR.Tn[9] 2.52282
R18076 XThR.Tn[9].n57 XThR.Tn[9] 2.52282
R18077 XThR.Tn[9].n62 XThR.Tn[9] 2.52282
R18078 XThR.Tn[9].n67 XThR.Tn[9] 2.52282
R18079 XThR.Tn[9].n72 XThR.Tn[9] 2.52282
R18080 XThR.Tn[9].n77 XThR.Tn[9] 2.52282
R18081 XThR.Tn[9].n82 XThR.Tn[9] 2.52282
R18082 XThR.Tn[9].n84 XThR.Tn[9] 2.2734
R18083 XThR.Tn[9] XThR.Tn[9].n88 1.50638
R18084 XThR.Tn[9].n80 XThR.Tn[9] 1.08677
R18085 XThR.Tn[9].n75 XThR.Tn[9] 1.08677
R18086 XThR.Tn[9].n70 XThR.Tn[9] 1.08677
R18087 XThR.Tn[9].n65 XThR.Tn[9] 1.08677
R18088 XThR.Tn[9].n60 XThR.Tn[9] 1.08677
R18089 XThR.Tn[9].n55 XThR.Tn[9] 1.08677
R18090 XThR.Tn[9].n50 XThR.Tn[9] 1.08677
R18091 XThR.Tn[9].n45 XThR.Tn[9] 1.08677
R18092 XThR.Tn[9].n40 XThR.Tn[9] 1.08677
R18093 XThR.Tn[9].n35 XThR.Tn[9] 1.08677
R18094 XThR.Tn[9].n30 XThR.Tn[9] 1.08677
R18095 XThR.Tn[9].n25 XThR.Tn[9] 1.08677
R18096 XThR.Tn[9].n20 XThR.Tn[9] 1.08677
R18097 XThR.Tn[9].n15 XThR.Tn[9] 1.08677
R18098 XThR.Tn[9].n10 XThR.Tn[9] 1.08677
R18099 XThR.Tn[9] XThR.Tn[9].n12 0.839786
R18100 XThR.Tn[9] XThR.Tn[9].n17 0.839786
R18101 XThR.Tn[9] XThR.Tn[9].n22 0.839786
R18102 XThR.Tn[9] XThR.Tn[9].n27 0.839786
R18103 XThR.Tn[9] XThR.Tn[9].n32 0.839786
R18104 XThR.Tn[9] XThR.Tn[9].n37 0.839786
R18105 XThR.Tn[9] XThR.Tn[9].n42 0.839786
R18106 XThR.Tn[9] XThR.Tn[9].n47 0.839786
R18107 XThR.Tn[9] XThR.Tn[9].n52 0.839786
R18108 XThR.Tn[9] XThR.Tn[9].n57 0.839786
R18109 XThR.Tn[9] XThR.Tn[9].n62 0.839786
R18110 XThR.Tn[9] XThR.Tn[9].n67 0.839786
R18111 XThR.Tn[9] XThR.Tn[9].n72 0.839786
R18112 XThR.Tn[9] XThR.Tn[9].n77 0.839786
R18113 XThR.Tn[9] XThR.Tn[9].n82 0.839786
R18114 XThR.Tn[9].n7 XThR.Tn[9] 0.499542
R18115 XThR.Tn[9].n81 XThR.Tn[9] 0.063
R18116 XThR.Tn[9].n76 XThR.Tn[9] 0.063
R18117 XThR.Tn[9].n71 XThR.Tn[9] 0.063
R18118 XThR.Tn[9].n66 XThR.Tn[9] 0.063
R18119 XThR.Tn[9].n61 XThR.Tn[9] 0.063
R18120 XThR.Tn[9].n56 XThR.Tn[9] 0.063
R18121 XThR.Tn[9].n51 XThR.Tn[9] 0.063
R18122 XThR.Tn[9].n46 XThR.Tn[9] 0.063
R18123 XThR.Tn[9].n41 XThR.Tn[9] 0.063
R18124 XThR.Tn[9].n36 XThR.Tn[9] 0.063
R18125 XThR.Tn[9].n31 XThR.Tn[9] 0.063
R18126 XThR.Tn[9].n26 XThR.Tn[9] 0.063
R18127 XThR.Tn[9].n21 XThR.Tn[9] 0.063
R18128 XThR.Tn[9].n16 XThR.Tn[9] 0.063
R18129 XThR.Tn[9].n11 XThR.Tn[9] 0.063
R18130 XThR.Tn[9].n83 XThR.Tn[9] 0.0540714
R18131 XThR.Tn[9] XThR.Tn[9].n83 0.038
R18132 XThR.Tn[9].n7 XThR.Tn[9] 0.0143889
R18133 XThR.Tn[9].n81 XThR.Tn[9].n80 0.00771154
R18134 XThR.Tn[9].n76 XThR.Tn[9].n75 0.00771154
R18135 XThR.Tn[9].n71 XThR.Tn[9].n70 0.00771154
R18136 XThR.Tn[9].n66 XThR.Tn[9].n65 0.00771154
R18137 XThR.Tn[9].n61 XThR.Tn[9].n60 0.00771154
R18138 XThR.Tn[9].n56 XThR.Tn[9].n55 0.00771154
R18139 XThR.Tn[9].n51 XThR.Tn[9].n50 0.00771154
R18140 XThR.Tn[9].n46 XThR.Tn[9].n45 0.00771154
R18141 XThR.Tn[9].n41 XThR.Tn[9].n40 0.00771154
R18142 XThR.Tn[9].n36 XThR.Tn[9].n35 0.00771154
R18143 XThR.Tn[9].n31 XThR.Tn[9].n30 0.00771154
R18144 XThR.Tn[9].n26 XThR.Tn[9].n25 0.00771154
R18145 XThR.Tn[9].n21 XThR.Tn[9].n20 0.00771154
R18146 XThR.Tn[9].n16 XThR.Tn[9].n15 0.00771154
R18147 XThR.Tn[9].n11 XThR.Tn[9].n10 0.00771154
R18148 XThC.Tn[5].n2 XThC.Tn[5].n1 332.332
R18149 XThC.Tn[5].n2 XThC.Tn[5].n0 296.493
R18150 XThC.Tn[5].n71 XThC.Tn[5].n69 161.365
R18151 XThC.Tn[5].n67 XThC.Tn[5].n65 161.365
R18152 XThC.Tn[5].n63 XThC.Tn[5].n61 161.365
R18153 XThC.Tn[5].n59 XThC.Tn[5].n57 161.365
R18154 XThC.Tn[5].n55 XThC.Tn[5].n53 161.365
R18155 XThC.Tn[5].n51 XThC.Tn[5].n49 161.365
R18156 XThC.Tn[5].n47 XThC.Tn[5].n45 161.365
R18157 XThC.Tn[5].n43 XThC.Tn[5].n41 161.365
R18158 XThC.Tn[5].n39 XThC.Tn[5].n37 161.365
R18159 XThC.Tn[5].n35 XThC.Tn[5].n33 161.365
R18160 XThC.Tn[5].n31 XThC.Tn[5].n29 161.365
R18161 XThC.Tn[5].n27 XThC.Tn[5].n25 161.365
R18162 XThC.Tn[5].n23 XThC.Tn[5].n21 161.365
R18163 XThC.Tn[5].n19 XThC.Tn[5].n17 161.365
R18164 XThC.Tn[5].n15 XThC.Tn[5].n13 161.365
R18165 XThC.Tn[5].n12 XThC.Tn[5].n10 161.365
R18166 XThC.Tn[5].n69 XThC.Tn[5].t41 161.202
R18167 XThC.Tn[5].n65 XThC.Tn[5].t30 161.202
R18168 XThC.Tn[5].n61 XThC.Tn[5].t18 161.202
R18169 XThC.Tn[5].n57 XThC.Tn[5].t16 161.202
R18170 XThC.Tn[5].n53 XThC.Tn[5].t39 161.202
R18171 XThC.Tn[5].n49 XThC.Tn[5].t26 161.202
R18172 XThC.Tn[5].n45 XThC.Tn[5].t25 161.202
R18173 XThC.Tn[5].n41 XThC.Tn[5].t37 161.202
R18174 XThC.Tn[5].n37 XThC.Tn[5].t35 161.202
R18175 XThC.Tn[5].n33 XThC.Tn[5].t27 161.202
R18176 XThC.Tn[5].n29 XThC.Tn[5].t14 161.202
R18177 XThC.Tn[5].n25 XThC.Tn[5].t13 161.202
R18178 XThC.Tn[5].n21 XThC.Tn[5].t24 161.202
R18179 XThC.Tn[5].n17 XThC.Tn[5].t23 161.202
R18180 XThC.Tn[5].n13 XThC.Tn[5].t19 161.202
R18181 XThC.Tn[5].n10 XThC.Tn[5].t33 161.202
R18182 XThC.Tn[5].n69 XThC.Tn[5].t22 145.137
R18183 XThC.Tn[5].n65 XThC.Tn[5].t12 145.137
R18184 XThC.Tn[5].n61 XThC.Tn[5].t32 145.137
R18185 XThC.Tn[5].n57 XThC.Tn[5].t31 145.137
R18186 XThC.Tn[5].n53 XThC.Tn[5].t21 145.137
R18187 XThC.Tn[5].n49 XThC.Tn[5].t42 145.137
R18188 XThC.Tn[5].n45 XThC.Tn[5].t40 145.137
R18189 XThC.Tn[5].n41 XThC.Tn[5].t20 145.137
R18190 XThC.Tn[5].n37 XThC.Tn[5].t17 145.137
R18191 XThC.Tn[5].n33 XThC.Tn[5].t43 145.137
R18192 XThC.Tn[5].n29 XThC.Tn[5].t29 145.137
R18193 XThC.Tn[5].n25 XThC.Tn[5].t28 145.137
R18194 XThC.Tn[5].n21 XThC.Tn[5].t38 145.137
R18195 XThC.Tn[5].n17 XThC.Tn[5].t36 145.137
R18196 XThC.Tn[5].n13 XThC.Tn[5].t34 145.137
R18197 XThC.Tn[5].n10 XThC.Tn[5].t15 145.137
R18198 XThC.Tn[5].n6 XThC.Tn[5].n4 135.249
R18199 XThC.Tn[5].n9 XThC.Tn[5].n3 98.981
R18200 XThC.Tn[5].n6 XThC.Tn[5].n5 98.981
R18201 XThC.Tn[5].n8 XThC.Tn[5].n7 98.981
R18202 XThC.Tn[5].n8 XThC.Tn[5].n6 36.2672
R18203 XThC.Tn[5].n9 XThC.Tn[5].n8 36.2672
R18204 XThC.Tn[5].n73 XThC.Tn[5].n9 32.6405
R18205 XThC.Tn[5].n1 XThC.Tn[5].t5 26.5955
R18206 XThC.Tn[5].n1 XThC.Tn[5].t4 26.5955
R18207 XThC.Tn[5].n0 XThC.Tn[5].t7 26.5955
R18208 XThC.Tn[5].n0 XThC.Tn[5].t6 26.5955
R18209 XThC.Tn[5].n3 XThC.Tn[5].t1 24.9236
R18210 XThC.Tn[5].n3 XThC.Tn[5].t0 24.9236
R18211 XThC.Tn[5].n4 XThC.Tn[5].t8 24.9236
R18212 XThC.Tn[5].n4 XThC.Tn[5].t11 24.9236
R18213 XThC.Tn[5].n5 XThC.Tn[5].t10 24.9236
R18214 XThC.Tn[5].n5 XThC.Tn[5].t9 24.9236
R18215 XThC.Tn[5].n7 XThC.Tn[5].t3 24.9236
R18216 XThC.Tn[5].n7 XThC.Tn[5].t2 24.9236
R18217 XThC.Tn[5] XThC.Tn[5].n2 23.3605
R18218 XThC.Tn[5] XThC.Tn[5].n12 8.0245
R18219 XThC.Tn[5].n72 XThC.Tn[5].n71 7.9105
R18220 XThC.Tn[5].n68 XThC.Tn[5].n67 7.9105
R18221 XThC.Tn[5].n64 XThC.Tn[5].n63 7.9105
R18222 XThC.Tn[5].n60 XThC.Tn[5].n59 7.9105
R18223 XThC.Tn[5].n56 XThC.Tn[5].n55 7.9105
R18224 XThC.Tn[5].n52 XThC.Tn[5].n51 7.9105
R18225 XThC.Tn[5].n48 XThC.Tn[5].n47 7.9105
R18226 XThC.Tn[5].n44 XThC.Tn[5].n43 7.9105
R18227 XThC.Tn[5].n40 XThC.Tn[5].n39 7.9105
R18228 XThC.Tn[5].n36 XThC.Tn[5].n35 7.9105
R18229 XThC.Tn[5].n32 XThC.Tn[5].n31 7.9105
R18230 XThC.Tn[5].n28 XThC.Tn[5].n27 7.9105
R18231 XThC.Tn[5].n24 XThC.Tn[5].n23 7.9105
R18232 XThC.Tn[5].n20 XThC.Tn[5].n19 7.9105
R18233 XThC.Tn[5].n16 XThC.Tn[5].n15 7.9105
R18234 XThC.Tn[5] XThC.Tn[5].n73 6.7205
R18235 XThC.Tn[5].n73 XThC.Tn[5] 5.69842
R18236 XThC.Tn[5].n16 XThC.Tn[5] 0.235138
R18237 XThC.Tn[5].n20 XThC.Tn[5] 0.235138
R18238 XThC.Tn[5].n24 XThC.Tn[5] 0.235138
R18239 XThC.Tn[5].n28 XThC.Tn[5] 0.235138
R18240 XThC.Tn[5].n32 XThC.Tn[5] 0.235138
R18241 XThC.Tn[5].n36 XThC.Tn[5] 0.235138
R18242 XThC.Tn[5].n40 XThC.Tn[5] 0.235138
R18243 XThC.Tn[5].n44 XThC.Tn[5] 0.235138
R18244 XThC.Tn[5].n48 XThC.Tn[5] 0.235138
R18245 XThC.Tn[5].n52 XThC.Tn[5] 0.235138
R18246 XThC.Tn[5].n56 XThC.Tn[5] 0.235138
R18247 XThC.Tn[5].n60 XThC.Tn[5] 0.235138
R18248 XThC.Tn[5].n64 XThC.Tn[5] 0.235138
R18249 XThC.Tn[5].n68 XThC.Tn[5] 0.235138
R18250 XThC.Tn[5].n72 XThC.Tn[5] 0.235138
R18251 XThC.Tn[5] XThC.Tn[5].n16 0.114505
R18252 XThC.Tn[5] XThC.Tn[5].n20 0.114505
R18253 XThC.Tn[5] XThC.Tn[5].n24 0.114505
R18254 XThC.Tn[5] XThC.Tn[5].n28 0.114505
R18255 XThC.Tn[5] XThC.Tn[5].n32 0.114505
R18256 XThC.Tn[5] XThC.Tn[5].n36 0.114505
R18257 XThC.Tn[5] XThC.Tn[5].n40 0.114505
R18258 XThC.Tn[5] XThC.Tn[5].n44 0.114505
R18259 XThC.Tn[5] XThC.Tn[5].n48 0.114505
R18260 XThC.Tn[5] XThC.Tn[5].n52 0.114505
R18261 XThC.Tn[5] XThC.Tn[5].n56 0.114505
R18262 XThC.Tn[5] XThC.Tn[5].n60 0.114505
R18263 XThC.Tn[5] XThC.Tn[5].n64 0.114505
R18264 XThC.Tn[5] XThC.Tn[5].n68 0.114505
R18265 XThC.Tn[5] XThC.Tn[5].n72 0.114505
R18266 XThC.Tn[5].n71 XThC.Tn[5].n70 0.0599512
R18267 XThC.Tn[5].n67 XThC.Tn[5].n66 0.0599512
R18268 XThC.Tn[5].n63 XThC.Tn[5].n62 0.0599512
R18269 XThC.Tn[5].n59 XThC.Tn[5].n58 0.0599512
R18270 XThC.Tn[5].n55 XThC.Tn[5].n54 0.0599512
R18271 XThC.Tn[5].n51 XThC.Tn[5].n50 0.0599512
R18272 XThC.Tn[5].n47 XThC.Tn[5].n46 0.0599512
R18273 XThC.Tn[5].n43 XThC.Tn[5].n42 0.0599512
R18274 XThC.Tn[5].n39 XThC.Tn[5].n38 0.0599512
R18275 XThC.Tn[5].n35 XThC.Tn[5].n34 0.0599512
R18276 XThC.Tn[5].n31 XThC.Tn[5].n30 0.0599512
R18277 XThC.Tn[5].n27 XThC.Tn[5].n26 0.0599512
R18278 XThC.Tn[5].n23 XThC.Tn[5].n22 0.0599512
R18279 XThC.Tn[5].n19 XThC.Tn[5].n18 0.0599512
R18280 XThC.Tn[5].n15 XThC.Tn[5].n14 0.0599512
R18281 XThC.Tn[5].n12 XThC.Tn[5].n11 0.0599512
R18282 XThC.Tn[5].n70 XThC.Tn[5] 0.0469286
R18283 XThC.Tn[5].n66 XThC.Tn[5] 0.0469286
R18284 XThC.Tn[5].n62 XThC.Tn[5] 0.0469286
R18285 XThC.Tn[5].n58 XThC.Tn[5] 0.0469286
R18286 XThC.Tn[5].n54 XThC.Tn[5] 0.0469286
R18287 XThC.Tn[5].n50 XThC.Tn[5] 0.0469286
R18288 XThC.Tn[5].n46 XThC.Tn[5] 0.0469286
R18289 XThC.Tn[5].n42 XThC.Tn[5] 0.0469286
R18290 XThC.Tn[5].n38 XThC.Tn[5] 0.0469286
R18291 XThC.Tn[5].n34 XThC.Tn[5] 0.0469286
R18292 XThC.Tn[5].n30 XThC.Tn[5] 0.0469286
R18293 XThC.Tn[5].n26 XThC.Tn[5] 0.0469286
R18294 XThC.Tn[5].n22 XThC.Tn[5] 0.0469286
R18295 XThC.Tn[5].n18 XThC.Tn[5] 0.0469286
R18296 XThC.Tn[5].n14 XThC.Tn[5] 0.0469286
R18297 XThC.Tn[5].n11 XThC.Tn[5] 0.0469286
R18298 XThC.Tn[5].n70 XThC.Tn[5] 0.0401341
R18299 XThC.Tn[5].n66 XThC.Tn[5] 0.0401341
R18300 XThC.Tn[5].n62 XThC.Tn[5] 0.0401341
R18301 XThC.Tn[5].n58 XThC.Tn[5] 0.0401341
R18302 XThC.Tn[5].n54 XThC.Tn[5] 0.0401341
R18303 XThC.Tn[5].n50 XThC.Tn[5] 0.0401341
R18304 XThC.Tn[5].n46 XThC.Tn[5] 0.0401341
R18305 XThC.Tn[5].n42 XThC.Tn[5] 0.0401341
R18306 XThC.Tn[5].n38 XThC.Tn[5] 0.0401341
R18307 XThC.Tn[5].n34 XThC.Tn[5] 0.0401341
R18308 XThC.Tn[5].n30 XThC.Tn[5] 0.0401341
R18309 XThC.Tn[5].n26 XThC.Tn[5] 0.0401341
R18310 XThC.Tn[5].n22 XThC.Tn[5] 0.0401341
R18311 XThC.Tn[5].n18 XThC.Tn[5] 0.0401341
R18312 XThC.Tn[5].n14 XThC.Tn[5] 0.0401341
R18313 XThC.Tn[5].n11 XThC.Tn[5] 0.0401341
R18314 XThC.Tn[9].n70 XThC.Tn[9].n69 265.341
R18315 XThC.Tn[9].n74 XThC.Tn[9].n72 243.68
R18316 XThC.Tn[9].n2 XThC.Tn[9].n0 241.847
R18317 XThC.Tn[9].n74 XThC.Tn[9].n73 205.28
R18318 XThC.Tn[9].n70 XThC.Tn[9].n68 202.094
R18319 XThC.Tn[9].n2 XThC.Tn[9].n1 185
R18320 XThC.Tn[9].n64 XThC.Tn[9].n62 161.365
R18321 XThC.Tn[9].n60 XThC.Tn[9].n58 161.365
R18322 XThC.Tn[9].n56 XThC.Tn[9].n54 161.365
R18323 XThC.Tn[9].n52 XThC.Tn[9].n50 161.365
R18324 XThC.Tn[9].n48 XThC.Tn[9].n46 161.365
R18325 XThC.Tn[9].n44 XThC.Tn[9].n42 161.365
R18326 XThC.Tn[9].n40 XThC.Tn[9].n38 161.365
R18327 XThC.Tn[9].n36 XThC.Tn[9].n34 161.365
R18328 XThC.Tn[9].n32 XThC.Tn[9].n30 161.365
R18329 XThC.Tn[9].n28 XThC.Tn[9].n26 161.365
R18330 XThC.Tn[9].n24 XThC.Tn[9].n22 161.365
R18331 XThC.Tn[9].n20 XThC.Tn[9].n18 161.365
R18332 XThC.Tn[9].n16 XThC.Tn[9].n14 161.365
R18333 XThC.Tn[9].n12 XThC.Tn[9].n10 161.365
R18334 XThC.Tn[9].n8 XThC.Tn[9].n6 161.365
R18335 XThC.Tn[9].n5 XThC.Tn[9].n3 161.365
R18336 XThC.Tn[9].n62 XThC.Tn[9].t20 161.202
R18337 XThC.Tn[9].n58 XThC.Tn[9].t41 161.202
R18338 XThC.Tn[9].n54 XThC.Tn[9].t29 161.202
R18339 XThC.Tn[9].n50 XThC.Tn[9].t27 161.202
R18340 XThC.Tn[9].n46 XThC.Tn[9].t18 161.202
R18341 XThC.Tn[9].n42 XThC.Tn[9].t37 161.202
R18342 XThC.Tn[9].n38 XThC.Tn[9].t36 161.202
R18343 XThC.Tn[9].n34 XThC.Tn[9].t16 161.202
R18344 XThC.Tn[9].n30 XThC.Tn[9].t14 161.202
R18345 XThC.Tn[9].n26 XThC.Tn[9].t38 161.202
R18346 XThC.Tn[9].n22 XThC.Tn[9].t25 161.202
R18347 XThC.Tn[9].n18 XThC.Tn[9].t24 161.202
R18348 XThC.Tn[9].n14 XThC.Tn[9].t35 161.202
R18349 XThC.Tn[9].n10 XThC.Tn[9].t34 161.202
R18350 XThC.Tn[9].n6 XThC.Tn[9].t30 161.202
R18351 XThC.Tn[9].n3 XThC.Tn[9].t12 161.202
R18352 XThC.Tn[9].n62 XThC.Tn[9].t33 145.137
R18353 XThC.Tn[9].n58 XThC.Tn[9].t23 145.137
R18354 XThC.Tn[9].n54 XThC.Tn[9].t43 145.137
R18355 XThC.Tn[9].n50 XThC.Tn[9].t42 145.137
R18356 XThC.Tn[9].n46 XThC.Tn[9].t32 145.137
R18357 XThC.Tn[9].n42 XThC.Tn[9].t21 145.137
R18358 XThC.Tn[9].n38 XThC.Tn[9].t19 145.137
R18359 XThC.Tn[9].n34 XThC.Tn[9].t31 145.137
R18360 XThC.Tn[9].n30 XThC.Tn[9].t28 145.137
R18361 XThC.Tn[9].n26 XThC.Tn[9].t22 145.137
R18362 XThC.Tn[9].n22 XThC.Tn[9].t40 145.137
R18363 XThC.Tn[9].n18 XThC.Tn[9].t39 145.137
R18364 XThC.Tn[9].n14 XThC.Tn[9].t17 145.137
R18365 XThC.Tn[9].n10 XThC.Tn[9].t15 145.137
R18366 XThC.Tn[9].n6 XThC.Tn[9].t13 145.137
R18367 XThC.Tn[9].n3 XThC.Tn[9].t26 145.137
R18368 XThC.Tn[9].n72 XThC.Tn[9].t1 26.5955
R18369 XThC.Tn[9].n72 XThC.Tn[9].t0 26.5955
R18370 XThC.Tn[9].n69 XThC.Tn[9].t6 26.5955
R18371 XThC.Tn[9].n69 XThC.Tn[9].t5 26.5955
R18372 XThC.Tn[9].n68 XThC.Tn[9].t4 26.5955
R18373 XThC.Tn[9].n68 XThC.Tn[9].t7 26.5955
R18374 XThC.Tn[9].n73 XThC.Tn[9].t3 26.5955
R18375 XThC.Tn[9].n73 XThC.Tn[9].t2 26.5955
R18376 XThC.Tn[9].n1 XThC.Tn[9].t10 24.9236
R18377 XThC.Tn[9].n1 XThC.Tn[9].t11 24.9236
R18378 XThC.Tn[9].n0 XThC.Tn[9].t9 24.9236
R18379 XThC.Tn[9].n0 XThC.Tn[9].t8 24.9236
R18380 XThC.Tn[9] XThC.Tn[9].n74 22.9652
R18381 XThC.Tn[9] XThC.Tn[9].n2 18.8943
R18382 XThC.Tn[9].n71 XThC.Tn[9].n70 13.9299
R18383 XThC.Tn[9] XThC.Tn[9].n71 13.9299
R18384 XThC.Tn[9] XThC.Tn[9].n5 8.0245
R18385 XThC.Tn[9].n65 XThC.Tn[9].n64 7.9105
R18386 XThC.Tn[9].n61 XThC.Tn[9].n60 7.9105
R18387 XThC.Tn[9].n57 XThC.Tn[9].n56 7.9105
R18388 XThC.Tn[9].n53 XThC.Tn[9].n52 7.9105
R18389 XThC.Tn[9].n49 XThC.Tn[9].n48 7.9105
R18390 XThC.Tn[9].n45 XThC.Tn[9].n44 7.9105
R18391 XThC.Tn[9].n41 XThC.Tn[9].n40 7.9105
R18392 XThC.Tn[9].n37 XThC.Tn[9].n36 7.9105
R18393 XThC.Tn[9].n33 XThC.Tn[9].n32 7.9105
R18394 XThC.Tn[9].n29 XThC.Tn[9].n28 7.9105
R18395 XThC.Tn[9].n25 XThC.Tn[9].n24 7.9105
R18396 XThC.Tn[9].n21 XThC.Tn[9].n20 7.9105
R18397 XThC.Tn[9].n17 XThC.Tn[9].n16 7.9105
R18398 XThC.Tn[9].n13 XThC.Tn[9].n12 7.9105
R18399 XThC.Tn[9].n9 XThC.Tn[9].n8 7.9105
R18400 XThC.Tn[9].n67 XThC.Tn[9].n66 7.44831
R18401 XThC.Tn[9].n67 XThC.Tn[9] 6.34069
R18402 XThC.Tn[9].n66 XThC.Tn[9] 4.25199
R18403 XThC.Tn[9] XThC.Tn[9].n67 1.79489
R18404 XThC.Tn[9].n71 XThC.Tn[9] 1.19676
R18405 XThC.Tn[9].n66 XThC.Tn[9] 0.657022
R18406 XThC.Tn[9].n9 XThC.Tn[9] 0.235138
R18407 XThC.Tn[9].n13 XThC.Tn[9] 0.235138
R18408 XThC.Tn[9].n17 XThC.Tn[9] 0.235138
R18409 XThC.Tn[9].n21 XThC.Tn[9] 0.235138
R18410 XThC.Tn[9].n25 XThC.Tn[9] 0.235138
R18411 XThC.Tn[9].n29 XThC.Tn[9] 0.235138
R18412 XThC.Tn[9].n33 XThC.Tn[9] 0.235138
R18413 XThC.Tn[9].n37 XThC.Tn[9] 0.235138
R18414 XThC.Tn[9].n41 XThC.Tn[9] 0.235138
R18415 XThC.Tn[9].n45 XThC.Tn[9] 0.235138
R18416 XThC.Tn[9].n49 XThC.Tn[9] 0.235138
R18417 XThC.Tn[9].n53 XThC.Tn[9] 0.235138
R18418 XThC.Tn[9].n57 XThC.Tn[9] 0.235138
R18419 XThC.Tn[9].n61 XThC.Tn[9] 0.235138
R18420 XThC.Tn[9].n65 XThC.Tn[9] 0.235138
R18421 XThC.Tn[9] XThC.Tn[9].n9 0.114505
R18422 XThC.Tn[9] XThC.Tn[9].n13 0.114505
R18423 XThC.Tn[9] XThC.Tn[9].n17 0.114505
R18424 XThC.Tn[9] XThC.Tn[9].n21 0.114505
R18425 XThC.Tn[9] XThC.Tn[9].n25 0.114505
R18426 XThC.Tn[9] XThC.Tn[9].n29 0.114505
R18427 XThC.Tn[9] XThC.Tn[9].n33 0.114505
R18428 XThC.Tn[9] XThC.Tn[9].n37 0.114505
R18429 XThC.Tn[9] XThC.Tn[9].n41 0.114505
R18430 XThC.Tn[9] XThC.Tn[9].n45 0.114505
R18431 XThC.Tn[9] XThC.Tn[9].n49 0.114505
R18432 XThC.Tn[9] XThC.Tn[9].n53 0.114505
R18433 XThC.Tn[9] XThC.Tn[9].n57 0.114505
R18434 XThC.Tn[9] XThC.Tn[9].n61 0.114505
R18435 XThC.Tn[9] XThC.Tn[9].n65 0.114505
R18436 XThC.Tn[9].n64 XThC.Tn[9].n63 0.0599512
R18437 XThC.Tn[9].n60 XThC.Tn[9].n59 0.0599512
R18438 XThC.Tn[9].n56 XThC.Tn[9].n55 0.0599512
R18439 XThC.Tn[9].n52 XThC.Tn[9].n51 0.0599512
R18440 XThC.Tn[9].n48 XThC.Tn[9].n47 0.0599512
R18441 XThC.Tn[9].n44 XThC.Tn[9].n43 0.0599512
R18442 XThC.Tn[9].n40 XThC.Tn[9].n39 0.0599512
R18443 XThC.Tn[9].n36 XThC.Tn[9].n35 0.0599512
R18444 XThC.Tn[9].n32 XThC.Tn[9].n31 0.0599512
R18445 XThC.Tn[9].n28 XThC.Tn[9].n27 0.0599512
R18446 XThC.Tn[9].n24 XThC.Tn[9].n23 0.0599512
R18447 XThC.Tn[9].n20 XThC.Tn[9].n19 0.0599512
R18448 XThC.Tn[9].n16 XThC.Tn[9].n15 0.0599512
R18449 XThC.Tn[9].n12 XThC.Tn[9].n11 0.0599512
R18450 XThC.Tn[9].n8 XThC.Tn[9].n7 0.0599512
R18451 XThC.Tn[9].n5 XThC.Tn[9].n4 0.0599512
R18452 XThC.Tn[9].n63 XThC.Tn[9] 0.0469286
R18453 XThC.Tn[9].n59 XThC.Tn[9] 0.0469286
R18454 XThC.Tn[9].n55 XThC.Tn[9] 0.0469286
R18455 XThC.Tn[9].n51 XThC.Tn[9] 0.0469286
R18456 XThC.Tn[9].n47 XThC.Tn[9] 0.0469286
R18457 XThC.Tn[9].n43 XThC.Tn[9] 0.0469286
R18458 XThC.Tn[9].n39 XThC.Tn[9] 0.0469286
R18459 XThC.Tn[9].n35 XThC.Tn[9] 0.0469286
R18460 XThC.Tn[9].n31 XThC.Tn[9] 0.0469286
R18461 XThC.Tn[9].n27 XThC.Tn[9] 0.0469286
R18462 XThC.Tn[9].n23 XThC.Tn[9] 0.0469286
R18463 XThC.Tn[9].n19 XThC.Tn[9] 0.0469286
R18464 XThC.Tn[9].n15 XThC.Tn[9] 0.0469286
R18465 XThC.Tn[9].n11 XThC.Tn[9] 0.0469286
R18466 XThC.Tn[9].n7 XThC.Tn[9] 0.0469286
R18467 XThC.Tn[9].n4 XThC.Tn[9] 0.0469286
R18468 XThC.Tn[9].n63 XThC.Tn[9] 0.0401341
R18469 XThC.Tn[9].n59 XThC.Tn[9] 0.0401341
R18470 XThC.Tn[9].n55 XThC.Tn[9] 0.0401341
R18471 XThC.Tn[9].n51 XThC.Tn[9] 0.0401341
R18472 XThC.Tn[9].n47 XThC.Tn[9] 0.0401341
R18473 XThC.Tn[9].n43 XThC.Tn[9] 0.0401341
R18474 XThC.Tn[9].n39 XThC.Tn[9] 0.0401341
R18475 XThC.Tn[9].n35 XThC.Tn[9] 0.0401341
R18476 XThC.Tn[9].n31 XThC.Tn[9] 0.0401341
R18477 XThC.Tn[9].n27 XThC.Tn[9] 0.0401341
R18478 XThC.Tn[9].n23 XThC.Tn[9] 0.0401341
R18479 XThC.Tn[9].n19 XThC.Tn[9] 0.0401341
R18480 XThC.Tn[9].n15 XThC.Tn[9] 0.0401341
R18481 XThC.Tn[9].n11 XThC.Tn[9] 0.0401341
R18482 XThC.Tn[9].n7 XThC.Tn[9] 0.0401341
R18483 XThC.Tn[9].n4 XThC.Tn[9] 0.0401341
R18484 XThC.Tn[11].n70 XThC.Tn[11].n69 265.341
R18485 XThC.Tn[11].n74 XThC.Tn[11].n73 243.68
R18486 XThC.Tn[11].n2 XThC.Tn[11].n0 241.847
R18487 XThC.Tn[11].n74 XThC.Tn[11].n72 205.28
R18488 XThC.Tn[11].n70 XThC.Tn[11].n68 202.094
R18489 XThC.Tn[11].n2 XThC.Tn[11].n1 185
R18490 XThC.Tn[11].n64 XThC.Tn[11].n62 161.365
R18491 XThC.Tn[11].n60 XThC.Tn[11].n58 161.365
R18492 XThC.Tn[11].n56 XThC.Tn[11].n54 161.365
R18493 XThC.Tn[11].n52 XThC.Tn[11].n50 161.365
R18494 XThC.Tn[11].n48 XThC.Tn[11].n46 161.365
R18495 XThC.Tn[11].n44 XThC.Tn[11].n42 161.365
R18496 XThC.Tn[11].n40 XThC.Tn[11].n38 161.365
R18497 XThC.Tn[11].n36 XThC.Tn[11].n34 161.365
R18498 XThC.Tn[11].n32 XThC.Tn[11].n30 161.365
R18499 XThC.Tn[11].n28 XThC.Tn[11].n26 161.365
R18500 XThC.Tn[11].n24 XThC.Tn[11].n22 161.365
R18501 XThC.Tn[11].n20 XThC.Tn[11].n18 161.365
R18502 XThC.Tn[11].n16 XThC.Tn[11].n14 161.365
R18503 XThC.Tn[11].n12 XThC.Tn[11].n10 161.365
R18504 XThC.Tn[11].n8 XThC.Tn[11].n6 161.365
R18505 XThC.Tn[11].n5 XThC.Tn[11].n3 161.365
R18506 XThC.Tn[11].n62 XThC.Tn[11].t24 161.202
R18507 XThC.Tn[11].n58 XThC.Tn[11].t14 161.202
R18508 XThC.Tn[11].n54 XThC.Tn[11].t33 161.202
R18509 XThC.Tn[11].n50 XThC.Tn[11].t30 161.202
R18510 XThC.Tn[11].n46 XThC.Tn[11].t22 161.202
R18511 XThC.Tn[11].n42 XThC.Tn[11].t41 161.202
R18512 XThC.Tn[11].n38 XThC.Tn[11].t40 161.202
R18513 XThC.Tn[11].n34 XThC.Tn[11].t21 161.202
R18514 XThC.Tn[11].n30 XThC.Tn[11].t19 161.202
R18515 XThC.Tn[11].n26 XThC.Tn[11].t42 161.202
R18516 XThC.Tn[11].n22 XThC.Tn[11].t29 161.202
R18517 XThC.Tn[11].n18 XThC.Tn[11].t28 161.202
R18518 XThC.Tn[11].n14 XThC.Tn[11].t39 161.202
R18519 XThC.Tn[11].n10 XThC.Tn[11].t37 161.202
R18520 XThC.Tn[11].n6 XThC.Tn[11].t35 161.202
R18521 XThC.Tn[11].n3 XThC.Tn[11].t18 161.202
R18522 XThC.Tn[11].n62 XThC.Tn[11].t27 145.137
R18523 XThC.Tn[11].n58 XThC.Tn[11].t17 145.137
R18524 XThC.Tn[11].n54 XThC.Tn[11].t36 145.137
R18525 XThC.Tn[11].n50 XThC.Tn[11].t34 145.137
R18526 XThC.Tn[11].n46 XThC.Tn[11].t26 145.137
R18527 XThC.Tn[11].n42 XThC.Tn[11].t15 145.137
R18528 XThC.Tn[11].n38 XThC.Tn[11].t13 145.137
R18529 XThC.Tn[11].n34 XThC.Tn[11].t25 145.137
R18530 XThC.Tn[11].n30 XThC.Tn[11].t23 145.137
R18531 XThC.Tn[11].n26 XThC.Tn[11].t16 145.137
R18532 XThC.Tn[11].n22 XThC.Tn[11].t32 145.137
R18533 XThC.Tn[11].n18 XThC.Tn[11].t31 145.137
R18534 XThC.Tn[11].n14 XThC.Tn[11].t12 145.137
R18535 XThC.Tn[11].n10 XThC.Tn[11].t43 145.137
R18536 XThC.Tn[11].n6 XThC.Tn[11].t38 145.137
R18537 XThC.Tn[11].n3 XThC.Tn[11].t20 145.137
R18538 XThC.Tn[11].n69 XThC.Tn[11].t4 26.5955
R18539 XThC.Tn[11].n69 XThC.Tn[11].t9 26.5955
R18540 XThC.Tn[11].n68 XThC.Tn[11].t6 26.5955
R18541 XThC.Tn[11].n68 XThC.Tn[11].t10 26.5955
R18542 XThC.Tn[11].n72 XThC.Tn[11].t2 26.5955
R18543 XThC.Tn[11].n72 XThC.Tn[11].t1 26.5955
R18544 XThC.Tn[11].n73 XThC.Tn[11].t0 26.5955
R18545 XThC.Tn[11].n73 XThC.Tn[11].t3 26.5955
R18546 XThC.Tn[11].n1 XThC.Tn[11].t7 24.9236
R18547 XThC.Tn[11].n1 XThC.Tn[11].t5 24.9236
R18548 XThC.Tn[11].n0 XThC.Tn[11].t8 24.9236
R18549 XThC.Tn[11].n0 XThC.Tn[11].t11 24.9236
R18550 XThC.Tn[11] XThC.Tn[11].n74 22.9652
R18551 XThC.Tn[11] XThC.Tn[11].n2 18.8943
R18552 XThC.Tn[11].n71 XThC.Tn[11].n70 13.9299
R18553 XThC.Tn[11] XThC.Tn[11].n71 13.9299
R18554 XThC.Tn[11] XThC.Tn[11].n5 8.0245
R18555 XThC.Tn[11].n65 XThC.Tn[11].n64 7.9105
R18556 XThC.Tn[11].n61 XThC.Tn[11].n60 7.9105
R18557 XThC.Tn[11].n57 XThC.Tn[11].n56 7.9105
R18558 XThC.Tn[11].n53 XThC.Tn[11].n52 7.9105
R18559 XThC.Tn[11].n49 XThC.Tn[11].n48 7.9105
R18560 XThC.Tn[11].n45 XThC.Tn[11].n44 7.9105
R18561 XThC.Tn[11].n41 XThC.Tn[11].n40 7.9105
R18562 XThC.Tn[11].n37 XThC.Tn[11].n36 7.9105
R18563 XThC.Tn[11].n33 XThC.Tn[11].n32 7.9105
R18564 XThC.Tn[11].n29 XThC.Tn[11].n28 7.9105
R18565 XThC.Tn[11].n25 XThC.Tn[11].n24 7.9105
R18566 XThC.Tn[11].n21 XThC.Tn[11].n20 7.9105
R18567 XThC.Tn[11].n17 XThC.Tn[11].n16 7.9105
R18568 XThC.Tn[11].n13 XThC.Tn[11].n12 7.9105
R18569 XThC.Tn[11].n9 XThC.Tn[11].n8 7.9105
R18570 XThC.Tn[11].n67 XThC.Tn[11].n66 7.44831
R18571 XThC.Tn[11].n67 XThC.Tn[11] 6.34069
R18572 XThC.Tn[11].n66 XThC.Tn[11] 4.37928
R18573 XThC.Tn[11] XThC.Tn[11].n67 1.79489
R18574 XThC.Tn[11].n71 XThC.Tn[11] 1.19676
R18575 XThC.Tn[11].n66 XThC.Tn[11] 1.0918
R18576 XThC.Tn[11].n9 XThC.Tn[11] 0.235138
R18577 XThC.Tn[11].n13 XThC.Tn[11] 0.235138
R18578 XThC.Tn[11].n17 XThC.Tn[11] 0.235138
R18579 XThC.Tn[11].n21 XThC.Tn[11] 0.235138
R18580 XThC.Tn[11].n25 XThC.Tn[11] 0.235138
R18581 XThC.Tn[11].n29 XThC.Tn[11] 0.235138
R18582 XThC.Tn[11].n33 XThC.Tn[11] 0.235138
R18583 XThC.Tn[11].n37 XThC.Tn[11] 0.235138
R18584 XThC.Tn[11].n41 XThC.Tn[11] 0.235138
R18585 XThC.Tn[11].n45 XThC.Tn[11] 0.235138
R18586 XThC.Tn[11].n49 XThC.Tn[11] 0.235138
R18587 XThC.Tn[11].n53 XThC.Tn[11] 0.235138
R18588 XThC.Tn[11].n57 XThC.Tn[11] 0.235138
R18589 XThC.Tn[11].n61 XThC.Tn[11] 0.235138
R18590 XThC.Tn[11].n65 XThC.Tn[11] 0.235138
R18591 XThC.Tn[11] XThC.Tn[11].n9 0.114505
R18592 XThC.Tn[11] XThC.Tn[11].n13 0.114505
R18593 XThC.Tn[11] XThC.Tn[11].n17 0.114505
R18594 XThC.Tn[11] XThC.Tn[11].n21 0.114505
R18595 XThC.Tn[11] XThC.Tn[11].n25 0.114505
R18596 XThC.Tn[11] XThC.Tn[11].n29 0.114505
R18597 XThC.Tn[11] XThC.Tn[11].n33 0.114505
R18598 XThC.Tn[11] XThC.Tn[11].n37 0.114505
R18599 XThC.Tn[11] XThC.Tn[11].n41 0.114505
R18600 XThC.Tn[11] XThC.Tn[11].n45 0.114505
R18601 XThC.Tn[11] XThC.Tn[11].n49 0.114505
R18602 XThC.Tn[11] XThC.Tn[11].n53 0.114505
R18603 XThC.Tn[11] XThC.Tn[11].n57 0.114505
R18604 XThC.Tn[11] XThC.Tn[11].n61 0.114505
R18605 XThC.Tn[11] XThC.Tn[11].n65 0.114505
R18606 XThC.Tn[11].n64 XThC.Tn[11].n63 0.0599512
R18607 XThC.Tn[11].n60 XThC.Tn[11].n59 0.0599512
R18608 XThC.Tn[11].n56 XThC.Tn[11].n55 0.0599512
R18609 XThC.Tn[11].n52 XThC.Tn[11].n51 0.0599512
R18610 XThC.Tn[11].n48 XThC.Tn[11].n47 0.0599512
R18611 XThC.Tn[11].n44 XThC.Tn[11].n43 0.0599512
R18612 XThC.Tn[11].n40 XThC.Tn[11].n39 0.0599512
R18613 XThC.Tn[11].n36 XThC.Tn[11].n35 0.0599512
R18614 XThC.Tn[11].n32 XThC.Tn[11].n31 0.0599512
R18615 XThC.Tn[11].n28 XThC.Tn[11].n27 0.0599512
R18616 XThC.Tn[11].n24 XThC.Tn[11].n23 0.0599512
R18617 XThC.Tn[11].n20 XThC.Tn[11].n19 0.0599512
R18618 XThC.Tn[11].n16 XThC.Tn[11].n15 0.0599512
R18619 XThC.Tn[11].n12 XThC.Tn[11].n11 0.0599512
R18620 XThC.Tn[11].n8 XThC.Tn[11].n7 0.0599512
R18621 XThC.Tn[11].n5 XThC.Tn[11].n4 0.0599512
R18622 XThC.Tn[11].n63 XThC.Tn[11] 0.0469286
R18623 XThC.Tn[11].n59 XThC.Tn[11] 0.0469286
R18624 XThC.Tn[11].n55 XThC.Tn[11] 0.0469286
R18625 XThC.Tn[11].n51 XThC.Tn[11] 0.0469286
R18626 XThC.Tn[11].n47 XThC.Tn[11] 0.0469286
R18627 XThC.Tn[11].n43 XThC.Tn[11] 0.0469286
R18628 XThC.Tn[11].n39 XThC.Tn[11] 0.0469286
R18629 XThC.Tn[11].n35 XThC.Tn[11] 0.0469286
R18630 XThC.Tn[11].n31 XThC.Tn[11] 0.0469286
R18631 XThC.Tn[11].n27 XThC.Tn[11] 0.0469286
R18632 XThC.Tn[11].n23 XThC.Tn[11] 0.0469286
R18633 XThC.Tn[11].n19 XThC.Tn[11] 0.0469286
R18634 XThC.Tn[11].n15 XThC.Tn[11] 0.0469286
R18635 XThC.Tn[11].n11 XThC.Tn[11] 0.0469286
R18636 XThC.Tn[11].n7 XThC.Tn[11] 0.0469286
R18637 XThC.Tn[11].n4 XThC.Tn[11] 0.0469286
R18638 XThC.Tn[11].n63 XThC.Tn[11] 0.0401341
R18639 XThC.Tn[11].n59 XThC.Tn[11] 0.0401341
R18640 XThC.Tn[11].n55 XThC.Tn[11] 0.0401341
R18641 XThC.Tn[11].n51 XThC.Tn[11] 0.0401341
R18642 XThC.Tn[11].n47 XThC.Tn[11] 0.0401341
R18643 XThC.Tn[11].n43 XThC.Tn[11] 0.0401341
R18644 XThC.Tn[11].n39 XThC.Tn[11] 0.0401341
R18645 XThC.Tn[11].n35 XThC.Tn[11] 0.0401341
R18646 XThC.Tn[11].n31 XThC.Tn[11] 0.0401341
R18647 XThC.Tn[11].n27 XThC.Tn[11] 0.0401341
R18648 XThC.Tn[11].n23 XThC.Tn[11] 0.0401341
R18649 XThC.Tn[11].n19 XThC.Tn[11] 0.0401341
R18650 XThC.Tn[11].n15 XThC.Tn[11] 0.0401341
R18651 XThC.Tn[11].n11 XThC.Tn[11] 0.0401341
R18652 XThC.Tn[11].n7 XThC.Tn[11] 0.0401341
R18653 XThC.Tn[11].n4 XThC.Tn[11] 0.0401341
R18654 XThC.Tn[12].n70 XThC.Tn[12].n69 256.103
R18655 XThC.Tn[12].n74 XThC.Tn[12].n72 243.68
R18656 XThC.Tn[12].n2 XThC.Tn[12].n0 241.847
R18657 XThC.Tn[12].n74 XThC.Tn[12].n73 205.28
R18658 XThC.Tn[12].n70 XThC.Tn[12].n68 202.095
R18659 XThC.Tn[12].n2 XThC.Tn[12].n1 185
R18660 XThC.Tn[12].n64 XThC.Tn[12].n62 161.365
R18661 XThC.Tn[12].n60 XThC.Tn[12].n58 161.365
R18662 XThC.Tn[12].n56 XThC.Tn[12].n54 161.365
R18663 XThC.Tn[12].n52 XThC.Tn[12].n50 161.365
R18664 XThC.Tn[12].n48 XThC.Tn[12].n46 161.365
R18665 XThC.Tn[12].n44 XThC.Tn[12].n42 161.365
R18666 XThC.Tn[12].n40 XThC.Tn[12].n38 161.365
R18667 XThC.Tn[12].n36 XThC.Tn[12].n34 161.365
R18668 XThC.Tn[12].n32 XThC.Tn[12].n30 161.365
R18669 XThC.Tn[12].n28 XThC.Tn[12].n26 161.365
R18670 XThC.Tn[12].n24 XThC.Tn[12].n22 161.365
R18671 XThC.Tn[12].n20 XThC.Tn[12].n18 161.365
R18672 XThC.Tn[12].n16 XThC.Tn[12].n14 161.365
R18673 XThC.Tn[12].n12 XThC.Tn[12].n10 161.365
R18674 XThC.Tn[12].n8 XThC.Tn[12].n6 161.365
R18675 XThC.Tn[12].n5 XThC.Tn[12].n3 161.365
R18676 XThC.Tn[12].n62 XThC.Tn[12].t41 161.202
R18677 XThC.Tn[12].n58 XThC.Tn[12].t31 161.202
R18678 XThC.Tn[12].n54 XThC.Tn[12].t18 161.202
R18679 XThC.Tn[12].n50 XThC.Tn[12].t15 161.202
R18680 XThC.Tn[12].n46 XThC.Tn[12].t39 161.202
R18681 XThC.Tn[12].n42 XThC.Tn[12].t26 161.202
R18682 XThC.Tn[12].n38 XThC.Tn[12].t25 161.202
R18683 XThC.Tn[12].n34 XThC.Tn[12].t38 161.202
R18684 XThC.Tn[12].n30 XThC.Tn[12].t36 161.202
R18685 XThC.Tn[12].n26 XThC.Tn[12].t27 161.202
R18686 XThC.Tn[12].n22 XThC.Tn[12].t14 161.202
R18687 XThC.Tn[12].n18 XThC.Tn[12].t13 161.202
R18688 XThC.Tn[12].n14 XThC.Tn[12].t24 161.202
R18689 XThC.Tn[12].n10 XThC.Tn[12].t22 161.202
R18690 XThC.Tn[12].n6 XThC.Tn[12].t20 161.202
R18691 XThC.Tn[12].n3 XThC.Tn[12].t35 161.202
R18692 XThC.Tn[12].n62 XThC.Tn[12].t12 145.137
R18693 XThC.Tn[12].n58 XThC.Tn[12].t34 145.137
R18694 XThC.Tn[12].n54 XThC.Tn[12].t21 145.137
R18695 XThC.Tn[12].n50 XThC.Tn[12].t19 145.137
R18696 XThC.Tn[12].n46 XThC.Tn[12].t43 145.137
R18697 XThC.Tn[12].n42 XThC.Tn[12].t32 145.137
R18698 XThC.Tn[12].n38 XThC.Tn[12].t30 145.137
R18699 XThC.Tn[12].n34 XThC.Tn[12].t42 145.137
R18700 XThC.Tn[12].n30 XThC.Tn[12].t40 145.137
R18701 XThC.Tn[12].n26 XThC.Tn[12].t33 145.137
R18702 XThC.Tn[12].n22 XThC.Tn[12].t17 145.137
R18703 XThC.Tn[12].n18 XThC.Tn[12].t16 145.137
R18704 XThC.Tn[12].n14 XThC.Tn[12].t29 145.137
R18705 XThC.Tn[12].n10 XThC.Tn[12].t28 145.137
R18706 XThC.Tn[12].n6 XThC.Tn[12].t23 145.137
R18707 XThC.Tn[12].n3 XThC.Tn[12].t37 145.137
R18708 XThC.Tn[12].n68 XThC.Tn[12].t1 26.5955
R18709 XThC.Tn[12].n68 XThC.Tn[12].t2 26.5955
R18710 XThC.Tn[12].n72 XThC.Tn[12].t9 26.5955
R18711 XThC.Tn[12].n72 XThC.Tn[12].t8 26.5955
R18712 XThC.Tn[12].n73 XThC.Tn[12].t11 26.5955
R18713 XThC.Tn[12].n73 XThC.Tn[12].t10 26.5955
R18714 XThC.Tn[12].n69 XThC.Tn[12].t0 26.5955
R18715 XThC.Tn[12].n69 XThC.Tn[12].t3 26.5955
R18716 XThC.Tn[12].n1 XThC.Tn[12].t5 24.9236
R18717 XThC.Tn[12].n1 XThC.Tn[12].t4 24.9236
R18718 XThC.Tn[12].n0 XThC.Tn[12].t7 24.9236
R18719 XThC.Tn[12].n0 XThC.Tn[12].t6 24.9236
R18720 XThC.Tn[12] XThC.Tn[12].n74 22.9652
R18721 XThC.Tn[12] XThC.Tn[12].n2 22.9615
R18722 XThC.Tn[12].n71 XThC.Tn[12].n70 13.9299
R18723 XThC.Tn[12] XThC.Tn[12].n71 13.9299
R18724 XThC.Tn[12] XThC.Tn[12].n5 8.0245
R18725 XThC.Tn[12].n65 XThC.Tn[12].n64 7.9105
R18726 XThC.Tn[12].n61 XThC.Tn[12].n60 7.9105
R18727 XThC.Tn[12].n57 XThC.Tn[12].n56 7.9105
R18728 XThC.Tn[12].n53 XThC.Tn[12].n52 7.9105
R18729 XThC.Tn[12].n49 XThC.Tn[12].n48 7.9105
R18730 XThC.Tn[12].n45 XThC.Tn[12].n44 7.9105
R18731 XThC.Tn[12].n41 XThC.Tn[12].n40 7.9105
R18732 XThC.Tn[12].n37 XThC.Tn[12].n36 7.9105
R18733 XThC.Tn[12].n33 XThC.Tn[12].n32 7.9105
R18734 XThC.Tn[12].n29 XThC.Tn[12].n28 7.9105
R18735 XThC.Tn[12].n25 XThC.Tn[12].n24 7.9105
R18736 XThC.Tn[12].n21 XThC.Tn[12].n20 7.9105
R18737 XThC.Tn[12].n17 XThC.Tn[12].n16 7.9105
R18738 XThC.Tn[12].n13 XThC.Tn[12].n12 7.9105
R18739 XThC.Tn[12].n9 XThC.Tn[12].n8 7.9105
R18740 XThC.Tn[12].n67 XThC.Tn[12].n66 7.4309
R18741 XThC.Tn[12].n66 XThC.Tn[12] 4.71945
R18742 XThC.Tn[12].n71 XThC.Tn[12].n67 2.99115
R18743 XThC.Tn[12].n71 XThC.Tn[12] 2.87153
R18744 XThC.Tn[12].n67 XThC.Tn[12] 2.2734
R18745 XThC.Tn[12].n66 XThC.Tn[12] 0.88175
R18746 XThC.Tn[12].n9 XThC.Tn[12] 0.235138
R18747 XThC.Tn[12].n13 XThC.Tn[12] 0.235138
R18748 XThC.Tn[12].n17 XThC.Tn[12] 0.235138
R18749 XThC.Tn[12].n21 XThC.Tn[12] 0.235138
R18750 XThC.Tn[12].n25 XThC.Tn[12] 0.235138
R18751 XThC.Tn[12].n29 XThC.Tn[12] 0.235138
R18752 XThC.Tn[12].n33 XThC.Tn[12] 0.235138
R18753 XThC.Tn[12].n37 XThC.Tn[12] 0.235138
R18754 XThC.Tn[12].n41 XThC.Tn[12] 0.235138
R18755 XThC.Tn[12].n45 XThC.Tn[12] 0.235138
R18756 XThC.Tn[12].n49 XThC.Tn[12] 0.235138
R18757 XThC.Tn[12].n53 XThC.Tn[12] 0.235138
R18758 XThC.Tn[12].n57 XThC.Tn[12] 0.235138
R18759 XThC.Tn[12].n61 XThC.Tn[12] 0.235138
R18760 XThC.Tn[12].n65 XThC.Tn[12] 0.235138
R18761 XThC.Tn[12] XThC.Tn[12].n9 0.114505
R18762 XThC.Tn[12] XThC.Tn[12].n13 0.114505
R18763 XThC.Tn[12] XThC.Tn[12].n17 0.114505
R18764 XThC.Tn[12] XThC.Tn[12].n21 0.114505
R18765 XThC.Tn[12] XThC.Tn[12].n25 0.114505
R18766 XThC.Tn[12] XThC.Tn[12].n29 0.114505
R18767 XThC.Tn[12] XThC.Tn[12].n33 0.114505
R18768 XThC.Tn[12] XThC.Tn[12].n37 0.114505
R18769 XThC.Tn[12] XThC.Tn[12].n41 0.114505
R18770 XThC.Tn[12] XThC.Tn[12].n45 0.114505
R18771 XThC.Tn[12] XThC.Tn[12].n49 0.114505
R18772 XThC.Tn[12] XThC.Tn[12].n53 0.114505
R18773 XThC.Tn[12] XThC.Tn[12].n57 0.114505
R18774 XThC.Tn[12] XThC.Tn[12].n61 0.114505
R18775 XThC.Tn[12] XThC.Tn[12].n65 0.114505
R18776 XThC.Tn[12].n64 XThC.Tn[12].n63 0.0599512
R18777 XThC.Tn[12].n60 XThC.Tn[12].n59 0.0599512
R18778 XThC.Tn[12].n56 XThC.Tn[12].n55 0.0599512
R18779 XThC.Tn[12].n52 XThC.Tn[12].n51 0.0599512
R18780 XThC.Tn[12].n48 XThC.Tn[12].n47 0.0599512
R18781 XThC.Tn[12].n44 XThC.Tn[12].n43 0.0599512
R18782 XThC.Tn[12].n40 XThC.Tn[12].n39 0.0599512
R18783 XThC.Tn[12].n36 XThC.Tn[12].n35 0.0599512
R18784 XThC.Tn[12].n32 XThC.Tn[12].n31 0.0599512
R18785 XThC.Tn[12].n28 XThC.Tn[12].n27 0.0599512
R18786 XThC.Tn[12].n24 XThC.Tn[12].n23 0.0599512
R18787 XThC.Tn[12].n20 XThC.Tn[12].n19 0.0599512
R18788 XThC.Tn[12].n16 XThC.Tn[12].n15 0.0599512
R18789 XThC.Tn[12].n12 XThC.Tn[12].n11 0.0599512
R18790 XThC.Tn[12].n8 XThC.Tn[12].n7 0.0599512
R18791 XThC.Tn[12].n5 XThC.Tn[12].n4 0.0599512
R18792 XThC.Tn[12].n63 XThC.Tn[12] 0.0469286
R18793 XThC.Tn[12].n59 XThC.Tn[12] 0.0469286
R18794 XThC.Tn[12].n55 XThC.Tn[12] 0.0469286
R18795 XThC.Tn[12].n51 XThC.Tn[12] 0.0469286
R18796 XThC.Tn[12].n47 XThC.Tn[12] 0.0469286
R18797 XThC.Tn[12].n43 XThC.Tn[12] 0.0469286
R18798 XThC.Tn[12].n39 XThC.Tn[12] 0.0469286
R18799 XThC.Tn[12].n35 XThC.Tn[12] 0.0469286
R18800 XThC.Tn[12].n31 XThC.Tn[12] 0.0469286
R18801 XThC.Tn[12].n27 XThC.Tn[12] 0.0469286
R18802 XThC.Tn[12].n23 XThC.Tn[12] 0.0469286
R18803 XThC.Tn[12].n19 XThC.Tn[12] 0.0469286
R18804 XThC.Tn[12].n15 XThC.Tn[12] 0.0469286
R18805 XThC.Tn[12].n11 XThC.Tn[12] 0.0469286
R18806 XThC.Tn[12].n7 XThC.Tn[12] 0.0469286
R18807 XThC.Tn[12].n4 XThC.Tn[12] 0.0469286
R18808 XThC.Tn[12].n63 XThC.Tn[12] 0.0401341
R18809 XThC.Tn[12].n59 XThC.Tn[12] 0.0401341
R18810 XThC.Tn[12].n55 XThC.Tn[12] 0.0401341
R18811 XThC.Tn[12].n51 XThC.Tn[12] 0.0401341
R18812 XThC.Tn[12].n47 XThC.Tn[12] 0.0401341
R18813 XThC.Tn[12].n43 XThC.Tn[12] 0.0401341
R18814 XThC.Tn[12].n39 XThC.Tn[12] 0.0401341
R18815 XThC.Tn[12].n35 XThC.Tn[12] 0.0401341
R18816 XThC.Tn[12].n31 XThC.Tn[12] 0.0401341
R18817 XThC.Tn[12].n27 XThC.Tn[12] 0.0401341
R18818 XThC.Tn[12].n23 XThC.Tn[12] 0.0401341
R18819 XThC.Tn[12].n19 XThC.Tn[12] 0.0401341
R18820 XThC.Tn[12].n15 XThC.Tn[12] 0.0401341
R18821 XThC.Tn[12].n11 XThC.Tn[12] 0.0401341
R18822 XThC.Tn[12].n7 XThC.Tn[12] 0.0401341
R18823 XThC.Tn[12].n4 XThC.Tn[12] 0.0401341
R18824 XThC.Tn[13].n70 XThC.Tn[13].n69 265.341
R18825 XThC.Tn[13].n74 XThC.Tn[13].n72 243.68
R18826 XThC.Tn[13].n2 XThC.Tn[13].n0 241.847
R18827 XThC.Tn[13].n74 XThC.Tn[13].n73 205.28
R18828 XThC.Tn[13].n70 XThC.Tn[13].n68 202.094
R18829 XThC.Tn[13].n2 XThC.Tn[13].n1 185
R18830 XThC.Tn[13].n64 XThC.Tn[13].n62 161.365
R18831 XThC.Tn[13].n60 XThC.Tn[13].n58 161.365
R18832 XThC.Tn[13].n56 XThC.Tn[13].n54 161.365
R18833 XThC.Tn[13].n52 XThC.Tn[13].n50 161.365
R18834 XThC.Tn[13].n48 XThC.Tn[13].n46 161.365
R18835 XThC.Tn[13].n44 XThC.Tn[13].n42 161.365
R18836 XThC.Tn[13].n40 XThC.Tn[13].n38 161.365
R18837 XThC.Tn[13].n36 XThC.Tn[13].n34 161.365
R18838 XThC.Tn[13].n32 XThC.Tn[13].n30 161.365
R18839 XThC.Tn[13].n28 XThC.Tn[13].n26 161.365
R18840 XThC.Tn[13].n24 XThC.Tn[13].n22 161.365
R18841 XThC.Tn[13].n20 XThC.Tn[13].n18 161.365
R18842 XThC.Tn[13].n16 XThC.Tn[13].n14 161.365
R18843 XThC.Tn[13].n12 XThC.Tn[13].n10 161.365
R18844 XThC.Tn[13].n8 XThC.Tn[13].n6 161.365
R18845 XThC.Tn[13].n5 XThC.Tn[13].n3 161.365
R18846 XThC.Tn[13].n62 XThC.Tn[13].t33 161.202
R18847 XThC.Tn[13].n58 XThC.Tn[13].t23 161.202
R18848 XThC.Tn[13].n54 XThC.Tn[13].t42 161.202
R18849 XThC.Tn[13].n50 XThC.Tn[13].t39 161.202
R18850 XThC.Tn[13].n46 XThC.Tn[13].t31 161.202
R18851 XThC.Tn[13].n42 XThC.Tn[13].t18 161.202
R18852 XThC.Tn[13].n38 XThC.Tn[13].t17 161.202
R18853 XThC.Tn[13].n34 XThC.Tn[13].t30 161.202
R18854 XThC.Tn[13].n30 XThC.Tn[13].t28 161.202
R18855 XThC.Tn[13].n26 XThC.Tn[13].t19 161.202
R18856 XThC.Tn[13].n22 XThC.Tn[13].t38 161.202
R18857 XThC.Tn[13].n18 XThC.Tn[13].t37 161.202
R18858 XThC.Tn[13].n14 XThC.Tn[13].t16 161.202
R18859 XThC.Tn[13].n10 XThC.Tn[13].t14 161.202
R18860 XThC.Tn[13].n6 XThC.Tn[13].t12 161.202
R18861 XThC.Tn[13].n3 XThC.Tn[13].t27 161.202
R18862 XThC.Tn[13].n62 XThC.Tn[13].t36 145.137
R18863 XThC.Tn[13].n58 XThC.Tn[13].t26 145.137
R18864 XThC.Tn[13].n54 XThC.Tn[13].t13 145.137
R18865 XThC.Tn[13].n50 XThC.Tn[13].t43 145.137
R18866 XThC.Tn[13].n46 XThC.Tn[13].t35 145.137
R18867 XThC.Tn[13].n42 XThC.Tn[13].t24 145.137
R18868 XThC.Tn[13].n38 XThC.Tn[13].t22 145.137
R18869 XThC.Tn[13].n34 XThC.Tn[13].t34 145.137
R18870 XThC.Tn[13].n30 XThC.Tn[13].t32 145.137
R18871 XThC.Tn[13].n26 XThC.Tn[13].t25 145.137
R18872 XThC.Tn[13].n22 XThC.Tn[13].t41 145.137
R18873 XThC.Tn[13].n18 XThC.Tn[13].t40 145.137
R18874 XThC.Tn[13].n14 XThC.Tn[13].t21 145.137
R18875 XThC.Tn[13].n10 XThC.Tn[13].t20 145.137
R18876 XThC.Tn[13].n6 XThC.Tn[13].t15 145.137
R18877 XThC.Tn[13].n3 XThC.Tn[13].t29 145.137
R18878 XThC.Tn[13].n72 XThC.Tn[13].t1 26.5955
R18879 XThC.Tn[13].n72 XThC.Tn[13].t0 26.5955
R18880 XThC.Tn[13].n69 XThC.Tn[13].t4 26.5955
R18881 XThC.Tn[13].n69 XThC.Tn[13].t7 26.5955
R18882 XThC.Tn[13].n68 XThC.Tn[13].t6 26.5955
R18883 XThC.Tn[13].n68 XThC.Tn[13].t5 26.5955
R18884 XThC.Tn[13].n73 XThC.Tn[13].t3 26.5955
R18885 XThC.Tn[13].n73 XThC.Tn[13].t2 26.5955
R18886 XThC.Tn[13].n1 XThC.Tn[13].t8 24.9236
R18887 XThC.Tn[13].n1 XThC.Tn[13].t10 24.9236
R18888 XThC.Tn[13].n0 XThC.Tn[13].t11 24.9236
R18889 XThC.Tn[13].n0 XThC.Tn[13].t9 24.9236
R18890 XThC.Tn[13] XThC.Tn[13].n74 22.9652
R18891 XThC.Tn[13] XThC.Tn[13].n2 18.8943
R18892 XThC.Tn[13].n71 XThC.Tn[13].n70 13.9299
R18893 XThC.Tn[13] XThC.Tn[13].n71 13.9299
R18894 XThC.Tn[13] XThC.Tn[13].n5 8.0245
R18895 XThC.Tn[13].n65 XThC.Tn[13].n64 7.9105
R18896 XThC.Tn[13].n61 XThC.Tn[13].n60 7.9105
R18897 XThC.Tn[13].n57 XThC.Tn[13].n56 7.9105
R18898 XThC.Tn[13].n53 XThC.Tn[13].n52 7.9105
R18899 XThC.Tn[13].n49 XThC.Tn[13].n48 7.9105
R18900 XThC.Tn[13].n45 XThC.Tn[13].n44 7.9105
R18901 XThC.Tn[13].n41 XThC.Tn[13].n40 7.9105
R18902 XThC.Tn[13].n37 XThC.Tn[13].n36 7.9105
R18903 XThC.Tn[13].n33 XThC.Tn[13].n32 7.9105
R18904 XThC.Tn[13].n29 XThC.Tn[13].n28 7.9105
R18905 XThC.Tn[13].n25 XThC.Tn[13].n24 7.9105
R18906 XThC.Tn[13].n21 XThC.Tn[13].n20 7.9105
R18907 XThC.Tn[13].n17 XThC.Tn[13].n16 7.9105
R18908 XThC.Tn[13].n13 XThC.Tn[13].n12 7.9105
R18909 XThC.Tn[13].n9 XThC.Tn[13].n8 7.9105
R18910 XThC.Tn[13].n67 XThC.Tn[13].n66 7.46054
R18911 XThC.Tn[13].n67 XThC.Tn[13] 6.34069
R18912 XThC.Tn[13].n66 XThC.Tn[13] 4.78838
R18913 XThC.Tn[13] XThC.Tn[13].n67 1.79489
R18914 XThC.Tn[13].n66 XThC.Tn[13] 1.51436
R18915 XThC.Tn[13].n71 XThC.Tn[13] 1.19676
R18916 XThC.Tn[13].n9 XThC.Tn[13] 0.235138
R18917 XThC.Tn[13].n13 XThC.Tn[13] 0.235138
R18918 XThC.Tn[13].n17 XThC.Tn[13] 0.235138
R18919 XThC.Tn[13].n21 XThC.Tn[13] 0.235138
R18920 XThC.Tn[13].n25 XThC.Tn[13] 0.235138
R18921 XThC.Tn[13].n29 XThC.Tn[13] 0.235138
R18922 XThC.Tn[13].n33 XThC.Tn[13] 0.235138
R18923 XThC.Tn[13].n37 XThC.Tn[13] 0.235138
R18924 XThC.Tn[13].n41 XThC.Tn[13] 0.235138
R18925 XThC.Tn[13].n45 XThC.Tn[13] 0.235138
R18926 XThC.Tn[13].n49 XThC.Tn[13] 0.235138
R18927 XThC.Tn[13].n53 XThC.Tn[13] 0.235138
R18928 XThC.Tn[13].n57 XThC.Tn[13] 0.235138
R18929 XThC.Tn[13].n61 XThC.Tn[13] 0.235138
R18930 XThC.Tn[13].n65 XThC.Tn[13] 0.235138
R18931 XThC.Tn[13] XThC.Tn[13].n9 0.114505
R18932 XThC.Tn[13] XThC.Tn[13].n13 0.114505
R18933 XThC.Tn[13] XThC.Tn[13].n17 0.114505
R18934 XThC.Tn[13] XThC.Tn[13].n21 0.114505
R18935 XThC.Tn[13] XThC.Tn[13].n25 0.114505
R18936 XThC.Tn[13] XThC.Tn[13].n29 0.114505
R18937 XThC.Tn[13] XThC.Tn[13].n33 0.114505
R18938 XThC.Tn[13] XThC.Tn[13].n37 0.114505
R18939 XThC.Tn[13] XThC.Tn[13].n41 0.114505
R18940 XThC.Tn[13] XThC.Tn[13].n45 0.114505
R18941 XThC.Tn[13] XThC.Tn[13].n49 0.114505
R18942 XThC.Tn[13] XThC.Tn[13].n53 0.114505
R18943 XThC.Tn[13] XThC.Tn[13].n57 0.114505
R18944 XThC.Tn[13] XThC.Tn[13].n61 0.114505
R18945 XThC.Tn[13] XThC.Tn[13].n65 0.114505
R18946 XThC.Tn[13].n64 XThC.Tn[13].n63 0.0599512
R18947 XThC.Tn[13].n60 XThC.Tn[13].n59 0.0599512
R18948 XThC.Tn[13].n56 XThC.Tn[13].n55 0.0599512
R18949 XThC.Tn[13].n52 XThC.Tn[13].n51 0.0599512
R18950 XThC.Tn[13].n48 XThC.Tn[13].n47 0.0599512
R18951 XThC.Tn[13].n44 XThC.Tn[13].n43 0.0599512
R18952 XThC.Tn[13].n40 XThC.Tn[13].n39 0.0599512
R18953 XThC.Tn[13].n36 XThC.Tn[13].n35 0.0599512
R18954 XThC.Tn[13].n32 XThC.Tn[13].n31 0.0599512
R18955 XThC.Tn[13].n28 XThC.Tn[13].n27 0.0599512
R18956 XThC.Tn[13].n24 XThC.Tn[13].n23 0.0599512
R18957 XThC.Tn[13].n20 XThC.Tn[13].n19 0.0599512
R18958 XThC.Tn[13].n16 XThC.Tn[13].n15 0.0599512
R18959 XThC.Tn[13].n12 XThC.Tn[13].n11 0.0599512
R18960 XThC.Tn[13].n8 XThC.Tn[13].n7 0.0599512
R18961 XThC.Tn[13].n5 XThC.Tn[13].n4 0.0599512
R18962 XThC.Tn[13].n63 XThC.Tn[13] 0.0469286
R18963 XThC.Tn[13].n59 XThC.Tn[13] 0.0469286
R18964 XThC.Tn[13].n55 XThC.Tn[13] 0.0469286
R18965 XThC.Tn[13].n51 XThC.Tn[13] 0.0469286
R18966 XThC.Tn[13].n47 XThC.Tn[13] 0.0469286
R18967 XThC.Tn[13].n43 XThC.Tn[13] 0.0469286
R18968 XThC.Tn[13].n39 XThC.Tn[13] 0.0469286
R18969 XThC.Tn[13].n35 XThC.Tn[13] 0.0469286
R18970 XThC.Tn[13].n31 XThC.Tn[13] 0.0469286
R18971 XThC.Tn[13].n27 XThC.Tn[13] 0.0469286
R18972 XThC.Tn[13].n23 XThC.Tn[13] 0.0469286
R18973 XThC.Tn[13].n19 XThC.Tn[13] 0.0469286
R18974 XThC.Tn[13].n15 XThC.Tn[13] 0.0469286
R18975 XThC.Tn[13].n11 XThC.Tn[13] 0.0469286
R18976 XThC.Tn[13].n7 XThC.Tn[13] 0.0469286
R18977 XThC.Tn[13].n4 XThC.Tn[13] 0.0469286
R18978 XThC.Tn[13].n63 XThC.Tn[13] 0.0401341
R18979 XThC.Tn[13].n59 XThC.Tn[13] 0.0401341
R18980 XThC.Tn[13].n55 XThC.Tn[13] 0.0401341
R18981 XThC.Tn[13].n51 XThC.Tn[13] 0.0401341
R18982 XThC.Tn[13].n47 XThC.Tn[13] 0.0401341
R18983 XThC.Tn[13].n43 XThC.Tn[13] 0.0401341
R18984 XThC.Tn[13].n39 XThC.Tn[13] 0.0401341
R18985 XThC.Tn[13].n35 XThC.Tn[13] 0.0401341
R18986 XThC.Tn[13].n31 XThC.Tn[13] 0.0401341
R18987 XThC.Tn[13].n27 XThC.Tn[13] 0.0401341
R18988 XThC.Tn[13].n23 XThC.Tn[13] 0.0401341
R18989 XThC.Tn[13].n19 XThC.Tn[13] 0.0401341
R18990 XThC.Tn[13].n15 XThC.Tn[13] 0.0401341
R18991 XThC.Tn[13].n11 XThC.Tn[13] 0.0401341
R18992 XThC.Tn[13].n7 XThC.Tn[13] 0.0401341
R18993 XThC.Tn[13].n4 XThC.Tn[13] 0.0401341
R18994 XThC.Tn[0].n2 XThC.Tn[0].n1 332.332
R18995 XThC.Tn[0].n2 XThC.Tn[0].n0 296.493
R18996 XThC.Tn[0].n71 XThC.Tn[0].n69 161.365
R18997 XThC.Tn[0].n67 XThC.Tn[0].n65 161.365
R18998 XThC.Tn[0].n63 XThC.Tn[0].n61 161.365
R18999 XThC.Tn[0].n59 XThC.Tn[0].n57 161.365
R19000 XThC.Tn[0].n55 XThC.Tn[0].n53 161.365
R19001 XThC.Tn[0].n51 XThC.Tn[0].n49 161.365
R19002 XThC.Tn[0].n47 XThC.Tn[0].n45 161.365
R19003 XThC.Tn[0].n43 XThC.Tn[0].n41 161.365
R19004 XThC.Tn[0].n39 XThC.Tn[0].n37 161.365
R19005 XThC.Tn[0].n35 XThC.Tn[0].n33 161.365
R19006 XThC.Tn[0].n31 XThC.Tn[0].n29 161.365
R19007 XThC.Tn[0].n27 XThC.Tn[0].n25 161.365
R19008 XThC.Tn[0].n23 XThC.Tn[0].n21 161.365
R19009 XThC.Tn[0].n19 XThC.Tn[0].n17 161.365
R19010 XThC.Tn[0].n15 XThC.Tn[0].n13 161.365
R19011 XThC.Tn[0].n12 XThC.Tn[0].n10 161.365
R19012 XThC.Tn[0].n69 XThC.Tn[0].t29 161.202
R19013 XThC.Tn[0].n65 XThC.Tn[0].t19 161.202
R19014 XThC.Tn[0].n61 XThC.Tn[0].t38 161.202
R19015 XThC.Tn[0].n57 XThC.Tn[0].t36 161.202
R19016 XThC.Tn[0].n53 XThC.Tn[0].t27 161.202
R19017 XThC.Tn[0].n49 XThC.Tn[0].t16 161.202
R19018 XThC.Tn[0].n45 XThC.Tn[0].t15 161.202
R19019 XThC.Tn[0].n41 XThC.Tn[0].t26 161.202
R19020 XThC.Tn[0].n37 XThC.Tn[0].t25 161.202
R19021 XThC.Tn[0].n33 XThC.Tn[0].t17 161.202
R19022 XThC.Tn[0].n29 XThC.Tn[0].t34 161.202
R19023 XThC.Tn[0].n25 XThC.Tn[0].t32 161.202
R19024 XThC.Tn[0].n21 XThC.Tn[0].t13 161.202
R19025 XThC.Tn[0].n17 XThC.Tn[0].t12 161.202
R19026 XThC.Tn[0].n13 XThC.Tn[0].t41 161.202
R19027 XThC.Tn[0].n10 XThC.Tn[0].t22 161.202
R19028 XThC.Tn[0].n69 XThC.Tn[0].t24 145.137
R19029 XThC.Tn[0].n65 XThC.Tn[0].t14 145.137
R19030 XThC.Tn[0].n61 XThC.Tn[0].t33 145.137
R19031 XThC.Tn[0].n57 XThC.Tn[0].t31 145.137
R19032 XThC.Tn[0].n53 XThC.Tn[0].t23 145.137
R19033 XThC.Tn[0].n49 XThC.Tn[0].t42 145.137
R19034 XThC.Tn[0].n45 XThC.Tn[0].t40 145.137
R19035 XThC.Tn[0].n41 XThC.Tn[0].t21 145.137
R19036 XThC.Tn[0].n37 XThC.Tn[0].t20 145.137
R19037 XThC.Tn[0].n33 XThC.Tn[0].t43 145.137
R19038 XThC.Tn[0].n29 XThC.Tn[0].t30 145.137
R19039 XThC.Tn[0].n25 XThC.Tn[0].t28 145.137
R19040 XThC.Tn[0].n21 XThC.Tn[0].t39 145.137
R19041 XThC.Tn[0].n17 XThC.Tn[0].t37 145.137
R19042 XThC.Tn[0].n13 XThC.Tn[0].t35 145.137
R19043 XThC.Tn[0].n10 XThC.Tn[0].t18 145.137
R19044 XThC.Tn[0].n7 XThC.Tn[0].n6 135.248
R19045 XThC.Tn[0].n9 XThC.Tn[0].n3 98.982
R19046 XThC.Tn[0].n8 XThC.Tn[0].n4 98.982
R19047 XThC.Tn[0].n7 XThC.Tn[0].n5 98.982
R19048 XThC.Tn[0].n9 XThC.Tn[0].n8 36.2672
R19049 XThC.Tn[0].n8 XThC.Tn[0].n7 36.2672
R19050 XThC.Tn[0].n74 XThC.Tn[0].n9 32.6405
R19051 XThC.Tn[0].n1 XThC.Tn[0].t10 26.5955
R19052 XThC.Tn[0].n1 XThC.Tn[0].t9 26.5955
R19053 XThC.Tn[0].n0 XThC.Tn[0].t8 26.5955
R19054 XThC.Tn[0].n0 XThC.Tn[0].t7 26.5955
R19055 XThC.Tn[0].n3 XThC.Tn[0].t4 24.9236
R19056 XThC.Tn[0].n3 XThC.Tn[0].t3 24.9236
R19057 XThC.Tn[0].n4 XThC.Tn[0].t6 24.9236
R19058 XThC.Tn[0].n4 XThC.Tn[0].t5 24.9236
R19059 XThC.Tn[0].n5 XThC.Tn[0].t1 24.9236
R19060 XThC.Tn[0].n5 XThC.Tn[0].t2 24.9236
R19061 XThC.Tn[0].n6 XThC.Tn[0].t11 24.9236
R19062 XThC.Tn[0].n6 XThC.Tn[0].t0 24.9236
R19063 XThC.Tn[0].n75 XThC.Tn[0].n2 18.5605
R19064 XThC.Tn[0].n73 XThC.Tn[0] 16.199
R19065 XThC.Tn[0].n75 XThC.Tn[0].n74 11.5205
R19066 XThC.Tn[0] XThC.Tn[0].n12 8.0245
R19067 XThC.Tn[0].n72 XThC.Tn[0].n71 7.9105
R19068 XThC.Tn[0].n68 XThC.Tn[0].n67 7.9105
R19069 XThC.Tn[0].n64 XThC.Tn[0].n63 7.9105
R19070 XThC.Tn[0].n60 XThC.Tn[0].n59 7.9105
R19071 XThC.Tn[0].n56 XThC.Tn[0].n55 7.9105
R19072 XThC.Tn[0].n52 XThC.Tn[0].n51 7.9105
R19073 XThC.Tn[0].n48 XThC.Tn[0].n47 7.9105
R19074 XThC.Tn[0].n44 XThC.Tn[0].n43 7.9105
R19075 XThC.Tn[0].n40 XThC.Tn[0].n39 7.9105
R19076 XThC.Tn[0].n36 XThC.Tn[0].n35 7.9105
R19077 XThC.Tn[0].n32 XThC.Tn[0].n31 7.9105
R19078 XThC.Tn[0].n28 XThC.Tn[0].n27 7.9105
R19079 XThC.Tn[0].n24 XThC.Tn[0].n23 7.9105
R19080 XThC.Tn[0].n20 XThC.Tn[0].n19 7.9105
R19081 XThC.Tn[0].n16 XThC.Tn[0].n15 7.9105
R19082 XThC.Tn[0].n74 XThC.Tn[0].n73 4.6005
R19083 XThC.Tn[0].n73 XThC.Tn[0] 1.84237
R19084 XThC.Tn[0] XThC.Tn[0].n75 0.6405
R19085 XThC.Tn[0].n16 XThC.Tn[0] 0.235138
R19086 XThC.Tn[0].n20 XThC.Tn[0] 0.235138
R19087 XThC.Tn[0].n24 XThC.Tn[0] 0.235138
R19088 XThC.Tn[0].n28 XThC.Tn[0] 0.235138
R19089 XThC.Tn[0].n32 XThC.Tn[0] 0.235138
R19090 XThC.Tn[0].n36 XThC.Tn[0] 0.235138
R19091 XThC.Tn[0].n40 XThC.Tn[0] 0.235138
R19092 XThC.Tn[0].n44 XThC.Tn[0] 0.235138
R19093 XThC.Tn[0].n48 XThC.Tn[0] 0.235138
R19094 XThC.Tn[0].n52 XThC.Tn[0] 0.235138
R19095 XThC.Tn[0].n56 XThC.Tn[0] 0.235138
R19096 XThC.Tn[0].n60 XThC.Tn[0] 0.235138
R19097 XThC.Tn[0].n64 XThC.Tn[0] 0.235138
R19098 XThC.Tn[0].n68 XThC.Tn[0] 0.235138
R19099 XThC.Tn[0].n72 XThC.Tn[0] 0.235138
R19100 XThC.Tn[0] XThC.Tn[0].n16 0.114505
R19101 XThC.Tn[0] XThC.Tn[0].n20 0.114505
R19102 XThC.Tn[0] XThC.Tn[0].n24 0.114505
R19103 XThC.Tn[0] XThC.Tn[0].n28 0.114505
R19104 XThC.Tn[0] XThC.Tn[0].n32 0.114505
R19105 XThC.Tn[0] XThC.Tn[0].n36 0.114505
R19106 XThC.Tn[0] XThC.Tn[0].n40 0.114505
R19107 XThC.Tn[0] XThC.Tn[0].n44 0.114505
R19108 XThC.Tn[0] XThC.Tn[0].n48 0.114505
R19109 XThC.Tn[0] XThC.Tn[0].n52 0.114505
R19110 XThC.Tn[0] XThC.Tn[0].n56 0.114505
R19111 XThC.Tn[0] XThC.Tn[0].n60 0.114505
R19112 XThC.Tn[0] XThC.Tn[0].n64 0.114505
R19113 XThC.Tn[0] XThC.Tn[0].n68 0.114505
R19114 XThC.Tn[0] XThC.Tn[0].n72 0.114505
R19115 XThC.Tn[0].n71 XThC.Tn[0].n70 0.0599512
R19116 XThC.Tn[0].n67 XThC.Tn[0].n66 0.0599512
R19117 XThC.Tn[0].n63 XThC.Tn[0].n62 0.0599512
R19118 XThC.Tn[0].n59 XThC.Tn[0].n58 0.0599512
R19119 XThC.Tn[0].n55 XThC.Tn[0].n54 0.0599512
R19120 XThC.Tn[0].n51 XThC.Tn[0].n50 0.0599512
R19121 XThC.Tn[0].n47 XThC.Tn[0].n46 0.0599512
R19122 XThC.Tn[0].n43 XThC.Tn[0].n42 0.0599512
R19123 XThC.Tn[0].n39 XThC.Tn[0].n38 0.0599512
R19124 XThC.Tn[0].n35 XThC.Tn[0].n34 0.0599512
R19125 XThC.Tn[0].n31 XThC.Tn[0].n30 0.0599512
R19126 XThC.Tn[0].n27 XThC.Tn[0].n26 0.0599512
R19127 XThC.Tn[0].n23 XThC.Tn[0].n22 0.0599512
R19128 XThC.Tn[0].n19 XThC.Tn[0].n18 0.0599512
R19129 XThC.Tn[0].n15 XThC.Tn[0].n14 0.0599512
R19130 XThC.Tn[0].n12 XThC.Tn[0].n11 0.0599512
R19131 XThC.Tn[0].n70 XThC.Tn[0] 0.0469286
R19132 XThC.Tn[0].n66 XThC.Tn[0] 0.0469286
R19133 XThC.Tn[0].n62 XThC.Tn[0] 0.0469286
R19134 XThC.Tn[0].n58 XThC.Tn[0] 0.0469286
R19135 XThC.Tn[0].n54 XThC.Tn[0] 0.0469286
R19136 XThC.Tn[0].n50 XThC.Tn[0] 0.0469286
R19137 XThC.Tn[0].n46 XThC.Tn[0] 0.0469286
R19138 XThC.Tn[0].n42 XThC.Tn[0] 0.0469286
R19139 XThC.Tn[0].n38 XThC.Tn[0] 0.0469286
R19140 XThC.Tn[0].n34 XThC.Tn[0] 0.0469286
R19141 XThC.Tn[0].n30 XThC.Tn[0] 0.0469286
R19142 XThC.Tn[0].n26 XThC.Tn[0] 0.0469286
R19143 XThC.Tn[0].n22 XThC.Tn[0] 0.0469286
R19144 XThC.Tn[0].n18 XThC.Tn[0] 0.0469286
R19145 XThC.Tn[0].n14 XThC.Tn[0] 0.0469286
R19146 XThC.Tn[0].n11 XThC.Tn[0] 0.0469286
R19147 XThC.Tn[0].n70 XThC.Tn[0] 0.0401341
R19148 XThC.Tn[0].n66 XThC.Tn[0] 0.0401341
R19149 XThC.Tn[0].n62 XThC.Tn[0] 0.0401341
R19150 XThC.Tn[0].n58 XThC.Tn[0] 0.0401341
R19151 XThC.Tn[0].n54 XThC.Tn[0] 0.0401341
R19152 XThC.Tn[0].n50 XThC.Tn[0] 0.0401341
R19153 XThC.Tn[0].n46 XThC.Tn[0] 0.0401341
R19154 XThC.Tn[0].n42 XThC.Tn[0] 0.0401341
R19155 XThC.Tn[0].n38 XThC.Tn[0] 0.0401341
R19156 XThC.Tn[0].n34 XThC.Tn[0] 0.0401341
R19157 XThC.Tn[0].n30 XThC.Tn[0] 0.0401341
R19158 XThC.Tn[0].n26 XThC.Tn[0] 0.0401341
R19159 XThC.Tn[0].n22 XThC.Tn[0] 0.0401341
R19160 XThC.Tn[0].n18 XThC.Tn[0] 0.0401341
R19161 XThC.Tn[0].n14 XThC.Tn[0] 0.0401341
R19162 XThC.Tn[0].n11 XThC.Tn[0] 0.0401341
R19163 XThC.XTB4.Y.n21 XThC.XTB4.Y.t0 235.56
R19164 XThC.XTB4.Y.n3 XThC.XTB4.Y.t3 212.081
R19165 XThC.XTB4.Y.n2 XThC.XTB4.Y.t2 212.081
R19166 XThC.XTB4.Y.n8 XThC.XTB4.Y.t17 212.081
R19167 XThC.XTB4.Y.n0 XThC.XTB4.Y.t13 212.081
R19168 XThC.XTB4.Y.n12 XThC.XTB4.Y.t8 212.081
R19169 XThC.XTB4.Y.n13 XThC.XTB4.Y.t12 212.081
R19170 XThC.XTB4.Y.n15 XThC.XTB4.Y.t6 212.081
R19171 XThC.XTB4.Y.n11 XThC.XTB4.Y.t16 212.081
R19172 XThC.XTB4.Y.n5 XThC.XTB4.Y.n4 173.761
R19173 XThC.XTB4.Y.n14 XThC.XTB4.Y 158.656
R19174 XThC.XTB4.Y.n7 XThC.XTB4.Y.n6 152
R19175 XThC.XTB4.Y.n5 XThC.XTB4.Y.n1 152
R19176 XThC.XTB4.Y.n10 XThC.XTB4.Y.n9 152
R19177 XThC.XTB4.Y.n17 XThC.XTB4.Y.n16 152
R19178 XThC.XTB4.Y.n3 XThC.XTB4.Y.t14 139.78
R19179 XThC.XTB4.Y.n2 XThC.XTB4.Y.t10 139.78
R19180 XThC.XTB4.Y.n8 XThC.XTB4.Y.t7 139.78
R19181 XThC.XTB4.Y.n0 XThC.XTB4.Y.t4 139.78
R19182 XThC.XTB4.Y.n12 XThC.XTB4.Y.t11 139.78
R19183 XThC.XTB4.Y.n13 XThC.XTB4.Y.t15 139.78
R19184 XThC.XTB4.Y.n15 XThC.XTB4.Y.t9 139.78
R19185 XThC.XTB4.Y.n11 XThC.XTB4.Y.t5 139.78
R19186 XThC.XTB4.Y.n20 XThC.XTB4.Y.t1 133.386
R19187 XThC.XTB4.Y.n19 XThC.XTB4.Y.n10 72.9296
R19188 XThC.XTB4.Y.n13 XThC.XTB4.Y.n12 61.346
R19189 XThC.XTB4.Y.n7 XThC.XTB4.Y.n1 49.6611
R19190 XThC.XTB4.Y.n9 XThC.XTB4.Y.n8 45.2793
R19191 XThC.XTB4.Y.n4 XThC.XTB4.Y.n2 42.3581
R19192 XThC.XTB4.Y.n19 XThC.XTB4.Y.n18 38.1854
R19193 XThC.XTB4.Y.n16 XThC.XTB4.Y.n11 30.6732
R19194 XThC.XTB4.Y.n16 XThC.XTB4.Y.n15 30.6732
R19195 XThC.XTB4.Y.n15 XThC.XTB4.Y.n14 30.6732
R19196 XThC.XTB4.Y.n14 XThC.XTB4.Y.n13 30.6732
R19197 XThC.XTB4.Y.n6 XThC.XTB4.Y.n5 21.7605
R19198 XThC.XTB4.Y XThC.XTB4.Y.n20 19.5051
R19199 XThC.XTB4.Y.n4 XThC.XTB4.Y.n3 18.9884
R19200 XThC.XTB4.Y.n9 XThC.XTB4.Y.n0 16.0672
R19201 XThC.XTB4.Y.n17 XThC.XTB4.Y 14.7905
R19202 XThC.XTB4.Y.n20 XThC.XTB4.Y.n19 11.994
R19203 XThC.XTB4.Y.n10 XThC.XTB4.Y 11.5205
R19204 XThC.XTB4.Y.n6 XThC.XTB4.Y 10.2405
R19205 XThC.XTB4.Y.n2 XThC.XTB4.Y.n1 7.30353
R19206 XThC.XTB4.Y.n18 XThC.XTB4.Y.n17 7.24578
R19207 XThC.XTB4.Y.n8 XThC.XTB4.Y.n7 4.38232
R19208 XThC.XTB4.Y.n21 XThC.XTB4.Y 2.22659
R19209 XThC.XTB4.Y XThC.XTB4.Y.n21 1.55202
R19210 XThC.XTB4.Y.n18 XThC.XTB4.Y 0.966538
R19211 XThR.Tn[3].n2 XThR.Tn[3].n1 332.332
R19212 XThR.Tn[3].n2 XThR.Tn[3].n0 296.493
R19213 XThR.Tn[3] XThR.Tn[3].n82 161.363
R19214 XThR.Tn[3] XThR.Tn[3].n77 161.363
R19215 XThR.Tn[3] XThR.Tn[3].n72 161.363
R19216 XThR.Tn[3] XThR.Tn[3].n67 161.363
R19217 XThR.Tn[3] XThR.Tn[3].n62 161.363
R19218 XThR.Tn[3] XThR.Tn[3].n57 161.363
R19219 XThR.Tn[3] XThR.Tn[3].n52 161.363
R19220 XThR.Tn[3] XThR.Tn[3].n47 161.363
R19221 XThR.Tn[3] XThR.Tn[3].n42 161.363
R19222 XThR.Tn[3] XThR.Tn[3].n37 161.363
R19223 XThR.Tn[3] XThR.Tn[3].n32 161.363
R19224 XThR.Tn[3] XThR.Tn[3].n27 161.363
R19225 XThR.Tn[3] XThR.Tn[3].n22 161.363
R19226 XThR.Tn[3] XThR.Tn[3].n17 161.363
R19227 XThR.Tn[3] XThR.Tn[3].n12 161.363
R19228 XThR.Tn[3] XThR.Tn[3].n10 161.363
R19229 XThR.Tn[3].n84 XThR.Tn[3].n83 161.3
R19230 XThR.Tn[3].n79 XThR.Tn[3].n78 161.3
R19231 XThR.Tn[3].n74 XThR.Tn[3].n73 161.3
R19232 XThR.Tn[3].n69 XThR.Tn[3].n68 161.3
R19233 XThR.Tn[3].n64 XThR.Tn[3].n63 161.3
R19234 XThR.Tn[3].n59 XThR.Tn[3].n58 161.3
R19235 XThR.Tn[3].n54 XThR.Tn[3].n53 161.3
R19236 XThR.Tn[3].n49 XThR.Tn[3].n48 161.3
R19237 XThR.Tn[3].n44 XThR.Tn[3].n43 161.3
R19238 XThR.Tn[3].n39 XThR.Tn[3].n38 161.3
R19239 XThR.Tn[3].n34 XThR.Tn[3].n33 161.3
R19240 XThR.Tn[3].n29 XThR.Tn[3].n28 161.3
R19241 XThR.Tn[3].n24 XThR.Tn[3].n23 161.3
R19242 XThR.Tn[3].n19 XThR.Tn[3].n18 161.3
R19243 XThR.Tn[3].n14 XThR.Tn[3].n13 161.3
R19244 XThR.Tn[3].n82 XThR.Tn[3].t46 161.106
R19245 XThR.Tn[3].n77 XThR.Tn[3].t53 161.106
R19246 XThR.Tn[3].n72 XThR.Tn[3].t34 161.106
R19247 XThR.Tn[3].n67 XThR.Tn[3].t17 161.106
R19248 XThR.Tn[3].n62 XThR.Tn[3].t44 161.106
R19249 XThR.Tn[3].n57 XThR.Tn[3].t69 161.106
R19250 XThR.Tn[3].n52 XThR.Tn[3].t51 161.106
R19251 XThR.Tn[3].n47 XThR.Tn[3].t31 161.106
R19252 XThR.Tn[3].n42 XThR.Tn[3].t14 161.106
R19253 XThR.Tn[3].n37 XThR.Tn[3].t20 161.106
R19254 XThR.Tn[3].n32 XThR.Tn[3].t68 161.106
R19255 XThR.Tn[3].n27 XThR.Tn[3].t33 161.106
R19256 XThR.Tn[3].n22 XThR.Tn[3].t67 161.106
R19257 XThR.Tn[3].n17 XThR.Tn[3].t49 161.106
R19258 XThR.Tn[3].n12 XThR.Tn[3].t70 161.106
R19259 XThR.Tn[3].n10 XThR.Tn[3].t57 161.106
R19260 XThR.Tn[3].n83 XThR.Tn[3].t27 159.978
R19261 XThR.Tn[3].n78 XThR.Tn[3].t32 159.978
R19262 XThR.Tn[3].n73 XThR.Tn[3].t15 159.978
R19263 XThR.Tn[3].n68 XThR.Tn[3].t63 159.978
R19264 XThR.Tn[3].n63 XThR.Tn[3].t25 159.978
R19265 XThR.Tn[3].n58 XThR.Tn[3].t50 159.978
R19266 XThR.Tn[3].n53 XThR.Tn[3].t30 159.978
R19267 XThR.Tn[3].n48 XThR.Tn[3].t73 159.978
R19268 XThR.Tn[3].n43 XThR.Tn[3].t61 159.978
R19269 XThR.Tn[3].n38 XThR.Tn[3].t66 159.978
R19270 XThR.Tn[3].n33 XThR.Tn[3].t48 159.978
R19271 XThR.Tn[3].n28 XThR.Tn[3].t13 159.978
R19272 XThR.Tn[3].n23 XThR.Tn[3].t47 159.978
R19273 XThR.Tn[3].n18 XThR.Tn[3].t29 159.978
R19274 XThR.Tn[3].n13 XThR.Tn[3].t55 159.978
R19275 XThR.Tn[3].n82 XThR.Tn[3].t36 145.038
R19276 XThR.Tn[3].n77 XThR.Tn[3].t60 145.038
R19277 XThR.Tn[3].n72 XThR.Tn[3].t40 145.038
R19278 XThR.Tn[3].n67 XThR.Tn[3].t21 145.038
R19279 XThR.Tn[3].n62 XThR.Tn[3].t54 145.038
R19280 XThR.Tn[3].n57 XThR.Tn[3].t35 145.038
R19281 XThR.Tn[3].n52 XThR.Tn[3].t41 145.038
R19282 XThR.Tn[3].n47 XThR.Tn[3].t22 145.038
R19283 XThR.Tn[3].n42 XThR.Tn[3].t19 145.038
R19284 XThR.Tn[3].n37 XThR.Tn[3].t52 145.038
R19285 XThR.Tn[3].n32 XThR.Tn[3].t72 145.038
R19286 XThR.Tn[3].n27 XThR.Tn[3].t39 145.038
R19287 XThR.Tn[3].n22 XThR.Tn[3].t71 145.038
R19288 XThR.Tn[3].n17 XThR.Tn[3].t59 145.038
R19289 XThR.Tn[3].n12 XThR.Tn[3].t18 145.038
R19290 XThR.Tn[3].n10 XThR.Tn[3].t64 145.038
R19291 XThR.Tn[3].n83 XThR.Tn[3].t38 143.911
R19292 XThR.Tn[3].n78 XThR.Tn[3].t65 143.911
R19293 XThR.Tn[3].n73 XThR.Tn[3].t43 143.911
R19294 XThR.Tn[3].n68 XThR.Tn[3].t26 143.911
R19295 XThR.Tn[3].n63 XThR.Tn[3].t58 143.911
R19296 XThR.Tn[3].n58 XThR.Tn[3].t37 143.911
R19297 XThR.Tn[3].n53 XThR.Tn[3].t45 143.911
R19298 XThR.Tn[3].n48 XThR.Tn[3].t28 143.911
R19299 XThR.Tn[3].n43 XThR.Tn[3].t23 143.911
R19300 XThR.Tn[3].n38 XThR.Tn[3].t56 143.911
R19301 XThR.Tn[3].n33 XThR.Tn[3].t16 143.911
R19302 XThR.Tn[3].n28 XThR.Tn[3].t42 143.911
R19303 XThR.Tn[3].n23 XThR.Tn[3].t12 143.911
R19304 XThR.Tn[3].n18 XThR.Tn[3].t62 143.911
R19305 XThR.Tn[3].n13 XThR.Tn[3].t24 143.911
R19306 XThR.Tn[3].n7 XThR.Tn[3].n6 135.249
R19307 XThR.Tn[3].n9 XThR.Tn[3].n3 98.981
R19308 XThR.Tn[3].n8 XThR.Tn[3].n4 98.981
R19309 XThR.Tn[3].n7 XThR.Tn[3].n5 98.981
R19310 XThR.Tn[3].n9 XThR.Tn[3].n8 36.2672
R19311 XThR.Tn[3].n8 XThR.Tn[3].n7 36.2672
R19312 XThR.Tn[3].n88 XThR.Tn[3].n9 32.6405
R19313 XThR.Tn[3].n1 XThR.Tn[3].t1 26.5955
R19314 XThR.Tn[3].n1 XThR.Tn[3].t4 26.5955
R19315 XThR.Tn[3].n0 XThR.Tn[3].t2 26.5955
R19316 XThR.Tn[3].n0 XThR.Tn[3].t3 26.5955
R19317 XThR.Tn[3].n3 XThR.Tn[3].t8 24.9236
R19318 XThR.Tn[3].n3 XThR.Tn[3].t5 24.9236
R19319 XThR.Tn[3].n4 XThR.Tn[3].t7 24.9236
R19320 XThR.Tn[3].n4 XThR.Tn[3].t6 24.9236
R19321 XThR.Tn[3].n5 XThR.Tn[3].t9 24.9236
R19322 XThR.Tn[3].n5 XThR.Tn[3].t10 24.9236
R19323 XThR.Tn[3].n6 XThR.Tn[3].t0 24.9236
R19324 XThR.Tn[3].n6 XThR.Tn[3].t11 24.9236
R19325 XThR.Tn[3].n89 XThR.Tn[3].n2 18.5605
R19326 XThR.Tn[3].n89 XThR.Tn[3].n88 11.5205
R19327 XThR.Tn[3].n88 XThR.Tn[3] 6.21508
R19328 XThR.Tn[3] XThR.Tn[3].n11 5.34038
R19329 XThR.Tn[3].n16 XThR.Tn[3].n15 4.5005
R19330 XThR.Tn[3].n21 XThR.Tn[3].n20 4.5005
R19331 XThR.Tn[3].n26 XThR.Tn[3].n25 4.5005
R19332 XThR.Tn[3].n31 XThR.Tn[3].n30 4.5005
R19333 XThR.Tn[3].n36 XThR.Tn[3].n35 4.5005
R19334 XThR.Tn[3].n41 XThR.Tn[3].n40 4.5005
R19335 XThR.Tn[3].n46 XThR.Tn[3].n45 4.5005
R19336 XThR.Tn[3].n51 XThR.Tn[3].n50 4.5005
R19337 XThR.Tn[3].n56 XThR.Tn[3].n55 4.5005
R19338 XThR.Tn[3].n61 XThR.Tn[3].n60 4.5005
R19339 XThR.Tn[3].n66 XThR.Tn[3].n65 4.5005
R19340 XThR.Tn[3].n71 XThR.Tn[3].n70 4.5005
R19341 XThR.Tn[3].n76 XThR.Tn[3].n75 4.5005
R19342 XThR.Tn[3].n81 XThR.Tn[3].n80 4.5005
R19343 XThR.Tn[3].n86 XThR.Tn[3].n85 4.5005
R19344 XThR.Tn[3].n87 XThR.Tn[3] 3.70586
R19345 XThR.Tn[3].n16 XThR.Tn[3] 2.52282
R19346 XThR.Tn[3].n21 XThR.Tn[3] 2.52282
R19347 XThR.Tn[3].n26 XThR.Tn[3] 2.52282
R19348 XThR.Tn[3].n31 XThR.Tn[3] 2.52282
R19349 XThR.Tn[3].n36 XThR.Tn[3] 2.52282
R19350 XThR.Tn[3].n41 XThR.Tn[3] 2.52282
R19351 XThR.Tn[3].n46 XThR.Tn[3] 2.52282
R19352 XThR.Tn[3].n51 XThR.Tn[3] 2.52282
R19353 XThR.Tn[3].n56 XThR.Tn[3] 2.52282
R19354 XThR.Tn[3].n61 XThR.Tn[3] 2.52282
R19355 XThR.Tn[3].n66 XThR.Tn[3] 2.52282
R19356 XThR.Tn[3].n71 XThR.Tn[3] 2.52282
R19357 XThR.Tn[3].n76 XThR.Tn[3] 2.52282
R19358 XThR.Tn[3].n81 XThR.Tn[3] 2.52282
R19359 XThR.Tn[3].n86 XThR.Tn[3] 2.52282
R19360 XThR.Tn[3].n84 XThR.Tn[3] 1.08677
R19361 XThR.Tn[3].n79 XThR.Tn[3] 1.08677
R19362 XThR.Tn[3].n74 XThR.Tn[3] 1.08677
R19363 XThR.Tn[3].n69 XThR.Tn[3] 1.08677
R19364 XThR.Tn[3].n64 XThR.Tn[3] 1.08677
R19365 XThR.Tn[3].n59 XThR.Tn[3] 1.08677
R19366 XThR.Tn[3].n54 XThR.Tn[3] 1.08677
R19367 XThR.Tn[3].n49 XThR.Tn[3] 1.08677
R19368 XThR.Tn[3].n44 XThR.Tn[3] 1.08677
R19369 XThR.Tn[3].n39 XThR.Tn[3] 1.08677
R19370 XThR.Tn[3].n34 XThR.Tn[3] 1.08677
R19371 XThR.Tn[3].n29 XThR.Tn[3] 1.08677
R19372 XThR.Tn[3].n24 XThR.Tn[3] 1.08677
R19373 XThR.Tn[3].n19 XThR.Tn[3] 1.08677
R19374 XThR.Tn[3].n14 XThR.Tn[3] 1.08677
R19375 XThR.Tn[3] XThR.Tn[3].n16 0.839786
R19376 XThR.Tn[3] XThR.Tn[3].n21 0.839786
R19377 XThR.Tn[3] XThR.Tn[3].n26 0.839786
R19378 XThR.Tn[3] XThR.Tn[3].n31 0.839786
R19379 XThR.Tn[3] XThR.Tn[3].n36 0.839786
R19380 XThR.Tn[3] XThR.Tn[3].n41 0.839786
R19381 XThR.Tn[3] XThR.Tn[3].n46 0.839786
R19382 XThR.Tn[3] XThR.Tn[3].n51 0.839786
R19383 XThR.Tn[3] XThR.Tn[3].n56 0.839786
R19384 XThR.Tn[3] XThR.Tn[3].n61 0.839786
R19385 XThR.Tn[3] XThR.Tn[3].n66 0.839786
R19386 XThR.Tn[3] XThR.Tn[3].n71 0.839786
R19387 XThR.Tn[3] XThR.Tn[3].n76 0.839786
R19388 XThR.Tn[3] XThR.Tn[3].n81 0.839786
R19389 XThR.Tn[3] XThR.Tn[3].n86 0.839786
R19390 XThR.Tn[3] XThR.Tn[3].n89 0.6405
R19391 XThR.Tn[3].n11 XThR.Tn[3] 0.499542
R19392 XThR.Tn[3].n85 XThR.Tn[3] 0.063
R19393 XThR.Tn[3].n80 XThR.Tn[3] 0.063
R19394 XThR.Tn[3].n75 XThR.Tn[3] 0.063
R19395 XThR.Tn[3].n70 XThR.Tn[3] 0.063
R19396 XThR.Tn[3].n65 XThR.Tn[3] 0.063
R19397 XThR.Tn[3].n60 XThR.Tn[3] 0.063
R19398 XThR.Tn[3].n55 XThR.Tn[3] 0.063
R19399 XThR.Tn[3].n50 XThR.Tn[3] 0.063
R19400 XThR.Tn[3].n45 XThR.Tn[3] 0.063
R19401 XThR.Tn[3].n40 XThR.Tn[3] 0.063
R19402 XThR.Tn[3].n35 XThR.Tn[3] 0.063
R19403 XThR.Tn[3].n30 XThR.Tn[3] 0.063
R19404 XThR.Tn[3].n25 XThR.Tn[3] 0.063
R19405 XThR.Tn[3].n20 XThR.Tn[3] 0.063
R19406 XThR.Tn[3].n15 XThR.Tn[3] 0.063
R19407 XThR.Tn[3].n87 XThR.Tn[3] 0.0540714
R19408 XThR.Tn[3] XThR.Tn[3].n87 0.038
R19409 XThR.Tn[3].n11 XThR.Tn[3] 0.0143889
R19410 XThR.Tn[3].n85 XThR.Tn[3].n84 0.00771154
R19411 XThR.Tn[3].n80 XThR.Tn[3].n79 0.00771154
R19412 XThR.Tn[3].n75 XThR.Tn[3].n74 0.00771154
R19413 XThR.Tn[3].n70 XThR.Tn[3].n69 0.00771154
R19414 XThR.Tn[3].n65 XThR.Tn[3].n64 0.00771154
R19415 XThR.Tn[3].n60 XThR.Tn[3].n59 0.00771154
R19416 XThR.Tn[3].n55 XThR.Tn[3].n54 0.00771154
R19417 XThR.Tn[3].n50 XThR.Tn[3].n49 0.00771154
R19418 XThR.Tn[3].n45 XThR.Tn[3].n44 0.00771154
R19419 XThR.Tn[3].n40 XThR.Tn[3].n39 0.00771154
R19420 XThR.Tn[3].n35 XThR.Tn[3].n34 0.00771154
R19421 XThR.Tn[3].n30 XThR.Tn[3].n29 0.00771154
R19422 XThR.Tn[3].n25 XThR.Tn[3].n24 0.00771154
R19423 XThR.Tn[3].n20 XThR.Tn[3].n19 0.00771154
R19424 XThR.Tn[3].n15 XThR.Tn[3].n14 0.00771154
R19425 XThR.Tn[5].n2 XThR.Tn[5].n1 332.332
R19426 XThR.Tn[5].n2 XThR.Tn[5].n0 296.493
R19427 XThR.Tn[5] XThR.Tn[5].n82 161.363
R19428 XThR.Tn[5] XThR.Tn[5].n77 161.363
R19429 XThR.Tn[5] XThR.Tn[5].n72 161.363
R19430 XThR.Tn[5] XThR.Tn[5].n67 161.363
R19431 XThR.Tn[5] XThR.Tn[5].n62 161.363
R19432 XThR.Tn[5] XThR.Tn[5].n57 161.363
R19433 XThR.Tn[5] XThR.Tn[5].n52 161.363
R19434 XThR.Tn[5] XThR.Tn[5].n47 161.363
R19435 XThR.Tn[5] XThR.Tn[5].n42 161.363
R19436 XThR.Tn[5] XThR.Tn[5].n37 161.363
R19437 XThR.Tn[5] XThR.Tn[5].n32 161.363
R19438 XThR.Tn[5] XThR.Tn[5].n27 161.363
R19439 XThR.Tn[5] XThR.Tn[5].n22 161.363
R19440 XThR.Tn[5] XThR.Tn[5].n17 161.363
R19441 XThR.Tn[5] XThR.Tn[5].n12 161.363
R19442 XThR.Tn[5] XThR.Tn[5].n10 161.363
R19443 XThR.Tn[5].n84 XThR.Tn[5].n83 161.3
R19444 XThR.Tn[5].n79 XThR.Tn[5].n78 161.3
R19445 XThR.Tn[5].n74 XThR.Tn[5].n73 161.3
R19446 XThR.Tn[5].n69 XThR.Tn[5].n68 161.3
R19447 XThR.Tn[5].n64 XThR.Tn[5].n63 161.3
R19448 XThR.Tn[5].n59 XThR.Tn[5].n58 161.3
R19449 XThR.Tn[5].n54 XThR.Tn[5].n53 161.3
R19450 XThR.Tn[5].n49 XThR.Tn[5].n48 161.3
R19451 XThR.Tn[5].n44 XThR.Tn[5].n43 161.3
R19452 XThR.Tn[5].n39 XThR.Tn[5].n38 161.3
R19453 XThR.Tn[5].n34 XThR.Tn[5].n33 161.3
R19454 XThR.Tn[5].n29 XThR.Tn[5].n28 161.3
R19455 XThR.Tn[5].n24 XThR.Tn[5].n23 161.3
R19456 XThR.Tn[5].n19 XThR.Tn[5].n18 161.3
R19457 XThR.Tn[5].n14 XThR.Tn[5].n13 161.3
R19458 XThR.Tn[5].n82 XThR.Tn[5].t62 161.106
R19459 XThR.Tn[5].n77 XThR.Tn[5].t70 161.106
R19460 XThR.Tn[5].n72 XThR.Tn[5].t52 161.106
R19461 XThR.Tn[5].n67 XThR.Tn[5].t35 161.106
R19462 XThR.Tn[5].n62 XThR.Tn[5].t60 161.106
R19463 XThR.Tn[5].n57 XThR.Tn[5].t24 161.106
R19464 XThR.Tn[5].n52 XThR.Tn[5].t68 161.106
R19465 XThR.Tn[5].n47 XThR.Tn[5].t49 161.106
R19466 XThR.Tn[5].n42 XThR.Tn[5].t32 161.106
R19467 XThR.Tn[5].n37 XThR.Tn[5].t40 161.106
R19468 XThR.Tn[5].n32 XThR.Tn[5].t22 161.106
R19469 XThR.Tn[5].n27 XThR.Tn[5].t51 161.106
R19470 XThR.Tn[5].n22 XThR.Tn[5].t21 161.106
R19471 XThR.Tn[5].n17 XThR.Tn[5].t66 161.106
R19472 XThR.Tn[5].n12 XThR.Tn[5].t26 161.106
R19473 XThR.Tn[5].n10 XThR.Tn[5].t72 161.106
R19474 XThR.Tn[5].n83 XThR.Tn[5].t59 159.978
R19475 XThR.Tn[5].n78 XThR.Tn[5].t64 159.978
R19476 XThR.Tn[5].n73 XThR.Tn[5].t47 159.978
R19477 XThR.Tn[5].n68 XThR.Tn[5].t31 159.978
R19478 XThR.Tn[5].n63 XThR.Tn[5].t57 159.978
R19479 XThR.Tn[5].n58 XThR.Tn[5].t20 159.978
R19480 XThR.Tn[5].n53 XThR.Tn[5].t63 159.978
R19481 XThR.Tn[5].n48 XThR.Tn[5].t45 159.978
R19482 XThR.Tn[5].n43 XThR.Tn[5].t29 159.978
R19483 XThR.Tn[5].n38 XThR.Tn[5].t37 159.978
R19484 XThR.Tn[5].n33 XThR.Tn[5].t19 159.978
R19485 XThR.Tn[5].n28 XThR.Tn[5].t46 159.978
R19486 XThR.Tn[5].n23 XThR.Tn[5].t18 159.978
R19487 XThR.Tn[5].n18 XThR.Tn[5].t61 159.978
R19488 XThR.Tn[5].n13 XThR.Tn[5].t23 159.978
R19489 XThR.Tn[5].n82 XThR.Tn[5].t54 145.038
R19490 XThR.Tn[5].n77 XThR.Tn[5].t12 145.038
R19491 XThR.Tn[5].n72 XThR.Tn[5].t56 145.038
R19492 XThR.Tn[5].n67 XThR.Tn[5].t41 145.038
R19493 XThR.Tn[5].n62 XThR.Tn[5].t71 145.038
R19494 XThR.Tn[5].n57 XThR.Tn[5].t53 145.038
R19495 XThR.Tn[5].n52 XThR.Tn[5].t58 145.038
R19496 XThR.Tn[5].n47 XThR.Tn[5].t42 145.038
R19497 XThR.Tn[5].n42 XThR.Tn[5].t38 145.038
R19498 XThR.Tn[5].n37 XThR.Tn[5].t69 145.038
R19499 XThR.Tn[5].n32 XThR.Tn[5].t30 145.038
R19500 XThR.Tn[5].n27 XThR.Tn[5].t55 145.038
R19501 XThR.Tn[5].n22 XThR.Tn[5].t28 145.038
R19502 XThR.Tn[5].n17 XThR.Tn[5].t73 145.038
R19503 XThR.Tn[5].n12 XThR.Tn[5].t39 145.038
R19504 XThR.Tn[5].n10 XThR.Tn[5].t17 145.038
R19505 XThR.Tn[5].n83 XThR.Tn[5].t27 143.911
R19506 XThR.Tn[5].n78 XThR.Tn[5].t50 143.911
R19507 XThR.Tn[5].n73 XThR.Tn[5].t34 143.911
R19508 XThR.Tn[5].n68 XThR.Tn[5].t15 143.911
R19509 XThR.Tn[5].n63 XThR.Tn[5].t44 143.911
R19510 XThR.Tn[5].n58 XThR.Tn[5].t25 143.911
R19511 XThR.Tn[5].n53 XThR.Tn[5].t36 143.911
R19512 XThR.Tn[5].n48 XThR.Tn[5].t16 143.911
R19513 XThR.Tn[5].n43 XThR.Tn[5].t14 143.911
R19514 XThR.Tn[5].n38 XThR.Tn[5].t43 143.911
R19515 XThR.Tn[5].n33 XThR.Tn[5].t67 143.911
R19516 XThR.Tn[5].n28 XThR.Tn[5].t33 143.911
R19517 XThR.Tn[5].n23 XThR.Tn[5].t65 143.911
R19518 XThR.Tn[5].n18 XThR.Tn[5].t48 143.911
R19519 XThR.Tn[5].n13 XThR.Tn[5].t13 143.911
R19520 XThR.Tn[5].n7 XThR.Tn[5].n5 135.249
R19521 XThR.Tn[5].n9 XThR.Tn[5].n3 98.981
R19522 XThR.Tn[5].n8 XThR.Tn[5].n4 98.981
R19523 XThR.Tn[5].n7 XThR.Tn[5].n6 98.981
R19524 XThR.Tn[5].n9 XThR.Tn[5].n8 36.2672
R19525 XThR.Tn[5].n8 XThR.Tn[5].n7 36.2672
R19526 XThR.Tn[5].n88 XThR.Tn[5].n9 32.6405
R19527 XThR.Tn[5].n1 XThR.Tn[5].t9 26.5955
R19528 XThR.Tn[5].n1 XThR.Tn[5].t8 26.5955
R19529 XThR.Tn[5].n0 XThR.Tn[5].t10 26.5955
R19530 XThR.Tn[5].n0 XThR.Tn[5].t11 26.5955
R19531 XThR.Tn[5].n3 XThR.Tn[5].t7 24.9236
R19532 XThR.Tn[5].n3 XThR.Tn[5].t4 24.9236
R19533 XThR.Tn[5].n4 XThR.Tn[5].t6 24.9236
R19534 XThR.Tn[5].n4 XThR.Tn[5].t5 24.9236
R19535 XThR.Tn[5].n5 XThR.Tn[5].t0 24.9236
R19536 XThR.Tn[5].n5 XThR.Tn[5].t1 24.9236
R19537 XThR.Tn[5].n6 XThR.Tn[5].t3 24.9236
R19538 XThR.Tn[5].n6 XThR.Tn[5].t2 24.9236
R19539 XThR.Tn[5].n89 XThR.Tn[5].n2 18.5605
R19540 XThR.Tn[5].n89 XThR.Tn[5].n88 11.5205
R19541 XThR.Tn[5].n88 XThR.Tn[5] 5.71508
R19542 XThR.Tn[5] XThR.Tn[5].n11 5.34038
R19543 XThR.Tn[5].n16 XThR.Tn[5].n15 4.5005
R19544 XThR.Tn[5].n21 XThR.Tn[5].n20 4.5005
R19545 XThR.Tn[5].n26 XThR.Tn[5].n25 4.5005
R19546 XThR.Tn[5].n31 XThR.Tn[5].n30 4.5005
R19547 XThR.Tn[5].n36 XThR.Tn[5].n35 4.5005
R19548 XThR.Tn[5].n41 XThR.Tn[5].n40 4.5005
R19549 XThR.Tn[5].n46 XThR.Tn[5].n45 4.5005
R19550 XThR.Tn[5].n51 XThR.Tn[5].n50 4.5005
R19551 XThR.Tn[5].n56 XThR.Tn[5].n55 4.5005
R19552 XThR.Tn[5].n61 XThR.Tn[5].n60 4.5005
R19553 XThR.Tn[5].n66 XThR.Tn[5].n65 4.5005
R19554 XThR.Tn[5].n71 XThR.Tn[5].n70 4.5005
R19555 XThR.Tn[5].n76 XThR.Tn[5].n75 4.5005
R19556 XThR.Tn[5].n81 XThR.Tn[5].n80 4.5005
R19557 XThR.Tn[5].n86 XThR.Tn[5].n85 4.5005
R19558 XThR.Tn[5].n87 XThR.Tn[5] 3.70586
R19559 XThR.Tn[5].n16 XThR.Tn[5] 2.52282
R19560 XThR.Tn[5].n21 XThR.Tn[5] 2.52282
R19561 XThR.Tn[5].n26 XThR.Tn[5] 2.52282
R19562 XThR.Tn[5].n31 XThR.Tn[5] 2.52282
R19563 XThR.Tn[5].n36 XThR.Tn[5] 2.52282
R19564 XThR.Tn[5].n41 XThR.Tn[5] 2.52282
R19565 XThR.Tn[5].n46 XThR.Tn[5] 2.52282
R19566 XThR.Tn[5].n51 XThR.Tn[5] 2.52282
R19567 XThR.Tn[5].n56 XThR.Tn[5] 2.52282
R19568 XThR.Tn[5].n61 XThR.Tn[5] 2.52282
R19569 XThR.Tn[5].n66 XThR.Tn[5] 2.52282
R19570 XThR.Tn[5].n71 XThR.Tn[5] 2.52282
R19571 XThR.Tn[5].n76 XThR.Tn[5] 2.52282
R19572 XThR.Tn[5].n81 XThR.Tn[5] 2.52282
R19573 XThR.Tn[5].n86 XThR.Tn[5] 2.52282
R19574 XThR.Tn[5].n84 XThR.Tn[5] 1.08677
R19575 XThR.Tn[5].n79 XThR.Tn[5] 1.08677
R19576 XThR.Tn[5].n74 XThR.Tn[5] 1.08677
R19577 XThR.Tn[5].n69 XThR.Tn[5] 1.08677
R19578 XThR.Tn[5].n64 XThR.Tn[5] 1.08677
R19579 XThR.Tn[5].n59 XThR.Tn[5] 1.08677
R19580 XThR.Tn[5].n54 XThR.Tn[5] 1.08677
R19581 XThR.Tn[5].n49 XThR.Tn[5] 1.08677
R19582 XThR.Tn[5].n44 XThR.Tn[5] 1.08677
R19583 XThR.Tn[5].n39 XThR.Tn[5] 1.08677
R19584 XThR.Tn[5].n34 XThR.Tn[5] 1.08677
R19585 XThR.Tn[5].n29 XThR.Tn[5] 1.08677
R19586 XThR.Tn[5].n24 XThR.Tn[5] 1.08677
R19587 XThR.Tn[5].n19 XThR.Tn[5] 1.08677
R19588 XThR.Tn[5].n14 XThR.Tn[5] 1.08677
R19589 XThR.Tn[5] XThR.Tn[5].n16 0.839786
R19590 XThR.Tn[5] XThR.Tn[5].n21 0.839786
R19591 XThR.Tn[5] XThR.Tn[5].n26 0.839786
R19592 XThR.Tn[5] XThR.Tn[5].n31 0.839786
R19593 XThR.Tn[5] XThR.Tn[5].n36 0.839786
R19594 XThR.Tn[5] XThR.Tn[5].n41 0.839786
R19595 XThR.Tn[5] XThR.Tn[5].n46 0.839786
R19596 XThR.Tn[5] XThR.Tn[5].n51 0.839786
R19597 XThR.Tn[5] XThR.Tn[5].n56 0.839786
R19598 XThR.Tn[5] XThR.Tn[5].n61 0.839786
R19599 XThR.Tn[5] XThR.Tn[5].n66 0.839786
R19600 XThR.Tn[5] XThR.Tn[5].n71 0.839786
R19601 XThR.Tn[5] XThR.Tn[5].n76 0.839786
R19602 XThR.Tn[5] XThR.Tn[5].n81 0.839786
R19603 XThR.Tn[5] XThR.Tn[5].n86 0.839786
R19604 XThR.Tn[5] XThR.Tn[5].n89 0.6405
R19605 XThR.Tn[5].n11 XThR.Tn[5] 0.499542
R19606 XThR.Tn[5].n85 XThR.Tn[5] 0.063
R19607 XThR.Tn[5].n80 XThR.Tn[5] 0.063
R19608 XThR.Tn[5].n75 XThR.Tn[5] 0.063
R19609 XThR.Tn[5].n70 XThR.Tn[5] 0.063
R19610 XThR.Tn[5].n65 XThR.Tn[5] 0.063
R19611 XThR.Tn[5].n60 XThR.Tn[5] 0.063
R19612 XThR.Tn[5].n55 XThR.Tn[5] 0.063
R19613 XThR.Tn[5].n50 XThR.Tn[5] 0.063
R19614 XThR.Tn[5].n45 XThR.Tn[5] 0.063
R19615 XThR.Tn[5].n40 XThR.Tn[5] 0.063
R19616 XThR.Tn[5].n35 XThR.Tn[5] 0.063
R19617 XThR.Tn[5].n30 XThR.Tn[5] 0.063
R19618 XThR.Tn[5].n25 XThR.Tn[5] 0.063
R19619 XThR.Tn[5].n20 XThR.Tn[5] 0.063
R19620 XThR.Tn[5].n15 XThR.Tn[5] 0.063
R19621 XThR.Tn[5].n87 XThR.Tn[5] 0.0540714
R19622 XThR.Tn[5] XThR.Tn[5].n87 0.038
R19623 XThR.Tn[5].n11 XThR.Tn[5] 0.0143889
R19624 XThR.Tn[5].n85 XThR.Tn[5].n84 0.00771154
R19625 XThR.Tn[5].n80 XThR.Tn[5].n79 0.00771154
R19626 XThR.Tn[5].n75 XThR.Tn[5].n74 0.00771154
R19627 XThR.Tn[5].n70 XThR.Tn[5].n69 0.00771154
R19628 XThR.Tn[5].n65 XThR.Tn[5].n64 0.00771154
R19629 XThR.Tn[5].n60 XThR.Tn[5].n59 0.00771154
R19630 XThR.Tn[5].n55 XThR.Tn[5].n54 0.00771154
R19631 XThR.Tn[5].n50 XThR.Tn[5].n49 0.00771154
R19632 XThR.Tn[5].n45 XThR.Tn[5].n44 0.00771154
R19633 XThR.Tn[5].n40 XThR.Tn[5].n39 0.00771154
R19634 XThR.Tn[5].n35 XThR.Tn[5].n34 0.00771154
R19635 XThR.Tn[5].n30 XThR.Tn[5].n29 0.00771154
R19636 XThR.Tn[5].n25 XThR.Tn[5].n24 0.00771154
R19637 XThR.Tn[5].n20 XThR.Tn[5].n19 0.00771154
R19638 XThR.Tn[5].n15 XThR.Tn[5].n14 0.00771154
R19639 XThC.Tn[4].n2 XThC.Tn[4].n1 332.332
R19640 XThC.Tn[4].n2 XThC.Tn[4].n0 296.493
R19641 XThC.Tn[4].n71 XThC.Tn[4].n69 161.365
R19642 XThC.Tn[4].n67 XThC.Tn[4].n65 161.365
R19643 XThC.Tn[4].n63 XThC.Tn[4].n61 161.365
R19644 XThC.Tn[4].n59 XThC.Tn[4].n57 161.365
R19645 XThC.Tn[4].n55 XThC.Tn[4].n53 161.365
R19646 XThC.Tn[4].n51 XThC.Tn[4].n49 161.365
R19647 XThC.Tn[4].n47 XThC.Tn[4].n45 161.365
R19648 XThC.Tn[4].n43 XThC.Tn[4].n41 161.365
R19649 XThC.Tn[4].n39 XThC.Tn[4].n37 161.365
R19650 XThC.Tn[4].n35 XThC.Tn[4].n33 161.365
R19651 XThC.Tn[4].n31 XThC.Tn[4].n29 161.365
R19652 XThC.Tn[4].n27 XThC.Tn[4].n25 161.365
R19653 XThC.Tn[4].n23 XThC.Tn[4].n21 161.365
R19654 XThC.Tn[4].n19 XThC.Tn[4].n17 161.365
R19655 XThC.Tn[4].n15 XThC.Tn[4].n13 161.365
R19656 XThC.Tn[4].n12 XThC.Tn[4].n10 161.365
R19657 XThC.Tn[4].n69 XThC.Tn[4].t32 161.202
R19658 XThC.Tn[4].n65 XThC.Tn[4].t22 161.202
R19659 XThC.Tn[4].n61 XThC.Tn[4].t41 161.202
R19660 XThC.Tn[4].n57 XThC.Tn[4].t38 161.202
R19661 XThC.Tn[4].n53 XThC.Tn[4].t30 161.202
R19662 XThC.Tn[4].n49 XThC.Tn[4].t17 161.202
R19663 XThC.Tn[4].n45 XThC.Tn[4].t16 161.202
R19664 XThC.Tn[4].n41 XThC.Tn[4].t29 161.202
R19665 XThC.Tn[4].n37 XThC.Tn[4].t27 161.202
R19666 XThC.Tn[4].n33 XThC.Tn[4].t18 161.202
R19667 XThC.Tn[4].n29 XThC.Tn[4].t37 161.202
R19668 XThC.Tn[4].n25 XThC.Tn[4].t36 161.202
R19669 XThC.Tn[4].n21 XThC.Tn[4].t15 161.202
R19670 XThC.Tn[4].n17 XThC.Tn[4].t13 161.202
R19671 XThC.Tn[4].n13 XThC.Tn[4].t43 161.202
R19672 XThC.Tn[4].n10 XThC.Tn[4].t26 161.202
R19673 XThC.Tn[4].n69 XThC.Tn[4].t35 145.137
R19674 XThC.Tn[4].n65 XThC.Tn[4].t25 145.137
R19675 XThC.Tn[4].n61 XThC.Tn[4].t12 145.137
R19676 XThC.Tn[4].n57 XThC.Tn[4].t42 145.137
R19677 XThC.Tn[4].n53 XThC.Tn[4].t34 145.137
R19678 XThC.Tn[4].n49 XThC.Tn[4].t23 145.137
R19679 XThC.Tn[4].n45 XThC.Tn[4].t21 145.137
R19680 XThC.Tn[4].n41 XThC.Tn[4].t33 145.137
R19681 XThC.Tn[4].n37 XThC.Tn[4].t31 145.137
R19682 XThC.Tn[4].n33 XThC.Tn[4].t24 145.137
R19683 XThC.Tn[4].n29 XThC.Tn[4].t40 145.137
R19684 XThC.Tn[4].n25 XThC.Tn[4].t39 145.137
R19685 XThC.Tn[4].n21 XThC.Tn[4].t20 145.137
R19686 XThC.Tn[4].n17 XThC.Tn[4].t19 145.137
R19687 XThC.Tn[4].n13 XThC.Tn[4].t14 145.137
R19688 XThC.Tn[4].n10 XThC.Tn[4].t28 145.137
R19689 XThC.Tn[4].n7 XThC.Tn[4].n6 135.248
R19690 XThC.Tn[4].n9 XThC.Tn[4].n3 98.982
R19691 XThC.Tn[4].n8 XThC.Tn[4].n4 98.982
R19692 XThC.Tn[4].n7 XThC.Tn[4].n5 98.982
R19693 XThC.Tn[4].n9 XThC.Tn[4].n8 36.2672
R19694 XThC.Tn[4].n8 XThC.Tn[4].n7 36.2672
R19695 XThC.Tn[4].n73 XThC.Tn[4].n9 32.6405
R19696 XThC.Tn[4].n1 XThC.Tn[4].t7 26.5955
R19697 XThC.Tn[4].n1 XThC.Tn[4].t6 26.5955
R19698 XThC.Tn[4].n0 XThC.Tn[4].t5 26.5955
R19699 XThC.Tn[4].n0 XThC.Tn[4].t4 26.5955
R19700 XThC.Tn[4].n3 XThC.Tn[4].t9 24.9236
R19701 XThC.Tn[4].n3 XThC.Tn[4].t8 24.9236
R19702 XThC.Tn[4].n4 XThC.Tn[4].t11 24.9236
R19703 XThC.Tn[4].n4 XThC.Tn[4].t10 24.9236
R19704 XThC.Tn[4].n5 XThC.Tn[4].t2 24.9236
R19705 XThC.Tn[4].n5 XThC.Tn[4].t1 24.9236
R19706 XThC.Tn[4].n6 XThC.Tn[4].t0 24.9236
R19707 XThC.Tn[4].n6 XThC.Tn[4].t3 24.9236
R19708 XThC.Tn[4].n74 XThC.Tn[4].n2 18.5605
R19709 XThC.Tn[4].n74 XThC.Tn[4].n73 11.5205
R19710 XThC.Tn[4] XThC.Tn[4].n12 8.0245
R19711 XThC.Tn[4].n72 XThC.Tn[4].n71 7.9105
R19712 XThC.Tn[4].n68 XThC.Tn[4].n67 7.9105
R19713 XThC.Tn[4].n64 XThC.Tn[4].n63 7.9105
R19714 XThC.Tn[4].n60 XThC.Tn[4].n59 7.9105
R19715 XThC.Tn[4].n56 XThC.Tn[4].n55 7.9105
R19716 XThC.Tn[4].n52 XThC.Tn[4].n51 7.9105
R19717 XThC.Tn[4].n48 XThC.Tn[4].n47 7.9105
R19718 XThC.Tn[4].n44 XThC.Tn[4].n43 7.9105
R19719 XThC.Tn[4].n40 XThC.Tn[4].n39 7.9105
R19720 XThC.Tn[4].n36 XThC.Tn[4].n35 7.9105
R19721 XThC.Tn[4].n32 XThC.Tn[4].n31 7.9105
R19722 XThC.Tn[4].n28 XThC.Tn[4].n27 7.9105
R19723 XThC.Tn[4].n24 XThC.Tn[4].n23 7.9105
R19724 XThC.Tn[4].n20 XThC.Tn[4].n19 7.9105
R19725 XThC.Tn[4].n16 XThC.Tn[4].n15 7.9105
R19726 XThC.Tn[4].n73 XThC.Tn[4] 5.77342
R19727 XThC.Tn[4] XThC.Tn[4].n74 0.6405
R19728 XThC.Tn[4].n16 XThC.Tn[4] 0.235138
R19729 XThC.Tn[4].n20 XThC.Tn[4] 0.235138
R19730 XThC.Tn[4].n24 XThC.Tn[4] 0.235138
R19731 XThC.Tn[4].n28 XThC.Tn[4] 0.235138
R19732 XThC.Tn[4].n32 XThC.Tn[4] 0.235138
R19733 XThC.Tn[4].n36 XThC.Tn[4] 0.235138
R19734 XThC.Tn[4].n40 XThC.Tn[4] 0.235138
R19735 XThC.Tn[4].n44 XThC.Tn[4] 0.235138
R19736 XThC.Tn[4].n48 XThC.Tn[4] 0.235138
R19737 XThC.Tn[4].n52 XThC.Tn[4] 0.235138
R19738 XThC.Tn[4].n56 XThC.Tn[4] 0.235138
R19739 XThC.Tn[4].n60 XThC.Tn[4] 0.235138
R19740 XThC.Tn[4].n64 XThC.Tn[4] 0.235138
R19741 XThC.Tn[4].n68 XThC.Tn[4] 0.235138
R19742 XThC.Tn[4].n72 XThC.Tn[4] 0.235138
R19743 XThC.Tn[4] XThC.Tn[4].n16 0.114505
R19744 XThC.Tn[4] XThC.Tn[4].n20 0.114505
R19745 XThC.Tn[4] XThC.Tn[4].n24 0.114505
R19746 XThC.Tn[4] XThC.Tn[4].n28 0.114505
R19747 XThC.Tn[4] XThC.Tn[4].n32 0.114505
R19748 XThC.Tn[4] XThC.Tn[4].n36 0.114505
R19749 XThC.Tn[4] XThC.Tn[4].n40 0.114505
R19750 XThC.Tn[4] XThC.Tn[4].n44 0.114505
R19751 XThC.Tn[4] XThC.Tn[4].n48 0.114505
R19752 XThC.Tn[4] XThC.Tn[4].n52 0.114505
R19753 XThC.Tn[4] XThC.Tn[4].n56 0.114505
R19754 XThC.Tn[4] XThC.Tn[4].n60 0.114505
R19755 XThC.Tn[4] XThC.Tn[4].n64 0.114505
R19756 XThC.Tn[4] XThC.Tn[4].n68 0.114505
R19757 XThC.Tn[4] XThC.Tn[4].n72 0.114505
R19758 XThC.Tn[4].n71 XThC.Tn[4].n70 0.0599512
R19759 XThC.Tn[4].n67 XThC.Tn[4].n66 0.0599512
R19760 XThC.Tn[4].n63 XThC.Tn[4].n62 0.0599512
R19761 XThC.Tn[4].n59 XThC.Tn[4].n58 0.0599512
R19762 XThC.Tn[4].n55 XThC.Tn[4].n54 0.0599512
R19763 XThC.Tn[4].n51 XThC.Tn[4].n50 0.0599512
R19764 XThC.Tn[4].n47 XThC.Tn[4].n46 0.0599512
R19765 XThC.Tn[4].n43 XThC.Tn[4].n42 0.0599512
R19766 XThC.Tn[4].n39 XThC.Tn[4].n38 0.0599512
R19767 XThC.Tn[4].n35 XThC.Tn[4].n34 0.0599512
R19768 XThC.Tn[4].n31 XThC.Tn[4].n30 0.0599512
R19769 XThC.Tn[4].n27 XThC.Tn[4].n26 0.0599512
R19770 XThC.Tn[4].n23 XThC.Tn[4].n22 0.0599512
R19771 XThC.Tn[4].n19 XThC.Tn[4].n18 0.0599512
R19772 XThC.Tn[4].n15 XThC.Tn[4].n14 0.0599512
R19773 XThC.Tn[4].n12 XThC.Tn[4].n11 0.0599512
R19774 XThC.Tn[4].n70 XThC.Tn[4] 0.0469286
R19775 XThC.Tn[4].n66 XThC.Tn[4] 0.0469286
R19776 XThC.Tn[4].n62 XThC.Tn[4] 0.0469286
R19777 XThC.Tn[4].n58 XThC.Tn[4] 0.0469286
R19778 XThC.Tn[4].n54 XThC.Tn[4] 0.0469286
R19779 XThC.Tn[4].n50 XThC.Tn[4] 0.0469286
R19780 XThC.Tn[4].n46 XThC.Tn[4] 0.0469286
R19781 XThC.Tn[4].n42 XThC.Tn[4] 0.0469286
R19782 XThC.Tn[4].n38 XThC.Tn[4] 0.0469286
R19783 XThC.Tn[4].n34 XThC.Tn[4] 0.0469286
R19784 XThC.Tn[4].n30 XThC.Tn[4] 0.0469286
R19785 XThC.Tn[4].n26 XThC.Tn[4] 0.0469286
R19786 XThC.Tn[4].n22 XThC.Tn[4] 0.0469286
R19787 XThC.Tn[4].n18 XThC.Tn[4] 0.0469286
R19788 XThC.Tn[4].n14 XThC.Tn[4] 0.0469286
R19789 XThC.Tn[4].n11 XThC.Tn[4] 0.0469286
R19790 XThC.Tn[4].n70 XThC.Tn[4] 0.0401341
R19791 XThC.Tn[4].n66 XThC.Tn[4] 0.0401341
R19792 XThC.Tn[4].n62 XThC.Tn[4] 0.0401341
R19793 XThC.Tn[4].n58 XThC.Tn[4] 0.0401341
R19794 XThC.Tn[4].n54 XThC.Tn[4] 0.0401341
R19795 XThC.Tn[4].n50 XThC.Tn[4] 0.0401341
R19796 XThC.Tn[4].n46 XThC.Tn[4] 0.0401341
R19797 XThC.Tn[4].n42 XThC.Tn[4] 0.0401341
R19798 XThC.Tn[4].n38 XThC.Tn[4] 0.0401341
R19799 XThC.Tn[4].n34 XThC.Tn[4] 0.0401341
R19800 XThC.Tn[4].n30 XThC.Tn[4] 0.0401341
R19801 XThC.Tn[4].n26 XThC.Tn[4] 0.0401341
R19802 XThC.Tn[4].n22 XThC.Tn[4] 0.0401341
R19803 XThC.Tn[4].n18 XThC.Tn[4] 0.0401341
R19804 XThC.Tn[4].n14 XThC.Tn[4] 0.0401341
R19805 XThC.Tn[4].n11 XThC.Tn[4] 0.0401341
R19806 XThC.Tn[2].n2 XThC.Tn[2].n1 332.332
R19807 XThC.Tn[2].n2 XThC.Tn[2].n0 296.493
R19808 XThC.Tn[2].n71 XThC.Tn[2].n69 161.365
R19809 XThC.Tn[2].n67 XThC.Tn[2].n65 161.365
R19810 XThC.Tn[2].n63 XThC.Tn[2].n61 161.365
R19811 XThC.Tn[2].n59 XThC.Tn[2].n57 161.365
R19812 XThC.Tn[2].n55 XThC.Tn[2].n53 161.365
R19813 XThC.Tn[2].n51 XThC.Tn[2].n49 161.365
R19814 XThC.Tn[2].n47 XThC.Tn[2].n45 161.365
R19815 XThC.Tn[2].n43 XThC.Tn[2].n41 161.365
R19816 XThC.Tn[2].n39 XThC.Tn[2].n37 161.365
R19817 XThC.Tn[2].n35 XThC.Tn[2].n33 161.365
R19818 XThC.Tn[2].n31 XThC.Tn[2].n29 161.365
R19819 XThC.Tn[2].n27 XThC.Tn[2].n25 161.365
R19820 XThC.Tn[2].n23 XThC.Tn[2].n21 161.365
R19821 XThC.Tn[2].n19 XThC.Tn[2].n17 161.365
R19822 XThC.Tn[2].n15 XThC.Tn[2].n13 161.365
R19823 XThC.Tn[2].n12 XThC.Tn[2].n10 161.365
R19824 XThC.Tn[2].n69 XThC.Tn[2].t24 161.202
R19825 XThC.Tn[2].n65 XThC.Tn[2].t14 161.202
R19826 XThC.Tn[2].n61 XThC.Tn[2].t33 161.202
R19827 XThC.Tn[2].n57 XThC.Tn[2].t30 161.202
R19828 XThC.Tn[2].n53 XThC.Tn[2].t22 161.202
R19829 XThC.Tn[2].n49 XThC.Tn[2].t41 161.202
R19830 XThC.Tn[2].n45 XThC.Tn[2].t40 161.202
R19831 XThC.Tn[2].n41 XThC.Tn[2].t21 161.202
R19832 XThC.Tn[2].n37 XThC.Tn[2].t19 161.202
R19833 XThC.Tn[2].n33 XThC.Tn[2].t42 161.202
R19834 XThC.Tn[2].n29 XThC.Tn[2].t29 161.202
R19835 XThC.Tn[2].n25 XThC.Tn[2].t28 161.202
R19836 XThC.Tn[2].n21 XThC.Tn[2].t39 161.202
R19837 XThC.Tn[2].n17 XThC.Tn[2].t37 161.202
R19838 XThC.Tn[2].n13 XThC.Tn[2].t35 161.202
R19839 XThC.Tn[2].n10 XThC.Tn[2].t18 161.202
R19840 XThC.Tn[2].n69 XThC.Tn[2].t27 145.137
R19841 XThC.Tn[2].n65 XThC.Tn[2].t17 145.137
R19842 XThC.Tn[2].n61 XThC.Tn[2].t36 145.137
R19843 XThC.Tn[2].n57 XThC.Tn[2].t34 145.137
R19844 XThC.Tn[2].n53 XThC.Tn[2].t26 145.137
R19845 XThC.Tn[2].n49 XThC.Tn[2].t15 145.137
R19846 XThC.Tn[2].n45 XThC.Tn[2].t13 145.137
R19847 XThC.Tn[2].n41 XThC.Tn[2].t25 145.137
R19848 XThC.Tn[2].n37 XThC.Tn[2].t23 145.137
R19849 XThC.Tn[2].n33 XThC.Tn[2].t16 145.137
R19850 XThC.Tn[2].n29 XThC.Tn[2].t32 145.137
R19851 XThC.Tn[2].n25 XThC.Tn[2].t31 145.137
R19852 XThC.Tn[2].n21 XThC.Tn[2].t12 145.137
R19853 XThC.Tn[2].n17 XThC.Tn[2].t43 145.137
R19854 XThC.Tn[2].n13 XThC.Tn[2].t38 145.137
R19855 XThC.Tn[2].n10 XThC.Tn[2].t20 145.137
R19856 XThC.Tn[2].n7 XThC.Tn[2].n6 135.248
R19857 XThC.Tn[2].n9 XThC.Tn[2].n3 98.982
R19858 XThC.Tn[2].n8 XThC.Tn[2].n4 98.982
R19859 XThC.Tn[2].n7 XThC.Tn[2].n5 98.982
R19860 XThC.Tn[2].n9 XThC.Tn[2].n8 36.2672
R19861 XThC.Tn[2].n8 XThC.Tn[2].n7 36.2672
R19862 XThC.Tn[2].n74 XThC.Tn[2].n9 32.6405
R19863 XThC.Tn[2].n1 XThC.Tn[2].t3 26.5955
R19864 XThC.Tn[2].n1 XThC.Tn[2].t2 26.5955
R19865 XThC.Tn[2].n0 XThC.Tn[2].t5 26.5955
R19866 XThC.Tn[2].n0 XThC.Tn[2].t4 26.5955
R19867 XThC.Tn[2].n3 XThC.Tn[2].t9 24.9236
R19868 XThC.Tn[2].n3 XThC.Tn[2].t8 24.9236
R19869 XThC.Tn[2].n4 XThC.Tn[2].t7 24.9236
R19870 XThC.Tn[2].n4 XThC.Tn[2].t6 24.9236
R19871 XThC.Tn[2].n5 XThC.Tn[2].t1 24.9236
R19872 XThC.Tn[2].n5 XThC.Tn[2].t10 24.9236
R19873 XThC.Tn[2].n6 XThC.Tn[2].t11 24.9236
R19874 XThC.Tn[2].n6 XThC.Tn[2].t0 24.9236
R19875 XThC.Tn[2].n75 XThC.Tn[2].n2 18.5605
R19876 XThC.Tn[2].n75 XThC.Tn[2].n74 11.5205
R19877 XThC.Tn[2] XThC.Tn[2].n12 8.0245
R19878 XThC.Tn[2].n72 XThC.Tn[2].n71 7.9105
R19879 XThC.Tn[2].n68 XThC.Tn[2].n67 7.9105
R19880 XThC.Tn[2].n64 XThC.Tn[2].n63 7.9105
R19881 XThC.Tn[2].n60 XThC.Tn[2].n59 7.9105
R19882 XThC.Tn[2].n56 XThC.Tn[2].n55 7.9105
R19883 XThC.Tn[2].n52 XThC.Tn[2].n51 7.9105
R19884 XThC.Tn[2].n48 XThC.Tn[2].n47 7.9105
R19885 XThC.Tn[2].n44 XThC.Tn[2].n43 7.9105
R19886 XThC.Tn[2].n40 XThC.Tn[2].n39 7.9105
R19887 XThC.Tn[2].n36 XThC.Tn[2].n35 7.9105
R19888 XThC.Tn[2].n32 XThC.Tn[2].n31 7.9105
R19889 XThC.Tn[2].n28 XThC.Tn[2].n27 7.9105
R19890 XThC.Tn[2].n24 XThC.Tn[2].n23 7.9105
R19891 XThC.Tn[2].n20 XThC.Tn[2].n19 7.9105
R19892 XThC.Tn[2].n16 XThC.Tn[2].n15 7.9105
R19893 XThC.Tn[2].n73 XThC.Tn[2] 5.58686
R19894 XThC.Tn[2].n74 XThC.Tn[2].n73 4.6005
R19895 XThC.Tn[2].n73 XThC.Tn[2] 1.83383
R19896 XThC.Tn[2] XThC.Tn[2].n75 0.6405
R19897 XThC.Tn[2].n16 XThC.Tn[2] 0.235138
R19898 XThC.Tn[2].n20 XThC.Tn[2] 0.235138
R19899 XThC.Tn[2].n24 XThC.Tn[2] 0.235138
R19900 XThC.Tn[2].n28 XThC.Tn[2] 0.235138
R19901 XThC.Tn[2].n32 XThC.Tn[2] 0.235138
R19902 XThC.Tn[2].n36 XThC.Tn[2] 0.235138
R19903 XThC.Tn[2].n40 XThC.Tn[2] 0.235138
R19904 XThC.Tn[2].n44 XThC.Tn[2] 0.235138
R19905 XThC.Tn[2].n48 XThC.Tn[2] 0.235138
R19906 XThC.Tn[2].n52 XThC.Tn[2] 0.235138
R19907 XThC.Tn[2].n56 XThC.Tn[2] 0.235138
R19908 XThC.Tn[2].n60 XThC.Tn[2] 0.235138
R19909 XThC.Tn[2].n64 XThC.Tn[2] 0.235138
R19910 XThC.Tn[2].n68 XThC.Tn[2] 0.235138
R19911 XThC.Tn[2].n72 XThC.Tn[2] 0.235138
R19912 XThC.Tn[2] XThC.Tn[2].n16 0.114505
R19913 XThC.Tn[2] XThC.Tn[2].n20 0.114505
R19914 XThC.Tn[2] XThC.Tn[2].n24 0.114505
R19915 XThC.Tn[2] XThC.Tn[2].n28 0.114505
R19916 XThC.Tn[2] XThC.Tn[2].n32 0.114505
R19917 XThC.Tn[2] XThC.Tn[2].n36 0.114505
R19918 XThC.Tn[2] XThC.Tn[2].n40 0.114505
R19919 XThC.Tn[2] XThC.Tn[2].n44 0.114505
R19920 XThC.Tn[2] XThC.Tn[2].n48 0.114505
R19921 XThC.Tn[2] XThC.Tn[2].n52 0.114505
R19922 XThC.Tn[2] XThC.Tn[2].n56 0.114505
R19923 XThC.Tn[2] XThC.Tn[2].n60 0.114505
R19924 XThC.Tn[2] XThC.Tn[2].n64 0.114505
R19925 XThC.Tn[2] XThC.Tn[2].n68 0.114505
R19926 XThC.Tn[2] XThC.Tn[2].n72 0.114505
R19927 XThC.Tn[2].n71 XThC.Tn[2].n70 0.0599512
R19928 XThC.Tn[2].n67 XThC.Tn[2].n66 0.0599512
R19929 XThC.Tn[2].n63 XThC.Tn[2].n62 0.0599512
R19930 XThC.Tn[2].n59 XThC.Tn[2].n58 0.0599512
R19931 XThC.Tn[2].n55 XThC.Tn[2].n54 0.0599512
R19932 XThC.Tn[2].n51 XThC.Tn[2].n50 0.0599512
R19933 XThC.Tn[2].n47 XThC.Tn[2].n46 0.0599512
R19934 XThC.Tn[2].n43 XThC.Tn[2].n42 0.0599512
R19935 XThC.Tn[2].n39 XThC.Tn[2].n38 0.0599512
R19936 XThC.Tn[2].n35 XThC.Tn[2].n34 0.0599512
R19937 XThC.Tn[2].n31 XThC.Tn[2].n30 0.0599512
R19938 XThC.Tn[2].n27 XThC.Tn[2].n26 0.0599512
R19939 XThC.Tn[2].n23 XThC.Tn[2].n22 0.0599512
R19940 XThC.Tn[2].n19 XThC.Tn[2].n18 0.0599512
R19941 XThC.Tn[2].n15 XThC.Tn[2].n14 0.0599512
R19942 XThC.Tn[2].n12 XThC.Tn[2].n11 0.0599512
R19943 XThC.Tn[2].n70 XThC.Tn[2] 0.0469286
R19944 XThC.Tn[2].n66 XThC.Tn[2] 0.0469286
R19945 XThC.Tn[2].n62 XThC.Tn[2] 0.0469286
R19946 XThC.Tn[2].n58 XThC.Tn[2] 0.0469286
R19947 XThC.Tn[2].n54 XThC.Tn[2] 0.0469286
R19948 XThC.Tn[2].n50 XThC.Tn[2] 0.0469286
R19949 XThC.Tn[2].n46 XThC.Tn[2] 0.0469286
R19950 XThC.Tn[2].n42 XThC.Tn[2] 0.0469286
R19951 XThC.Tn[2].n38 XThC.Tn[2] 0.0469286
R19952 XThC.Tn[2].n34 XThC.Tn[2] 0.0469286
R19953 XThC.Tn[2].n30 XThC.Tn[2] 0.0469286
R19954 XThC.Tn[2].n26 XThC.Tn[2] 0.0469286
R19955 XThC.Tn[2].n22 XThC.Tn[2] 0.0469286
R19956 XThC.Tn[2].n18 XThC.Tn[2] 0.0469286
R19957 XThC.Tn[2].n14 XThC.Tn[2] 0.0469286
R19958 XThC.Tn[2].n11 XThC.Tn[2] 0.0469286
R19959 XThC.Tn[2].n70 XThC.Tn[2] 0.0401341
R19960 XThC.Tn[2].n66 XThC.Tn[2] 0.0401341
R19961 XThC.Tn[2].n62 XThC.Tn[2] 0.0401341
R19962 XThC.Tn[2].n58 XThC.Tn[2] 0.0401341
R19963 XThC.Tn[2].n54 XThC.Tn[2] 0.0401341
R19964 XThC.Tn[2].n50 XThC.Tn[2] 0.0401341
R19965 XThC.Tn[2].n46 XThC.Tn[2] 0.0401341
R19966 XThC.Tn[2].n42 XThC.Tn[2] 0.0401341
R19967 XThC.Tn[2].n38 XThC.Tn[2] 0.0401341
R19968 XThC.Tn[2].n34 XThC.Tn[2] 0.0401341
R19969 XThC.Tn[2].n30 XThC.Tn[2] 0.0401341
R19970 XThC.Tn[2].n26 XThC.Tn[2] 0.0401341
R19971 XThC.Tn[2].n22 XThC.Tn[2] 0.0401341
R19972 XThC.Tn[2].n18 XThC.Tn[2] 0.0401341
R19973 XThC.Tn[2].n14 XThC.Tn[2] 0.0401341
R19974 XThC.Tn[2].n11 XThC.Tn[2] 0.0401341
R19975 Vbias.n512 Vbias.t5 651.571
R19976 Vbias.n512 Vbias.t2 651.571
R19977 Vbias.n513 Vbias.t3 651.571
R19978 Vbias.n513 Vbias.t4 651.571
R19979 Vbias.n509 Vbias.t181 119.309
R19980 Vbias.n507 Vbias.t24 119.309
R19981 Vbias.n505 Vbias.t12 119.309
R19982 Vbias.n503 Vbias.t248 119.309
R19983 Vbias.n501 Vbias.t95 119.309
R19984 Vbias.n499 Vbias.t75 119.309
R19985 Vbias.n497 Vbias.t246 119.309
R19986 Vbias.n495 Vbias.t169 119.309
R19987 Vbias.n493 Vbias.t147 119.309
R19988 Vbias.n491 Vbias.t60 119.309
R19989 Vbias.n489 Vbias.t227 119.309
R19990 Vbias.n487 Vbias.t141 119.309
R19991 Vbias.n485 Vbias.t56 119.309
R19992 Vbias.n483 Vbias.t41 119.309
R19993 Vbias.n481 Vbias.t201 119.309
R19994 Vbias.n480 Vbias.t129 119.309
R19995 Vbias.n477 Vbias.t110 119.309
R19996 Vbias.n475 Vbias.t210 119.309
R19997 Vbias.n473 Vbias.t193 119.309
R19998 Vbias.n471 Vbias.t173 119.309
R19999 Vbias.n469 Vbias.t25 119.309
R20000 Vbias.n467 Vbias.t258 119.309
R20001 Vbias.n465 Vbias.t171 119.309
R20002 Vbias.n463 Vbias.t96 119.309
R20003 Vbias.n461 Vbias.t76 119.309
R20004 Vbias.n459 Vbias.t247 119.309
R20005 Vbias.n457 Vbias.t156 119.309
R20006 Vbias.n455 Vbias.t69 119.309
R20007 Vbias.n453 Vbias.t242 119.309
R20008 Vbias.n451 Vbias.t229 119.309
R20009 Vbias.n449 Vbias.t130 119.309
R20010 Vbias.n448 Vbias.t57 119.309
R20011 Vbias.n445 Vbias.t146 119.309
R20012 Vbias.n443 Vbias.t238 119.309
R20013 Vbias.n441 Vbias.t225 119.309
R20014 Vbias.n439 Vbias.t205 119.309
R20015 Vbias.n437 Vbias.t52 119.309
R20016 Vbias.n435 Vbias.t32 119.309
R20017 Vbias.n433 Vbias.t199 119.309
R20018 Vbias.n431 Vbias.t125 119.309
R20019 Vbias.n429 Vbias.t102 119.309
R20020 Vbias.n427 Vbias.t18 119.309
R20021 Vbias.n425 Vbias.t183 119.309
R20022 Vbias.n423 Vbias.t99 119.309
R20023 Vbias.n421 Vbias.t14 119.309
R20024 Vbias.n419 Vbias.t261 119.309
R20025 Vbias.n417 Vbias.t160 119.309
R20026 Vbias.n416 Vbias.t87 119.309
R20027 Vbias.n413 Vbias.t73 119.309
R20028 Vbias.n411 Vbias.t165 119.309
R20029 Vbias.n409 Vbias.t153 119.309
R20030 Vbias.n407 Vbias.t133 119.309
R20031 Vbias.n405 Vbias.t239 119.309
R20032 Vbias.n403 Vbias.t217 119.309
R20033 Vbias.n401 Vbias.t126 119.309
R20034 Vbias.n399 Vbias.t53 119.309
R20035 Vbias.n397 Vbias.t33 119.309
R20036 Vbias.n395 Vbias.t200 119.309
R20037 Vbias.n393 Vbias.t112 119.309
R20038 Vbias.n391 Vbias.t29 119.309
R20039 Vbias.n389 Vbias.t196 119.309
R20040 Vbias.n387 Vbias.t185 119.309
R20041 Vbias.n385 Vbias.t88 119.309
R20042 Vbias.n384 Vbias.t16 119.309
R20043 Vbias.n381 Vbias.t255 119.309
R20044 Vbias.n379 Vbias.t92 119.309
R20045 Vbias.n377 Vbias.t81 119.309
R20046 Vbias.n375 Vbias.t62 119.309
R20047 Vbias.n373 Vbias.t166 119.309
R20048 Vbias.n371 Vbias.t144 119.309
R20049 Vbias.n369 Vbias.t54 119.309
R20050 Vbias.n367 Vbias.t240 119.309
R20051 Vbias.n365 Vbias.t219 119.309
R20052 Vbias.n363 Vbias.t127 119.309
R20053 Vbias.n361 Vbias.t40 119.309
R20054 Vbias.n359 Vbias.t213 119.309
R20055 Vbias.n357 Vbias.t124 119.309
R20056 Vbias.n355 Vbias.t113 119.309
R20057 Vbias.n353 Vbias.t17 119.309
R20058 Vbias.n352 Vbias.t198 119.309
R20059 Vbias.n349 Vbias.t176 119.309
R20060 Vbias.n347 Vbias.t20 119.309
R20061 Vbias.n345 Vbias.t7 119.309
R20062 Vbias.n343 Vbias.t243 119.309
R20063 Vbias.n341 Vbias.t90 119.309
R20064 Vbias.n339 Vbias.t65 119.309
R20065 Vbias.n337 Vbias.t236 119.309
R20066 Vbias.n335 Vbias.t163 119.309
R20067 Vbias.n333 Vbias.t138 119.309
R20068 Vbias.n331 Vbias.t50 119.309
R20069 Vbias.n329 Vbias.t221 119.309
R20070 Vbias.n327 Vbias.t135 119.309
R20071 Vbias.n325 Vbias.t48 119.309
R20072 Vbias.n323 Vbias.t37 119.309
R20073 Vbias.n321 Vbias.t195 119.309
R20074 Vbias.n320 Vbias.t121 119.309
R20075 Vbias.n317 Vbias.t105 119.309
R20076 Vbias.n315 Vbias.t204 119.309
R20077 Vbias.n313 Vbias.t187 119.309
R20078 Vbias.n311 Vbias.t168 119.309
R20079 Vbias.n309 Vbias.t21 119.309
R20080 Vbias.n307 Vbias.t251 119.309
R20081 Vbias.n305 Vbias.t164 119.309
R20082 Vbias.n303 Vbias.t91 119.309
R20083 Vbias.n301 Vbias.t68 119.309
R20084 Vbias.n299 Vbias.t237 119.309
R20085 Vbias.n297 Vbias.t150 119.309
R20086 Vbias.n295 Vbias.t63 119.309
R20087 Vbias.n293 Vbias.t235 119.309
R20088 Vbias.n291 Vbias.t222 119.309
R20089 Vbias.n289 Vbias.t122 119.309
R20090 Vbias.n288 Vbias.t49 119.309
R20091 Vbias.n285 Vbias.t137 119.309
R20092 Vbias.n283 Vbias.t232 119.309
R20093 Vbias.n281 Vbias.t220 119.309
R20094 Vbias.n279 Vbias.t197 119.309
R20095 Vbias.n277 Vbias.t44 119.309
R20096 Vbias.n275 Vbias.t27 119.309
R20097 Vbias.n273 Vbias.t190 119.309
R20098 Vbias.n271 Vbias.t118 119.309
R20099 Vbias.n269 Vbias.t98 119.309
R20100 Vbias.n267 Vbias.t11 119.309
R20101 Vbias.n265 Vbias.t179 119.309
R20102 Vbias.n263 Vbias.t93 119.309
R20103 Vbias.n261 Vbias.t8 119.309
R20104 Vbias.n259 Vbias.t257 119.309
R20105 Vbias.n257 Vbias.t154 119.309
R20106 Vbias.n256 Vbias.t82 119.309
R20107 Vbias.n253 Vbias.t64 119.309
R20108 Vbias.n251 Vbias.t161 119.309
R20109 Vbias.n249 Vbias.t149 119.309
R20110 Vbias.n247 Vbias.t123 119.309
R20111 Vbias.n245 Vbias.t233 119.309
R20112 Vbias.n243 Vbias.t211 119.309
R20113 Vbias.n241 Vbias.t119 119.309
R20114 Vbias.n239 Vbias.t45 119.309
R20115 Vbias.n237 Vbias.t28 119.309
R20116 Vbias.n235 Vbias.t192 119.309
R20117 Vbias.n233 Vbias.t107 119.309
R20118 Vbias.n231 Vbias.t23 119.309
R20119 Vbias.n229 Vbias.t188 119.309
R20120 Vbias.n227 Vbias.t180 119.309
R20121 Vbias.n225 Vbias.t83 119.309
R20122 Vbias.n224 Vbias.t9 119.309
R20123 Vbias.n221 Vbias.t250 119.309
R20124 Vbias.n219 Vbias.t89 119.309
R20125 Vbias.n217 Vbias.t80 119.309
R20126 Vbias.n215 Vbias.t51 119.309
R20127 Vbias.n213 Vbias.t162 119.309
R20128 Vbias.n211 Vbias.t136 119.309
R20129 Vbias.n209 Vbias.t46 119.309
R20130 Vbias.n207 Vbias.t234 119.309
R20131 Vbias.n205 Vbias.t212 119.309
R20132 Vbias.n203 Vbias.t120 119.309
R20133 Vbias.n201 Vbias.t36 119.309
R20134 Vbias.n199 Vbias.t208 119.309
R20135 Vbias.n197 Vbias.t117 119.309
R20136 Vbias.n195 Vbias.t108 119.309
R20137 Vbias.n193 Vbias.t10 119.309
R20138 Vbias.n192 Vbias.t189 119.309
R20139 Vbias.n189 Vbias.t109 119.309
R20140 Vbias.n187 Vbias.t207 119.309
R20141 Vbias.n185 Vbias.t191 119.309
R20142 Vbias.n183 Vbias.t172 119.309
R20143 Vbias.n181 Vbias.t22 119.309
R20144 Vbias.n179 Vbias.t256 119.309
R20145 Vbias.n177 Vbias.t167 119.309
R20146 Vbias.n175 Vbias.t94 119.309
R20147 Vbias.n173 Vbias.t74 119.309
R20148 Vbias.n171 Vbias.t244 119.309
R20149 Vbias.n169 Vbias.t155 119.309
R20150 Vbias.n167 Vbias.t66 119.309
R20151 Vbias.n165 Vbias.t241 119.309
R20152 Vbias.n163 Vbias.t226 119.309
R20153 Vbias.n161 Vbias.t128 119.309
R20154 Vbias.n160 Vbias.t55 119.309
R20155 Vbias.n157 Vbias.t249 119.309
R20156 Vbias.n155 Vbias.t85 119.309
R20157 Vbias.n153 Vbias.t78 119.309
R20158 Vbias.n151 Vbias.t47 119.309
R20159 Vbias.n149 Vbias.t159 119.309
R20160 Vbias.n147 Vbias.t134 119.309
R20161 Vbias.n145 Vbias.t43 119.309
R20162 Vbias.n143 Vbias.t231 119.309
R20163 Vbias.n141 Vbias.t209 119.309
R20164 Vbias.n139 Vbias.t116 119.309
R20165 Vbias.n137 Vbias.t34 119.309
R20166 Vbias.n135 Vbias.t206 119.309
R20167 Vbias.n133 Vbias.t115 119.309
R20168 Vbias.n131 Vbias.t103 119.309
R20169 Vbias.n129 Vbias.t6 119.309
R20170 Vbias.n128 Vbias.t186 119.309
R20171 Vbias.n125 Vbias.t86 119.309
R20172 Vbias.n123 Vbias.t175 119.309
R20173 Vbias.n121 Vbias.t170 119.309
R20174 Vbias.n119 Vbias.t148 119.309
R20175 Vbias.n117 Vbias.t252 119.309
R20176 Vbias.n115 Vbias.t228 119.309
R20177 Vbias.n113 Vbias.t143 119.309
R20178 Vbias.n111 Vbias.t70 119.309
R20179 Vbias.n109 Vbias.t42 119.309
R20180 Vbias.n107 Vbias.t218 119.309
R20181 Vbias.n105 Vbias.t131 119.309
R20182 Vbias.n103 Vbias.t38 119.309
R20183 Vbias.n101 Vbias.t214 119.309
R20184 Vbias.n99 Vbias.t203 119.309
R20185 Vbias.n97 Vbias.t100 119.309
R20186 Vbias.n96 Vbias.t30 119.309
R20187 Vbias.n93 Vbias.t13 119.309
R20188 Vbias.n91 Vbias.t104 119.309
R20189 Vbias.n89 Vbias.t97 119.309
R20190 Vbias.n87 Vbias.t77 119.309
R20191 Vbias.n85 Vbias.t177 119.309
R20192 Vbias.n83 Vbias.t157 119.309
R20193 Vbias.n81 Vbias.t71 119.309
R20194 Vbias.n79 Vbias.t253 119.309
R20195 Vbias.n77 Vbias.t230 119.309
R20196 Vbias.n75 Vbias.t145 119.309
R20197 Vbias.n73 Vbias.t58 119.309
R20198 Vbias.n71 Vbias.t224 119.309
R20199 Vbias.n69 Vbias.t139 119.309
R20200 Vbias.n67 Vbias.t132 119.309
R20201 Vbias.n65 Vbias.t31 119.309
R20202 Vbias.n64 Vbias.t215 119.309
R20203 Vbias.n61 Vbias.t194 119.309
R20204 Vbias.n59 Vbias.t35 119.309
R20205 Vbias.n57 Vbias.t26 119.309
R20206 Vbias.n55 Vbias.t259 119.309
R20207 Vbias.n53 Vbias.t106 119.309
R20208 Vbias.n51 Vbias.t84 119.309
R20209 Vbias.n49 Vbias.t254 119.309
R20210 Vbias.n47 Vbias.t178 119.309
R20211 Vbias.n45 Vbias.t158 119.309
R20212 Vbias.n43 Vbias.t72 119.309
R20213 Vbias.n41 Vbias.t245 119.309
R20214 Vbias.n39 Vbias.t152 119.309
R20215 Vbias.n37 Vbias.t67 119.309
R20216 Vbias.n35 Vbias.t59 119.309
R20217 Vbias.n33 Vbias.t216 119.309
R20218 Vbias.n32 Vbias.t140 119.309
R20219 Vbias.n29 Vbias.t61 119.309
R20220 Vbias.n27 Vbias.t151 119.309
R20221 Vbias.n25 Vbias.t142 119.309
R20222 Vbias.n23 Vbias.t114 119.309
R20223 Vbias.n21 Vbias.t223 119.309
R20224 Vbias.n19 Vbias.t202 119.309
R20225 Vbias.n17 Vbias.t111 119.309
R20226 Vbias.n15 Vbias.t39 119.309
R20227 Vbias.n13 Vbias.t19 119.309
R20228 Vbias.n11 Vbias.t184 119.309
R20229 Vbias.n9 Vbias.t101 119.309
R20230 Vbias.n7 Vbias.t15 119.309
R20231 Vbias.n5 Vbias.t182 119.309
R20232 Vbias.n3 Vbias.t174 119.309
R20233 Vbias.n1 Vbias.t79 119.309
R20234 Vbias.n0 Vbias.t260 119.309
R20235 Vbias.n515 Vbias.t0 77.1775
R20236 Vbias.n515 Vbias.t1 34.3847
R20237 Vbias Vbias.n480 8.00727
R20238 Vbias Vbias.n448 8.00727
R20239 Vbias Vbias.n416 8.00727
R20240 Vbias Vbias.n384 8.00727
R20241 Vbias Vbias.n352 8.00727
R20242 Vbias Vbias.n320 8.00727
R20243 Vbias Vbias.n288 8.00727
R20244 Vbias Vbias.n256 8.00727
R20245 Vbias Vbias.n224 8.00727
R20246 Vbias Vbias.n192 8.00727
R20247 Vbias Vbias.n160 8.00727
R20248 Vbias Vbias.n128 8.00727
R20249 Vbias Vbias.n96 8.00727
R20250 Vbias Vbias.n64 8.00727
R20251 Vbias Vbias.n32 8.00727
R20252 Vbias Vbias.n0 8.00727
R20253 Vbias.n510 Vbias.n509 7.9105
R20254 Vbias.n508 Vbias.n507 7.9105
R20255 Vbias.n506 Vbias.n505 7.9105
R20256 Vbias.n504 Vbias.n503 7.9105
R20257 Vbias.n502 Vbias.n501 7.9105
R20258 Vbias.n500 Vbias.n499 7.9105
R20259 Vbias.n498 Vbias.n497 7.9105
R20260 Vbias.n496 Vbias.n495 7.9105
R20261 Vbias.n494 Vbias.n493 7.9105
R20262 Vbias.n492 Vbias.n491 7.9105
R20263 Vbias.n490 Vbias.n489 7.9105
R20264 Vbias.n488 Vbias.n487 7.9105
R20265 Vbias.n486 Vbias.n485 7.9105
R20266 Vbias.n484 Vbias.n483 7.9105
R20267 Vbias.n482 Vbias.n481 7.9105
R20268 Vbias.n478 Vbias.n477 7.9105
R20269 Vbias.n476 Vbias.n475 7.9105
R20270 Vbias.n474 Vbias.n473 7.9105
R20271 Vbias.n472 Vbias.n471 7.9105
R20272 Vbias.n470 Vbias.n469 7.9105
R20273 Vbias.n468 Vbias.n467 7.9105
R20274 Vbias.n466 Vbias.n465 7.9105
R20275 Vbias.n464 Vbias.n463 7.9105
R20276 Vbias.n462 Vbias.n461 7.9105
R20277 Vbias.n460 Vbias.n459 7.9105
R20278 Vbias.n458 Vbias.n457 7.9105
R20279 Vbias.n456 Vbias.n455 7.9105
R20280 Vbias.n454 Vbias.n453 7.9105
R20281 Vbias.n452 Vbias.n451 7.9105
R20282 Vbias.n450 Vbias.n449 7.9105
R20283 Vbias.n446 Vbias.n445 7.9105
R20284 Vbias.n444 Vbias.n443 7.9105
R20285 Vbias.n442 Vbias.n441 7.9105
R20286 Vbias.n440 Vbias.n439 7.9105
R20287 Vbias.n438 Vbias.n437 7.9105
R20288 Vbias.n436 Vbias.n435 7.9105
R20289 Vbias.n434 Vbias.n433 7.9105
R20290 Vbias.n432 Vbias.n431 7.9105
R20291 Vbias.n430 Vbias.n429 7.9105
R20292 Vbias.n428 Vbias.n427 7.9105
R20293 Vbias.n426 Vbias.n425 7.9105
R20294 Vbias.n424 Vbias.n423 7.9105
R20295 Vbias.n422 Vbias.n421 7.9105
R20296 Vbias.n420 Vbias.n419 7.9105
R20297 Vbias.n418 Vbias.n417 7.9105
R20298 Vbias.n414 Vbias.n413 7.9105
R20299 Vbias.n412 Vbias.n411 7.9105
R20300 Vbias.n410 Vbias.n409 7.9105
R20301 Vbias.n408 Vbias.n407 7.9105
R20302 Vbias.n406 Vbias.n405 7.9105
R20303 Vbias.n404 Vbias.n403 7.9105
R20304 Vbias.n402 Vbias.n401 7.9105
R20305 Vbias.n400 Vbias.n399 7.9105
R20306 Vbias.n398 Vbias.n397 7.9105
R20307 Vbias.n396 Vbias.n395 7.9105
R20308 Vbias.n394 Vbias.n393 7.9105
R20309 Vbias.n392 Vbias.n391 7.9105
R20310 Vbias.n390 Vbias.n389 7.9105
R20311 Vbias.n388 Vbias.n387 7.9105
R20312 Vbias.n386 Vbias.n385 7.9105
R20313 Vbias.n382 Vbias.n381 7.9105
R20314 Vbias.n380 Vbias.n379 7.9105
R20315 Vbias.n378 Vbias.n377 7.9105
R20316 Vbias.n376 Vbias.n375 7.9105
R20317 Vbias.n374 Vbias.n373 7.9105
R20318 Vbias.n372 Vbias.n371 7.9105
R20319 Vbias.n370 Vbias.n369 7.9105
R20320 Vbias.n368 Vbias.n367 7.9105
R20321 Vbias.n366 Vbias.n365 7.9105
R20322 Vbias.n364 Vbias.n363 7.9105
R20323 Vbias.n362 Vbias.n361 7.9105
R20324 Vbias.n360 Vbias.n359 7.9105
R20325 Vbias.n358 Vbias.n357 7.9105
R20326 Vbias.n356 Vbias.n355 7.9105
R20327 Vbias.n354 Vbias.n353 7.9105
R20328 Vbias.n350 Vbias.n349 7.9105
R20329 Vbias.n348 Vbias.n347 7.9105
R20330 Vbias.n346 Vbias.n345 7.9105
R20331 Vbias.n344 Vbias.n343 7.9105
R20332 Vbias.n342 Vbias.n341 7.9105
R20333 Vbias.n340 Vbias.n339 7.9105
R20334 Vbias.n338 Vbias.n337 7.9105
R20335 Vbias.n336 Vbias.n335 7.9105
R20336 Vbias.n334 Vbias.n333 7.9105
R20337 Vbias.n332 Vbias.n331 7.9105
R20338 Vbias.n330 Vbias.n329 7.9105
R20339 Vbias.n328 Vbias.n327 7.9105
R20340 Vbias.n326 Vbias.n325 7.9105
R20341 Vbias.n324 Vbias.n323 7.9105
R20342 Vbias.n322 Vbias.n321 7.9105
R20343 Vbias.n318 Vbias.n317 7.9105
R20344 Vbias.n316 Vbias.n315 7.9105
R20345 Vbias.n314 Vbias.n313 7.9105
R20346 Vbias.n312 Vbias.n311 7.9105
R20347 Vbias.n310 Vbias.n309 7.9105
R20348 Vbias.n308 Vbias.n307 7.9105
R20349 Vbias.n306 Vbias.n305 7.9105
R20350 Vbias.n304 Vbias.n303 7.9105
R20351 Vbias.n302 Vbias.n301 7.9105
R20352 Vbias.n300 Vbias.n299 7.9105
R20353 Vbias.n298 Vbias.n297 7.9105
R20354 Vbias.n296 Vbias.n295 7.9105
R20355 Vbias.n294 Vbias.n293 7.9105
R20356 Vbias.n292 Vbias.n291 7.9105
R20357 Vbias.n290 Vbias.n289 7.9105
R20358 Vbias.n286 Vbias.n285 7.9105
R20359 Vbias.n284 Vbias.n283 7.9105
R20360 Vbias.n282 Vbias.n281 7.9105
R20361 Vbias.n280 Vbias.n279 7.9105
R20362 Vbias.n278 Vbias.n277 7.9105
R20363 Vbias.n276 Vbias.n275 7.9105
R20364 Vbias.n274 Vbias.n273 7.9105
R20365 Vbias.n272 Vbias.n271 7.9105
R20366 Vbias.n270 Vbias.n269 7.9105
R20367 Vbias.n268 Vbias.n267 7.9105
R20368 Vbias.n266 Vbias.n265 7.9105
R20369 Vbias.n264 Vbias.n263 7.9105
R20370 Vbias.n262 Vbias.n261 7.9105
R20371 Vbias.n260 Vbias.n259 7.9105
R20372 Vbias.n258 Vbias.n257 7.9105
R20373 Vbias.n254 Vbias.n253 7.9105
R20374 Vbias.n252 Vbias.n251 7.9105
R20375 Vbias.n250 Vbias.n249 7.9105
R20376 Vbias.n248 Vbias.n247 7.9105
R20377 Vbias.n246 Vbias.n245 7.9105
R20378 Vbias.n244 Vbias.n243 7.9105
R20379 Vbias.n242 Vbias.n241 7.9105
R20380 Vbias.n240 Vbias.n239 7.9105
R20381 Vbias.n238 Vbias.n237 7.9105
R20382 Vbias.n236 Vbias.n235 7.9105
R20383 Vbias.n234 Vbias.n233 7.9105
R20384 Vbias.n232 Vbias.n231 7.9105
R20385 Vbias.n230 Vbias.n229 7.9105
R20386 Vbias.n228 Vbias.n227 7.9105
R20387 Vbias.n226 Vbias.n225 7.9105
R20388 Vbias.n222 Vbias.n221 7.9105
R20389 Vbias.n220 Vbias.n219 7.9105
R20390 Vbias.n218 Vbias.n217 7.9105
R20391 Vbias.n216 Vbias.n215 7.9105
R20392 Vbias.n214 Vbias.n213 7.9105
R20393 Vbias.n212 Vbias.n211 7.9105
R20394 Vbias.n210 Vbias.n209 7.9105
R20395 Vbias.n208 Vbias.n207 7.9105
R20396 Vbias.n206 Vbias.n205 7.9105
R20397 Vbias.n204 Vbias.n203 7.9105
R20398 Vbias.n202 Vbias.n201 7.9105
R20399 Vbias.n200 Vbias.n199 7.9105
R20400 Vbias.n198 Vbias.n197 7.9105
R20401 Vbias.n196 Vbias.n195 7.9105
R20402 Vbias.n194 Vbias.n193 7.9105
R20403 Vbias.n190 Vbias.n189 7.9105
R20404 Vbias.n188 Vbias.n187 7.9105
R20405 Vbias.n186 Vbias.n185 7.9105
R20406 Vbias.n184 Vbias.n183 7.9105
R20407 Vbias.n182 Vbias.n181 7.9105
R20408 Vbias.n180 Vbias.n179 7.9105
R20409 Vbias.n178 Vbias.n177 7.9105
R20410 Vbias.n176 Vbias.n175 7.9105
R20411 Vbias.n174 Vbias.n173 7.9105
R20412 Vbias.n172 Vbias.n171 7.9105
R20413 Vbias.n170 Vbias.n169 7.9105
R20414 Vbias.n168 Vbias.n167 7.9105
R20415 Vbias.n166 Vbias.n165 7.9105
R20416 Vbias.n164 Vbias.n163 7.9105
R20417 Vbias.n162 Vbias.n161 7.9105
R20418 Vbias.n158 Vbias.n157 7.9105
R20419 Vbias.n156 Vbias.n155 7.9105
R20420 Vbias.n154 Vbias.n153 7.9105
R20421 Vbias.n152 Vbias.n151 7.9105
R20422 Vbias.n150 Vbias.n149 7.9105
R20423 Vbias.n148 Vbias.n147 7.9105
R20424 Vbias.n146 Vbias.n145 7.9105
R20425 Vbias.n144 Vbias.n143 7.9105
R20426 Vbias.n142 Vbias.n141 7.9105
R20427 Vbias.n140 Vbias.n139 7.9105
R20428 Vbias.n138 Vbias.n137 7.9105
R20429 Vbias.n136 Vbias.n135 7.9105
R20430 Vbias.n134 Vbias.n133 7.9105
R20431 Vbias.n132 Vbias.n131 7.9105
R20432 Vbias.n130 Vbias.n129 7.9105
R20433 Vbias.n126 Vbias.n125 7.9105
R20434 Vbias.n124 Vbias.n123 7.9105
R20435 Vbias.n122 Vbias.n121 7.9105
R20436 Vbias.n120 Vbias.n119 7.9105
R20437 Vbias.n118 Vbias.n117 7.9105
R20438 Vbias.n116 Vbias.n115 7.9105
R20439 Vbias.n114 Vbias.n113 7.9105
R20440 Vbias.n112 Vbias.n111 7.9105
R20441 Vbias.n110 Vbias.n109 7.9105
R20442 Vbias.n108 Vbias.n107 7.9105
R20443 Vbias.n106 Vbias.n105 7.9105
R20444 Vbias.n104 Vbias.n103 7.9105
R20445 Vbias.n102 Vbias.n101 7.9105
R20446 Vbias.n100 Vbias.n99 7.9105
R20447 Vbias.n98 Vbias.n97 7.9105
R20448 Vbias.n94 Vbias.n93 7.9105
R20449 Vbias.n92 Vbias.n91 7.9105
R20450 Vbias.n90 Vbias.n89 7.9105
R20451 Vbias.n88 Vbias.n87 7.9105
R20452 Vbias.n86 Vbias.n85 7.9105
R20453 Vbias.n84 Vbias.n83 7.9105
R20454 Vbias.n82 Vbias.n81 7.9105
R20455 Vbias.n80 Vbias.n79 7.9105
R20456 Vbias.n78 Vbias.n77 7.9105
R20457 Vbias.n76 Vbias.n75 7.9105
R20458 Vbias.n74 Vbias.n73 7.9105
R20459 Vbias.n72 Vbias.n71 7.9105
R20460 Vbias.n70 Vbias.n69 7.9105
R20461 Vbias.n68 Vbias.n67 7.9105
R20462 Vbias.n66 Vbias.n65 7.9105
R20463 Vbias.n62 Vbias.n61 7.9105
R20464 Vbias.n60 Vbias.n59 7.9105
R20465 Vbias.n58 Vbias.n57 7.9105
R20466 Vbias.n56 Vbias.n55 7.9105
R20467 Vbias.n54 Vbias.n53 7.9105
R20468 Vbias.n52 Vbias.n51 7.9105
R20469 Vbias.n50 Vbias.n49 7.9105
R20470 Vbias.n48 Vbias.n47 7.9105
R20471 Vbias.n46 Vbias.n45 7.9105
R20472 Vbias.n44 Vbias.n43 7.9105
R20473 Vbias.n42 Vbias.n41 7.9105
R20474 Vbias.n40 Vbias.n39 7.9105
R20475 Vbias.n38 Vbias.n37 7.9105
R20476 Vbias.n36 Vbias.n35 7.9105
R20477 Vbias.n34 Vbias.n33 7.9105
R20478 Vbias.n30 Vbias.n29 7.9105
R20479 Vbias.n28 Vbias.n27 7.9105
R20480 Vbias.n26 Vbias.n25 7.9105
R20481 Vbias.n24 Vbias.n23 7.9105
R20482 Vbias.n22 Vbias.n21 7.9105
R20483 Vbias.n20 Vbias.n19 7.9105
R20484 Vbias.n18 Vbias.n17 7.9105
R20485 Vbias.n16 Vbias.n15 7.9105
R20486 Vbias.n14 Vbias.n13 7.9105
R20487 Vbias.n12 Vbias.n11 7.9105
R20488 Vbias.n10 Vbias.n9 7.9105
R20489 Vbias.n8 Vbias.n7 7.9105
R20490 Vbias.n6 Vbias.n5 7.9105
R20491 Vbias.n4 Vbias.n3 7.9105
R20492 Vbias.n2 Vbias.n1 7.9105
R20493 Vbias.n514 Vbias.n512 4.78773
R20494 Vbias.n514 Vbias.n513 4.78773
R20495 Vbias.n516 Vbias.n514 2.09636
R20496 Vbias.n511 Vbias 1.6647
R20497 Vbias.n479 Vbias 1.6647
R20498 Vbias.n447 Vbias 1.6647
R20499 Vbias.n415 Vbias 1.6647
R20500 Vbias.n383 Vbias 1.6647
R20501 Vbias.n351 Vbias 1.6647
R20502 Vbias.n319 Vbias 1.6647
R20503 Vbias.n287 Vbias 1.6647
R20504 Vbias.n255 Vbias 1.6647
R20505 Vbias.n223 Vbias 1.6647
R20506 Vbias.n191 Vbias 1.6647
R20507 Vbias.n159 Vbias 1.6647
R20508 Vbias.n127 Vbias 1.6647
R20509 Vbias.n95 Vbias 1.6647
R20510 Vbias.n63 Vbias 1.6647
R20511 Vbias.n31 Vbias 1.6647
R20512 Vbias.n517 Vbias 1.34721
R20513 Vbias Vbias.n516 0.752103
R20514 Vbias.n517 Vbias.n511 0.5692
R20515 Vbias.n516 Vbias.n515 0.515506
R20516 Vbias.n63 Vbias.n31 0.410967
R20517 Vbias.n95 Vbias.n63 0.410967
R20518 Vbias.n127 Vbias.n95 0.410967
R20519 Vbias.n159 Vbias.n127 0.410967
R20520 Vbias.n191 Vbias.n159 0.410967
R20521 Vbias.n223 Vbias.n191 0.410967
R20522 Vbias.n255 Vbias.n223 0.410967
R20523 Vbias.n287 Vbias.n255 0.410967
R20524 Vbias.n319 Vbias.n287 0.410967
R20525 Vbias.n351 Vbias.n319 0.410967
R20526 Vbias.n383 Vbias.n351 0.410967
R20527 Vbias.n415 Vbias.n383 0.410967
R20528 Vbias.n447 Vbias.n415 0.410967
R20529 Vbias.n479 Vbias.n447 0.410967
R20530 Vbias.n511 Vbias.n479 0.410967
R20531 Vbias.n31 Vbias 0.383811
R20532 Vbias.n482 Vbias 0.252372
R20533 Vbias.n484 Vbias 0.252372
R20534 Vbias.n486 Vbias 0.252372
R20535 Vbias.n488 Vbias 0.252372
R20536 Vbias.n490 Vbias 0.252372
R20537 Vbias.n492 Vbias 0.252372
R20538 Vbias.n494 Vbias 0.252372
R20539 Vbias.n496 Vbias 0.252372
R20540 Vbias.n498 Vbias 0.252372
R20541 Vbias.n500 Vbias 0.252372
R20542 Vbias.n502 Vbias 0.252372
R20543 Vbias.n504 Vbias 0.252372
R20544 Vbias.n506 Vbias 0.252372
R20545 Vbias.n508 Vbias 0.252372
R20546 Vbias.n510 Vbias 0.252372
R20547 Vbias.n450 Vbias 0.252372
R20548 Vbias.n452 Vbias 0.252372
R20549 Vbias.n454 Vbias 0.252372
R20550 Vbias.n456 Vbias 0.252372
R20551 Vbias.n458 Vbias 0.252372
R20552 Vbias.n460 Vbias 0.252372
R20553 Vbias.n462 Vbias 0.252372
R20554 Vbias.n464 Vbias 0.252372
R20555 Vbias.n466 Vbias 0.252372
R20556 Vbias.n468 Vbias 0.252372
R20557 Vbias.n470 Vbias 0.252372
R20558 Vbias.n472 Vbias 0.252372
R20559 Vbias.n474 Vbias 0.252372
R20560 Vbias.n476 Vbias 0.252372
R20561 Vbias.n478 Vbias 0.252372
R20562 Vbias.n418 Vbias 0.252372
R20563 Vbias.n420 Vbias 0.252372
R20564 Vbias.n422 Vbias 0.252372
R20565 Vbias.n424 Vbias 0.252372
R20566 Vbias.n426 Vbias 0.252372
R20567 Vbias.n428 Vbias 0.252372
R20568 Vbias.n430 Vbias 0.252372
R20569 Vbias.n432 Vbias 0.252372
R20570 Vbias.n434 Vbias 0.252372
R20571 Vbias.n436 Vbias 0.252372
R20572 Vbias.n438 Vbias 0.252372
R20573 Vbias.n440 Vbias 0.252372
R20574 Vbias.n442 Vbias 0.252372
R20575 Vbias.n444 Vbias 0.252372
R20576 Vbias.n446 Vbias 0.252372
R20577 Vbias.n386 Vbias 0.252372
R20578 Vbias.n388 Vbias 0.252372
R20579 Vbias.n390 Vbias 0.252372
R20580 Vbias.n392 Vbias 0.252372
R20581 Vbias.n394 Vbias 0.252372
R20582 Vbias.n396 Vbias 0.252372
R20583 Vbias.n398 Vbias 0.252372
R20584 Vbias.n400 Vbias 0.252372
R20585 Vbias.n402 Vbias 0.252372
R20586 Vbias.n404 Vbias 0.252372
R20587 Vbias.n406 Vbias 0.252372
R20588 Vbias.n408 Vbias 0.252372
R20589 Vbias.n410 Vbias 0.252372
R20590 Vbias.n412 Vbias 0.252372
R20591 Vbias.n414 Vbias 0.252372
R20592 Vbias.n354 Vbias 0.252372
R20593 Vbias.n356 Vbias 0.252372
R20594 Vbias.n358 Vbias 0.252372
R20595 Vbias.n360 Vbias 0.252372
R20596 Vbias.n362 Vbias 0.252372
R20597 Vbias.n364 Vbias 0.252372
R20598 Vbias.n366 Vbias 0.252372
R20599 Vbias.n368 Vbias 0.252372
R20600 Vbias.n370 Vbias 0.252372
R20601 Vbias.n372 Vbias 0.252372
R20602 Vbias.n374 Vbias 0.252372
R20603 Vbias.n376 Vbias 0.252372
R20604 Vbias.n378 Vbias 0.252372
R20605 Vbias.n380 Vbias 0.252372
R20606 Vbias.n382 Vbias 0.252372
R20607 Vbias.n322 Vbias 0.252372
R20608 Vbias.n324 Vbias 0.252372
R20609 Vbias.n326 Vbias 0.252372
R20610 Vbias.n328 Vbias 0.252372
R20611 Vbias.n330 Vbias 0.252372
R20612 Vbias.n332 Vbias 0.252372
R20613 Vbias.n334 Vbias 0.252372
R20614 Vbias.n336 Vbias 0.252372
R20615 Vbias.n338 Vbias 0.252372
R20616 Vbias.n340 Vbias 0.252372
R20617 Vbias.n342 Vbias 0.252372
R20618 Vbias.n344 Vbias 0.252372
R20619 Vbias.n346 Vbias 0.252372
R20620 Vbias.n348 Vbias 0.252372
R20621 Vbias.n350 Vbias 0.252372
R20622 Vbias.n290 Vbias 0.252372
R20623 Vbias.n292 Vbias 0.252372
R20624 Vbias.n294 Vbias 0.252372
R20625 Vbias.n296 Vbias 0.252372
R20626 Vbias.n298 Vbias 0.252372
R20627 Vbias.n300 Vbias 0.252372
R20628 Vbias.n302 Vbias 0.252372
R20629 Vbias.n304 Vbias 0.252372
R20630 Vbias.n306 Vbias 0.252372
R20631 Vbias.n308 Vbias 0.252372
R20632 Vbias.n310 Vbias 0.252372
R20633 Vbias.n312 Vbias 0.252372
R20634 Vbias.n314 Vbias 0.252372
R20635 Vbias.n316 Vbias 0.252372
R20636 Vbias.n318 Vbias 0.252372
R20637 Vbias.n258 Vbias 0.252372
R20638 Vbias.n260 Vbias 0.252372
R20639 Vbias.n262 Vbias 0.252372
R20640 Vbias.n264 Vbias 0.252372
R20641 Vbias.n266 Vbias 0.252372
R20642 Vbias.n268 Vbias 0.252372
R20643 Vbias.n270 Vbias 0.252372
R20644 Vbias.n272 Vbias 0.252372
R20645 Vbias.n274 Vbias 0.252372
R20646 Vbias.n276 Vbias 0.252372
R20647 Vbias.n278 Vbias 0.252372
R20648 Vbias.n280 Vbias 0.252372
R20649 Vbias.n282 Vbias 0.252372
R20650 Vbias.n284 Vbias 0.252372
R20651 Vbias.n286 Vbias 0.252372
R20652 Vbias.n226 Vbias 0.252372
R20653 Vbias.n228 Vbias 0.252372
R20654 Vbias.n230 Vbias 0.252372
R20655 Vbias.n232 Vbias 0.252372
R20656 Vbias.n234 Vbias 0.252372
R20657 Vbias.n236 Vbias 0.252372
R20658 Vbias.n238 Vbias 0.252372
R20659 Vbias.n240 Vbias 0.252372
R20660 Vbias.n242 Vbias 0.252372
R20661 Vbias.n244 Vbias 0.252372
R20662 Vbias.n246 Vbias 0.252372
R20663 Vbias.n248 Vbias 0.252372
R20664 Vbias.n250 Vbias 0.252372
R20665 Vbias.n252 Vbias 0.252372
R20666 Vbias.n254 Vbias 0.252372
R20667 Vbias.n194 Vbias 0.252372
R20668 Vbias.n196 Vbias 0.252372
R20669 Vbias.n198 Vbias 0.252372
R20670 Vbias.n200 Vbias 0.252372
R20671 Vbias.n202 Vbias 0.252372
R20672 Vbias.n204 Vbias 0.252372
R20673 Vbias.n206 Vbias 0.252372
R20674 Vbias.n208 Vbias 0.252372
R20675 Vbias.n210 Vbias 0.252372
R20676 Vbias.n212 Vbias 0.252372
R20677 Vbias.n214 Vbias 0.252372
R20678 Vbias.n216 Vbias 0.252372
R20679 Vbias.n218 Vbias 0.252372
R20680 Vbias.n220 Vbias 0.252372
R20681 Vbias.n222 Vbias 0.252372
R20682 Vbias.n162 Vbias 0.252372
R20683 Vbias.n164 Vbias 0.252372
R20684 Vbias.n166 Vbias 0.252372
R20685 Vbias.n168 Vbias 0.252372
R20686 Vbias.n170 Vbias 0.252372
R20687 Vbias.n172 Vbias 0.252372
R20688 Vbias.n174 Vbias 0.252372
R20689 Vbias.n176 Vbias 0.252372
R20690 Vbias.n178 Vbias 0.252372
R20691 Vbias.n180 Vbias 0.252372
R20692 Vbias.n182 Vbias 0.252372
R20693 Vbias.n184 Vbias 0.252372
R20694 Vbias.n186 Vbias 0.252372
R20695 Vbias.n188 Vbias 0.252372
R20696 Vbias.n190 Vbias 0.252372
R20697 Vbias.n130 Vbias 0.252372
R20698 Vbias.n132 Vbias 0.252372
R20699 Vbias.n134 Vbias 0.252372
R20700 Vbias.n136 Vbias 0.252372
R20701 Vbias.n138 Vbias 0.252372
R20702 Vbias.n140 Vbias 0.252372
R20703 Vbias.n142 Vbias 0.252372
R20704 Vbias.n144 Vbias 0.252372
R20705 Vbias.n146 Vbias 0.252372
R20706 Vbias.n148 Vbias 0.252372
R20707 Vbias.n150 Vbias 0.252372
R20708 Vbias.n152 Vbias 0.252372
R20709 Vbias.n154 Vbias 0.252372
R20710 Vbias.n156 Vbias 0.252372
R20711 Vbias.n158 Vbias 0.252372
R20712 Vbias.n98 Vbias 0.252372
R20713 Vbias.n100 Vbias 0.252372
R20714 Vbias.n102 Vbias 0.252372
R20715 Vbias.n104 Vbias 0.252372
R20716 Vbias.n106 Vbias 0.252372
R20717 Vbias.n108 Vbias 0.252372
R20718 Vbias.n110 Vbias 0.252372
R20719 Vbias.n112 Vbias 0.252372
R20720 Vbias.n114 Vbias 0.252372
R20721 Vbias.n116 Vbias 0.252372
R20722 Vbias.n118 Vbias 0.252372
R20723 Vbias.n120 Vbias 0.252372
R20724 Vbias.n122 Vbias 0.252372
R20725 Vbias.n124 Vbias 0.252372
R20726 Vbias.n126 Vbias 0.252372
R20727 Vbias.n66 Vbias 0.252372
R20728 Vbias.n68 Vbias 0.252372
R20729 Vbias.n70 Vbias 0.252372
R20730 Vbias.n72 Vbias 0.252372
R20731 Vbias.n74 Vbias 0.252372
R20732 Vbias.n76 Vbias 0.252372
R20733 Vbias.n78 Vbias 0.252372
R20734 Vbias.n80 Vbias 0.252372
R20735 Vbias.n82 Vbias 0.252372
R20736 Vbias.n84 Vbias 0.252372
R20737 Vbias.n86 Vbias 0.252372
R20738 Vbias.n88 Vbias 0.252372
R20739 Vbias.n90 Vbias 0.252372
R20740 Vbias.n92 Vbias 0.252372
R20741 Vbias.n94 Vbias 0.252372
R20742 Vbias.n34 Vbias 0.252372
R20743 Vbias.n36 Vbias 0.252372
R20744 Vbias.n38 Vbias 0.252372
R20745 Vbias.n40 Vbias 0.252372
R20746 Vbias.n42 Vbias 0.252372
R20747 Vbias.n44 Vbias 0.252372
R20748 Vbias.n46 Vbias 0.252372
R20749 Vbias.n48 Vbias 0.252372
R20750 Vbias.n50 Vbias 0.252372
R20751 Vbias.n52 Vbias 0.252372
R20752 Vbias.n54 Vbias 0.252372
R20753 Vbias.n56 Vbias 0.252372
R20754 Vbias.n58 Vbias 0.252372
R20755 Vbias.n60 Vbias 0.252372
R20756 Vbias.n62 Vbias 0.252372
R20757 Vbias.n2 Vbias 0.252372
R20758 Vbias.n4 Vbias 0.252372
R20759 Vbias.n6 Vbias 0.252372
R20760 Vbias.n8 Vbias 0.252372
R20761 Vbias.n10 Vbias 0.252372
R20762 Vbias.n12 Vbias 0.252372
R20763 Vbias.n14 Vbias 0.252372
R20764 Vbias.n16 Vbias 0.252372
R20765 Vbias.n18 Vbias 0.252372
R20766 Vbias.n20 Vbias 0.252372
R20767 Vbias.n22 Vbias 0.252372
R20768 Vbias.n24 Vbias 0.252372
R20769 Vbias.n26 Vbias 0.252372
R20770 Vbias.n28 Vbias 0.252372
R20771 Vbias.n30 Vbias 0.252372
R20772 Vbias Vbias.n517 0.237067
R20773 Vbias Vbias.n482 0.0972718
R20774 Vbias Vbias.n484 0.0972718
R20775 Vbias Vbias.n486 0.0972718
R20776 Vbias Vbias.n488 0.0972718
R20777 Vbias Vbias.n490 0.0972718
R20778 Vbias Vbias.n492 0.0972718
R20779 Vbias Vbias.n494 0.0972718
R20780 Vbias Vbias.n496 0.0972718
R20781 Vbias Vbias.n498 0.0972718
R20782 Vbias Vbias.n500 0.0972718
R20783 Vbias Vbias.n502 0.0972718
R20784 Vbias Vbias.n504 0.0972718
R20785 Vbias Vbias.n506 0.0972718
R20786 Vbias Vbias.n508 0.0972718
R20787 Vbias Vbias.n510 0.0972718
R20788 Vbias Vbias.n450 0.0972718
R20789 Vbias Vbias.n452 0.0972718
R20790 Vbias Vbias.n454 0.0972718
R20791 Vbias Vbias.n456 0.0972718
R20792 Vbias Vbias.n458 0.0972718
R20793 Vbias Vbias.n460 0.0972718
R20794 Vbias Vbias.n462 0.0972718
R20795 Vbias Vbias.n464 0.0972718
R20796 Vbias Vbias.n466 0.0972718
R20797 Vbias Vbias.n468 0.0972718
R20798 Vbias Vbias.n470 0.0972718
R20799 Vbias Vbias.n472 0.0972718
R20800 Vbias Vbias.n474 0.0972718
R20801 Vbias Vbias.n476 0.0972718
R20802 Vbias Vbias.n478 0.0972718
R20803 Vbias Vbias.n418 0.0972718
R20804 Vbias Vbias.n420 0.0972718
R20805 Vbias Vbias.n422 0.0972718
R20806 Vbias Vbias.n424 0.0972718
R20807 Vbias Vbias.n426 0.0972718
R20808 Vbias Vbias.n428 0.0972718
R20809 Vbias Vbias.n430 0.0972718
R20810 Vbias Vbias.n432 0.0972718
R20811 Vbias Vbias.n434 0.0972718
R20812 Vbias Vbias.n436 0.0972718
R20813 Vbias Vbias.n438 0.0972718
R20814 Vbias Vbias.n440 0.0972718
R20815 Vbias Vbias.n442 0.0972718
R20816 Vbias Vbias.n444 0.0972718
R20817 Vbias Vbias.n446 0.0972718
R20818 Vbias Vbias.n386 0.0972718
R20819 Vbias Vbias.n388 0.0972718
R20820 Vbias Vbias.n390 0.0972718
R20821 Vbias Vbias.n392 0.0972718
R20822 Vbias Vbias.n394 0.0972718
R20823 Vbias Vbias.n396 0.0972718
R20824 Vbias Vbias.n398 0.0972718
R20825 Vbias Vbias.n400 0.0972718
R20826 Vbias Vbias.n402 0.0972718
R20827 Vbias Vbias.n404 0.0972718
R20828 Vbias Vbias.n406 0.0972718
R20829 Vbias Vbias.n408 0.0972718
R20830 Vbias Vbias.n410 0.0972718
R20831 Vbias Vbias.n412 0.0972718
R20832 Vbias Vbias.n414 0.0972718
R20833 Vbias Vbias.n354 0.0972718
R20834 Vbias Vbias.n356 0.0972718
R20835 Vbias Vbias.n358 0.0972718
R20836 Vbias Vbias.n360 0.0972718
R20837 Vbias Vbias.n362 0.0972718
R20838 Vbias Vbias.n364 0.0972718
R20839 Vbias Vbias.n366 0.0972718
R20840 Vbias Vbias.n368 0.0972718
R20841 Vbias Vbias.n370 0.0972718
R20842 Vbias Vbias.n372 0.0972718
R20843 Vbias Vbias.n374 0.0972718
R20844 Vbias Vbias.n376 0.0972718
R20845 Vbias Vbias.n378 0.0972718
R20846 Vbias Vbias.n380 0.0972718
R20847 Vbias Vbias.n382 0.0972718
R20848 Vbias Vbias.n322 0.0972718
R20849 Vbias Vbias.n324 0.0972718
R20850 Vbias Vbias.n326 0.0972718
R20851 Vbias Vbias.n328 0.0972718
R20852 Vbias Vbias.n330 0.0972718
R20853 Vbias Vbias.n332 0.0972718
R20854 Vbias Vbias.n334 0.0972718
R20855 Vbias Vbias.n336 0.0972718
R20856 Vbias Vbias.n338 0.0972718
R20857 Vbias Vbias.n340 0.0972718
R20858 Vbias Vbias.n342 0.0972718
R20859 Vbias Vbias.n344 0.0972718
R20860 Vbias Vbias.n346 0.0972718
R20861 Vbias Vbias.n348 0.0972718
R20862 Vbias Vbias.n350 0.0972718
R20863 Vbias Vbias.n290 0.0972718
R20864 Vbias Vbias.n292 0.0972718
R20865 Vbias Vbias.n294 0.0972718
R20866 Vbias Vbias.n296 0.0972718
R20867 Vbias Vbias.n298 0.0972718
R20868 Vbias Vbias.n300 0.0972718
R20869 Vbias Vbias.n302 0.0972718
R20870 Vbias Vbias.n304 0.0972718
R20871 Vbias Vbias.n306 0.0972718
R20872 Vbias Vbias.n308 0.0972718
R20873 Vbias Vbias.n310 0.0972718
R20874 Vbias Vbias.n312 0.0972718
R20875 Vbias Vbias.n314 0.0972718
R20876 Vbias Vbias.n316 0.0972718
R20877 Vbias Vbias.n318 0.0972718
R20878 Vbias Vbias.n258 0.0972718
R20879 Vbias Vbias.n260 0.0972718
R20880 Vbias Vbias.n262 0.0972718
R20881 Vbias Vbias.n264 0.0972718
R20882 Vbias Vbias.n266 0.0972718
R20883 Vbias Vbias.n268 0.0972718
R20884 Vbias Vbias.n270 0.0972718
R20885 Vbias Vbias.n272 0.0972718
R20886 Vbias Vbias.n274 0.0972718
R20887 Vbias Vbias.n276 0.0972718
R20888 Vbias Vbias.n278 0.0972718
R20889 Vbias Vbias.n280 0.0972718
R20890 Vbias Vbias.n282 0.0972718
R20891 Vbias Vbias.n284 0.0972718
R20892 Vbias Vbias.n286 0.0972718
R20893 Vbias Vbias.n226 0.0972718
R20894 Vbias Vbias.n228 0.0972718
R20895 Vbias Vbias.n230 0.0972718
R20896 Vbias Vbias.n232 0.0972718
R20897 Vbias Vbias.n234 0.0972718
R20898 Vbias Vbias.n236 0.0972718
R20899 Vbias Vbias.n238 0.0972718
R20900 Vbias Vbias.n240 0.0972718
R20901 Vbias Vbias.n242 0.0972718
R20902 Vbias Vbias.n244 0.0972718
R20903 Vbias Vbias.n246 0.0972718
R20904 Vbias Vbias.n248 0.0972718
R20905 Vbias Vbias.n250 0.0972718
R20906 Vbias Vbias.n252 0.0972718
R20907 Vbias Vbias.n254 0.0972718
R20908 Vbias Vbias.n194 0.0972718
R20909 Vbias Vbias.n196 0.0972718
R20910 Vbias Vbias.n198 0.0972718
R20911 Vbias Vbias.n200 0.0972718
R20912 Vbias Vbias.n202 0.0972718
R20913 Vbias Vbias.n204 0.0972718
R20914 Vbias Vbias.n206 0.0972718
R20915 Vbias Vbias.n208 0.0972718
R20916 Vbias Vbias.n210 0.0972718
R20917 Vbias Vbias.n212 0.0972718
R20918 Vbias Vbias.n214 0.0972718
R20919 Vbias Vbias.n216 0.0972718
R20920 Vbias Vbias.n218 0.0972718
R20921 Vbias Vbias.n220 0.0972718
R20922 Vbias Vbias.n222 0.0972718
R20923 Vbias Vbias.n162 0.0972718
R20924 Vbias Vbias.n164 0.0972718
R20925 Vbias Vbias.n166 0.0972718
R20926 Vbias Vbias.n168 0.0972718
R20927 Vbias Vbias.n170 0.0972718
R20928 Vbias Vbias.n172 0.0972718
R20929 Vbias Vbias.n174 0.0972718
R20930 Vbias Vbias.n176 0.0972718
R20931 Vbias Vbias.n178 0.0972718
R20932 Vbias Vbias.n180 0.0972718
R20933 Vbias Vbias.n182 0.0972718
R20934 Vbias Vbias.n184 0.0972718
R20935 Vbias Vbias.n186 0.0972718
R20936 Vbias Vbias.n188 0.0972718
R20937 Vbias Vbias.n190 0.0972718
R20938 Vbias Vbias.n130 0.0972718
R20939 Vbias Vbias.n132 0.0972718
R20940 Vbias Vbias.n134 0.0972718
R20941 Vbias Vbias.n136 0.0972718
R20942 Vbias Vbias.n138 0.0972718
R20943 Vbias Vbias.n140 0.0972718
R20944 Vbias Vbias.n142 0.0972718
R20945 Vbias Vbias.n144 0.0972718
R20946 Vbias Vbias.n146 0.0972718
R20947 Vbias Vbias.n148 0.0972718
R20948 Vbias Vbias.n150 0.0972718
R20949 Vbias Vbias.n152 0.0972718
R20950 Vbias Vbias.n154 0.0972718
R20951 Vbias Vbias.n156 0.0972718
R20952 Vbias Vbias.n158 0.0972718
R20953 Vbias Vbias.n98 0.0972718
R20954 Vbias Vbias.n100 0.0972718
R20955 Vbias Vbias.n102 0.0972718
R20956 Vbias Vbias.n104 0.0972718
R20957 Vbias Vbias.n106 0.0972718
R20958 Vbias Vbias.n108 0.0972718
R20959 Vbias Vbias.n110 0.0972718
R20960 Vbias Vbias.n112 0.0972718
R20961 Vbias Vbias.n114 0.0972718
R20962 Vbias Vbias.n116 0.0972718
R20963 Vbias Vbias.n118 0.0972718
R20964 Vbias Vbias.n120 0.0972718
R20965 Vbias Vbias.n122 0.0972718
R20966 Vbias Vbias.n124 0.0972718
R20967 Vbias Vbias.n126 0.0972718
R20968 Vbias Vbias.n66 0.0972718
R20969 Vbias Vbias.n68 0.0972718
R20970 Vbias Vbias.n70 0.0972718
R20971 Vbias Vbias.n72 0.0972718
R20972 Vbias Vbias.n74 0.0972718
R20973 Vbias Vbias.n76 0.0972718
R20974 Vbias Vbias.n78 0.0972718
R20975 Vbias Vbias.n80 0.0972718
R20976 Vbias Vbias.n82 0.0972718
R20977 Vbias Vbias.n84 0.0972718
R20978 Vbias Vbias.n86 0.0972718
R20979 Vbias Vbias.n88 0.0972718
R20980 Vbias Vbias.n90 0.0972718
R20981 Vbias Vbias.n92 0.0972718
R20982 Vbias Vbias.n94 0.0972718
R20983 Vbias Vbias.n34 0.0972718
R20984 Vbias Vbias.n36 0.0972718
R20985 Vbias Vbias.n38 0.0972718
R20986 Vbias Vbias.n40 0.0972718
R20987 Vbias Vbias.n42 0.0972718
R20988 Vbias Vbias.n44 0.0972718
R20989 Vbias Vbias.n46 0.0972718
R20990 Vbias Vbias.n48 0.0972718
R20991 Vbias Vbias.n50 0.0972718
R20992 Vbias Vbias.n52 0.0972718
R20993 Vbias Vbias.n54 0.0972718
R20994 Vbias Vbias.n56 0.0972718
R20995 Vbias Vbias.n58 0.0972718
R20996 Vbias Vbias.n60 0.0972718
R20997 Vbias Vbias.n62 0.0972718
R20998 Vbias Vbias.n2 0.0972718
R20999 Vbias Vbias.n4 0.0972718
R21000 Vbias Vbias.n6 0.0972718
R21001 Vbias Vbias.n8 0.0972718
R21002 Vbias Vbias.n10 0.0972718
R21003 Vbias Vbias.n12 0.0972718
R21004 Vbias Vbias.n14 0.0972718
R21005 Vbias Vbias.n16 0.0972718
R21006 Vbias Vbias.n18 0.0972718
R21007 Vbias Vbias.n20 0.0972718
R21008 Vbias Vbias.n22 0.0972718
R21009 Vbias Vbias.n24 0.0972718
R21010 Vbias Vbias.n26 0.0972718
R21011 Vbias Vbias.n28 0.0972718
R21012 Vbias Vbias.n30 0.0972718
R21013 Vbias.n509 Vbias 0.0489375
R21014 Vbias.n507 Vbias 0.0489375
R21015 Vbias.n505 Vbias 0.0489375
R21016 Vbias.n503 Vbias 0.0489375
R21017 Vbias.n501 Vbias 0.0489375
R21018 Vbias.n499 Vbias 0.0489375
R21019 Vbias.n497 Vbias 0.0489375
R21020 Vbias.n495 Vbias 0.0489375
R21021 Vbias.n493 Vbias 0.0489375
R21022 Vbias.n491 Vbias 0.0489375
R21023 Vbias.n489 Vbias 0.0489375
R21024 Vbias.n487 Vbias 0.0489375
R21025 Vbias.n485 Vbias 0.0489375
R21026 Vbias.n483 Vbias 0.0489375
R21027 Vbias.n481 Vbias 0.0489375
R21028 Vbias.n480 Vbias 0.0489375
R21029 Vbias.n477 Vbias 0.0489375
R21030 Vbias.n475 Vbias 0.0489375
R21031 Vbias.n473 Vbias 0.0489375
R21032 Vbias.n471 Vbias 0.0489375
R21033 Vbias.n469 Vbias 0.0489375
R21034 Vbias.n467 Vbias 0.0489375
R21035 Vbias.n465 Vbias 0.0489375
R21036 Vbias.n463 Vbias 0.0489375
R21037 Vbias.n461 Vbias 0.0489375
R21038 Vbias.n459 Vbias 0.0489375
R21039 Vbias.n457 Vbias 0.0489375
R21040 Vbias.n455 Vbias 0.0489375
R21041 Vbias.n453 Vbias 0.0489375
R21042 Vbias.n451 Vbias 0.0489375
R21043 Vbias.n449 Vbias 0.0489375
R21044 Vbias.n448 Vbias 0.0489375
R21045 Vbias.n445 Vbias 0.0489375
R21046 Vbias.n443 Vbias 0.0489375
R21047 Vbias.n441 Vbias 0.0489375
R21048 Vbias.n439 Vbias 0.0489375
R21049 Vbias.n437 Vbias 0.0489375
R21050 Vbias.n435 Vbias 0.0489375
R21051 Vbias.n433 Vbias 0.0489375
R21052 Vbias.n431 Vbias 0.0489375
R21053 Vbias.n429 Vbias 0.0489375
R21054 Vbias.n427 Vbias 0.0489375
R21055 Vbias.n425 Vbias 0.0489375
R21056 Vbias.n423 Vbias 0.0489375
R21057 Vbias.n421 Vbias 0.0489375
R21058 Vbias.n419 Vbias 0.0489375
R21059 Vbias.n417 Vbias 0.0489375
R21060 Vbias.n416 Vbias 0.0489375
R21061 Vbias.n413 Vbias 0.0489375
R21062 Vbias.n411 Vbias 0.0489375
R21063 Vbias.n409 Vbias 0.0489375
R21064 Vbias.n407 Vbias 0.0489375
R21065 Vbias.n405 Vbias 0.0489375
R21066 Vbias.n403 Vbias 0.0489375
R21067 Vbias.n401 Vbias 0.0489375
R21068 Vbias.n399 Vbias 0.0489375
R21069 Vbias.n397 Vbias 0.0489375
R21070 Vbias.n395 Vbias 0.0489375
R21071 Vbias.n393 Vbias 0.0489375
R21072 Vbias.n391 Vbias 0.0489375
R21073 Vbias.n389 Vbias 0.0489375
R21074 Vbias.n387 Vbias 0.0489375
R21075 Vbias.n385 Vbias 0.0489375
R21076 Vbias.n384 Vbias 0.0489375
R21077 Vbias.n381 Vbias 0.0489375
R21078 Vbias.n379 Vbias 0.0489375
R21079 Vbias.n377 Vbias 0.0489375
R21080 Vbias.n375 Vbias 0.0489375
R21081 Vbias.n373 Vbias 0.0489375
R21082 Vbias.n371 Vbias 0.0489375
R21083 Vbias.n369 Vbias 0.0489375
R21084 Vbias.n367 Vbias 0.0489375
R21085 Vbias.n365 Vbias 0.0489375
R21086 Vbias.n363 Vbias 0.0489375
R21087 Vbias.n361 Vbias 0.0489375
R21088 Vbias.n359 Vbias 0.0489375
R21089 Vbias.n357 Vbias 0.0489375
R21090 Vbias.n355 Vbias 0.0489375
R21091 Vbias.n353 Vbias 0.0489375
R21092 Vbias.n352 Vbias 0.0489375
R21093 Vbias.n349 Vbias 0.0489375
R21094 Vbias.n347 Vbias 0.0489375
R21095 Vbias.n345 Vbias 0.0489375
R21096 Vbias.n343 Vbias 0.0489375
R21097 Vbias.n341 Vbias 0.0489375
R21098 Vbias.n339 Vbias 0.0489375
R21099 Vbias.n337 Vbias 0.0489375
R21100 Vbias.n335 Vbias 0.0489375
R21101 Vbias.n333 Vbias 0.0489375
R21102 Vbias.n331 Vbias 0.0489375
R21103 Vbias.n329 Vbias 0.0489375
R21104 Vbias.n327 Vbias 0.0489375
R21105 Vbias.n325 Vbias 0.0489375
R21106 Vbias.n323 Vbias 0.0489375
R21107 Vbias.n321 Vbias 0.0489375
R21108 Vbias.n320 Vbias 0.0489375
R21109 Vbias.n317 Vbias 0.0489375
R21110 Vbias.n315 Vbias 0.0489375
R21111 Vbias.n313 Vbias 0.0489375
R21112 Vbias.n311 Vbias 0.0489375
R21113 Vbias.n309 Vbias 0.0489375
R21114 Vbias.n307 Vbias 0.0489375
R21115 Vbias.n305 Vbias 0.0489375
R21116 Vbias.n303 Vbias 0.0489375
R21117 Vbias.n301 Vbias 0.0489375
R21118 Vbias.n299 Vbias 0.0489375
R21119 Vbias.n297 Vbias 0.0489375
R21120 Vbias.n295 Vbias 0.0489375
R21121 Vbias.n293 Vbias 0.0489375
R21122 Vbias.n291 Vbias 0.0489375
R21123 Vbias.n289 Vbias 0.0489375
R21124 Vbias.n288 Vbias 0.0489375
R21125 Vbias.n285 Vbias 0.0489375
R21126 Vbias.n283 Vbias 0.0489375
R21127 Vbias.n281 Vbias 0.0489375
R21128 Vbias.n279 Vbias 0.0489375
R21129 Vbias.n277 Vbias 0.0489375
R21130 Vbias.n275 Vbias 0.0489375
R21131 Vbias.n273 Vbias 0.0489375
R21132 Vbias.n271 Vbias 0.0489375
R21133 Vbias.n269 Vbias 0.0489375
R21134 Vbias.n267 Vbias 0.0489375
R21135 Vbias.n265 Vbias 0.0489375
R21136 Vbias.n263 Vbias 0.0489375
R21137 Vbias.n261 Vbias 0.0489375
R21138 Vbias.n259 Vbias 0.0489375
R21139 Vbias.n257 Vbias 0.0489375
R21140 Vbias.n256 Vbias 0.0489375
R21141 Vbias.n253 Vbias 0.0489375
R21142 Vbias.n251 Vbias 0.0489375
R21143 Vbias.n249 Vbias 0.0489375
R21144 Vbias.n247 Vbias 0.0489375
R21145 Vbias.n245 Vbias 0.0489375
R21146 Vbias.n243 Vbias 0.0489375
R21147 Vbias.n241 Vbias 0.0489375
R21148 Vbias.n239 Vbias 0.0489375
R21149 Vbias.n237 Vbias 0.0489375
R21150 Vbias.n235 Vbias 0.0489375
R21151 Vbias.n233 Vbias 0.0489375
R21152 Vbias.n231 Vbias 0.0489375
R21153 Vbias.n229 Vbias 0.0489375
R21154 Vbias.n227 Vbias 0.0489375
R21155 Vbias.n225 Vbias 0.0489375
R21156 Vbias.n224 Vbias 0.0489375
R21157 Vbias.n221 Vbias 0.0489375
R21158 Vbias.n219 Vbias 0.0489375
R21159 Vbias.n217 Vbias 0.0489375
R21160 Vbias.n215 Vbias 0.0489375
R21161 Vbias.n213 Vbias 0.0489375
R21162 Vbias.n211 Vbias 0.0489375
R21163 Vbias.n209 Vbias 0.0489375
R21164 Vbias.n207 Vbias 0.0489375
R21165 Vbias.n205 Vbias 0.0489375
R21166 Vbias.n203 Vbias 0.0489375
R21167 Vbias.n201 Vbias 0.0489375
R21168 Vbias.n199 Vbias 0.0489375
R21169 Vbias.n197 Vbias 0.0489375
R21170 Vbias.n195 Vbias 0.0489375
R21171 Vbias.n193 Vbias 0.0489375
R21172 Vbias.n192 Vbias 0.0489375
R21173 Vbias.n189 Vbias 0.0489375
R21174 Vbias.n187 Vbias 0.0489375
R21175 Vbias.n185 Vbias 0.0489375
R21176 Vbias.n183 Vbias 0.0489375
R21177 Vbias.n181 Vbias 0.0489375
R21178 Vbias.n179 Vbias 0.0489375
R21179 Vbias.n177 Vbias 0.0489375
R21180 Vbias.n175 Vbias 0.0489375
R21181 Vbias.n173 Vbias 0.0489375
R21182 Vbias.n171 Vbias 0.0489375
R21183 Vbias.n169 Vbias 0.0489375
R21184 Vbias.n167 Vbias 0.0489375
R21185 Vbias.n165 Vbias 0.0489375
R21186 Vbias.n163 Vbias 0.0489375
R21187 Vbias.n161 Vbias 0.0489375
R21188 Vbias.n160 Vbias 0.0489375
R21189 Vbias.n157 Vbias 0.0489375
R21190 Vbias.n155 Vbias 0.0489375
R21191 Vbias.n153 Vbias 0.0489375
R21192 Vbias.n151 Vbias 0.0489375
R21193 Vbias.n149 Vbias 0.0489375
R21194 Vbias.n147 Vbias 0.0489375
R21195 Vbias.n145 Vbias 0.0489375
R21196 Vbias.n143 Vbias 0.0489375
R21197 Vbias.n141 Vbias 0.0489375
R21198 Vbias.n139 Vbias 0.0489375
R21199 Vbias.n137 Vbias 0.0489375
R21200 Vbias.n135 Vbias 0.0489375
R21201 Vbias.n133 Vbias 0.0489375
R21202 Vbias.n131 Vbias 0.0489375
R21203 Vbias.n129 Vbias 0.0489375
R21204 Vbias.n128 Vbias 0.0489375
R21205 Vbias.n125 Vbias 0.0489375
R21206 Vbias.n123 Vbias 0.0489375
R21207 Vbias.n121 Vbias 0.0489375
R21208 Vbias.n119 Vbias 0.0489375
R21209 Vbias.n117 Vbias 0.0489375
R21210 Vbias.n115 Vbias 0.0489375
R21211 Vbias.n113 Vbias 0.0489375
R21212 Vbias.n111 Vbias 0.0489375
R21213 Vbias.n109 Vbias 0.0489375
R21214 Vbias.n107 Vbias 0.0489375
R21215 Vbias.n105 Vbias 0.0489375
R21216 Vbias.n103 Vbias 0.0489375
R21217 Vbias.n101 Vbias 0.0489375
R21218 Vbias.n99 Vbias 0.0489375
R21219 Vbias.n97 Vbias 0.0489375
R21220 Vbias.n96 Vbias 0.0489375
R21221 Vbias.n93 Vbias 0.0489375
R21222 Vbias.n91 Vbias 0.0489375
R21223 Vbias.n89 Vbias 0.0489375
R21224 Vbias.n87 Vbias 0.0489375
R21225 Vbias.n85 Vbias 0.0489375
R21226 Vbias.n83 Vbias 0.0489375
R21227 Vbias.n81 Vbias 0.0489375
R21228 Vbias.n79 Vbias 0.0489375
R21229 Vbias.n77 Vbias 0.0489375
R21230 Vbias.n75 Vbias 0.0489375
R21231 Vbias.n73 Vbias 0.0489375
R21232 Vbias.n71 Vbias 0.0489375
R21233 Vbias.n69 Vbias 0.0489375
R21234 Vbias.n67 Vbias 0.0489375
R21235 Vbias.n65 Vbias 0.0489375
R21236 Vbias.n64 Vbias 0.0489375
R21237 Vbias.n61 Vbias 0.0489375
R21238 Vbias.n59 Vbias 0.0489375
R21239 Vbias.n57 Vbias 0.0489375
R21240 Vbias.n55 Vbias 0.0489375
R21241 Vbias.n53 Vbias 0.0489375
R21242 Vbias.n51 Vbias 0.0489375
R21243 Vbias.n49 Vbias 0.0489375
R21244 Vbias.n47 Vbias 0.0489375
R21245 Vbias.n45 Vbias 0.0489375
R21246 Vbias.n43 Vbias 0.0489375
R21247 Vbias.n41 Vbias 0.0489375
R21248 Vbias.n39 Vbias 0.0489375
R21249 Vbias.n37 Vbias 0.0489375
R21250 Vbias.n35 Vbias 0.0489375
R21251 Vbias.n33 Vbias 0.0489375
R21252 Vbias.n32 Vbias 0.0489375
R21253 Vbias.n29 Vbias 0.0489375
R21254 Vbias.n27 Vbias 0.0489375
R21255 Vbias.n25 Vbias 0.0489375
R21256 Vbias.n23 Vbias 0.0489375
R21257 Vbias.n21 Vbias 0.0489375
R21258 Vbias.n19 Vbias 0.0489375
R21259 Vbias.n17 Vbias 0.0489375
R21260 Vbias.n15 Vbias 0.0489375
R21261 Vbias.n13 Vbias 0.0489375
R21262 Vbias.n11 Vbias 0.0489375
R21263 Vbias.n9 Vbias 0.0489375
R21264 Vbias.n7 Vbias 0.0489375
R21265 Vbias.n5 Vbias 0.0489375
R21266 Vbias.n3 Vbias 0.0489375
R21267 Vbias.n1 Vbias 0.0489375
R21268 Vbias.n0 Vbias 0.0489375
R21269 XThC.Tn[1].n2 XThC.Tn[1].n1 332.332
R21270 XThC.Tn[1].n2 XThC.Tn[1].n0 296.493
R21271 XThC.Tn[1].n71 XThC.Tn[1].n69 161.365
R21272 XThC.Tn[1].n67 XThC.Tn[1].n65 161.365
R21273 XThC.Tn[1].n63 XThC.Tn[1].n61 161.365
R21274 XThC.Tn[1].n59 XThC.Tn[1].n57 161.365
R21275 XThC.Tn[1].n55 XThC.Tn[1].n53 161.365
R21276 XThC.Tn[1].n51 XThC.Tn[1].n49 161.365
R21277 XThC.Tn[1].n47 XThC.Tn[1].n45 161.365
R21278 XThC.Tn[1].n43 XThC.Tn[1].n41 161.365
R21279 XThC.Tn[1].n39 XThC.Tn[1].n37 161.365
R21280 XThC.Tn[1].n35 XThC.Tn[1].n33 161.365
R21281 XThC.Tn[1].n31 XThC.Tn[1].n29 161.365
R21282 XThC.Tn[1].n27 XThC.Tn[1].n25 161.365
R21283 XThC.Tn[1].n23 XThC.Tn[1].n21 161.365
R21284 XThC.Tn[1].n19 XThC.Tn[1].n17 161.365
R21285 XThC.Tn[1].n15 XThC.Tn[1].n13 161.365
R21286 XThC.Tn[1].n12 XThC.Tn[1].n10 161.365
R21287 XThC.Tn[1].n69 XThC.Tn[1].t35 161.202
R21288 XThC.Tn[1].n65 XThC.Tn[1].t25 161.202
R21289 XThC.Tn[1].n61 XThC.Tn[1].t12 161.202
R21290 XThC.Tn[1].n57 XThC.Tn[1].t41 161.202
R21291 XThC.Tn[1].n53 XThC.Tn[1].t33 161.202
R21292 XThC.Tn[1].n49 XThC.Tn[1].t20 161.202
R21293 XThC.Tn[1].n45 XThC.Tn[1].t19 161.202
R21294 XThC.Tn[1].n41 XThC.Tn[1].t32 161.202
R21295 XThC.Tn[1].n37 XThC.Tn[1].t30 161.202
R21296 XThC.Tn[1].n33 XThC.Tn[1].t21 161.202
R21297 XThC.Tn[1].n29 XThC.Tn[1].t40 161.202
R21298 XThC.Tn[1].n25 XThC.Tn[1].t39 161.202
R21299 XThC.Tn[1].n21 XThC.Tn[1].t18 161.202
R21300 XThC.Tn[1].n17 XThC.Tn[1].t16 161.202
R21301 XThC.Tn[1].n13 XThC.Tn[1].t14 161.202
R21302 XThC.Tn[1].n10 XThC.Tn[1].t29 161.202
R21303 XThC.Tn[1].n69 XThC.Tn[1].t38 145.137
R21304 XThC.Tn[1].n65 XThC.Tn[1].t28 145.137
R21305 XThC.Tn[1].n61 XThC.Tn[1].t15 145.137
R21306 XThC.Tn[1].n57 XThC.Tn[1].t13 145.137
R21307 XThC.Tn[1].n53 XThC.Tn[1].t37 145.137
R21308 XThC.Tn[1].n49 XThC.Tn[1].t26 145.137
R21309 XThC.Tn[1].n45 XThC.Tn[1].t24 145.137
R21310 XThC.Tn[1].n41 XThC.Tn[1].t36 145.137
R21311 XThC.Tn[1].n37 XThC.Tn[1].t34 145.137
R21312 XThC.Tn[1].n33 XThC.Tn[1].t27 145.137
R21313 XThC.Tn[1].n29 XThC.Tn[1].t43 145.137
R21314 XThC.Tn[1].n25 XThC.Tn[1].t42 145.137
R21315 XThC.Tn[1].n21 XThC.Tn[1].t23 145.137
R21316 XThC.Tn[1].n17 XThC.Tn[1].t22 145.137
R21317 XThC.Tn[1].n13 XThC.Tn[1].t17 145.137
R21318 XThC.Tn[1].n10 XThC.Tn[1].t31 145.137
R21319 XThC.Tn[1].n5 XThC.Tn[1].n3 135.249
R21320 XThC.Tn[1].n5 XThC.Tn[1].n4 98.981
R21321 XThC.Tn[1].n7 XThC.Tn[1].n6 98.981
R21322 XThC.Tn[1].n9 XThC.Tn[1].n8 98.981
R21323 XThC.Tn[1].n7 XThC.Tn[1].n5 36.2672
R21324 XThC.Tn[1].n9 XThC.Tn[1].n7 36.2672
R21325 XThC.Tn[1].n74 XThC.Tn[1].n9 32.6405
R21326 XThC.Tn[1].n1 XThC.Tn[1].t1 26.5955
R21327 XThC.Tn[1].n1 XThC.Tn[1].t0 26.5955
R21328 XThC.Tn[1].n0 XThC.Tn[1].t3 26.5955
R21329 XThC.Tn[1].n0 XThC.Tn[1].t2 26.5955
R21330 XThC.Tn[1].n3 XThC.Tn[1].t11 24.9236
R21331 XThC.Tn[1].n3 XThC.Tn[1].t10 24.9236
R21332 XThC.Tn[1].n4 XThC.Tn[1].t9 24.9236
R21333 XThC.Tn[1].n4 XThC.Tn[1].t8 24.9236
R21334 XThC.Tn[1].n6 XThC.Tn[1].t7 24.9236
R21335 XThC.Tn[1].n6 XThC.Tn[1].t6 24.9236
R21336 XThC.Tn[1].n8 XThC.Tn[1].t5 24.9236
R21337 XThC.Tn[1].n8 XThC.Tn[1].t4 24.9236
R21338 XThC.Tn[1] XThC.Tn[1].n2 23.3605
R21339 XThC.Tn[1] XThC.Tn[1].n12 8.0245
R21340 XThC.Tn[1].n72 XThC.Tn[1].n71 7.9105
R21341 XThC.Tn[1].n68 XThC.Tn[1].n67 7.9105
R21342 XThC.Tn[1].n64 XThC.Tn[1].n63 7.9105
R21343 XThC.Tn[1].n60 XThC.Tn[1].n59 7.9105
R21344 XThC.Tn[1].n56 XThC.Tn[1].n55 7.9105
R21345 XThC.Tn[1].n52 XThC.Tn[1].n51 7.9105
R21346 XThC.Tn[1].n48 XThC.Tn[1].n47 7.9105
R21347 XThC.Tn[1].n44 XThC.Tn[1].n43 7.9105
R21348 XThC.Tn[1].n40 XThC.Tn[1].n39 7.9105
R21349 XThC.Tn[1].n36 XThC.Tn[1].n35 7.9105
R21350 XThC.Tn[1].n32 XThC.Tn[1].n31 7.9105
R21351 XThC.Tn[1].n28 XThC.Tn[1].n27 7.9105
R21352 XThC.Tn[1].n24 XThC.Tn[1].n23 7.9105
R21353 XThC.Tn[1].n20 XThC.Tn[1].n19 7.9105
R21354 XThC.Tn[1].n16 XThC.Tn[1].n15 7.9105
R21355 XThC.Tn[1] XThC.Tn[1].n74 6.7205
R21356 XThC.Tn[1].n73 XThC.Tn[1] 6.08068
R21357 XThC.Tn[1].n74 XThC.Tn[1].n73 4.65249
R21358 XThC.Tn[1].n73 XThC.Tn[1] 1.8942
R21359 XThC.Tn[1].n16 XThC.Tn[1] 0.235138
R21360 XThC.Tn[1].n20 XThC.Tn[1] 0.235138
R21361 XThC.Tn[1].n24 XThC.Tn[1] 0.235138
R21362 XThC.Tn[1].n28 XThC.Tn[1] 0.235138
R21363 XThC.Tn[1].n32 XThC.Tn[1] 0.235138
R21364 XThC.Tn[1].n36 XThC.Tn[1] 0.235138
R21365 XThC.Tn[1].n40 XThC.Tn[1] 0.235138
R21366 XThC.Tn[1].n44 XThC.Tn[1] 0.235138
R21367 XThC.Tn[1].n48 XThC.Tn[1] 0.235138
R21368 XThC.Tn[1].n52 XThC.Tn[1] 0.235138
R21369 XThC.Tn[1].n56 XThC.Tn[1] 0.235138
R21370 XThC.Tn[1].n60 XThC.Tn[1] 0.235138
R21371 XThC.Tn[1].n64 XThC.Tn[1] 0.235138
R21372 XThC.Tn[1].n68 XThC.Tn[1] 0.235138
R21373 XThC.Tn[1].n72 XThC.Tn[1] 0.235138
R21374 XThC.Tn[1] XThC.Tn[1].n16 0.114505
R21375 XThC.Tn[1] XThC.Tn[1].n20 0.114505
R21376 XThC.Tn[1] XThC.Tn[1].n24 0.114505
R21377 XThC.Tn[1] XThC.Tn[1].n28 0.114505
R21378 XThC.Tn[1] XThC.Tn[1].n32 0.114505
R21379 XThC.Tn[1] XThC.Tn[1].n36 0.114505
R21380 XThC.Tn[1] XThC.Tn[1].n40 0.114505
R21381 XThC.Tn[1] XThC.Tn[1].n44 0.114505
R21382 XThC.Tn[1] XThC.Tn[1].n48 0.114505
R21383 XThC.Tn[1] XThC.Tn[1].n52 0.114505
R21384 XThC.Tn[1] XThC.Tn[1].n56 0.114505
R21385 XThC.Tn[1] XThC.Tn[1].n60 0.114505
R21386 XThC.Tn[1] XThC.Tn[1].n64 0.114505
R21387 XThC.Tn[1] XThC.Tn[1].n68 0.114505
R21388 XThC.Tn[1] XThC.Tn[1].n72 0.114505
R21389 XThC.Tn[1].n71 XThC.Tn[1].n70 0.0599512
R21390 XThC.Tn[1].n67 XThC.Tn[1].n66 0.0599512
R21391 XThC.Tn[1].n63 XThC.Tn[1].n62 0.0599512
R21392 XThC.Tn[1].n59 XThC.Tn[1].n58 0.0599512
R21393 XThC.Tn[1].n55 XThC.Tn[1].n54 0.0599512
R21394 XThC.Tn[1].n51 XThC.Tn[1].n50 0.0599512
R21395 XThC.Tn[1].n47 XThC.Tn[1].n46 0.0599512
R21396 XThC.Tn[1].n43 XThC.Tn[1].n42 0.0599512
R21397 XThC.Tn[1].n39 XThC.Tn[1].n38 0.0599512
R21398 XThC.Tn[1].n35 XThC.Tn[1].n34 0.0599512
R21399 XThC.Tn[1].n31 XThC.Tn[1].n30 0.0599512
R21400 XThC.Tn[1].n27 XThC.Tn[1].n26 0.0599512
R21401 XThC.Tn[1].n23 XThC.Tn[1].n22 0.0599512
R21402 XThC.Tn[1].n19 XThC.Tn[1].n18 0.0599512
R21403 XThC.Tn[1].n15 XThC.Tn[1].n14 0.0599512
R21404 XThC.Tn[1].n12 XThC.Tn[1].n11 0.0599512
R21405 XThC.Tn[1].n70 XThC.Tn[1] 0.0469286
R21406 XThC.Tn[1].n66 XThC.Tn[1] 0.0469286
R21407 XThC.Tn[1].n62 XThC.Tn[1] 0.0469286
R21408 XThC.Tn[1].n58 XThC.Tn[1] 0.0469286
R21409 XThC.Tn[1].n54 XThC.Tn[1] 0.0469286
R21410 XThC.Tn[1].n50 XThC.Tn[1] 0.0469286
R21411 XThC.Tn[1].n46 XThC.Tn[1] 0.0469286
R21412 XThC.Tn[1].n42 XThC.Tn[1] 0.0469286
R21413 XThC.Tn[1].n38 XThC.Tn[1] 0.0469286
R21414 XThC.Tn[1].n34 XThC.Tn[1] 0.0469286
R21415 XThC.Tn[1].n30 XThC.Tn[1] 0.0469286
R21416 XThC.Tn[1].n26 XThC.Tn[1] 0.0469286
R21417 XThC.Tn[1].n22 XThC.Tn[1] 0.0469286
R21418 XThC.Tn[1].n18 XThC.Tn[1] 0.0469286
R21419 XThC.Tn[1].n14 XThC.Tn[1] 0.0469286
R21420 XThC.Tn[1].n11 XThC.Tn[1] 0.0469286
R21421 XThC.Tn[1].n70 XThC.Tn[1] 0.0401341
R21422 XThC.Tn[1].n66 XThC.Tn[1] 0.0401341
R21423 XThC.Tn[1].n62 XThC.Tn[1] 0.0401341
R21424 XThC.Tn[1].n58 XThC.Tn[1] 0.0401341
R21425 XThC.Tn[1].n54 XThC.Tn[1] 0.0401341
R21426 XThC.Tn[1].n50 XThC.Tn[1] 0.0401341
R21427 XThC.Tn[1].n46 XThC.Tn[1] 0.0401341
R21428 XThC.Tn[1].n42 XThC.Tn[1] 0.0401341
R21429 XThC.Tn[1].n38 XThC.Tn[1] 0.0401341
R21430 XThC.Tn[1].n34 XThC.Tn[1] 0.0401341
R21431 XThC.Tn[1].n30 XThC.Tn[1] 0.0401341
R21432 XThC.Tn[1].n26 XThC.Tn[1] 0.0401341
R21433 XThC.Tn[1].n22 XThC.Tn[1] 0.0401341
R21434 XThC.Tn[1].n18 XThC.Tn[1] 0.0401341
R21435 XThC.Tn[1].n14 XThC.Tn[1] 0.0401341
R21436 XThC.Tn[1].n11 XThC.Tn[1] 0.0401341
R21437 XThC.Tn[3].n2 XThC.Tn[3].n1 332.332
R21438 XThC.Tn[3].n2 XThC.Tn[3].n0 296.493
R21439 XThC.Tn[3].n71 XThC.Tn[3].n69 161.365
R21440 XThC.Tn[3].n67 XThC.Tn[3].n65 161.365
R21441 XThC.Tn[3].n63 XThC.Tn[3].n61 161.365
R21442 XThC.Tn[3].n59 XThC.Tn[3].n57 161.365
R21443 XThC.Tn[3].n55 XThC.Tn[3].n53 161.365
R21444 XThC.Tn[3].n51 XThC.Tn[3].n49 161.365
R21445 XThC.Tn[3].n47 XThC.Tn[3].n45 161.365
R21446 XThC.Tn[3].n43 XThC.Tn[3].n41 161.365
R21447 XThC.Tn[3].n39 XThC.Tn[3].n37 161.365
R21448 XThC.Tn[3].n35 XThC.Tn[3].n33 161.365
R21449 XThC.Tn[3].n31 XThC.Tn[3].n29 161.365
R21450 XThC.Tn[3].n27 XThC.Tn[3].n25 161.365
R21451 XThC.Tn[3].n23 XThC.Tn[3].n21 161.365
R21452 XThC.Tn[3].n19 XThC.Tn[3].n17 161.365
R21453 XThC.Tn[3].n15 XThC.Tn[3].n13 161.365
R21454 XThC.Tn[3].n12 XThC.Tn[3].n10 161.365
R21455 XThC.Tn[3].n69 XThC.Tn[3].t16 161.202
R21456 XThC.Tn[3].n65 XThC.Tn[3].t38 161.202
R21457 XThC.Tn[3].n61 XThC.Tn[3].t25 161.202
R21458 XThC.Tn[3].n57 XThC.Tn[3].t22 161.202
R21459 XThC.Tn[3].n53 XThC.Tn[3].t14 161.202
R21460 XThC.Tn[3].n49 XThC.Tn[3].t33 161.202
R21461 XThC.Tn[3].n45 XThC.Tn[3].t32 161.202
R21462 XThC.Tn[3].n41 XThC.Tn[3].t13 161.202
R21463 XThC.Tn[3].n37 XThC.Tn[3].t43 161.202
R21464 XThC.Tn[3].n33 XThC.Tn[3].t34 161.202
R21465 XThC.Tn[3].n29 XThC.Tn[3].t21 161.202
R21466 XThC.Tn[3].n25 XThC.Tn[3].t20 161.202
R21467 XThC.Tn[3].n21 XThC.Tn[3].t31 161.202
R21468 XThC.Tn[3].n17 XThC.Tn[3].t29 161.202
R21469 XThC.Tn[3].n13 XThC.Tn[3].t27 161.202
R21470 XThC.Tn[3].n10 XThC.Tn[3].t42 161.202
R21471 XThC.Tn[3].n69 XThC.Tn[3].t19 145.137
R21472 XThC.Tn[3].n65 XThC.Tn[3].t41 145.137
R21473 XThC.Tn[3].n61 XThC.Tn[3].t28 145.137
R21474 XThC.Tn[3].n57 XThC.Tn[3].t26 145.137
R21475 XThC.Tn[3].n53 XThC.Tn[3].t18 145.137
R21476 XThC.Tn[3].n49 XThC.Tn[3].t39 145.137
R21477 XThC.Tn[3].n45 XThC.Tn[3].t37 145.137
R21478 XThC.Tn[3].n41 XThC.Tn[3].t17 145.137
R21479 XThC.Tn[3].n37 XThC.Tn[3].t15 145.137
R21480 XThC.Tn[3].n33 XThC.Tn[3].t40 145.137
R21481 XThC.Tn[3].n29 XThC.Tn[3].t24 145.137
R21482 XThC.Tn[3].n25 XThC.Tn[3].t23 145.137
R21483 XThC.Tn[3].n21 XThC.Tn[3].t36 145.137
R21484 XThC.Tn[3].n17 XThC.Tn[3].t35 145.137
R21485 XThC.Tn[3].n13 XThC.Tn[3].t30 145.137
R21486 XThC.Tn[3].n10 XThC.Tn[3].t12 145.137
R21487 XThC.Tn[3].n6 XThC.Tn[3].n4 135.249
R21488 XThC.Tn[3].n9 XThC.Tn[3].n3 98.981
R21489 XThC.Tn[3].n6 XThC.Tn[3].n5 98.981
R21490 XThC.Tn[3].n8 XThC.Tn[3].n7 98.981
R21491 XThC.Tn[3].n8 XThC.Tn[3].n6 36.2672
R21492 XThC.Tn[3].n9 XThC.Tn[3].n8 36.2672
R21493 XThC.Tn[3].n74 XThC.Tn[3].n9 32.6405
R21494 XThC.Tn[3].n1 XThC.Tn[3].t7 26.5955
R21495 XThC.Tn[3].n1 XThC.Tn[3].t6 26.5955
R21496 XThC.Tn[3].n0 XThC.Tn[3].t5 26.5955
R21497 XThC.Tn[3].n0 XThC.Tn[3].t4 26.5955
R21498 XThC.Tn[3].n3 XThC.Tn[3].t1 24.9236
R21499 XThC.Tn[3].n3 XThC.Tn[3].t0 24.9236
R21500 XThC.Tn[3].n4 XThC.Tn[3].t11 24.9236
R21501 XThC.Tn[3].n4 XThC.Tn[3].t10 24.9236
R21502 XThC.Tn[3].n5 XThC.Tn[3].t9 24.9236
R21503 XThC.Tn[3].n5 XThC.Tn[3].t8 24.9236
R21504 XThC.Tn[3].n7 XThC.Tn[3].t3 24.9236
R21505 XThC.Tn[3].n7 XThC.Tn[3].t2 24.9236
R21506 XThC.Tn[3] XThC.Tn[3].n2 23.3605
R21507 XThC.Tn[3] XThC.Tn[3].n12 8.0245
R21508 XThC.Tn[3].n72 XThC.Tn[3].n71 7.9105
R21509 XThC.Tn[3].n68 XThC.Tn[3].n67 7.9105
R21510 XThC.Tn[3].n64 XThC.Tn[3].n63 7.9105
R21511 XThC.Tn[3].n60 XThC.Tn[3].n59 7.9105
R21512 XThC.Tn[3].n56 XThC.Tn[3].n55 7.9105
R21513 XThC.Tn[3].n52 XThC.Tn[3].n51 7.9105
R21514 XThC.Tn[3].n48 XThC.Tn[3].n47 7.9105
R21515 XThC.Tn[3].n44 XThC.Tn[3].n43 7.9105
R21516 XThC.Tn[3].n40 XThC.Tn[3].n39 7.9105
R21517 XThC.Tn[3].n36 XThC.Tn[3].n35 7.9105
R21518 XThC.Tn[3].n32 XThC.Tn[3].n31 7.9105
R21519 XThC.Tn[3].n28 XThC.Tn[3].n27 7.9105
R21520 XThC.Tn[3].n24 XThC.Tn[3].n23 7.9105
R21521 XThC.Tn[3].n20 XThC.Tn[3].n19 7.9105
R21522 XThC.Tn[3].n16 XThC.Tn[3].n15 7.9105
R21523 XThC.Tn[3].n73 XThC.Tn[3] 7.48718
R21524 XThC.Tn[3] XThC.Tn[3].n74 6.7205
R21525 XThC.Tn[3].n74 XThC.Tn[3].n73 5.06464
R21526 XThC.Tn[3].n73 XThC.Tn[3] 1.18175
R21527 XThC.Tn[3].n16 XThC.Tn[3] 0.235138
R21528 XThC.Tn[3].n20 XThC.Tn[3] 0.235138
R21529 XThC.Tn[3].n24 XThC.Tn[3] 0.235138
R21530 XThC.Tn[3].n28 XThC.Tn[3] 0.235138
R21531 XThC.Tn[3].n32 XThC.Tn[3] 0.235138
R21532 XThC.Tn[3].n36 XThC.Tn[3] 0.235138
R21533 XThC.Tn[3].n40 XThC.Tn[3] 0.235138
R21534 XThC.Tn[3].n44 XThC.Tn[3] 0.235138
R21535 XThC.Tn[3].n48 XThC.Tn[3] 0.235138
R21536 XThC.Tn[3].n52 XThC.Tn[3] 0.235138
R21537 XThC.Tn[3].n56 XThC.Tn[3] 0.235138
R21538 XThC.Tn[3].n60 XThC.Tn[3] 0.235138
R21539 XThC.Tn[3].n64 XThC.Tn[3] 0.235138
R21540 XThC.Tn[3].n68 XThC.Tn[3] 0.235138
R21541 XThC.Tn[3].n72 XThC.Tn[3] 0.235138
R21542 XThC.Tn[3] XThC.Tn[3].n16 0.114505
R21543 XThC.Tn[3] XThC.Tn[3].n20 0.114505
R21544 XThC.Tn[3] XThC.Tn[3].n24 0.114505
R21545 XThC.Tn[3] XThC.Tn[3].n28 0.114505
R21546 XThC.Tn[3] XThC.Tn[3].n32 0.114505
R21547 XThC.Tn[3] XThC.Tn[3].n36 0.114505
R21548 XThC.Tn[3] XThC.Tn[3].n40 0.114505
R21549 XThC.Tn[3] XThC.Tn[3].n44 0.114505
R21550 XThC.Tn[3] XThC.Tn[3].n48 0.114505
R21551 XThC.Tn[3] XThC.Tn[3].n52 0.114505
R21552 XThC.Tn[3] XThC.Tn[3].n56 0.114505
R21553 XThC.Tn[3] XThC.Tn[3].n60 0.114505
R21554 XThC.Tn[3] XThC.Tn[3].n64 0.114505
R21555 XThC.Tn[3] XThC.Tn[3].n68 0.114505
R21556 XThC.Tn[3] XThC.Tn[3].n72 0.114505
R21557 XThC.Tn[3].n71 XThC.Tn[3].n70 0.0599512
R21558 XThC.Tn[3].n67 XThC.Tn[3].n66 0.0599512
R21559 XThC.Tn[3].n63 XThC.Tn[3].n62 0.0599512
R21560 XThC.Tn[3].n59 XThC.Tn[3].n58 0.0599512
R21561 XThC.Tn[3].n55 XThC.Tn[3].n54 0.0599512
R21562 XThC.Tn[3].n51 XThC.Tn[3].n50 0.0599512
R21563 XThC.Tn[3].n47 XThC.Tn[3].n46 0.0599512
R21564 XThC.Tn[3].n43 XThC.Tn[3].n42 0.0599512
R21565 XThC.Tn[3].n39 XThC.Tn[3].n38 0.0599512
R21566 XThC.Tn[3].n35 XThC.Tn[3].n34 0.0599512
R21567 XThC.Tn[3].n31 XThC.Tn[3].n30 0.0599512
R21568 XThC.Tn[3].n27 XThC.Tn[3].n26 0.0599512
R21569 XThC.Tn[3].n23 XThC.Tn[3].n22 0.0599512
R21570 XThC.Tn[3].n19 XThC.Tn[3].n18 0.0599512
R21571 XThC.Tn[3].n15 XThC.Tn[3].n14 0.0599512
R21572 XThC.Tn[3].n12 XThC.Tn[3].n11 0.0599512
R21573 XThC.Tn[3].n70 XThC.Tn[3] 0.0469286
R21574 XThC.Tn[3].n66 XThC.Tn[3] 0.0469286
R21575 XThC.Tn[3].n62 XThC.Tn[3] 0.0469286
R21576 XThC.Tn[3].n58 XThC.Tn[3] 0.0469286
R21577 XThC.Tn[3].n54 XThC.Tn[3] 0.0469286
R21578 XThC.Tn[3].n50 XThC.Tn[3] 0.0469286
R21579 XThC.Tn[3].n46 XThC.Tn[3] 0.0469286
R21580 XThC.Tn[3].n42 XThC.Tn[3] 0.0469286
R21581 XThC.Tn[3].n38 XThC.Tn[3] 0.0469286
R21582 XThC.Tn[3].n34 XThC.Tn[3] 0.0469286
R21583 XThC.Tn[3].n30 XThC.Tn[3] 0.0469286
R21584 XThC.Tn[3].n26 XThC.Tn[3] 0.0469286
R21585 XThC.Tn[3].n22 XThC.Tn[3] 0.0469286
R21586 XThC.Tn[3].n18 XThC.Tn[3] 0.0469286
R21587 XThC.Tn[3].n14 XThC.Tn[3] 0.0469286
R21588 XThC.Tn[3].n11 XThC.Tn[3] 0.0469286
R21589 XThC.Tn[3].n70 XThC.Tn[3] 0.0401341
R21590 XThC.Tn[3].n66 XThC.Tn[3] 0.0401341
R21591 XThC.Tn[3].n62 XThC.Tn[3] 0.0401341
R21592 XThC.Tn[3].n58 XThC.Tn[3] 0.0401341
R21593 XThC.Tn[3].n54 XThC.Tn[3] 0.0401341
R21594 XThC.Tn[3].n50 XThC.Tn[3] 0.0401341
R21595 XThC.Tn[3].n46 XThC.Tn[3] 0.0401341
R21596 XThC.Tn[3].n42 XThC.Tn[3] 0.0401341
R21597 XThC.Tn[3].n38 XThC.Tn[3] 0.0401341
R21598 XThC.Tn[3].n34 XThC.Tn[3] 0.0401341
R21599 XThC.Tn[3].n30 XThC.Tn[3] 0.0401341
R21600 XThC.Tn[3].n26 XThC.Tn[3] 0.0401341
R21601 XThC.Tn[3].n22 XThC.Tn[3] 0.0401341
R21602 XThC.Tn[3].n18 XThC.Tn[3] 0.0401341
R21603 XThC.Tn[3].n14 XThC.Tn[3] 0.0401341
R21604 XThC.Tn[3].n11 XThC.Tn[3] 0.0401341
R21605 XThR.Tn[10].n87 XThR.Tn[10].n86 256.103
R21606 XThR.Tn[10].n2 XThR.Tn[10].n0 243.68
R21607 XThR.Tn[10].n5 XThR.Tn[10].n3 241.847
R21608 XThR.Tn[10].n2 XThR.Tn[10].n1 205.28
R21609 XThR.Tn[10].n87 XThR.Tn[10].n85 202.095
R21610 XThR.Tn[10].n5 XThR.Tn[10].n4 185
R21611 XThR.Tn[10] XThR.Tn[10].n78 161.363
R21612 XThR.Tn[10] XThR.Tn[10].n73 161.363
R21613 XThR.Tn[10] XThR.Tn[10].n68 161.363
R21614 XThR.Tn[10] XThR.Tn[10].n63 161.363
R21615 XThR.Tn[10] XThR.Tn[10].n58 161.363
R21616 XThR.Tn[10] XThR.Tn[10].n53 161.363
R21617 XThR.Tn[10] XThR.Tn[10].n48 161.363
R21618 XThR.Tn[10] XThR.Tn[10].n43 161.363
R21619 XThR.Tn[10] XThR.Tn[10].n38 161.363
R21620 XThR.Tn[10] XThR.Tn[10].n33 161.363
R21621 XThR.Tn[10] XThR.Tn[10].n28 161.363
R21622 XThR.Tn[10] XThR.Tn[10].n23 161.363
R21623 XThR.Tn[10] XThR.Tn[10].n18 161.363
R21624 XThR.Tn[10] XThR.Tn[10].n13 161.363
R21625 XThR.Tn[10] XThR.Tn[10].n8 161.363
R21626 XThR.Tn[10] XThR.Tn[10].n6 161.363
R21627 XThR.Tn[10].n80 XThR.Tn[10].n79 161.3
R21628 XThR.Tn[10].n75 XThR.Tn[10].n74 161.3
R21629 XThR.Tn[10].n70 XThR.Tn[10].n69 161.3
R21630 XThR.Tn[10].n65 XThR.Tn[10].n64 161.3
R21631 XThR.Tn[10].n60 XThR.Tn[10].n59 161.3
R21632 XThR.Tn[10].n55 XThR.Tn[10].n54 161.3
R21633 XThR.Tn[10].n50 XThR.Tn[10].n49 161.3
R21634 XThR.Tn[10].n45 XThR.Tn[10].n44 161.3
R21635 XThR.Tn[10].n40 XThR.Tn[10].n39 161.3
R21636 XThR.Tn[10].n35 XThR.Tn[10].n34 161.3
R21637 XThR.Tn[10].n30 XThR.Tn[10].n29 161.3
R21638 XThR.Tn[10].n25 XThR.Tn[10].n24 161.3
R21639 XThR.Tn[10].n20 XThR.Tn[10].n19 161.3
R21640 XThR.Tn[10].n15 XThR.Tn[10].n14 161.3
R21641 XThR.Tn[10].n10 XThR.Tn[10].n9 161.3
R21642 XThR.Tn[10].n78 XThR.Tn[10].t37 161.106
R21643 XThR.Tn[10].n73 XThR.Tn[10].t45 161.106
R21644 XThR.Tn[10].n68 XThR.Tn[10].t27 161.106
R21645 XThR.Tn[10].n63 XThR.Tn[10].t72 161.106
R21646 XThR.Tn[10].n58 XThR.Tn[10].t35 161.106
R21647 XThR.Tn[10].n53 XThR.Tn[10].t61 161.106
R21648 XThR.Tn[10].n48 XThR.Tn[10].t43 161.106
R21649 XThR.Tn[10].n43 XThR.Tn[10].t24 161.106
R21650 XThR.Tn[10].n38 XThR.Tn[10].t69 161.106
R21651 XThR.Tn[10].n33 XThR.Tn[10].t15 161.106
R21652 XThR.Tn[10].n28 XThR.Tn[10].t59 161.106
R21653 XThR.Tn[10].n23 XThR.Tn[10].t26 161.106
R21654 XThR.Tn[10].n18 XThR.Tn[10].t58 161.106
R21655 XThR.Tn[10].n13 XThR.Tn[10].t41 161.106
R21656 XThR.Tn[10].n8 XThR.Tn[10].t63 161.106
R21657 XThR.Tn[10].n6 XThR.Tn[10].t47 161.106
R21658 XThR.Tn[10].n79 XThR.Tn[10].t34 159.978
R21659 XThR.Tn[10].n74 XThR.Tn[10].t39 159.978
R21660 XThR.Tn[10].n69 XThR.Tn[10].t22 159.978
R21661 XThR.Tn[10].n64 XThR.Tn[10].t68 159.978
R21662 XThR.Tn[10].n59 XThR.Tn[10].t32 159.978
R21663 XThR.Tn[10].n54 XThR.Tn[10].t57 159.978
R21664 XThR.Tn[10].n49 XThR.Tn[10].t38 159.978
R21665 XThR.Tn[10].n44 XThR.Tn[10].t20 159.978
R21666 XThR.Tn[10].n39 XThR.Tn[10].t66 159.978
R21667 XThR.Tn[10].n34 XThR.Tn[10].t12 159.978
R21668 XThR.Tn[10].n29 XThR.Tn[10].t56 159.978
R21669 XThR.Tn[10].n24 XThR.Tn[10].t21 159.978
R21670 XThR.Tn[10].n19 XThR.Tn[10].t55 159.978
R21671 XThR.Tn[10].n14 XThR.Tn[10].t36 159.978
R21672 XThR.Tn[10].n9 XThR.Tn[10].t60 159.978
R21673 XThR.Tn[10].n78 XThR.Tn[10].t29 145.038
R21674 XThR.Tn[10].n73 XThR.Tn[10].t49 145.038
R21675 XThR.Tn[10].n68 XThR.Tn[10].t31 145.038
R21676 XThR.Tn[10].n63 XThR.Tn[10].t16 145.038
R21677 XThR.Tn[10].n58 XThR.Tn[10].t46 145.038
R21678 XThR.Tn[10].n53 XThR.Tn[10].t28 145.038
R21679 XThR.Tn[10].n48 XThR.Tn[10].t33 145.038
R21680 XThR.Tn[10].n43 XThR.Tn[10].t17 145.038
R21681 XThR.Tn[10].n38 XThR.Tn[10].t14 145.038
R21682 XThR.Tn[10].n33 XThR.Tn[10].t44 145.038
R21683 XThR.Tn[10].n28 XThR.Tn[10].t67 145.038
R21684 XThR.Tn[10].n23 XThR.Tn[10].t30 145.038
R21685 XThR.Tn[10].n18 XThR.Tn[10].t65 145.038
R21686 XThR.Tn[10].n13 XThR.Tn[10].t48 145.038
R21687 XThR.Tn[10].n8 XThR.Tn[10].t13 145.038
R21688 XThR.Tn[10].n6 XThR.Tn[10].t54 145.038
R21689 XThR.Tn[10].n79 XThR.Tn[10].t64 143.911
R21690 XThR.Tn[10].n74 XThR.Tn[10].t25 143.911
R21691 XThR.Tn[10].n69 XThR.Tn[10].t71 143.911
R21692 XThR.Tn[10].n64 XThR.Tn[10].t52 143.911
R21693 XThR.Tn[10].n59 XThR.Tn[10].t19 143.911
R21694 XThR.Tn[10].n54 XThR.Tn[10].t62 143.911
R21695 XThR.Tn[10].n49 XThR.Tn[10].t73 143.911
R21696 XThR.Tn[10].n44 XThR.Tn[10].t53 143.911
R21697 XThR.Tn[10].n39 XThR.Tn[10].t51 143.911
R21698 XThR.Tn[10].n34 XThR.Tn[10].t18 143.911
R21699 XThR.Tn[10].n29 XThR.Tn[10].t42 143.911
R21700 XThR.Tn[10].n24 XThR.Tn[10].t70 143.911
R21701 XThR.Tn[10].n19 XThR.Tn[10].t40 143.911
R21702 XThR.Tn[10].n14 XThR.Tn[10].t23 143.911
R21703 XThR.Tn[10].n9 XThR.Tn[10].t50 143.911
R21704 XThR.Tn[10] XThR.Tn[10].n2 35.7652
R21705 XThR.Tn[10].n85 XThR.Tn[10].t4 26.5955
R21706 XThR.Tn[10].n85 XThR.Tn[10].t5 26.5955
R21707 XThR.Tn[10].n0 XThR.Tn[10].t10 26.5955
R21708 XThR.Tn[10].n0 XThR.Tn[10].t8 26.5955
R21709 XThR.Tn[10].n1 XThR.Tn[10].t11 26.5955
R21710 XThR.Tn[10].n1 XThR.Tn[10].t9 26.5955
R21711 XThR.Tn[10].n86 XThR.Tn[10].t1 26.5955
R21712 XThR.Tn[10].n86 XThR.Tn[10].t0 26.5955
R21713 XThR.Tn[10].n4 XThR.Tn[10].t2 24.9236
R21714 XThR.Tn[10].n4 XThR.Tn[10].t3 24.9236
R21715 XThR.Tn[10].n3 XThR.Tn[10].t7 24.9236
R21716 XThR.Tn[10].n3 XThR.Tn[10].t6 24.9236
R21717 XThR.Tn[10] XThR.Tn[10].n5 18.8943
R21718 XThR.Tn[10].n88 XThR.Tn[10].n87 13.5534
R21719 XThR.Tn[10].n84 XThR.Tn[10] 7.84567
R21720 XThR.Tn[10].n84 XThR.Tn[10] 6.34069
R21721 XThR.Tn[10] XThR.Tn[10].n7 5.34038
R21722 XThR.Tn[10].n12 XThR.Tn[10].n11 4.5005
R21723 XThR.Tn[10].n17 XThR.Tn[10].n16 4.5005
R21724 XThR.Tn[10].n22 XThR.Tn[10].n21 4.5005
R21725 XThR.Tn[10].n27 XThR.Tn[10].n26 4.5005
R21726 XThR.Tn[10].n32 XThR.Tn[10].n31 4.5005
R21727 XThR.Tn[10].n37 XThR.Tn[10].n36 4.5005
R21728 XThR.Tn[10].n42 XThR.Tn[10].n41 4.5005
R21729 XThR.Tn[10].n47 XThR.Tn[10].n46 4.5005
R21730 XThR.Tn[10].n52 XThR.Tn[10].n51 4.5005
R21731 XThR.Tn[10].n57 XThR.Tn[10].n56 4.5005
R21732 XThR.Tn[10].n62 XThR.Tn[10].n61 4.5005
R21733 XThR.Tn[10].n67 XThR.Tn[10].n66 4.5005
R21734 XThR.Tn[10].n72 XThR.Tn[10].n71 4.5005
R21735 XThR.Tn[10].n77 XThR.Tn[10].n76 4.5005
R21736 XThR.Tn[10].n82 XThR.Tn[10].n81 4.5005
R21737 XThR.Tn[10].n83 XThR.Tn[10] 3.70586
R21738 XThR.Tn[10].n12 XThR.Tn[10] 2.52282
R21739 XThR.Tn[10].n17 XThR.Tn[10] 2.52282
R21740 XThR.Tn[10].n22 XThR.Tn[10] 2.52282
R21741 XThR.Tn[10].n27 XThR.Tn[10] 2.52282
R21742 XThR.Tn[10].n32 XThR.Tn[10] 2.52282
R21743 XThR.Tn[10].n37 XThR.Tn[10] 2.52282
R21744 XThR.Tn[10].n42 XThR.Tn[10] 2.52282
R21745 XThR.Tn[10].n47 XThR.Tn[10] 2.52282
R21746 XThR.Tn[10].n52 XThR.Tn[10] 2.52282
R21747 XThR.Tn[10].n57 XThR.Tn[10] 2.52282
R21748 XThR.Tn[10].n62 XThR.Tn[10] 2.52282
R21749 XThR.Tn[10].n67 XThR.Tn[10] 2.52282
R21750 XThR.Tn[10].n72 XThR.Tn[10] 2.52282
R21751 XThR.Tn[10].n77 XThR.Tn[10] 2.52282
R21752 XThR.Tn[10].n82 XThR.Tn[10] 2.52282
R21753 XThR.Tn[10] XThR.Tn[10].n84 1.79489
R21754 XThR.Tn[10] XThR.Tn[10].n88 1.50638
R21755 XThR.Tn[10].n88 XThR.Tn[10] 1.19676
R21756 XThR.Tn[10].n80 XThR.Tn[10] 1.08677
R21757 XThR.Tn[10].n75 XThR.Tn[10] 1.08677
R21758 XThR.Tn[10].n70 XThR.Tn[10] 1.08677
R21759 XThR.Tn[10].n65 XThR.Tn[10] 1.08677
R21760 XThR.Tn[10].n60 XThR.Tn[10] 1.08677
R21761 XThR.Tn[10].n55 XThR.Tn[10] 1.08677
R21762 XThR.Tn[10].n50 XThR.Tn[10] 1.08677
R21763 XThR.Tn[10].n45 XThR.Tn[10] 1.08677
R21764 XThR.Tn[10].n40 XThR.Tn[10] 1.08677
R21765 XThR.Tn[10].n35 XThR.Tn[10] 1.08677
R21766 XThR.Tn[10].n30 XThR.Tn[10] 1.08677
R21767 XThR.Tn[10].n25 XThR.Tn[10] 1.08677
R21768 XThR.Tn[10].n20 XThR.Tn[10] 1.08677
R21769 XThR.Tn[10].n15 XThR.Tn[10] 1.08677
R21770 XThR.Tn[10].n10 XThR.Tn[10] 1.08677
R21771 XThR.Tn[10] XThR.Tn[10].n12 0.839786
R21772 XThR.Tn[10] XThR.Tn[10].n17 0.839786
R21773 XThR.Tn[10] XThR.Tn[10].n22 0.839786
R21774 XThR.Tn[10] XThR.Tn[10].n27 0.839786
R21775 XThR.Tn[10] XThR.Tn[10].n32 0.839786
R21776 XThR.Tn[10] XThR.Tn[10].n37 0.839786
R21777 XThR.Tn[10] XThR.Tn[10].n42 0.839786
R21778 XThR.Tn[10] XThR.Tn[10].n47 0.839786
R21779 XThR.Tn[10] XThR.Tn[10].n52 0.839786
R21780 XThR.Tn[10] XThR.Tn[10].n57 0.839786
R21781 XThR.Tn[10] XThR.Tn[10].n62 0.839786
R21782 XThR.Tn[10] XThR.Tn[10].n67 0.839786
R21783 XThR.Tn[10] XThR.Tn[10].n72 0.839786
R21784 XThR.Tn[10] XThR.Tn[10].n77 0.839786
R21785 XThR.Tn[10] XThR.Tn[10].n82 0.839786
R21786 XThR.Tn[10].n7 XThR.Tn[10] 0.499542
R21787 XThR.Tn[10].n81 XThR.Tn[10] 0.063
R21788 XThR.Tn[10].n76 XThR.Tn[10] 0.063
R21789 XThR.Tn[10].n71 XThR.Tn[10] 0.063
R21790 XThR.Tn[10].n66 XThR.Tn[10] 0.063
R21791 XThR.Tn[10].n61 XThR.Tn[10] 0.063
R21792 XThR.Tn[10].n56 XThR.Tn[10] 0.063
R21793 XThR.Tn[10].n51 XThR.Tn[10] 0.063
R21794 XThR.Tn[10].n46 XThR.Tn[10] 0.063
R21795 XThR.Tn[10].n41 XThR.Tn[10] 0.063
R21796 XThR.Tn[10].n36 XThR.Tn[10] 0.063
R21797 XThR.Tn[10].n31 XThR.Tn[10] 0.063
R21798 XThR.Tn[10].n26 XThR.Tn[10] 0.063
R21799 XThR.Tn[10].n21 XThR.Tn[10] 0.063
R21800 XThR.Tn[10].n16 XThR.Tn[10] 0.063
R21801 XThR.Tn[10].n11 XThR.Tn[10] 0.063
R21802 XThR.Tn[10].n83 XThR.Tn[10] 0.0540714
R21803 XThR.Tn[10] XThR.Tn[10].n83 0.038
R21804 XThR.Tn[10].n7 XThR.Tn[10] 0.0143889
R21805 XThR.Tn[10].n81 XThR.Tn[10].n80 0.00771154
R21806 XThR.Tn[10].n76 XThR.Tn[10].n75 0.00771154
R21807 XThR.Tn[10].n71 XThR.Tn[10].n70 0.00771154
R21808 XThR.Tn[10].n66 XThR.Tn[10].n65 0.00771154
R21809 XThR.Tn[10].n61 XThR.Tn[10].n60 0.00771154
R21810 XThR.Tn[10].n56 XThR.Tn[10].n55 0.00771154
R21811 XThR.Tn[10].n51 XThR.Tn[10].n50 0.00771154
R21812 XThR.Tn[10].n46 XThR.Tn[10].n45 0.00771154
R21813 XThR.Tn[10].n41 XThR.Tn[10].n40 0.00771154
R21814 XThR.Tn[10].n36 XThR.Tn[10].n35 0.00771154
R21815 XThR.Tn[10].n31 XThR.Tn[10].n30 0.00771154
R21816 XThR.Tn[10].n26 XThR.Tn[10].n25 0.00771154
R21817 XThR.Tn[10].n21 XThR.Tn[10].n20 0.00771154
R21818 XThR.Tn[10].n16 XThR.Tn[10].n15 0.00771154
R21819 XThR.Tn[10].n11 XThR.Tn[10].n10 0.00771154
R21820 XThC.Tn[14].n70 XThC.Tn[14].n69 256.104
R21821 XThC.Tn[14].n74 XThC.Tn[14].n73 243.679
R21822 XThC.Tn[14].n2 XThC.Tn[14].n0 241.847
R21823 XThC.Tn[14].n74 XThC.Tn[14].n72 205.28
R21824 XThC.Tn[14].n70 XThC.Tn[14].n68 202.095
R21825 XThC.Tn[14].n2 XThC.Tn[14].n1 185
R21826 XThC.Tn[14].n64 XThC.Tn[14].n62 161.365
R21827 XThC.Tn[14].n60 XThC.Tn[14].n58 161.365
R21828 XThC.Tn[14].n56 XThC.Tn[14].n54 161.365
R21829 XThC.Tn[14].n52 XThC.Tn[14].n50 161.365
R21830 XThC.Tn[14].n48 XThC.Tn[14].n46 161.365
R21831 XThC.Tn[14].n44 XThC.Tn[14].n42 161.365
R21832 XThC.Tn[14].n40 XThC.Tn[14].n38 161.365
R21833 XThC.Tn[14].n36 XThC.Tn[14].n34 161.365
R21834 XThC.Tn[14].n32 XThC.Tn[14].n30 161.365
R21835 XThC.Tn[14].n28 XThC.Tn[14].n26 161.365
R21836 XThC.Tn[14].n24 XThC.Tn[14].n22 161.365
R21837 XThC.Tn[14].n20 XThC.Tn[14].n18 161.365
R21838 XThC.Tn[14].n16 XThC.Tn[14].n14 161.365
R21839 XThC.Tn[14].n12 XThC.Tn[14].n10 161.365
R21840 XThC.Tn[14].n8 XThC.Tn[14].n6 161.365
R21841 XThC.Tn[14].n5 XThC.Tn[14].n3 161.365
R21842 XThC.Tn[14].n62 XThC.Tn[14].t12 161.202
R21843 XThC.Tn[14].n58 XThC.Tn[14].t33 161.202
R21844 XThC.Tn[14].n54 XThC.Tn[14].t21 161.202
R21845 XThC.Tn[14].n50 XThC.Tn[14].t19 161.202
R21846 XThC.Tn[14].n46 XThC.Tn[14].t42 161.202
R21847 XThC.Tn[14].n42 XThC.Tn[14].t30 161.202
R21848 XThC.Tn[14].n38 XThC.Tn[14].t27 161.202
R21849 XThC.Tn[14].n34 XThC.Tn[14].t41 161.202
R21850 XThC.Tn[14].n30 XThC.Tn[14].t39 161.202
R21851 XThC.Tn[14].n26 XThC.Tn[14].t31 161.202
R21852 XThC.Tn[14].n22 XThC.Tn[14].t17 161.202
R21853 XThC.Tn[14].n18 XThC.Tn[14].t14 161.202
R21854 XThC.Tn[14].n14 XThC.Tn[14].t26 161.202
R21855 XThC.Tn[14].n10 XThC.Tn[14].t25 161.202
R21856 XThC.Tn[14].n6 XThC.Tn[14].t22 161.202
R21857 XThC.Tn[14].n3 XThC.Tn[14].t38 161.202
R21858 XThC.Tn[14].n62 XThC.Tn[14].t18 145.137
R21859 XThC.Tn[14].n58 XThC.Tn[14].t40 145.137
R21860 XThC.Tn[14].n54 XThC.Tn[14].t28 145.137
R21861 XThC.Tn[14].n50 XThC.Tn[14].t24 145.137
R21862 XThC.Tn[14].n46 XThC.Tn[14].t16 145.137
R21863 XThC.Tn[14].n42 XThC.Tn[14].t36 145.137
R21864 XThC.Tn[14].n38 XThC.Tn[14].t35 145.137
R21865 XThC.Tn[14].n34 XThC.Tn[14].t15 145.137
R21866 XThC.Tn[14].n30 XThC.Tn[14].t13 145.137
R21867 XThC.Tn[14].n26 XThC.Tn[14].t37 145.137
R21868 XThC.Tn[14].n22 XThC.Tn[14].t23 145.137
R21869 XThC.Tn[14].n18 XThC.Tn[14].t20 145.137
R21870 XThC.Tn[14].n14 XThC.Tn[14].t34 145.137
R21871 XThC.Tn[14].n10 XThC.Tn[14].t32 145.137
R21872 XThC.Tn[14].n6 XThC.Tn[14].t29 145.137
R21873 XThC.Tn[14].n3 XThC.Tn[14].t43 145.137
R21874 XThC.Tn[14].n68 XThC.Tn[14].t4 26.5955
R21875 XThC.Tn[14].n68 XThC.Tn[14].t5 26.5955
R21876 XThC.Tn[14].n69 XThC.Tn[14].t7 26.5955
R21877 XThC.Tn[14].n69 XThC.Tn[14].t6 26.5955
R21878 XThC.Tn[14].n72 XThC.Tn[14].t1 26.5955
R21879 XThC.Tn[14].n72 XThC.Tn[14].t0 26.5955
R21880 XThC.Tn[14].n73 XThC.Tn[14].t3 26.5955
R21881 XThC.Tn[14].n73 XThC.Tn[14].t2 26.5955
R21882 XThC.Tn[14].n1 XThC.Tn[14].t9 24.9236
R21883 XThC.Tn[14].n1 XThC.Tn[14].t11 24.9236
R21884 XThC.Tn[14].n0 XThC.Tn[14].t8 24.9236
R21885 XThC.Tn[14].n0 XThC.Tn[14].t10 24.9236
R21886 XThC.Tn[14] XThC.Tn[14].n74 22.9652
R21887 XThC.Tn[14] XThC.Tn[14].n2 22.9615
R21888 XThC.Tn[14].n71 XThC.Tn[14].n70 13.9299
R21889 XThC.Tn[14] XThC.Tn[14].n71 13.9299
R21890 XThC.Tn[14] XThC.Tn[14].n5 8.0245
R21891 XThC.Tn[14].n65 XThC.Tn[14].n64 7.9105
R21892 XThC.Tn[14].n61 XThC.Tn[14].n60 7.9105
R21893 XThC.Tn[14].n57 XThC.Tn[14].n56 7.9105
R21894 XThC.Tn[14].n53 XThC.Tn[14].n52 7.9105
R21895 XThC.Tn[14].n49 XThC.Tn[14].n48 7.9105
R21896 XThC.Tn[14].n45 XThC.Tn[14].n44 7.9105
R21897 XThC.Tn[14].n41 XThC.Tn[14].n40 7.9105
R21898 XThC.Tn[14].n37 XThC.Tn[14].n36 7.9105
R21899 XThC.Tn[14].n33 XThC.Tn[14].n32 7.9105
R21900 XThC.Tn[14].n29 XThC.Tn[14].n28 7.9105
R21901 XThC.Tn[14].n25 XThC.Tn[14].n24 7.9105
R21902 XThC.Tn[14].n21 XThC.Tn[14].n20 7.9105
R21903 XThC.Tn[14].n17 XThC.Tn[14].n16 7.9105
R21904 XThC.Tn[14].n13 XThC.Tn[14].n12 7.9105
R21905 XThC.Tn[14].n9 XThC.Tn[14].n8 7.9105
R21906 XThC.Tn[14].n67 XThC.Tn[14].n66 7.51947
R21907 XThC.Tn[14].n66 XThC.Tn[14] 5.85107
R21908 XThC.Tn[14].n71 XThC.Tn[14].n67 2.99115
R21909 XThC.Tn[14].n71 XThC.Tn[14] 2.87153
R21910 XThC.Tn[14].n67 XThC.Tn[14] 2.2734
R21911 XThC.Tn[14].n66 XThC.Tn[14] 1.06164
R21912 XThC.Tn[14].n9 XThC.Tn[14] 0.235138
R21913 XThC.Tn[14].n13 XThC.Tn[14] 0.235138
R21914 XThC.Tn[14].n17 XThC.Tn[14] 0.235138
R21915 XThC.Tn[14].n21 XThC.Tn[14] 0.235138
R21916 XThC.Tn[14].n25 XThC.Tn[14] 0.235138
R21917 XThC.Tn[14].n29 XThC.Tn[14] 0.235138
R21918 XThC.Tn[14].n33 XThC.Tn[14] 0.235138
R21919 XThC.Tn[14].n37 XThC.Tn[14] 0.235138
R21920 XThC.Tn[14].n41 XThC.Tn[14] 0.235138
R21921 XThC.Tn[14].n45 XThC.Tn[14] 0.235138
R21922 XThC.Tn[14].n49 XThC.Tn[14] 0.235138
R21923 XThC.Tn[14].n53 XThC.Tn[14] 0.235138
R21924 XThC.Tn[14].n57 XThC.Tn[14] 0.235138
R21925 XThC.Tn[14].n61 XThC.Tn[14] 0.235138
R21926 XThC.Tn[14].n65 XThC.Tn[14] 0.235138
R21927 XThC.Tn[14] XThC.Tn[14].n9 0.114505
R21928 XThC.Tn[14] XThC.Tn[14].n13 0.114505
R21929 XThC.Tn[14] XThC.Tn[14].n17 0.114505
R21930 XThC.Tn[14] XThC.Tn[14].n21 0.114505
R21931 XThC.Tn[14] XThC.Tn[14].n25 0.114505
R21932 XThC.Tn[14] XThC.Tn[14].n29 0.114505
R21933 XThC.Tn[14] XThC.Tn[14].n33 0.114505
R21934 XThC.Tn[14] XThC.Tn[14].n37 0.114505
R21935 XThC.Tn[14] XThC.Tn[14].n41 0.114505
R21936 XThC.Tn[14] XThC.Tn[14].n45 0.114505
R21937 XThC.Tn[14] XThC.Tn[14].n49 0.114505
R21938 XThC.Tn[14] XThC.Tn[14].n53 0.114505
R21939 XThC.Tn[14] XThC.Tn[14].n57 0.114505
R21940 XThC.Tn[14] XThC.Tn[14].n61 0.114505
R21941 XThC.Tn[14] XThC.Tn[14].n65 0.114505
R21942 XThC.Tn[14].n64 XThC.Tn[14].n63 0.0599512
R21943 XThC.Tn[14].n60 XThC.Tn[14].n59 0.0599512
R21944 XThC.Tn[14].n56 XThC.Tn[14].n55 0.0599512
R21945 XThC.Tn[14].n52 XThC.Tn[14].n51 0.0599512
R21946 XThC.Tn[14].n48 XThC.Tn[14].n47 0.0599512
R21947 XThC.Tn[14].n44 XThC.Tn[14].n43 0.0599512
R21948 XThC.Tn[14].n40 XThC.Tn[14].n39 0.0599512
R21949 XThC.Tn[14].n36 XThC.Tn[14].n35 0.0599512
R21950 XThC.Tn[14].n32 XThC.Tn[14].n31 0.0599512
R21951 XThC.Tn[14].n28 XThC.Tn[14].n27 0.0599512
R21952 XThC.Tn[14].n24 XThC.Tn[14].n23 0.0599512
R21953 XThC.Tn[14].n20 XThC.Tn[14].n19 0.0599512
R21954 XThC.Tn[14].n16 XThC.Tn[14].n15 0.0599512
R21955 XThC.Tn[14].n12 XThC.Tn[14].n11 0.0599512
R21956 XThC.Tn[14].n8 XThC.Tn[14].n7 0.0599512
R21957 XThC.Tn[14].n5 XThC.Tn[14].n4 0.0599512
R21958 XThC.Tn[14].n63 XThC.Tn[14] 0.0469286
R21959 XThC.Tn[14].n59 XThC.Tn[14] 0.0469286
R21960 XThC.Tn[14].n55 XThC.Tn[14] 0.0469286
R21961 XThC.Tn[14].n51 XThC.Tn[14] 0.0469286
R21962 XThC.Tn[14].n47 XThC.Tn[14] 0.0469286
R21963 XThC.Tn[14].n43 XThC.Tn[14] 0.0469286
R21964 XThC.Tn[14].n39 XThC.Tn[14] 0.0469286
R21965 XThC.Tn[14].n35 XThC.Tn[14] 0.0469286
R21966 XThC.Tn[14].n31 XThC.Tn[14] 0.0469286
R21967 XThC.Tn[14].n27 XThC.Tn[14] 0.0469286
R21968 XThC.Tn[14].n23 XThC.Tn[14] 0.0469286
R21969 XThC.Tn[14].n19 XThC.Tn[14] 0.0469286
R21970 XThC.Tn[14].n15 XThC.Tn[14] 0.0469286
R21971 XThC.Tn[14].n11 XThC.Tn[14] 0.0469286
R21972 XThC.Tn[14].n7 XThC.Tn[14] 0.0469286
R21973 XThC.Tn[14].n4 XThC.Tn[14] 0.0469286
R21974 XThC.Tn[14].n63 XThC.Tn[14] 0.0401341
R21975 XThC.Tn[14].n59 XThC.Tn[14] 0.0401341
R21976 XThC.Tn[14].n55 XThC.Tn[14] 0.0401341
R21977 XThC.Tn[14].n51 XThC.Tn[14] 0.0401341
R21978 XThC.Tn[14].n47 XThC.Tn[14] 0.0401341
R21979 XThC.Tn[14].n43 XThC.Tn[14] 0.0401341
R21980 XThC.Tn[14].n39 XThC.Tn[14] 0.0401341
R21981 XThC.Tn[14].n35 XThC.Tn[14] 0.0401341
R21982 XThC.Tn[14].n31 XThC.Tn[14] 0.0401341
R21983 XThC.Tn[14].n27 XThC.Tn[14] 0.0401341
R21984 XThC.Tn[14].n23 XThC.Tn[14] 0.0401341
R21985 XThC.Tn[14].n19 XThC.Tn[14] 0.0401341
R21986 XThC.Tn[14].n15 XThC.Tn[14] 0.0401341
R21987 XThC.Tn[14].n11 XThC.Tn[14] 0.0401341
R21988 XThC.Tn[14].n7 XThC.Tn[14] 0.0401341
R21989 XThC.Tn[14].n4 XThC.Tn[14] 0.0401341
R21990 XThC.XTB1.Y.n6 XThC.XTB1.Y.t11 212.081
R21991 XThC.XTB1.Y.n5 XThC.XTB1.Y.t8 212.081
R21992 XThC.XTB1.Y.n11 XThC.XTB1.Y.t6 212.081
R21993 XThC.XTB1.Y.n3 XThC.XTB1.Y.t17 212.081
R21994 XThC.XTB1.Y.n15 XThC.XTB1.Y.t10 212.081
R21995 XThC.XTB1.Y.n16 XThC.XTB1.Y.t14 212.081
R21996 XThC.XTB1.Y.n18 XThC.XTB1.Y.t7 212.081
R21997 XThC.XTB1.Y.n14 XThC.XTB1.Y.t18 212.081
R21998 XThC.XTB1.Y.n22 XThC.XTB1.Y.n2 201.288
R21999 XThC.XTB1.Y.n8 XThC.XTB1.Y.n7 173.761
R22000 XThC.XTB1.Y.n17 XThC.XTB1.Y 158.656
R22001 XThC.XTB1.Y.n10 XThC.XTB1.Y.n9 152
R22002 XThC.XTB1.Y.n8 XThC.XTB1.Y.n4 152
R22003 XThC.XTB1.Y.n13 XThC.XTB1.Y.n12 152
R22004 XThC.XTB1.Y.n20 XThC.XTB1.Y.n19 152
R22005 XThC.XTB1.Y.n6 XThC.XTB1.Y.t16 139.78
R22006 XThC.XTB1.Y.n5 XThC.XTB1.Y.t13 139.78
R22007 XThC.XTB1.Y.n11 XThC.XTB1.Y.t12 139.78
R22008 XThC.XTB1.Y.n3 XThC.XTB1.Y.t5 139.78
R22009 XThC.XTB1.Y.n15 XThC.XTB1.Y.t4 139.78
R22010 XThC.XTB1.Y.n16 XThC.XTB1.Y.t3 139.78
R22011 XThC.XTB1.Y.n18 XThC.XTB1.Y.t15 139.78
R22012 XThC.XTB1.Y.n14 XThC.XTB1.Y.t9 139.78
R22013 XThC.XTB1.Y.n0 XThC.XTB1.Y.t2 132.067
R22014 XThC.XTB1.Y.n21 XThC.XTB1.Y 83.4676
R22015 XThC.XTB1.Y.n21 XThC.XTB1.Y.n13 61.4091
R22016 XThC.XTB1.Y.n16 XThC.XTB1.Y.n15 61.346
R22017 XThC.XTB1.Y.n10 XThC.XTB1.Y.n4 49.6611
R22018 XThC.XTB1.Y.n12 XThC.XTB1.Y.n11 45.2793
R22019 XThC.XTB1.Y.n7 XThC.XTB1.Y.n5 42.3581
R22020 XThC.XTB1.Y.n19 XThC.XTB1.Y.n14 30.6732
R22021 XThC.XTB1.Y.n19 XThC.XTB1.Y.n18 30.6732
R22022 XThC.XTB1.Y.n18 XThC.XTB1.Y.n17 30.6732
R22023 XThC.XTB1.Y.n17 XThC.XTB1.Y.n16 30.6732
R22024 XThC.XTB1.Y.n2 XThC.XTB1.Y.t1 26.5955
R22025 XThC.XTB1.Y.n2 XThC.XTB1.Y.t0 26.5955
R22026 XThC.XTB1.Y XThC.XTB1.Y.n22 23.489
R22027 XThC.XTB1.Y.n9 XThC.XTB1.Y.n8 21.7605
R22028 XThC.XTB1.Y.n7 XThC.XTB1.Y.n6 18.9884
R22029 XThC.XTB1.Y.n12 XThC.XTB1.Y.n3 16.0672
R22030 XThC.XTB1.Y.n20 XThC.XTB1.Y 14.8485
R22031 XThC.XTB1.Y.n13 XThC.XTB1.Y 11.5205
R22032 XThC.XTB1.Y.n22 XThC.XTB1.Y.n21 10.7939
R22033 XThC.XTB1.Y.n9 XThC.XTB1.Y 10.2405
R22034 XThC.XTB1.Y XThC.XTB1.Y.n20 8.7045
R22035 XThC.XTB1.Y.n5 XThC.XTB1.Y.n4 7.30353
R22036 XThC.XTB1.Y.n11 XThC.XTB1.Y.n10 4.38232
R22037 XThC.XTB1.Y.n1 XThC.XTB1.Y.n0 4.15748
R22038 XThC.XTB1.Y XThC.XTB1.Y.n1 3.76521
R22039 XThC.XTB1.Y.n0 XThC.XTB1.Y 1.17559
R22040 XThC.XTB1.Y.n1 XThC.XTB1.Y 0.921363
R22041 XThC.Tn[8].n71 XThC.Tn[8].n70 256.104
R22042 XThC.Tn[8].n75 XThC.Tn[8].n74 243.679
R22043 XThC.Tn[8].n2 XThC.Tn[8].n0 241.847
R22044 XThC.Tn[8].n75 XThC.Tn[8].n73 205.28
R22045 XThC.Tn[8].n71 XThC.Tn[8].n69 202.095
R22046 XThC.Tn[8].n2 XThC.Tn[8].n1 185
R22047 XThC.Tn[8].n65 XThC.Tn[8].n63 161.365
R22048 XThC.Tn[8].n61 XThC.Tn[8].n59 161.365
R22049 XThC.Tn[8].n57 XThC.Tn[8].n55 161.365
R22050 XThC.Tn[8].n53 XThC.Tn[8].n51 161.365
R22051 XThC.Tn[8].n49 XThC.Tn[8].n47 161.365
R22052 XThC.Tn[8].n45 XThC.Tn[8].n43 161.365
R22053 XThC.Tn[8].n41 XThC.Tn[8].n39 161.365
R22054 XThC.Tn[8].n37 XThC.Tn[8].n35 161.365
R22055 XThC.Tn[8].n33 XThC.Tn[8].n31 161.365
R22056 XThC.Tn[8].n29 XThC.Tn[8].n27 161.365
R22057 XThC.Tn[8].n25 XThC.Tn[8].n23 161.365
R22058 XThC.Tn[8].n21 XThC.Tn[8].n19 161.365
R22059 XThC.Tn[8].n17 XThC.Tn[8].n15 161.365
R22060 XThC.Tn[8].n13 XThC.Tn[8].n11 161.365
R22061 XThC.Tn[8].n9 XThC.Tn[8].n7 161.365
R22062 XThC.Tn[8].n6 XThC.Tn[8].n4 161.365
R22063 XThC.Tn[8].n63 XThC.Tn[8].t15 161.202
R22064 XThC.Tn[8].n59 XThC.Tn[8].t37 161.202
R22065 XThC.Tn[8].n55 XThC.Tn[8].t24 161.202
R22066 XThC.Tn[8].n51 XThC.Tn[8].t21 161.202
R22067 XThC.Tn[8].n47 XThC.Tn[8].t13 161.202
R22068 XThC.Tn[8].n43 XThC.Tn[8].t32 161.202
R22069 XThC.Tn[8].n39 XThC.Tn[8].t31 161.202
R22070 XThC.Tn[8].n35 XThC.Tn[8].t12 161.202
R22071 XThC.Tn[8].n31 XThC.Tn[8].t42 161.202
R22072 XThC.Tn[8].n27 XThC.Tn[8].t33 161.202
R22073 XThC.Tn[8].n23 XThC.Tn[8].t20 161.202
R22074 XThC.Tn[8].n19 XThC.Tn[8].t19 161.202
R22075 XThC.Tn[8].n15 XThC.Tn[8].t30 161.202
R22076 XThC.Tn[8].n11 XThC.Tn[8].t28 161.202
R22077 XThC.Tn[8].n7 XThC.Tn[8].t26 161.202
R22078 XThC.Tn[8].n4 XThC.Tn[8].t41 161.202
R22079 XThC.Tn[8].n63 XThC.Tn[8].t18 145.137
R22080 XThC.Tn[8].n59 XThC.Tn[8].t40 145.137
R22081 XThC.Tn[8].n55 XThC.Tn[8].t27 145.137
R22082 XThC.Tn[8].n51 XThC.Tn[8].t25 145.137
R22083 XThC.Tn[8].n47 XThC.Tn[8].t17 145.137
R22084 XThC.Tn[8].n43 XThC.Tn[8].t38 145.137
R22085 XThC.Tn[8].n39 XThC.Tn[8].t36 145.137
R22086 XThC.Tn[8].n35 XThC.Tn[8].t16 145.137
R22087 XThC.Tn[8].n31 XThC.Tn[8].t14 145.137
R22088 XThC.Tn[8].n27 XThC.Tn[8].t39 145.137
R22089 XThC.Tn[8].n23 XThC.Tn[8].t23 145.137
R22090 XThC.Tn[8].n19 XThC.Tn[8].t22 145.137
R22091 XThC.Tn[8].n15 XThC.Tn[8].t35 145.137
R22092 XThC.Tn[8].n11 XThC.Tn[8].t34 145.137
R22093 XThC.Tn[8].n7 XThC.Tn[8].t29 145.137
R22094 XThC.Tn[8].n4 XThC.Tn[8].t43 145.137
R22095 XThC.Tn[8].n69 XThC.Tn[8].t5 26.5955
R22096 XThC.Tn[8].n69 XThC.Tn[8].t6 26.5955
R22097 XThC.Tn[8].n70 XThC.Tn[8].t4 26.5955
R22098 XThC.Tn[8].n70 XThC.Tn[8].t7 26.5955
R22099 XThC.Tn[8].n73 XThC.Tn[8].t2 26.5955
R22100 XThC.Tn[8].n73 XThC.Tn[8].t1 26.5955
R22101 XThC.Tn[8].n74 XThC.Tn[8].t0 26.5955
R22102 XThC.Tn[8].n74 XThC.Tn[8].t3 26.5955
R22103 XThC.Tn[8].n1 XThC.Tn[8].t11 24.9236
R22104 XThC.Tn[8].n1 XThC.Tn[8].t10 24.9236
R22105 XThC.Tn[8].n0 XThC.Tn[8].t9 24.9236
R22106 XThC.Tn[8].n0 XThC.Tn[8].t8 24.9236
R22107 XThC.Tn[8] XThC.Tn[8].n75 22.9652
R22108 XThC.Tn[8] XThC.Tn[8].n2 22.9615
R22109 XThC.Tn[8].n72 XThC.Tn[8].n71 13.9299
R22110 XThC.Tn[8] XThC.Tn[8].n72 13.9299
R22111 XThC.Tn[8] XThC.Tn[8].n6 8.0245
R22112 XThC.Tn[8].n66 XThC.Tn[8].n65 7.9105
R22113 XThC.Tn[8].n62 XThC.Tn[8].n61 7.9105
R22114 XThC.Tn[8].n58 XThC.Tn[8].n57 7.9105
R22115 XThC.Tn[8].n54 XThC.Tn[8].n53 7.9105
R22116 XThC.Tn[8].n50 XThC.Tn[8].n49 7.9105
R22117 XThC.Tn[8].n46 XThC.Tn[8].n45 7.9105
R22118 XThC.Tn[8].n42 XThC.Tn[8].n41 7.9105
R22119 XThC.Tn[8].n38 XThC.Tn[8].n37 7.9105
R22120 XThC.Tn[8].n34 XThC.Tn[8].n33 7.9105
R22121 XThC.Tn[8].n30 XThC.Tn[8].n29 7.9105
R22122 XThC.Tn[8].n26 XThC.Tn[8].n25 7.9105
R22123 XThC.Tn[8].n22 XThC.Tn[8].n21 7.9105
R22124 XThC.Tn[8].n18 XThC.Tn[8].n17 7.9105
R22125 XThC.Tn[8].n14 XThC.Tn[8].n13 7.9105
R22126 XThC.Tn[8].n10 XThC.Tn[8].n9 7.9105
R22127 XThC.Tn[8].n68 XThC.Tn[8].n67 7.42331
R22128 XThC.Tn[8].n67 XThC.Tn[8] 4.24005
R22129 XThC.Tn[8].n72 XThC.Tn[8].n68 2.99115
R22130 XThC.Tn[8].n72 XThC.Tn[8] 2.87153
R22131 XThC.Tn[8].n68 XThC.Tn[8] 2.2734
R22132 XThC.Tn[8].n3 XThC.Tn[8] 0.672375
R22133 XThC.Tn[8].n10 XThC.Tn[8] 0.235138
R22134 XThC.Tn[8].n14 XThC.Tn[8] 0.235138
R22135 XThC.Tn[8].n18 XThC.Tn[8] 0.235138
R22136 XThC.Tn[8].n22 XThC.Tn[8] 0.235138
R22137 XThC.Tn[8].n26 XThC.Tn[8] 0.235138
R22138 XThC.Tn[8].n30 XThC.Tn[8] 0.235138
R22139 XThC.Tn[8].n34 XThC.Tn[8] 0.235138
R22140 XThC.Tn[8].n38 XThC.Tn[8] 0.235138
R22141 XThC.Tn[8].n42 XThC.Tn[8] 0.235138
R22142 XThC.Tn[8].n46 XThC.Tn[8] 0.235138
R22143 XThC.Tn[8].n50 XThC.Tn[8] 0.235138
R22144 XThC.Tn[8].n54 XThC.Tn[8] 0.235138
R22145 XThC.Tn[8].n58 XThC.Tn[8] 0.235138
R22146 XThC.Tn[8].n62 XThC.Tn[8] 0.235138
R22147 XThC.Tn[8].n66 XThC.Tn[8] 0.235138
R22148 XThC.Tn[8].n67 XThC.Tn[8].n3 0.220435
R22149 XThC.Tn[8].n3 XThC.Tn[8] 0.168469
R22150 XThC.Tn[8] XThC.Tn[8].n10 0.114505
R22151 XThC.Tn[8] XThC.Tn[8].n14 0.114505
R22152 XThC.Tn[8] XThC.Tn[8].n18 0.114505
R22153 XThC.Tn[8] XThC.Tn[8].n22 0.114505
R22154 XThC.Tn[8] XThC.Tn[8].n26 0.114505
R22155 XThC.Tn[8] XThC.Tn[8].n30 0.114505
R22156 XThC.Tn[8] XThC.Tn[8].n34 0.114505
R22157 XThC.Tn[8] XThC.Tn[8].n38 0.114505
R22158 XThC.Tn[8] XThC.Tn[8].n42 0.114505
R22159 XThC.Tn[8] XThC.Tn[8].n46 0.114505
R22160 XThC.Tn[8] XThC.Tn[8].n50 0.114505
R22161 XThC.Tn[8] XThC.Tn[8].n54 0.114505
R22162 XThC.Tn[8] XThC.Tn[8].n58 0.114505
R22163 XThC.Tn[8] XThC.Tn[8].n62 0.114505
R22164 XThC.Tn[8] XThC.Tn[8].n66 0.114505
R22165 XThC.Tn[8].n65 XThC.Tn[8].n64 0.0599512
R22166 XThC.Tn[8].n61 XThC.Tn[8].n60 0.0599512
R22167 XThC.Tn[8].n57 XThC.Tn[8].n56 0.0599512
R22168 XThC.Tn[8].n53 XThC.Tn[8].n52 0.0599512
R22169 XThC.Tn[8].n49 XThC.Tn[8].n48 0.0599512
R22170 XThC.Tn[8].n45 XThC.Tn[8].n44 0.0599512
R22171 XThC.Tn[8].n41 XThC.Tn[8].n40 0.0599512
R22172 XThC.Tn[8].n37 XThC.Tn[8].n36 0.0599512
R22173 XThC.Tn[8].n33 XThC.Tn[8].n32 0.0599512
R22174 XThC.Tn[8].n29 XThC.Tn[8].n28 0.0599512
R22175 XThC.Tn[8].n25 XThC.Tn[8].n24 0.0599512
R22176 XThC.Tn[8].n21 XThC.Tn[8].n20 0.0599512
R22177 XThC.Tn[8].n17 XThC.Tn[8].n16 0.0599512
R22178 XThC.Tn[8].n13 XThC.Tn[8].n12 0.0599512
R22179 XThC.Tn[8].n9 XThC.Tn[8].n8 0.0599512
R22180 XThC.Tn[8].n6 XThC.Tn[8].n5 0.0599512
R22181 XThC.Tn[8].n64 XThC.Tn[8] 0.0469286
R22182 XThC.Tn[8].n60 XThC.Tn[8] 0.0469286
R22183 XThC.Tn[8].n56 XThC.Tn[8] 0.0469286
R22184 XThC.Tn[8].n52 XThC.Tn[8] 0.0469286
R22185 XThC.Tn[8].n48 XThC.Tn[8] 0.0469286
R22186 XThC.Tn[8].n44 XThC.Tn[8] 0.0469286
R22187 XThC.Tn[8].n40 XThC.Tn[8] 0.0469286
R22188 XThC.Tn[8].n36 XThC.Tn[8] 0.0469286
R22189 XThC.Tn[8].n32 XThC.Tn[8] 0.0469286
R22190 XThC.Tn[8].n28 XThC.Tn[8] 0.0469286
R22191 XThC.Tn[8].n24 XThC.Tn[8] 0.0469286
R22192 XThC.Tn[8].n20 XThC.Tn[8] 0.0469286
R22193 XThC.Tn[8].n16 XThC.Tn[8] 0.0469286
R22194 XThC.Tn[8].n12 XThC.Tn[8] 0.0469286
R22195 XThC.Tn[8].n8 XThC.Tn[8] 0.0469286
R22196 XThC.Tn[8].n5 XThC.Tn[8] 0.0469286
R22197 XThC.Tn[8].n64 XThC.Tn[8] 0.0401341
R22198 XThC.Tn[8].n60 XThC.Tn[8] 0.0401341
R22199 XThC.Tn[8].n56 XThC.Tn[8] 0.0401341
R22200 XThC.Tn[8].n52 XThC.Tn[8] 0.0401341
R22201 XThC.Tn[8].n48 XThC.Tn[8] 0.0401341
R22202 XThC.Tn[8].n44 XThC.Tn[8] 0.0401341
R22203 XThC.Tn[8].n40 XThC.Tn[8] 0.0401341
R22204 XThC.Tn[8].n36 XThC.Tn[8] 0.0401341
R22205 XThC.Tn[8].n32 XThC.Tn[8] 0.0401341
R22206 XThC.Tn[8].n28 XThC.Tn[8] 0.0401341
R22207 XThC.Tn[8].n24 XThC.Tn[8] 0.0401341
R22208 XThC.Tn[8].n20 XThC.Tn[8] 0.0401341
R22209 XThC.Tn[8].n16 XThC.Tn[8] 0.0401341
R22210 XThC.Tn[8].n12 XThC.Tn[8] 0.0401341
R22211 XThC.Tn[8].n8 XThC.Tn[8] 0.0401341
R22212 XThC.Tn[8].n5 XThC.Tn[8] 0.0401341
R22213 XThR.Tn[1].n2 XThR.Tn[1].n1 332.332
R22214 XThR.Tn[1].n2 XThR.Tn[1].n0 296.493
R22215 XThR.Tn[1] XThR.Tn[1].n82 161.363
R22216 XThR.Tn[1] XThR.Tn[1].n77 161.363
R22217 XThR.Tn[1] XThR.Tn[1].n72 161.363
R22218 XThR.Tn[1] XThR.Tn[1].n67 161.363
R22219 XThR.Tn[1] XThR.Tn[1].n62 161.363
R22220 XThR.Tn[1] XThR.Tn[1].n57 161.363
R22221 XThR.Tn[1] XThR.Tn[1].n52 161.363
R22222 XThR.Tn[1] XThR.Tn[1].n47 161.363
R22223 XThR.Tn[1] XThR.Tn[1].n42 161.363
R22224 XThR.Tn[1] XThR.Tn[1].n37 161.363
R22225 XThR.Tn[1] XThR.Tn[1].n32 161.363
R22226 XThR.Tn[1] XThR.Tn[1].n27 161.363
R22227 XThR.Tn[1] XThR.Tn[1].n22 161.363
R22228 XThR.Tn[1] XThR.Tn[1].n17 161.363
R22229 XThR.Tn[1] XThR.Tn[1].n12 161.363
R22230 XThR.Tn[1] XThR.Tn[1].n10 161.363
R22231 XThR.Tn[1].n84 XThR.Tn[1].n83 161.3
R22232 XThR.Tn[1].n79 XThR.Tn[1].n78 161.3
R22233 XThR.Tn[1].n74 XThR.Tn[1].n73 161.3
R22234 XThR.Tn[1].n69 XThR.Tn[1].n68 161.3
R22235 XThR.Tn[1].n64 XThR.Tn[1].n63 161.3
R22236 XThR.Tn[1].n59 XThR.Tn[1].n58 161.3
R22237 XThR.Tn[1].n54 XThR.Tn[1].n53 161.3
R22238 XThR.Tn[1].n49 XThR.Tn[1].n48 161.3
R22239 XThR.Tn[1].n44 XThR.Tn[1].n43 161.3
R22240 XThR.Tn[1].n39 XThR.Tn[1].n38 161.3
R22241 XThR.Tn[1].n34 XThR.Tn[1].n33 161.3
R22242 XThR.Tn[1].n29 XThR.Tn[1].n28 161.3
R22243 XThR.Tn[1].n24 XThR.Tn[1].n23 161.3
R22244 XThR.Tn[1].n19 XThR.Tn[1].n18 161.3
R22245 XThR.Tn[1].n14 XThR.Tn[1].n13 161.3
R22246 XThR.Tn[1].n82 XThR.Tn[1].t70 161.106
R22247 XThR.Tn[1].n77 XThR.Tn[1].t14 161.106
R22248 XThR.Tn[1].n72 XThR.Tn[1].t56 161.106
R22249 XThR.Tn[1].n67 XThR.Tn[1].t42 161.106
R22250 XThR.Tn[1].n62 XThR.Tn[1].t68 161.106
R22251 XThR.Tn[1].n57 XThR.Tn[1].t31 161.106
R22252 XThR.Tn[1].n52 XThR.Tn[1].t12 161.106
R22253 XThR.Tn[1].n47 XThR.Tn[1].t54 161.106
R22254 XThR.Tn[1].n42 XThR.Tn[1].t41 161.106
R22255 XThR.Tn[1].n37 XThR.Tn[1].t46 161.106
R22256 XThR.Tn[1].n32 XThR.Tn[1].t29 161.106
R22257 XThR.Tn[1].n27 XThR.Tn[1].t55 161.106
R22258 XThR.Tn[1].n22 XThR.Tn[1].t28 161.106
R22259 XThR.Tn[1].n17 XThR.Tn[1].t73 161.106
R22260 XThR.Tn[1].n12 XThR.Tn[1].t34 161.106
R22261 XThR.Tn[1].n10 XThR.Tn[1].t18 161.106
R22262 XThR.Tn[1].n83 XThR.Tn[1].t66 159.978
R22263 XThR.Tn[1].n78 XThR.Tn[1].t72 159.978
R22264 XThR.Tn[1].n73 XThR.Tn[1].t52 159.978
R22265 XThR.Tn[1].n68 XThR.Tn[1].t39 159.978
R22266 XThR.Tn[1].n63 XThR.Tn[1].t63 159.978
R22267 XThR.Tn[1].n58 XThR.Tn[1].t27 159.978
R22268 XThR.Tn[1].n53 XThR.Tn[1].t71 159.978
R22269 XThR.Tn[1].n48 XThR.Tn[1].t49 159.978
R22270 XThR.Tn[1].n43 XThR.Tn[1].t36 159.978
R22271 XThR.Tn[1].n38 XThR.Tn[1].t43 159.978
R22272 XThR.Tn[1].n33 XThR.Tn[1].t26 159.978
R22273 XThR.Tn[1].n28 XThR.Tn[1].t51 159.978
R22274 XThR.Tn[1].n23 XThR.Tn[1].t25 159.978
R22275 XThR.Tn[1].n18 XThR.Tn[1].t69 159.978
R22276 XThR.Tn[1].n13 XThR.Tn[1].t30 159.978
R22277 XThR.Tn[1].n82 XThR.Tn[1].t58 145.038
R22278 XThR.Tn[1].n77 XThR.Tn[1].t20 145.038
R22279 XThR.Tn[1].n72 XThR.Tn[1].t62 145.038
R22280 XThR.Tn[1].n67 XThR.Tn[1].t47 145.038
R22281 XThR.Tn[1].n62 XThR.Tn[1].t15 145.038
R22282 XThR.Tn[1].n57 XThR.Tn[1].t57 145.038
R22283 XThR.Tn[1].n52 XThR.Tn[1].t64 145.038
R22284 XThR.Tn[1].n47 XThR.Tn[1].t48 145.038
R22285 XThR.Tn[1].n42 XThR.Tn[1].t45 145.038
R22286 XThR.Tn[1].n37 XThR.Tn[1].t13 145.038
R22287 XThR.Tn[1].n32 XThR.Tn[1].t37 145.038
R22288 XThR.Tn[1].n27 XThR.Tn[1].t59 145.038
R22289 XThR.Tn[1].n22 XThR.Tn[1].t35 145.038
R22290 XThR.Tn[1].n17 XThR.Tn[1].t19 145.038
R22291 XThR.Tn[1].n12 XThR.Tn[1].t44 145.038
R22292 XThR.Tn[1].n10 XThR.Tn[1].t24 145.038
R22293 XThR.Tn[1].n83 XThR.Tn[1].t17 143.911
R22294 XThR.Tn[1].n78 XThR.Tn[1].t40 143.911
R22295 XThR.Tn[1].n73 XThR.Tn[1].t22 143.911
R22296 XThR.Tn[1].n68 XThR.Tn[1].t65 143.911
R22297 XThR.Tn[1].n63 XThR.Tn[1].t33 143.911
R22298 XThR.Tn[1].n58 XThR.Tn[1].t16 143.911
R22299 XThR.Tn[1].n53 XThR.Tn[1].t23 143.911
R22300 XThR.Tn[1].n48 XThR.Tn[1].t67 143.911
R22301 XThR.Tn[1].n43 XThR.Tn[1].t60 143.911
R22302 XThR.Tn[1].n38 XThR.Tn[1].t32 143.911
R22303 XThR.Tn[1].n33 XThR.Tn[1].t53 143.911
R22304 XThR.Tn[1].n28 XThR.Tn[1].t21 143.911
R22305 XThR.Tn[1].n23 XThR.Tn[1].t50 143.911
R22306 XThR.Tn[1].n18 XThR.Tn[1].t38 143.911
R22307 XThR.Tn[1].n13 XThR.Tn[1].t61 143.911
R22308 XThR.Tn[1].n7 XThR.Tn[1].n6 135.249
R22309 XThR.Tn[1].n9 XThR.Tn[1].n3 98.981
R22310 XThR.Tn[1].n8 XThR.Tn[1].n4 98.981
R22311 XThR.Tn[1].n7 XThR.Tn[1].n5 98.981
R22312 XThR.Tn[1].n9 XThR.Tn[1].n8 36.2672
R22313 XThR.Tn[1].n8 XThR.Tn[1].n7 36.2672
R22314 XThR.Tn[1].n88 XThR.Tn[1].n9 32.6405
R22315 XThR.Tn[1].n1 XThR.Tn[1].t7 26.5955
R22316 XThR.Tn[1].n1 XThR.Tn[1].t6 26.5955
R22317 XThR.Tn[1].n0 XThR.Tn[1].t4 26.5955
R22318 XThR.Tn[1].n0 XThR.Tn[1].t5 26.5955
R22319 XThR.Tn[1].n3 XThR.Tn[1].t11 24.9236
R22320 XThR.Tn[1].n3 XThR.Tn[1].t8 24.9236
R22321 XThR.Tn[1].n4 XThR.Tn[1].t10 24.9236
R22322 XThR.Tn[1].n4 XThR.Tn[1].t9 24.9236
R22323 XThR.Tn[1].n5 XThR.Tn[1].t2 24.9236
R22324 XThR.Tn[1].n5 XThR.Tn[1].t1 24.9236
R22325 XThR.Tn[1].n6 XThR.Tn[1].t3 24.9236
R22326 XThR.Tn[1].n6 XThR.Tn[1].t0 24.9236
R22327 XThR.Tn[1].n89 XThR.Tn[1].n2 18.5605
R22328 XThR.Tn[1].n89 XThR.Tn[1].n88 11.5205
R22329 XThR.Tn[1].n88 XThR.Tn[1] 6.42118
R22330 XThR.Tn[1] XThR.Tn[1].n11 5.34038
R22331 XThR.Tn[1].n16 XThR.Tn[1].n15 4.5005
R22332 XThR.Tn[1].n21 XThR.Tn[1].n20 4.5005
R22333 XThR.Tn[1].n26 XThR.Tn[1].n25 4.5005
R22334 XThR.Tn[1].n31 XThR.Tn[1].n30 4.5005
R22335 XThR.Tn[1].n36 XThR.Tn[1].n35 4.5005
R22336 XThR.Tn[1].n41 XThR.Tn[1].n40 4.5005
R22337 XThR.Tn[1].n46 XThR.Tn[1].n45 4.5005
R22338 XThR.Tn[1].n51 XThR.Tn[1].n50 4.5005
R22339 XThR.Tn[1].n56 XThR.Tn[1].n55 4.5005
R22340 XThR.Tn[1].n61 XThR.Tn[1].n60 4.5005
R22341 XThR.Tn[1].n66 XThR.Tn[1].n65 4.5005
R22342 XThR.Tn[1].n71 XThR.Tn[1].n70 4.5005
R22343 XThR.Tn[1].n76 XThR.Tn[1].n75 4.5005
R22344 XThR.Tn[1].n81 XThR.Tn[1].n80 4.5005
R22345 XThR.Tn[1].n86 XThR.Tn[1].n85 4.5005
R22346 XThR.Tn[1].n87 XThR.Tn[1] 3.70586
R22347 XThR.Tn[1].n16 XThR.Tn[1] 2.52282
R22348 XThR.Tn[1].n21 XThR.Tn[1] 2.52282
R22349 XThR.Tn[1].n26 XThR.Tn[1] 2.52282
R22350 XThR.Tn[1].n31 XThR.Tn[1] 2.52282
R22351 XThR.Tn[1].n36 XThR.Tn[1] 2.52282
R22352 XThR.Tn[1].n41 XThR.Tn[1] 2.52282
R22353 XThR.Tn[1].n46 XThR.Tn[1] 2.52282
R22354 XThR.Tn[1].n51 XThR.Tn[1] 2.52282
R22355 XThR.Tn[1].n56 XThR.Tn[1] 2.52282
R22356 XThR.Tn[1].n61 XThR.Tn[1] 2.52282
R22357 XThR.Tn[1].n66 XThR.Tn[1] 2.52282
R22358 XThR.Tn[1].n71 XThR.Tn[1] 2.52282
R22359 XThR.Tn[1].n76 XThR.Tn[1] 2.52282
R22360 XThR.Tn[1].n81 XThR.Tn[1] 2.52282
R22361 XThR.Tn[1].n86 XThR.Tn[1] 2.52282
R22362 XThR.Tn[1].n84 XThR.Tn[1] 1.08677
R22363 XThR.Tn[1].n79 XThR.Tn[1] 1.08677
R22364 XThR.Tn[1].n74 XThR.Tn[1] 1.08677
R22365 XThR.Tn[1].n69 XThR.Tn[1] 1.08677
R22366 XThR.Tn[1].n64 XThR.Tn[1] 1.08677
R22367 XThR.Tn[1].n59 XThR.Tn[1] 1.08677
R22368 XThR.Tn[1].n54 XThR.Tn[1] 1.08677
R22369 XThR.Tn[1].n49 XThR.Tn[1] 1.08677
R22370 XThR.Tn[1].n44 XThR.Tn[1] 1.08677
R22371 XThR.Tn[1].n39 XThR.Tn[1] 1.08677
R22372 XThR.Tn[1].n34 XThR.Tn[1] 1.08677
R22373 XThR.Tn[1].n29 XThR.Tn[1] 1.08677
R22374 XThR.Tn[1].n24 XThR.Tn[1] 1.08677
R22375 XThR.Tn[1].n19 XThR.Tn[1] 1.08677
R22376 XThR.Tn[1].n14 XThR.Tn[1] 1.08677
R22377 XThR.Tn[1] XThR.Tn[1].n16 0.839786
R22378 XThR.Tn[1] XThR.Tn[1].n21 0.839786
R22379 XThR.Tn[1] XThR.Tn[1].n26 0.839786
R22380 XThR.Tn[1] XThR.Tn[1].n31 0.839786
R22381 XThR.Tn[1] XThR.Tn[1].n36 0.839786
R22382 XThR.Tn[1] XThR.Tn[1].n41 0.839786
R22383 XThR.Tn[1] XThR.Tn[1].n46 0.839786
R22384 XThR.Tn[1] XThR.Tn[1].n51 0.839786
R22385 XThR.Tn[1] XThR.Tn[1].n56 0.839786
R22386 XThR.Tn[1] XThR.Tn[1].n61 0.839786
R22387 XThR.Tn[1] XThR.Tn[1].n66 0.839786
R22388 XThR.Tn[1] XThR.Tn[1].n71 0.839786
R22389 XThR.Tn[1] XThR.Tn[1].n76 0.839786
R22390 XThR.Tn[1] XThR.Tn[1].n81 0.839786
R22391 XThR.Tn[1] XThR.Tn[1].n86 0.839786
R22392 XThR.Tn[1] XThR.Tn[1].n89 0.6405
R22393 XThR.Tn[1].n11 XThR.Tn[1] 0.499542
R22394 XThR.Tn[1].n85 XThR.Tn[1] 0.063
R22395 XThR.Tn[1].n80 XThR.Tn[1] 0.063
R22396 XThR.Tn[1].n75 XThR.Tn[1] 0.063
R22397 XThR.Tn[1].n70 XThR.Tn[1] 0.063
R22398 XThR.Tn[1].n65 XThR.Tn[1] 0.063
R22399 XThR.Tn[1].n60 XThR.Tn[1] 0.063
R22400 XThR.Tn[1].n55 XThR.Tn[1] 0.063
R22401 XThR.Tn[1].n50 XThR.Tn[1] 0.063
R22402 XThR.Tn[1].n45 XThR.Tn[1] 0.063
R22403 XThR.Tn[1].n40 XThR.Tn[1] 0.063
R22404 XThR.Tn[1].n35 XThR.Tn[1] 0.063
R22405 XThR.Tn[1].n30 XThR.Tn[1] 0.063
R22406 XThR.Tn[1].n25 XThR.Tn[1] 0.063
R22407 XThR.Tn[1].n20 XThR.Tn[1] 0.063
R22408 XThR.Tn[1].n15 XThR.Tn[1] 0.063
R22409 XThR.Tn[1].n87 XThR.Tn[1] 0.0540714
R22410 XThR.Tn[1] XThR.Tn[1].n87 0.038
R22411 XThR.Tn[1].n11 XThR.Tn[1] 0.0143889
R22412 XThR.Tn[1].n85 XThR.Tn[1].n84 0.00771154
R22413 XThR.Tn[1].n80 XThR.Tn[1].n79 0.00771154
R22414 XThR.Tn[1].n75 XThR.Tn[1].n74 0.00771154
R22415 XThR.Tn[1].n70 XThR.Tn[1].n69 0.00771154
R22416 XThR.Tn[1].n65 XThR.Tn[1].n64 0.00771154
R22417 XThR.Tn[1].n60 XThR.Tn[1].n59 0.00771154
R22418 XThR.Tn[1].n55 XThR.Tn[1].n54 0.00771154
R22419 XThR.Tn[1].n50 XThR.Tn[1].n49 0.00771154
R22420 XThR.Tn[1].n45 XThR.Tn[1].n44 0.00771154
R22421 XThR.Tn[1].n40 XThR.Tn[1].n39 0.00771154
R22422 XThR.Tn[1].n35 XThR.Tn[1].n34 0.00771154
R22423 XThR.Tn[1].n30 XThR.Tn[1].n29 0.00771154
R22424 XThR.Tn[1].n25 XThR.Tn[1].n24 0.00771154
R22425 XThR.Tn[1].n20 XThR.Tn[1].n19 0.00771154
R22426 XThR.Tn[1].n15 XThR.Tn[1].n14 0.00771154
R22427 XThC.Tn[7].n5 XThC.Tn[7].n4 255.096
R22428 XThC.Tn[7].n2 XThC.Tn[7].n0 236.589
R22429 XThC.Tn[7].n5 XThC.Tn[7].n3 201.845
R22430 XThC.Tn[7].n2 XThC.Tn[7].n1 200.321
R22431 XThC.Tn[7].n67 XThC.Tn[7].n65 161.365
R22432 XThC.Tn[7].n63 XThC.Tn[7].n61 161.365
R22433 XThC.Tn[7].n59 XThC.Tn[7].n57 161.365
R22434 XThC.Tn[7].n55 XThC.Tn[7].n53 161.365
R22435 XThC.Tn[7].n51 XThC.Tn[7].n49 161.365
R22436 XThC.Tn[7].n47 XThC.Tn[7].n45 161.365
R22437 XThC.Tn[7].n43 XThC.Tn[7].n41 161.365
R22438 XThC.Tn[7].n39 XThC.Tn[7].n37 161.365
R22439 XThC.Tn[7].n35 XThC.Tn[7].n33 161.365
R22440 XThC.Tn[7].n31 XThC.Tn[7].n29 161.365
R22441 XThC.Tn[7].n27 XThC.Tn[7].n25 161.365
R22442 XThC.Tn[7].n23 XThC.Tn[7].n21 161.365
R22443 XThC.Tn[7].n19 XThC.Tn[7].n17 161.365
R22444 XThC.Tn[7].n15 XThC.Tn[7].n13 161.365
R22445 XThC.Tn[7].n11 XThC.Tn[7].n9 161.365
R22446 XThC.Tn[7].n8 XThC.Tn[7].n6 161.365
R22447 XThC.Tn[7].n65 XThC.Tn[7].t19 161.202
R22448 XThC.Tn[7].n61 XThC.Tn[7].t9 161.202
R22449 XThC.Tn[7].n57 XThC.Tn[7].t28 161.202
R22450 XThC.Tn[7].n53 XThC.Tn[7].t26 161.202
R22451 XThC.Tn[7].n49 XThC.Tn[7].t17 161.202
R22452 XThC.Tn[7].n45 XThC.Tn[7].t38 161.202
R22453 XThC.Tn[7].n41 XThC.Tn[7].t36 161.202
R22454 XThC.Tn[7].n37 XThC.Tn[7].t16 161.202
R22455 XThC.Tn[7].n33 XThC.Tn[7].t14 161.202
R22456 XThC.Tn[7].n29 XThC.Tn[7].t39 161.202
R22457 XThC.Tn[7].n25 XThC.Tn[7].t23 161.202
R22458 XThC.Tn[7].n21 XThC.Tn[7].t22 161.202
R22459 XThC.Tn[7].n17 XThC.Tn[7].t35 161.202
R22460 XThC.Tn[7].n13 XThC.Tn[7].t34 161.202
R22461 XThC.Tn[7].n9 XThC.Tn[7].t30 161.202
R22462 XThC.Tn[7].n6 XThC.Tn[7].t11 161.202
R22463 XThC.Tn[7].n65 XThC.Tn[7].t15 145.137
R22464 XThC.Tn[7].n61 XThC.Tn[7].t37 145.137
R22465 XThC.Tn[7].n57 XThC.Tn[7].t24 145.137
R22466 XThC.Tn[7].n53 XThC.Tn[7].t21 145.137
R22467 XThC.Tn[7].n49 XThC.Tn[7].t13 145.137
R22468 XThC.Tn[7].n45 XThC.Tn[7].t32 145.137
R22469 XThC.Tn[7].n41 XThC.Tn[7].t31 145.137
R22470 XThC.Tn[7].n37 XThC.Tn[7].t12 145.137
R22471 XThC.Tn[7].n33 XThC.Tn[7].t10 145.137
R22472 XThC.Tn[7].n29 XThC.Tn[7].t33 145.137
R22473 XThC.Tn[7].n25 XThC.Tn[7].t20 145.137
R22474 XThC.Tn[7].n21 XThC.Tn[7].t18 145.137
R22475 XThC.Tn[7].n17 XThC.Tn[7].t29 145.137
R22476 XThC.Tn[7].n13 XThC.Tn[7].t27 145.137
R22477 XThC.Tn[7].n9 XThC.Tn[7].t25 145.137
R22478 XThC.Tn[7].n6 XThC.Tn[7].t8 145.137
R22479 XThC.Tn[7].n4 XThC.Tn[7].t2 26.5955
R22480 XThC.Tn[7].n4 XThC.Tn[7].t1 26.5955
R22481 XThC.Tn[7].n3 XThC.Tn[7].t0 26.5955
R22482 XThC.Tn[7].n3 XThC.Tn[7].t3 26.5955
R22483 XThC.Tn[7] XThC.Tn[7].n5 26.4992
R22484 XThC.Tn[7].n0 XThC.Tn[7].t6 24.9236
R22485 XThC.Tn[7].n0 XThC.Tn[7].t5 24.9236
R22486 XThC.Tn[7].n1 XThC.Tn[7].t4 24.9236
R22487 XThC.Tn[7].n1 XThC.Tn[7].t7 24.9236
R22488 XThC.Tn[7].n70 XThC.Tn[7].n2 12.0894
R22489 XThC.Tn[7].n70 XThC.Tn[7] 9.64206
R22490 XThC.Tn[7].n69 XThC.Tn[7] 8.14595
R22491 XThC.Tn[7] XThC.Tn[7].n8 8.0245
R22492 XThC.Tn[7].n68 XThC.Tn[7].n67 7.9105
R22493 XThC.Tn[7].n64 XThC.Tn[7].n63 7.9105
R22494 XThC.Tn[7].n60 XThC.Tn[7].n59 7.9105
R22495 XThC.Tn[7].n56 XThC.Tn[7].n55 7.9105
R22496 XThC.Tn[7].n52 XThC.Tn[7].n51 7.9105
R22497 XThC.Tn[7].n48 XThC.Tn[7].n47 7.9105
R22498 XThC.Tn[7].n44 XThC.Tn[7].n43 7.9105
R22499 XThC.Tn[7].n40 XThC.Tn[7].n39 7.9105
R22500 XThC.Tn[7].n36 XThC.Tn[7].n35 7.9105
R22501 XThC.Tn[7].n32 XThC.Tn[7].n31 7.9105
R22502 XThC.Tn[7].n28 XThC.Tn[7].n27 7.9105
R22503 XThC.Tn[7].n24 XThC.Tn[7].n23 7.9105
R22504 XThC.Tn[7].n20 XThC.Tn[7].n19 7.9105
R22505 XThC.Tn[7].n16 XThC.Tn[7].n15 7.9105
R22506 XThC.Tn[7].n12 XThC.Tn[7].n11 7.9105
R22507 XThC.Tn[7].n69 XThC.Tn[7] 5.30358
R22508 XThC.Tn[7] XThC.Tn[7].n69 3.15894
R22509 XThC.Tn[7] XThC.Tn[7].n70 1.66284
R22510 XThC.Tn[7].n12 XThC.Tn[7] 0.235138
R22511 XThC.Tn[7].n16 XThC.Tn[7] 0.235138
R22512 XThC.Tn[7].n20 XThC.Tn[7] 0.235138
R22513 XThC.Tn[7].n24 XThC.Tn[7] 0.235138
R22514 XThC.Tn[7].n28 XThC.Tn[7] 0.235138
R22515 XThC.Tn[7].n32 XThC.Tn[7] 0.235138
R22516 XThC.Tn[7].n36 XThC.Tn[7] 0.235138
R22517 XThC.Tn[7].n40 XThC.Tn[7] 0.235138
R22518 XThC.Tn[7].n44 XThC.Tn[7] 0.235138
R22519 XThC.Tn[7].n48 XThC.Tn[7] 0.235138
R22520 XThC.Tn[7].n52 XThC.Tn[7] 0.235138
R22521 XThC.Tn[7].n56 XThC.Tn[7] 0.235138
R22522 XThC.Tn[7].n60 XThC.Tn[7] 0.235138
R22523 XThC.Tn[7].n64 XThC.Tn[7] 0.235138
R22524 XThC.Tn[7].n68 XThC.Tn[7] 0.235138
R22525 XThC.Tn[7] XThC.Tn[7].n12 0.114505
R22526 XThC.Tn[7] XThC.Tn[7].n16 0.114505
R22527 XThC.Tn[7] XThC.Tn[7].n20 0.114505
R22528 XThC.Tn[7] XThC.Tn[7].n24 0.114505
R22529 XThC.Tn[7] XThC.Tn[7].n28 0.114505
R22530 XThC.Tn[7] XThC.Tn[7].n32 0.114505
R22531 XThC.Tn[7] XThC.Tn[7].n36 0.114505
R22532 XThC.Tn[7] XThC.Tn[7].n40 0.114505
R22533 XThC.Tn[7] XThC.Tn[7].n44 0.114505
R22534 XThC.Tn[7] XThC.Tn[7].n48 0.114505
R22535 XThC.Tn[7] XThC.Tn[7].n52 0.114505
R22536 XThC.Tn[7] XThC.Tn[7].n56 0.114505
R22537 XThC.Tn[7] XThC.Tn[7].n60 0.114505
R22538 XThC.Tn[7] XThC.Tn[7].n64 0.114505
R22539 XThC.Tn[7] XThC.Tn[7].n68 0.114505
R22540 XThC.Tn[7].n67 XThC.Tn[7].n66 0.0599512
R22541 XThC.Tn[7].n63 XThC.Tn[7].n62 0.0599512
R22542 XThC.Tn[7].n59 XThC.Tn[7].n58 0.0599512
R22543 XThC.Tn[7].n55 XThC.Tn[7].n54 0.0599512
R22544 XThC.Tn[7].n51 XThC.Tn[7].n50 0.0599512
R22545 XThC.Tn[7].n47 XThC.Tn[7].n46 0.0599512
R22546 XThC.Tn[7].n43 XThC.Tn[7].n42 0.0599512
R22547 XThC.Tn[7].n39 XThC.Tn[7].n38 0.0599512
R22548 XThC.Tn[7].n35 XThC.Tn[7].n34 0.0599512
R22549 XThC.Tn[7].n31 XThC.Tn[7].n30 0.0599512
R22550 XThC.Tn[7].n27 XThC.Tn[7].n26 0.0599512
R22551 XThC.Tn[7].n23 XThC.Tn[7].n22 0.0599512
R22552 XThC.Tn[7].n19 XThC.Tn[7].n18 0.0599512
R22553 XThC.Tn[7].n15 XThC.Tn[7].n14 0.0599512
R22554 XThC.Tn[7].n11 XThC.Tn[7].n10 0.0599512
R22555 XThC.Tn[7].n8 XThC.Tn[7].n7 0.0599512
R22556 XThC.Tn[7].n66 XThC.Tn[7] 0.0469286
R22557 XThC.Tn[7].n62 XThC.Tn[7] 0.0469286
R22558 XThC.Tn[7].n58 XThC.Tn[7] 0.0469286
R22559 XThC.Tn[7].n54 XThC.Tn[7] 0.0469286
R22560 XThC.Tn[7].n50 XThC.Tn[7] 0.0469286
R22561 XThC.Tn[7].n46 XThC.Tn[7] 0.0469286
R22562 XThC.Tn[7].n42 XThC.Tn[7] 0.0469286
R22563 XThC.Tn[7].n38 XThC.Tn[7] 0.0469286
R22564 XThC.Tn[7].n34 XThC.Tn[7] 0.0469286
R22565 XThC.Tn[7].n30 XThC.Tn[7] 0.0469286
R22566 XThC.Tn[7].n26 XThC.Tn[7] 0.0469286
R22567 XThC.Tn[7].n22 XThC.Tn[7] 0.0469286
R22568 XThC.Tn[7].n18 XThC.Tn[7] 0.0469286
R22569 XThC.Tn[7].n14 XThC.Tn[7] 0.0469286
R22570 XThC.Tn[7].n10 XThC.Tn[7] 0.0469286
R22571 XThC.Tn[7].n7 XThC.Tn[7] 0.0469286
R22572 XThC.Tn[7].n66 XThC.Tn[7] 0.0401341
R22573 XThC.Tn[7].n62 XThC.Tn[7] 0.0401341
R22574 XThC.Tn[7].n58 XThC.Tn[7] 0.0401341
R22575 XThC.Tn[7].n54 XThC.Tn[7] 0.0401341
R22576 XThC.Tn[7].n50 XThC.Tn[7] 0.0401341
R22577 XThC.Tn[7].n46 XThC.Tn[7] 0.0401341
R22578 XThC.Tn[7].n42 XThC.Tn[7] 0.0401341
R22579 XThC.Tn[7].n38 XThC.Tn[7] 0.0401341
R22580 XThC.Tn[7].n34 XThC.Tn[7] 0.0401341
R22581 XThC.Tn[7].n30 XThC.Tn[7] 0.0401341
R22582 XThC.Tn[7].n26 XThC.Tn[7] 0.0401341
R22583 XThC.Tn[7].n22 XThC.Tn[7] 0.0401341
R22584 XThC.Tn[7].n18 XThC.Tn[7] 0.0401341
R22585 XThC.Tn[7].n14 XThC.Tn[7] 0.0401341
R22586 XThC.Tn[7].n10 XThC.Tn[7] 0.0401341
R22587 XThC.Tn[7].n7 XThC.Tn[7] 0.0401341
R22588 XThR.Tn[4].n2 XThR.Tn[4].n1 332.332
R22589 XThR.Tn[4].n2 XThR.Tn[4].n0 296.493
R22590 XThR.Tn[4] XThR.Tn[4].n82 161.363
R22591 XThR.Tn[4] XThR.Tn[4].n77 161.363
R22592 XThR.Tn[4] XThR.Tn[4].n72 161.363
R22593 XThR.Tn[4] XThR.Tn[4].n67 161.363
R22594 XThR.Tn[4] XThR.Tn[4].n62 161.363
R22595 XThR.Tn[4] XThR.Tn[4].n57 161.363
R22596 XThR.Tn[4] XThR.Tn[4].n52 161.363
R22597 XThR.Tn[4] XThR.Tn[4].n47 161.363
R22598 XThR.Tn[4] XThR.Tn[4].n42 161.363
R22599 XThR.Tn[4] XThR.Tn[4].n37 161.363
R22600 XThR.Tn[4] XThR.Tn[4].n32 161.363
R22601 XThR.Tn[4] XThR.Tn[4].n27 161.363
R22602 XThR.Tn[4] XThR.Tn[4].n22 161.363
R22603 XThR.Tn[4] XThR.Tn[4].n17 161.363
R22604 XThR.Tn[4] XThR.Tn[4].n12 161.363
R22605 XThR.Tn[4] XThR.Tn[4].n10 161.363
R22606 XThR.Tn[4].n84 XThR.Tn[4].n83 161.3
R22607 XThR.Tn[4].n79 XThR.Tn[4].n78 161.3
R22608 XThR.Tn[4].n74 XThR.Tn[4].n73 161.3
R22609 XThR.Tn[4].n69 XThR.Tn[4].n68 161.3
R22610 XThR.Tn[4].n64 XThR.Tn[4].n63 161.3
R22611 XThR.Tn[4].n59 XThR.Tn[4].n58 161.3
R22612 XThR.Tn[4].n54 XThR.Tn[4].n53 161.3
R22613 XThR.Tn[4].n49 XThR.Tn[4].n48 161.3
R22614 XThR.Tn[4].n44 XThR.Tn[4].n43 161.3
R22615 XThR.Tn[4].n39 XThR.Tn[4].n38 161.3
R22616 XThR.Tn[4].n34 XThR.Tn[4].n33 161.3
R22617 XThR.Tn[4].n29 XThR.Tn[4].n28 161.3
R22618 XThR.Tn[4].n24 XThR.Tn[4].n23 161.3
R22619 XThR.Tn[4].n19 XThR.Tn[4].n18 161.3
R22620 XThR.Tn[4].n14 XThR.Tn[4].n13 161.3
R22621 XThR.Tn[4].n82 XThR.Tn[4].t28 161.106
R22622 XThR.Tn[4].n77 XThR.Tn[4].t34 161.106
R22623 XThR.Tn[4].n72 XThR.Tn[4].t14 161.106
R22624 XThR.Tn[4].n67 XThR.Tn[4].t62 161.106
R22625 XThR.Tn[4].n62 XThR.Tn[4].t26 161.106
R22626 XThR.Tn[4].n57 XThR.Tn[4].t51 161.106
R22627 XThR.Tn[4].n52 XThR.Tn[4].t32 161.106
R22628 XThR.Tn[4].n47 XThR.Tn[4].t12 161.106
R22629 XThR.Tn[4].n42 XThR.Tn[4].t61 161.106
R22630 XThR.Tn[4].n37 XThR.Tn[4].t66 161.106
R22631 XThR.Tn[4].n32 XThR.Tn[4].t49 161.106
R22632 XThR.Tn[4].n27 XThR.Tn[4].t13 161.106
R22633 XThR.Tn[4].n22 XThR.Tn[4].t48 161.106
R22634 XThR.Tn[4].n17 XThR.Tn[4].t31 161.106
R22635 XThR.Tn[4].n12 XThR.Tn[4].t54 161.106
R22636 XThR.Tn[4].n10 XThR.Tn[4].t38 161.106
R22637 XThR.Tn[4].n83 XThR.Tn[4].t24 159.978
R22638 XThR.Tn[4].n78 XThR.Tn[4].t30 159.978
R22639 XThR.Tn[4].n73 XThR.Tn[4].t72 159.978
R22640 XThR.Tn[4].n68 XThR.Tn[4].t59 159.978
R22641 XThR.Tn[4].n63 XThR.Tn[4].t21 159.978
R22642 XThR.Tn[4].n58 XThR.Tn[4].t47 159.978
R22643 XThR.Tn[4].n53 XThR.Tn[4].t29 159.978
R22644 XThR.Tn[4].n48 XThR.Tn[4].t69 159.978
R22645 XThR.Tn[4].n43 XThR.Tn[4].t56 159.978
R22646 XThR.Tn[4].n38 XThR.Tn[4].t63 159.978
R22647 XThR.Tn[4].n33 XThR.Tn[4].t46 159.978
R22648 XThR.Tn[4].n28 XThR.Tn[4].t71 159.978
R22649 XThR.Tn[4].n23 XThR.Tn[4].t45 159.978
R22650 XThR.Tn[4].n18 XThR.Tn[4].t27 159.978
R22651 XThR.Tn[4].n13 XThR.Tn[4].t50 159.978
R22652 XThR.Tn[4].n82 XThR.Tn[4].t16 145.038
R22653 XThR.Tn[4].n77 XThR.Tn[4].t40 145.038
R22654 XThR.Tn[4].n72 XThR.Tn[4].t20 145.038
R22655 XThR.Tn[4].n67 XThR.Tn[4].t67 145.038
R22656 XThR.Tn[4].n62 XThR.Tn[4].t35 145.038
R22657 XThR.Tn[4].n57 XThR.Tn[4].t15 145.038
R22658 XThR.Tn[4].n52 XThR.Tn[4].t22 145.038
R22659 XThR.Tn[4].n47 XThR.Tn[4].t68 145.038
R22660 XThR.Tn[4].n42 XThR.Tn[4].t64 145.038
R22661 XThR.Tn[4].n37 XThR.Tn[4].t33 145.038
R22662 XThR.Tn[4].n32 XThR.Tn[4].t57 145.038
R22663 XThR.Tn[4].n27 XThR.Tn[4].t17 145.038
R22664 XThR.Tn[4].n22 XThR.Tn[4].t55 145.038
R22665 XThR.Tn[4].n17 XThR.Tn[4].t39 145.038
R22666 XThR.Tn[4].n12 XThR.Tn[4].t65 145.038
R22667 XThR.Tn[4].n10 XThR.Tn[4].t44 145.038
R22668 XThR.Tn[4].n83 XThR.Tn[4].t37 143.911
R22669 XThR.Tn[4].n78 XThR.Tn[4].t60 143.911
R22670 XThR.Tn[4].n73 XThR.Tn[4].t42 143.911
R22671 XThR.Tn[4].n68 XThR.Tn[4].t23 143.911
R22672 XThR.Tn[4].n63 XThR.Tn[4].t53 143.911
R22673 XThR.Tn[4].n58 XThR.Tn[4].t36 143.911
R22674 XThR.Tn[4].n53 XThR.Tn[4].t43 143.911
R22675 XThR.Tn[4].n48 XThR.Tn[4].t25 143.911
R22676 XThR.Tn[4].n43 XThR.Tn[4].t18 143.911
R22677 XThR.Tn[4].n38 XThR.Tn[4].t52 143.911
R22678 XThR.Tn[4].n33 XThR.Tn[4].t73 143.911
R22679 XThR.Tn[4].n28 XThR.Tn[4].t41 143.911
R22680 XThR.Tn[4].n23 XThR.Tn[4].t70 143.911
R22681 XThR.Tn[4].n18 XThR.Tn[4].t58 143.911
R22682 XThR.Tn[4].n13 XThR.Tn[4].t19 143.911
R22683 XThR.Tn[4].n7 XThR.Tn[4].n5 135.249
R22684 XThR.Tn[4].n9 XThR.Tn[4].n3 98.982
R22685 XThR.Tn[4].n8 XThR.Tn[4].n4 98.982
R22686 XThR.Tn[4].n7 XThR.Tn[4].n6 98.982
R22687 XThR.Tn[4].n9 XThR.Tn[4].n8 36.2672
R22688 XThR.Tn[4].n8 XThR.Tn[4].n7 36.2672
R22689 XThR.Tn[4].n88 XThR.Tn[4].n9 32.6405
R22690 XThR.Tn[4].n1 XThR.Tn[4].t4 26.5955
R22691 XThR.Tn[4].n1 XThR.Tn[4].t7 26.5955
R22692 XThR.Tn[4].n0 XThR.Tn[4].t5 26.5955
R22693 XThR.Tn[4].n0 XThR.Tn[4].t6 26.5955
R22694 XThR.Tn[4].n3 XThR.Tn[4].t11 24.9236
R22695 XThR.Tn[4].n3 XThR.Tn[4].t8 24.9236
R22696 XThR.Tn[4].n4 XThR.Tn[4].t10 24.9236
R22697 XThR.Tn[4].n4 XThR.Tn[4].t9 24.9236
R22698 XThR.Tn[4].n5 XThR.Tn[4].t0 24.9236
R22699 XThR.Tn[4].n5 XThR.Tn[4].t1 24.9236
R22700 XThR.Tn[4].n6 XThR.Tn[4].t3 24.9236
R22701 XThR.Tn[4].n6 XThR.Tn[4].t2 24.9236
R22702 XThR.Tn[4] XThR.Tn[4].n2 23.3605
R22703 XThR.Tn[4] XThR.Tn[4].n88 6.7205
R22704 XThR.Tn[4].n88 XThR.Tn[4] 5.80883
R22705 XThR.Tn[4] XThR.Tn[4].n11 5.34038
R22706 XThR.Tn[4].n16 XThR.Tn[4].n15 4.5005
R22707 XThR.Tn[4].n21 XThR.Tn[4].n20 4.5005
R22708 XThR.Tn[4].n26 XThR.Tn[4].n25 4.5005
R22709 XThR.Tn[4].n31 XThR.Tn[4].n30 4.5005
R22710 XThR.Tn[4].n36 XThR.Tn[4].n35 4.5005
R22711 XThR.Tn[4].n41 XThR.Tn[4].n40 4.5005
R22712 XThR.Tn[4].n46 XThR.Tn[4].n45 4.5005
R22713 XThR.Tn[4].n51 XThR.Tn[4].n50 4.5005
R22714 XThR.Tn[4].n56 XThR.Tn[4].n55 4.5005
R22715 XThR.Tn[4].n61 XThR.Tn[4].n60 4.5005
R22716 XThR.Tn[4].n66 XThR.Tn[4].n65 4.5005
R22717 XThR.Tn[4].n71 XThR.Tn[4].n70 4.5005
R22718 XThR.Tn[4].n76 XThR.Tn[4].n75 4.5005
R22719 XThR.Tn[4].n81 XThR.Tn[4].n80 4.5005
R22720 XThR.Tn[4].n86 XThR.Tn[4].n85 4.5005
R22721 XThR.Tn[4].n87 XThR.Tn[4] 3.70586
R22722 XThR.Tn[4].n16 XThR.Tn[4] 2.52282
R22723 XThR.Tn[4].n21 XThR.Tn[4] 2.52282
R22724 XThR.Tn[4].n26 XThR.Tn[4] 2.52282
R22725 XThR.Tn[4].n31 XThR.Tn[4] 2.52282
R22726 XThR.Tn[4].n36 XThR.Tn[4] 2.52282
R22727 XThR.Tn[4].n41 XThR.Tn[4] 2.52282
R22728 XThR.Tn[4].n46 XThR.Tn[4] 2.52282
R22729 XThR.Tn[4].n51 XThR.Tn[4] 2.52282
R22730 XThR.Tn[4].n56 XThR.Tn[4] 2.52282
R22731 XThR.Tn[4].n61 XThR.Tn[4] 2.52282
R22732 XThR.Tn[4].n66 XThR.Tn[4] 2.52282
R22733 XThR.Tn[4].n71 XThR.Tn[4] 2.52282
R22734 XThR.Tn[4].n76 XThR.Tn[4] 2.52282
R22735 XThR.Tn[4].n81 XThR.Tn[4] 2.52282
R22736 XThR.Tn[4].n86 XThR.Tn[4] 2.52282
R22737 XThR.Tn[4].n84 XThR.Tn[4] 1.08677
R22738 XThR.Tn[4].n79 XThR.Tn[4] 1.08677
R22739 XThR.Tn[4].n74 XThR.Tn[4] 1.08677
R22740 XThR.Tn[4].n69 XThR.Tn[4] 1.08677
R22741 XThR.Tn[4].n64 XThR.Tn[4] 1.08677
R22742 XThR.Tn[4].n59 XThR.Tn[4] 1.08677
R22743 XThR.Tn[4].n54 XThR.Tn[4] 1.08677
R22744 XThR.Tn[4].n49 XThR.Tn[4] 1.08677
R22745 XThR.Tn[4].n44 XThR.Tn[4] 1.08677
R22746 XThR.Tn[4].n39 XThR.Tn[4] 1.08677
R22747 XThR.Tn[4].n34 XThR.Tn[4] 1.08677
R22748 XThR.Tn[4].n29 XThR.Tn[4] 1.08677
R22749 XThR.Tn[4].n24 XThR.Tn[4] 1.08677
R22750 XThR.Tn[4].n19 XThR.Tn[4] 1.08677
R22751 XThR.Tn[4].n14 XThR.Tn[4] 1.08677
R22752 XThR.Tn[4] XThR.Tn[4].n16 0.839786
R22753 XThR.Tn[4] XThR.Tn[4].n21 0.839786
R22754 XThR.Tn[4] XThR.Tn[4].n26 0.839786
R22755 XThR.Tn[4] XThR.Tn[4].n31 0.839786
R22756 XThR.Tn[4] XThR.Tn[4].n36 0.839786
R22757 XThR.Tn[4] XThR.Tn[4].n41 0.839786
R22758 XThR.Tn[4] XThR.Tn[4].n46 0.839786
R22759 XThR.Tn[4] XThR.Tn[4].n51 0.839786
R22760 XThR.Tn[4] XThR.Tn[4].n56 0.839786
R22761 XThR.Tn[4] XThR.Tn[4].n61 0.839786
R22762 XThR.Tn[4] XThR.Tn[4].n66 0.839786
R22763 XThR.Tn[4] XThR.Tn[4].n71 0.839786
R22764 XThR.Tn[4] XThR.Tn[4].n76 0.839786
R22765 XThR.Tn[4] XThR.Tn[4].n81 0.839786
R22766 XThR.Tn[4] XThR.Tn[4].n86 0.839786
R22767 XThR.Tn[4].n11 XThR.Tn[4] 0.499542
R22768 XThR.Tn[4].n85 XThR.Tn[4] 0.063
R22769 XThR.Tn[4].n80 XThR.Tn[4] 0.063
R22770 XThR.Tn[4].n75 XThR.Tn[4] 0.063
R22771 XThR.Tn[4].n70 XThR.Tn[4] 0.063
R22772 XThR.Tn[4].n65 XThR.Tn[4] 0.063
R22773 XThR.Tn[4].n60 XThR.Tn[4] 0.063
R22774 XThR.Tn[4].n55 XThR.Tn[4] 0.063
R22775 XThR.Tn[4].n50 XThR.Tn[4] 0.063
R22776 XThR.Tn[4].n45 XThR.Tn[4] 0.063
R22777 XThR.Tn[4].n40 XThR.Tn[4] 0.063
R22778 XThR.Tn[4].n35 XThR.Tn[4] 0.063
R22779 XThR.Tn[4].n30 XThR.Tn[4] 0.063
R22780 XThR.Tn[4].n25 XThR.Tn[4] 0.063
R22781 XThR.Tn[4].n20 XThR.Tn[4] 0.063
R22782 XThR.Tn[4].n15 XThR.Tn[4] 0.063
R22783 XThR.Tn[4].n87 XThR.Tn[4] 0.0540714
R22784 XThR.Tn[4] XThR.Tn[4].n87 0.038
R22785 XThR.Tn[4].n11 XThR.Tn[4] 0.0143889
R22786 XThR.Tn[4].n85 XThR.Tn[4].n84 0.00771154
R22787 XThR.Tn[4].n80 XThR.Tn[4].n79 0.00771154
R22788 XThR.Tn[4].n75 XThR.Tn[4].n74 0.00771154
R22789 XThR.Tn[4].n70 XThR.Tn[4].n69 0.00771154
R22790 XThR.Tn[4].n65 XThR.Tn[4].n64 0.00771154
R22791 XThR.Tn[4].n60 XThR.Tn[4].n59 0.00771154
R22792 XThR.Tn[4].n55 XThR.Tn[4].n54 0.00771154
R22793 XThR.Tn[4].n50 XThR.Tn[4].n49 0.00771154
R22794 XThR.Tn[4].n45 XThR.Tn[4].n44 0.00771154
R22795 XThR.Tn[4].n40 XThR.Tn[4].n39 0.00771154
R22796 XThR.Tn[4].n35 XThR.Tn[4].n34 0.00771154
R22797 XThR.Tn[4].n30 XThR.Tn[4].n29 0.00771154
R22798 XThR.Tn[4].n25 XThR.Tn[4].n24 0.00771154
R22799 XThR.Tn[4].n20 XThR.Tn[4].n19 0.00771154
R22800 XThR.Tn[4].n15 XThR.Tn[4].n14 0.00771154
R22801 XThR.Tn[11].n8 XThR.Tn[11].n7 256.104
R22802 XThR.Tn[11].n5 XThR.Tn[11].n3 243.68
R22803 XThR.Tn[11].n2 XThR.Tn[11].n1 241.847
R22804 XThR.Tn[11].n5 XThR.Tn[11].n4 205.28
R22805 XThR.Tn[11].n8 XThR.Tn[11].n6 202.094
R22806 XThR.Tn[11].n2 XThR.Tn[11].n0 185
R22807 XThR.Tn[11] XThR.Tn[11].n82 161.363
R22808 XThR.Tn[11] XThR.Tn[11].n77 161.363
R22809 XThR.Tn[11] XThR.Tn[11].n72 161.363
R22810 XThR.Tn[11] XThR.Tn[11].n67 161.363
R22811 XThR.Tn[11] XThR.Tn[11].n62 161.363
R22812 XThR.Tn[11] XThR.Tn[11].n57 161.363
R22813 XThR.Tn[11] XThR.Tn[11].n52 161.363
R22814 XThR.Tn[11] XThR.Tn[11].n47 161.363
R22815 XThR.Tn[11] XThR.Tn[11].n42 161.363
R22816 XThR.Tn[11] XThR.Tn[11].n37 161.363
R22817 XThR.Tn[11] XThR.Tn[11].n32 161.363
R22818 XThR.Tn[11] XThR.Tn[11].n27 161.363
R22819 XThR.Tn[11] XThR.Tn[11].n22 161.363
R22820 XThR.Tn[11] XThR.Tn[11].n17 161.363
R22821 XThR.Tn[11] XThR.Tn[11].n12 161.363
R22822 XThR.Tn[11] XThR.Tn[11].n10 161.363
R22823 XThR.Tn[11].n84 XThR.Tn[11].n83 161.3
R22824 XThR.Tn[11].n79 XThR.Tn[11].n78 161.3
R22825 XThR.Tn[11].n74 XThR.Tn[11].n73 161.3
R22826 XThR.Tn[11].n69 XThR.Tn[11].n68 161.3
R22827 XThR.Tn[11].n64 XThR.Tn[11].n63 161.3
R22828 XThR.Tn[11].n59 XThR.Tn[11].n58 161.3
R22829 XThR.Tn[11].n54 XThR.Tn[11].n53 161.3
R22830 XThR.Tn[11].n49 XThR.Tn[11].n48 161.3
R22831 XThR.Tn[11].n44 XThR.Tn[11].n43 161.3
R22832 XThR.Tn[11].n39 XThR.Tn[11].n38 161.3
R22833 XThR.Tn[11].n34 XThR.Tn[11].n33 161.3
R22834 XThR.Tn[11].n29 XThR.Tn[11].n28 161.3
R22835 XThR.Tn[11].n24 XThR.Tn[11].n23 161.3
R22836 XThR.Tn[11].n19 XThR.Tn[11].n18 161.3
R22837 XThR.Tn[11].n14 XThR.Tn[11].n13 161.3
R22838 XThR.Tn[11].n82 XThR.Tn[11].t40 161.106
R22839 XThR.Tn[11].n77 XThR.Tn[11].t46 161.106
R22840 XThR.Tn[11].n72 XThR.Tn[11].t24 161.106
R22841 XThR.Tn[11].n67 XThR.Tn[11].t73 161.106
R22842 XThR.Tn[11].n62 XThR.Tn[11].t39 161.106
R22843 XThR.Tn[11].n57 XThR.Tn[11].t63 161.106
R22844 XThR.Tn[11].n52 XThR.Tn[11].t43 161.106
R22845 XThR.Tn[11].n47 XThR.Tn[11].t22 161.106
R22846 XThR.Tn[11].n42 XThR.Tn[11].t71 161.106
R22847 XThR.Tn[11].n37 XThR.Tn[11].t14 161.106
R22848 XThR.Tn[11].n32 XThR.Tn[11].t62 161.106
R22849 XThR.Tn[11].n27 XThR.Tn[11].t23 161.106
R22850 XThR.Tn[11].n22 XThR.Tn[11].t60 161.106
R22851 XThR.Tn[11].n17 XThR.Tn[11].t41 161.106
R22852 XThR.Tn[11].n12 XThR.Tn[11].t67 161.106
R22853 XThR.Tn[11].n10 XThR.Tn[11].t48 161.106
R22854 XThR.Tn[11].n83 XThR.Tn[11].t31 159.978
R22855 XThR.Tn[11].n78 XThR.Tn[11].t38 159.978
R22856 XThR.Tn[11].n73 XThR.Tn[11].t20 159.978
R22857 XThR.Tn[11].n68 XThR.Tn[11].t66 159.978
R22858 XThR.Tn[11].n63 XThR.Tn[11].t29 159.978
R22859 XThR.Tn[11].n58 XThR.Tn[11].t57 159.978
R22860 XThR.Tn[11].n53 XThR.Tn[11].t37 159.978
R22861 XThR.Tn[11].n48 XThR.Tn[11].t17 159.978
R22862 XThR.Tn[11].n43 XThR.Tn[11].t64 159.978
R22863 XThR.Tn[11].n38 XThR.Tn[11].t72 159.978
R22864 XThR.Tn[11].n33 XThR.Tn[11].t55 159.978
R22865 XThR.Tn[11].n28 XThR.Tn[11].t19 159.978
R22866 XThR.Tn[11].n23 XThR.Tn[11].t54 159.978
R22867 XThR.Tn[11].n18 XThR.Tn[11].t36 159.978
R22868 XThR.Tn[11].n13 XThR.Tn[11].t58 159.978
R22869 XThR.Tn[11].n82 XThR.Tn[11].t26 145.038
R22870 XThR.Tn[11].n77 XThR.Tn[11].t53 145.038
R22871 XThR.Tn[11].n72 XThR.Tn[11].t34 145.038
R22872 XThR.Tn[11].n67 XThR.Tn[11].t15 145.038
R22873 XThR.Tn[11].n62 XThR.Tn[11].t47 145.038
R22874 XThR.Tn[11].n57 XThR.Tn[11].t25 145.038
R22875 XThR.Tn[11].n52 XThR.Tn[11].t35 145.038
R22876 XThR.Tn[11].n47 XThR.Tn[11].t16 145.038
R22877 XThR.Tn[11].n42 XThR.Tn[11].t13 145.038
R22878 XThR.Tn[11].n37 XThR.Tn[11].t44 145.038
R22879 XThR.Tn[11].n32 XThR.Tn[11].t70 145.038
R22880 XThR.Tn[11].n27 XThR.Tn[11].t33 145.038
R22881 XThR.Tn[11].n22 XThR.Tn[11].t68 145.038
R22882 XThR.Tn[11].n17 XThR.Tn[11].t49 145.038
R22883 XThR.Tn[11].n12 XThR.Tn[11].t12 145.038
R22884 XThR.Tn[11].n10 XThR.Tn[11].t56 145.038
R22885 XThR.Tn[11].n83 XThR.Tn[11].t45 143.911
R22886 XThR.Tn[11].n78 XThR.Tn[11].t69 143.911
R22887 XThR.Tn[11].n73 XThR.Tn[11].t51 143.911
R22888 XThR.Tn[11].n68 XThR.Tn[11].t30 143.911
R22889 XThR.Tn[11].n63 XThR.Tn[11].t61 143.911
R22890 XThR.Tn[11].n58 XThR.Tn[11].t42 143.911
R22891 XThR.Tn[11].n53 XThR.Tn[11].t52 143.911
R22892 XThR.Tn[11].n48 XThR.Tn[11].t32 143.911
R22893 XThR.Tn[11].n43 XThR.Tn[11].t28 143.911
R22894 XThR.Tn[11].n38 XThR.Tn[11].t59 143.911
R22895 XThR.Tn[11].n33 XThR.Tn[11].t21 143.911
R22896 XThR.Tn[11].n28 XThR.Tn[11].t50 143.911
R22897 XThR.Tn[11].n23 XThR.Tn[11].t18 143.911
R22898 XThR.Tn[11].n18 XThR.Tn[11].t65 143.911
R22899 XThR.Tn[11].n13 XThR.Tn[11].t27 143.911
R22900 XThR.Tn[11] XThR.Tn[11].n5 35.7652
R22901 XThR.Tn[11].n6 XThR.Tn[11].t3 26.5955
R22902 XThR.Tn[11].n6 XThR.Tn[11].t9 26.5955
R22903 XThR.Tn[11].n7 XThR.Tn[11].t1 26.5955
R22904 XThR.Tn[11].n7 XThR.Tn[11].t8 26.5955
R22905 XThR.Tn[11].n3 XThR.Tn[11].t4 26.5955
R22906 XThR.Tn[11].n3 XThR.Tn[11].t6 26.5955
R22907 XThR.Tn[11].n4 XThR.Tn[11].t5 26.5955
R22908 XThR.Tn[11].n4 XThR.Tn[11].t7 26.5955
R22909 XThR.Tn[11].n0 XThR.Tn[11].t11 24.9236
R22910 XThR.Tn[11].n0 XThR.Tn[11].t2 24.9236
R22911 XThR.Tn[11].n1 XThR.Tn[11].t10 24.9236
R22912 XThR.Tn[11].n1 XThR.Tn[11].t0 24.9236
R22913 XThR.Tn[11] XThR.Tn[11].n2 22.9615
R22914 XThR.Tn[11].n9 XThR.Tn[11].n8 13.5534
R22915 XThR.Tn[11].n88 XThR.Tn[11] 8.41462
R22916 XThR.Tn[11] XThR.Tn[11].n11 5.34038
R22917 XThR.Tn[11].n16 XThR.Tn[11].n15 4.5005
R22918 XThR.Tn[11].n21 XThR.Tn[11].n20 4.5005
R22919 XThR.Tn[11].n26 XThR.Tn[11].n25 4.5005
R22920 XThR.Tn[11].n31 XThR.Tn[11].n30 4.5005
R22921 XThR.Tn[11].n36 XThR.Tn[11].n35 4.5005
R22922 XThR.Tn[11].n41 XThR.Tn[11].n40 4.5005
R22923 XThR.Tn[11].n46 XThR.Tn[11].n45 4.5005
R22924 XThR.Tn[11].n51 XThR.Tn[11].n50 4.5005
R22925 XThR.Tn[11].n56 XThR.Tn[11].n55 4.5005
R22926 XThR.Tn[11].n61 XThR.Tn[11].n60 4.5005
R22927 XThR.Tn[11].n66 XThR.Tn[11].n65 4.5005
R22928 XThR.Tn[11].n71 XThR.Tn[11].n70 4.5005
R22929 XThR.Tn[11].n76 XThR.Tn[11].n75 4.5005
R22930 XThR.Tn[11].n81 XThR.Tn[11].n80 4.5005
R22931 XThR.Tn[11].n86 XThR.Tn[11].n85 4.5005
R22932 XThR.Tn[11].n87 XThR.Tn[11] 3.70586
R22933 XThR.Tn[11].n88 XThR.Tn[11].n9 2.99115
R22934 XThR.Tn[11].n9 XThR.Tn[11] 2.87153
R22935 XThR.Tn[11].n16 XThR.Tn[11] 2.52282
R22936 XThR.Tn[11].n21 XThR.Tn[11] 2.52282
R22937 XThR.Tn[11].n26 XThR.Tn[11] 2.52282
R22938 XThR.Tn[11].n31 XThR.Tn[11] 2.52282
R22939 XThR.Tn[11].n36 XThR.Tn[11] 2.52282
R22940 XThR.Tn[11].n41 XThR.Tn[11] 2.52282
R22941 XThR.Tn[11].n46 XThR.Tn[11] 2.52282
R22942 XThR.Tn[11].n51 XThR.Tn[11] 2.52282
R22943 XThR.Tn[11].n56 XThR.Tn[11] 2.52282
R22944 XThR.Tn[11].n61 XThR.Tn[11] 2.52282
R22945 XThR.Tn[11].n66 XThR.Tn[11] 2.52282
R22946 XThR.Tn[11].n71 XThR.Tn[11] 2.52282
R22947 XThR.Tn[11].n76 XThR.Tn[11] 2.52282
R22948 XThR.Tn[11].n81 XThR.Tn[11] 2.52282
R22949 XThR.Tn[11].n86 XThR.Tn[11] 2.52282
R22950 XThR.Tn[11] XThR.Tn[11].n88 2.2734
R22951 XThR.Tn[11].n9 XThR.Tn[11] 1.50638
R22952 XThR.Tn[11].n84 XThR.Tn[11] 1.08677
R22953 XThR.Tn[11].n79 XThR.Tn[11] 1.08677
R22954 XThR.Tn[11].n74 XThR.Tn[11] 1.08677
R22955 XThR.Tn[11].n69 XThR.Tn[11] 1.08677
R22956 XThR.Tn[11].n64 XThR.Tn[11] 1.08677
R22957 XThR.Tn[11].n59 XThR.Tn[11] 1.08677
R22958 XThR.Tn[11].n54 XThR.Tn[11] 1.08677
R22959 XThR.Tn[11].n49 XThR.Tn[11] 1.08677
R22960 XThR.Tn[11].n44 XThR.Tn[11] 1.08677
R22961 XThR.Tn[11].n39 XThR.Tn[11] 1.08677
R22962 XThR.Tn[11].n34 XThR.Tn[11] 1.08677
R22963 XThR.Tn[11].n29 XThR.Tn[11] 1.08677
R22964 XThR.Tn[11].n24 XThR.Tn[11] 1.08677
R22965 XThR.Tn[11].n19 XThR.Tn[11] 1.08677
R22966 XThR.Tn[11].n14 XThR.Tn[11] 1.08677
R22967 XThR.Tn[11] XThR.Tn[11].n16 0.839786
R22968 XThR.Tn[11] XThR.Tn[11].n21 0.839786
R22969 XThR.Tn[11] XThR.Tn[11].n26 0.839786
R22970 XThR.Tn[11] XThR.Tn[11].n31 0.839786
R22971 XThR.Tn[11] XThR.Tn[11].n36 0.839786
R22972 XThR.Tn[11] XThR.Tn[11].n41 0.839786
R22973 XThR.Tn[11] XThR.Tn[11].n46 0.839786
R22974 XThR.Tn[11] XThR.Tn[11].n51 0.839786
R22975 XThR.Tn[11] XThR.Tn[11].n56 0.839786
R22976 XThR.Tn[11] XThR.Tn[11].n61 0.839786
R22977 XThR.Tn[11] XThR.Tn[11].n66 0.839786
R22978 XThR.Tn[11] XThR.Tn[11].n71 0.839786
R22979 XThR.Tn[11] XThR.Tn[11].n76 0.839786
R22980 XThR.Tn[11] XThR.Tn[11].n81 0.839786
R22981 XThR.Tn[11] XThR.Tn[11].n86 0.839786
R22982 XThR.Tn[11].n11 XThR.Tn[11] 0.499542
R22983 XThR.Tn[11].n85 XThR.Tn[11] 0.063
R22984 XThR.Tn[11].n80 XThR.Tn[11] 0.063
R22985 XThR.Tn[11].n75 XThR.Tn[11] 0.063
R22986 XThR.Tn[11].n70 XThR.Tn[11] 0.063
R22987 XThR.Tn[11].n65 XThR.Tn[11] 0.063
R22988 XThR.Tn[11].n60 XThR.Tn[11] 0.063
R22989 XThR.Tn[11].n55 XThR.Tn[11] 0.063
R22990 XThR.Tn[11].n50 XThR.Tn[11] 0.063
R22991 XThR.Tn[11].n45 XThR.Tn[11] 0.063
R22992 XThR.Tn[11].n40 XThR.Tn[11] 0.063
R22993 XThR.Tn[11].n35 XThR.Tn[11] 0.063
R22994 XThR.Tn[11].n30 XThR.Tn[11] 0.063
R22995 XThR.Tn[11].n25 XThR.Tn[11] 0.063
R22996 XThR.Tn[11].n20 XThR.Tn[11] 0.063
R22997 XThR.Tn[11].n15 XThR.Tn[11] 0.063
R22998 XThR.Tn[11].n87 XThR.Tn[11] 0.0540714
R22999 XThR.Tn[11] XThR.Tn[11].n87 0.038
R23000 XThR.Tn[11].n11 XThR.Tn[11] 0.0143889
R23001 XThR.Tn[11].n85 XThR.Tn[11].n84 0.00771154
R23002 XThR.Tn[11].n80 XThR.Tn[11].n79 0.00771154
R23003 XThR.Tn[11].n75 XThR.Tn[11].n74 0.00771154
R23004 XThR.Tn[11].n70 XThR.Tn[11].n69 0.00771154
R23005 XThR.Tn[11].n65 XThR.Tn[11].n64 0.00771154
R23006 XThR.Tn[11].n60 XThR.Tn[11].n59 0.00771154
R23007 XThR.Tn[11].n55 XThR.Tn[11].n54 0.00771154
R23008 XThR.Tn[11].n50 XThR.Tn[11].n49 0.00771154
R23009 XThR.Tn[11].n45 XThR.Tn[11].n44 0.00771154
R23010 XThR.Tn[11].n40 XThR.Tn[11].n39 0.00771154
R23011 XThR.Tn[11].n35 XThR.Tn[11].n34 0.00771154
R23012 XThR.Tn[11].n30 XThR.Tn[11].n29 0.00771154
R23013 XThR.Tn[11].n25 XThR.Tn[11].n24 0.00771154
R23014 XThR.Tn[11].n20 XThR.Tn[11].n19 0.00771154
R23015 XThR.Tn[11].n15 XThR.Tn[11].n14 0.00771154
R23016 XThR.Tn[7].n5 XThR.Tn[7].n3 244.067
R23017 XThR.Tn[7].n2 XThR.Tn[7].n0 236.589
R23018 XThR.Tn[7].n5 XThR.Tn[7].n4 204.893
R23019 XThR.Tn[7].n2 XThR.Tn[7].n1 200.321
R23020 XThR.Tn[7] XThR.Tn[7].n79 161.363
R23021 XThR.Tn[7] XThR.Tn[7].n74 161.363
R23022 XThR.Tn[7] XThR.Tn[7].n69 161.363
R23023 XThR.Tn[7] XThR.Tn[7].n64 161.363
R23024 XThR.Tn[7] XThR.Tn[7].n59 161.363
R23025 XThR.Tn[7] XThR.Tn[7].n54 161.363
R23026 XThR.Tn[7] XThR.Tn[7].n49 161.363
R23027 XThR.Tn[7] XThR.Tn[7].n44 161.363
R23028 XThR.Tn[7] XThR.Tn[7].n39 161.363
R23029 XThR.Tn[7] XThR.Tn[7].n34 161.363
R23030 XThR.Tn[7] XThR.Tn[7].n29 161.363
R23031 XThR.Tn[7] XThR.Tn[7].n24 161.363
R23032 XThR.Tn[7] XThR.Tn[7].n19 161.363
R23033 XThR.Tn[7] XThR.Tn[7].n14 161.363
R23034 XThR.Tn[7] XThR.Tn[7].n9 161.363
R23035 XThR.Tn[7] XThR.Tn[7].n7 161.363
R23036 XThR.Tn[7].n81 XThR.Tn[7].n80 161.3
R23037 XThR.Tn[7].n76 XThR.Tn[7].n75 161.3
R23038 XThR.Tn[7].n71 XThR.Tn[7].n70 161.3
R23039 XThR.Tn[7].n66 XThR.Tn[7].n65 161.3
R23040 XThR.Tn[7].n61 XThR.Tn[7].n60 161.3
R23041 XThR.Tn[7].n56 XThR.Tn[7].n55 161.3
R23042 XThR.Tn[7].n51 XThR.Tn[7].n50 161.3
R23043 XThR.Tn[7].n46 XThR.Tn[7].n45 161.3
R23044 XThR.Tn[7].n41 XThR.Tn[7].n40 161.3
R23045 XThR.Tn[7].n36 XThR.Tn[7].n35 161.3
R23046 XThR.Tn[7].n31 XThR.Tn[7].n30 161.3
R23047 XThR.Tn[7].n26 XThR.Tn[7].n25 161.3
R23048 XThR.Tn[7].n21 XThR.Tn[7].n20 161.3
R23049 XThR.Tn[7].n16 XThR.Tn[7].n15 161.3
R23050 XThR.Tn[7].n11 XThR.Tn[7].n10 161.3
R23051 XThR.Tn[7].n79 XThR.Tn[7].t35 161.106
R23052 XThR.Tn[7].n74 XThR.Tn[7].t41 161.106
R23053 XThR.Tn[7].n69 XThR.Tn[7].t22 161.106
R23054 XThR.Tn[7].n64 XThR.Tn[7].t69 161.106
R23055 XThR.Tn[7].n59 XThR.Tn[7].t33 161.106
R23056 XThR.Tn[7].n54 XThR.Tn[7].t57 161.106
R23057 XThR.Tn[7].n49 XThR.Tn[7].t39 161.106
R23058 XThR.Tn[7].n44 XThR.Tn[7].t20 161.106
R23059 XThR.Tn[7].n39 XThR.Tn[7].t68 161.106
R23060 XThR.Tn[7].n34 XThR.Tn[7].t11 161.106
R23061 XThR.Tn[7].n29 XThR.Tn[7].t56 161.106
R23062 XThR.Tn[7].n24 XThR.Tn[7].t21 161.106
R23063 XThR.Tn[7].n19 XThR.Tn[7].t55 161.106
R23064 XThR.Tn[7].n14 XThR.Tn[7].t37 161.106
R23065 XThR.Tn[7].n9 XThR.Tn[7].t60 161.106
R23066 XThR.Tn[7].n7 XThR.Tn[7].t45 161.106
R23067 XThR.Tn[7].n80 XThR.Tn[7].t13 159.978
R23068 XThR.Tn[7].n75 XThR.Tn[7].t17 159.978
R23069 XThR.Tn[7].n70 XThR.Tn[7].t64 159.978
R23070 XThR.Tn[7].n65 XThR.Tn[7].t48 159.978
R23071 XThR.Tn[7].n60 XThR.Tn[7].t10 159.978
R23072 XThR.Tn[7].n55 XThR.Tn[7].t36 159.978
R23073 XThR.Tn[7].n50 XThR.Tn[7].t16 159.978
R23074 XThR.Tn[7].n45 XThR.Tn[7].t61 159.978
R23075 XThR.Tn[7].n40 XThR.Tn[7].t46 159.978
R23076 XThR.Tn[7].n35 XThR.Tn[7].t54 159.978
R23077 XThR.Tn[7].n30 XThR.Tn[7].t34 159.978
R23078 XThR.Tn[7].n25 XThR.Tn[7].t63 159.978
R23079 XThR.Tn[7].n20 XThR.Tn[7].t32 159.978
R23080 XThR.Tn[7].n15 XThR.Tn[7].t15 159.978
R23081 XThR.Tn[7].n10 XThR.Tn[7].t38 159.978
R23082 XThR.Tn[7].n79 XThR.Tn[7].t24 145.038
R23083 XThR.Tn[7].n74 XThR.Tn[7].t49 145.038
R23084 XThR.Tn[7].n69 XThR.Tn[7].t28 145.038
R23085 XThR.Tn[7].n64 XThR.Tn[7].t12 145.038
R23086 XThR.Tn[7].n59 XThR.Tn[7].t42 145.038
R23087 XThR.Tn[7].n54 XThR.Tn[7].t23 145.038
R23088 XThR.Tn[7].n49 XThR.Tn[7].t29 145.038
R23089 XThR.Tn[7].n44 XThR.Tn[7].t14 145.038
R23090 XThR.Tn[7].n39 XThR.Tn[7].t9 145.038
R23091 XThR.Tn[7].n34 XThR.Tn[7].t40 145.038
R23092 XThR.Tn[7].n29 XThR.Tn[7].t65 145.038
R23093 XThR.Tn[7].n24 XThR.Tn[7].t25 145.038
R23094 XThR.Tn[7].n19 XThR.Tn[7].t62 145.038
R23095 XThR.Tn[7].n14 XThR.Tn[7].t47 145.038
R23096 XThR.Tn[7].n9 XThR.Tn[7].t8 145.038
R23097 XThR.Tn[7].n7 XThR.Tn[7].t53 145.038
R23098 XThR.Tn[7].n80 XThR.Tn[7].t44 143.911
R23099 XThR.Tn[7].n75 XThR.Tn[7].t67 143.911
R23100 XThR.Tn[7].n70 XThR.Tn[7].t51 143.911
R23101 XThR.Tn[7].n65 XThR.Tn[7].t30 143.911
R23102 XThR.Tn[7].n60 XThR.Tn[7].t59 143.911
R23103 XThR.Tn[7].n55 XThR.Tn[7].t43 143.911
R23104 XThR.Tn[7].n50 XThR.Tn[7].t52 143.911
R23105 XThR.Tn[7].n45 XThR.Tn[7].t31 143.911
R23106 XThR.Tn[7].n40 XThR.Tn[7].t27 143.911
R23107 XThR.Tn[7].n35 XThR.Tn[7].t58 143.911
R23108 XThR.Tn[7].n30 XThR.Tn[7].t19 143.911
R23109 XThR.Tn[7].n25 XThR.Tn[7].t50 143.911
R23110 XThR.Tn[7].n20 XThR.Tn[7].t18 143.911
R23111 XThR.Tn[7].n15 XThR.Tn[7].t66 143.911
R23112 XThR.Tn[7].n10 XThR.Tn[7].t26 143.911
R23113 XThR.Tn[7].n4 XThR.Tn[7].t1 26.5955
R23114 XThR.Tn[7].n4 XThR.Tn[7].t0 26.5955
R23115 XThR.Tn[7].n3 XThR.Tn[7].t2 26.5955
R23116 XThR.Tn[7].n3 XThR.Tn[7].t3 26.5955
R23117 XThR.Tn[7].n0 XThR.Tn[7].t7 24.9236
R23118 XThR.Tn[7].n0 XThR.Tn[7].t4 24.9236
R23119 XThR.Tn[7].n1 XThR.Tn[7].t6 24.9236
R23120 XThR.Tn[7].n1 XThR.Tn[7].t5 24.9236
R23121 XThR.Tn[7] XThR.Tn[7].n2 16.079
R23122 XThR.Tn[7].n6 XThR.Tn[7].n5 11.4531
R23123 XThR.Tn[7] XThR.Tn[7].n6 10.4732
R23124 XThR.Tn[7] XThR.Tn[7].n85 8.81089
R23125 XThR.Tn[7] XThR.Tn[7].n8 5.34038
R23126 XThR.Tn[7].n85 XThR.Tn[7] 5.25732
R23127 XThR.Tn[7].n13 XThR.Tn[7].n12 4.5005
R23128 XThR.Tn[7].n18 XThR.Tn[7].n17 4.5005
R23129 XThR.Tn[7].n23 XThR.Tn[7].n22 4.5005
R23130 XThR.Tn[7].n28 XThR.Tn[7].n27 4.5005
R23131 XThR.Tn[7].n33 XThR.Tn[7].n32 4.5005
R23132 XThR.Tn[7].n38 XThR.Tn[7].n37 4.5005
R23133 XThR.Tn[7].n43 XThR.Tn[7].n42 4.5005
R23134 XThR.Tn[7].n48 XThR.Tn[7].n47 4.5005
R23135 XThR.Tn[7].n53 XThR.Tn[7].n52 4.5005
R23136 XThR.Tn[7].n58 XThR.Tn[7].n57 4.5005
R23137 XThR.Tn[7].n63 XThR.Tn[7].n62 4.5005
R23138 XThR.Tn[7].n68 XThR.Tn[7].n67 4.5005
R23139 XThR.Tn[7].n73 XThR.Tn[7].n72 4.5005
R23140 XThR.Tn[7].n78 XThR.Tn[7].n77 4.5005
R23141 XThR.Tn[7].n83 XThR.Tn[7].n82 4.5005
R23142 XThR.Tn[7].n84 XThR.Tn[7] 3.70586
R23143 XThR.Tn[7].n13 XThR.Tn[7] 2.52282
R23144 XThR.Tn[7].n18 XThR.Tn[7] 2.52282
R23145 XThR.Tn[7].n23 XThR.Tn[7] 2.52282
R23146 XThR.Tn[7].n28 XThR.Tn[7] 2.52282
R23147 XThR.Tn[7].n33 XThR.Tn[7] 2.52282
R23148 XThR.Tn[7].n38 XThR.Tn[7] 2.52282
R23149 XThR.Tn[7].n43 XThR.Tn[7] 2.52282
R23150 XThR.Tn[7].n48 XThR.Tn[7] 2.52282
R23151 XThR.Tn[7].n53 XThR.Tn[7] 2.52282
R23152 XThR.Tn[7].n58 XThR.Tn[7] 2.52282
R23153 XThR.Tn[7].n63 XThR.Tn[7] 2.52282
R23154 XThR.Tn[7].n68 XThR.Tn[7] 2.52282
R23155 XThR.Tn[7].n73 XThR.Tn[7] 2.52282
R23156 XThR.Tn[7].n78 XThR.Tn[7] 2.52282
R23157 XThR.Tn[7].n83 XThR.Tn[7] 2.52282
R23158 XThR.Tn[7].n85 XThR.Tn[7] 2.49401
R23159 XThR.Tn[7].n81 XThR.Tn[7] 1.08677
R23160 XThR.Tn[7].n76 XThR.Tn[7] 1.08677
R23161 XThR.Tn[7].n71 XThR.Tn[7] 1.08677
R23162 XThR.Tn[7].n66 XThR.Tn[7] 1.08677
R23163 XThR.Tn[7].n61 XThR.Tn[7] 1.08677
R23164 XThR.Tn[7].n56 XThR.Tn[7] 1.08677
R23165 XThR.Tn[7].n51 XThR.Tn[7] 1.08677
R23166 XThR.Tn[7].n46 XThR.Tn[7] 1.08677
R23167 XThR.Tn[7].n41 XThR.Tn[7] 1.08677
R23168 XThR.Tn[7].n36 XThR.Tn[7] 1.08677
R23169 XThR.Tn[7].n31 XThR.Tn[7] 1.08677
R23170 XThR.Tn[7].n26 XThR.Tn[7] 1.08677
R23171 XThR.Tn[7].n21 XThR.Tn[7] 1.08677
R23172 XThR.Tn[7].n16 XThR.Tn[7] 1.08677
R23173 XThR.Tn[7].n11 XThR.Tn[7] 1.08677
R23174 XThR.Tn[7] XThR.Tn[7].n13 0.839786
R23175 XThR.Tn[7] XThR.Tn[7].n18 0.839786
R23176 XThR.Tn[7] XThR.Tn[7].n23 0.839786
R23177 XThR.Tn[7] XThR.Tn[7].n28 0.839786
R23178 XThR.Tn[7] XThR.Tn[7].n33 0.839786
R23179 XThR.Tn[7] XThR.Tn[7].n38 0.839786
R23180 XThR.Tn[7] XThR.Tn[7].n43 0.839786
R23181 XThR.Tn[7] XThR.Tn[7].n48 0.839786
R23182 XThR.Tn[7] XThR.Tn[7].n53 0.839786
R23183 XThR.Tn[7] XThR.Tn[7].n58 0.839786
R23184 XThR.Tn[7] XThR.Tn[7].n63 0.839786
R23185 XThR.Tn[7] XThR.Tn[7].n68 0.839786
R23186 XThR.Tn[7] XThR.Tn[7].n73 0.839786
R23187 XThR.Tn[7] XThR.Tn[7].n78 0.839786
R23188 XThR.Tn[7] XThR.Tn[7].n83 0.839786
R23189 XThR.Tn[7].n6 XThR.Tn[7] 0.830612
R23190 XThR.Tn[7].n8 XThR.Tn[7] 0.499542
R23191 XThR.Tn[7].n82 XThR.Tn[7] 0.063
R23192 XThR.Tn[7].n77 XThR.Tn[7] 0.063
R23193 XThR.Tn[7].n72 XThR.Tn[7] 0.063
R23194 XThR.Tn[7].n67 XThR.Tn[7] 0.063
R23195 XThR.Tn[7].n62 XThR.Tn[7] 0.063
R23196 XThR.Tn[7].n57 XThR.Tn[7] 0.063
R23197 XThR.Tn[7].n52 XThR.Tn[7] 0.063
R23198 XThR.Tn[7].n47 XThR.Tn[7] 0.063
R23199 XThR.Tn[7].n42 XThR.Tn[7] 0.063
R23200 XThR.Tn[7].n37 XThR.Tn[7] 0.063
R23201 XThR.Tn[7].n32 XThR.Tn[7] 0.063
R23202 XThR.Tn[7].n27 XThR.Tn[7] 0.063
R23203 XThR.Tn[7].n22 XThR.Tn[7] 0.063
R23204 XThR.Tn[7].n17 XThR.Tn[7] 0.063
R23205 XThR.Tn[7].n12 XThR.Tn[7] 0.063
R23206 XThR.Tn[7].n84 XThR.Tn[7] 0.0540714
R23207 XThR.Tn[7] XThR.Tn[7].n84 0.038
R23208 XThR.Tn[7].n8 XThR.Tn[7] 0.0143889
R23209 XThR.Tn[7].n82 XThR.Tn[7].n81 0.00771154
R23210 XThR.Tn[7].n77 XThR.Tn[7].n76 0.00771154
R23211 XThR.Tn[7].n72 XThR.Tn[7].n71 0.00771154
R23212 XThR.Tn[7].n67 XThR.Tn[7].n66 0.00771154
R23213 XThR.Tn[7].n62 XThR.Tn[7].n61 0.00771154
R23214 XThR.Tn[7].n57 XThR.Tn[7].n56 0.00771154
R23215 XThR.Tn[7].n52 XThR.Tn[7].n51 0.00771154
R23216 XThR.Tn[7].n47 XThR.Tn[7].n46 0.00771154
R23217 XThR.Tn[7].n42 XThR.Tn[7].n41 0.00771154
R23218 XThR.Tn[7].n37 XThR.Tn[7].n36 0.00771154
R23219 XThR.Tn[7].n32 XThR.Tn[7].n31 0.00771154
R23220 XThR.Tn[7].n27 XThR.Tn[7].n26 0.00771154
R23221 XThR.Tn[7].n22 XThR.Tn[7].n21 0.00771154
R23222 XThR.Tn[7].n17 XThR.Tn[7].n16 0.00771154
R23223 XThR.Tn[7].n12 XThR.Tn[7].n11 0.00771154
R23224 XThR.Tn[0].n2 XThR.Tn[0].n1 332.332
R23225 XThR.Tn[0].n2 XThR.Tn[0].n0 296.493
R23226 XThR.Tn[0] XThR.Tn[0].n82 161.363
R23227 XThR.Tn[0] XThR.Tn[0].n77 161.363
R23228 XThR.Tn[0] XThR.Tn[0].n72 161.363
R23229 XThR.Tn[0] XThR.Tn[0].n67 161.363
R23230 XThR.Tn[0] XThR.Tn[0].n62 161.363
R23231 XThR.Tn[0] XThR.Tn[0].n57 161.363
R23232 XThR.Tn[0] XThR.Tn[0].n52 161.363
R23233 XThR.Tn[0] XThR.Tn[0].n47 161.363
R23234 XThR.Tn[0] XThR.Tn[0].n42 161.363
R23235 XThR.Tn[0] XThR.Tn[0].n37 161.363
R23236 XThR.Tn[0] XThR.Tn[0].n32 161.363
R23237 XThR.Tn[0] XThR.Tn[0].n27 161.363
R23238 XThR.Tn[0] XThR.Tn[0].n22 161.363
R23239 XThR.Tn[0] XThR.Tn[0].n17 161.363
R23240 XThR.Tn[0] XThR.Tn[0].n12 161.363
R23241 XThR.Tn[0] XThR.Tn[0].n10 161.363
R23242 XThR.Tn[0].n84 XThR.Tn[0].n83 161.3
R23243 XThR.Tn[0].n79 XThR.Tn[0].n78 161.3
R23244 XThR.Tn[0].n74 XThR.Tn[0].n73 161.3
R23245 XThR.Tn[0].n69 XThR.Tn[0].n68 161.3
R23246 XThR.Tn[0].n64 XThR.Tn[0].n63 161.3
R23247 XThR.Tn[0].n59 XThR.Tn[0].n58 161.3
R23248 XThR.Tn[0].n54 XThR.Tn[0].n53 161.3
R23249 XThR.Tn[0].n49 XThR.Tn[0].n48 161.3
R23250 XThR.Tn[0].n44 XThR.Tn[0].n43 161.3
R23251 XThR.Tn[0].n39 XThR.Tn[0].n38 161.3
R23252 XThR.Tn[0].n34 XThR.Tn[0].n33 161.3
R23253 XThR.Tn[0].n29 XThR.Tn[0].n28 161.3
R23254 XThR.Tn[0].n24 XThR.Tn[0].n23 161.3
R23255 XThR.Tn[0].n19 XThR.Tn[0].n18 161.3
R23256 XThR.Tn[0].n14 XThR.Tn[0].n13 161.3
R23257 XThR.Tn[0].n82 XThR.Tn[0].t32 161.106
R23258 XThR.Tn[0].n77 XThR.Tn[0].t36 161.106
R23259 XThR.Tn[0].n72 XThR.Tn[0].t16 161.106
R23260 XThR.Tn[0].n67 XThR.Tn[0].t65 161.106
R23261 XThR.Tn[0].n62 XThR.Tn[0].t31 161.106
R23262 XThR.Tn[0].n57 XThR.Tn[0].t53 161.106
R23263 XThR.Tn[0].n52 XThR.Tn[0].t34 161.106
R23264 XThR.Tn[0].n47 XThR.Tn[0].t14 161.106
R23265 XThR.Tn[0].n42 XThR.Tn[0].t63 161.106
R23266 XThR.Tn[0].n37 XThR.Tn[0].t68 161.106
R23267 XThR.Tn[0].n32 XThR.Tn[0].t52 161.106
R23268 XThR.Tn[0].n27 XThR.Tn[0].t15 161.106
R23269 XThR.Tn[0].n22 XThR.Tn[0].t51 161.106
R23270 XThR.Tn[0].n17 XThR.Tn[0].t33 161.106
R23271 XThR.Tn[0].n12 XThR.Tn[0].t58 161.106
R23272 XThR.Tn[0].n10 XThR.Tn[0].t40 161.106
R23273 XThR.Tn[0].n83 XThR.Tn[0].t20 159.978
R23274 XThR.Tn[0].n78 XThR.Tn[0].t30 159.978
R23275 XThR.Tn[0].n73 XThR.Tn[0].t73 159.978
R23276 XThR.Tn[0].n68 XThR.Tn[0].t57 159.978
R23277 XThR.Tn[0].n63 XThR.Tn[0].t19 159.978
R23278 XThR.Tn[0].n58 XThR.Tn[0].t49 159.978
R23279 XThR.Tn[0].n53 XThR.Tn[0].t29 159.978
R23280 XThR.Tn[0].n48 XThR.Tn[0].t71 159.978
R23281 XThR.Tn[0].n43 XThR.Tn[0].t55 159.978
R23282 XThR.Tn[0].n38 XThR.Tn[0].t64 159.978
R23283 XThR.Tn[0].n33 XThR.Tn[0].t46 159.978
R23284 XThR.Tn[0].n28 XThR.Tn[0].t72 159.978
R23285 XThR.Tn[0].n23 XThR.Tn[0].t44 159.978
R23286 XThR.Tn[0].n18 XThR.Tn[0].t26 159.978
R23287 XThR.Tn[0].n13 XThR.Tn[0].t50 159.978
R23288 XThR.Tn[0].n82 XThR.Tn[0].t18 145.038
R23289 XThR.Tn[0].n77 XThR.Tn[0].t42 145.038
R23290 XThR.Tn[0].n72 XThR.Tn[0].t22 145.038
R23291 XThR.Tn[0].n67 XThR.Tn[0].t69 145.038
R23292 XThR.Tn[0].n62 XThR.Tn[0].t37 145.038
R23293 XThR.Tn[0].n57 XThR.Tn[0].t17 145.038
R23294 XThR.Tn[0].n52 XThR.Tn[0].t25 145.038
R23295 XThR.Tn[0].n47 XThR.Tn[0].t70 145.038
R23296 XThR.Tn[0].n42 XThR.Tn[0].t66 145.038
R23297 XThR.Tn[0].n37 XThR.Tn[0].t35 145.038
R23298 XThR.Tn[0].n32 XThR.Tn[0].t60 145.038
R23299 XThR.Tn[0].n27 XThR.Tn[0].t21 145.038
R23300 XThR.Tn[0].n22 XThR.Tn[0].t59 145.038
R23301 XThR.Tn[0].n17 XThR.Tn[0].t41 145.038
R23302 XThR.Tn[0].n12 XThR.Tn[0].t67 145.038
R23303 XThR.Tn[0].n10 XThR.Tn[0].t48 145.038
R23304 XThR.Tn[0].n83 XThR.Tn[0].t39 143.911
R23305 XThR.Tn[0].n78 XThR.Tn[0].t62 143.911
R23306 XThR.Tn[0].n73 XThR.Tn[0].t45 143.911
R23307 XThR.Tn[0].n68 XThR.Tn[0].t27 143.911
R23308 XThR.Tn[0].n63 XThR.Tn[0].t56 143.911
R23309 XThR.Tn[0].n58 XThR.Tn[0].t38 143.911
R23310 XThR.Tn[0].n53 XThR.Tn[0].t47 143.911
R23311 XThR.Tn[0].n48 XThR.Tn[0].t28 143.911
R23312 XThR.Tn[0].n43 XThR.Tn[0].t23 143.911
R23313 XThR.Tn[0].n38 XThR.Tn[0].t54 143.911
R23314 XThR.Tn[0].n33 XThR.Tn[0].t13 143.911
R23315 XThR.Tn[0].n28 XThR.Tn[0].t43 143.911
R23316 XThR.Tn[0].n23 XThR.Tn[0].t12 143.911
R23317 XThR.Tn[0].n18 XThR.Tn[0].t61 143.911
R23318 XThR.Tn[0].n13 XThR.Tn[0].t24 143.911
R23319 XThR.Tn[0].n7 XThR.Tn[0].n5 135.249
R23320 XThR.Tn[0].n9 XThR.Tn[0].n3 98.982
R23321 XThR.Tn[0].n8 XThR.Tn[0].n4 98.982
R23322 XThR.Tn[0].n7 XThR.Tn[0].n6 98.982
R23323 XThR.Tn[0].n9 XThR.Tn[0].n8 36.2672
R23324 XThR.Tn[0].n8 XThR.Tn[0].n7 36.2672
R23325 XThR.Tn[0].n88 XThR.Tn[0].n9 32.6405
R23326 XThR.Tn[0].n1 XThR.Tn[0].t3 26.5955
R23327 XThR.Tn[0].n1 XThR.Tn[0].t2 26.5955
R23328 XThR.Tn[0].n0 XThR.Tn[0].t4 26.5955
R23329 XThR.Tn[0].n0 XThR.Tn[0].t5 26.5955
R23330 XThR.Tn[0].n3 XThR.Tn[0].t7 24.9236
R23331 XThR.Tn[0].n3 XThR.Tn[0].t8 24.9236
R23332 XThR.Tn[0].n4 XThR.Tn[0].t6 24.9236
R23333 XThR.Tn[0].n4 XThR.Tn[0].t9 24.9236
R23334 XThR.Tn[0].n5 XThR.Tn[0].t11 24.9236
R23335 XThR.Tn[0].n5 XThR.Tn[0].t10 24.9236
R23336 XThR.Tn[0].n6 XThR.Tn[0].t1 24.9236
R23337 XThR.Tn[0].n6 XThR.Tn[0].t0 24.9236
R23338 XThR.Tn[0] XThR.Tn[0].n2 23.3605
R23339 XThR.Tn[0] XThR.Tn[0].n88 6.7205
R23340 XThR.Tn[0].n88 XThR.Tn[0] 6.36522
R23341 XThR.Tn[0] XThR.Tn[0].n11 5.34038
R23342 XThR.Tn[0].n16 XThR.Tn[0].n15 4.5005
R23343 XThR.Tn[0].n21 XThR.Tn[0].n20 4.5005
R23344 XThR.Tn[0].n26 XThR.Tn[0].n25 4.5005
R23345 XThR.Tn[0].n31 XThR.Tn[0].n30 4.5005
R23346 XThR.Tn[0].n36 XThR.Tn[0].n35 4.5005
R23347 XThR.Tn[0].n41 XThR.Tn[0].n40 4.5005
R23348 XThR.Tn[0].n46 XThR.Tn[0].n45 4.5005
R23349 XThR.Tn[0].n51 XThR.Tn[0].n50 4.5005
R23350 XThR.Tn[0].n56 XThR.Tn[0].n55 4.5005
R23351 XThR.Tn[0].n61 XThR.Tn[0].n60 4.5005
R23352 XThR.Tn[0].n66 XThR.Tn[0].n65 4.5005
R23353 XThR.Tn[0].n71 XThR.Tn[0].n70 4.5005
R23354 XThR.Tn[0].n76 XThR.Tn[0].n75 4.5005
R23355 XThR.Tn[0].n81 XThR.Tn[0].n80 4.5005
R23356 XThR.Tn[0].n86 XThR.Tn[0].n85 4.5005
R23357 XThR.Tn[0].n87 XThR.Tn[0] 3.70586
R23358 XThR.Tn[0].n16 XThR.Tn[0] 2.52282
R23359 XThR.Tn[0].n21 XThR.Tn[0] 2.52282
R23360 XThR.Tn[0].n26 XThR.Tn[0] 2.52282
R23361 XThR.Tn[0].n31 XThR.Tn[0] 2.52282
R23362 XThR.Tn[0].n36 XThR.Tn[0] 2.52282
R23363 XThR.Tn[0].n41 XThR.Tn[0] 2.52282
R23364 XThR.Tn[0].n46 XThR.Tn[0] 2.52282
R23365 XThR.Tn[0].n51 XThR.Tn[0] 2.52282
R23366 XThR.Tn[0].n56 XThR.Tn[0] 2.52282
R23367 XThR.Tn[0].n61 XThR.Tn[0] 2.52282
R23368 XThR.Tn[0].n66 XThR.Tn[0] 2.52282
R23369 XThR.Tn[0].n71 XThR.Tn[0] 2.52282
R23370 XThR.Tn[0].n76 XThR.Tn[0] 2.52282
R23371 XThR.Tn[0].n81 XThR.Tn[0] 2.52282
R23372 XThR.Tn[0].n86 XThR.Tn[0] 2.52282
R23373 XThR.Tn[0].n84 XThR.Tn[0] 1.08677
R23374 XThR.Tn[0].n79 XThR.Tn[0] 1.08677
R23375 XThR.Tn[0].n74 XThR.Tn[0] 1.08677
R23376 XThR.Tn[0].n69 XThR.Tn[0] 1.08677
R23377 XThR.Tn[0].n64 XThR.Tn[0] 1.08677
R23378 XThR.Tn[0].n59 XThR.Tn[0] 1.08677
R23379 XThR.Tn[0].n54 XThR.Tn[0] 1.08677
R23380 XThR.Tn[0].n49 XThR.Tn[0] 1.08677
R23381 XThR.Tn[0].n44 XThR.Tn[0] 1.08677
R23382 XThR.Tn[0].n39 XThR.Tn[0] 1.08677
R23383 XThR.Tn[0].n34 XThR.Tn[0] 1.08677
R23384 XThR.Tn[0].n29 XThR.Tn[0] 1.08677
R23385 XThR.Tn[0].n24 XThR.Tn[0] 1.08677
R23386 XThR.Tn[0].n19 XThR.Tn[0] 1.08677
R23387 XThR.Tn[0].n14 XThR.Tn[0] 1.08677
R23388 XThR.Tn[0] XThR.Tn[0].n16 0.839786
R23389 XThR.Tn[0] XThR.Tn[0].n21 0.839786
R23390 XThR.Tn[0] XThR.Tn[0].n26 0.839786
R23391 XThR.Tn[0] XThR.Tn[0].n31 0.839786
R23392 XThR.Tn[0] XThR.Tn[0].n36 0.839786
R23393 XThR.Tn[0] XThR.Tn[0].n41 0.839786
R23394 XThR.Tn[0] XThR.Tn[0].n46 0.839786
R23395 XThR.Tn[0] XThR.Tn[0].n51 0.839786
R23396 XThR.Tn[0] XThR.Tn[0].n56 0.839786
R23397 XThR.Tn[0] XThR.Tn[0].n61 0.839786
R23398 XThR.Tn[0] XThR.Tn[0].n66 0.839786
R23399 XThR.Tn[0] XThR.Tn[0].n71 0.839786
R23400 XThR.Tn[0] XThR.Tn[0].n76 0.839786
R23401 XThR.Tn[0] XThR.Tn[0].n81 0.839786
R23402 XThR.Tn[0] XThR.Tn[0].n86 0.839786
R23403 XThR.Tn[0].n11 XThR.Tn[0] 0.499542
R23404 XThR.Tn[0].n85 XThR.Tn[0] 0.063
R23405 XThR.Tn[0].n80 XThR.Tn[0] 0.063
R23406 XThR.Tn[0].n75 XThR.Tn[0] 0.063
R23407 XThR.Tn[0].n70 XThR.Tn[0] 0.063
R23408 XThR.Tn[0].n65 XThR.Tn[0] 0.063
R23409 XThR.Tn[0].n60 XThR.Tn[0] 0.063
R23410 XThR.Tn[0].n55 XThR.Tn[0] 0.063
R23411 XThR.Tn[0].n50 XThR.Tn[0] 0.063
R23412 XThR.Tn[0].n45 XThR.Tn[0] 0.063
R23413 XThR.Tn[0].n40 XThR.Tn[0] 0.063
R23414 XThR.Tn[0].n35 XThR.Tn[0] 0.063
R23415 XThR.Tn[0].n30 XThR.Tn[0] 0.063
R23416 XThR.Tn[0].n25 XThR.Tn[0] 0.063
R23417 XThR.Tn[0].n20 XThR.Tn[0] 0.063
R23418 XThR.Tn[0].n15 XThR.Tn[0] 0.063
R23419 XThR.Tn[0].n87 XThR.Tn[0] 0.0540714
R23420 XThR.Tn[0] XThR.Tn[0].n87 0.038
R23421 XThR.Tn[0].n11 XThR.Tn[0] 0.0143889
R23422 XThR.Tn[0].n85 XThR.Tn[0].n84 0.00771154
R23423 XThR.Tn[0].n80 XThR.Tn[0].n79 0.00771154
R23424 XThR.Tn[0].n75 XThR.Tn[0].n74 0.00771154
R23425 XThR.Tn[0].n70 XThR.Tn[0].n69 0.00771154
R23426 XThR.Tn[0].n65 XThR.Tn[0].n64 0.00771154
R23427 XThR.Tn[0].n60 XThR.Tn[0].n59 0.00771154
R23428 XThR.Tn[0].n55 XThR.Tn[0].n54 0.00771154
R23429 XThR.Tn[0].n50 XThR.Tn[0].n49 0.00771154
R23430 XThR.Tn[0].n45 XThR.Tn[0].n44 0.00771154
R23431 XThR.Tn[0].n40 XThR.Tn[0].n39 0.00771154
R23432 XThR.Tn[0].n35 XThR.Tn[0].n34 0.00771154
R23433 XThR.Tn[0].n30 XThR.Tn[0].n29 0.00771154
R23434 XThR.Tn[0].n25 XThR.Tn[0].n24 0.00771154
R23435 XThR.Tn[0].n20 XThR.Tn[0].n19 0.00771154
R23436 XThR.Tn[0].n15 XThR.Tn[0].n14 0.00771154
R23437 XThR.Tn[8].n87 XThR.Tn[8].n86 256.103
R23438 XThR.Tn[8].n2 XThR.Tn[8].n0 243.68
R23439 XThR.Tn[8].n5 XThR.Tn[8].n3 241.847
R23440 XThR.Tn[8].n2 XThR.Tn[8].n1 205.28
R23441 XThR.Tn[8].n87 XThR.Tn[8].n85 202.095
R23442 XThR.Tn[8].n5 XThR.Tn[8].n4 185
R23443 XThR.Tn[8] XThR.Tn[8].n78 161.363
R23444 XThR.Tn[8] XThR.Tn[8].n73 161.363
R23445 XThR.Tn[8] XThR.Tn[8].n68 161.363
R23446 XThR.Tn[8] XThR.Tn[8].n63 161.363
R23447 XThR.Tn[8] XThR.Tn[8].n58 161.363
R23448 XThR.Tn[8] XThR.Tn[8].n53 161.363
R23449 XThR.Tn[8] XThR.Tn[8].n48 161.363
R23450 XThR.Tn[8] XThR.Tn[8].n43 161.363
R23451 XThR.Tn[8] XThR.Tn[8].n38 161.363
R23452 XThR.Tn[8] XThR.Tn[8].n33 161.363
R23453 XThR.Tn[8] XThR.Tn[8].n28 161.363
R23454 XThR.Tn[8] XThR.Tn[8].n23 161.363
R23455 XThR.Tn[8] XThR.Tn[8].n18 161.363
R23456 XThR.Tn[8] XThR.Tn[8].n13 161.363
R23457 XThR.Tn[8] XThR.Tn[8].n8 161.363
R23458 XThR.Tn[8] XThR.Tn[8].n6 161.363
R23459 XThR.Tn[8].n80 XThR.Tn[8].n79 161.3
R23460 XThR.Tn[8].n75 XThR.Tn[8].n74 161.3
R23461 XThR.Tn[8].n70 XThR.Tn[8].n69 161.3
R23462 XThR.Tn[8].n65 XThR.Tn[8].n64 161.3
R23463 XThR.Tn[8].n60 XThR.Tn[8].n59 161.3
R23464 XThR.Tn[8].n55 XThR.Tn[8].n54 161.3
R23465 XThR.Tn[8].n50 XThR.Tn[8].n49 161.3
R23466 XThR.Tn[8].n45 XThR.Tn[8].n44 161.3
R23467 XThR.Tn[8].n40 XThR.Tn[8].n39 161.3
R23468 XThR.Tn[8].n35 XThR.Tn[8].n34 161.3
R23469 XThR.Tn[8].n30 XThR.Tn[8].n29 161.3
R23470 XThR.Tn[8].n25 XThR.Tn[8].n24 161.3
R23471 XThR.Tn[8].n20 XThR.Tn[8].n19 161.3
R23472 XThR.Tn[8].n15 XThR.Tn[8].n14 161.3
R23473 XThR.Tn[8].n10 XThR.Tn[8].n9 161.3
R23474 XThR.Tn[8].n78 XThR.Tn[8].t23 161.106
R23475 XThR.Tn[8].n73 XThR.Tn[8].t29 161.106
R23476 XThR.Tn[8].n68 XThR.Tn[8].t71 161.106
R23477 XThR.Tn[8].n63 XThR.Tn[8].t57 161.106
R23478 XThR.Tn[8].n58 XThR.Tn[8].t21 161.106
R23479 XThR.Tn[8].n53 XThR.Tn[8].t46 161.106
R23480 XThR.Tn[8].n48 XThR.Tn[8].t27 161.106
R23481 XThR.Tn[8].n43 XThR.Tn[8].t69 161.106
R23482 XThR.Tn[8].n38 XThR.Tn[8].t56 161.106
R23483 XThR.Tn[8].n33 XThR.Tn[8].t61 161.106
R23484 XThR.Tn[8].n28 XThR.Tn[8].t44 161.106
R23485 XThR.Tn[8].n23 XThR.Tn[8].t70 161.106
R23486 XThR.Tn[8].n18 XThR.Tn[8].t43 161.106
R23487 XThR.Tn[8].n13 XThR.Tn[8].t26 161.106
R23488 XThR.Tn[8].n8 XThR.Tn[8].t49 161.106
R23489 XThR.Tn[8].n6 XThR.Tn[8].t33 161.106
R23490 XThR.Tn[8].n79 XThR.Tn[8].t19 159.978
R23491 XThR.Tn[8].n74 XThR.Tn[8].t25 159.978
R23492 XThR.Tn[8].n69 XThR.Tn[8].t67 159.978
R23493 XThR.Tn[8].n64 XThR.Tn[8].t54 159.978
R23494 XThR.Tn[8].n59 XThR.Tn[8].t16 159.978
R23495 XThR.Tn[8].n54 XThR.Tn[8].t42 159.978
R23496 XThR.Tn[8].n49 XThR.Tn[8].t24 159.978
R23497 XThR.Tn[8].n44 XThR.Tn[8].t64 159.978
R23498 XThR.Tn[8].n39 XThR.Tn[8].t51 159.978
R23499 XThR.Tn[8].n34 XThR.Tn[8].t58 159.978
R23500 XThR.Tn[8].n29 XThR.Tn[8].t41 159.978
R23501 XThR.Tn[8].n24 XThR.Tn[8].t66 159.978
R23502 XThR.Tn[8].n19 XThR.Tn[8].t40 159.978
R23503 XThR.Tn[8].n14 XThR.Tn[8].t22 159.978
R23504 XThR.Tn[8].n9 XThR.Tn[8].t45 159.978
R23505 XThR.Tn[8].n78 XThR.Tn[8].t73 145.038
R23506 XThR.Tn[8].n73 XThR.Tn[8].t35 145.038
R23507 XThR.Tn[8].n68 XThR.Tn[8].t15 145.038
R23508 XThR.Tn[8].n63 XThR.Tn[8].t62 145.038
R23509 XThR.Tn[8].n58 XThR.Tn[8].t30 145.038
R23510 XThR.Tn[8].n53 XThR.Tn[8].t72 145.038
R23511 XThR.Tn[8].n48 XThR.Tn[8].t17 145.038
R23512 XThR.Tn[8].n43 XThR.Tn[8].t63 145.038
R23513 XThR.Tn[8].n38 XThR.Tn[8].t60 145.038
R23514 XThR.Tn[8].n33 XThR.Tn[8].t28 145.038
R23515 XThR.Tn[8].n28 XThR.Tn[8].t52 145.038
R23516 XThR.Tn[8].n23 XThR.Tn[8].t12 145.038
R23517 XThR.Tn[8].n18 XThR.Tn[8].t50 145.038
R23518 XThR.Tn[8].n13 XThR.Tn[8].t34 145.038
R23519 XThR.Tn[8].n8 XThR.Tn[8].t59 145.038
R23520 XThR.Tn[8].n6 XThR.Tn[8].t39 145.038
R23521 XThR.Tn[8].n79 XThR.Tn[8].t32 143.911
R23522 XThR.Tn[8].n74 XThR.Tn[8].t55 143.911
R23523 XThR.Tn[8].n69 XThR.Tn[8].t37 143.911
R23524 XThR.Tn[8].n64 XThR.Tn[8].t18 143.911
R23525 XThR.Tn[8].n59 XThR.Tn[8].t48 143.911
R23526 XThR.Tn[8].n54 XThR.Tn[8].t31 143.911
R23527 XThR.Tn[8].n49 XThR.Tn[8].t38 143.911
R23528 XThR.Tn[8].n44 XThR.Tn[8].t20 143.911
R23529 XThR.Tn[8].n39 XThR.Tn[8].t14 143.911
R23530 XThR.Tn[8].n34 XThR.Tn[8].t47 143.911
R23531 XThR.Tn[8].n29 XThR.Tn[8].t68 143.911
R23532 XThR.Tn[8].n24 XThR.Tn[8].t36 143.911
R23533 XThR.Tn[8].n19 XThR.Tn[8].t65 143.911
R23534 XThR.Tn[8].n14 XThR.Tn[8].t53 143.911
R23535 XThR.Tn[8].n9 XThR.Tn[8].t13 143.911
R23536 XThR.Tn[8] XThR.Tn[8].n2 35.7652
R23537 XThR.Tn[8].n85 XThR.Tn[8].t9 26.5955
R23538 XThR.Tn[8].n85 XThR.Tn[8].t11 26.5955
R23539 XThR.Tn[8].n0 XThR.Tn[8].t7 26.5955
R23540 XThR.Tn[8].n0 XThR.Tn[8].t5 26.5955
R23541 XThR.Tn[8].n1 XThR.Tn[8].t8 26.5955
R23542 XThR.Tn[8].n1 XThR.Tn[8].t6 26.5955
R23543 XThR.Tn[8].n86 XThR.Tn[8].t0 26.5955
R23544 XThR.Tn[8].n86 XThR.Tn[8].t10 26.5955
R23545 XThR.Tn[8].n4 XThR.Tn[8].t2 24.9236
R23546 XThR.Tn[8].n4 XThR.Tn[8].t4 24.9236
R23547 XThR.Tn[8].n3 XThR.Tn[8].t1 24.9236
R23548 XThR.Tn[8].n3 XThR.Tn[8].t3 24.9236
R23549 XThR.Tn[8] XThR.Tn[8].n5 18.8943
R23550 XThR.Tn[8].n88 XThR.Tn[8].n87 13.5534
R23551 XThR.Tn[8].n84 XThR.Tn[8] 7.82692
R23552 XThR.Tn[8].n84 XThR.Tn[8] 6.34069
R23553 XThR.Tn[8] XThR.Tn[8].n7 5.34038
R23554 XThR.Tn[8].n12 XThR.Tn[8].n11 4.5005
R23555 XThR.Tn[8].n17 XThR.Tn[8].n16 4.5005
R23556 XThR.Tn[8].n22 XThR.Tn[8].n21 4.5005
R23557 XThR.Tn[8].n27 XThR.Tn[8].n26 4.5005
R23558 XThR.Tn[8].n32 XThR.Tn[8].n31 4.5005
R23559 XThR.Tn[8].n37 XThR.Tn[8].n36 4.5005
R23560 XThR.Tn[8].n42 XThR.Tn[8].n41 4.5005
R23561 XThR.Tn[8].n47 XThR.Tn[8].n46 4.5005
R23562 XThR.Tn[8].n52 XThR.Tn[8].n51 4.5005
R23563 XThR.Tn[8].n57 XThR.Tn[8].n56 4.5005
R23564 XThR.Tn[8].n62 XThR.Tn[8].n61 4.5005
R23565 XThR.Tn[8].n67 XThR.Tn[8].n66 4.5005
R23566 XThR.Tn[8].n72 XThR.Tn[8].n71 4.5005
R23567 XThR.Tn[8].n77 XThR.Tn[8].n76 4.5005
R23568 XThR.Tn[8].n82 XThR.Tn[8].n81 4.5005
R23569 XThR.Tn[8].n83 XThR.Tn[8] 3.70586
R23570 XThR.Tn[8].n12 XThR.Tn[8] 2.52282
R23571 XThR.Tn[8].n17 XThR.Tn[8] 2.52282
R23572 XThR.Tn[8].n22 XThR.Tn[8] 2.52282
R23573 XThR.Tn[8].n27 XThR.Tn[8] 2.52282
R23574 XThR.Tn[8].n32 XThR.Tn[8] 2.52282
R23575 XThR.Tn[8].n37 XThR.Tn[8] 2.52282
R23576 XThR.Tn[8].n42 XThR.Tn[8] 2.52282
R23577 XThR.Tn[8].n47 XThR.Tn[8] 2.52282
R23578 XThR.Tn[8].n52 XThR.Tn[8] 2.52282
R23579 XThR.Tn[8].n57 XThR.Tn[8] 2.52282
R23580 XThR.Tn[8].n62 XThR.Tn[8] 2.52282
R23581 XThR.Tn[8].n67 XThR.Tn[8] 2.52282
R23582 XThR.Tn[8].n72 XThR.Tn[8] 2.52282
R23583 XThR.Tn[8].n77 XThR.Tn[8] 2.52282
R23584 XThR.Tn[8].n82 XThR.Tn[8] 2.52282
R23585 XThR.Tn[8] XThR.Tn[8].n84 1.79489
R23586 XThR.Tn[8] XThR.Tn[8].n88 1.50638
R23587 XThR.Tn[8].n88 XThR.Tn[8] 1.19676
R23588 XThR.Tn[8].n80 XThR.Tn[8] 1.08677
R23589 XThR.Tn[8].n75 XThR.Tn[8] 1.08677
R23590 XThR.Tn[8].n70 XThR.Tn[8] 1.08677
R23591 XThR.Tn[8].n65 XThR.Tn[8] 1.08677
R23592 XThR.Tn[8].n60 XThR.Tn[8] 1.08677
R23593 XThR.Tn[8].n55 XThR.Tn[8] 1.08677
R23594 XThR.Tn[8].n50 XThR.Tn[8] 1.08677
R23595 XThR.Tn[8].n45 XThR.Tn[8] 1.08677
R23596 XThR.Tn[8].n40 XThR.Tn[8] 1.08677
R23597 XThR.Tn[8].n35 XThR.Tn[8] 1.08677
R23598 XThR.Tn[8].n30 XThR.Tn[8] 1.08677
R23599 XThR.Tn[8].n25 XThR.Tn[8] 1.08677
R23600 XThR.Tn[8].n20 XThR.Tn[8] 1.08677
R23601 XThR.Tn[8].n15 XThR.Tn[8] 1.08677
R23602 XThR.Tn[8].n10 XThR.Tn[8] 1.08677
R23603 XThR.Tn[8] XThR.Tn[8].n12 0.839786
R23604 XThR.Tn[8] XThR.Tn[8].n17 0.839786
R23605 XThR.Tn[8] XThR.Tn[8].n22 0.839786
R23606 XThR.Tn[8] XThR.Tn[8].n27 0.839786
R23607 XThR.Tn[8] XThR.Tn[8].n32 0.839786
R23608 XThR.Tn[8] XThR.Tn[8].n37 0.839786
R23609 XThR.Tn[8] XThR.Tn[8].n42 0.839786
R23610 XThR.Tn[8] XThR.Tn[8].n47 0.839786
R23611 XThR.Tn[8] XThR.Tn[8].n52 0.839786
R23612 XThR.Tn[8] XThR.Tn[8].n57 0.839786
R23613 XThR.Tn[8] XThR.Tn[8].n62 0.839786
R23614 XThR.Tn[8] XThR.Tn[8].n67 0.839786
R23615 XThR.Tn[8] XThR.Tn[8].n72 0.839786
R23616 XThR.Tn[8] XThR.Tn[8].n77 0.839786
R23617 XThR.Tn[8] XThR.Tn[8].n82 0.839786
R23618 XThR.Tn[8].n7 XThR.Tn[8] 0.499542
R23619 XThR.Tn[8].n81 XThR.Tn[8] 0.063
R23620 XThR.Tn[8].n76 XThR.Tn[8] 0.063
R23621 XThR.Tn[8].n71 XThR.Tn[8] 0.063
R23622 XThR.Tn[8].n66 XThR.Tn[8] 0.063
R23623 XThR.Tn[8].n61 XThR.Tn[8] 0.063
R23624 XThR.Tn[8].n56 XThR.Tn[8] 0.063
R23625 XThR.Tn[8].n51 XThR.Tn[8] 0.063
R23626 XThR.Tn[8].n46 XThR.Tn[8] 0.063
R23627 XThR.Tn[8].n41 XThR.Tn[8] 0.063
R23628 XThR.Tn[8].n36 XThR.Tn[8] 0.063
R23629 XThR.Tn[8].n31 XThR.Tn[8] 0.063
R23630 XThR.Tn[8].n26 XThR.Tn[8] 0.063
R23631 XThR.Tn[8].n21 XThR.Tn[8] 0.063
R23632 XThR.Tn[8].n16 XThR.Tn[8] 0.063
R23633 XThR.Tn[8].n11 XThR.Tn[8] 0.063
R23634 XThR.Tn[8].n83 XThR.Tn[8] 0.0540714
R23635 XThR.Tn[8] XThR.Tn[8].n83 0.038
R23636 XThR.Tn[8].n7 XThR.Tn[8] 0.0143889
R23637 XThR.Tn[8].n81 XThR.Tn[8].n80 0.00771154
R23638 XThR.Tn[8].n76 XThR.Tn[8].n75 0.00771154
R23639 XThR.Tn[8].n71 XThR.Tn[8].n70 0.00771154
R23640 XThR.Tn[8].n66 XThR.Tn[8].n65 0.00771154
R23641 XThR.Tn[8].n61 XThR.Tn[8].n60 0.00771154
R23642 XThR.Tn[8].n56 XThR.Tn[8].n55 0.00771154
R23643 XThR.Tn[8].n51 XThR.Tn[8].n50 0.00771154
R23644 XThR.Tn[8].n46 XThR.Tn[8].n45 0.00771154
R23645 XThR.Tn[8].n41 XThR.Tn[8].n40 0.00771154
R23646 XThR.Tn[8].n36 XThR.Tn[8].n35 0.00771154
R23647 XThR.Tn[8].n31 XThR.Tn[8].n30 0.00771154
R23648 XThR.Tn[8].n26 XThR.Tn[8].n25 0.00771154
R23649 XThR.Tn[8].n21 XThR.Tn[8].n20 0.00771154
R23650 XThR.Tn[8].n16 XThR.Tn[8].n15 0.00771154
R23651 XThR.Tn[8].n11 XThR.Tn[8].n10 0.00771154
R23652 XThC.XTB3.Y.n6 XThC.XTB3.Y.t3 212.081
R23653 XThC.XTB3.Y.n5 XThC.XTB3.Y.t15 212.081
R23654 XThC.XTB3.Y.n11 XThC.XTB3.Y.t14 212.081
R23655 XThC.XTB3.Y.n3 XThC.XTB3.Y.t10 212.081
R23656 XThC.XTB3.Y.n15 XThC.XTB3.Y.t11 212.081
R23657 XThC.XTB3.Y.n16 XThC.XTB3.Y.t12 212.081
R23658 XThC.XTB3.Y.n18 XThC.XTB3.Y.t4 212.081
R23659 XThC.XTB3.Y.n14 XThC.XTB3.Y.t16 212.081
R23660 XThC.XTB3.Y.n22 XThC.XTB3.Y.n2 201.288
R23661 XThC.XTB3.Y.n8 XThC.XTB3.Y.n7 173.761
R23662 XThC.XTB3.Y.n17 XThC.XTB3.Y 158.656
R23663 XThC.XTB3.Y.n10 XThC.XTB3.Y.n9 152
R23664 XThC.XTB3.Y.n8 XThC.XTB3.Y.n4 152
R23665 XThC.XTB3.Y.n13 XThC.XTB3.Y.n12 152
R23666 XThC.XTB3.Y.n20 XThC.XTB3.Y.n19 152
R23667 XThC.XTB3.Y.n6 XThC.XTB3.Y.t9 139.78
R23668 XThC.XTB3.Y.n5 XThC.XTB3.Y.t6 139.78
R23669 XThC.XTB3.Y.n11 XThC.XTB3.Y.t5 139.78
R23670 XThC.XTB3.Y.n3 XThC.XTB3.Y.t17 139.78
R23671 XThC.XTB3.Y.n15 XThC.XTB3.Y.t8 139.78
R23672 XThC.XTB3.Y.n16 XThC.XTB3.Y.t18 139.78
R23673 XThC.XTB3.Y.n18 XThC.XTB3.Y.t13 139.78
R23674 XThC.XTB3.Y.n14 XThC.XTB3.Y.t7 139.78
R23675 XThC.XTB3.Y.n0 XThC.XTB3.Y.t1 132.067
R23676 XThC.XTB3.Y.n21 XThC.XTB3.Y.n13 61.4096
R23677 XThC.XTB3.Y.n16 XThC.XTB3.Y.n15 61.346
R23678 XThC.XTB3.Y.n21 XThC.XTB3.Y 54.2785
R23679 XThC.XTB3.Y.n10 XThC.XTB3.Y.n4 49.6611
R23680 XThC.XTB3.Y.n12 XThC.XTB3.Y.n11 45.2793
R23681 XThC.XTB3.Y.n7 XThC.XTB3.Y.n5 42.3581
R23682 XThC.XTB3.Y.n19 XThC.XTB3.Y.n14 30.6732
R23683 XThC.XTB3.Y.n19 XThC.XTB3.Y.n18 30.6732
R23684 XThC.XTB3.Y.n18 XThC.XTB3.Y.n17 30.6732
R23685 XThC.XTB3.Y.n17 XThC.XTB3.Y.n16 30.6732
R23686 XThC.XTB3.Y.n2 XThC.XTB3.Y.t0 26.5955
R23687 XThC.XTB3.Y.n2 XThC.XTB3.Y.t2 26.5955
R23688 XThC.XTB3.Y XThC.XTB3.Y.n22 23.489
R23689 XThC.XTB3.Y.n9 XThC.XTB3.Y.n8 21.7605
R23690 XThC.XTB3.Y.n7 XThC.XTB3.Y.n6 18.9884
R23691 XThC.XTB3.Y.n12 XThC.XTB3.Y.n3 16.0672
R23692 XThC.XTB3.Y.n20 XThC.XTB3.Y 14.8485
R23693 XThC.XTB3.Y.n13 XThC.XTB3.Y 11.5205
R23694 XThC.XTB3.Y.n22 XThC.XTB3.Y.n21 10.8207
R23695 XThC.XTB3.Y.n9 XThC.XTB3.Y 10.2405
R23696 XThC.XTB3.Y XThC.XTB3.Y.n20 8.7045
R23697 XThC.XTB3.Y.n5 XThC.XTB3.Y.n4 7.30353
R23698 XThC.XTB3.Y.n11 XThC.XTB3.Y.n10 4.38232
R23699 XThC.XTB3.Y.n1 XThC.XTB3.Y.n0 4.15748
R23700 XThC.XTB3.Y XThC.XTB3.Y.n1 3.76521
R23701 XThC.XTB3.Y.n0 XThC.XTB3.Y 1.17559
R23702 XThC.XTB3.Y.n1 XThC.XTB3.Y 0.921363
R23703 data[4].n3 data[4].t0 231.835
R23704 data[4].n0 data[4].t3 230.155
R23705 data[4].n0 data[4].t1 157.856
R23706 data[4].n3 data[4].t2 157.07
R23707 data[4].n1 data[4].n0 152
R23708 data[4].n4 data[4].n3 152
R23709 data[4].n2 data[4].n1 25.6681
R23710 data[4].n4 data[4].n2 10.7642
R23711 data[4].n2 data[4] 2.763
R23712 data[4].n1 data[4] 2.10199
R23713 data[4] data[4].n4 2.01193
R23714 XThR.Tn[13].n87 XThR.Tn[13].n86 256.103
R23715 XThR.Tn[13].n2 XThR.Tn[13].n0 243.68
R23716 XThR.Tn[13].n5 XThR.Tn[13].n3 241.847
R23717 XThR.Tn[13].n2 XThR.Tn[13].n1 205.28
R23718 XThR.Tn[13].n87 XThR.Tn[13].n85 202.094
R23719 XThR.Tn[13].n5 XThR.Tn[13].n4 185
R23720 XThR.Tn[13] XThR.Tn[13].n78 161.363
R23721 XThR.Tn[13] XThR.Tn[13].n73 161.363
R23722 XThR.Tn[13] XThR.Tn[13].n68 161.363
R23723 XThR.Tn[13] XThR.Tn[13].n63 161.363
R23724 XThR.Tn[13] XThR.Tn[13].n58 161.363
R23725 XThR.Tn[13] XThR.Tn[13].n53 161.363
R23726 XThR.Tn[13] XThR.Tn[13].n48 161.363
R23727 XThR.Tn[13] XThR.Tn[13].n43 161.363
R23728 XThR.Tn[13] XThR.Tn[13].n38 161.363
R23729 XThR.Tn[13] XThR.Tn[13].n33 161.363
R23730 XThR.Tn[13] XThR.Tn[13].n28 161.363
R23731 XThR.Tn[13] XThR.Tn[13].n23 161.363
R23732 XThR.Tn[13] XThR.Tn[13].n18 161.363
R23733 XThR.Tn[13] XThR.Tn[13].n13 161.363
R23734 XThR.Tn[13] XThR.Tn[13].n8 161.363
R23735 XThR.Tn[13] XThR.Tn[13].n6 161.363
R23736 XThR.Tn[13].n80 XThR.Tn[13].n79 161.3
R23737 XThR.Tn[13].n75 XThR.Tn[13].n74 161.3
R23738 XThR.Tn[13].n70 XThR.Tn[13].n69 161.3
R23739 XThR.Tn[13].n65 XThR.Tn[13].n64 161.3
R23740 XThR.Tn[13].n60 XThR.Tn[13].n59 161.3
R23741 XThR.Tn[13].n55 XThR.Tn[13].n54 161.3
R23742 XThR.Tn[13].n50 XThR.Tn[13].n49 161.3
R23743 XThR.Tn[13].n45 XThR.Tn[13].n44 161.3
R23744 XThR.Tn[13].n40 XThR.Tn[13].n39 161.3
R23745 XThR.Tn[13].n35 XThR.Tn[13].n34 161.3
R23746 XThR.Tn[13].n30 XThR.Tn[13].n29 161.3
R23747 XThR.Tn[13].n25 XThR.Tn[13].n24 161.3
R23748 XThR.Tn[13].n20 XThR.Tn[13].n19 161.3
R23749 XThR.Tn[13].n15 XThR.Tn[13].n14 161.3
R23750 XThR.Tn[13].n10 XThR.Tn[13].n9 161.3
R23751 XThR.Tn[13].n78 XThR.Tn[13].t56 161.106
R23752 XThR.Tn[13].n73 XThR.Tn[13].t62 161.106
R23753 XThR.Tn[13].n68 XThR.Tn[13].t40 161.106
R23754 XThR.Tn[13].n63 XThR.Tn[13].t27 161.106
R23755 XThR.Tn[13].n58 XThR.Tn[13].t55 161.106
R23756 XThR.Tn[13].n53 XThR.Tn[13].t17 161.106
R23757 XThR.Tn[13].n48 XThR.Tn[13].t59 161.106
R23758 XThR.Tn[13].n43 XThR.Tn[13].t38 161.106
R23759 XThR.Tn[13].n38 XThR.Tn[13].t25 161.106
R23760 XThR.Tn[13].n33 XThR.Tn[13].t30 161.106
R23761 XThR.Tn[13].n28 XThR.Tn[13].t16 161.106
R23762 XThR.Tn[13].n23 XThR.Tn[13].t39 161.106
R23763 XThR.Tn[13].n18 XThR.Tn[13].t14 161.106
R23764 XThR.Tn[13].n13 XThR.Tn[13].t57 161.106
R23765 XThR.Tn[13].n8 XThR.Tn[13].t21 161.106
R23766 XThR.Tn[13].n6 XThR.Tn[13].t64 161.106
R23767 XThR.Tn[13].n79 XThR.Tn[13].t47 159.978
R23768 XThR.Tn[13].n74 XThR.Tn[13].t54 159.978
R23769 XThR.Tn[13].n69 XThR.Tn[13].t36 159.978
R23770 XThR.Tn[13].n64 XThR.Tn[13].t20 159.978
R23771 XThR.Tn[13].n59 XThR.Tn[13].t45 159.978
R23772 XThR.Tn[13].n54 XThR.Tn[13].t73 159.978
R23773 XThR.Tn[13].n49 XThR.Tn[13].t53 159.978
R23774 XThR.Tn[13].n44 XThR.Tn[13].t33 159.978
R23775 XThR.Tn[13].n39 XThR.Tn[13].t18 159.978
R23776 XThR.Tn[13].n34 XThR.Tn[13].t26 159.978
R23777 XThR.Tn[13].n29 XThR.Tn[13].t71 159.978
R23778 XThR.Tn[13].n24 XThR.Tn[13].t35 159.978
R23779 XThR.Tn[13].n19 XThR.Tn[13].t70 159.978
R23780 XThR.Tn[13].n14 XThR.Tn[13].t52 159.978
R23781 XThR.Tn[13].n9 XThR.Tn[13].t12 159.978
R23782 XThR.Tn[13].n78 XThR.Tn[13].t42 145.038
R23783 XThR.Tn[13].n73 XThR.Tn[13].t69 145.038
R23784 XThR.Tn[13].n68 XThR.Tn[13].t50 145.038
R23785 XThR.Tn[13].n63 XThR.Tn[13].t31 145.038
R23786 XThR.Tn[13].n58 XThR.Tn[13].t63 145.038
R23787 XThR.Tn[13].n53 XThR.Tn[13].t41 145.038
R23788 XThR.Tn[13].n48 XThR.Tn[13].t51 145.038
R23789 XThR.Tn[13].n43 XThR.Tn[13].t32 145.038
R23790 XThR.Tn[13].n38 XThR.Tn[13].t29 145.038
R23791 XThR.Tn[13].n33 XThR.Tn[13].t60 145.038
R23792 XThR.Tn[13].n28 XThR.Tn[13].t24 145.038
R23793 XThR.Tn[13].n23 XThR.Tn[13].t49 145.038
R23794 XThR.Tn[13].n18 XThR.Tn[13].t22 145.038
R23795 XThR.Tn[13].n13 XThR.Tn[13].t65 145.038
R23796 XThR.Tn[13].n8 XThR.Tn[13].t28 145.038
R23797 XThR.Tn[13].n6 XThR.Tn[13].t72 145.038
R23798 XThR.Tn[13].n79 XThR.Tn[13].t61 143.911
R23799 XThR.Tn[13].n74 XThR.Tn[13].t23 143.911
R23800 XThR.Tn[13].n69 XThR.Tn[13].t67 143.911
R23801 XThR.Tn[13].n64 XThR.Tn[13].t46 143.911
R23802 XThR.Tn[13].n59 XThR.Tn[13].t15 143.911
R23803 XThR.Tn[13].n54 XThR.Tn[13].t58 143.911
R23804 XThR.Tn[13].n49 XThR.Tn[13].t68 143.911
R23805 XThR.Tn[13].n44 XThR.Tn[13].t48 143.911
R23806 XThR.Tn[13].n39 XThR.Tn[13].t43 143.911
R23807 XThR.Tn[13].n34 XThR.Tn[13].t13 143.911
R23808 XThR.Tn[13].n29 XThR.Tn[13].t37 143.911
R23809 XThR.Tn[13].n24 XThR.Tn[13].t66 143.911
R23810 XThR.Tn[13].n19 XThR.Tn[13].t34 143.911
R23811 XThR.Tn[13].n14 XThR.Tn[13].t19 143.911
R23812 XThR.Tn[13].n9 XThR.Tn[13].t44 143.911
R23813 XThR.Tn[13] XThR.Tn[13].n2 35.7652
R23814 XThR.Tn[13].n85 XThR.Tn[13].t2 26.5955
R23815 XThR.Tn[13].n85 XThR.Tn[13].t0 26.5955
R23816 XThR.Tn[13].n0 XThR.Tn[13].t9 26.5955
R23817 XThR.Tn[13].n0 XThR.Tn[13].t11 26.5955
R23818 XThR.Tn[13].n1 XThR.Tn[13].t10 26.5955
R23819 XThR.Tn[13].n1 XThR.Tn[13].t8 26.5955
R23820 XThR.Tn[13].n86 XThR.Tn[13].t3 26.5955
R23821 XThR.Tn[13].n86 XThR.Tn[13].t1 26.5955
R23822 XThR.Tn[13].n4 XThR.Tn[13].t6 24.9236
R23823 XThR.Tn[13].n4 XThR.Tn[13].t4 24.9236
R23824 XThR.Tn[13].n3 XThR.Tn[13].t7 24.9236
R23825 XThR.Tn[13].n3 XThR.Tn[13].t5 24.9236
R23826 XThR.Tn[13] XThR.Tn[13].n5 22.9615
R23827 XThR.Tn[13].n88 XThR.Tn[13].n87 13.5534
R23828 XThR.Tn[13].n84 XThR.Tn[13] 8.8494
R23829 XThR.Tn[13] XThR.Tn[13].n7 5.34038
R23830 XThR.Tn[13].n12 XThR.Tn[13].n11 4.5005
R23831 XThR.Tn[13].n17 XThR.Tn[13].n16 4.5005
R23832 XThR.Tn[13].n22 XThR.Tn[13].n21 4.5005
R23833 XThR.Tn[13].n27 XThR.Tn[13].n26 4.5005
R23834 XThR.Tn[13].n32 XThR.Tn[13].n31 4.5005
R23835 XThR.Tn[13].n37 XThR.Tn[13].n36 4.5005
R23836 XThR.Tn[13].n42 XThR.Tn[13].n41 4.5005
R23837 XThR.Tn[13].n47 XThR.Tn[13].n46 4.5005
R23838 XThR.Tn[13].n52 XThR.Tn[13].n51 4.5005
R23839 XThR.Tn[13].n57 XThR.Tn[13].n56 4.5005
R23840 XThR.Tn[13].n62 XThR.Tn[13].n61 4.5005
R23841 XThR.Tn[13].n67 XThR.Tn[13].n66 4.5005
R23842 XThR.Tn[13].n72 XThR.Tn[13].n71 4.5005
R23843 XThR.Tn[13].n77 XThR.Tn[13].n76 4.5005
R23844 XThR.Tn[13].n82 XThR.Tn[13].n81 4.5005
R23845 XThR.Tn[13].n83 XThR.Tn[13] 3.70586
R23846 XThR.Tn[13].n88 XThR.Tn[13].n84 2.99115
R23847 XThR.Tn[13].n88 XThR.Tn[13] 2.87153
R23848 XThR.Tn[13].n12 XThR.Tn[13] 2.52282
R23849 XThR.Tn[13].n17 XThR.Tn[13] 2.52282
R23850 XThR.Tn[13].n22 XThR.Tn[13] 2.52282
R23851 XThR.Tn[13].n27 XThR.Tn[13] 2.52282
R23852 XThR.Tn[13].n32 XThR.Tn[13] 2.52282
R23853 XThR.Tn[13].n37 XThR.Tn[13] 2.52282
R23854 XThR.Tn[13].n42 XThR.Tn[13] 2.52282
R23855 XThR.Tn[13].n47 XThR.Tn[13] 2.52282
R23856 XThR.Tn[13].n52 XThR.Tn[13] 2.52282
R23857 XThR.Tn[13].n57 XThR.Tn[13] 2.52282
R23858 XThR.Tn[13].n62 XThR.Tn[13] 2.52282
R23859 XThR.Tn[13].n67 XThR.Tn[13] 2.52282
R23860 XThR.Tn[13].n72 XThR.Tn[13] 2.52282
R23861 XThR.Tn[13].n77 XThR.Tn[13] 2.52282
R23862 XThR.Tn[13].n82 XThR.Tn[13] 2.52282
R23863 XThR.Tn[13].n84 XThR.Tn[13] 2.2734
R23864 XThR.Tn[13] XThR.Tn[13].n88 1.50638
R23865 XThR.Tn[13].n80 XThR.Tn[13] 1.08677
R23866 XThR.Tn[13].n75 XThR.Tn[13] 1.08677
R23867 XThR.Tn[13].n70 XThR.Tn[13] 1.08677
R23868 XThR.Tn[13].n65 XThR.Tn[13] 1.08677
R23869 XThR.Tn[13].n60 XThR.Tn[13] 1.08677
R23870 XThR.Tn[13].n55 XThR.Tn[13] 1.08677
R23871 XThR.Tn[13].n50 XThR.Tn[13] 1.08677
R23872 XThR.Tn[13].n45 XThR.Tn[13] 1.08677
R23873 XThR.Tn[13].n40 XThR.Tn[13] 1.08677
R23874 XThR.Tn[13].n35 XThR.Tn[13] 1.08677
R23875 XThR.Tn[13].n30 XThR.Tn[13] 1.08677
R23876 XThR.Tn[13].n25 XThR.Tn[13] 1.08677
R23877 XThR.Tn[13].n20 XThR.Tn[13] 1.08677
R23878 XThR.Tn[13].n15 XThR.Tn[13] 1.08677
R23879 XThR.Tn[13].n10 XThR.Tn[13] 1.08677
R23880 XThR.Tn[13] XThR.Tn[13].n12 0.839786
R23881 XThR.Tn[13] XThR.Tn[13].n17 0.839786
R23882 XThR.Tn[13] XThR.Tn[13].n22 0.839786
R23883 XThR.Tn[13] XThR.Tn[13].n27 0.839786
R23884 XThR.Tn[13] XThR.Tn[13].n32 0.839786
R23885 XThR.Tn[13] XThR.Tn[13].n37 0.839786
R23886 XThR.Tn[13] XThR.Tn[13].n42 0.839786
R23887 XThR.Tn[13] XThR.Tn[13].n47 0.839786
R23888 XThR.Tn[13] XThR.Tn[13].n52 0.839786
R23889 XThR.Tn[13] XThR.Tn[13].n57 0.839786
R23890 XThR.Tn[13] XThR.Tn[13].n62 0.839786
R23891 XThR.Tn[13] XThR.Tn[13].n67 0.839786
R23892 XThR.Tn[13] XThR.Tn[13].n72 0.839786
R23893 XThR.Tn[13] XThR.Tn[13].n77 0.839786
R23894 XThR.Tn[13] XThR.Tn[13].n82 0.839786
R23895 XThR.Tn[13].n7 XThR.Tn[13] 0.499542
R23896 XThR.Tn[13].n81 XThR.Tn[13] 0.063
R23897 XThR.Tn[13].n76 XThR.Tn[13] 0.063
R23898 XThR.Tn[13].n71 XThR.Tn[13] 0.063
R23899 XThR.Tn[13].n66 XThR.Tn[13] 0.063
R23900 XThR.Tn[13].n61 XThR.Tn[13] 0.063
R23901 XThR.Tn[13].n56 XThR.Tn[13] 0.063
R23902 XThR.Tn[13].n51 XThR.Tn[13] 0.063
R23903 XThR.Tn[13].n46 XThR.Tn[13] 0.063
R23904 XThR.Tn[13].n41 XThR.Tn[13] 0.063
R23905 XThR.Tn[13].n36 XThR.Tn[13] 0.063
R23906 XThR.Tn[13].n31 XThR.Tn[13] 0.063
R23907 XThR.Tn[13].n26 XThR.Tn[13] 0.063
R23908 XThR.Tn[13].n21 XThR.Tn[13] 0.063
R23909 XThR.Tn[13].n16 XThR.Tn[13] 0.063
R23910 XThR.Tn[13].n11 XThR.Tn[13] 0.063
R23911 XThR.Tn[13].n83 XThR.Tn[13] 0.0540714
R23912 XThR.Tn[13] XThR.Tn[13].n83 0.038
R23913 XThR.Tn[13].n7 XThR.Tn[13] 0.0143889
R23914 XThR.Tn[13].n81 XThR.Tn[13].n80 0.00771154
R23915 XThR.Tn[13].n76 XThR.Tn[13].n75 0.00771154
R23916 XThR.Tn[13].n71 XThR.Tn[13].n70 0.00771154
R23917 XThR.Tn[13].n66 XThR.Tn[13].n65 0.00771154
R23918 XThR.Tn[13].n61 XThR.Tn[13].n60 0.00771154
R23919 XThR.Tn[13].n56 XThR.Tn[13].n55 0.00771154
R23920 XThR.Tn[13].n51 XThR.Tn[13].n50 0.00771154
R23921 XThR.Tn[13].n46 XThR.Tn[13].n45 0.00771154
R23922 XThR.Tn[13].n41 XThR.Tn[13].n40 0.00771154
R23923 XThR.Tn[13].n36 XThR.Tn[13].n35 0.00771154
R23924 XThR.Tn[13].n31 XThR.Tn[13].n30 0.00771154
R23925 XThR.Tn[13].n26 XThR.Tn[13].n25 0.00771154
R23926 XThR.Tn[13].n21 XThR.Tn[13].n20 0.00771154
R23927 XThR.Tn[13].n16 XThR.Tn[13].n15 0.00771154
R23928 XThR.Tn[13].n11 XThR.Tn[13].n10 0.00771154
R23929 data[0].n1 data[0].t0 230.155
R23930 data[0].n0 data[0].t2 228.463
R23931 data[0].n1 data[0].t1 157.856
R23932 data[0].n0 data[0].t3 157.07
R23933 data[0].n2 data[0].n1 152.768
R23934 data[0].n4 data[0].n0 152.256
R23935 data[0].n3 data[0].n2 24.1398
R23936 data[0].n4 data[0].n3 9.48418
R23937 data[0] data[0].n4 6.1445
R23938 data[0].n2 data[0] 5.6325
R23939 data[0].n3 data[0] 2.638
R23940 XThR.XTB4.Y XThR.XTB4.Y.t0 230.518
R23941 XThR.XTB4.Y.n10 XThR.XTB4.Y.t12 212.081
R23942 XThR.XTB4.Y.n11 XThR.XTB4.Y.t2 212.081
R23943 XThR.XTB4.Y.n16 XThR.XTB4.Y.t7 212.081
R23944 XThR.XTB4.Y.n17 XThR.XTB4.Y.t6 212.081
R23945 XThR.XTB4.Y.n0 XThR.XTB4.Y.t17 212.081
R23946 XThR.XTB4.Y.n1 XThR.XTB4.Y.t5 212.081
R23947 XThR.XTB4.Y.n3 XThR.XTB4.Y.t15 212.081
R23948 XThR.XTB4.Y.n4 XThR.XTB4.Y.t4 212.081
R23949 XThR.XTB4.Y.n13 XThR.XTB4.Y.n12 173.761
R23950 XThR.XTB4.Y.n2 XThR.XTB4.Y 167.361
R23951 XThR.XTB4.Y.n19 XThR.XTB4.Y.n18 152
R23952 XThR.XTB4.Y.n15 XThR.XTB4.Y.n14 152
R23953 XThR.XTB4.Y.n13 XThR.XTB4.Y.n9 152
R23954 XThR.XTB4.Y.n6 XThR.XTB4.Y.n5 152
R23955 XThR.XTB4.Y.n10 XThR.XTB4.Y.t3 139.78
R23956 XThR.XTB4.Y.n11 XThR.XTB4.Y.t9 139.78
R23957 XThR.XTB4.Y.n16 XThR.XTB4.Y.t14 139.78
R23958 XThR.XTB4.Y.n17 XThR.XTB4.Y.t11 139.78
R23959 XThR.XTB4.Y.n0 XThR.XTB4.Y.t10 139.78
R23960 XThR.XTB4.Y.n1 XThR.XTB4.Y.t16 139.78
R23961 XThR.XTB4.Y.n3 XThR.XTB4.Y.t8 139.78
R23962 XThR.XTB4.Y.n4 XThR.XTB4.Y.t13 139.78
R23963 XThR.XTB4.Y.n21 XThR.XTB4.Y.t1 133.386
R23964 XThR.XTB4.Y.n20 XThR.XTB4.Y.n19 72.9296
R23965 XThR.XTB4.Y.n1 XThR.XTB4.Y.n0 61.346
R23966 XThR.XTB4.Y.n15 XThR.XTB4.Y.n9 49.6611
R23967 XThR.XTB4.Y.n18 XThR.XTB4.Y.n16 45.2793
R23968 XThR.XTB4.Y.n12 XThR.XTB4.Y.n11 42.3581
R23969 XThR.XTB4.Y.n20 XThR.XTB4.Y.n8 38.1854
R23970 XThR.XTB4.Y.n2 XThR.XTB4.Y.n1 30.6732
R23971 XThR.XTB4.Y.n3 XThR.XTB4.Y.n2 30.6732
R23972 XThR.XTB4.Y.n5 XThR.XTB4.Y.n3 30.6732
R23973 XThR.XTB4.Y.n5 XThR.XTB4.Y.n4 30.6732
R23974 XThR.XTB4.Y XThR.XTB4.Y.n21 28.966
R23975 XThR.XTB4.Y.n14 XThR.XTB4.Y.n13 21.7605
R23976 XThR.XTB4.Y.n14 XThR.XTB4.Y 21.1205
R23977 XThR.XTB4.Y.n12 XThR.XTB4.Y.n10 18.9884
R23978 XThR.XTB4.Y.n18 XThR.XTB4.Y.n17 16.0672
R23979 XThR.XTB4.Y.n21 XThR.XTB4.Y.n20 11.994
R23980 XThR.XTB4.Y.n22 XThR.XTB4.Y 11.6875
R23981 XThR.XTB4.Y.n8 XThR.XTB4.Y.n7 8.21182
R23982 XThR.XTB4.Y.n11 XThR.XTB4.Y.n9 7.30353
R23983 XThR.XTB4.Y.n8 XThR.XTB4.Y.n6 7.24578
R23984 XThR.XTB4.Y.n22 XThR.XTB4.Y 7.23528
R23985 XThR.XTB4.Y.n6 XThR.XTB4.Y 6.08654
R23986 XThR.XTB4.Y XThR.XTB4.Y.n22 5.04292
R23987 XThR.XTB4.Y.n16 XThR.XTB4.Y.n15 4.38232
R23988 XThR.XTB4.Y.n7 XThR.XTB4.Y 1.79489
R23989 XThR.XTB4.Y.n7 XThR.XTB4.Y 0.966538
R23990 XThR.XTB4.Y.n19 XThR.XTB4.Y 0.6405
R23991 XThR.XTB1.Y.n9 XThR.XTB1.Y.t12 212.081
R23992 XThR.XTB1.Y.n10 XThR.XTB1.Y.t17 212.081
R23993 XThR.XTB1.Y.n15 XThR.XTB1.Y.t6 212.081
R23994 XThR.XTB1.Y.n16 XThR.XTB1.Y.t3 212.081
R23995 XThR.XTB1.Y.n1 XThR.XTB1.Y.t10 212.081
R23996 XThR.XTB1.Y.n2 XThR.XTB1.Y.t14 212.081
R23997 XThR.XTB1.Y.n4 XThR.XTB1.Y.t8 212.081
R23998 XThR.XTB1.Y.n5 XThR.XTB1.Y.t13 212.081
R23999 XThR.XTB1.Y.n21 XThR.XTB1.Y.n20 201.288
R24000 XThR.XTB1.Y.n12 XThR.XTB1.Y.n11 173.761
R24001 XThR.XTB1.Y.n3 XThR.XTB1.Y 167.361
R24002 XThR.XTB1.Y.n18 XThR.XTB1.Y.n17 152
R24003 XThR.XTB1.Y.n14 XThR.XTB1.Y.n13 152
R24004 XThR.XTB1.Y.n12 XThR.XTB1.Y.n8 152
R24005 XThR.XTB1.Y.n7 XThR.XTB1.Y.n6 152
R24006 XThR.XTB1.Y.n9 XThR.XTB1.Y.t16 139.78
R24007 XThR.XTB1.Y.n10 XThR.XTB1.Y.t5 139.78
R24008 XThR.XTB1.Y.n15 XThR.XTB1.Y.t11 139.78
R24009 XThR.XTB1.Y.n16 XThR.XTB1.Y.t9 139.78
R24010 XThR.XTB1.Y.n1 XThR.XTB1.Y.t18 139.78
R24011 XThR.XTB1.Y.n2 XThR.XTB1.Y.t7 139.78
R24012 XThR.XTB1.Y.n4 XThR.XTB1.Y.t15 139.78
R24013 XThR.XTB1.Y.n5 XThR.XTB1.Y.t4 139.78
R24014 XThR.XTB1.Y.n0 XThR.XTB1.Y.t1 130.548
R24015 XThR.XTB1.Y.n19 XThR.XTB1.Y 74.7655
R24016 XThR.XTB1.Y.n19 XThR.XTB1.Y.n18 61.4072
R24017 XThR.XTB1.Y.n2 XThR.XTB1.Y.n1 61.346
R24018 XThR.XTB1.Y.n14 XThR.XTB1.Y.n8 49.6611
R24019 XThR.XTB1.Y.n17 XThR.XTB1.Y.n15 45.2793
R24020 XThR.XTB1.Y.n11 XThR.XTB1.Y.n10 42.3581
R24021 XThR.XTB1.Y XThR.XTB1.Y.n21 36.289
R24022 XThR.XTB1.Y.n3 XThR.XTB1.Y.n2 30.6732
R24023 XThR.XTB1.Y.n4 XThR.XTB1.Y.n3 30.6732
R24024 XThR.XTB1.Y.n6 XThR.XTB1.Y.n4 30.6732
R24025 XThR.XTB1.Y.n6 XThR.XTB1.Y.n5 30.6732
R24026 XThR.XTB1.Y.n20 XThR.XTB1.Y.t2 26.5955
R24027 XThR.XTB1.Y.n20 XThR.XTB1.Y.t0 26.5955
R24028 XThR.XTB1.Y.n13 XThR.XTB1.Y.n12 21.7605
R24029 XThR.XTB1.Y.n13 XThR.XTB1.Y 21.1205
R24030 XThR.XTB1.Y.n11 XThR.XTB1.Y.n9 18.9884
R24031 XThR.XTB1.Y XThR.XTB1.Y.n7 17.4085
R24032 XThR.XTB1.Y.n22 XThR.XTB1.Y 16.5652
R24033 XThR.XTB1.Y.n17 XThR.XTB1.Y.n16 16.0672
R24034 XThR.XTB1.Y.n21 XThR.XTB1.Y.n19 10.8571
R24035 XThR.XTB1.Y XThR.XTB1.Y.n22 9.03579
R24036 XThR.XTB1.Y.n10 XThR.XTB1.Y.n8 7.30353
R24037 XThR.XTB1.Y.n7 XThR.XTB1.Y 6.1445
R24038 XThR.XTB1.Y.n15 XThR.XTB1.Y.n14 4.38232
R24039 XThR.XTB1.Y XThR.XTB1.Y.n0 3.46739
R24040 XThR.XTB1.Y.n0 XThR.XTB1.Y 2.74112
R24041 XThR.XTB1.Y.n22 XThR.XTB1.Y 2.21057
R24042 XThR.XTB1.Y.n18 XThR.XTB1.Y 0.6405
R24043 XThR.XTB3.Y.n9 XThR.XTB3.Y.t7 212.081
R24044 XThR.XTB3.Y.n10 XThR.XTB3.Y.t11 212.081
R24045 XThR.XTB3.Y.n15 XThR.XTB3.Y.t18 212.081
R24046 XThR.XTB3.Y.n16 XThR.XTB3.Y.t14 212.081
R24047 XThR.XTB3.Y.n1 XThR.XTB3.Y.t9 212.081
R24048 XThR.XTB3.Y.n2 XThR.XTB3.Y.t13 212.081
R24049 XThR.XTB3.Y.n4 XThR.XTB3.Y.t8 212.081
R24050 XThR.XTB3.Y.n5 XThR.XTB3.Y.t12 212.081
R24051 XThR.XTB3.Y.n21 XThR.XTB3.Y.n20 201.288
R24052 XThR.XTB3.Y.n12 XThR.XTB3.Y.n11 173.761
R24053 XThR.XTB3.Y.n3 XThR.XTB3.Y 167.361
R24054 XThR.XTB3.Y.n18 XThR.XTB3.Y.n17 152
R24055 XThR.XTB3.Y.n14 XThR.XTB3.Y.n13 152
R24056 XThR.XTB3.Y.n12 XThR.XTB3.Y.n8 152
R24057 XThR.XTB3.Y.n7 XThR.XTB3.Y.n6 152
R24058 XThR.XTB3.Y.n9 XThR.XTB3.Y.t10 139.78
R24059 XThR.XTB3.Y.n10 XThR.XTB3.Y.t16 139.78
R24060 XThR.XTB3.Y.n15 XThR.XTB3.Y.t5 139.78
R24061 XThR.XTB3.Y.n16 XThR.XTB3.Y.t3 139.78
R24062 XThR.XTB3.Y.n1 XThR.XTB3.Y.t17 139.78
R24063 XThR.XTB3.Y.n2 XThR.XTB3.Y.t6 139.78
R24064 XThR.XTB3.Y.n4 XThR.XTB3.Y.t15 139.78
R24065 XThR.XTB3.Y.n5 XThR.XTB3.Y.t4 139.78
R24066 XThR.XTB3.Y.n0 XThR.XTB3.Y.t1 130.548
R24067 XThR.XTB3.Y.n19 XThR.XTB3.Y.n18 61.4096
R24068 XThR.XTB3.Y.n2 XThR.XTB3.Y.n1 61.346
R24069 XThR.XTB3.Y.n14 XThR.XTB3.Y.n8 49.6611
R24070 XThR.XTB3.Y.n19 XThR.XTB3.Y 45.5863
R24071 XThR.XTB3.Y.n17 XThR.XTB3.Y.n15 45.2793
R24072 XThR.XTB3.Y.n11 XThR.XTB3.Y.n10 42.3581
R24073 XThR.XTB3.Y XThR.XTB3.Y.n21 36.289
R24074 XThR.XTB3.Y.n3 XThR.XTB3.Y.n2 30.6732
R24075 XThR.XTB3.Y.n4 XThR.XTB3.Y.n3 30.6732
R24076 XThR.XTB3.Y.n6 XThR.XTB3.Y.n4 30.6732
R24077 XThR.XTB3.Y.n6 XThR.XTB3.Y.n5 30.6732
R24078 XThR.XTB3.Y.n20 XThR.XTB3.Y.t2 26.5955
R24079 XThR.XTB3.Y.n20 XThR.XTB3.Y.t0 26.5955
R24080 XThR.XTB3.Y.n13 XThR.XTB3.Y.n12 21.7605
R24081 XThR.XTB3.Y.n13 XThR.XTB3.Y 21.1205
R24082 XThR.XTB3.Y.n11 XThR.XTB3.Y.n9 18.9884
R24083 XThR.XTB3.Y XThR.XTB3.Y.n7 17.4085
R24084 XThR.XTB3.Y.n22 XThR.XTB3.Y 16.5652
R24085 XThR.XTB3.Y.n17 XThR.XTB3.Y.n16 16.0672
R24086 XThR.XTB3.Y.n21 XThR.XTB3.Y.n19 10.8207
R24087 XThR.XTB3.Y XThR.XTB3.Y.n22 9.03579
R24088 XThR.XTB3.Y.n10 XThR.XTB3.Y.n8 7.30353
R24089 XThR.XTB3.Y.n7 XThR.XTB3.Y 6.1445
R24090 XThR.XTB3.Y.n15 XThR.XTB3.Y.n14 4.38232
R24091 XThR.XTB3.Y XThR.XTB3.Y.n0 3.46739
R24092 XThR.XTB3.Y.n0 XThR.XTB3.Y 2.74112
R24093 XThR.XTB3.Y.n22 XThR.XTB3.Y 2.21057
R24094 XThR.XTB3.Y.n18 XThR.XTB3.Y 0.6405
R24095 data[6].n0 data[6].t0 230.576
R24096 data[6].n0 data[6].t1 158.275
R24097 data[6].n1 data[6].n0 152
R24098 data[6].n1 data[6] 11.9995
R24099 data[6] data[6].n1 6.66717
R24100 data[1].n4 data[1].t2 230.576
R24101 data[1].n1 data[1].t0 230.363
R24102 data[1].n0 data[1].t4 229.369
R24103 data[1].n4 data[1].t5 158.275
R24104 data[1].n1 data[1].t3 158.064
R24105 data[1].n0 data[1].t1 157.07
R24106 data[1].n2 data[1].n1 153.28
R24107 data[1].n7 data[1].n0 153.147
R24108 data[1].n5 data[1].n4 152
R24109 data[1].n7 data[1].n6 16.3874
R24110 data[1].n6 data[1].n5 14.9641
R24111 data[1].n3 data[1].n2 9.3005
R24112 data[1].n6 data[1].n3 6.49639
R24113 data[1] data[1].n7 3.24826
R24114 data[1].n2 data[1] 2.92621
R24115 data[1].n3 data[1] 2.15819
R24116 data[1].n5 data[1] 2.13383
R24117 data[2].n0 data[2].t0 230.576
R24118 data[2].n0 data[2].t1 158.275
R24119 data[2].n1 data[2].n0 152
R24120 data[2].n1 data[2] 12.7714
R24121 data[2] data[2].n1 2.13383
R24122 data[5].n4 data[5].t2 230.576
R24123 data[5].n1 data[5].t0 230.363
R24124 data[5].n0 data[5].t1 229.369
R24125 data[5].n4 data[5].t5 158.275
R24126 data[5].n1 data[5].t3 158.064
R24127 data[5].n0 data[5].t4 157.07
R24128 data[5].n2 data[5].n1 152.256
R24129 data[5].n7 data[5].n0 152.238
R24130 data[5].n5 data[5].n4 152
R24131 data[5].n7 data[5].n6 16.3874
R24132 data[5].n6 data[5].n5 14.6005
R24133 data[5].n3 data[5].n2 9.3005
R24134 data[5].n5 data[5] 6.66717
R24135 data[5].n6 data[5].n3 6.49639
R24136 data[5].n2 data[5] 6.1445
R24137 data[5] data[5].n7 5.68939
R24138 data[5].n3 data[5] 2.28319
R24139 bias[0] bias[0].t0 12.1467
R24140 bias[2].n0 bias[2].t0 56.8043
R24141 bias[2].n0 bias[2] 6.35112
R24142 bias[2] bias[2].n0 0.828709
R24143 data[3].n0 data[3].t1 230.576
R24144 data[3].n0 data[3].t0 158.275
R24145 data[3].n1 data[3].n0 153.553
R24146 data[3].n1 data[3] 11.6078
R24147 data[3] data[3].n1 2.90959
R24148 data[7].n0 data[7].t0 230.576
R24149 data[7].n0 data[7].t1 158.275
R24150 data[7].n1 data[7].n0 152
R24151 data[7].n1 data[7] 11.9995
R24152 data[7] data[7].n1 6.66717
R24153 bias[1] bias[1].t0 23.8076
C0 XThR.Tn[14] XA.XIR[14].XIC[12].icell.Ien 0.15202f
C1 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.Ien 0.04854f
C2 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PDM 0.02765f
C3 XA.XIR[6].XIC[11].icell.Ien Iout 0.06821f
C4 XA.XIR[14].XIC_15.icell.PUM VPWR 0.01655f
C5 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR 0.08209f
C6 XA.XIR[7].XIC[5].icell.PUM VPWR 0.01015f
C7 XThC.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.03184f
C8 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.PDM 0.02104f
C9 XA.XIR[14].XIC[9].icell.Ien VPWR 0.19845f
C10 Vbias bias[0] 0.21039f
C11 bias[1] bias[2] 0.16429f
C12 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.Ien 0.04854f
C13 a_4861_9615# XThC.Tn[3] 0.27012f
C14 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.Ien 0.04854f
C15 XA.XIR[14].XIC[5].icell.Ien Iout 0.06821f
C16 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR 0.38903f
C17 XThR.Tn[3] XA.XIR[3].XIC[2].icell.Ien 0.15202f
C18 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR 0.35722f
C19 XA.XIR[13].XIC[7].icell.Ien Iout 0.06821f
C20 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0222f
C21 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.PDM 0.02104f
C22 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.Ien 0.04854f
C23 XA.XIR[6].XIC_dummy_right.icell.Iout VPWR 0.11567f
C24 XA.XIR[15].XIC[1].icell.Ien Vbias 0.15966f
C25 XA.XIR[11].XIC[11].icell.PUM VPWR 0.01015f
C26 XA.XIR[14].XIC_dummy_right.icell.Iout XA.XIR[15].XIC_dummy_right.icell.Iout 0.04047f
C27 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PDM 0.04035f
C28 XA.XIR[11].XIC[2].icell.PDM Vbias 0.03922f
C29 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PDM 0.02765f
C30 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PDM 0.04035f
C31 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.PDM 0.02104f
C32 XA.XIR[10].XIC[6].icell.PDM Vbias 0.03922f
C33 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.02765f
C34 XThC.Tn[2] XThR.Tn[14] 0.29362f
C35 XThC.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.03605f
C36 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.02765f
C37 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PDM 0.04035f
C38 XThR.Tn[4] VPWR 8.2593f
C39 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.PDM 0.02104f
C40 XThC.Tn[10] XA.XIR[2].XIC[10].icell.Ien 0.03605f
C41 XA.XIR[15].XIC[6].icell.Ien Vbias 0.15966f
C42 XA.XIR[2].XIC[14].icell.Ien Iout 0.06821f
C43 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.Ien 0.04854f
C44 a_n1049_7493# VPWR 0.72084f
C45 XThR.Tn[8] XA.XIR[8].XIC_15.icell.Ien 0.13564f
C46 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.Ien 0.04854f
C47 XA.XIR[11].XIC[12].icell.Ien VPWR 0.1979f
C48 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.PDM 0.02104f
C49 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.Ien 0.04854f
C50 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PDM 0.02765f
C51 XA.XIR[4].XIC[9].icell.Ien Vbias 0.19161f
C52 XA.XIR[14].XIC[0].icell.Ien Iout 0.06814f
C53 XA.XIR[0].XIC[0].icell.Ien Vbias 0.19207f
C54 XThR.Tn[14] XA.XIR[14].XIC[10].icell.Ien 0.15202f
C55 XThR.XTB6.Y VPWR 1.05512f
C56 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.PDM 0.02104f
C57 XThR.Tn[13] Iout 1.19576f
C58 XA.XIR[14].XIC[13].icell.PUM VPWR 0.01015f
C59 XA.XIR[8].XIC[3].icell.Ien Vbias 0.19161f
C60 XThC.Tn[13] VPWR 7.4336f
C61 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.PDM 0.02104f
C62 XThR.Tn[5] XA.XIR[5].XIC[14].icell.Ien 0.15202f
C63 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.Ien 0.04854f
C64 XA.XIR[15].XIC[8].icell.PUM VPWR 0.01015f
C65 XA.XIR[0].XIC[14].icell.PDM Vbias 0.03943f
C66 XA.XIR[5].XIC[8].icell.Ien VPWR 0.1979f
C67 XA.XIR[8].XIC_dummy_right.icell.Iout XA.XIR[9].XIC_dummy_right.icell.Iout 0.04047f
C68 XA.XIR[10].XIC_dummy_left.icell.Iout VPWR 0.11267f
C69 XA.XIR[9].XIC[12].icell.Ien Vbias 0.19161f
C70 XThC.Tn[8] XA.XIR[14].XIC[8].icell.Ien 0.03605f
C71 XThC.Tn[0] XA.XIR[11].XIC[0].icell.Ien 0.03605f
C72 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.PDM 0.02104f
C73 XA.XIR[4].XIC[11].icell.PUM VPWR 0.01015f
C74 XA.XIR[5].XIC[4].icell.Ien Iout 0.06821f
C75 XThC.XTB6.A XThC.XTB7.Y 0.01596f
C76 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.PDM 0.02104f
C77 XA.XIR[0].XIC[5].icell.Ien Vbias 0.19209f
C78 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PDM 0.02765f
C79 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.PDM 0.02104f
C80 XA.XIR[8].XIC[5].icell.PUM VPWR 0.01015f
C81 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PDM 0.02765f
C82 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.PDM 0.02104f
C83 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PDM 0.02765f
C84 XA.XIR[12].XIC[3].icell.Ien VPWR 0.1979f
C85 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PDM 0.02816f
C86 XA.XIR[14].XIC[14].icell.Ien VPWR 0.19851f
C87 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.Ien 0.04854f
C88 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PDM 0.04035f
C89 XA.XIR[7].XIC[8].icell.Ien Vbias 0.19161f
C90 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PDM 0.02765f
C91 XThC.Tn[4] XThR.Tn[13] 0.29362f
C92 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PDM 0.02765f
C93 XA.XIR[9].XIC[14].icell.PUM VPWR 0.01015f
C94 XThR.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.15202f
C95 XA.XIR[1].XIC_dummy_left.icell.Iout Iout 0.0353f
C96 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.PDM 0.02104f
C97 XThC.XTB2.Y a_3773_9615# 0.2342f
C98 XThC.Tn[7] Iout 0.84285f
C99 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.PDM 0.02104f
C100 XThC.Tn[7] XThR.Tn[9] 0.29362f
C101 XThC.Tn[3] XThR.Tn[8] 0.29362f
C102 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.0404f
C103 XThC.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.03605f
C104 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.Ien 0.04854f
C105 XThR.Tn[10] XA.XIR[10].XIC[13].icell.Ien 0.15202f
C106 XA.XIR[7].XIC[10].icell.PUM VPWR 0.01015f
C107 XA.XIR[11].XIC[10].icell.Ien VPWR 0.1979f
C108 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.PDM 0.02104f
C109 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PDM 0.04035f
C110 XA.XIR[10].XIC[0].icell.Ien Vbias 0.19149f
C111 XA.XIR[14].XIC[11].icell.PUM VPWR 0.01015f
C112 XA.XIR[6].XIC[5].icell.PDM Vbias 0.03922f
C113 VPWR data[3] 0.20846f
C114 XThR.Tn[12] XA.XIR[12].XIC[2].icell.Ien 0.15202f
C115 XThC.XTBN.A VPWR 0.88811f
C116 XA.XIR[14].XIC[2].icell.PDM Vbias 0.03922f
C117 XThR.Tn[3] XA.XIR[3].XIC[7].icell.Ien 0.15202f
C118 XA.XIR[5].XIC[12].icell.PDM Vbias 0.03922f
C119 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.PDM 0.02104f
C120 XA.XIR[2].XIC[1].icell.PUM VPWR 0.01015f
C121 XThC.Tn[0] XThC.Tn[2] 0.12858f
C122 XA.XIR[13].XIC[6].icell.PDM Vbias 0.03922f
C123 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.PDM 0.02104f
C124 XA.XIR[11].XIC[0].icell.Ien VPWR 0.1979f
C125 XThC.Tn[5] XThC.Tn[6] 0.30991f
C126 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PDM 0.04035f
C127 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PDM 0.02765f
C128 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR 0.08221f
C129 XA.XIR[10].XIC[2].icell.PUM VPWR 0.01015f
C130 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.PDM 0.02104f
C131 XThR.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.15202f
C132 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR 0.35722f
C133 XThR.Tn[14] XA.XIR[14].XIC_15.icell.Ien 0.13564f
C134 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.PDM 0.02104f
C135 XA.XIR[15].XIC[0].icell.PDM VPWR 0.01334f
C136 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.Ien 0.04854f
C137 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR 0.08209f
C138 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.PDM 0.02104f
C139 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.PDM 0.02104f
C140 XA.XIR[14].XIC[12].icell.Ien VPWR 0.19845f
C141 XA.XIR[3].XIC[5].icell.Ien Vbias 0.19161f
C142 XThC.Tn[2] XA.XIR[9].XIC[2].icell.Ien 0.03605f
C143 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.PDM 0.02104f
C144 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PDM 0.02765f
C145 XThC.Tn[9] XA.XIR[0].XIC[9].icell.Ien 0.03754f
C146 XA.XIR[6].XIC_dummy_left.icell.Iout Iout 0.0353f
C147 XThC.XTB7.Y XThC.Tn[8] 0.07806f
C148 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.Ien 0.04854f
C149 XThC.Tn[12] Vbias 1.17777f
C150 XA.XIR[9].XIC[4].icell.Ien VPWR 0.1979f
C151 XThR.Tn[0] XThR.Tn[1] 0.25949f
C152 XThC.Tn[3] XA.XIR[1].XIC[3].icell.Ien 0.03605f
C153 XA.XIR[3].XIC[7].icell.PDM Vbias 0.03922f
C154 XA.XIR[4].XIC[14].icell.Ien Vbias 0.19161f
C155 XA.XIR[8].XIC[9].icell.PDM Vbias 0.03922f
C156 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.Ien 0.04854f
C157 XA.XIR[13].XIC_dummy_left.icell.Iout VPWR 0.11153f
C158 XA.XIR[2].XIC[13].icell.PDM Vbias 0.03922f
C159 XThR.Tn[10] XA.XIR[10].XIC[11].icell.Ien 0.15202f
C160 XA.XIR[8].XIC[8].icell.Ien Vbias 0.19161f
C161 XThR.XTB7.A XThR.XTB5.Y 0.11935f
C162 XA.XIR[3].XIC[7].icell.PUM VPWR 0.01015f
C163 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PDM 0.02765f
C164 XA.XIR[10].XIC_15.icell.PDM Vbias 0.03927f
C165 XThC.Tn[11] XA.XIR[4].XIC[11].icell.Ien 0.03605f
C166 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Iout 0.01728f
C167 XA.XIR[5].XIC[13].icell.Ien VPWR 0.1979f
C168 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.PDM 0.02104f
C169 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Iout 0.01728f
C170 XThC.XTB3.Y VPWR 1.07065f
C171 XA.XIR[5].XIC[9].icell.Ien Iout 0.06821f
C172 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR 0.01691f
C173 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.02765f
C174 XThC.XTB1.Y XThC.Tn[0] 0.18574f
C175 XThC.Tn[14] XThR.Tn[3] 0.29368f
C176 XThC.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.03605f
C177 XThC.Tn[2] VPWR 6.49267f
C178 XA.XIR[0].XIC[10].icell.Ien Vbias 0.19209f
C179 XThC.XTBN.A a_9827_9569# 0.09118f
C180 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PDM 0.04035f
C181 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PDM 0.04035f
C182 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.PDM 0.02104f
C183 XA.XIR[8].XIC[10].icell.PUM VPWR 0.01015f
C184 XA.XIR[11].XIC_15.icell.PDM VPWR 0.07527f
C185 XA.XIR[11].XIC_15.icell.Ien VPWR 0.26829f
C186 XA.XIR[12].XIC[8].icell.Ien VPWR 0.1979f
C187 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.Ien 0.04854f
C188 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR 0.35722f
C189 XThC.Tn[8] XThR.Tn[0] 0.29427f
C190 XA.XIR[12].XIC[4].icell.Ien Iout 0.06821f
C191 XThC.Tn[10] XThR.Tn[5] 0.29362f
C192 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.Ien 0.04854f
C193 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.PDM 0.02104f
C194 XA.XIR[7].XIC[13].icell.Ien Vbias 0.19161f
C195 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.Ien 0.04854f
C196 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.PDM 0.02104f
C197 XThR.Tn[4] XA.XIR[4].XIC[9].icell.Ien 0.15202f
C198 XThC.Tn[0] XA.XIR[7].XIC[0].icell.Ien 0.03605f
C199 XA.XIR[14].XIC[10].icell.Ien VPWR 0.19845f
C200 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.Ien 0.04854f
C201 XThC.XTB5.Y a_5155_9615# 0.24821f
C202 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.Ien 0.04854f
C203 XA.XIR[13].XIC[0].icell.Ien Vbias 0.19149f
C204 XThC.XTB7.A a_4067_9615# 0.0127f
C205 XThR.XTB1.Y XThR.XTB7.A 0.48957f
C206 XThC.XTBN.A XThC.XTB7.B 0.35142f
C207 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PDM 0.04056f
C208 XA.XIR[11].XIC_dummy_right.icell.Iout VPWR 0.11567f
C209 XThC.Tn[3] XA.XIR[6].XIC[3].icell.Ien 0.03605f
C210 XA.XIR[7].XIC_15.icell.PUM VPWR 0.01655f
C211 XThR.Tn[7] XA.XIR[7].XIC[2].icell.Ien 0.15202f
C212 XA.XIR[7].XIC[13].icell.PDM Vbias 0.03922f
C213 XThC.Tn[9] XA.XIR[3].XIC[9].icell.Ien 0.03605f
C214 XA.XIR[4].XIC[1].icell.Ien VPWR 0.1979f
C215 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR 0.08252f
C216 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.Ien 0.04854f
C217 XThC.Tn[4] XA.XIR[12].XIC[4].icell.Ien 0.03605f
C218 XA.XIR[13].XIC[2].icell.PUM VPWR 0.01015f
C219 XThR.Tn[12] XA.XIR[12].XIC[7].icell.Ien 0.15202f
C220 XThC.XTBN.Y a_5155_9615# 0.07602f
C221 XThR.Tn[3] XA.XIR[3].XIC[12].icell.Ien 0.15202f
C222 XThC.XTB1.Y VPWR 1.1176f
C223 XA.XIR[9].XIC[9].icell.PDM Vbias 0.03922f
C224 XThC.XTB5.Y XThC.XTB6.Y 2.12831f
C225 XA.XIR[0].XIC[1].icell.PDM Vbias 0.03943f
C226 XA.XIR[15].XIC[3].icell.Ien VPWR 0.33655f
C227 XThR.Tn[7] Iout 1.19572f
C228 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PDM 0.02765f
C229 XA.XIR[10].XIC_dummy_right.icell.Iout XA.XIR[11].XIC_dummy_right.icell.Iout 0.04047f
C230 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.02765f
C231 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PDM 0.02765f
C232 XThR.Tn[2] XA.XIR[2].XIC[7].icell.Ien 0.15202f
C233 XA.XIR[4].XIC[6].icell.Ien VPWR 0.1979f
C234 XThC.XTB7.A XThC.Tn[3] 0.03065f
C235 XThR.Tn[1] XA.XIR[1].XIC[0].icell.Ien 0.1525f
C236 XA.XIR[14].XIC_dummy_left.icell.Ien XThR.Tn[14] 0.01432f
C237 XA.XIR[4].XIC[2].icell.Ien Iout 0.06821f
C238 XThR.XTB7.B XThR.XTB5.Y 0.30227f
C239 a_2979_9615# XThC.Tn[0] 0.2829f
C240 VPWR bias[2] 1.20331f
C241 XA.XIR[3].XIC[10].icell.Ien Vbias 0.19161f
C242 XA.XIR[1].XIC[14].icell.PDM Vbias 0.03922f
C243 XA.XIR[10].XIC[14].icell.PDM Vbias 0.03922f
C244 XThC.Tn[12] XThR.Tn[6] 0.29362f
C245 XA.XIR[7].XIC[0].icell.Ien VPWR 0.1979f
C246 XA.XIR[0].XIC[5].icell.PDM VPWR 0.01101f
C247 XThC.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.03605f
C248 XA.XIR[2].XIC[3].icell.Ien Vbias 0.19161f
C249 XA.XIR[4].XIC[14].icell.PDM Vbias 0.03922f
C250 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.Ien 0.04854f
C251 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.PDM 0.02104f
C252 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.PDM 0.02104f
C253 XThC.XTB6.Y XThC.XTBN.Y 0.18947f
C254 XA.XIR[1].XIC[2].icell.PUM VPWR 0.01015f
C255 XA.XIR[13].XIC_15.icell.PDM Vbias 0.03927f
C256 XA.XIR[9].XIC[9].icell.Ien VPWR 0.1979f
C257 XA.XIR[10].XIC[3].icell.PUM VPWR 0.01015f
C258 XA.XIR[1].XIC[5].icell.Ien Vbias 0.19173f
C259 XThC.Tn[14] XThR.Tn[11] 0.29368f
C260 XA.XIR[9].XIC[5].icell.Ien Iout 0.06821f
C261 XThR.Tn[9] XA.XIR[9].XIC[5].icell.Ien 0.15202f
C262 XThC.XTB3.Y XThC.XTB7.B 0.23315f
C263 XThC.XTB4.Y XThC.XTB5.Y 2.06459f
C264 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PDM 0.04035f
C265 XA.XIR[0].XIC[2].icell.Ien VPWR 0.19726f
C266 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.Ien 0.04854f
C267 XThC.Tn[4] XThR.Tn[7] 0.29362f
C268 XA.XIR[11].XIC[14].icell.PDM VPWR 0.01002f
C269 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PDM 0.04035f
C270 XA.XIR[8].XIC[13].icell.Ien Vbias 0.19161f
C271 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PDM 0.04035f
C272 XA.XIR[3].XIC[12].icell.PUM VPWR 0.01015f
C273 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.02774f
C274 XThC.XTB7.Y XThC.Tn[6] 0.2144f
C275 XThC.Tn[1] Vbias 1.09737f
C276 XA.XIR[14].XIC_15.icell.PDM VPWR 0.07527f
C277 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.PDM 0.02104f
C278 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PDM 0.02765f
C279 XA.XIR[14].XIC_15.icell.Ien VPWR 0.26861f
C280 XA.XIR[2].XIC[5].icell.PUM VPWR 0.01015f
C281 XA.XIR[7].XIC[5].icell.Ien VPWR 0.1979f
C282 XThC.XTB6.Y XThC.Tn[10] 0.02461f
C283 XThC.Tn[10] XA.XIR[5].XIC[10].icell.Ien 0.03605f
C284 XA.XIR[5].XIC[14].icell.Ien Iout 0.06821f
C285 XA.XIR[1].XIC[7].icell.PUM VPWR 0.01015f
C286 XThC.Tn[8] XThR.Tn[1] 0.29362f
C287 XThR.Tn[0] XA.XIR[0].XIC[1].icell.Ien 0.15202f
C288 XA.XIR[0].XIC_15.icell.Ien Vbias 0.19241f
C289 XThR.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.15202f
C290 XThR.XTB7.B XThR.XTB1.Y 1.61695f
C291 XA.XIR[8].XIC_15.icell.PUM VPWR 0.01655f
C292 XThC.Tn[8] XThR.Tn[12] 0.29362f
C293 XThC.XTB4.Y XThC.XTBN.Y 0.15636f
C294 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PDM 0.02765f
C295 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.Ien 0.04854f
C296 XA.XIR[12].XIC[9].icell.Ien Iout 0.06821f
C297 XA.XIR[6].XIC[0].icell.Ien Vbias 0.19149f
C298 XThC.Tn[3] XThR.Tn[3] 0.29362f
C299 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.PDM 0.02104f
C300 XA.XIR[14].XIC[0].icell.PUM VPWR 0.01015f
C301 XThC.Tn[12] XThR.Tn[4] 0.29362f
C302 XA.XIR[14].XIC_dummy_right.icell.Iout VPWR 0.11567f
C303 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PDM 0.04056f
C304 XThC.Tn[14] XA.XIR[10].XIC[14].icell.Ien 0.03605f
C305 XThR.Tn[4] XA.XIR[4].XIC[14].icell.Ien 0.15202f
C306 a_2979_9615# VPWR 0.70527f
C307 XA.XIR[9].XIC[0].icell.Ien Iout 0.06814f
C308 XA.XIR[11].XIC[4].icell.PDM Vbias 0.03922f
C309 XThR.Tn[0] XA.XIR[0].XIC[6].icell.Ien 0.15202f
C310 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9] 0.15202f
C311 XThR.Tn[10] XA.XIR[10].XIC[5].icell.Ien 0.15202f
C312 XThC.XTB4.Y XThC.Tn[10] 0.01391f
C313 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PDM 0.04035f
C314 XA.XIR[10].XIC[8].icell.PDM Vbias 0.03922f
C315 XThC.Tn[12] XA.XIR[11].XIC[12].icell.Ien 0.03605f
C316 XThC.Tn[6] XThR.Tn[0] 0.29373f
C317 XThC.XTB4.Y a_4861_9615# 0.23756f
C318 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PDM 0.02765f
C319 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PDM 0.0404f
C320 XA.XIR[6].XIC[2].icell.PUM VPWR 0.01015f
C321 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.Ien 0.04854f
C322 XThR.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.15202f
C323 XA.XIR[6].XIC[5].icell.Ien Vbias 0.19161f
C324 XThC.Tn[12] XThC.Tn[13] 0.23689f
C325 XThC.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.03605f
C326 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PDM 0.02765f
C327 XThC.XTB2.Y XThC.XTB5.Y 0.0451f
C328 XThC.XTB1.Y XThC.XTB7.B 1.61695f
C329 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PDM 0.02765f
C330 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.02765f
C331 XThR.XTBN.Y XThR.XTB5.Y 0.16186f
C332 XA.XIR[2].XIC[0].icell.PDM Vbias 0.03915f
C333 XThC.Tn[9] XA.XIR[1].XIC[9].icell.Ien 0.03605f
C334 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PDM 0.04042f
C335 XA.XIR[3].XIC[2].icell.Ien VPWR 0.1979f
C336 XA.XIR[10].XIC[13].icell.PDM Vbias 0.03922f
C337 XA.XIR[6].XIC[7].icell.PUM VPWR 0.01015f
C338 XThC.Tn[0] XA.XIR[8].XIC[0].icell.Ien 0.03605f
C339 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.PDM 0.02104f
C340 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PDM 0.02765f
C341 XA.XIR[15].XIC[8].icell.Ien VPWR 0.33655f
C342 XA.XIR[11].XIC[4].icell.Ien Vbias 0.19161f
C343 XThC.XTBN.Y a_7875_9569# 0.229f
C344 XA.XIR[13].XIC[14].icell.PDM Vbias 0.03922f
C345 XThR.Tn[2] XA.XIR[2].XIC[12].icell.Ien 0.15202f
C346 XA.XIR[15].XIC[4].icell.Ien Iout 0.07211f
C347 XThR.Tn[13] XA.XIR[13].XIC[11].icell.Ien 0.15202f
C348 XA.XIR[4].XIC[11].icell.Ien VPWR 0.1979f
C349 XA.XIR[10].XIC[6].icell.Ien Vbias 0.19161f
C350 XThC.XTB2.Y XThC.XTBN.Y 0.2075f
C351 XThC.Tn[5] XThR.Tn[2] 0.29362f
C352 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.PDM 0.02104f
C353 XThR.XTB4.Y XThR.XTB5.Y 2.06459f
C354 XA.XIR[4].XIC[7].icell.Ien Iout 0.06821f
C355 XA.XIR[13].XIC[3].icell.PUM VPWR 0.01015f
C356 XThC.Tn[14] XThR.Tn[14] 0.29368f
C357 XA.XIR[8].XIC[5].icell.Ien VPWR 0.1979f
C358 XA.XIR[3].XIC_15.icell.Ien Vbias 0.19195f
C359 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Iout 0.01728f
C360 XThR.XTB5.Y XThR.Tn[10] 0.01742f
C361 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.Ien 0.04854f
C362 XThC.Tn[13] XA.XIR[7].XIC[13].icell.Ien 0.03605f
C363 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.Ien 0.04854f
C364 XA.XIR[14].XIC[14].icell.PDM VPWR 0.01002f
C365 XA.XIR[11].XIC[6].icell.PUM VPWR 0.01015f
C366 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PDM 0.04035f
C367 XA.XIR[2].XIC[8].icell.Ien Vbias 0.19161f
C368 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout 0.06446f
C369 XA.XIR[7].XIC[1].icell.Ien Iout 0.06821f
C370 XA.XIR[9].XIC[14].icell.Ien VPWR 0.19796f
C371 XA.XIR[1].XIC[10].icell.Ien Vbias 0.19173f
C372 XA.XIR[10].XIC[8].icell.PUM VPWR 0.01015f
C373 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.PDM 0.02104f
C374 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PDM 0.02765f
C375 XA.XIR[9].XIC[10].icell.Ien Iout 0.06821f
C376 XThR.Tn[9] XA.XIR[9].XIC[10].icell.Ien 0.15202f
C377 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.Ien 0.04854f
C378 XThR.XTB1.Y XThR.XTBN.Y 0.20262f
C379 XA.XIR[0].XIC[7].icell.Ien VPWR 0.19725f
C380 XA.XIR[12].XIC[14].icell.Ien Iout 0.06821f
C381 XThC.Tn[1] XThR.Tn[6] 0.29362f
C382 XA.XIR[0].XIC[3].icell.Ien Iout 0.06775f
C383 XThC.Tn[4] XA.XIR[15].XIC[4].icell.Ien 0.03184f
C384 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PDM 0.04035f
C385 XThC.XTBN.A XThC.Tn[12] 0.22686f
C386 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR 0.35722f
C387 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.PDM 0.02104f
C388 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.04035f
C389 XThR.Tn[5] a_n1049_5611# 0.27042f
C390 XA.XIR[2].XIC[10].icell.PUM VPWR 0.01015f
C391 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PDM 0.02765f
C392 XA.XIR[7].XIC[10].icell.Ien VPWR 0.1979f
C393 XA.XIR[0].XIC_dummy_right.icell.Iout XA.XIR[1].XIC_dummy_right.icell.Iout 0.04047f
C394 XThC.Tn[3] XThR.Tn[11] 0.29362f
C395 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR 0.38903f
C396 XA.XIR[7].XIC[6].icell.Ien Iout 0.06821f
C397 XA.XIR[1].XIC[12].icell.PUM VPWR 0.01015f
C398 XThC.Tn[5] XA.XIR[11].XIC[5].icell.Ien 0.03605f
C399 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PDM 0.04035f
C400 XA.XIR[7].XIC[0].icell.PDM Vbias 0.03915f
C401 XThC.Tn[9] XA.XIR[6].XIC[9].icell.Ien 0.03605f
C402 XThR.XTB1.Y XThR.XTB4.Y 0.05121f
C403 XA.XIR[6].XIC[7].icell.PDM Vbias 0.03922f
C404 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.Ien 0.04854f
C405 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.PDM 0.02104f
C406 XThR.Tn[6] XA.XIR[6].XIC[0].icell.Ien 0.15202f
C407 XA.XIR[8].XIC[0].icell.Ien VPWR 0.1979f
C408 XThC.Tn[14] XA.XIR[13].XIC[14].icell.Ien 0.03605f
C409 XA.XIR[14].XIC[4].icell.PDM Vbias 0.03922f
C410 XA.XIR[5].XIC[14].icell.PDM Vbias 0.03922f
C411 a_10915_9569# XThC.Tn[13] 0.01061f
C412 XThC.XTB5.Y XThC.Tn[4] 0.19958f
C413 XThC.Tn[12] XA.XIR[14].XIC[12].icell.Ien 0.03605f
C414 XA.XIR[13].XIC[8].icell.PDM Vbias 0.03922f
C415 XThR.Tn[11] XA.XIR[11].XIC[6].icell.Ien 0.15202f
C416 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.Ien 0.04854f
C417 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PDM 0.04035f
C418 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PDM 0.02765f
C419 XThC.Tn[6] XThR.Tn[1] 0.29364f
C420 XThR.XTB6.A XThR.XTB7.A 0.44014f
C421 XThC.Tn[10] Iout 0.84085f
C422 XA.XIR[12].XIC_dummy_left.icell.Iout XA.XIR[13].XIC_dummy_left.icell.Iout 0.03665f
C423 XThC.Tn[10] XThR.Tn[9] 0.29362f
C424 XA.XIR[15].XIC[2].icell.PDM VPWR 0.01334f
C425 XThR.Tn[0] XA.XIR[0].XIC[11].icell.Ien 0.15202f
C426 XThC.Tn[6] XThR.Tn[12] 0.29362f
C427 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PDM 0.02765f
C428 XThR.Tn[6] XA.XIR[6].XIC[5].icell.Ien 0.15202f
C429 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.Ien 0.04854f
C430 XThR.XTB5.Y a_n997_1803# 0.06458f
C431 XA.XIR[13].XIC_dummy_right.icell.Iout XA.XIR[14].XIC_dummy_right.icell.Iout 0.04047f
C432 XA.XIR[10].XIC[12].icell.PDM Vbias 0.03922f
C433 XA.XIR[1].XIC[1].icell.PDM Vbias 0.03922f
C434 XThC.Tn[1] XThR.Tn[4] 0.29362f
C435 XThC.XTBN.Y XThC.Tn[4] 0.61061f
C436 XA.XIR[6].XIC[10].icell.Ien Vbias 0.19161f
C437 XThR.Tn[7] XA.XIR[7].XIC[12].icell.Ien 0.15202f
C438 XA.XIR[13].XIC[13].icell.PDM Vbias 0.03922f
C439 XA.XIR[4].XIC[1].icell.PDM Vbias 0.03922f
C440 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR 0.08221f
C441 XA.XIR[12].XIC[12].icell.Ien Iout 0.06821f
C442 XA.XIR[3].XIC[9].icell.PDM Vbias 0.03922f
C443 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PDM 0.02765f
C444 XA.XIR[8].XIC[11].icell.PDM Vbias 0.03922f
C445 XA.XIR[14].XIC[4].icell.Ien Vbias 0.19161f
C446 XThC.Tn[13] XA.XIR[8].XIC[13].icell.Ien 0.03605f
C447 XThC.Tn[5] XThR.Tn[10] 0.29362f
C448 XThC.Tn[0] XA.XIR[5].XIC[0].icell.Ien 0.03605f
C449 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.Ien 0.04854f
C450 XA.XIR[2].XIC_15.icell.PDM Vbias 0.03927f
C451 XA.XIR[13].XIC[6].icell.Ien Vbias 0.19161f
C452 XA.XIR[3].XIC[7].icell.Ien VPWR 0.1979f
C453 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.Ien 0.04854f
C454 XA.XIR[8].XIC[1].icell.Ien Iout 0.06821f
C455 XA.XIR[6].XIC[12].icell.PUM VPWR 0.01015f
C456 XA.XIR[3].XIC[3].icell.Ien Iout 0.06821f
C457 XA.XIR[11].XIC[9].icell.Ien Vbias 0.19161f
C458 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PDM 0.04035f
C459 XA.XIR[15].XIC[9].icell.Ien Iout 0.07211f
C460 XA.XIR[1].XIC[2].icell.Ien VPWR 0.1979f
C461 XA.XIR[8].XIC_15.icell.PDM VPWR 0.07527f
C462 XA.XIR[14].XIC[6].icell.PUM VPWR 0.01015f
C463 XThC.Tn[7] XA.XIR[2].XIC[7].icell.Ien 0.03605f
C464 XA.XIR[4].XIC[12].icell.Ien Iout 0.06821f
C465 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PDM 0.04035f
C466 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PDM 0.04035f
C467 XA.XIR[13].XIC[8].icell.PUM VPWR 0.01015f
C468 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.PDM 0.02104f
C469 XA.XIR[8].XIC[10].icell.Ien VPWR 0.1979f
C470 XA.XIR[8].XIC[6].icell.Ien Iout 0.06821f
C471 XA.XIR[2].XIC[13].icell.Ien Vbias 0.19161f
C472 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR 0.01604f
C473 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR 0.35722f
C474 XA.XIR[1].XIC_15.icell.Ien Vbias 0.19206f
C475 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PDM 0.04035f
C476 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.PDM 0.02104f
C477 XThC.Tn[3] XThR.Tn[14] 0.29362f
C478 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.PDM 0.02104f
C479 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PDM 0.02765f
C480 XA.XIR[9].XIC_15.icell.Ien Iout 0.0694f
C481 XThR.Tn[9] XA.XIR[9].XIC_15.icell.Ien 0.13564f
C482 XA.XIR[0].XIC[12].icell.Ien VPWR 0.19971f
C483 XThC.Tn[5] XA.XIR[14].XIC[5].icell.Ien 0.03605f
C484 XThC.XTB7.A a_5155_9615# 0.02287f
C485 XA.XIR[0].XIC[8].icell.Ien Iout 0.06775f
C486 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.PDM 0.02104f
C487 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.PDM 0.02104f
C488 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PDM 0.04039f
C489 XA.XIR[2].XIC_15.icell.PUM VPWR 0.01655f
C490 XA.XIR[7].XIC_15.icell.Ien VPWR 0.26829f
C491 XA.XIR[12].XIC[10].icell.Ien Iout 0.06821f
C492 XThR.Tn[13] XA.XIR[13].XIC[5].icell.Ien 0.15202f
C493 XA.XIR[5].XIC[0].icell.Ien VPWR 0.1979f
C494 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.PDM 0.02104f
C495 XA.XIR[5].XIC[3].icell.Ien Vbias 0.19161f
C496 XA.XIR[7].XIC_15.icell.PDM Vbias 0.03927f
C497 XThR.XTB7.B XThR.XTB6.A 1.47641f
C498 XThR.XTB5.A XThR.XTB2.Y 0.02203f
C499 XA.XIR[7].XIC[11].icell.Ien Iout 0.06821f
C500 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.Ien 0.04854f
C501 XA.XIR[14].XIC[1].icell.PUM VPWR 0.01015f
C502 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.PDM 0.02104f
C503 XA.XIR[4].XIC_dummy_left.icell.Iout VPWR 0.1106f
C504 XThC.Tn[14] VPWR 7.41153f
C505 XThC.XTBN.Y a_6243_9615# 0.07731f
C506 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PDM 0.02765f
C507 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.PDM 0.02104f
C508 XA.XIR[9].XIC_dummy_right.icell.Iout Iout 0.01732f
C509 XA.XIR[10].XIC[11].icell.PDM Vbias 0.03922f
C510 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout 0.06446f
C511 XA.XIR[3].XIC[0].icell.Ien Iout 0.06814f
C512 XThR.Tn[8] Iout 1.19572f
C513 XThR.Tn[8] XThR.Tn[9] 0.09382f
C514 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.Ien 0.04854f
C515 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR 0.08221f
C516 XA.XIR[6].XIC[2].icell.Ien VPWR 0.1979f
C517 XA.XIR[9].XIC[11].icell.PDM Vbias 0.03922f
C518 XA.XIR[13].XIC[12].icell.PDM Vbias 0.03922f
C519 XA.XIR[0].XIC[3].icell.PDM Vbias 0.03938f
C520 XA.XIR[11].XIC[1].icell.Ien Iout 0.06821f
C521 XA.XIR[5].XIC[5].icell.PUM VPWR 0.01015f
C522 XA.XIR[7].XIC_dummy_right.icell.Iout VPWR 0.11567f
C523 XThC.XTB7.A XThC.XTB6.Y 0.19112f
C524 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Ien 0.01734f
C525 XA.XIR[10].XIC_dummy_left.icell.Ien XThR.Tn[10] 0.01432f
C526 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Ien 0.01785f
C527 XThR.Tn[6] XA.XIR[6].XIC[10].icell.Ien 0.15202f
C528 XThR.XTB2.Y data[5] 0.017f
C529 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.PDM 0.02104f
C530 XA.XIR[11].XIC[14].icell.Ien Vbias 0.19161f
C531 XThR.Tn[6] Vbias 1.44824f
C532 XThC.Tn[5] XThR.Tn[13] 0.29362f
C533 XA.XIR[15].XIC[14].icell.Ien Iout 0.07211f
C534 XA.XIR[6].XIC_15.icell.Ien Vbias 0.19195f
C535 XA.XIR[9].XIC_15.icell.PDM VPWR 0.07527f
C536 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.Ien 0.04854f
C537 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.Ien 0.04854f
C538 XA.XIR[10].XIC[3].icell.Ien VPWR 0.1979f
C539 XThC.Tn[4] XThR.Tn[8] 0.29362f
C540 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.PDM 0.02104f
C541 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.Ien 0.04854f
C542 XA.XIR[14].XIC[9].icell.Ien Vbias 0.19161f
C543 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.PDM 0.02104f
C544 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PDM 0.04035f
C545 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PDM 0.04056f
C546 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PDM 0.04035f
C547 XThC.XTB7.A XThC.XTB4.Y 0.14536f
C548 XA.XIR[3].XIC[12].icell.Ien VPWR 0.1979f
C549 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.PDM 0.02104f
C550 XA.XIR[3].XIC[8].icell.Ien Iout 0.06821f
C551 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.Ien 0.04854f
C552 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.Ien 0.04854f
C553 XA.XIR[2].XIC[5].icell.Ien VPWR 0.1979f
C554 XA.XIR[9].XIC[0].icell.PUM VPWR 0.01015f
C555 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.PDM 0.02104f
C556 XA.XIR[1].XIC[7].icell.Ien VPWR 0.1979f
C557 XThC.XTB6.Y a_5949_9615# 0.26831f
C558 XThR.Tn[8] XA.XIR[8].XIC[2].icell.Ien 0.15202f
C559 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.Ien 0.04854f
C560 XThC.Tn[6] XA.XIR[0].XIC[6].icell.Ien 0.03691f
C561 XThC.Tn[0] XThC.Tn[3] 0.12428f
C562 XThC.Tn[1] XThC.Tn[2] 0.72045f
C563 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.04494f
C564 XA.XIR[1].XIC[3].icell.Ien Iout 0.06821f
C565 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PDM 0.02765f
C566 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.Ien 0.04854f
C567 XA.XIR[8].XIC_15.icell.Ien VPWR 0.26829f
C568 XThR.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.15202f
C569 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PDM 0.02765f
C570 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PDM 0.02765f
C571 XA.XIR[12].XIC_15.icell.Ien Iout 0.0694f
C572 XA.XIR[5].XIC[1].icell.PDM Vbias 0.03922f
C573 XThR.XTB7.A a_n1049_5317# 0.02018f
C574 XA.XIR[8].XIC[11].icell.Ien Iout 0.06821f
C575 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.PDM 0.02104f
C576 XThR.Tn[4] Vbias 1.44824f
C577 XThR.XTBN.Y XThR.XTB6.A 0.03867f
C578 XA.XIR[12].XIC[0].icell.PDM Vbias 0.03915f
C579 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.PDM 0.02104f
C580 a_4067_9615# VPWR 0.70648f
C581 XA.XIR[11].XIC[6].icell.PDM Vbias 0.03922f
C582 a_n997_3755# XThR.Tn[9] 0.19352f
C583 XA.XIR[11].XIC[12].icell.Ien Vbias 0.19161f
C584 XThR.XTB2.Y XThR.Tn[9] 0.292f
C585 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PDM 0.04035f
C586 XA.XIR[15].XIC[12].icell.Ien Iout 0.07211f
C587 XThR.Tn[1] XA.XIR[1].XIC[6].icell.Ien 0.15202f
C588 XThC.XTB7.Y XThC.Tn[9] 0.07413f
C589 XA.XIR[10].XIC[10].icell.PDM Vbias 0.03922f
C590 XThR.Tn[14] XA.XIR[14].XIC[6].icell.Ien 0.15202f
C591 XA.XIR[0].XIC[13].icell.Ien Iout 0.06775f
C592 XThC.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.03605f
C593 XThR.XTBN.Y XThR.Tn[0] 0.55717f
C594 XA.XIR[8].XIC_dummy_right.icell.Iout VPWR 0.11567f
C595 XThC.Tn[13] Vbias 1.09272f
C596 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PDM 0.02765f
C597 XA.XIR[12].XIC_dummy_right.icell.Iout Iout 0.01732f
C598 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.PDM 0.02104f
C599 XA.XIR[13].XIC[11].icell.PDM Vbias 0.03922f
C600 XThR.XTB6.A XThR.XTB4.Y 0.04137f
C601 XA.XIR[5].XIC[8].icell.Ien Vbias 0.19161f
C602 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.Ien 0.04854f
C603 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.Ien 0.04854f
C604 XThC.Tn[1] XA.XIR[4].XIC[1].icell.Ien 0.03605f
C605 XThC.XTB2.Y XThC.XTB7.A 0.2319f
C606 XThC.XTB5.A XThC.XTB4.Y 0.02767f
C607 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.PDM 0.02104f
C608 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.Ien 0.04854f
C609 XA.XIR[14].XIC[1].icell.Ien Iout 0.06821f
C610 XA.XIR[2].XIC[2].icell.PDM Vbias 0.03922f
C611 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PDM 0.04035f
C612 XA.XIR[12].XIC[3].icell.Ien Vbias 0.19161f
C613 XThC.XTB1.Y XThC.Tn[1] 0.02048f
C614 XA.XIR[6].XIC[7].icell.Ien VPWR 0.1979f
C615 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.Ien 0.04854f
C616 XThR.XTB7.A a_n1049_6405# 0.02287f
C617 XA.XIR[14].XIC[14].icell.Ien Vbias 0.19161f
C618 XA.XIR[6].XIC[3].icell.Ien Iout 0.06821f
C619 XThC.Tn[3] VPWR 6.46374f
C620 XA.XIR[5].XIC[10].icell.PUM VPWR 0.01015f
C621 XThC.XTBN.Y a_8963_9569# 0.22784f
C622 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PDM 0.02765f
C623 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.PDM 0.02104f
C624 XA.XIR[12].XIC[14].icell.PUM VPWR 0.01015f
C625 XA.XIR[4].XIC_dummy_left.icell.Iout XA.XIR[5].XIC_dummy_left.icell.Iout 0.03665f
C626 XThR.XTB5.A data[4] 0.14415f
C627 XThC.Tn[9] XThR.Tn[0] 0.29432f
C628 XThC.Tn[11] XThR.Tn[5] 0.29362f
C629 XThR.Tn[6] XA.XIR[6].XIC_15.icell.Ien 0.13564f
C630 XThC.Tn[6] XA.XIR[3].XIC[6].icell.Ien 0.03605f
C631 XThR.Tn[1] XThR.Tn[2] 0.14094f
C632 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.PDM 0.02104f
C633 XA.XIR[13].XIC[3].icell.Ien VPWR 0.1979f
C634 XThR.XTB1.Y a_n997_3979# 0.06353f
C635 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.PDM 0.02104f
C636 XThC.Tn[13] XA.XIR[2].XIC[13].icell.Ien 0.03605f
C637 XA.XIR[12].XIC[5].icell.PUM VPWR 0.01015f
C638 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.Ien 0.04854f
C639 XA.XIR[11].XIC[6].icell.Ien VPWR 0.1979f
C640 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PDM 0.04035f
C641 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR 0.38914f
C642 XA.XIR[2].XIC[1].icell.Ien Iout 0.06821f
C643 XA.XIR[11].XIC[10].icell.Ien Vbias 0.19161f
C644 XA.XIR[7].XIC_dummy_left.icell.Iout Iout 0.0353f
C645 XA.XIR[10].XIC[8].icell.Ien VPWR 0.1979f
C646 XA.XIR[11].XIC[2].icell.Ien Iout 0.06821f
C647 XA.XIR[15].XIC[10].icell.Ien Iout 0.07211f
C648 XA.XIR[10].XIC[4].icell.Ien Iout 0.06821f
C649 XThC.XTBN.A Vbias 0.01661f
C650 XThR.XTB7.B a_n1049_5317# 0.01743f
C651 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PDM 0.04035f
C652 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PDM 0.02765f
C653 data[5] data[4] 0.64735f
C654 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.PDM 0.02104f
C655 XA.XIR[3].XIC[13].icell.Ien Iout 0.06821f
C656 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.Ien 0.04854f
C657 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PDM 0.04035f
C658 VPWR data[6] 0.21221f
C659 XThR.Tn[11] XA.XIR[11].XIC_dummy_left.icell.Iout 0.0404f
C660 XThR.Tn[5] XA.XIR[5].XIC[1].icell.Ien 0.15202f
C661 XA.XIR[2].XIC[10].icell.Ien VPWR 0.1979f
C662 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.PDM 0.02104f
C663 XA.XIR[11].XIC[0].icell.Ien Vbias 0.19149f
C664 XThC.XTB5.A XThC.XTB2.Y 0.02203f
C665 XThC.Tn[8] XThR.Tn[2] 0.29362f
C666 XA.XIR[2].XIC[6].icell.Ien Iout 0.06821f
C667 XThR.Tn[8] XA.XIR[8].XIC[7].icell.Ien 0.15202f
C668 XA.XIR[1].XIC[12].icell.Ien VPWR 0.1979f
C669 XA.XIR[7].XIC[2].icell.PDM Vbias 0.03922f
C670 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PDM 0.04035f
C671 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.Ien 0.04854f
C672 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.Ien 0.04854f
C673 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PDM 0.02765f
C674 XA.XIR[1].XIC[8].icell.Ien Iout 0.06821f
C675 XA.XIR[6].XIC[9].icell.PDM Vbias 0.03922f
C676 XA.XIR[15].XIC[0].icell.PDM Vbias 0.03915f
C677 XA.XIR[14].XIC[6].icell.PDM Vbias 0.03922f
C678 XA.XIR[14].XIC[12].icell.Ien Vbias 0.19161f
C679 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.PDM 0.02104f
C680 XA.XIR[13].XIC[10].icell.PDM Vbias 0.03922f
C681 XThC.XTB7.A XThC.Tn[4] 0.0274f
C682 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.PDM 0.02104f
C683 XThC.Tn[4] XA.XIR[10].XIC[4].icell.Ien 0.03605f
C684 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PDM 0.02765f
C685 XThR.Tn[5] XA.XIR[5].XIC[6].icell.Ien 0.15202f
C686 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PDM 0.04035f
C687 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR 0.35722f
C688 XThR.XTB6.Y XThR.XTBN.A 0.06405f
C689 XA.XIR[12].XIC[12].icell.PUM VPWR 0.01015f
C690 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.PDM 0.02104f
C691 XThR.XTBN.Y XThR.Tn[1] 0.61094f
C692 a_2979_9615# XThC.Tn[1] 0.01205f
C693 XA.XIR[9].XIC[4].icell.Ien Vbias 0.19161f
C694 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.Ien 0.04854f
C695 XA.XIR[4].XIC[3].icell.PUM VPWR 0.01015f
C696 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.Ien 0.04854f
C697 XA.XIR[15].XIC[4].icell.PDM VPWR 0.01334f
C698 XThC.Tn[7] XA.XIR[5].XIC[7].icell.Ien 0.03605f
C699 XThC.Tn[13] XThR.Tn[6] 0.29363f
C700 XThR.XTBN.Y XThR.Tn[12] 0.50762f
C701 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.PDM 0.02104f
C702 XThR.Tn[1] XA.XIR[1].XIC[11].icell.Ien 0.15202f
C703 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.PDM 0.02104f
C704 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PDM 0.02765f
C705 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.PDM 0.02104f
C706 XA.XIR[1].XIC[3].icell.PDM Vbias 0.03922f
C707 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.PDM 0.02104f
C708 XA.XIR[13].XIC_dummy_left.icell.Ien XThR.Tn[13] 0.01432f
C709 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.Ien 0.04854f
C710 XA.XIR[4].XIC[3].icell.PDM Vbias 0.03922f
C711 XThC.Tn[3] XA.XIR[7].XIC[3].icell.Ien 0.03605f
C712 XA.XIR[5].XIC[13].icell.Ien Vbias 0.19161f
C713 XThC.Tn[5] XThR.Tn[7] 0.29362f
C714 XThR.Tn[3] Iout 1.19576f
C715 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.PDM 0.02104f
C716 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR 0.08221f
C717 XA.XIR[9].XIC[6].icell.PUM VPWR 0.01015f
C718 XThC.XTB3.Y Vbias 0.01225f
C719 XA.XIR[12].XIC[13].icell.Ien VPWR 0.1979f
C720 XA.XIR[3].XIC[11].icell.PDM Vbias 0.03922f
C721 XA.XIR[8].XIC[13].icell.PDM Vbias 0.03922f
C722 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PDM 0.02765f
C723 XThC.XTB7.Y XThC.Tn[7] 0.0835f
C724 XThC.Tn[2] Vbias 1.30848f
C725 XThC.XTB6.Y XThC.Tn[11] 0.02513f
C726 XThR.XTB7.Y XThR.Tn[9] 0.07413f
C727 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PDM 0.04035f
C728 XA.XIR[11].XIC_15.icell.PDM Vbias 0.03927f
C729 XA.XIR[11].XIC_15.icell.Ien Vbias 0.19195f
C730 XA.XIR[8].XIC_dummy_left.icell.Iout Iout 0.0353f
C731 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Iout 0.01728f
C732 XA.XIR[6].XIC[12].icell.Ien VPWR 0.1979f
C733 XA.XIR[12].XIC[8].icell.Ien Vbias 0.19161f
C734 XThC.Tn[9] XThR.Tn[1] 0.29362f
C735 XA.XIR[15].XIC_15.icell.Ien Iout 0.0733f
C736 XA.XIR[6].XIC[8].icell.Ien Iout 0.06821f
C737 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.PDM 0.02104f
C738 XA.XIR[5].XIC_15.icell.PUM VPWR 0.01655f
C739 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PDM 0.04035f
C740 XThC.Tn[9] XThR.Tn[12] 0.29362f
C741 XA.XIR[3].XIC_15.icell.PDM VPWR 0.07527f
C742 XA.XIR[14].XIC[6].icell.Ien VPWR 0.19845f
C743 XA.XIR[14].XIC[10].icell.Ien Vbias 0.19161f
C744 XThR.XTBN.Y a_n1049_5317# 0.07731f
C745 XThC.Tn[5] XA.XIR[9].XIC[5].icell.Ien 0.03605f
C746 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PDM 0.04035f
C747 XA.XIR[14].XIC[2].icell.Ien Iout 0.06821f
C748 XA.XIR[13].XIC[8].icell.Ien VPWR 0.1979f
C749 XThC.Tn[4] XThR.Tn[3] 0.29362f
C750 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout 0.06446f
C751 XThC.Tn[12] XA.XIR[0].XIC[12].icell.Ien 0.03728f
C752 XA.XIR[12].XIC[10].icell.PUM VPWR 0.01015f
C753 XA.XIR[13].XIC[4].icell.Ien Iout 0.06821f
C754 XThC.Tn[13] XThR.Tn[4] 0.29363f
C755 XThC.Tn[11] XA.XIR[15].XIC[11].icell.Ien 0.03184f
C756 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.Ien 0.04854f
C757 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.PDM 0.02104f
C758 XThC.XTB4.Y XThC.Tn[11] 0.30582f
C759 XThC.Tn[6] XA.XIR[1].XIC[6].icell.Ien 0.03605f
C760 XA.XIR[15].XIC_dummy_right.icell.Iout Iout 0.01732f
C761 XThC.Tn[8] XThR.Tn[10] 0.29362f
C762 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.01728f
C763 XA.XIR[11].XIC[7].icell.Ien Iout 0.06821f
C764 XA.XIR[9].XIC[1].icell.PUM VPWR 0.01015f
C765 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.Ien 0.04854f
C766 XThC.Tn[0] XThR.Tn[5] 0.29369f
C767 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PDM 0.04035f
C768 XThC.Tn[7] XThR.Tn[0] 0.29461f
C769 XA.XIR[4].XIC[1].icell.Ien Vbias 0.19161f
C770 XA.XIR[10].XIC[9].icell.Ien Iout 0.06821f
C771 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.Ien 0.04854f
C772 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.Ien 0.04854f
C773 XThC.Tn[8] XThC.Tn[9] 0.05322f
C774 XA.XIR[3].XIC[0].icell.PUM VPWR 0.01015f
C775 XThC.XTB7.A a_6243_9615# 0.02018f
C776 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR 0.35722f
C777 XThC.Tn[12] XThC.Tn[14] 0.03994f
C778 XThC.Tn[14] XA.XIR[4].XIC[14].icell.Ien 0.03605f
C779 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PDM 0.04035f
C780 XA.XIR[2].XIC_15.icell.Ien VPWR 0.26829f
C781 XA.XIR[12].XIC[11].icell.Ien VPWR 0.1979f
C782 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.Ien 0.04854f
C783 XThC.XTB1.Y Vbias 0.01234f
C784 XA.XIR[2].XIC[11].icell.Ien Iout 0.06821f
C785 XA.XIR[15].XIC[3].icell.Ien Vbias 0.15966f
C786 XThR.Tn[8] XA.XIR[8].XIC[12].icell.Ien 0.15202f
C787 XThC.Tn[4] XA.XIR[13].XIC[4].icell.Ien 0.03605f
C788 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PDM 0.02765f
C789 XA.XIR[1].XIC[13].icell.Ien Iout 0.06821f
C790 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.Ien 0.04854f
C791 XA.XIR[4].XIC[6].icell.Ien Vbias 0.19161f
C792 XA.XIR[15].XIC[14].icell.PUM VPWR 0.01015f
C793 XThC.Tn[3] XA.XIR[8].XIC[3].icell.Ien 0.03605f
C794 Vbias bias[2] 0.06133f
C795 XThR.XTBN.Y a_n1049_6405# 0.07602f
C796 XThR.Tn[12] a_n997_1803# 0.18719f
C797 XA.XIR[12].XIC[0].icell.Ien Iout 0.06814f
C798 XThR.Tn[5] XA.XIR[5].XIC[11].icell.Ien 0.15202f
C799 XA.XIR[9].XIC[13].icell.PDM Vbias 0.03922f
C800 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PDM 0.02765f
C801 XThC.Tn[6] XThR.Tn[2] 0.29362f
C802 XA.XIR[7].XIC[0].icell.Ien Vbias 0.19149f
C803 XA.XIR[0].XIC[5].icell.PDM Vbias 0.03936f
C804 XA.XIR[15].XIC[5].icell.PUM VPWR 0.01015f
C805 XThR.Tn[11] Iout 1.19575f
C806 XA.XIR[5].XIC[5].icell.Ien VPWR 0.1979f
C807 XA.XIR[2].XIC_dummy_right.icell.Iout VPWR 0.11567f
C808 XA.XIR[9].XIC[9].icell.Ien Vbias 0.19161f
C809 XA.XIR[4].XIC[8].icell.PUM VPWR 0.01015f
C810 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.Ien 0.04854f
C811 XA.XIR[0].XIC[2].icell.Ien Vbias 0.19209f
C812 XA.XIR[11].XIC[14].icell.PDM Vbias 0.03922f
C813 XThC.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.03605f
C814 XThR.XTB4.Y a_n1049_6405# 0.01546f
C815 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PDM 0.02765f
C816 XThR.Tn[5] VPWR 8.25724f
C817 XThC.Tn[12] XA.XIR[3].XIC[12].icell.Ien 0.03605f
C818 XThR.Tn[2] XA.XIR[2].XIC[0].icell.Ien 0.1525f
C819 XA.XIR[0].XIC[9].icell.PDM VPWR 0.01287f
C820 XA.XIR[7].XIC[2].icell.PUM VPWR 0.01015f
C821 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.PDM 0.02104f
C822 XA.XIR[14].XIC_15.icell.PDM Vbias 0.03927f
C823 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.Ien 0.04854f
C824 XA.XIR[14].XIC_15.icell.Ien Vbias 0.19195f
C825 XA.XIR[7].XIC[5].icell.Ien Vbias 0.19161f
C826 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.PDM 0.02104f
C827 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PDM 0.02765f
C828 XThC.Tn[7] XA.XIR[12].XIC[7].icell.Ien 0.03605f
C829 XThC.Tn[2] XThR.Tn[6] 0.29362f
C830 XA.XIR[9].XIC[11].icell.PUM VPWR 0.01015f
C831 XThR.Tn[12] XThR.Tn[13] 0.09917f
C832 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.Ien 0.04854f
C833 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.Ien 0.04854f
C834 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PDM 0.04035f
C835 XThC.Tn[4] XThR.Tn[11] 0.29362f
C836 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PDM 0.04035f
C837 XA.XIR[6].XIC[13].icell.Ien Iout 0.06821f
C838 XA.XIR[7].XIC[7].icell.PUM VPWR 0.01015f
C839 XA.XIR[10].XIC[14].icell.Ien Iout 0.06821f
C840 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.02765f
C841 XThC.XTB5.Y XThC.Tn[5] 0.01095f
C842 XA.XIR[15].XIC[12].icell.PUM VPWR 0.01015f
C843 a_10915_9569# XThC.Tn[14] 0.20278f
C844 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR 0.38999f
C845 XThC.Tn[8] XThR.Tn[13] 0.29362f
C846 XA.XIR[14].XIC[7].icell.Ien Iout 0.06821f
C847 XThR.Tn[14] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0404f
C848 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Iout 0.04498f
C849 XA.XIR[5].XIC[3].icell.PDM Vbias 0.03922f
C850 XThR.Tn[3] XA.XIR[3].XIC[4].icell.Ien 0.15202f
C851 XA.XIR[13].XIC[9].icell.Ien Iout 0.06821f
C852 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.Ien 0.04854f
C853 XThC.Tn[7] XThR.Tn[1] 0.294f
C854 XThC.Tn[11] XThR.Tn[9] 0.29362f
C855 XThC.Tn[11] Iout 0.84391f
C856 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout 0.06446f
C857 XThC.XTB2.Y data[1] 0.017f
C858 XThC.Tn[7] XThR.Tn[12] 0.29362f
C859 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PDM 0.02765f
C860 XA.XIR[12].XIC[2].icell.PDM Vbias 0.03922f
C861 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PDM 0.02765f
C862 a_5155_9615# VPWR 0.7051f
C863 XA.XIR[11].XIC[8].icell.PDM Vbias 0.03922f
C864 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PDM 0.04056f
C865 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PDM 0.02765f
C866 XThC.XTBN.Y XThC.Tn[5] 0.60785f
C867 XThC.Tn[2] XThR.Tn[4] 0.29362f
C868 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PDM 0.04035f
C869 XA.XIR[15].XIC[13].icell.Ien VPWR 0.33655f
C870 XA.XIR[3].XIC[2].icell.Ien Vbias 0.19161f
C871 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.Ien 0.04854f
C872 XThC.Tn[13] XA.XIR[5].XIC[13].icell.Ien 0.03605f
C873 XThC.Tn[6] XThR.Tn[10] 0.29362f
C874 XThR.XTB7.B XThR.XTB7.A 0.35833f
C875 XThR.XTB5.A XThR.XTB3.Y 0.01152f
C876 XThC.XTBN.A data[3] 0.07741f
C877 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PDM 0.02765f
C878 XA.XIR[15].XIC[8].icell.Ien Vbias 0.15966f
C879 XThC.XTB7.A data[0] 0.86893f
C880 XA.XIR[5].XIC[1].icell.Ien Iout 0.06821f
C881 XThC.Tn[7] XThC.Tn[8] 0.07597f
C882 XA.XIR[4].XIC[11].icell.Ien Vbias 0.19161f
C883 XA.XIR[8].XIC[0].icell.PDM Vbias 0.03915f
C884 XThR.Tn[14] Iout 1.19574f
C885 XThC.Tn[9] XA.XIR[7].XIC[9].icell.Ien 0.03605f
C886 XA.XIR[11].XIC[13].icell.PDM Vbias 0.03922f
C887 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout 0.06446f
C888 XA.XIR[2].XIC[4].icell.PDM Vbias 0.03922f
C889 XA.XIR[8].XIC[2].icell.PUM VPWR 0.01015f
C890 XA.XIR[8].XIC[5].icell.Ien Vbias 0.19161f
C891 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PDM 0.04035f
C892 XA.XIR[3].XIC[4].icell.PUM VPWR 0.01015f
C893 XA.XIR[10].XIC[12].icell.Ien Iout 0.06821f
C894 XThC.XTB6.Y VPWR 1.03148f
C895 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.Ien 0.04854f
C896 XA.XIR[14].XIC[14].icell.PDM Vbias 0.03922f
C897 XA.XIR[11].XIC_dummy_left.icell.Iout VPWR 0.1106f
C898 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.PDM 0.02104f
C899 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.02765f
C900 XA.XIR[15].XIC[10].icell.PUM VPWR 0.01015f
C901 XA.XIR[5].XIC[10].icell.Ien VPWR 0.1979f
C902 XThC.XTBN.Y a_10051_9569# 0.23006f
C903 XA.XIR[9].XIC[14].icell.Ien Vbias 0.19161f
C904 XThR.XTB7.A XThR.Tn[2] 0.12549f
C905 XThR.XTB5.Y XThR.Tn[8] 0.01728f
C906 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.Ien 0.04854f
C907 XThR.Tn[4] XA.XIR[4].XIC[1].icell.Ien 0.15202f
C908 XA.XIR[5].XIC[6].icell.Ien Iout 0.06821f
C909 XA.XIR[4].XIC[13].icell.PUM VPWR 0.01015f
C910 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PDM 0.02765f
C911 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10] 0.15202f
C912 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PDM 0.02765f
C913 XThR.Tn[3] XA.XIR[3].XIC[1].icell.Ien 0.15202f
C914 XA.XIR[0].XIC[7].icell.Ien Vbias 0.19212f
C915 XA.XIR[8].XIC[7].icell.PUM VPWR 0.01015f
C916 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PDM 0.02765f
C917 XA.XIR[12].XIC[5].icell.Ien VPWR 0.1979f
C918 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.Ien 0.04854f
C919 XThC.Tn[11] XA.XIR[9].XIC[11].icell.Ien 0.03605f
C920 XThC.Tn[4] XThR.Tn[14] 0.29362f
C921 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.Ien 0.04854f
C922 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PDM 0.04035f
C923 XA.XIR[7].XIC[10].icell.Ien Vbias 0.19161f
C924 XA.XIR[2].XIC_dummy_left.icell.Iout Iout 0.0353f
C925 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PDM 0.02765f
C926 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR 0.01691f
C927 XA.XIR[15].XIC[11].icell.Ien VPWR 0.33655f
C928 XThR.Tn[4] XA.XIR[4].XIC[6].icell.Ien 0.15202f
C929 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PDM 0.02765f
C930 XA.XIR[13].XIC[14].icell.Ien Iout 0.06821f
C931 XThC.XTB4.Y VPWR 0.91479f
C932 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.Ien 0.04854f
C933 XThC.Tn[12] XA.XIR[1].XIC[12].icell.Ien 0.03611f
C934 XA.XIR[8].XIC[0].icell.Ien Vbias 0.19149f
C935 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PDM 0.04035f
C936 XThC.XTB3.Y XThC.XTBN.A 0.03907f
C937 XA.XIR[8].XIC_dummy_left.icell.Iout XA.XIR[9].XIC_dummy_left.icell.Iout 0.03665f
C938 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PDM 0.04035f
C939 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout 0.06446f
C940 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Iout 0.04591f
C941 XThR.XTB5.A VPWR 0.83125f
C942 XThC.XTB5.A data[0] 0.14415f
C943 XA.XIR[7].XIC[12].icell.PUM VPWR 0.01015f
C944 XA.XIR[7].XIC[4].icell.PDM Vbias 0.03922f
C945 XThR.XTB1.Y XThR.Tn[8] 0.29191f
C946 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PDM 0.04035f
C947 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PDM 0.0404f
C948 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR 0.08221f
C949 XA.XIR[15].XIC[2].icell.PDM Vbias 0.03922f
C950 XA.XIR[6].XIC[11].icell.PDM Vbias 0.03922f
C951 XA.XIR[10].XIC[10].icell.Ien Iout 0.06821f
C952 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.PDM 0.02104f
C953 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PDM 0.02765f
C954 XThR.Tn[12] XA.XIR[12].XIC[4].icell.Ien 0.15202f
C955 XA.XIR[3].XIC[1].icell.PUM VPWR 0.01015f
C956 XA.XIR[14].XIC[8].icell.PDM Vbias 0.03922f
C957 XThR.Tn[3] XA.XIR[3].XIC[9].icell.Ien 0.15202f
C958 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PDM 0.02765f
C959 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PDM 0.02765f
C960 XThR.XTBN.Y XThR.XTB7.A 0.59539f
C961 XA.XIR[11].XIC[2].icell.PUM VPWR 0.01015f
C962 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.Ien 0.04854f
C963 XA.XIR[9].XIC[0].icell.PDM Vbias 0.03915f
C964 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PDM 0.04035f
C965 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR 0.35722f
C966 XThC.Tn[9] XA.XIR[8].XIC[9].icell.Ien 0.03605f
C967 XA.XIR[9].XIC[1].icell.Ien VPWR 0.1979f
C968 XThR.Tn[2] XA.XIR[2].XIC[4].icell.Ien 0.15202f
C969 XThC.Tn[6] XThR.Tn[13] 0.29362f
C970 VPWR data[5] 0.4402f
C971 XA.XIR[4].XIC[3].icell.Ien VPWR 0.1979f
C972 XA.XIR[15].XIC[6].icell.PDM VPWR 0.01334f
C973 XA.XIR[6].XIC_15.icell.PDM VPWR 0.07527f
C974 XThC.Tn[7] XA.XIR[15].XIC[7].icell.Ien 0.03184f
C975 XThC.Tn[0] Iout 0.82184f
C976 XA.XIR[11].XIC[12].icell.PDM Vbias 0.03922f
C977 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout 0.06446f
C978 XThC.Tn[0] XThR.Tn[9] 0.29367f
C979 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.PDM 0.02104f
C980 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.Ien 0.04854f
C981 XA.XIR[1].XIC[5].icell.PDM Vbias 0.03922f
C982 XThC.Tn[5] XThR.Tn[8] 0.29362f
C983 XA.XIR[3].XIC[7].icell.Ien Vbias 0.19161f
C984 XThR.XTB2.Y XThR.XTB5.Y 0.0451f
C985 XThR.XTB7.A XThR.XTB4.Y 0.14536f
C986 XA.XIR[14].XIC[13].icell.PDM Vbias 0.03922f
C987 XA.XIR[13].XIC[12].icell.Ien Iout 0.06821f
C988 XThC.Tn[12] XA.XIR[6].XIC[12].icell.Ien 0.03605f
C989 XThC.Tn[3] XA.XIR[2].XIC[3].icell.Ien 0.03605f
C990 XA.XIR[4].XIC[5].icell.PDM Vbias 0.03922f
C991 XThC.XTB2.Y VPWR 0.97668f
C992 XThC.XTB5.Y XThC.XTB7.Y 0.036f
C993 XThC.XTB7.B XThC.XTB6.Y 0.30244f
C994 XA.XIR[14].XIC_dummy_left.icell.Iout VPWR 0.1106f
C995 XA.XIR[9].XIC[6].icell.Ien VPWR 0.1979f
C996 XA.XIR[1].XIC[2].icell.Ien Vbias 0.19173f
C997 XA.XIR[8].XIC_15.icell.PDM Vbias 0.03927f
C998 XA.XIR[3].XIC[13].icell.PDM Vbias 0.03922f
C999 XThC.Tn[0] XA.XIR[15].XIC[0].icell.Ien 0.03184f
C1000 XA.XIR[9].XIC[2].icell.Ien Iout 0.06821f
C1001 XThR.Tn[9] XA.XIR[9].XIC[2].icell.Ien 0.15202f
C1002 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.Ien 0.04854f
C1003 XThC.XTB1.Y XThC.XTBN.A 0.12307f
C1004 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PDM 0.04035f
C1005 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PDM 0.02765f
C1006 XA.XIR[8].XIC[10].icell.Ien Vbias 0.19161f
C1007 XA.XIR[3].XIC[9].icell.PUM VPWR 0.01015f
C1008 XThC.XTB3.Y XThC.Tn[2] 0.1864f
C1009 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PDM 0.02855f
C1010 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.Ien 0.04854f
C1011 XThC.Tn[1] XThC.Tn[3] 0.10977f
C1012 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PDM 0.02765f
C1013 XA.XIR[7].XIC[2].icell.Ien VPWR 0.1979f
C1014 XA.XIR[5].XIC_15.icell.Ien VPWR 0.26829f
C1015 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PDM 0.04035f
C1016 XThC.Tn[6] XThC.Tn[7] 0.16021f
C1017 XA.XIR[1].XIC[4].icell.PUM VPWR 0.01015f
C1018 XA.XIR[5].XIC[11].icell.Ien Iout 0.06821f
C1019 XThC.XTB7.Y XThC.XTBN.Y 0.50018f
C1020 XA.XIR[12].XIC_15.icell.PDM VPWR 0.07527f
C1021 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.Ien 0.04854f
C1022 XA.XIR[0].XIC[12].icell.Ien Vbias 0.19209f
C1023 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1024 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PDM 0.02765f
C1025 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.04035f
C1026 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.PDM 0.02104f
C1027 XA.XIR[8].XIC[12].icell.PUM VPWR 0.01015f
C1028 XThC.XTB4.Y XThC.XTB7.B 0.33064f
C1029 XThC.Tn[8] XThR.Tn[7] 0.29362f
C1030 XThR.XTB1.Y XThR.XTB2.Y 2.14864f
C1031 XA.XIR[12].XIC[6].icell.Ien Iout 0.06821f
C1032 XA.XIR[7].XIC_15.icell.Ien Vbias 0.19195f
C1033 XA.XIR[10].XIC_15.icell.Ien Iout 0.0694f
C1034 XThC.XTB7.Y XThC.Tn[10] 0.07406f
C1035 VPWR Iout 56.251f
C1036 XA.XIR[5].XIC[0].icell.Ien Vbias 0.19149f
C1037 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PDM 0.04035f
C1038 XThR.Tn[9] VPWR 9.19311f
C1039 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.PDM 0.02104f
C1040 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.04035f
C1041 XThR.Tn[4] XA.XIR[4].XIC[11].icell.Ien 0.15202f
C1042 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.PDM 0.02104f
C1043 XA.XIR[5].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1044 XThC.Tn[14] Vbias 1.14968f
C1045 XThR.Tn[10] XA.XIR[10].XIC[2].icell.Ien 0.15202f
C1046 XThR.Tn[0] XA.XIR[0].XIC[3].icell.Ien 0.15202f
C1047 XA.XIR[12].XIC[0].icell.PUM VPWR 0.01015f
C1048 XThR.XTB7.B XThR.XTBN.Y 0.3875f
C1049 XA.XIR[13].XIC[10].icell.Ien Iout 0.06821f
C1050 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PDM 0.04035f
C1051 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.04056f
C1052 XA.XIR[6].XIC[2].icell.Ien Vbias 0.19161f
C1053 XThR.Tn[7] XA.XIR[7].XIC[4].icell.Ien 0.15202f
C1054 XA.XIR[15].XIC[0].icell.Ien VPWR 0.33655f
C1055 XThC.Tn[11] XA.XIR[10].XIC[11].icell.Ien 0.03605f
C1056 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.PDM 0.02104f
C1057 XA.XIR[14].XIC[2].icell.PUM VPWR 0.01015f
C1058 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.Ien 0.04854f
C1059 XThC.XTB1.Y XThC.XTB3.Y 0.04033f
C1060 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PDM 0.02765f
C1061 XA.XIR[10].XIC_dummy_right.icell.Iout Iout 0.01732f
C1062 XA.XIR[11].XIC[11].icell.PDM Vbias 0.03922f
C1063 XThR.Tn[12] XA.XIR[12].XIC[9].icell.Ien 0.15202f
C1064 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.PDM 0.02104f
C1065 XThC.Tn[4] VPWR 6.44479f
C1066 XThR.Tn[3] XA.XIR[3].XIC[14].icell.Ien 0.15202f
C1067 XThR.XTB7.B XThR.XTB4.Y 0.33064f
C1068 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.Ien 0.04854f
C1069 XA.XIR[14].XIC[12].icell.PDM Vbias 0.03922f
C1070 XA.XIR[6].XIC[4].icell.PUM VPWR 0.01015f
C1071 XA.XIR[9].XIC_15.icell.PDM Vbias 0.03927f
C1072 XThC.Tn[10] XThR.Tn[0] 0.2938f
C1073 XThR.XTBN.Y XThR.Tn[2] 0.6189f
C1074 XA.XIR[15].XIC[5].icell.Ien VPWR 0.33655f
C1075 XA.XIR[0].XIC[7].icell.PDM Vbias 0.03939f
C1076 XThC.Tn[12] XThR.Tn[5] 0.29362f
C1077 XThR.XTB7.B XThR.Tn[10] 0.06102f
C1078 XThC.XTB7.B a_7875_9569# 0.01174f
C1079 XThR.Tn[2] XA.XIR[2].XIC[9].icell.Ien 0.15202f
C1080 XA.XIR[10].XIC[3].icell.Ien Vbias 0.19161f
C1081 XA.XIR[4].XIC[8].icell.Ien VPWR 0.1979f
C1082 XThC.XTB6.A XThC.XTB5.Y 0.01866f
C1083 XThC.XTB2.Y XThC.XTB7.B 0.22599f
C1084 XA.XIR[4].XIC[4].icell.Ien Iout 0.06821f
C1085 a_8963_9569# XThC.Tn[11] 0.19413f
C1086 XA.XIR[8].XIC[2].icell.Ien VPWR 0.1979f
C1087 XA.XIR[3].XIC[12].icell.Ien Vbias 0.19161f
C1088 XA.XIR[10].XIC[14].icell.PUM VPWR 0.01015f
C1089 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.Ien 0.04854f
C1090 XA.XIR[2].XIC[2].icell.PUM VPWR 0.01015f
C1091 XThC.Tn[2] XA.XIR[0].XIC[2].icell.Ien 0.03784f
C1092 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13] 0.15202f
C1093 XA.XIR[11].XIC[3].icell.PUM VPWR 0.01015f
C1094 XA.XIR[2].XIC[5].icell.Ien Vbias 0.19161f
C1095 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.Ien 0.04854f
C1096 XA.XIR[9].XIC[11].icell.Ien VPWR 0.1979f
C1097 XA.XIR[1].XIC[7].icell.Ien Vbias 0.19173f
C1098 XA.XIR[10].XIC[5].icell.PUM VPWR 0.01015f
C1099 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.PDM 0.02104f
C1100 XA.XIR[12].XIC[14].icell.PDM VPWR 0.01002f
C1101 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.PDM 0.02104f
C1102 XA.XIR[9].XIC[7].icell.Ien Iout 0.06821f
C1103 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PDM 0.02765f
C1104 XThR.Tn[9] XA.XIR[9].XIC[7].icell.Ien 0.15202f
C1105 XThC.XTB6.A XThC.XTBN.Y 0.03867f
C1106 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PDM 0.04035f
C1107 XA.XIR[0].XIC[4].icell.Ien VPWR 0.19742f
C1108 XA.XIR[8].XIC_15.icell.Ien Vbias 0.19195f
C1109 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PDM 0.04035f
C1110 XA.XIR[3].XIC[14].icell.PUM VPWR 0.01015f
C1111 XThC.Tn[9] XThR.Tn[2] 0.29362f
C1112 XA.XIR[15].XIC_15.icell.PDM VPWR 0.07867f
C1113 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PDM 0.02765f
C1114 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.PDM 0.02104f
C1115 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.Ien 0.04854f
C1116 XA.XIR[2].XIC[7].icell.PUM VPWR 0.01015f
C1117 XThC.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.03605f
C1118 XA.XIR[7].XIC[7].icell.Ien VPWR 0.1979f
C1119 XThR.XTB5.Y XThR.XTB7.Y 0.036f
C1120 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.04035f
C1121 XA.XIR[7].XIC_dummy_left.icell.Ien XThR.Tn[7] 0.01444f
C1122 XA.XIR[1].XIC[9].icell.PUM VPWR 0.01015f
C1123 XA.XIR[7].XIC[3].icell.Ien Iout 0.06821f
C1124 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.PDM 0.02104f
C1125 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.Ien 0.04854f
C1126 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PDM 0.02765f
C1127 XA.XIR[13].XIC_15.icell.Ien Iout 0.0694f
C1128 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.Ien 0.04854f
C1129 XThC.XTB7.A XThC.Tn[5] 0.02758f
C1130 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR 0.38922f
C1131 XA.XIR[5].XIC[5].icell.PDM Vbias 0.03922f
C1132 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.PDM 0.02104f
C1133 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PDM 0.0404f
C1134 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.Ien 0.04854f
C1135 data[1] data[0] 0.64735f
C1136 XThC.Tn[14] XA.XIR[11].XIC[14].icell.Ien 0.03605f
C1137 XThR.Tn[11] XA.XIR[11].XIC[3].icell.Ien 0.15202f
C1138 XThC.Tn[14] XThR.Tn[6] 0.29368f
C1139 XA.XIR[12].XIC[4].icell.PDM Vbias 0.03922f
C1140 XThR.Tn[12] XA.XIR[12].XIC[14].icell.Ien 0.15202f
C1141 XA.XIR[11].XIC[10].icell.PDM Vbias 0.03922f
C1142 a_6243_9615# VPWR 0.70553f
C1143 XThR.Tn[0] XA.XIR[0].XIC[8].icell.Ien 0.15202f
C1144 XThC.Tn[11] XA.XIR[13].XIC[11].icell.Ien 0.03605f
C1145 XThR.Tn[10] XA.XIR[10].XIC[7].icell.Ien 0.15202f
C1146 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PDM 0.04035f
C1147 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.Ien 0.04854f
C1148 XA.XIR[10].XIC[12].icell.PUM VPWR 0.01015f
C1149 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.Ien 0.04854f
C1150 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PDM 0.02765f
C1151 XThR.XTBN.Y XThR.XTB4.Y 0.15627f
C1152 XThR.Tn[6] XA.XIR[6].XIC[2].icell.Ien 0.15202f
C1153 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.02765f
C1154 XA.XIR[13].XIC_dummy_right.icell.Iout Iout 0.01732f
C1155 XThC.Tn[6] XThR.Tn[7] 0.29362f
C1156 XA.XIR[14].XIC[11].icell.PDM Vbias 0.03922f
C1157 XA.XIR[11].XIC_dummy_left.icell.Iout XA.XIR[12].XIC_dummy_left.icell.Iout 0.03665f
C1158 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PDM 0.02844f
C1159 XThR.Tn[7] XA.XIR[7].XIC[9].icell.Ien 0.15202f
C1160 XA.XIR[6].XIC[7].icell.Ien Vbias 0.19161f
C1161 XThR.XTBN.Y XThR.Tn[10] 0.46535f
C1162 XThC.XTB5.Y XThC.Tn[8] 0.01728f
C1163 XThR.XTB1.Y data[4] 0.06453f
C1164 XThR.XTB1.Y XThR.XTB7.Y 0.05211f
C1165 XThC.Tn[3] Vbias 1.14954f
C1166 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PDM 0.02765f
C1167 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.Ien 0.04854f
C1168 XThC.XTB6.Y XThC.Tn[12] 0.02863f
C1169 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.Ien 0.04854f
C1170 XA.XIR[15].XIC[1].icell.Ien Iout 0.07211f
C1171 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.Ien 0.04854f
C1172 XA.XIR[5].XIC_dummy_left.icell.Iout Iout 0.0353f
C1173 XThC.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.03605f
C1174 XA.XIR[3].XIC[0].icell.PDM Vbias 0.03915f
C1175 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.Ien 0.04854f
C1176 XA.XIR[8].XIC[2].icell.PDM Vbias 0.03922f
C1177 XThC.Tn[10] XThR.Tn[1] 0.29362f
C1178 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PDM 0.02765f
C1179 XThC.Tn[9] XA.XIR[2].XIC[9].icell.Ien 0.03605f
C1180 XA.XIR[2].XIC[6].icell.PDM Vbias 0.03922f
C1181 a_5949_9615# XThC.Tn[5] 0.27124f
C1182 XA.XIR[13].XIC[3].icell.Ien Vbias 0.19161f
C1183 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PDM 0.04035f
C1184 XA.XIR[10].XIC[13].icell.Ien VPWR 0.1979f
C1185 XA.XIR[3].XIC[4].icell.Ien VPWR 0.1979f
C1186 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1187 XThC.Tn[10] XThR.Tn[12] 0.29362f
C1188 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.02765f
C1189 XA.XIR[6].XIC[9].icell.PUM VPWR 0.01015f
C1190 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.PDM 0.02104f
C1191 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.Ien 0.04854f
C1192 XThR.XTB4.Y XThR.Tn[10] 0.01391f
C1193 XA.XIR[11].XIC[6].icell.Ien Vbias 0.19161f
C1194 XA.XIR[13].XIC[14].icell.PUM VPWR 0.01015f
C1195 XThR.Tn[2] XA.XIR[2].XIC[14].icell.Ien 0.15202f
C1196 XThC.Tn[5] XThR.Tn[3] 0.29362f
C1197 XThC.XTBN.Y XThC.Tn[8] 0.50311f
C1198 XA.XIR[15].XIC[6].icell.Ien Iout 0.07211f
C1199 XA.XIR[6].XIC_dummy_right.icell.Iout XA.XIR[7].XIC_dummy_right.icell.Iout 0.04047f
C1200 XA.XIR[10].XIC[8].icell.Ien Vbias 0.19161f
C1201 XA.XIR[4].XIC[13].icell.Ien VPWR 0.1979f
C1202 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.PDM 0.02104f
C1203 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Iout 0.04563f
C1204 XThC.XTB1.Y a_2979_9615# 0.21263f
C1205 XA.XIR[14].XIC[3].icell.PUM VPWR 0.01015f
C1206 XThC.Tn[14] XThR.Tn[4] 0.29368f
C1207 XA.XIR[4].XIC[9].icell.Ien Iout 0.06821f
C1208 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Iout 0.04498f
C1209 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.PDM 0.02104f
C1210 XA.XIR[13].XIC[5].icell.PUM VPWR 0.01015f
C1211 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PDM 0.02765f
C1212 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PDM 0.04041f
C1213 XA.XIR[0].XIC[0].icell.Ien Iout 0.06768f
C1214 XThR.XTB5.Y XThR.Tn[11] 0.02067f
C1215 XA.XIR[15].XIC[14].icell.PDM VPWR 0.01343f
C1216 XA.XIR[8].XIC[7].icell.Ien VPWR 0.1979f
C1217 XThC.Tn[9] XThR.Tn[10] 0.29362f
C1218 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.PDM 0.02104f
C1219 XThC.Tn[1] XThR.Tn[5] 0.29362f
C1220 XA.XIR[8].XIC[3].icell.Ien Iout 0.06821f
C1221 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PDM 0.02765f
C1222 XThR.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.15202f
C1223 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.Ien 0.04854f
C1224 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PDM 0.02765f
C1225 XA.XIR[11].XIC[8].icell.PUM VPWR 0.01015f
C1226 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.Ien 0.04854f
C1227 XA.XIR[2].XIC[10].icell.Ien Vbias 0.19161f
C1228 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PDM 0.04035f
C1229 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1230 XThC.Tn[13] XThC.Tn[14] 0.38789f
C1231 XA.XIR[10].XIC[10].icell.PUM VPWR 0.01015f
C1232 XA.XIR[1].XIC[12].icell.Ien Vbias 0.19173f
C1233 XA.XIR[9].XIC[12].icell.Ien Iout 0.06821f
C1234 XThR.Tn[9] XA.XIR[9].XIC[12].icell.Ien 0.15202f
C1235 XA.XIR[0].XIC[9].icell.Ien VPWR 0.19875f
C1236 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1237 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PDM 0.02765f
C1238 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.PDM 0.02104f
C1239 XA.XIR[0].XIC[5].icell.Ien Iout 0.06775f
C1240 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PDM 0.04035f
C1241 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PDM 0.04035f
C1242 XThR.XTBN.Y a_n997_1803# 0.22873f
C1243 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PDM 0.04035f
C1244 XA.XIR[2].XIC[12].icell.PUM VPWR 0.01015f
C1245 XA.XIR[7].XIC[12].icell.Ien VPWR 0.1979f
C1246 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.PDM 0.02104f
C1247 XThR.Tn[13] XA.XIR[13].XIC[2].icell.Ien 0.15202f
C1248 XA.XIR[7].XIC[8].icell.Ien Iout 0.06821f
C1249 XA.XIR[1].XIC[14].icell.PUM VPWR 0.01015f
C1250 XThC.Tn[3] XA.XIR[5].XIC[3].icell.Ien 0.03605f
C1251 XA.XIR[7].XIC[6].icell.PDM Vbias 0.03922f
C1252 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PDM 0.04035f
C1253 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.Ien 0.04854f
C1254 XThC.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.03605f
C1255 XA.XIR[15].XIC[4].icell.PDM Vbias 0.03922f
C1256 XThR.XTB6.A XThR.XTB2.Y 0.18237f
C1257 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.Ien 0.04854f
C1258 XA.XIR[10].XIC[11].icell.Ien VPWR 0.1979f
C1259 XA.XIR[6].XIC[13].icell.PDM Vbias 0.03922f
C1260 XA.XIR[3].XIC[1].icell.Ien VPWR 0.1979f
C1261 XThC.Tn[7] XThR.Tn[2] 0.29372f
C1262 XThC.XTB7.B a_6243_9615# 0.01743f
C1263 XA.XIR[14].XIC[10].icell.PDM Vbias 0.03922f
C1264 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PDM 0.02765f
C1265 XA.XIR[12].XIC[1].icell.PUM VPWR 0.01015f
C1266 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.PDM 0.02104f
C1267 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout 0.06446f
C1268 XA.XIR[13].XIC[12].icell.PUM VPWR 0.01015f
C1269 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PDM 0.02765f
C1270 XThR.Tn[11] XA.XIR[11].XIC[8].icell.Ien 0.15202f
C1271 XA.XIR[9].XIC[2].icell.PDM Vbias 0.03922f
C1272 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PDM 0.0404f
C1273 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PDM 0.02802f
C1274 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.PDM 0.02104f
C1275 XA.XIR[9].XIC_dummy_left.icell.Iout VPWR 0.1106f
C1276 XThR.XTBN.Y XThR.Tn[13] 0.56841f
C1277 XA.XIR[12].XIC[13].icell.Ien Vbias 0.19161f
C1278 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PDM 0.02765f
C1279 XA.XIR[15].XIC[8].icell.PDM VPWR 0.01334f
C1280 XA.XIR[10].XIC[0].icell.Ien Iout 0.06814f
C1281 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.PDM 0.02104f
C1282 XThR.Tn[0] XA.XIR[0].XIC[13].icell.Ien 0.15202f
C1283 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.PDM 0.02104f
C1284 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.Ien 0.04854f
C1285 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.PDM 0.02104f
C1286 XThR.Tn[6] XA.XIR[6].XIC[7].icell.Ien 0.15202f
C1287 XThR.Tn[12] XA.XIR[12].XIC[10].icell.Ien 0.15202f
C1288 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.PDM 0.02104f
C1289 XA.XIR[0].XIC_dummy_left.icell.Iout XA.XIR[1].XIC_dummy_left.icell.Iout 0.03665f
C1290 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.PDM 0.02104f
C1291 XThC.Tn[3] XThR.Tn[6] 0.29362f
C1292 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PDM 0.02765f
C1293 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.PDM 0.02104f
C1294 XA.XIR[1].XIC[7].icell.PDM Vbias 0.03922f
C1295 XThR.Tn[7] XA.XIR[7].XIC[14].icell.Ien 0.15202f
C1296 XA.XIR[6].XIC[12].icell.Ien Vbias 0.19161f
C1297 VPWR data[0] 0.52929f
C1298 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.Ien 0.04854f
C1299 XA.XIR[13].XIC[13].icell.Ien VPWR 0.1979f
C1300 XA.XIR[4].XIC[7].icell.PDM Vbias 0.03922f
C1301 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PDM 0.02765f
C1302 XThC.Tn[5] XThR.Tn[11] 0.29362f
C1303 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.Ien 0.04854f
C1304 XA.XIR[3].XIC_15.icell.PDM Vbias 0.03927f
C1305 XThC.XTB7.A XThC.XTB7.Y 0.37429f
C1306 XA.XIR[14].XIC[6].icell.Ien Vbias 0.19161f
C1307 XThC.Tn[8] XA.XIR[0].XIC[8].icell.Ien 0.03758f
C1308 XA.XIR[13].XIC[8].icell.Ien Vbias 0.19161f
C1309 XA.XIR[15].XIC[13].icell.PDM VPWR 0.01334f
C1310 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PDM 0.04035f
C1311 XThC.Tn[7] XA.XIR[10].XIC[7].icell.Ien 0.03605f
C1312 XA.XIR[3].XIC[9].icell.Ien VPWR 0.1979f
C1313 XThC.Tn[2] XA.XIR[1].XIC[2].icell.Ien 0.0362f
C1314 XA.XIR[6].XIC[14].icell.PUM VPWR 0.01015f
C1315 XA.XIR[12].XIC_dummy_left.icell.Iout Iout 0.0353f
C1316 XA.XIR[3].XIC[5].icell.Ien Iout 0.06821f
C1317 XThC.Tn[9] XThR.Tn[13] 0.29362f
C1318 XA.XIR[2].XIC[2].icell.Ien VPWR 0.1979f
C1319 XA.XIR[2].XIC_dummy_right.icell.Iout XA.XIR[3].XIC_dummy_right.icell.Iout 0.04047f
C1320 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PDM 0.04035f
C1321 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.PDM 0.02104f
C1322 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PDM 0.02765f
C1323 XA.XIR[1].XIC[4].icell.Ien VPWR 0.1979f
C1324 XA.XIR[14].XIC[8].icell.PUM VPWR 0.01015f
C1325 XThC.Tn[12] Iout 0.84555f
C1326 XThC.Tn[10] XA.XIR[4].XIC[10].icell.Ien 0.03605f
C1327 XThC.Tn[12] XThR.Tn[9] 0.29362f
C1328 XA.XIR[4].XIC[14].icell.Ien Iout 0.06821f
C1329 XThC.Tn[8] XThR.Tn[8] 0.29362f
C1330 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PDM 0.04035f
C1331 XA.XIR[13].XIC[10].icell.PUM VPWR 0.01015f
C1332 XA.XIR[8].XIC[12].icell.Ien VPWR 0.1979f
C1333 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PDM 0.04035f
C1334 XA.XIR[8].XIC[8].icell.Ien Iout 0.06821f
C1335 XThC.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.03605f
C1336 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.PDM 0.02104f
C1337 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.Ien 0.04854f
C1338 XA.XIR[2].XIC_15.icell.Ien Vbias 0.19195f
C1339 XThC.XTBN.Y XThC.Tn[6] 0.61358f
C1340 XThC.Tn[3] XThR.Tn[4] 0.29362f
C1341 XA.XIR[12].XIC[11].icell.Ien Vbias 0.19161f
C1342 XThR.XTB7.B a_n997_3979# 0.01152f
C1343 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.Ien 0.04854f
C1344 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PDM 0.04035f
C1345 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.Ien 0.04854f
C1346 XA.XIR[0].XIC[14].icell.Ien VPWR 0.19732f
C1347 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.Ien 0.04854f
C1348 XThC.Tn[7] XThR.Tn[10] 0.29362f
C1349 XThR.Tn[1] XA.XIR[1].XIC[3].icell.Ien 0.15202f
C1350 XA.XIR[10].XIC[1].icell.PDM Vbias 0.03922f
C1351 XThR.Tn[14] XA.XIR[14].XIC[3].icell.Ien 0.15202f
C1352 XA.XIR[0].XIC[10].icell.Ien Iout 0.06775f
C1353 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.PDM 0.02104f
C1354 XA.XIR[13].XIC[11].icell.Ien VPWR 0.1979f
C1355 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.04035f
C1356 a_7651_9569# XThC.Tn[8] 0.1927f
C1357 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PDM 0.02765f
C1358 XA.XIR[5].XIC[2].icell.PUM VPWR 0.01015f
C1359 XThR.Tn[13] XA.XIR[13].XIC[7].icell.Ien 0.15202f
C1360 XA.XIR[5].XIC[5].icell.Ien Vbias 0.19161f
C1361 XA.XIR[7].XIC[13].icell.Ien Iout 0.06821f
C1362 XThR.Tn[12] XA.XIR[12].XIC_15.icell.Ien 0.13564f
C1363 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.Ien 0.04854f
C1364 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PDM 0.02765f
C1365 XThC.Tn[2] XA.XIR[6].XIC[2].icell.Ien 0.03605f
C1366 XThR.XTB2.Y XThR.Tn[1] 0.17876f
C1367 XA.XIR[13].XIC[0].icell.Ien Iout 0.06814f
C1368 XThC.Tn[8] XA.XIR[3].XIC[8].icell.Ien 0.03605f
C1369 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PDM 0.02774f
C1370 XThR.Tn[5] Vbias 1.44824f
C1371 XThR.XTB7.B XThR.Tn[7] 0.07415f
C1372 XThC.Tn[3] XA.XIR[12].XIC[3].icell.Ien 0.03605f
C1373 XA.XIR[6].XIC[4].icell.Ien VPWR 0.1979f
C1374 XThR.XTB7.B a_n997_2891# 0.0168f
C1375 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PDM 0.02765f
C1376 XA.XIR[0].XIC[9].icell.PDM Vbias 0.03943f
C1377 XA.XIR[5].XIC[7].icell.PUM VPWR 0.01015f
C1378 XThC.Tn[1] XA.XIR[9].XIC[1].icell.Ien 0.03605f
C1379 XThC.XTB7.B a_8963_9569# 0.02071f
C1380 XThC.XTB7.B data[0] 0.0138f
C1381 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.Ien 0.04854f
C1382 XThC.Tn[5] XThR.Tn[14] 0.29362f
C1383 XThR.Tn[6] XA.XIR[6].XIC[12].icell.Ien 0.15202f
C1384 XA.XIR[15].XIC[12].icell.PDM VPWR 0.01334f
C1385 XThC.XTB6.A XThC.XTB7.A 0.44014f
C1386 XThR.XTB6.A data[4] 0.48493f
C1387 XThR.XTB6.A XThR.XTB7.Y 0.01596f
C1388 XThR.XTB3.Y XThR.XTB5.Y 0.04438f
C1389 XThC.Tn[7] XA.XIR[13].XIC[7].icell.Ien 0.03605f
C1390 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.PDM 0.02104f
C1391 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.Ien 0.04854f
C1392 XA.XIR[11].XIC[3].icell.Ien VPWR 0.1979f
C1393 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.PDM 0.02104f
C1394 XThC.XTB2.Y XThC.Tn[1] 0.17879f
C1395 XA.XIR[10].XIC[5].icell.Ien VPWR 0.1979f
C1396 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout 0.06446f
C1397 XThC.Tn[6] XA.XIR[8].XIC[6].icell.Ien 0.03605f
C1398 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PDM 0.04035f
C1399 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.Ien 0.04854f
C1400 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PDM 0.04035f
C1401 XA.XIR[3].XIC[14].icell.Ien VPWR 0.19796f
C1402 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PDM 0.02765f
C1403 XA.XIR[3].XIC[10].icell.Ien Iout 0.06821f
C1404 XThR.XTBN.Y a_n997_3979# 0.23021f
C1405 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.Ien 0.04854f
C1406 XA.XIR[2].XIC[7].icell.Ien VPWR 0.1979f
C1407 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PDM 0.04056f
C1408 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.PDM 0.02104f
C1409 XA.XIR[2].XIC[3].icell.Ien Iout 0.06821f
C1410 XA.XIR[1].XIC[9].icell.Ien VPWR 0.1979f
C1411 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PDM 0.02765f
C1412 XThR.Tn[8] XA.XIR[8].XIC[4].icell.Ien 0.15202f
C1413 XA.XIR[14].XIC_dummy_left.icell.Iout XA.XIR[15].XIC_dummy_left.icell.Iout 0.03665f
C1414 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PDM 0.02765f
C1415 XA.XIR[1].XIC[5].icell.Ien Iout 0.06821f
C1416 XA.XIR[6].XIC[0].icell.PDM Vbias 0.03915f
C1417 XA.XIR[2].XIC_dummy_left.icell.Iout XA.XIR[3].XIC_dummy_left.icell.Iout 0.03665f
C1418 XA.XIR[15].XIC[13].icell.Ien Vbias 0.15966f
C1419 XA.XIR[1].XIC_dummy_right.icell.Iout XA.XIR[2].XIC_dummy_right.icell.Iout 0.04047f
C1420 XThC.Tn[9] XA.XIR[5].XIC[9].icell.Ien 0.03605f
C1421 XThC.XTB3.Y a_4067_9615# 0.23056f
C1422 XThR.XTB1.Y XThR.XTB3.Y 0.04033f
C1423 XA.XIR[5].XIC[7].icell.PDM Vbias 0.03922f
C1424 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.Ien 0.04854f
C1425 XA.XIR[8].XIC[13].icell.Ien Iout 0.06821f
C1426 a_4067_9615# XThC.Tn[2] 0.27699f
C1427 XThC.Tn[7] XThR.Tn[13] 0.29362f
C1428 XA.XIR[13].XIC[1].icell.PDM Vbias 0.03922f
C1429 XThR.Tn[5] XA.XIR[5].XIC[3].icell.Ien 0.15202f
C1430 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PDM 0.02765f
C1431 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PDM 0.0404f
C1432 XThC.Tn[1] Iout 0.84477f
C1433 XThC.Tn[13] XA.XIR[12].XIC[13].icell.Ien 0.03605f
C1434 XA.XIR[12].XIC[6].icell.PDM Vbias 0.03922f
C1435 XThC.Tn[1] XThR.Tn[9] 0.29362f
C1436 XThC.XTB5.A XThC.XTB6.A 1.80461f
C1437 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout 0.06446f
C1438 XThC.Tn[6] XThR.Tn[8] 0.29362f
C1439 XThR.XTB7.A a_n1049_6699# 0.02294f
C1440 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PDM 0.04056f
C1441 XA.XIR[0].XIC_15.icell.Ien Iout 0.06774f
C1442 XThR.Tn[14] XA.XIR[14].XIC[8].icell.Ien 0.15202f
C1443 XThR.Tn[1] XA.XIR[1].XIC[8].icell.Ien 0.15202f
C1444 XThR.XTB5.Y VPWR 1.0269f
C1445 XThR.XTBN.Y XThR.Tn[7] 0.89996f
C1446 XThR.XTBN.Y a_n997_2891# 0.22804f
C1447 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PDM 0.02765f
C1448 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.Ien 0.04854f
C1449 XThC.XTB6.Y Vbias 0.01503f
C1450 XA.XIR[6].XIC[0].icell.Ien Iout 0.06814f
C1451 XA.XIR[5].XIC[10].icell.Ien Vbias 0.19161f
C1452 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.02765f
C1453 XA.XIR[15].XIC_dummy_left.icell.Iout Iout 0.0353f
C1454 XA.XIR[9].XIC[3].icell.PUM VPWR 0.01015f
C1455 XThC.XTB3.Y XThC.Tn[3] 0.01287f
C1456 XA.XIR[3].XIC[2].icell.PDM Vbias 0.03922f
C1457 XA.XIR[8].XIC[4].icell.PDM Vbias 0.03922f
C1458 XA.XIR[15].XIC[11].icell.PDM VPWR 0.01334f
C1459 XThR.Tn[5] XThR.Tn[6] 0.10245f
C1460 XA.XIR[2].XIC[8].icell.PDM Vbias 0.03922f
C1461 XThC.Tn[2] XThC.Tn[3] 0.33669f
C1462 XThR.XTB4.Y XThR.Tn[7] 0.01797f
C1463 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PDM 0.04035f
C1464 XA.XIR[0].XIC_dummy_right.icell.Iout Iout 0.01732f
C1465 XA.XIR[12].XIC[5].icell.Ien Vbias 0.19161f
C1466 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PDM 0.02765f
C1467 XA.XIR[6].XIC[9].icell.Ien VPWR 0.1979f
C1468 XA.XIR[5].XIC[12].icell.PUM VPWR 0.01015f
C1469 XA.XIR[6].XIC[5].icell.Ien Iout 0.06821f
C1470 XThR.Tn[10] a_n997_2891# 0.1927f
C1471 XThC.Tn[8] XA.XIR[1].XIC[8].icell.Ien 0.03605f
C1472 XA.XIR[15].XIC[11].icell.Ien Vbias 0.15966f
C1473 XA.XIR[14].XIC[3].icell.Ien VPWR 0.19845f
C1474 XThC.Tn[9] XThR.Tn[7] 0.29362f
C1475 XThC.XTB4.Y Vbias 0.01548f
C1476 XA.XIR[13].XIC[5].icell.Ien VPWR 0.1979f
C1477 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.PDM 0.02104f
C1478 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PDM 0.04035f
C1479 XThC.XTB2.Y a_3523_10575# 0.01006f
C1480 XThR.XTB1.Y VPWR 1.13148f
C1481 XThC.XTB7.Y XThC.Tn[11] 0.07471f
C1482 XA.XIR[12].XIC[7].icell.PUM VPWR 0.01015f
C1483 XThR.XTB6.Y a_n1319_5611# 0.01283f
C1484 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.Ien 0.04854f
C1485 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.PDM 0.02104f
C1486 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PDM 0.0404f
C1487 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1488 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PDM 0.02765f
C1489 XA.XIR[11].XIC[8].icell.Ien VPWR 0.1979f
C1490 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PDM 0.02765f
C1491 XThR.XTB7.Y XThR.Tn[12] 0.07066f
C1492 XA.XIR[11].XIC[4].icell.Ien Iout 0.06821f
C1493 XThC.Tn[12] XA.XIR[7].XIC[12].icell.Ien 0.03605f
C1494 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.02787f
C1495 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.Ien 0.04854f
C1496 XA.XIR[10].XIC[6].icell.Ien Iout 0.06821f
C1497 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PDM 0.02765f
C1498 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PDM 0.02765f
C1499 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PDM 0.04035f
C1500 XA.XIR[3].XIC_15.icell.Ien Iout 0.0694f
C1501 XThR.Tn[4] XThR.Tn[5] 0.10984f
C1502 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PDM 0.04035f
C1503 XThC.Tn[8] XThR.Tn[3] 0.29362f
C1504 XA.XIR[2].XIC[12].icell.Ien VPWR 0.1979f
C1505 XA.XIR[10].XIC[0].icell.PUM VPWR 0.01015f
C1506 XA.XIR[2].XIC[8].icell.Ien Iout 0.06821f
C1507 XThC.Tn[3] XA.XIR[15].XIC[3].icell.Ien 0.03184f
C1508 XA.XIR[7].XIC[8].icell.PDM Vbias 0.03922f
C1509 XThC.Tn[5] VPWR 6.45659f
C1510 XA.XIR[1].XIC[14].icell.Ien VPWR 0.19796f
C1511 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PDM 0.04056f
C1512 XThR.Tn[8] XA.XIR[8].XIC[9].icell.Ien 0.15202f
C1513 XA.XIR[9].XIC[1].icell.Ien Vbias 0.19161f
C1514 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PDM 0.02765f
C1515 XA.XIR[1].XIC[10].icell.Ien Iout 0.06821f
C1516 XA.XIR[6].XIC_15.icell.PDM Vbias 0.03927f
C1517 XA.XIR[4].XIC[3].icell.Ien Vbias 0.19161f
C1518 XA.XIR[15].XIC[6].icell.PDM Vbias 0.03922f
C1519 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.PDM 0.02104f
C1520 XThR.XTB6.Y XThR.Tn[5] 0.20186f
C1521 XA.XIR[3].XIC_dummy_left.icell.Iout VPWR 0.11336f
C1522 XThC.Tn[14] XA.XIR[9].XIC[14].icell.Ien 0.03605f
C1523 XThC.Tn[11] XThR.Tn[0] 0.29385f
C1524 XThC.Tn[13] XThR.Tn[5] 0.29363f
C1525 XThC.Tn[4] XA.XIR[11].XIC[4].icell.Ien 0.03605f
C1526 XA.XIR[12].XIC[1].icell.Ien VPWR 0.1979f
C1527 XThC.Tn[8] XA.XIR[6].XIC[8].icell.Ien 0.03605f
C1528 XThR.Tn[5] XA.XIR[5].XIC[8].icell.Ien 0.15202f
C1529 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.Ien 0.04854f
C1530 XA.XIR[9].XIC[4].icell.PDM Vbias 0.03922f
C1531 XThR.XTBN.Y a_n997_1579# 0.23006f
C1532 XA.XIR[3].XIC_dummy_right.icell.Iout Iout 0.01732f
C1533 XA.XIR[5].XIC[2].icell.Ien VPWR 0.1979f
C1534 XThR.XTB7.Y a_n1049_5317# 0.27822f
C1535 XThC.XTB2.Y Vbias 0.0123f
C1536 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout 0.06446f
C1537 XThC.Tn[9] XA.XIR[12].XIC[9].icell.Ien 0.03605f
C1538 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.PDM 0.02104f
C1539 XA.XIR[9].XIC[6].icell.Ien Vbias 0.19161f
C1540 XA.XIR[15].XIC[10].icell.PDM VPWR 0.01334f
C1541 XA.XIR[4].XIC[5].icell.PUM VPWR 0.01015f
C1542 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PDM 0.02765f
C1543 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PDM 0.02765f
C1544 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.Ien 0.04854f
C1545 XThR.Tn[1] XA.XIR[1].XIC[13].icell.Ien 0.15202f
C1546 XA.XIR[1].XIC[9].icell.PDM Vbias 0.03922f
C1547 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.Ien 0.04854f
C1548 XA.XIR[7].XIC[2].icell.Ien Vbias 0.19161f
C1549 XA.XIR[4].XIC[9].icell.PDM Vbias 0.03922f
C1550 XA.XIR[5].XIC_15.icell.Ien Vbias 0.19195f
C1551 XA.XIR[9].XIC[8].icell.PUM VPWR 0.01015f
C1552 XThC.Tn[10] XThR.Tn[2] 0.29362f
C1553 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12] 0.15202f
C1554 XA.XIR[12].XIC_15.icell.PDM Vbias 0.03927f
C1555 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.Ien 0.04854f
C1556 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PDM 0.04035f
C1557 XThR.Tn[11] XThR.Tn[12] 0.15074f
C1558 XA.XIR[6].XIC[14].icell.Ien VPWR 0.19796f
C1559 XThC.Tn[12] XA.XIR[8].XIC[12].icell.Ien 0.03605f
C1560 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PDM 0.04035f
C1561 XThC.XTB7.A XThC.Tn[6] 0.10589f
C1562 XA.XIR[6].XIC[10].icell.Ien Iout 0.06821f
C1563 XA.XIR[7].XIC[4].icell.PUM VPWR 0.01015f
C1564 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PDM 0.04035f
C1565 Vbias Iout 74.00211f
C1566 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PDM 0.02765f
C1567 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1568 XThR.Tn[9] Vbias 1.4483f
C1569 XA.XIR[14].XIC[8].icell.Ien VPWR 0.19845f
C1570 XThC.Tn[13] XA.XIR[15].XIC[13].icell.Ien 0.03184f
C1571 XThR.XTB5.A XThR.XTBN.A 0.06303f
C1572 XA.XIR[14].XIC[4].icell.Ien Iout 0.06821f
C1573 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PDM 0.04035f
C1574 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.PDM 0.02104f
C1575 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PDM 0.02765f
C1576 XA.XIR[13].XIC[6].icell.Ien Iout 0.06821f
C1577 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.PDM 0.02104f
C1578 XThC.Tn[6] XA.XIR[2].XIC[6].icell.Ien 0.03605f
C1579 XThC.Tn[8] XThR.Tn[11] 0.29362f
C1580 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR 0.39006f
C1581 XA.XIR[15].XIC[0].icell.Ien Vbias 0.15953f
C1582 XA.XIR[11].XIC[9].icell.Ien Iout 0.06821f
C1583 XThR.XTBN.Y a_n1049_6699# 0.07601f
C1584 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PDM 0.04035f
C1585 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.PDM 0.02104f
C1586 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.PDM 0.02104f
C1587 XThC.Tn[7] XThR.Tn[7] 0.29362f
C1588 XA.XIR[13].XIC[0].icell.PUM VPWR 0.01015f
C1589 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PDM 0.04035f
C1590 XThC.XTB5.Y XThC.Tn[9] 0.01732f
C1591 XA.XIR[10].XIC[3].icell.PDM Vbias 0.03922f
C1592 XThC.Tn[4] Vbias 1.17728f
C1593 XThC.XTB6.Y XThC.Tn[13] 0.32552f
C1594 XThR.XTBN.A data[5] 0.0148f
C1595 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PDM 0.04035f
C1596 XThC.Tn[4] XA.XIR[14].XIC[4].icell.Ien 0.03605f
C1597 XThC.Tn[11] XThR.Tn[1] 0.29369f
C1598 XA.XIR[15].XIC[2].icell.PUM VPWR 0.01015f
C1599 XA.XIR[15].XIC[5].icell.Ien Vbias 0.15966f
C1600 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.PDM 0.02104f
C1601 XA.XIR[2].XIC[13].icell.Ien Iout 0.06821f
C1602 XThC.XTB6.A data[1] 0.37233f
C1603 XThR.Tn[8] XA.XIR[8].XIC[14].icell.Ien 0.15202f
C1604 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.Ien 0.04854f
C1605 XThR.XTB4.Y a_n1049_6699# 0.23756f
C1606 XA.XIR[10].XIC_dummy_left.icell.Iout XA.XIR[11].XIC_dummy_left.icell.Iout 0.03665f
C1607 XThR.XTB2.Y XThR.XTB7.A 0.2319f
C1608 XThR.XTB6.A XThR.XTB3.Y 0.03869f
C1609 XA.XIR[1].XIC_15.icell.Ien Iout 0.0694f
C1610 XThC.Tn[11] XThR.Tn[12] 0.29362f
C1611 XA.XIR[4].XIC[8].icell.Ien Vbias 0.19161f
C1612 XThC.Tn[1] XA.XIR[3].XIC[1].icell.Ien 0.03605f
C1613 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.Ien 0.04854f
C1614 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.PDM 0.02104f
C1615 XThR.XTB7.B XThR.Tn[8] 0.05091f
C1616 XThC.XTBN.Y XThC.Tn[9] 0.49746f
C1617 XA.XIR[8].XIC[2].icell.Ien Vbias 0.19161f
C1618 XThC.Tn[6] XThR.Tn[3] 0.29362f
C1619 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PDM 0.02765f
C1620 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.Ien 0.04854f
C1621 XThR.Tn[5] XA.XIR[5].XIC[13].icell.Ien 0.15202f
C1622 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR 0.08547f
C1623 XA.XIR[15].XIC[7].icell.PUM VPWR 0.01015f
C1624 XA.XIR[0].XIC[11].icell.PDM Vbias 0.03943f
C1625 XA.XIR[5].XIC[7].icell.Ien VPWR 0.1979f
C1626 XThR.XTB7.A a_n1049_5611# 0.01824f
C1627 XA.XIR[9].XIC[11].icell.Ien Vbias 0.19161f
C1628 XA.XIR[5].XIC[3].icell.Ien Iout 0.06821f
C1629 XThC.Tn[10] XThR.Tn[10] 0.29362f
C1630 XThC.Tn[0] XThR.Tn[0] 0.29747f
C1631 XThC.Tn[2] XThR.Tn[5] 0.29362f
C1632 XA.XIR[4].XIC[10].icell.PUM VPWR 0.01015f
C1633 XA.XIR[12].XIC[14].icell.PDM Vbias 0.03922f
C1634 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PDM 0.02765f
C1635 XA.XIR[1].XIC_dummy_right.icell.Iout Iout 0.01732f
C1636 XA.XIR[0].XIC[4].icell.Ien Vbias 0.19205f
C1637 XThC.Tn[9] XThC.Tn[10] 0.07959f
C1638 XA.XIR[8].XIC[4].icell.PUM VPWR 0.01015f
C1639 XThR.Tn[13] a_n997_1579# 0.19413f
C1640 XA.XIR[15].XIC_15.icell.PDM Vbias 0.03927f
C1641 XA.XIR[12].XIC[2].icell.Ien VPWR 0.1979f
C1642 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PDM 0.04035f
C1643 XA.XIR[0].XIC_15.icell.PDM VPWR 0.07389f
C1644 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.PDM 0.02104f
C1645 XThC.XTB7.Y VPWR 1.07717f
C1646 XA.XIR[7].XIC[7].icell.Ien Vbias 0.19161f
C1647 XA.XIR[9].XIC[13].icell.PUM VPWR 0.01015f
C1648 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.PDM 0.02104f
C1649 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.PDM 0.02104f
C1650 XThR.Tn[4] XA.XIR[4].XIC[3].icell.Ien 0.15202f
C1651 XThC.XTBN.A XThC.XTB6.Y 0.06405f
C1652 XThR.XTBN.A XThR.Tn[9] 0.12398f
C1653 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.PDM 0.02104f
C1654 XThR.Tn[6] Iout 1.19569f
C1655 XA.XIR[11].XIC[14].icell.Ien Iout 0.06821f
C1656 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.Ien 0.04854f
C1657 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1658 XA.XIR[6].XIC_15.icell.Ien Iout 0.0694f
C1659 XA.XIR[7].XIC[9].icell.PUM VPWR 0.01015f
C1660 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.02765f
C1661 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.PDM 0.02104f
C1662 XThC.Tn[8] XThR.Tn[14] 0.29362f
C1663 XThR.XTB6.A VPWR 0.68638f
C1664 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PDM 0.04035f
C1665 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.Ien 0.04854f
C1666 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Iout 0.01728f
C1667 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR 0.39003f
C1668 a_6243_9615# Vbias 0.01017f
C1669 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PDM 0.02765f
C1670 XA.XIR[6].XIC[2].icell.PDM Vbias 0.03922f
C1671 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.Ien 0.04854f
C1672 XA.XIR[14].XIC[9].icell.Ien Iout 0.06821f
C1673 XThC.Tn[9] XA.XIR[15].XIC[9].icell.Ien 0.03184f
C1674 XThR.XTB1.Y a_n1049_8581# 0.21263f
C1675 XA.XIR[5].XIC[9].icell.PDM Vbias 0.03922f
C1676 XThR.Tn[3] XA.XIR[3].XIC[6].icell.Ien 0.15202f
C1677 XThC.Tn[5] XA.XIR[0].XIC[5].icell.Ien 0.037f
C1678 XA.XIR[6].XIC[0].icell.PUM VPWR 0.01015f
C1679 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.PDM 0.02104f
C1680 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.Ien 0.04854f
C1681 XThR.Tn[0] VPWR 8.31136f
C1682 XA.XIR[13].XIC[3].icell.PDM Vbias 0.03922f
C1683 XThC.XTB4.Y XThC.XTBN.A 0.03415f
C1684 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PDM 0.04035f
C1685 XA.XIR[12].XIC[8].icell.PDM Vbias 0.03922f
C1686 XThR.XTB7.B XThR.XTB2.Y 0.22599f
C1687 XA.XIR[10].XIC[1].icell.PUM VPWR 0.01015f
C1688 XThR.XTB7.B a_n997_3755# 0.01174f
C1689 XA.XIR[6].XIC_dummy_right.icell.Iout Iout 0.01732f
C1690 XThC.Tn[4] XThR.Tn[6] 0.29362f
C1691 XA.XIR[5].XIC_dummy_right.icell.Iout XA.XIR[6].XIC_dummy_right.icell.Iout 0.04047f
C1692 XThR.XTBN.Y XThR.Tn[8] 0.47831f
C1693 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.Ien 0.04854f
C1694 XThC.Tn[7] XA.XIR[4].XIC[7].icell.Ien 0.03605f
C1695 XThC.Tn[6] XThR.Tn[11] 0.29362f
C1696 XA.XIR[10].XIC[13].icell.Ien Vbias 0.19161f
C1697 XA.XIR[3].XIC[4].icell.Ien Vbias 0.19161f
C1698 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.PDM 0.02104f
C1699 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.PDM 0.02104f
C1700 XThR.Tn[4] Iout 1.19572f
C1701 XThC.XTB3.Y XThC.XTB6.Y 0.04428f
C1702 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.Ien 0.04854f
C1703 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.Ien 0.04854f
C1704 XA.XIR[9].XIC[3].icell.Ien VPWR 0.1979f
C1705 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PDM 0.02765f
C1706 XA.XIR[8].XIC[6].icell.PDM Vbias 0.03922f
C1707 XA.XIR[3].XIC[4].icell.PDM Vbias 0.03922f
C1708 XA.XIR[12].XIC[13].icell.PDM Vbias 0.03922f
C1709 XA.XIR[4].XIC[13].icell.Ien Vbias 0.19161f
C1710 XThR.XTB4.Y XThR.Tn[8] 0.01306f
C1711 XThC.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.03605f
C1712 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.Ien 0.04854f
C1713 XA.XIR[11].XIC[12].icell.Ien Iout 0.06821f
C1714 XA.XIR[2].XIC[10].icell.PDM Vbias 0.03922f
C1715 XThC.Tn[10] XThR.Tn[13] 0.29362f
C1716 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.02765f
C1717 XThC.Tn[0] XA.XIR[4].XIC[0].icell.Ien 0.03605f
C1718 XA.XIR[8].XIC[7].icell.Ien Vbias 0.19161f
C1719 XThC.Tn[0] XThR.Tn[1] 0.29406f
C1720 XA.XIR[15].XIC[14].icell.PDM Vbias 0.03922f
C1721 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PDM 0.02765f
C1722 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PDM 0.04035f
C1723 XA.XIR[3].XIC[6].icell.PUM VPWR 0.01015f
C1724 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.02765f
C1725 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.PDM 0.02104f
C1726 XThR.XTB6.Y XThR.Tn[9] 0.0246f
C1727 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.Ien 0.04854f
C1728 XThR.XTB7.A XThR.Tn[3] 0.0306f
C1729 XThC.Tn[13] Iout 0.84487f
C1730 XThC.Tn[13] XThR.Tn[9] 0.29363f
C1731 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.PDM 0.02104f
C1732 XA.XIR[5].XIC[12].icell.Ien VPWR 0.1979f
C1733 XThC.Tn[0] XThR.Tn[12] 0.29366f
C1734 XThC.Tn[9] XThR.Tn[8] 0.29362f
C1735 XA.XIR[5].XIC[8].icell.Ien Iout 0.06821f
C1736 XThC.XTB6.A VPWR 0.68179f
C1737 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.PDM 0.02104f
C1738 XA.XIR[4].XIC_15.icell.PUM VPWR 0.01655f
C1739 XThC.XTB7.B XThC.XTB7.Y 0.33493f
C1740 XA.XIR[10].XIC_dummy_left.icell.Iout Iout 0.0353f
C1741 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Iout 0.01779f
C1742 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.PDM 0.02104f
C1743 XThR.XTB7.A data[4] 0.8689f
C1744 XThR.XTB7.A XThR.XTB7.Y 0.37429f
C1745 XThC.XTBN.A a_7875_9569# 0.01939f
C1746 XA.XIR[2].XIC[14].icell.PDM VPWR 0.01002f
C1747 XA.XIR[0].XIC[9].icell.Ien Vbias 0.19209f
C1748 XThC.XTBN.Y XThC.Tn[7] 0.91493f
C1749 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PDM 0.04035f
C1750 XThC.Tn[4] XThR.Tn[4] 0.29362f
C1751 XA.XIR[8].XIC[9].icell.PUM VPWR 0.01015f
C1752 XThC.XTB2.Y XThC.XTBN.A 0.04716f
C1753 XThC.XTB3.Y XThC.XTB4.Y 2.13136f
C1754 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.PDM 0.02104f
C1755 XA.XIR[12].XIC[7].icell.Ien VPWR 0.1979f
C1756 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1757 XA.XIR[7].XIC_dummy_right.icell.Iout XA.XIR[8].XIC_dummy_right.icell.Iout 0.04047f
C1758 XA.XIR[12].XIC[3].icell.Ien Iout 0.06821f
C1759 XThC.Tn[5] XA.XIR[3].XIC[5].icell.Ien 0.03605f
C1760 XA.XIR[7].XIC[12].icell.Ien Vbias 0.19161f
C1761 XA.XIR[14].XIC[14].icell.Ien Iout 0.06821f
C1762 XThC.Tn[12] XA.XIR[2].XIC[12].icell.Ien 0.03605f
C1763 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR 0.01669f
C1764 XThR.Tn[4] XA.XIR[4].XIC[8].icell.Ien 0.15202f
C1765 XThR.Tn[11] XA.XIR[11].XIC[13].icell.Ien 0.15202f
C1766 XA.XIR[10].XIC[11].icell.Ien Vbias 0.19161f
C1767 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.PDM 0.02104f
C1768 XA.XIR[3].XIC[1].icell.Ien Vbias 0.19161f
C1769 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR 0.38996f
C1770 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PDM 0.04035f
C1771 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PDM 0.04035f
C1772 XThC.XTB1.Y XThC.XTB6.Y 0.05752f
C1773 XA.XIR[7].XIC[14].icell.PUM VPWR 0.01015f
C1774 XA.XIR[1].XIC[0].icell.Ien VPWR 0.1979f
C1775 XThR.XTBN.Y XThR.XTB2.Y 0.2075f
C1776 XThR.XTBN.Y a_n997_3755# 0.229f
C1777 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.PDM 0.02104f
C1778 XThR.Tn[2] XA.XIR[2].XIC[1].icell.Ien 0.15202f
C1779 XA.XIR[7].XIC[10].icell.PDM Vbias 0.03922f
C1780 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.Ien 0.04854f
C1781 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.Ien 0.04854f
C1782 XA.XIR[11].XIC[10].icell.Ien Iout 0.06821f
C1783 XThR.Tn[1] VPWR 8.31638f
C1784 XA.XIR[4].XIC[0].icell.Ien VPWR 0.1979f
C1785 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PDM 0.02765f
C1786 XA.XIR[15].XIC[8].icell.PDM Vbias 0.03922f
C1787 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.Ien 0.04854f
C1788 XA.XIR[13].XIC[1].icell.PUM VPWR 0.01015f
C1789 XThR.Tn[12] XA.XIR[12].XIC[6].icell.Ien 0.15202f
C1790 XThC.XTBN.Y a_3773_9615# 0.08456f
C1791 XThR.Tn[3] XA.XIR[3].XIC[11].icell.Ien 0.15202f
C1792 XThR.Tn[12] VPWR 9.21906f
C1793 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.PDM 0.02104f
C1794 XA.XIR[13].XIC_dummy_left.icell.Iout XA.XIR[14].XIC_dummy_left.icell.Iout 0.03665f
C1795 XThR.XTBN.Y a_n1049_5611# 0.0768f
C1796 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.Ien 0.04854f
C1797 XA.XIR[9].XIC[6].icell.PDM Vbias 0.03922f
C1798 XThR.XTB2.Y XThR.XTB4.Y 0.04006f
C1799 XThC.Tn[6] XThR.Tn[14] 0.29362f
C1800 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.Ien 0.04854f
C1801 XA.XIR[13].XIC[13].icell.Ien Vbias 0.19161f
C1802 XA.XIR[15].XIC[2].icell.Ien VPWR 0.33655f
C1803 XA.XIR[11].XIC[0].icell.Ien Iout 0.06814f
C1804 XA.XIR[7].XIC[14].icell.PDM VPWR 0.01002f
C1805 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.PDM 0.02104f
C1806 XThR.Tn[2] XA.XIR[2].XIC[6].icell.Ien 0.15202f
C1807 XA.XIR[12].XIC[12].icell.PDM Vbias 0.03922f
C1808 XThC.Tn[3] XA.XIR[10].XIC[3].icell.Ien 0.03605f
C1809 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.PDM 0.02104f
C1810 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.Ien 0.04854f
C1811 XThC.XTB1.Y XThC.XTB4.Y 0.05121f
C1812 XThC.XTB2.Y XThC.XTB3.Y 2.04808f
C1813 XA.XIR[4].XIC[5].icell.Ien VPWR 0.1979f
C1814 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PDM 0.02765f
C1815 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.PDM 0.02104f
C1816 XThC.XTB2.Y XThC.Tn[2] 0.01113f
C1817 XA.XIR[15].XIC[13].icell.PDM Vbias 0.03922f
C1818 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1819 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.PDM 0.02104f
C1820 XA.XIR[3].XIC[9].icell.Ien Vbias 0.19161f
C1821 XA.XIR[1].XIC[11].icell.PDM Vbias 0.03922f
C1822 XA.XIR[14].XIC[12].icell.Ien Iout 0.06821f
C1823 XThC.Tn[6] XA.XIR[5].XIC[6].icell.Ien 0.03605f
C1824 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PDM 0.02765f
C1825 XThC.Tn[8] VPWR 7.39788f
C1826 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1827 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.Ien 0.04854f
C1828 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PDM 0.02765f
C1829 XA.XIR[2].XIC[2].icell.Ien Vbias 0.19161f
C1830 XA.XIR[4].XIC[11].icell.PDM Vbias 0.03922f
C1831 XThR.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.15202f
C1832 XA.XIR[9].XIC[8].icell.Ien VPWR 0.1979f
C1833 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.Ien 0.04854f
C1834 XA.XIR[1].XIC[4].icell.Ien Vbias 0.19173f
C1835 XA.XIR[7].XIC[0].icell.PUM VPWR 0.01015f
C1836 XThR.XTB7.B data[4] 0.01382f
C1837 XThR.XTB7.B XThR.XTB7.Y 0.33493f
C1838 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.Ien 0.04854f
C1839 XThR.Tn[9] XA.XIR[9].XIC[4].icell.Ien 0.15202f
C1840 XA.XIR[9].XIC[4].icell.Ien Iout 0.06821f
C1841 XThC.XTB6.A XThC.XTB7.B 1.47641f
C1842 XThC.Tn[2] XA.XIR[7].XIC[2].icell.Ien 0.03605f
C1843 XThR.XTB5.Y a_n1319_6405# 0.01188f
C1844 XA.XIR[8].XIC[12].icell.Ien Vbias 0.19161f
C1845 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PDM 0.04035f
C1846 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.PDM 0.02104f
C1847 a_n1049_5317# VPWR 0.72036f
C1848 XA.XIR[13].XIC_dummy_left.icell.Iout Iout 0.0353f
C1849 XA.XIR[3].XIC[11].icell.PUM VPWR 0.01015f
C1850 XA.XIR[1].XIC_15.icell.PDM VPWR 0.07527f
C1851 XA.XIR[2].XIC[4].icell.PUM VPWR 0.01015f
C1852 XA.XIR[7].XIC[4].icell.Ien VPWR 0.1979f
C1853 XA.XIR[4].XIC_15.icell.PDM VPWR 0.07527f
C1854 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.Ien 0.04854f
C1855 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.PDM 0.02104f
C1856 XThR.Tn[2] XThR.Tn[3] 0.1415f
C1857 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1858 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.PDM 0.02104f
C1859 XA.XIR[5].XIC[13].icell.Ien Iout 0.06821f
C1860 XA.XIR[1].XIC[6].icell.PUM VPWR 0.01015f
C1861 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout 0.06446f
C1862 XThR.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.1525f
C1863 XA.XIR[0].XIC[14].icell.Ien Vbias 0.19209f
C1864 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PDM 0.04056f
C1865 XA.XIR[8].XIC[14].icell.PUM VPWR 0.01015f
C1866 XThC.Tn[2] Iout 0.85054f
C1867 XThC.Tn[2] XThR.Tn[9] 0.29362f
C1868 XA.XIR[13].XIC[11].icell.Ien Vbias 0.19161f
C1869 XThR.XTBN.Y a_n997_715# 0.21503f
C1870 XThR.Tn[7] XA.XIR[7].XIC[1].icell.Ien 0.15202f
C1871 XA.XIR[11].XIC_15.icell.Ien Iout 0.0694f
C1872 XThC.Tn[4] XA.XIR[9].XIC[4].icell.Ien 0.03605f
C1873 VPWR data[7] 0.212f
C1874 XA.XIR[12].XIC[8].icell.Ien Iout 0.06821f
C1875 XThC.Tn[7] XThR.Tn[8] 0.29362f
C1876 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.Ien 0.04854f
C1877 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.PDM 0.02104f
C1878 XThC.XTB1.Y XThC.XTB2.Y 2.14864f
C1879 XThC.Tn[11] XA.XIR[0].XIC[11].icell.Ien 0.03728f
C1880 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PDM 0.04035f
C1881 XThR.Tn[4] XA.XIR[4].XIC[13].icell.Ien 0.15202f
C1882 XA.XIR[11].XIC[1].icell.PDM Vbias 0.03922f
C1883 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR 0.01499f
C1884 XThR.Tn[0] XA.XIR[0].XIC[5].icell.Ien 0.15202f
C1885 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.Ien 0.04854f
C1886 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PDM 0.04035f
C1887 XThR.Tn[10] XA.XIR[10].XIC[4].icell.Ien 0.15202f
C1888 XThR.XTB7.B a_n997_2667# 0.02071f
C1889 XThC.Tn[5] XA.XIR[1].XIC[5].icell.Ien 0.03605f
C1890 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PDM 0.02765f
C1891 XA.XIR[14].XIC[10].icell.Ien Iout 0.06821f
C1892 XThC.Tn[13] XA.XIR[10].XIC[13].icell.Ien 0.03605f
C1893 XA.XIR[10].XIC[5].icell.PDM Vbias 0.03922f
C1894 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.PDM 0.02104f
C1895 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PDM 0.04035f
C1896 XA.XIR[6].XIC[1].icell.PUM VPWR 0.01015f
C1897 XThC.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.03605f
C1898 a_n1049_6405# VPWR 0.72095f
C1899 XThR.Tn[7] XA.XIR[7].XIC[6].icell.Ien 0.15202f
C1900 XA.XIR[6].XIC[4].icell.Ien Vbias 0.19161f
C1901 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.Ien 0.04854f
C1902 XA.XIR[8].XIC_dummy_left.icell.Ien XThR.Tn[8] 0.01438f
C1903 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.Ien 0.04854f
C1904 XA.XIR[11].XIC_dummy_right.icell.Iout Iout 0.01732f
C1905 XThC.Tn[2] XThC.Tn[4] 0.02725f
C1906 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PDM 0.02765f
C1907 XThC.Tn[13] XA.XIR[4].XIC[13].icell.Ien 0.03605f
C1908 XA.XIR[12].XIC[11].icell.PDM Vbias 0.03922f
C1909 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.PDM 0.02104f
C1910 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.Ien 0.04854f
C1911 XA.XIR[4].XIC[1].icell.Ien Iout 0.06821f
C1912 XA.XIR[15].XIC[12].icell.PDM Vbias 0.03922f
C1913 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.Ien 0.04854f
C1914 XThC.Tn[1] XA.XIR[12].XIC[1].icell.Ien 0.03605f
C1915 XThC.Tn[3] XA.XIR[13].XIC[3].icell.Ien 0.03605f
C1916 XThR.XTBN.Y XThR.Tn[3] 0.62502f
C1917 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.PDM 0.02104f
C1918 XA.XIR[11].XIC_dummy_left.icell.Ien XThR.Tn[11] 0.01432f
C1919 a_n1049_8581# XThR.Tn[0] 0.2685f
C1920 XA.XIR[6].XIC[6].icell.PUM VPWR 0.01015f
C1921 XThR.XTB7.B XThR.Tn[11] 0.03888f
C1922 XThC.Tn[10] XThR.Tn[7] 0.29362f
C1923 XA.XIR[0].XIC[13].icell.PDM Vbias 0.03943f
C1924 XA.XIR[15].XIC[7].icell.Ien VPWR 0.33655f
C1925 XA.XIR[11].XIC[3].icell.Ien Vbias 0.19161f
C1926 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.Ien 0.04854f
C1927 XThC.XTB7.B XThC.Tn[8] 0.09736f
C1928 XThC.Tn[2] XA.XIR[8].XIC[2].icell.Ien 0.03605f
C1929 XThC.Tn[0] XA.XIR[2].XIC[0].icell.Ien 0.03605f
C1930 XThR.Tn[2] XA.XIR[2].XIC[11].icell.Ien 0.15202f
C1931 XA.XIR[15].XIC[3].icell.Ien Iout 0.07211f
C1932 XThR.XTBN.Y XThR.XTB7.Y 0.50018f
C1933 XA.XIR[10].XIC[5].icell.Ien Vbias 0.19161f
C1934 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR 0.38903f
C1935 XThC.XTB7.Y XThC.Tn[12] 0.07222f
C1936 XA.XIR[4].XIC[10].icell.Ien VPWR 0.1979f
C1937 XA.XIR[0].XIC[1].icell.Ien VPWR 0.19726f
C1938 XA.XIR[4].XIC[6].icell.Ien Iout 0.06821f
C1939 XA.XIR[11].XIC[14].icell.PUM VPWR 0.01015f
C1940 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.PDM 0.02104f
C1941 XA.XIR[8].XIC[4].icell.Ien VPWR 0.1979f
C1942 XThR.XTB4.Y XThR.Tn[3] 0.1895f
C1943 XA.XIR[3].XIC[14].icell.Ien Vbias 0.19161f
C1944 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.PDM 0.02104f
C1945 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.Ien 0.04854f
C1946 XA.XIR[11].XIC[5].icell.PUM VPWR 0.01015f
C1947 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PDM 0.04035f
C1948 XA.XIR[2].XIC[7].icell.Ien Vbias 0.19161f
C1949 XThC.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.03605f
C1950 XA.XIR[7].XIC[0].icell.Ien Iout 0.06814f
C1951 XA.XIR[9].XIC[13].icell.Ien VPWR 0.1979f
C1952 XThR.XTB4.Y XThR.XTB7.Y 0.03475f
C1953 XA.XIR[10].XIC[7].icell.PUM VPWR 0.01015f
C1954 XA.XIR[1].XIC[9].icell.Ien Vbias 0.19173f
C1955 XA.XIR[9].XIC[9].icell.Ien Iout 0.06821f
C1956 XThC.Tn[11] XA.XIR[3].XIC[11].icell.Ien 0.03605f
C1957 XThR.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.15202f
C1958 XThC.Tn[9] XThR.Tn[3] 0.29362f
C1959 XA.XIR[0].XIC[6].icell.Ien VPWR 0.19733f
C1960 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.Ien 0.04854f
C1961 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1962 XThC.Tn[6] XA.XIR[12].XIC[6].icell.Ien 0.03605f
C1963 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1964 XThR.XTB7.Y XThR.Tn[10] 0.07406f
C1965 XA.XIR[0].XIC[2].icell.Ien Iout 0.06775f
C1966 XThC.Tn[6] VPWR 6.46044f
C1967 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.Ien 0.04854f
C1968 XA.XIR[2].XIC[9].icell.PUM VPWR 0.01015f
C1969 XThR.Tn[5] XA.XIR[5].XIC[0].icell.Ien 0.15228f
C1970 XA.XIR[7].XIC[9].icell.Ien VPWR 0.1979f
C1971 XThR.Tn[14] XA.XIR[14].XIC[13].icell.Ien 0.15202f
C1972 XThC.Tn[12] XThR.Tn[0] 0.29452f
C1973 XA.XIR[14].XIC_15.icell.Ien Iout 0.0694f
C1974 XA.XIR[1].XIC[11].icell.PUM VPWR 0.01015f
C1975 XA.XIR[7].XIC[5].icell.Ien Iout 0.06821f
C1976 XThC.Tn[14] XThR.Tn[5] 0.29368f
C1977 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PDM 0.04035f
C1978 XThR.XTBN.Y a_n997_2667# 0.22784f
C1979 XA.XIR[9].XIC_dummy_left.icell.Iout XA.XIR[10].XIC_dummy_left.icell.Iout 0.03665f
C1980 XA.XIR[6].XIC[4].icell.PDM Vbias 0.03922f
C1981 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1982 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.PDM 0.02104f
C1983 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.PDM 0.02104f
C1984 XThR.Tn[8] a_n997_3979# 0.1927f
C1985 XA.XIR[5].XIC[11].icell.PDM Vbias 0.03922f
C1986 XA.XIR[14].XIC[1].icell.PDM Vbias 0.03922f
C1987 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.Ien 0.04854f
C1988 XA.XIR[2].XIC[0].icell.Ien VPWR 0.1979f
C1989 XThC.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.03605f
C1990 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PDM 0.02765f
C1991 XA.XIR[13].XIC[5].icell.PDM Vbias 0.03922f
C1992 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PDM 0.04035f
C1993 XThR.Tn[11] XA.XIR[11].XIC[5].icell.Ien 0.15202f
C1994 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PDM 0.02765f
C1995 XA.XIR[12].XIC[10].icell.PDM Vbias 0.03922f
C1996 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Ien 0.01746f
C1997 XThC.Tn[11] XA.XIR[14].XIC[11].icell.Ien 0.03605f
C1998 XA.XIR[10].XIC[1].icell.Ien VPWR 0.1979f
C1999 XA.XIR[11].XIC[12].icell.PUM VPWR 0.01015f
C2000 XThR.XTB4.Y a_n997_2667# 0.07199f
C2001 XA.XIR[14].XIC_dummy_right.icell.Iout Iout 0.01732f
C2002 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PDM 0.02765f
C2003 XThR.Tn[0] XA.XIR[0].XIC[10].icell.Ien 0.15202f
C2004 XThR.Tn[10] XA.XIR[10].XIC[9].icell.Ien 0.15202f
C2005 XA.XIR[15].XIC[11].icell.PDM Vbias 0.03922f
C2006 XA.XIR[5].XIC_15.icell.PDM VPWR 0.07527f
C2007 XThR.Tn[6] XA.XIR[6].XIC[4].icell.Ien 0.15202f
C2008 XThC.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.03605f
C2009 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.Ien 0.04854f
C2010 XThR.XTBN.Y XThR.Tn[11] 0.52268f
C2011 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.Ien 0.04854f
C2012 XThC.Tn[11] XThR.Tn[2] 0.29362f
C2013 XA.XIR[6].XIC[9].icell.Ien Vbias 0.19161f
C2014 XThR.Tn[7] XA.XIR[7].XIC[11].icell.Ien 0.15202f
C2015 XThC.XTB7.Y a_10915_9569# 0.06874f
C2016 XThR.XTB7.A XThR.XTB3.Y 0.57441f
C2017 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2018 XThC.Tn[12] XA.XIR[5].XIC[12].icell.Ien 0.03605f
C2019 XA.XIR[8].XIC[8].icell.PDM Vbias 0.03922f
C2020 XA.XIR[3].XIC[6].icell.PDM Vbias 0.03922f
C2021 XA.XIR[14].XIC[3].icell.Ien Vbias 0.19161f
C2022 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout 0.06446f
C2023 XThR.Tn[7] XThR.Tn[8] 0.11022f
C2024 XA.XIR[11].XIC[13].icell.Ien VPWR 0.1979f
C2025 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.PDM 0.02104f
C2026 XA.XIR[2].XIC[12].icell.PDM Vbias 0.03922f
C2027 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.Ien 0.04854f
C2028 XA.XIR[13].XIC[5].icell.Ien Vbias 0.19161f
C2029 XA.XIR[3].XIC[6].icell.Ien VPWR 0.1979f
C2030 XThR.Tn[14] XA.XIR[14].XIC[11].icell.Ien 0.15202f
C2031 XThR.XTB4.Y XThR.Tn[11] 0.3042f
C2032 XA.XIR[14].XIC[14].icell.PUM VPWR 0.01015f
C2033 XA.XIR[6].XIC[11].icell.PUM VPWR 0.01015f
C2034 XThC.Tn[8] XA.XIR[7].XIC[8].icell.Ien 0.03605f
C2035 XA.XIR[3].XIC[2].icell.Ien Iout 0.06821f
C2036 XA.XIR[11].XIC[8].icell.Ien Vbias 0.19161f
C2037 XThR.Tn[10] XThR.Tn[11] 0.09505f
C2038 XA.XIR[15].XIC[8].icell.Ien Iout 0.07211f
C2039 XA.XIR[4].XIC_15.icell.Ien VPWR 0.26829f
C2040 XA.XIR[14].XIC[5].icell.PUM VPWR 0.01015f
C2041 XThC.XTB5.Y XThC.XTBN.Y 0.162f
C2042 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout 0.06446f
C2043 XThC.Tn[9] XThR.Tn[11] 0.29362f
C2044 XThC.XTBN.A a_8963_9569# 0.01679f
C2045 XA.XIR[4].XIC[11].icell.Ien Iout 0.06821f
C2046 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2047 XA.XIR[13].XIC[7].icell.PUM VPWR 0.01015f
C2048 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PDM 0.04035f
C2049 XThC.XTBN.A data[0] 0.02545f
C2050 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PDM 0.04035f
C2051 XA.XIR[8].XIC[9].icell.Ien VPWR 0.1979f
C2052 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PDM 0.02765f
C2053 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.Ien 0.04854f
C2054 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.Ien 0.04854f
C2055 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.PDM 0.02104f
C2056 XA.XIR[8].XIC[5].icell.Ien Iout 0.06821f
C2057 XThR.XTB7.Y XThR.Tn[13] 0.10781f
C2058 XA.XIR[11].XIC[10].icell.PUM VPWR 0.01015f
C2059 XThC.XTB7.B XThC.Tn[6] 0.05039f
C2060 XA.XIR[2].XIC[12].icell.Ien Vbias 0.19161f
C2061 XThC.XTB5.Y XThC.Tn[10] 0.01742f
C2062 XA.XIR[1].XIC[14].icell.Ien Vbias 0.19173f
C2063 XThC.Tn[5] Vbias 1.00831f
C2064 XThC.Tn[10] XA.XIR[9].XIC[10].icell.Ien 0.03605f
C2065 XA.XIR[9].XIC[14].icell.Ien Iout 0.06821f
C2066 XThR.Tn[9] XA.XIR[9].XIC[14].icell.Ien 0.15202f
C2067 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.Ien 0.04854f
C2068 XA.XIR[0].XIC[11].icell.Ien VPWR 0.19832f
C2069 XA.XIR[4].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2070 XThR.Tn[12] XA.XIR[12].XIC_dummy_left.icell.Iout 0.0404f
C2071 XThC.Tn[12] XThR.Tn[1] 0.29369f
C2072 XA.XIR[0].XIC[7].icell.Ien Iout 0.06775f
C2073 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PDM 0.04056f
C2074 XA.XIR[12].XIC[1].icell.Ien Vbias 0.19161f
C2075 XA.XIR[6].XIC_dummy_left.icell.Iout XA.XIR[7].XIC_dummy_left.icell.Iout 0.03665f
C2076 XA.XIR[11].XIC[0].icell.PUM VPWR 0.01015f
C2077 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PDM 0.0404f
C2078 XThC.Tn[11] XA.XIR[1].XIC[11].icell.Ien 0.03611f
C2079 XA.XIR[2].XIC[14].icell.PUM VPWR 0.01015f
C2080 XThR.XTB5.Y XThR.XTBN.A 0.10854f
C2081 XA.XIR[7].XIC[14].icell.Ien VPWR 0.19796f
C2082 XThC.Tn[12] XThR.Tn[12] 0.29362f
C2083 XThR.XTB7.A VPWR 0.88595f
C2084 XThR.Tn[13] XA.XIR[13].XIC[4].icell.Ien 0.15202f
C2085 XThR.Tn[10] XA.XIR[10].XIC[14].icell.Ien 0.15202f
C2086 XA.XIR[7].XIC[10].icell.Ien Iout 0.06821f
C2087 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2088 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PDM 0.02765f
C2089 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Iout 0.04497f
C2090 XA.XIR[5].XIC[2].icell.Ien Vbias 0.19161f
C2091 XA.XIR[11].XIC[11].icell.Ien VPWR 0.1979f
C2092 XA.XIR[7].XIC[12].icell.PDM Vbias 0.03922f
C2093 XThC.XTBN.Y XThC.Tn[10] 0.51405f
C2094 XThC.Tn[7] XThR.Tn[3] 0.29362f
C2095 XA.XIR[15].XIC[10].icell.PDM Vbias 0.03922f
C2096 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PDM 0.02765f
C2097 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.PDM 0.02104f
C2098 XA.XIR[13].XIC[1].icell.Ien VPWR 0.1979f
C2099 XThC.XTBN.Y a_4861_9615# 0.07601f
C2100 XA.XIR[14].XIC[12].icell.PUM VPWR 0.01015f
C2101 XA.XIR[8].XIC[0].icell.Ien Iout 0.06814f
C2102 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PDM 0.02765f
C2103 XThC.Tn[1] XThR.Tn[0] 0.29448f
C2104 XThC.Tn[11] XThR.Tn[10] 0.29362f
C2105 XThC.Tn[3] XThR.Tn[5] 0.29362f
C2106 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.Ien 0.04854f
C2107 XA.XIR[9].XIC[8].icell.PDM Vbias 0.03922f
C2108 XThC.XTB5.Y a_5155_10571# 0.01188f
C2109 XThR.XTB7.B XThR.XTB3.Y 0.23315f
C2110 XThC.Tn[9] XA.XIR[13].XIC[9].icell.Ien 0.03605f
C2111 XA.XIR[0].XIC[0].icell.PDM Vbias 0.03935f
C2112 XThR.XTBN.Y XThR.Tn[14] 0.47807f
C2113 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.Ien 0.04854f
C2114 XA.XIR[5].XIC[4].icell.PUM VPWR 0.01015f
C2115 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2116 XThC.XTB3.Y data[0] 0.03253f
C2117 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PDM 0.02765f
C2118 XThR.Tn[0] XA.XIR[0].XIC_15.icell.Ien 0.13564f
C2119 XThR.Tn[6] XA.XIR[6].XIC[9].icell.Ien 0.15202f
C2120 XThC.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.03605f
C2121 XA.XIR[14].XIC[13].icell.Ien VPWR 0.19845f
C2122 XA.XIR[1].XIC[13].icell.PDM Vbias 0.03922f
C2123 XA.XIR[6].XIC[14].icell.Ien Vbias 0.19161f
C2124 XThC.Tn[6] XA.XIR[15].XIC[6].icell.Ien 0.03184f
C2125 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.PDM 0.02104f
C2126 XThR.XTB1.Y XThR.XTBN.A 0.12307f
C2127 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout 0.06446f
C2128 XA.XIR[4].XIC[13].icell.PDM Vbias 0.03922f
C2129 XA.XIR[1].XIC[1].icell.Ien VPWR 0.1979f
C2130 XThR.XTB3.Y XThR.Tn[2] 0.18254f
C2131 XA.XIR[10].XIC[2].icell.Ien VPWR 0.1979f
C2132 XA.XIR[14].XIC[8].icell.Ien Vbias 0.19161f
C2133 XThC.Tn[7] XA.XIR[11].XIC[7].icell.Ien 0.03605f
C2134 XThC.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.03605f
C2135 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.Ien 0.04854f
C2136 XThC.Tn[11] XA.XIR[6].XIC[11].icell.Ien 0.03605f
C2137 XThC.Tn[0] XThR.Tn[2] 0.29389f
C2138 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PDM 0.04035f
C2139 XThR.XTB5.Y XThR.Tn[4] 0.19957f
C2140 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PDM 0.04035f
C2141 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PDM 0.04035f
C2142 XA.XIR[3].XIC[11].icell.Ien VPWR 0.1979f
C2143 XThC.Tn[9] XThR.Tn[14] 0.29362f
C2144 XThR.Tn[10] XA.XIR[10].XIC[12].icell.Ien 0.15202f
C2145 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PDM 0.02765f
C2146 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2147 XA.XIR[3].XIC[7].icell.Ien Iout 0.06821f
C2148 XA.XIR[2].XIC[4].icell.Ien VPWR 0.1979f
C2149 XThR.Tn[1] a_n1049_7787# 0.26879f
C2150 XA.XIR[1].XIC[6].icell.Ien VPWR 0.1979f
C2151 XA.XIR[14].XIC[10].icell.PUM VPWR 0.01015f
C2152 XThR.XTB5.Y XThR.XTB6.Y 2.12831f
C2153 XA.XIR[1].XIC[2].icell.Ien Iout 0.06821f
C2154 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.PDM 0.02104f
C2155 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.Ien 0.04854f
C2156 XA.XIR[8].XIC[14].icell.Ien VPWR 0.19796f
C2157 XA.XIR[8].XIC[10].icell.Ien Iout 0.06821f
C2158 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR 0.38915f
C2159 XThC.Tn[5] XThR.Tn[6] 0.29362f
C2160 XThR.Tn[7] XA.XIR[7].XIC_dummy_left.icell.Iout 0.04675f
C2161 XThR.XTB7.B VPWR 1.67447f
C2162 XThC.XTB1.Y data[0] 0.06453f
C2163 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.PDM 0.02104f
C2164 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.PDM 0.02104f
C2165 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PDM 0.0404f
C2166 XThC.Tn[7] XThR.Tn[11] 0.29362f
C2167 XA.XIR[11].XIC[3].icell.PDM Vbias 0.03922f
C2168 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PDM 0.04035f
C2169 XA.XIR[14].XIC[11].icell.Ien VPWR 0.19845f
C2170 XA.XIR[10].XIC[7].icell.PDM Vbias 0.03922f
C2171 XA.XIR[0].XIC[12].icell.Ien Iout 0.06775f
C2172 XThR.Tn[14] XA.XIR[14].XIC[5].icell.Ien 0.15202f
C2173 XThR.Tn[1] XA.XIR[1].XIC[5].icell.Ien 0.15202f
C2174 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PDM 0.02765f
C2175 XA.XIR[6].XIC[1].icell.Ien VPWR 0.1979f
C2176 XThR.XTBN.Y XThR.XTB3.Y 0.17246f
C2177 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PDM 0.04035f
C2178 XThC.Tn[10] XA.XIR[12].XIC[10].icell.Ien 0.03605f
C2179 XThR.Tn[13] XA.XIR[13].XIC[9].icell.Ien 0.15202f
C2180 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.PDM 0.02104f
C2181 XA.XIR[7].XIC_15.icell.Ien Iout 0.0694f
C2182 XThC.Tn[11] XThR.Tn[13] 0.29362f
C2183 XThR.Tn[2] VPWR 8.27233f
C2184 XA.XIR[5].XIC[7].icell.Ien Vbias 0.19161f
C2185 XA.XIR[5].XIC[0].icell.Ien Iout 0.06814f
C2186 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.PDM 0.02104f
C2187 XThC.Tn[1] XThR.Tn[1] 0.29362f
C2188 XThR.XTB1.Y XThR.XTB6.Y 0.05751f
C2189 XA.XIR[4].XIC_dummy_left.icell.Iout Iout 0.0353f
C2190 XThR.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.15202f
C2191 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.PDM 0.02104f
C2192 XThC.Tn[14] Iout 0.84533f
C2193 XThC.Tn[14] XThR.Tn[9] 0.29368f
C2194 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PDM 0.02765f
C2195 XThC.Tn[1] XThR.Tn[12] 0.29362f
C2196 XThC.Tn[10] XThR.Tn[8] 0.29362f
C2197 XA.XIR[6].XIC[6].icell.Ien VPWR 0.1979f
C2198 XThR.XTB3.Y XThR.XTB4.Y 2.13136f
C2199 XA.XIR[12].XIC[2].icell.Ien Vbias 0.19161f
C2200 XA.XIR[0].XIC_15.icell.PDM Vbias 0.03947f
C2201 XA.XIR[6].XIC[2].icell.Ien Iout 0.06821f
C2202 XA.XIR[5].XIC[9].icell.PUM VPWR 0.01015f
C2203 XThC.XTB7.Y Vbias 0.01727f
C2204 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.PDM 0.02104f
C2205 XThC.XTBN.Y a_7651_9569# 0.23021f
C2206 XThR.XTB3.Y XThR.Tn[10] 0.29462f
C2207 XThC.Tn[5] XThR.Tn[4] 0.29362f
C2208 XA.XIR[7].XIC_dummy_right.icell.Iout Iout 0.01732f
C2209 XA.XIR[0].XIC_dummy_left.icell.Iout VPWR 0.11857f
C2210 XThC.XTB4.Y XThC.Tn[3] 0.18952f
C2211 XThC.Tn[0] XThR.Tn[10] 0.2936f
C2212 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14] 0.15202f
C2213 XThR.Tn[6] XA.XIR[6].XIC[14].icell.Ien 0.15202f
C2214 XA.XIR[13].XIC[2].icell.Ien VPWR 0.1979f
C2215 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.Ien 0.04854f
C2216 XThC.Tn[7] XA.XIR[14].XIC[7].icell.Ien 0.03605f
C2217 XThR.Tn[13] XThR.Tn[14] 0.19161f
C2218 XA.XIR[12].XIC[4].icell.PUM VPWR 0.01015f
C2219 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PDM 0.04035f
C2220 XA.XIR[11].XIC[5].icell.Ien VPWR 0.1979f
C2221 XThR.Tn[8] XA.XIR[8].XIC[1].icell.Ien 0.15202f
C2222 XA.XIR[10].XIC[7].icell.Ien VPWR 0.1979f
C2223 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.PDM 0.02104f
C2224 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2225 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.PDM 0.02104f
C2226 XThR.XTB7.Y XThR.Tn[7] 0.0835f
C2227 XA.XIR[10].XIC[3].icell.Ien Iout 0.06821f
C2228 XThC.XTB2.Y a_4067_9615# 0.02133f
C2229 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Iout 0.01728f
C2230 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PDM 0.02765f
C2231 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.PDM 0.02104f
C2232 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PDM 0.04035f
C2233 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2234 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.PDM 0.02104f
C2235 XThR.XTBN.Y VPWR 4.54375f
C2236 XA.XIR[3].XIC[12].icell.Ien Iout 0.06821f
C2237 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PDM 0.0404f
C2238 XA.XIR[2].XIC[9].icell.Ien VPWR 0.1979f
C2239 XThR.Tn[0] Vbias 1.46106f
C2240 XA.XIR[2].XIC[5].icell.Ien Iout 0.06821f
C2241 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.PDM 0.02104f
C2242 XA.XIR[1].XIC[11].icell.Ien VPWR 0.1979f
C2243 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.Ien 0.04854f
C2244 XThR.Tn[8] XA.XIR[8].XIC[6].icell.Ien 0.15202f
C2245 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PDM 0.04035f
C2246 XA.XIR[1].XIC[7].icell.Ien Iout 0.06821f
C2247 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.Ien 0.04854f
C2248 XThC.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.03605f
C2249 XA.XIR[6].XIC[6].icell.PDM Vbias 0.03922f
C2250 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PDM 0.02765f
C2251 XThC.Tn[7] XThR.Tn[14] 0.29362f
C2252 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.PDM 0.02104f
C2253 XA.XIR[14].XIC[3].icell.PDM Vbias 0.03922f
C2254 XThR.Tn[13] XA.XIR[13].XIC[14].icell.Ien 0.15202f
C2255 XA.XIR[5].XIC[13].icell.PDM Vbias 0.03922f
C2256 a_10051_9569# XThC.Tn[13] 0.19413f
C2257 XA.XIR[8].XIC_15.icell.Ien Iout 0.0694f
C2258 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PDM 0.02765f
C2259 XThR.XTB4.Y VPWR 0.92827f
C2260 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.PDM 0.02104f
C2261 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.Ien 0.04854f
C2262 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PDM 0.04056f
C2263 XA.XIR[13].XIC[7].icell.PDM Vbias 0.03922f
C2264 XA.XIR[11].XIC[1].icell.PUM VPWR 0.01015f
C2265 XThR.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.15202f
C2266 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PDM 0.04035f
C2267 XThR.Tn[10] XA.XIR[10].XIC_15.icell.Ien 0.13564f
C2268 XThR.Tn[10] VPWR 9.1748f
C2269 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Ien 0.01745f
C2270 XA.XIR[9].XIC[3].icell.Ien Vbias 0.19161f
C2271 XA.XIR[15].XIC[1].icell.PDM VPWR 0.01334f
C2272 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.Ien 0.04854f
C2273 XThC.Tn[9] VPWR 7.38691f
C2274 XThR.XTB5.A a_n1335_4229# 0.01243f
C2275 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PDM 0.02765f
C2276 XThR.Tn[1] XA.XIR[1].XIC[10].icell.Ien 0.15202f
C2277 XA.XIR[1].XIC[0].icell.PDM Vbias 0.03915f
C2278 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PDM 0.02765f
C2279 XA.XIR[8].XIC_dummy_right.icell.Iout Iout 0.01732f
C2280 XA.XIR[4].XIC[0].icell.PDM Vbias 0.03915f
C2281 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.Ien 0.04854f
C2282 XA.XIR[5].XIC[12].icell.Ien Vbias 0.19161f
C2283 XA.XIR[1].XIC_dummy_left.icell.Iout XA.XIR[2].XIC_dummy_left.icell.Iout 0.03665f
C2284 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.Ien 0.04854f
C2285 XA.XIR[9].XIC[5].icell.PUM VPWR 0.01015f
C2286 XA.XIR[3].XIC[8].icell.PDM Vbias 0.03922f
C2287 data[5] data[6] 0.01513f
C2288 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.Ien 0.04854f
C2289 XThC.XTB7.A XThC.XTB5.Y 0.11935f
C2290 XA.XIR[8].XIC[10].icell.PDM Vbias 0.03922f
C2291 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.PDM 0.02104f
C2292 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PDM 0.02765f
C2293 XA.XIR[2].XIC[14].icell.PDM Vbias 0.03922f
C2294 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.Ien 0.04854f
C2295 XThC.Tn[0] XA.XIR[14].XIC[0].icell.Ien 0.03605f
C2296 XA.XIR[6].XIC[11].icell.Ien VPWR 0.1979f
C2297 XThC.Tn[0] XThR.Tn[13] 0.29372f
C2298 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.PDM 0.02104f
C2299 XA.XIR[12].XIC[7].icell.Ien Vbias 0.19161f
C2300 XThC.Tn[8] XA.XIR[2].XIC[8].icell.Ien 0.03605f
C2301 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.Ien 0.04854f
C2302 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.Ien 0.04854f
C2303 XA.XIR[5].XIC[14].icell.PUM VPWR 0.01015f
C2304 XA.XIR[6].XIC[7].icell.Ien Iout 0.06821f
C2305 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PDM 0.04042f
C2306 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.Ien 0.04854f
C2307 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.Ien 0.04854f
C2308 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.PDM 0.02104f
C2309 XThC.Tn[3] Iout 0.84089f
C2310 XThC.Tn[3] XThR.Tn[9] 0.29362f
C2311 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout 0.06446f
C2312 XA.XIR[8].XIC[14].icell.PDM VPWR 0.01002f
C2313 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.Ien 0.04854f
C2314 XA.XIR[14].XIC[5].icell.Ien VPWR 0.19845f
C2315 XThC.Tn[1] XA.XIR[0].XIC[1].icell.Ien 0.0378f
C2316 XThR.Tn[13] XA.XIR[13].XIC[12].icell.Ien 0.15202f
C2317 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.02765f
C2318 XThC.XTB7.A XThC.XTBN.Y 0.59539f
C2319 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PDM 0.04035f
C2320 XA.XIR[13].XIC[7].icell.Ien VPWR 0.1979f
C2321 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PDM 0.04035f
C2322 XThR.XTB6.A XThR.XTBN.A 0.0512f
C2323 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2324 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.PDM 0.02104f
C2325 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2326 XThR.XTB7.Y a_n997_1579# 0.013f
C2327 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PDM 0.02765f
C2328 XA.XIR[13].XIC[3].icell.Ien Iout 0.06821f
C2329 XA.XIR[12].XIC[9].icell.PUM VPWR 0.01015f
C2330 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PDM 0.02765f
C2331 a_n997_1803# VPWR 0.01991f
C2332 XA.XIR[1].XIC[0].icell.Ien Vbias 0.1916f
C2333 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PDM 0.02765f
C2334 XA.XIR[11].XIC[6].icell.Ien Iout 0.06821f
C2335 XThC.Tn[10] XA.XIR[15].XIC[10].icell.Ien 0.03184f
C2336 XA.XIR[9].XIC_dummy_left.icell.Ien XThR.Tn[9] 0.01432f
C2337 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PDM 0.0404f
C2338 XA.XIR[4].XIC[0].icell.Ien Vbias 0.19149f
C2339 XThR.Tn[1] Vbias 1.4485f
C2340 XA.XIR[10].XIC[8].icell.Ien Iout 0.06821f
C2341 XA.XIR[8].XIC[0].icell.PUM VPWR 0.01015f
C2342 XThC.XTB7.A a_4861_9615# 0.02294f
C2343 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PDM 0.02765f
C2344 XThC.Tn[3] XThC.Tn[4] 0.49877f
C2345 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PDM 0.02765f
C2346 XThR.Tn[12] Vbias 1.44829f
C2347 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PDM 0.0404f
C2348 XA.XIR[2].XIC[14].icell.Ien VPWR 0.19796f
C2349 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.PDM 0.02104f
C2350 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.02765f
C2351 XThC.XTB5.A XThC.XTB5.Y 0.0538f
C2352 XA.XIR[2].XIC[10].icell.Ien Iout 0.06821f
C2353 XA.XIR[15].XIC[2].icell.Ien Vbias 0.15966f
C2354 XThR.Tn[8] XA.XIR[8].XIC[11].icell.Ien 0.15202f
C2355 XA.XIR[7].XIC[14].icell.PDM Vbias 0.03922f
C2356 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.Ien 0.04854f
C2357 XA.XIR[14].XIC[0].icell.Ien VPWR 0.19845f
C2358 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.Ien 0.04854f
C2359 XA.XIR[4].XIC[2].icell.PUM VPWR 0.01015f
C2360 XA.XIR[1].XIC[12].icell.Ien Iout 0.06821f
C2361 XA.XIR[4].XIC[5].icell.Ien Vbias 0.19161f
C2362 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.Ien 0.04854f
C2363 XThR.Tn[13] VPWR 9.25617f
C2364 XThC.Tn[11] XThR.Tn[7] 0.29362f
C2365 XThC.XTBN.Y a_5949_9615# 0.0768f
C2366 XThC.Tn[2] XA.XIR[5].XIC[2].icell.Ien 0.03605f
C2367 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.PDM 0.02104f
C2368 XThC.XTB7.B XThC.Tn[9] 0.09571f
C2369 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.PDM 0.02104f
C2370 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.PDM 0.02104f
C2371 XThC.XTB7.Y XThC.Tn[13] 0.11626f
C2372 XThR.Tn[5] XA.XIR[5].XIC[10].icell.Ien 0.15202f
C2373 XThC.Tn[8] Vbias 0.9946f
C2374 XA.XIR[9].XIC[10].icell.PDM Vbias 0.03922f
C2375 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.Ien 0.04854f
C2376 XA.XIR[15].XIC[4].icell.PUM VPWR 0.01015f
C2377 XA.XIR[0].XIC[2].icell.PDM Vbias 0.03943f
C2378 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PDM 0.02765f
C2379 XA.XIR[5].XIC[4].icell.Ien VPWR 0.1979f
C2380 XThC.Tn[1] XA.XIR[10].XIC[1].icell.Ien 0.03605f
C2381 XThR.Tn[13] XA.XIR[13].XIC[10].icell.Ien 0.15202f
C2382 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PDM 0.02765f
C2383 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.PDM 0.02104f
C2384 XA.XIR[9].XIC[8].icell.Ien Vbias 0.19161f
C2385 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.PDM 0.02104f
C2386 XA.XIR[4].XIC[7].icell.PUM VPWR 0.01015f
C2387 XThR.Tn[3] a_n1049_6699# 0.27008f
C2388 XThR.Tn[1] XA.XIR[1].XIC_15.icell.Ien 0.13564f
C2389 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.PDM 0.02104f
C2390 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.02765f
C2391 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.PDM 0.02104f
C2392 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.PDM 0.02104f
C2393 XA.XIR[1].XIC_15.icell.PDM Vbias 0.03927f
C2394 XA.XIR[9].XIC[14].icell.PDM VPWR 0.01002f
C2395 XThR.XTB6.A XThR.XTB6.Y 0.10153f
C2396 XA.XIR[7].XIC[1].icell.PUM VPWR 0.01015f
C2397 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.PDM 0.02104f
C2398 XThC.Tn[10] XThR.Tn[3] 0.29362f
C2399 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.Ien 0.04854f
C2400 XA.XIR[4].XIC_15.icell.PDM Vbias 0.03927f
C2401 XA.XIR[7].XIC[4].icell.Ien Vbias 0.19161f
C2402 XA.XIR[1].XIC_dummy_left.icell.Iout VPWR 0.11154f
C2403 XA.XIR[9].XIC[10].icell.PUM VPWR 0.01015f
C2404 XThC.Tn[7] VPWR 6.847f
C2405 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.Ien 0.04854f
C2406 XA.XIR[12].XIC[13].icell.Ien Iout 0.06821f
C2407 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PDM 0.04035f
C2408 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PDM 0.0404f
C2409 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PDM 0.04035f
C2410 XThC.Tn[13] XThR.Tn[0] 0.29454f
C2411 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.PDM 0.02104f
C2412 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.PDM 0.02104f
C2413 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2414 XA.XIR[7].XIC[6].icell.PUM VPWR 0.01015f
C2415 XA.XIR[6].XIC[12].icell.Ien Iout 0.06821f
C2416 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2417 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PDM 0.02765f
C2418 XThC.Tn[6] XA.XIR[10].XIC[6].icell.Ien 0.03605f
C2419 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.PDM 0.02104f
C2420 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout 0.06446f
C2421 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PDM 0.0283f
C2422 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Ien 0.01451f
C2423 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.Ien 0.04854f
C2424 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR 0.38999f
C2425 XA.XIR[14].XIC[6].icell.Ien Iout 0.06821f
C2426 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PDM 0.02765f
C2427 XThC.XTBN.A XThC.XTB7.Y 1.11562f
C2428 XA.XIR[5].XIC[0].icell.PDM Vbias 0.03915f
C2429 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.04035f
C2430 XA.XIR[13].XIC[8].icell.Ien Iout 0.06821f
C2431 XThR.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.15202f
C2432 XThC.Tn[9] XA.XIR[4].XIC[9].icell.Ien 0.03605f
C2433 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PDM 0.02765f
C2434 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.Ien 0.04854f
C2435 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.PDM 0.02104f
C2436 XA.XIR[5].XIC[0].icell.PUM VPWR 0.01015f
C2437 XThR.XTBN.A XThR.Tn[12] 0.22096f
C2438 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.PDM 0.02104f
C2439 XThC.Tn[5] XA.XIR[7].XIC[5].icell.Ien 0.03605f
C2440 a_3773_9615# VPWR 0.70508f
C2441 XA.XIR[11].XIC[5].icell.PDM Vbias 0.03922f
C2442 XThC.Tn[12] XThR.Tn[2] 0.29362f
C2443 XThR.XTB2.Y a_n997_3755# 0.06476f
C2444 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.Ien 0.04854f
C2445 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PDM 0.04035f
C2446 XA.XIR[10].XIC[9].icell.PDM Vbias 0.03922f
C2447 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.PDM 0.02104f
C2448 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.PDM 0.02104f
C2449 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout 0.06446f
C2450 XThR.XTBN.Y a_n1049_8581# 0.0607f
C2451 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.PDM 0.02104f
C2452 XThR.Tn[13] XA.XIR[13].XIC_15.icell.Ien 0.13564f
C2453 XThC.XTB4.Y a_5155_9615# 0.01546f
C2454 XA.XIR[6].XIC_dummy_left.icell.Iout VPWR 0.11115f
C2455 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PDM 0.04056f
C2456 XA.XIR[15].XIC[7].icell.Ien Vbias 0.15966f
C2457 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.Ien 0.04854f
C2458 XA.XIR[2].XIC_15.icell.Ien Iout 0.0694f
C2459 XA.XIR[12].XIC[11].icell.Ien Iout 0.06821f
C2460 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.PDM 0.02104f
C2461 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.Ien 0.04854f
C2462 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PDM 0.02765f
C2463 XA.XIR[4].XIC[10].icell.Ien Vbias 0.19161f
C2464 XThC.Tn[1] XA.XIR[13].XIC[1].icell.Ien 0.03605f
C2465 XA.XIR[0].XIC[1].icell.Ien Vbias 0.19209f
C2466 XA.XIR[2].XIC[1].icell.PDM Vbias 0.03922f
C2467 XThC.Tn[8] XThR.Tn[6] 0.29362f
C2468 XThC.Tn[7] XA.XIR[9].XIC[7].icell.Ien 0.03605f
C2469 XA.XIR[8].XIC[4].icell.Ien Vbias 0.19161f
C2470 XA.XIR[3].XIC[3].icell.PUM VPWR 0.01015f
C2471 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PDM 0.04035f
C2472 XThC.Tn[14] XA.XIR[0].XIC[14].icell.Ien 0.03731f
C2473 XThR.Tn[5] XA.XIR[5].XIC_15.icell.Ien 0.13564f
C2474 XThR.XTB3.Y a_n997_2891# 0.07285f
C2475 XA.XIR[15].XIC[9].icell.PUM VPWR 0.01015f
C2476 XThC.Tn[10] XThR.Tn[11] 0.29362f
C2477 XA.XIR[5].XIC[9].icell.Ien VPWR 0.1979f
C2478 XThC.XTBN.Y a_8739_9569# 0.22804f
C2479 XThC.Tn[0] XThR.Tn[7] 0.29363f
C2480 XA.XIR[9].XIC[13].icell.Ien Vbias 0.19161f
C2481 XA.XIR[5].XIC[5].icell.Ien Iout 0.06821f
C2482 XThC.XTB4.Y XThC.XTB6.Y 0.04273f
C2483 XA.XIR[2].XIC_dummy_right.icell.Iout Iout 0.01732f
C2484 XThC.Tn[2] XA.XIR[12].XIC[2].icell.Ien 0.03605f
C2485 XThR.Tn[4] XA.XIR[4].XIC[0].icell.Ien 0.15228f
C2486 XA.XIR[4].XIC[12].icell.PUM VPWR 0.01015f
C2487 XThC.XTB3.Y XThC.XTB7.Y 0.03772f
C2488 a_n1049_5317# XThR.Tn[6] 0.26047f
C2489 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10] 0.15202f
C2490 XThR.Tn[3] XA.XIR[3].XIC[0].icell.Ien 0.1525f
C2491 XA.XIR[0].XIC[6].icell.Ien Vbias 0.19212f
C2492 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout 0.06446f
C2493 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.PDM 0.02104f
C2494 XA.XIR[8].XIC[6].icell.PUM VPWR 0.01015f
C2495 XThC.XTB7.B XThC.Tn[7] 0.08407f
C2496 XThC.XTB5.Y XThC.Tn[11] 0.02206f
C2497 XA.XIR[12].XIC[4].icell.Ien VPWR 0.1979f
C2498 XThC.Tn[6] Vbias 0.92065f
C2499 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout 0.06446f
C2500 XThR.Tn[5] Iout 1.19572f
C2501 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.Ien 0.04854f
C2502 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.PDM 0.02104f
C2503 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PDM 0.04035f
C2504 XThR.Tn[8] data[4] 0.01643f
C2505 XThR.XTB7.Y XThR.Tn[8] 0.07806f
C2506 a_8739_9569# XThC.Tn[10] 0.19671f
C2507 a_n997_3979# VPWR 0.01662f
C2508 XA.XIR[7].XIC[9].icell.Ien Vbias 0.19161f
C2509 XThC.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.03605f
C2510 XA.XIR[9].XIC_15.icell.PUM VPWR 0.01655f
C2511 XThC.Tn[13] XThR.Tn[1] 0.29363f
C2512 XThR.Tn[8] XA.XIR[8].XIC_dummy_left.icell.Iout 0.04617f
C2513 XThR.XTBN.A data[7] 0.07741f
C2514 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2515 XThC.Tn[6] XA.XIR[13].XIC[6].icell.Ien 0.03605f
C2516 XThR.Tn[4] XA.XIR[4].XIC[5].icell.Ien 0.15202f
C2517 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.Ien 0.04854f
C2518 XThR.XTB6.Y XThR.Tn[12] 0.02431f
C2519 XThC.Tn[13] XThR.Tn[12] 0.29363f
C2520 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.Ien 0.04854f
C2521 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PDM 0.04035f
C2522 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.PDM 0.02104f
C2523 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PDM 0.04035f
C2524 XThC.XTB6.A XThC.XTBN.A 0.0513f
C2525 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PDM 0.02765f
C2526 XA.XIR[2].XIC[0].icell.Ien Vbias 0.19149f
C2527 XThC.XTBN.Y XThC.Tn[11] 0.53369f
C2528 XThC.Tn[8] XThR.Tn[4] 0.29362f
C2529 XThC.Tn[5] XA.XIR[8].XIC[5].icell.Ien 0.03605f
C2530 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PDM 0.04035f
C2531 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR 0.38939f
C2532 XA.XIR[7].XIC[11].icell.PUM VPWR 0.01015f
C2533 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PDM 0.02765f
C2534 XA.XIR[7].XIC[1].icell.PDM Vbias 0.03922f
C2535 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.04035f
C2536 XA.XIR[10].XIC[1].icell.Ien Vbias 0.19161f
C2537 XThC.Tn[12] XThR.Tn[10] 0.29362f
C2538 XThC.Tn[2] XThR.Tn[0] 0.29628f
C2539 XA.XIR[6].XIC[8].icell.PDM Vbias 0.03922f
C2540 XThC.Tn[4] XThR.Tn[5] 0.29362f
C2541 XThR.Tn[12] XA.XIR[12].XIC[3].icell.Ien 0.15202f
C2542 XA.XIR[8].XIC[1].icell.PUM VPWR 0.01015f
C2543 XA.XIR[5].XIC_15.icell.PDM Vbias 0.03927f
C2544 XA.XIR[14].XIC[5].icell.PDM Vbias 0.03922f
C2545 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.Ien 0.04854f
C2546 XThR.Tn[3] XA.XIR[3].XIC[8].icell.Ien 0.15202f
C2547 XThC.Tn[10] XThC.Tn[11] 0.09949f
C2548 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PDM 0.02765f
C2549 XThR.Tn[7] VPWR 8.62165f
C2550 XA.XIR[13].XIC[9].icell.PDM Vbias 0.03922f
C2551 a_n997_2891# VPWR 0.01347f
C2552 XThC.XTB1.Y XThC.XTB7.Y 0.05222f
C2553 XThC.Tn[8] XA.XIR[5].XIC[8].icell.Ien 0.03605f
C2554 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PDM 0.04035f
C2555 XThC.XTB2.Y XThC.XTB6.Y 0.04959f
C2556 XThC.Tn[14] XA.XIR[3].XIC[14].icell.Ien 0.03605f
C2557 XThR.Tn[2] XA.XIR[2].XIC[3].icell.Ien 0.15202f
C2558 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout 0.06446f
C2559 XThR.XTB6.Y a_n1049_5317# 0.01199f
C2560 XA.XIR[15].XIC[3].icell.PDM VPWR 0.01334f
C2561 XA.XIR[4].XIC[2].icell.Ien VPWR 0.1979f
C2562 XA.XIR[3].XIC_dummy_right.icell.Iout XA.XIR[4].XIC_dummy_right.icell.Iout 0.04047f
C2563 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.Ien 0.04854f
C2564 XThC.Tn[0] XA.XIR[9].XIC[0].icell.Ien 0.03605f
C2565 XA.XIR[11].XIC[13].icell.Ien Vbias 0.19161f
C2566 XA.XIR[15].XIC[13].icell.Ien Iout 0.07211f
C2567 XThC.Tn[1] XA.XIR[6].XIC[1].icell.Ien 0.03605f
C2568 XA.XIR[3].XIC[6].icell.Ien Vbias 0.19161f
C2569 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.Ien 0.04854f
C2570 XA.XIR[1].XIC[2].icell.PDM Vbias 0.03922f
C2571 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PDM 0.02765f
C2572 XThC.Tn[1] XThR.Tn[2] 0.29362f
C2573 XA.XIR[4].XIC[2].icell.PDM Vbias 0.03922f
C2574 XA.XIR[9].XIC[5].icell.Ien VPWR 0.1979f
C2575 XThR.XTB5.A data[5] 0.11096f
C2576 XA.XIR[8].XIC[12].icell.PDM Vbias 0.03922f
C2577 XA.XIR[3].XIC[10].icell.PDM Vbias 0.03922f
C2578 XThC.Tn[10] XThR.Tn[14] 0.29362f
C2579 XA.XIR[4].XIC_15.icell.Ien Vbias 0.19195f
C2580 XThC.XTB2.Y XThC.XTB4.Y 0.04006f
C2581 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PDM 0.02765f
C2582 XThR.XTBN.Y a_n1049_7787# 0.08456f
C2583 XThC.XTB6.A XThC.XTB3.Y 0.03869f
C2584 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.Ien 0.04854f
C2585 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PDM 0.0404f
C2586 XA.XIR[8].XIC[9].icell.Ien Vbias 0.19161f
C2587 XThR.XTB2.Y XThR.XTB7.Y 0.0437f
C2588 XA.XIR[3].XIC[8].icell.PUM VPWR 0.01015f
C2589 XA.XIR[5].XIC_dummy_left.icell.Iout XA.XIR[6].XIC_dummy_left.icell.Iout 0.03665f
C2590 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PDM 0.02765f
C2591 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11] 0.15202f
C2592 a_5155_9615# XThC.Tn[4] 0.26653f
C2593 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2594 a_n1049_6405# XThR.Tn[4] 0.26564f
C2595 XA.XIR[5].XIC[14].icell.Ien VPWR 0.19796f
C2596 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PDM 0.04035f
C2597 XA.XIR[11].XIC_dummy_left.icell.Iout Iout 0.0353f
C2598 XA.XIR[5].XIC[10].icell.Ien Iout 0.06821f
C2599 XA.XIR[1].XIC[3].icell.PUM VPWR 0.01015f
C2600 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2601 XA.XIR[3].XIC[14].icell.PDM VPWR 0.01002f
C2602 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.PDM 0.02104f
C2603 XThC.Tn[6] XThR.Tn[6] 0.29362f
C2604 XThC.XTBN.A XThC.Tn[8] 0.1369f
C2605 XA.XIR[12].XIC_15.icell.PUM VPWR 0.01655f
C2606 XA.XIR[0].XIC[11].icell.Ien Vbias 0.19209f
C2607 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PDM 0.04035f
C2608 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PDM 0.04035f
C2609 XA.XIR[8].XIC[11].icell.PUM VPWR 0.01015f
C2610 XA.XIR[12].XIC[9].icell.Ien VPWR 0.1979f
C2611 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.Ien 0.04854f
C2612 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2613 XA.XIR[12].XIC[5].icell.Ien Iout 0.06821f
C2614 XA.XIR[7].XIC[14].icell.Ien Vbias 0.19161f
C2615 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PDM 0.02765f
C2616 XA.XIR[9].XIC[0].icell.Ien VPWR 0.1979f
C2617 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Iout 0.01828f
C2618 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PDM 0.02765f
C2619 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PDM 0.04035f
C2620 XA.XIR[11].XIC[11].icell.Ien Vbias 0.19161f
C2621 XThR.Tn[4] XA.XIR[4].XIC[10].icell.Ien 0.15202f
C2622 XA.XIR[15].XIC[11].icell.Ien Iout 0.07211f
C2623 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PDM 0.02765f
C2624 XThR.Tn[0] XA.XIR[0].XIC[2].icell.Ien 0.15202f
C2625 XA.XIR[13].XIC[1].icell.Ien Vbias 0.19161f
C2626 XThC.XTB7.A a_5949_9615# 0.01824f
C2627 XThC.Tn[11] XA.XIR[7].XIC[11].icell.Ien 0.03605f
C2628 XThC.Tn[12] XThR.Tn[13] 0.29362f
C2629 XThC.Tn[2] XThR.Tn[1] 0.29434f
C2630 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PDM 0.04035f
C2631 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.Ien 0.04854f
C2632 XThR.Tn[7] XA.XIR[7].XIC[3].icell.Ien 0.15202f
C2633 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PDM 0.02765f
C2634 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2635 XThC.XTB2.Y a_7875_9569# 0.06476f
C2636 XA.XIR[5].XIC[1].icell.PUM VPWR 0.01015f
C2637 XThC.XTB1.Y XThC.XTB6.A 0.01609f
C2638 XThC.Tn[2] XThR.Tn[12] 0.29362f
C2639 XThC.XTB5.A XThC.XTB7.A 0.07824f
C2640 XThC.Tn[11] XThR.Tn[8] 0.29362f
C2641 a_n997_1579# VPWR 0.02417f
C2642 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout 0.06446f
C2643 XThC.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.03605f
C2644 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.PDM 0.02104f
C2645 XThR.Tn[12] XA.XIR[12].XIC[8].icell.Ien 0.15202f
C2646 XThC.XTBN.Y XThC.Tn[0] 0.52915f
C2647 XA.XIR[7].XIC_dummy_left.icell.Iout XA.XIR[8].XIC_dummy_left.icell.Iout 0.03665f
C2648 XThC.Tn[2] XA.XIR[15].XIC[2].icell.Ien 0.03184f
C2649 XThR.Tn[3] XA.XIR[3].XIC[13].icell.Ien 0.15202f
C2650 XThC.Tn[6] XThR.Tn[4] 0.29362f
C2651 XA.XIR[14].XIC[13].icell.Ien Vbias 0.19161f
C2652 XA.XIR[6].XIC[3].icell.PUM VPWR 0.01015f
C2653 XA.XIR[9].XIC[12].icell.PDM Vbias 0.03922f
C2654 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.Ien 0.04854f
C2655 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.Ien 0.04854f
C2656 XThC.Tn[13] XA.XIR[9].XIC[13].icell.Ien 0.03605f
C2657 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout 0.06446f
C2658 XA.XIR[15].XIC[4].icell.Ien VPWR 0.33655f
C2659 XA.XIR[0].XIC[4].icell.PDM Vbias 0.03932f
C2660 XThC.Tn[1] XThR.Tn[10] 0.29362f
C2661 XThC.Tn[3] XA.XIR[11].XIC[3].icell.Ien 0.03605f
C2662 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PDM 0.02765f
C2663 XThR.Tn[2] XA.XIR[2].XIC[8].icell.Ien 0.15202f
C2664 XA.XIR[12].XIC[13].icell.PUM VPWR 0.01015f
C2665 XA.XIR[1].XIC[1].icell.Ien Vbias 0.19173f
C2666 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PDM 0.02765f
C2667 XA.XIR[4].XIC[7].icell.Ien VPWR 0.1979f
C2668 XA.XIR[10].XIC[2].icell.Ien Vbias 0.19161f
C2669 XA.XIR[9].XIC[1].icell.Ien Iout 0.06821f
C2670 XThR.Tn[9] XA.XIR[9].XIC[1].icell.Ien 0.15202f
C2671 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PDM 0.02827f
C2672 XThR.XTB7.Y a_n997_715# 0.06874f
C2673 XA.XIR[4].XIC[3].icell.Ien Iout 0.06821f
C2674 XThC.Tn[14] XA.XIR[1].XIC[14].icell.Ien 0.0361f
C2675 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PDM 0.02765f
C2676 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PDM 0.02765f
C2677 XThC.Tn[8] XA.XIR[12].XIC[8].icell.Ien 0.03605f
C2678 XA.XIR[3].XIC[11].icell.Ien Vbias 0.19161f
C2679 XA.XIR[3].XIC_dummy_left.icell.Iout XA.XIR[4].XIC_dummy_left.icell.Iout 0.03665f
C2680 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2681 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13] 0.15202f
C2682 XA.XIR[7].XIC[1].icell.Ien VPWR 0.1979f
C2683 XA.XIR[0].XIC[8].icell.PDM VPWR 0.01287f
C2684 XA.XIR[2].XIC[4].icell.Ien Vbias 0.19161f
C2685 XThC.XTB5.Y VPWR 1.01191f
C2686 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PDM 0.02765f
C2687 XA.XIR[9].XIC[10].icell.Ien VPWR 0.1979f
C2688 XA.XIR[10].XIC[4].icell.PUM VPWR 0.01015f
C2689 XA.XIR[1].XIC[6].icell.Ien Vbias 0.19173f
C2690 XA.XIR[12].XIC[14].icell.Ien VPWR 0.19796f
C2691 XA.XIR[9].XIC[6].icell.Ien Iout 0.06821f
C2692 XA.XIR[14].XIC_dummy_left.icell.Iout Iout 0.0353f
C2693 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.Ien 0.04854f
C2694 XThR.Tn[9] XA.XIR[9].XIC[6].icell.Ien 0.15202f
C2695 XA.XIR[0].XIC[3].icell.Ien VPWR 0.19726f
C2696 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PDM 0.04035f
C2697 XA.XIR[8].XIC[14].icell.Ien Vbias 0.19161f
C2698 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PDM 0.04035f
C2699 XA.XIR[3].XIC[13].icell.PUM VPWR 0.01015f
C2700 XA.XIR[7].XIC[6].icell.Ien VPWR 0.1979f
C2701 XA.XIR[2].XIC[6].icell.PUM VPWR 0.01015f
C2702 XA.XIR[5].XIC_15.icell.Ien Iout 0.0694f
C2703 XThC.XTBN.Y VPWR 4.08851f
C2704 XA.XIR[7].XIC[2].icell.Ien Iout 0.06821f
C2705 XA.XIR[1].XIC[8].icell.PUM VPWR 0.01015f
C2706 XThC.XTB6.Y a_6243_9615# 0.01199f
C2707 XThC.Tn[11] XA.XIR[8].XIC[11].icell.Ien 0.03605f
C2708 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.PDM 0.02104f
C2709 a_n1049_6699# VPWR 0.72162f
C2710 XThR.XTB7.A XThR.XTBN.A 0.19736f
C2711 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.PDM 0.02104f
C2712 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PDM 0.02765f
C2713 XA.XIR[14].XIC[11].icell.Ien Vbias 0.19161f
C2714 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2715 XA.XIR[5].XIC[2].icell.PDM Vbias 0.03922f
C2716 XThR.XTB7.A XThR.Tn[6] 0.1056f
C2717 XThC.XTB1.Y XThC.Tn[8] 0.29191f
C2718 XA.XIR[6].XIC[1].icell.Ien Vbias 0.19161f
C2719 XA.XIR[12].XIC[11].icell.PUM VPWR 0.01015f
C2720 XThR.Tn[11] XA.XIR[11].XIC[2].icell.Ien 0.15202f
C2721 XThC.Tn[10] VPWR 7.39238f
C2722 XA.XIR[12].XIC[1].icell.PDM Vbias 0.03922f
C2723 XThC.Tn[14] XA.XIR[6].XIC[14].icell.Ien 0.03605f
C2724 XThR.Tn[2] Vbias 1.44825f
C2725 XThC.Tn[5] XA.XIR[2].XIC[5].icell.Ien 0.03605f
C2726 XThR.Tn[4] XA.XIR[4].XIC_15.icell.Ien 0.13564f
C2727 a_4861_9615# VPWR 0.70525f
C2728 XThC.Tn[13] XA.XIR[11].XIC[13].icell.Ien 0.03605f
C2729 XThR.Tn[9] Iout 1.19574f
C2730 XA.XIR[11].XIC[7].icell.PDM Vbias 0.03922f
C2731 XA.XIR[5].XIC_dummy_right.icell.Iout Iout 0.01732f
C2732 XThR.Tn[0] XA.XIR[0].XIC[7].icell.Ien 0.15202f
C2733 XThR.Tn[10] XA.XIR[10].XIC[6].icell.Ien 0.15202f
C2734 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PDM 0.04035f
C2735 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2736 XThC.Tn[10] XA.XIR[13].XIC[10].icell.Ien 0.03605f
C2737 XThR.Tn[7] XA.XIR[7].XIC[8].icell.Ien 0.15202f
C2738 XA.XIR[6].XIC[6].icell.Ien Vbias 0.19161f
C2739 XThC.XTB5.Y a_9827_9569# 0.06458f
C2740 XA.XIR[12].XIC[12].icell.Ien VPWR 0.1979f
C2741 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.PDM 0.02104f
C2742 XA.XIR[15].XIC[0].icell.Ien Iout 0.07204f
C2743 XThC.Tn[3] XA.XIR[14].XIC[3].icell.Ien 0.03605f
C2744 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PDM 0.02765f
C2745 XThC.Tn[1] XThR.Tn[13] 0.29362f
C2746 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.Ien 0.04854f
C2747 XA.XIR[2].XIC[3].icell.PDM Vbias 0.03922f
C2748 XA.XIR[8].XIC[1].icell.Ien VPWR 0.1979f
C2749 XA.XIR[13].XIC[2].icell.Ien Vbias 0.19161f
C2750 XA.XIR[15].XIC_15.icell.PUM VPWR 0.01655f
C2751 XA.XIR[3].XIC[3].icell.Ien VPWR 0.1979f
C2752 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PDM 0.04035f
C2753 XThC.Tn[4] Iout 0.84166f
C2754 XThC.Tn[4] XThR.Tn[9] 0.29362f
C2755 XA.XIR[6].XIC[8].icell.PUM VPWR 0.01015f
C2756 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PDM 0.02765f
C2757 XThC.Tn[0] XThR.Tn[8] 0.29364f
C2758 XThC.Tn[0] XA.XIR[3].XIC[0].icell.Ien 0.03605f
C2759 XThR.XTB7.A XThR.Tn[4] 0.02736f
C2760 XA.XIR[15].XIC[9].icell.Ien VPWR 0.33655f
C2761 XA.XIR[11].XIC[5].icell.Ien Vbias 0.19161f
C2762 XThR.Tn[2] XA.XIR[2].XIC[13].icell.Ien 0.15202f
C2763 XThC.XTBN.Y a_9827_9569# 0.22873f
C2764 XThR.XTB7.A a_n1049_7493# 0.0127f
C2765 XA.XIR[15].XIC[5].icell.Ien Iout 0.07211f
C2766 XA.XIR[4].XIC[12].icell.Ien VPWR 0.1979f
C2767 XThC.XTB5.Y XThC.XTB7.B 0.30234f
C2768 XA.XIR[10].XIC[7].icell.Ien Vbias 0.19161f
C2769 data[1] data[2] 0.01393f
C2770 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14] 0.15202f
C2771 XA.XIR[4].XIC[8].icell.Ien Iout 0.06821f
C2772 XA.XIR[13].XIC[4].icell.PUM VPWR 0.01015f
C2773 XA.XIR[8].XIC[6].icell.Ien VPWR 0.1979f
C2774 XThR.XTB7.A XThR.XTB6.Y 0.19112f
C2775 XA.XIR[8].XIC[2].icell.Ien Iout 0.06821f
C2776 XA.XIR[11].XIC[7].icell.PUM VPWR 0.01015f
C2777 XA.XIR[2].XIC[9].icell.Ien Vbias 0.19161f
C2778 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PDM 0.04035f
C2779 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.Ien 0.04854f
C2780 XA.XIR[9].XIC_15.icell.Ien VPWR 0.26829f
C2781 XA.XIR[10].XIC[9].icell.PUM VPWR 0.01015f
C2782 XA.XIR[1].XIC[11].icell.Ien Vbias 0.19173f
C2783 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.PDM 0.02104f
C2784 XThR.XTB7.B XThR.XTBN.A 0.35142f
C2785 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.PDM 0.02104f
C2786 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2787 XThR.XTB7.Y XThR.Tn[11] 0.07412f
C2788 XA.XIR[9].XIC[11].icell.Ien Iout 0.06821f
C2789 XThR.Tn[9] XA.XIR[9].XIC[11].icell.Ien 0.15202f
C2790 XThC.XTB7.B XThC.XTBN.Y 0.38751f
C2791 XA.XIR[0].XIC[8].icell.Ien VPWR 0.19909f
C2792 XThR.XTB7.B XThR.Tn[6] 0.04822f
C2793 XA.XIR[0].XIC[4].icell.Ien Iout 0.06775f
C2794 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.PDM 0.02104f
C2795 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PDM 0.04035f
C2796 XA.XIR[12].XIC[10].icell.Ien VPWR 0.1979f
C2797 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PDM 0.04035f
C2798 XA.XIR[2].XIC[11].icell.PUM VPWR 0.01015f
C2799 XA.XIR[7].XIC[11].icell.Ien VPWR 0.1979f
C2800 XThC.Tn[12] XThR.Tn[7] 0.29362f
C2801 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.Ien 0.04854f
C2802 XA.XIR[7].XIC[7].icell.Ien Iout 0.06821f
C2803 XA.XIR[1].XIC[13].icell.PUM VPWR 0.01015f
C2804 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PDM 0.04035f
C2805 XA.XIR[7].XIC[3].icell.PDM Vbias 0.03922f
C2806 XThR.Tn[10] Vbias 1.4483f
C2807 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.Ien 0.04854f
C2808 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PDM 0.02765f
C2809 XThC.XTB7.B XThC.Tn[10] 0.14845f
C2810 XA.XIR[9].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2811 XA.XIR[6].XIC[10].icell.PDM Vbias 0.03922f
C2812 XA.XIR[15].XIC[1].icell.PDM Vbias 0.03922f
C2813 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.Ien 0.04854f
C2814 XThC.XTB7.Y XThC.Tn[14] 0.4237f
C2815 XA.XIR[15].XIC[13].icell.PUM VPWR 0.01015f
C2816 XThR.Tn[6] XA.XIR[6].XIC[1].icell.Ien 0.15202f
C2817 XThC.Tn[9] Vbias 0.99569f
C2818 XThR.Tn[8] VPWR 9.15728f
C2819 XA.XIR[3].XIC[0].icell.Ien VPWR 0.1979f
C2820 XThC.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.03605f
C2821 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.PDM 0.02104f
C2822 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PDM 0.02765f
C2823 XA.XIR[14].XIC[7].icell.PDM Vbias 0.03922f
C2824 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.PDM 0.02104f
C2825 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2826 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.PDM 0.02104f
C2827 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PDM 0.02765f
C2828 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.Ien 0.04854f
C2829 XA.XIR[11].XIC[1].icell.Ien VPWR 0.1979f
C2830 XThC.Tn[8] XA.XIR[15].XIC[8].icell.Ien 0.03184f
C2831 XThR.Tn[11] XA.XIR[11].XIC[7].icell.Ien 0.15202f
C2832 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PDM 0.04035f
C2833 XThC.XTB7.A data[1] 0.06544f
C2834 XThC.Tn[4] XA.XIR[0].XIC[4].icell.Ien 0.03708f
C2835 a_3773_9615# XThC.Tn[1] 0.27139f
C2836 XThR.XTB2.Y XThR.XTB3.Y 2.04808f
C2837 XThR.Tn[14] a_n997_715# 0.1927f
C2838 XThR.Tn[0] XA.XIR[0].XIC[12].icell.Ien 0.15202f
C2839 XA.XIR[15].XIC[5].icell.PDM VPWR 0.01334f
C2840 XA.XIR[6].XIC[14].icell.PDM VPWR 0.01002f
C2841 XThR.Tn[11] a_n997_2667# 0.19413f
C2842 XThC.Tn[9] XA.XIR[11].XIC[9].icell.Ien 0.03605f
C2843 XThR.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.15202f
C2844 XA.XIR[9].XIC_dummy_right.icell.Iout XA.XIR[10].XIC_dummy_right.icell.Iout 0.04047f
C2845 XThC.Tn[11] XThR.Tn[3] 0.29362f
C2846 XA.XIR[15].XIC[14].icell.Ien VPWR 0.33661f
C2847 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Ien 0.01757f
C2848 XA.XIR[1].XIC[4].icell.PDM Vbias 0.03922f
C2849 XA.XIR[6].XIC[11].icell.Ien Vbias 0.19161f
C2850 XThR.Tn[7] XA.XIR[7].XIC[13].icell.Ien 0.15202f
C2851 XA.XIR[4].XIC[4].icell.PDM Vbias 0.03922f
C2852 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.Ien 0.04854f
C2853 XThC.Tn[6] XA.XIR[4].XIC[6].icell.Ien 0.03605f
C2854 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.Ien 0.04854f
C2855 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PDM 0.02791f
C2856 XThC.XTB4.Y a_8963_9569# 0.07199f
C2857 XA.XIR[3].XIC[12].icell.PDM Vbias 0.03922f
C2858 XThC.Tn[14] XThR.Tn[0] 0.29421f
C2859 XA.XIR[8].XIC[14].icell.PDM Vbias 0.03922f
C2860 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.PDM 0.02104f
C2861 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.PDM 0.02104f
C2862 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.Ien 0.04854f
C2863 XA.XIR[14].XIC[5].icell.Ien Vbias 0.19161f
C2864 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.PDM 0.02104f
C2865 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PDM 0.02765f
C2866 XA.XIR[13].XIC[7].icell.Ien Vbias 0.19161f
C2867 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PDM 0.04035f
C2868 XThR.XTB7.B XThR.XTB6.Y 0.30244f
C2869 XA.XIR[3].XIC[8].icell.Ien VPWR 0.1979f
C2870 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.Ien 0.04854f
C2871 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.PDM 0.02104f
C2872 XA.XIR[6].XIC[13].icell.PUM VPWR 0.01015f
C2873 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.Ien 0.04854f
C2874 XA.XIR[3].XIC[4].icell.Ien Iout 0.06821f
C2875 XA.XIR[10].XIC[13].icell.Ien Iout 0.06821f
C2876 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout 0.06446f
C2877 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PDM 0.04035f
C2878 XThR.XTBN.Y XThR.XTBN.A 0.77119f
C2879 XA.XIR[15].XIC[11].icell.PUM VPWR 0.01015f
C2880 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PDM 0.02765f
C2881 XA.XIR[1].XIC[3].icell.Ien VPWR 0.1979f
C2882 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2883 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.PDM 0.02104f
C2884 XThC.XTB7.Y a_6243_10571# 0.01283f
C2885 XA.XIR[14].XIC[7].icell.PUM VPWR 0.01015f
C2886 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.Ien 0.04854f
C2887 a_n1049_7493# XThR.Tn[2] 0.26564f
C2888 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.Ien 0.04854f
C2889 XA.XIR[12].XIC_15.icell.Ien VPWR 0.26829f
C2890 XA.XIR[4].XIC[13].icell.Ien Iout 0.06821f
C2891 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.Ien 0.04854f
C2892 XThR.XTBN.Y XThR.Tn[6] 0.59899f
C2893 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PDM 0.04035f
C2894 XA.XIR[13].XIC[9].icell.PUM VPWR 0.01015f
C2895 XA.XIR[8].XIC[11].icell.Ien VPWR 0.1979f
C2896 XThR.XTB7.Y XThR.Tn[14] 0.4222f
C2897 XA.XIR[8].XIC[7].icell.Ien Iout 0.06821f
C2898 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.PDM 0.02104f
C2899 XThC.XTB5.A data[1] 0.11102f
C2900 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.Ien 0.04854f
C2901 XA.XIR[2].XIC[14].icell.Ien Vbias 0.19161f
C2902 XThC.Tn[13] XThR.Tn[2] 0.29363f
C2903 XThR.XTB2.Y VPWR 0.98845f
C2904 a_n997_3755# VPWR 0.0133f
C2905 XThR.XTB4.Y XThR.XTBN.A 0.03415f
C2906 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PDM 0.04035f
C2907 XA.XIR[14].XIC[0].icell.Ien Vbias 0.19149f
C2908 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PDM 0.02765f
C2909 XA.XIR[15].XIC[12].icell.Ien VPWR 0.33655f
C2910 XA.XIR[0].XIC[13].icell.Ien VPWR 0.19726f
C2911 XThC.Tn[4] XA.XIR[3].XIC[4].icell.Ien 0.03605f
C2912 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout 0.06446f
C2913 XThR.XTB5.Y XThR.Tn[5] 0.01094f
C2914 VPWR data[2] 0.21031f
C2915 XThR.XTBN.A XThR.Tn[10] 0.12147f
C2916 XThR.Tn[13] Vbias 1.4483f
C2917 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PDM 0.02765f
C2918 XThR.Tn[14] XA.XIR[14].XIC[2].icell.Ien 0.15202f
C2919 XThR.Tn[1] XA.XIR[1].XIC[2].icell.Ien 0.15202f
C2920 XA.XIR[0].XIC[9].icell.Ien Iout 0.06775f
C2921 XThC.Tn[11] XA.XIR[2].XIC[11].icell.Ien 0.03605f
C2922 XA.XIR[12].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2923 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PDM 0.02765f
C2924 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PDM 0.04035f
C2925 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PDM 0.02765f
C2926 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2927 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PDM 0.02765f
C2928 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.PDM 0.02104f
C2929 XThR.Tn[13] XA.XIR[13].XIC[6].icell.Ien 0.15202f
C2930 a_n1049_5611# VPWR 0.71817f
C2931 XA.XIR[7].XIC[12].icell.Ien Iout 0.06821f
C2932 XA.XIR[5].XIC[4].icell.Ien Vbias 0.19161f
C2933 XThC.Tn[9] XThR.Tn[6] 0.29362f
C2934 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.Ien 0.04854f
C2935 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.Ien 0.04854f
C2936 XA.XIR[14].XIC[1].icell.Ien VPWR 0.19845f
C2937 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.Ien 0.04854f
C2938 XA.XIR[10].XIC[11].icell.Ien Iout 0.06821f
C2939 XThC.Tn[11] XThR.Tn[11] 0.29362f
C2940 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.PDM 0.02104f
C2941 XA.XIR[3].XIC[1].icell.Ien Iout 0.06821f
C2942 XThR.XTBN.Y XThR.Tn[4] 0.60351f
C2943 XThC.Tn[9] XA.XIR[14].XIC[9].icell.Ien 0.03605f
C2944 XThC.Tn[1] XThR.Tn[7] 0.29362f
C2945 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.PDM 0.02104f
C2946 XA.XIR[6].XIC[3].icell.Ien VPWR 0.1979f
C2947 XA.XIR[9].XIC[14].icell.PDM Vbias 0.03922f
C2948 XThR.XTBN.Y a_n1049_7493# 0.08456f
C2949 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.Ien 0.04854f
C2950 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.PDM 0.02104f
C2951 XA.XIR[0].XIC[6].icell.PDM Vbias 0.03943f
C2952 XA.XIR[5].XIC[6].icell.PUM VPWR 0.01015f
C2953 XThC.XTB7.B a_7651_9569# 0.01152f
C2954 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.PDM 0.02104f
C2955 XThC.XTB5.Y XThC.Tn[12] 0.32495f
C2956 XA.XIR[9].XIC_dummy_left.icell.Iout Iout 0.0353f
C2957 XThR.Tn[9] XA.XIR[9].XIC_dummy_left.icell.Iout 0.04041f
C2958 XThC.Tn[7] Vbias 0.98016f
C2959 XThR.XTBN.Y XThR.XTB6.Y 0.1894f
C2960 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.PDM 0.02104f
C2961 XThR.Tn[6] XA.XIR[6].XIC[11].icell.Ien 0.15202f
C2962 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.PDM 0.02104f
C2963 XThC.Tn[2] XA.XIR[10].XIC[2].icell.Ien 0.03605f
C2964 XThC.Tn[14] XThR.Tn[1] 0.29381f
C2965 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout 0.06446f
C2966 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PDM 0.02765f
C2967 XA.XIR[2].XIC[1].icell.Ien VPWR 0.1979f
C2968 XA.XIR[7].XIC_dummy_left.icell.Iout VPWR 0.1106f
C2969 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.Ien 0.04854f
C2970 XThR.XTB3.Y XThR.Tn[3] 0.01287f
C2971 XA.XIR[11].XIC[2].icell.Ien VPWR 0.1979f
C2972 XA.XIR[15].XIC[10].icell.Ien VPWR 0.33655f
C2973 XThC.Tn[14] XThR.Tn[12] 0.29368f
C2974 XA.XIR[13].XIC[13].icell.Ien Iout 0.06821f
C2975 XA.XIR[10].XIC[4].icell.Ien VPWR 0.1979f
C2976 XThC.XTB7.A VPWR 0.87301f
C2977 XThC.Tn[0] XThR.Tn[3] 0.29373f
C2978 XThC.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.03605f
C2979 XThR.XTBN.A a_n997_1803# 0.09118f
C2980 XThC.XTBN.Y XThC.Tn[12] 0.56523f
C2981 XThR.XTB3.Y XThR.XTB7.Y 0.03772f
C2982 XThR.XTB4.Y XThR.XTB6.Y 0.04273f
C2983 XThR.XTB3.Y data[4] 0.03253f
C2984 XThC.Tn[9] XThR.Tn[4] 0.29362f
C2985 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PDM 0.02765f
C2986 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PDM 0.04035f
C2987 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PDM 0.04035f
C2988 XA.XIR[3].XIC[13].icell.Ien VPWR 0.1979f
C2989 XA.XIR[3].XIC[9].icell.Ien Iout 0.06821f
C2990 XThR.XTB6.Y XThR.Tn[10] 0.02461f
C2991 XThC.Tn[3] XThR.Tn[0] 0.29366f
C2992 XA.XIR[2].XIC[6].icell.Ien VPWR 0.1979f
C2993 XThC.Tn[13] XThR.Tn[10] 0.29363f
C2994 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.PDM 0.02104f
C2995 XThC.Tn[5] XThR.Tn[5] 0.29362f
C2996 a_n997_715# VPWR 0.02818f
C2997 XA.XIR[1].XIC[8].icell.Ien VPWR 0.1979f
C2998 XA.XIR[2].XIC[2].icell.Ien Iout 0.06821f
C2999 XThR.Tn[8] XA.XIR[8].XIC[3].icell.Ien 0.15202f
C3000 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3001 XThR.Tn[10] XA.XIR[10].XIC_dummy_left.icell.Iout 0.0404f
C3002 XA.XIR[1].XIC[4].icell.Ien Iout 0.06821f
C3003 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PDM 0.02765f
C3004 XA.XIR[5].XIC[4].icell.PDM Vbias 0.03922f
C3005 XA.XIR[8].XIC[12].icell.Ien Iout 0.06821f
C3006 XThC.XTB7.B data[2] 0.07481f
C3007 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.PDM 0.02104f
C3008 XA.XIR[15].XIC[0].icell.PUM VPWR 0.01015f
C3009 XThR.Tn[5] XA.XIR[5].XIC[2].icell.Ien 0.15202f
C3010 XA.XIR[12].XIC[3].icell.PDM Vbias 0.03922f
C3011 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PDM 0.02765f
C3012 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.PDM 0.02104f
C3013 XThC.Tn[3] XA.XIR[9].XIC[3].icell.Ien 0.03605f
C3014 XA.XIR[11].XIC[9].icell.PDM Vbias 0.03922f
C3015 a_5949_9615# VPWR 0.7053f
C3016 XThC.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.03605f
C3017 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.Ien 0.04854f
C3018 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PDM 0.04035f
C3019 XThC.Tn[10] XA.XIR[0].XIC[10].icell.Ien 0.03735f
C3020 XThR.Tn[14] XA.XIR[14].XIC[7].icell.Ien 0.15202f
C3021 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.PDM 0.02104f
C3022 XA.XIR[0].XIC[14].icell.Ien Iout 0.06775f
C3023 XThR.Tn[1] XA.XIR[1].XIC[7].icell.Ien 0.15202f
C3024 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.PDM 0.02104f
C3025 XThC.Tn[2] XThR.Tn[2] 0.29362f
C3026 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.PDM 0.02104f
C3027 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.PDM 0.02104f
C3028 XThC.Tn[4] XA.XIR[1].XIC[4].icell.Ien 0.03605f
C3029 XThC.Tn[11] XThR.Tn[14] 0.29362f
C3030 XThR.Tn[3] VPWR 8.28824f
C3031 XA.XIR[13].XIC[11].icell.Ien Iout 0.06821f
C3032 XThC.XTB5.A VPWR 0.82807f
C3033 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.PDM 0.02104f
C3034 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout 0.06446f
C3035 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.Ien 0.04854f
C3036 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.Ien 0.04854f
C3037 XA.XIR[5].XIC[9].icell.Ien Vbias 0.19161f
C3038 XA.XIR[12].XIC_dummy_right.icell.Iout XA.XIR[13].XIC_dummy_right.icell.Iout 0.04047f
C3039 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.Ien 0.04854f
C3040 XA.XIR[8].XIC[1].icell.PDM Vbias 0.03922f
C3041 VPWR data[4] 0.5303f
C3042 XThR.XTB7.Y VPWR 1.14768f
C3043 XThC.Tn[12] XA.XIR[4].XIC[12].icell.Ien 0.03605f
C3044 XA.XIR[2].XIC[5].icell.PDM Vbias 0.03922f
C3045 XThR.XTB5.A XThR.XTB5.Y 0.0538f
C3046 XA.XIR[8].XIC_dummy_left.icell.Iout VPWR 0.11107f
C3047 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.Ien 0.04854f
C3048 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.Ien 0.04854f
C3049 XA.XIR[15].XIC_15.icell.Ien VPWR 0.37868f
C3050 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PDM 0.04035f
C3051 XA.XIR[12].XIC[4].icell.Ien Vbias 0.19161f
C3052 XA.XIR[6].XIC[8].icell.Ien VPWR 0.1979f
C3053 XThC.Tn[0] XA.XIR[12].XIC[0].icell.Ien 0.03605f
C3054 XThC.XTBN.A XThC.Tn[9] 0.12399f
C3055 XA.XIR[6].XIC[4].icell.Ien Iout 0.06821f
C3056 XThC.Tn[7] XThR.Tn[6] 0.29362f
C3057 XA.XIR[5].XIC[11].icell.PUM VPWR 0.01015f
C3058 XThC.Tn[2] XA.XIR[13].XIC[2].icell.Ien 0.03605f
C3059 XThC.XTBN.Y a_10915_9569# 0.21503f
C3060 XThC.Tn[0] XThR.Tn[11] 0.2937f
C3061 XA.XIR[14].XIC[2].icell.Ien VPWR 0.19845f
C3062 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.Ien 0.04854f
C3063 XThC.XTB7.A XThC.XTB7.B 0.35844f
C3064 XA.XIR[13].XIC[4].icell.Ien VPWR 0.1979f
C3065 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.PDM 0.02104f
C3066 XA.XIR[12].XIC[6].icell.PUM VPWR 0.01015f
C3067 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PDM 0.02765f
C3068 XThC.Tn[1] XA.XIR[7].XIC[1].icell.Ien 0.03605f
C3069 XA.XIR[10].XIC_15.icell.PUM VPWR 0.01655f
C3070 XA.XIR[15].XIC_dummy_right.icell.Iout VPWR 0.21463f
C3071 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.PDM 0.02104f
C3072 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.Ien 0.04854f
C3073 XA.XIR[11].XIC[7].icell.Ien VPWR 0.1979f
C3074 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PDM 0.04035f
C3075 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.PDM 0.02104f
C3076 XThC.XTB6.Y XThC.Tn[5] 0.20189f
C3077 XThR.XTB6.Y XThR.Tn[13] 0.32265f
C3078 XA.XIR[11].XIC[3].icell.Ien Iout 0.06821f
C3079 XA.XIR[10].XIC[9].icell.Ien VPWR 0.1979f
C3080 XThC.Tn[13] XThR.Tn[13] 0.29363f
C3081 XThC.Tn[3] XThR.Tn[1] 0.29363f
C3082 XA.XIR[10].XIC[5].icell.Ien Iout 0.06821f
C3083 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.Ien 0.04854f
C3084 a_n997_2667# VPWR 0.01642f
C3085 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3086 XThC.Tn[4] XA.XIR[6].XIC[4].icell.Ien 0.03605f
C3087 XThR.XTB5.A XThR.XTB1.Y 0.1098f
C3088 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PDM 0.04035f
C3089 XThC.Tn[3] XThR.Tn[12] 0.29362f
C3090 XThC.Tn[10] XA.XIR[3].XIC[10].icell.Ien 0.03605f
C3091 XThC.Tn[12] XThR.Tn[8] 0.29362f
C3092 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR 0.38711f
C3093 XA.XIR[3].XIC[14].icell.Ien Iout 0.06821f
C3094 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PDM 0.04035f
C3095 XThR.Tn[7] Vbias 1.44824f
C3096 XA.XIR[2].XIC[11].icell.Ien VPWR 0.1979f
C3097 XThC.Tn[5] XA.XIR[12].XIC[5].icell.Ien 0.03605f
C3098 XThC.XTBN.Y XThC.Tn[1] 0.73206f
C3099 XA.XIR[2].XIC[7].icell.Ien Iout 0.06821f
C3100 XA.XIR[1].XIC[13].icell.Ien VPWR 0.1979f
C3101 XA.XIR[7].XIC[5].icell.PDM Vbias 0.03922f
C3102 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PDM 0.04035f
C3103 XThR.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.15202f
C3104 XThC.Tn[7] XThR.Tn[4] 0.29362f
C3105 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.Ien 0.04854f
C3106 XA.XIR[1].XIC[9].icell.Ien Iout 0.06821f
C3107 XA.XIR[6].XIC[12].icell.PDM Vbias 0.03922f
C3108 XA.XIR[15].XIC[3].icell.PDM Vbias 0.03922f
C3109 XA.XIR[4].XIC[2].icell.Ien Vbias 0.19161f
C3110 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Iout 0.04432f
C3111 VPWR bias[1] 1.33312f
C3112 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.Ien 0.04854f
C3113 XA.XIR[14].XIC[9].icell.PDM Vbias 0.03922f
C3114 XThC.Tn[2] XThR.Tn[10] 0.29362f
C3115 XA.XIR[12].XIC[0].icell.Ien VPWR 0.1979f
C3116 XThC.XTB6.Y a_10051_9569# 0.07626f
C3117 XThR.Tn[11] VPWR 9.22686f
C3118 XThR.Tn[5] XA.XIR[5].XIC[7].icell.Ien 0.15202f
C3119 XA.XIR[9].XIC[1].icell.PDM Vbias 0.03922f
C3120 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PDM 0.04035f
C3121 XA.XIR[9].XIC[2].icell.PUM VPWR 0.01015f
C3122 XThC.XTB5.A XThC.XTB7.B 0.30355f
C3123 XA.XIR[9].XIC[5].icell.Ien Vbias 0.19161f
C3124 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3125 XA.XIR[4].XIC[4].icell.PUM VPWR 0.01015f
C3126 XA.XIR[15].XIC[7].icell.PDM VPWR 0.01334f
C3127 XThR.Tn[1] XA.XIR[1].XIC[12].icell.Ien 0.15202f
C3128 XA.XIR[10].XIC[13].icell.PUM VPWR 0.01015f
C3129 XA.XIR[1].XIC[6].icell.PDM Vbias 0.03922f
C3130 XThR.XTB5.Y XThR.Tn[9] 0.01732f
C3131 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.Ien 0.04854f
C3132 XA.XIR[4].XIC[6].icell.PDM Vbias 0.03922f
C3133 XA.XIR[5].XIC[14].icell.Ien Vbias 0.19161f
C3134 XThC.Tn[8] XA.XIR[10].XIC[8].icell.Ien 0.03605f
C3135 XA.XIR[9].XIC[7].icell.PUM VPWR 0.01015f
C3136 XA.XIR[3].XIC[14].icell.PDM Vbias 0.03922f
C3137 XThR.XTBN.A a_n997_3979# 0.02087f
C3138 XThC.Tn[1] XA.XIR[8].XIC[1].icell.Ien 0.03605f
C3139 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.PDM 0.02104f
C3140 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.Ien 0.04854f
C3141 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.Ien 0.04854f
C3142 XThC.Tn[0] XThR.Tn[14] 0.29368f
C3143 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.04035f
C3144 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PDM 0.02765f
C3145 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.PDM 0.02104f
C3146 XThC.Tn[11] XA.XIR[5].XIC[11].icell.Ien 0.03605f
C3147 XA.XIR[12].XIC[9].icell.Ien Vbias 0.19161f
C3148 XA.XIR[6].XIC[13].icell.Ien VPWR 0.1979f
C3149 XA.XIR[10].XIC[14].icell.Ien VPWR 0.19796f
C3150 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3151 XA.XIR[6].XIC[9].icell.Ien Iout 0.06821f
C3152 XA.XIR[7].XIC[3].icell.PUM VPWR 0.01015f
C3153 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PDM 0.02765f
C3154 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PDM 0.04035f
C3155 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PDM 0.02765f
C3156 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PDM 0.02765f
C3157 XA.XIR[9].XIC[0].icell.Ien Vbias 0.19149f
C3158 XA.XIR[13].XIC_15.icell.PUM VPWR 0.01655f
C3159 XA.XIR[14].XIC[7].icell.Ien VPWR 0.19845f
C3160 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3161 XA.XIR[14].XIC[3].icell.Ien Iout 0.06821f
C3162 XA.XIR[13].XIC[9].icell.Ien VPWR 0.1979f
C3163 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PDM 0.04035f
C3164 XThC.Tn[12] XA.XIR[15].XIC[12].icell.Ien 0.03184f
C3165 XThC.Tn[11] VPWR 7.42185f
C3166 XA.XIR[13].XIC[5].icell.Ien Iout 0.06821f
C3167 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.Ien 0.04854f
C3168 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR 0.01604f
C3169 XThC.XTBN.A XThC.Tn[7] 0.01439f
C3170 XThR.Tn[12] XA.XIR[12].XIC[13].icell.Ien 0.15202f
C3171 XThR.Tn[13] XA.XIR[13].XIC_dummy_left.icell.Iout 0.0404f
C3172 XA.XIR[11].XIC[8].icell.Ien Iout 0.06821f
C3173 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PDM 0.04035f
C3174 XThR.XTBN.A XThR.Tn[7] 0.01439f
C3175 XThR.XTBN.A a_n997_2891# 0.01719f
C3176 XA.XIR[10].XIC[11].icell.PUM VPWR 0.01015f
C3177 XThR.Tn[6] XThR.Tn[7] 0.10214f
C3178 XA.XIR[10].XIC[0].icell.PDM Vbias 0.03915f
C3179 XThC.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.03605f
C3180 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PDM 0.04056f
C3181 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PDM 0.04035f
C3182 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.Ien 0.04854f
C3183 data[6] data[7] 0.04128f
C3184 XThC.Tn[2] XThR.Tn[13] 0.29362f
C3185 XA.XIR[15].XIC[1].icell.PUM VPWR 0.01015f
C3186 XA.XIR[5].XIC[1].icell.Ien VPWR 0.1979f
C3187 XA.XIR[2].XIC[12].icell.Ien Iout 0.06821f
C3188 XA.XIR[15].XIC[4].icell.Ien Vbias 0.15966f
C3189 XThR.Tn[8] XA.XIR[8].XIC[13].icell.Ien 0.15202f
C3190 XThR.Tn[14] VPWR 9.46534f
C3191 XThC.Tn[10] XA.XIR[1].XIC[10].icell.Ien 0.03605f
C3192 XA.XIR[1].XIC[14].icell.Ien Iout 0.06821f
C3193 XThC.Tn[5] Iout 0.84205f
C3194 XThC.Tn[5] XThR.Tn[9] 0.29362f
C3195 XA.XIR[4].XIC[7].icell.Ien Vbias 0.19161f
C3196 XThC.Tn[1] XThR.Tn[8] 0.29362f
C3197 XThR.XTB2.Y a_n1335_8107# 0.01006f
C3198 XA.XIR[10].XIC[12].icell.Ien VPWR 0.1979f
C3199 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.Ien 0.04854f
C3200 XA.XIR[3].XIC_dummy_left.icell.Iout Iout 0.0353f
C3201 bias[1] bias[0] 0.56718f
C3202 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PDM 0.02765f
C3203 XThC.Tn[1] XA.XIR[11].XIC[1].icell.Ien 0.03605f
C3204 XA.XIR[12].XIC[1].icell.Ien Iout 0.06821f
C3205 XThR.Tn[5] XA.XIR[5].XIC[12].icell.Ien 0.15202f
C3206 VPWR data[1] 0.44103f
C3207 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.Ien 0.04854f
C3208 XA.XIR[13].XIC[13].icell.PUM VPWR 0.01015f
C3209 XThC.XTB6.Y XThC.XTB7.Y 2.05133f
C3210 XA.XIR[7].XIC[1].icell.Ien Vbias 0.19161f
C3211 XA.XIR[0].XIC[8].icell.PDM Vbias 0.03943f
C3212 XA.XIR[15].XIC[6].icell.PUM VPWR 0.01015f
C3213 XA.XIR[5].XIC[6].icell.Ien VPWR 0.1979f
C3214 XThC.XTB5.Y Vbias 0.01575f
C3215 XThC.XTB7.B a_8739_9569# 0.0168f
C3216 XA.XIR[9].XIC[10].icell.Ien Vbias 0.19161f
C3217 XA.XIR[4].XIC[9].icell.PUM VPWR 0.01015f
C3218 XA.XIR[5].XIC[2].icell.Ien Iout 0.06821f
C3219 XThC.Tn[14] XA.XIR[7].XIC[14].icell.Ien 0.03605f
C3220 XA.XIR[12].XIC[14].icell.Ien Vbias 0.19161f
C3221 XThC.Tn[8] XA.XIR[13].XIC[8].icell.Ien 0.03605f
C3222 XA.XIR[0].XIC[3].icell.Ien Vbias 0.19206f
C3223 XA.XIR[8].XIC[3].icell.PUM VPWR 0.01015f
C3224 XThR.Tn[12] XA.XIR[12].XIC[11].icell.Ien 0.15202f
C3225 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR 0.3367f
C3226 XThC.Tn[4] XThC.Tn[5] 0.4169f
C3227 XThR.XTB2.Y a_n1049_7787# 0.2342f
C3228 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PDM 0.02765f
C3229 XA.XIR[2].XIC_dummy_left.icell.Iout VPWR 0.1106f
C3230 XA.XIR[0].XIC[12].icell.PDM VPWR 0.01293f
C3231 XA.XIR[7].XIC[6].icell.Ien Vbias 0.19161f
C3232 XA.XIR[13].XIC[14].icell.Ien VPWR 0.19796f
C3233 XA.XIR[9].XIC[12].icell.PUM VPWR 0.01015f
C3234 XThC.XTBN.Y Vbias 0.16301f
C3235 XThC.Tn[5] XA.XIR[15].XIC[5].icell.Ien 0.03184f
C3236 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PDM 0.02765f
C3237 XThR.Tn[4] XA.XIR[4].XIC[2].icell.Ien 0.15202f
C3238 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.Ien 0.04854f
C3239 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PDM 0.04035f
C3240 XThC.XTB4.Y XThC.XTB7.Y 0.03475f
C3241 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.Ien 0.04854f
C3242 XThR.XTB6.Y XThR.Tn[7] 0.01462f
C3243 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PDM 0.04035f
C3244 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.PDM 0.02104f
C3245 XThC.Tn[13] XThR.Tn[7] 0.29363f
C3246 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR 0.0824f
C3247 XThC.Tn[6] XA.XIR[11].XIC[6].icell.Ien 0.03605f
C3248 XThC.XTB7.B XThC.Tn[11] 0.03903f
C3249 XThC.Tn[10] XA.XIR[6].XIC[10].icell.Ien 0.03605f
C3250 XA.XIR[6].XIC[14].icell.Ien Iout 0.06821f
C3251 XA.XIR[7].XIC[8].icell.PUM VPWR 0.01015f
C3252 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.PDM 0.02104f
C3253 XThC.Tn[10] Vbias 1.05697f
C3254 XA.XIR[10].XIC[10].icell.Ien VPWR 0.1979f
C3255 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.PDM 0.02104f
C3256 XA.XIR[14].XIC[8].icell.Ien Iout 0.06821f
C3257 XA.XIR[5].XIC[6].icell.PDM Vbias 0.03922f
C3258 XA.XIR[13].XIC[11].icell.PUM VPWR 0.01015f
C3259 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PDM 0.0404f
C3260 XThR.Tn[3] XA.XIR[3].XIC[5].icell.Ien 0.15202f
C3261 a_3773_9615# XThC.Tn[2] 0.01175f
C3262 XA.XIR[13].XIC[0].icell.PDM Vbias 0.03915f
C3263 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.Ien 0.04854f
C3264 XThR.XTB3.Y VPWR 1.07975f
C3265 XA.XIR[12].XIC[5].icell.PDM Vbias 0.03922f
C3266 XA.XIR[12].XIC[12].icell.Ien Vbias 0.19161f
C3267 XThC.Tn[12] XThR.Tn[3] 0.29362f
C3268 XThR.XTB5.A XThR.XTB6.A 1.80461f
C3269 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3270 XThC.Tn[0] VPWR 6.52685f
C3271 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PDM 0.0404f
C3272 XA.XIR[8].XIC[1].icell.Ien Vbias 0.19161f
C3273 XA.XIR[3].XIC[3].icell.Ien Vbias 0.19161f
C3274 XThC.Tn[8] XThR.Tn[5] 0.29362f
C3275 XA.XIR[13].XIC[12].icell.Ien VPWR 0.1979f
C3276 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.02765f
C3277 XThC.Tn[14] XA.XIR[8].XIC[14].icell.Ien 0.03605f
C3278 XA.XIR[15].XIC[9].icell.Ien Vbias 0.15966f
C3279 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.PDM 0.02104f
C3280 XThC.Tn[1] XA.XIR[14].XIC[1].icell.Ien 0.03605f
C3281 XThC.XTB2.Y XThC.XTB7.Y 0.0437f
C3282 XThC.XTB6.A XThC.XTB6.Y 0.10153f
C3283 XA.XIR[9].XIC[2].icell.Ien VPWR 0.1979f
C3284 XA.XIR[4].XIC[12].icell.Ien Vbias 0.19161f
C3285 XA.XIR[3].XIC[1].icell.PDM Vbias 0.03922f
C3286 XA.XIR[8].XIC[3].icell.PDM Vbias 0.03922f
C3287 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.Ien 0.04854f
C3288 XA.XIR[2].XIC[7].icell.PDM Vbias 0.03922f
C3289 XThR.XTB6.A data[5] 0.37233f
C3290 XA.XIR[8].XIC[6].icell.Ien Vbias 0.19161f
C3291 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PDM 0.04035f
C3292 XA.XIR[3].XIC[5].icell.PUM VPWR 0.01015f
C3293 XA.XIR[5].XIC[11].icell.Ien VPWR 0.1979f
C3294 XA.XIR[9].XIC_15.icell.Ien Vbias 0.19195f
C3295 XA.XIR[5].XIC[7].icell.Ien Iout 0.06821f
C3296 XA.XIR[4].XIC[14].icell.PUM VPWR 0.01015f
C3297 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.PDM 0.02104f
C3298 XA.XIR[0].XIC[8].icell.Ien Vbias 0.19209f
C3299 XThC.Tn[14] XThR.Tn[2] 0.29368f
C3300 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.PDM 0.02104f
C3301 XA.XIR[8].XIC[8].icell.PUM VPWR 0.01015f
C3302 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PDM 0.04035f
C3303 XThC.XTB6.A XThC.XTB4.Y 0.04137f
C3304 XA.XIR[12].XIC[6].icell.Ien VPWR 0.1979f
C3305 XThC.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.03605f
C3306 XA.XIR[12].XIC[10].icell.Ien Vbias 0.19161f
C3307 XThR.XTB6.Y a_n997_1579# 0.07626f
C3308 XA.XIR[10].XIC_15.icell.Ien VPWR 0.26829f
C3309 XA.XIR[12].XIC[2].icell.Ien Iout 0.06821f
C3310 XA.XIR[7].XIC[11].icell.Ien Vbias 0.19161f
C3311 XThC.Tn[6] XA.XIR[14].XIC[6].icell.Ien 0.03605f
C3312 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.PDM 0.02104f
C3313 XThR.Tn[4] XA.XIR[4].XIC[7].icell.Ien 0.15202f
C3314 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.PDM 0.02104f
C3315 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.Ien 0.04854f
C3316 XA.XIR[13].XIC[10].icell.Ien VPWR 0.1979f
C3317 XA.XIR[3].XIC[0].icell.Ien Vbias 0.19149f
C3318 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PDM 0.04035f
C3319 XThR.Tn[8] Vbias 1.44824f
C3320 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PDM 0.04035f
C3321 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Iout 0.02485f
C3322 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.PDM 0.02104f
C3323 XThC.Tn[10] XThR.Tn[6] 0.29362f
C3324 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PDM 0.04035f
C3325 XA.XIR[7].XIC[13].icell.PUM VPWR 0.01015f
C3326 XA.XIR[11].XIC[1].icell.Ien Vbias 0.19161f
C3327 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.PDM 0.02104f
C3328 XThC.Tn[12] XThR.Tn[11] 0.29362f
C3329 XA.XIR[10].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3330 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.Ien 0.04854f
C3331 XA.XIR[7].XIC[7].icell.PDM Vbias 0.03922f
C3332 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PDM 0.0404f
C3333 XThC.Tn[2] XThR.Tn[7] 0.29362f
C3334 XA.XIR[15].XIC[5].icell.PDM Vbias 0.03922f
C3335 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PDM 0.04056f
C3336 XA.XIR[6].XIC[14].icell.PDM Vbias 0.03922f
C3337 XThR.Tn[12] XA.XIR[12].XIC[5].icell.Ien 0.15202f
C3338 XA.XIR[3].XIC[2].icell.PUM VPWR 0.01015f
C3339 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3340 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.PDM 0.02104f
C3341 XThR.Tn[3] XA.XIR[3].XIC[10].icell.Ien 0.15202f
C3342 XA.XIR[15].XIC[14].icell.Ien Vbias 0.15966f
C3343 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.PDM 0.02104f
C3344 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.Ien 0.04854f
C3345 XThC.XTB6.Y XThC.Tn[8] 0.02461f
C3346 XThC.Tn[2] XA.XIR[4].XIC[2].icell.Ien 0.03605f
C3347 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PDM 0.04056f
C3348 XA.XIR[9].XIC[3].icell.PDM Vbias 0.03922f
C3349 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.Ien 0.04854f
C3350 XThR.Tn[0] Iout 1.19579f
C3351 XThR.XTB7.Y a_n1319_5317# 0.01283f
C3352 XThR.Tn[2] XA.XIR[2].XIC[5].icell.Ien 0.15202f
C3353 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PDM 0.02765f
C3354 XA.XIR[15].XIC[9].icell.PDM VPWR 0.01334f
C3355 XA.XIR[4].XIC[4].icell.Ien VPWR 0.1979f
C3356 XThC.XTB2.Y XThC.XTB6.A 0.18237f
C3357 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PDM 0.02765f
C3358 XA.XIR[3].XIC[8].icell.Ien Vbias 0.19161f
C3359 XA.XIR[1].XIC[8].icell.PDM Vbias 0.03922f
C3360 XThC.Tn[1] XThR.Tn[3] 0.29362f
C3361 XThC.XTBN.Y XThC.Tn[13] 0.62331f
C3362 XThC.Tn[10] XThR.Tn[4] 0.29362f
C3363 XA.XIR[4].XIC[8].icell.PDM Vbias 0.03922f
C3364 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.Ien 0.04854f
C3365 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.Ien 0.04854f
C3366 XA.XIR[9].XIC[7].icell.Ien VPWR 0.1979f
C3367 XA.XIR[1].XIC[3].icell.Ien Vbias 0.19173f
C3368 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.Ien 0.04854f
C3369 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.PDM 0.02104f
C3370 XThC.XTB4.Y XThC.Tn[8] 0.01306f
C3371 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.PDM 0.02104f
C3372 XA.XIR[9].XIC[3].icell.Ien Iout 0.06821f
C3373 XThR.Tn[9] XA.XIR[9].XIC[3].icell.Ien 0.15202f
C3374 XA.XIR[12].XIC_15.icell.Ien Vbias 0.19195f
C3375 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.PDM 0.02104f
C3376 XThC.Tn[14] XThR.Tn[10] 0.29368f
C3377 XThC.Tn[4] XThR.Tn[0] 0.29364f
C3378 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PDM 0.02765f
C3379 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PDM 0.04035f
C3380 XThC.Tn[6] XThR.Tn[5] 0.29362f
C3381 XA.XIR[8].XIC[11].icell.Ien Vbias 0.19161f
C3382 XA.XIR[3].XIC[10].icell.PUM VPWR 0.01015f
C3383 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.PDM 0.02104f
C3384 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.Ien 0.04854f
C3385 XThC.Tn[7] XA.XIR[0].XIC[7].icell.Ien 0.03684f
C3386 XThC.Tn[11] XThC.Tn[12] 0.22144f
C3387 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.Ien 0.04854f
C3388 XA.XIR[2].XIC[3].icell.PUM VPWR 0.01015f
C3389 XA.XIR[7].XIC[3].icell.Ien VPWR 0.1979f
C3390 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PDM 0.04035f
C3391 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.Ien 0.04854f
C3392 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.Ien 0.04854f
C3393 XThC.XTB7.B VPWR 1.32988f
C3394 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.PDM 0.02104f
C3395 XA.XIR[5].XIC[12].icell.Ien Iout 0.06821f
C3396 XA.XIR[1].XIC[5].icell.PUM VPWR 0.01015f
C3397 XA.XIR[13].XIC_15.icell.Ien VPWR 0.26829f
C3398 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.Ien 0.04854f
C3399 XA.XIR[15].XIC[12].icell.Ien Vbias 0.15966f
C3400 XA.XIR[0].XIC[13].icell.Ien Vbias 0.19209f
C3401 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.Ien 0.04854f
C3402 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PDM 0.04035f
C3403 XA.XIR[8].XIC[13].icell.PUM VPWR 0.01015f
C3404 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PDM 0.04035f
C3405 XThC.XTBN.A XThC.XTB5.Y 0.10854f
C3406 XThC.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.03699f
C3407 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.PDM 0.02104f
C3408 XThR.Tn[7] XA.XIR[7].XIC[0].icell.Ien 0.15202f
C3409 XA.XIR[12].XIC[7].icell.Ien Iout 0.06821f
C3410 XThR.XTBN.A XThR.Tn[8] 0.1369f
C3411 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PDM 0.02765f
C3412 VPWR bias[0] 2.10172f
C3413 XThC.Tn[3] XThR.Tn[2] 0.29362f
C3414 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PDM 0.04035f
C3415 XThR.Tn[4] XA.XIR[4].XIC[12].icell.Ien 0.15202f
C3416 XA.XIR[14].XIC[1].icell.Ien Vbias 0.19161f
C3417 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.0404f
C3418 XThC.XTB7.Y a_6243_9615# 0.27822f
C3419 XThR.Tn[0] XA.XIR[0].XIC[4].icell.Ien 0.15202f
C3420 XA.XIR[0].XIC_15.icell.PUM VPWR 0.01577f
C3421 XThR.Tn[10] XA.XIR[10].XIC[3].icell.Ien 0.15202f
C3422 XThC.Tn[12] XThR.Tn[14] 0.29362f
C3423 XA.XIR[13].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3424 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PDM 0.0404f
C3425 XA.XIR[10].XIC[2].icell.PDM Vbias 0.03922f
C3426 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PDM 0.02765f
C3427 XThC.XTBN.A XThC.XTBN.Y 0.77125f
C3428 XThC.Tn[12] XA.XIR[10].XIC[12].icell.Ien 0.03605f
C3429 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PDM 0.04035f
C3430 XA.XIR[6].XIC[3].icell.Ien Vbias 0.19161f
C3431 XThR.XTB7.B data[6] 0.07481f
C3432 XThR.Tn[7] XA.XIR[7].XIC[5].icell.Ien 0.15202f
C3433 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.PDM 0.02104f
C3434 XA.XIR[15].XIC[1].icell.Ien VPWR 0.33655f
C3435 XA.XIR[5].XIC_dummy_left.icell.Iout VPWR 0.11117f
C3436 XThC.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.03605f
C3437 XA.XIR[1].XIC[0].icell.Ien Iout 0.06814f
C3438 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.Ien 0.04854f
C3439 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.Ien 0.04854f
C3440 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.Ien 0.04854f
C3441 XA.XIR[4].XIC[0].icell.Ien Iout 0.06814f
C3442 XThR.Tn[1] Iout 1.19576f
C3443 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PDM 0.02765f
C3444 XThR.Tn[3] XA.XIR[3].XIC_15.icell.Ien 0.13564f
C3445 XThC.XTBN.A XThC.Tn[10] 0.12148f
C3446 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.PDM 0.02104f
C3447 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PDM 0.02765f
C3448 XA.XIR[6].XIC[5].icell.PUM VPWR 0.01015f
C3449 XThC.Tn[1] XThR.Tn[11] 0.29362f
C3450 XThR.Tn[12] Iout 1.19574f
C3451 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout 0.06446f
C3452 XA.XIR[2].XIC[1].icell.Ien Vbias 0.19161f
C3453 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.Ien 0.04854f
C3454 XA.XIR[15].XIC[6].icell.Ien VPWR 0.33655f
C3455 XA.XIR[0].XIC[10].icell.PDM Vbias 0.03943f
C3456 XA.XIR[11].XIC[2].icell.Ien Vbias 0.19161f
C3457 XThC.Tn[7] XA.XIR[3].XIC[7].icell.Ien 0.03605f
C3458 XThR.Tn[2] XA.XIR[2].XIC[10].icell.Ien 0.15202f
C3459 XA.XIR[15].XIC[10].icell.Ien Vbias 0.15966f
C3460 XA.XIR[15].XIC[2].icell.Ien Iout 0.07211f
C3461 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PDM 0.02765f
C3462 XThC.XTB7.A Vbias 0.0149f
C3463 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.PDM 0.02104f
C3464 XA.XIR[10].XIC[4].icell.Ien Vbias 0.19161f
C3465 XThC.Tn[14] XA.XIR[2].XIC[14].icell.Ien 0.03605f
C3466 XThC.XTB3.Y XThC.XTB5.Y 0.04438f
C3467 XA.XIR[4].XIC[9].icell.Ien VPWR 0.1979f
C3468 XA.XIR[0].XIC[0].icell.Ien VPWR 0.19726f
C3469 XA.XIR[4].XIC[5].icell.Ien Iout 0.06821f
C3470 XThC.Tn[0] XA.XIR[10].XIC[0].icell.Ien 0.03605f
C3471 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.PDM 0.02104f
C3472 XA.XIR[8].XIC[3].icell.Ien VPWR 0.1979f
C3473 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.Ien 0.04854f
C3474 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.Ien 0.04854f
C3475 XA.XIR[3].XIC[13].icell.Ien Vbias 0.19161f
C3476 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.PDM 0.02104f
C3477 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PDM 0.02765f
C3478 XThC.Tn[14] XThR.Tn[13] 0.29368f
C3479 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PDM 0.02765f
C3480 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.Ien 0.04854f
C3481 XThC.Tn[4] XThR.Tn[1] 0.29363f
C3482 XA.XIR[2].XIC[6].icell.Ien Vbias 0.19161f
C3483 XA.XIR[11].XIC[4].icell.PUM VPWR 0.01015f
C3484 XThC.Tn[8] Iout 0.84039f
C3485 XThC.Tn[8] XThR.Tn[9] 0.29362f
C3486 XA.XIR[9].XIC[12].icell.Ien VPWR 0.1979f
C3487 XA.XIR[10].XIC[6].icell.PUM VPWR 0.01015f
C3488 XA.XIR[1].XIC[8].icell.Ien Vbias 0.19173f
C3489 XThR.XTB6.Y XThR.Tn[8] 0.02461f
C3490 XThC.Tn[4] XThR.Tn[12] 0.29362f
C3491 XThC.Tn[13] XThR.Tn[8] 0.29363f
C3492 XA.XIR[9].XIC[8].icell.Ien Iout 0.06821f
C3493 XThR.Tn[9] XA.XIR[9].XIC[8].icell.Ien 0.15202f
C3494 XThC.XTB3.Y XThC.XTBN.Y 0.17246f
C3495 XA.XIR[0].XIC[5].icell.Ien VPWR 0.19747f
C3496 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.04035f
C3497 XThR.XTB2.Y XThR.XTBN.A 0.04716f
C3498 XThR.XTBN.A a_n997_3755# 0.01939f
C3499 XThC.XTBN.Y XThC.Tn[2] 0.64352f
C3500 XA.XIR[3].XIC_15.icell.PUM VPWR 0.01655f
C3501 XThR.XTB7.A XThR.Tn[5] 0.02751f
C3502 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3503 XA.XIR[7].XIC[8].icell.Ien VPWR 0.1979f
C3504 XA.XIR[2].XIC[8].icell.PUM VPWR 0.01015f
C3505 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.Ien 0.04854f
C3506 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.PDM 0.02104f
C3507 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.Ien 0.04854f
C3508 XA.XIR[1].XIC[10].icell.PUM VPWR 0.01015f
C3509 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PDM 0.02765f
C3510 XA.XIR[7].XIC[4].icell.Ien Iout 0.06821f
C3511 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PDM 0.0404f
C3512 XThC.Tn[3] XThR.Tn[10] 0.29362f
C3513 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PDM 0.04035f
C3514 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PDM 0.02765f
C3515 XThC.XTB3.Y XThC.Tn[10] 0.29462f
C3516 XA.XIR[6].XIC[1].icell.PDM Vbias 0.03922f
C3517 XThC.Tn[5] XA.XIR[10].XIC[5].icell.Ien 0.03605f
C3518 XA.XIR[5].XIC[8].icell.PDM Vbias 0.03922f
C3519 a_n1049_8581# VPWR 0.71707f
C3520 XA.XIR[13].XIC[2].icell.PDM Vbias 0.03922f
C3521 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.PDM 0.02104f
C3522 XThR.Tn[3] Vbias 1.44825f
C3523 XThR.Tn[11] XA.XIR[11].XIC[4].icell.Ien 0.15202f
C3524 XThC.XTB1.Y XThC.XTB5.Y 0.05054f
C3525 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PDM 0.04035f
C3526 XA.XIR[12].XIC[7].icell.PDM Vbias 0.03922f
C3527 XThC.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.03605f
C3528 XA.XIR[10].XIC[0].icell.Ien VPWR 0.1979f
C3529 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.PDM 0.02104f
C3530 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout 0.06446f
C3531 XThC.Tn[8] XA.XIR[4].XIC[8].icell.Ien 0.03605f
C3532 XThR.XTB1.Y XThR.XTB5.Y 0.05054f
C3533 XThR.Tn[0] XA.XIR[0].XIC[9].icell.Ien 0.15202f
C3534 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.Ien 0.04854f
C3535 XThR.Tn[10] XA.XIR[10].XIC[8].icell.Ien 0.15202f
C3536 XThC.Tn[10] XA.XIR[14].XIC[10].icell.Ien 0.03605f
C3537 XThR.Tn[6] XA.XIR[6].XIC[3].icell.Ien 0.15202f
C3538 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.PDM 0.02104f
C3539 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.PDM 0.02104f
C3540 XThC.Tn[4] XA.XIR[7].XIC[4].icell.Ien 0.03605f
C3541 XA.XIR[15].XIC_15.icell.Ien Vbias 0.15966f
C3542 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.PDM 0.02104f
C3543 XThR.Tn[7] XA.XIR[7].XIC[10].icell.Ien 0.15202f
C3544 XA.XIR[6].XIC[8].icell.Ien Vbias 0.19161f
C3545 XThC.Tn[1] XA.XIR[5].XIC[1].icell.Ien 0.03605f
C3546 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.Ien 0.04854f
C3547 XThC.XTB1.Y XThC.XTBN.Y 0.1979f
C3548 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PDM 0.02765f
C3549 XThC.Tn[1] XThR.Tn[14] 0.29362f
C3550 XA.XIR[12].XIC_dummy_left.icell.Ien XThR.Tn[12] 0.01432f
C3551 XA.XIR[3].XIC[3].icell.PDM Vbias 0.03922f
C3552 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.PDM 0.02104f
C3553 XA.XIR[8].XIC[5].icell.PDM Vbias 0.03922f
C3554 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PDM 0.02896f
C3555 XA.XIR[14].XIC[2].icell.Ien Vbias 0.19161f
C3556 XThR.XTB2.Y a_n1049_7493# 0.02133f
C3557 XA.XIR[2].XIC[9].icell.PDM Vbias 0.03922f
C3558 XA.XIR[13].XIC[4].icell.Ien Vbias 0.19161f
C3559 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Iout 0.01728f
C3560 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.PDM 0.02104f
C3561 XA.XIR[12].XIC_dummy_left.icell.Iout VPWR 0.11103f
C3562 XA.XIR[3].XIC[5].icell.Ien VPWR 0.1979f
C3563 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.04035f
C3564 XThC.Tn[0] XA.XIR[13].XIC[0].icell.Ien 0.03605f
C3565 XA.XIR[6].XIC[10].icell.PUM VPWR 0.01015f
C3566 XThR.XTB2.Y XThR.XTB6.Y 0.04959f
C3567 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PDM 0.02765f
C3568 XThC.Tn[6] XA.XIR[9].XIC[6].icell.Ien 0.03605f
C3569 XA.XIR[11].XIC[7].icell.Ien Vbias 0.19161f
C3570 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.PDM 0.02104f
C3571 XThR.Tn[2] XA.XIR[2].XIC_15.icell.Ien 0.13564f
C3572 XThC.Tn[12] VPWR 7.41403f
C3573 XA.XIR[15].XIC[7].icell.Ien Iout 0.07211f
C3574 XThC.Tn[13] XA.XIR[0].XIC[13].icell.Ien 0.0373f
C3575 XA.XIR[10].XIC[9].icell.Ien Vbias 0.19161f
C3576 XA.XIR[4].XIC[14].icell.Ien VPWR 0.19796f
C3577 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Iout 0.0203f
C3578 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.Ien 0.04854f
C3579 XA.XIR[14].XIC[4].icell.PUM VPWR 0.01015f
C3580 XThC.XTBN.A a_7651_9569# 0.02087f
C3581 XA.XIR[4].XIC[10].icell.Ien Iout 0.06821f
C3582 XA.XIR[13].XIC[6].icell.PUM VPWR 0.01015f
C3583 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PDM 0.04035f
C3584 XA.XIR[0].XIC[1].icell.Ien Iout 0.06775f
C3585 XThC.Tn[7] XA.XIR[1].XIC[7].icell.Ien 0.03606f
C3586 XA.XIR[8].XIC[8].icell.Ien VPWR 0.1979f
C3587 XThR.XTB6.Y a_n1049_5611# 0.26831f
C3588 XA.XIR[8].XIC[4].icell.Ien Iout 0.06821f
C3589 XA.XIR[10].XIC_15.icell.PDM VPWR 0.07527f
C3590 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.Ien 0.04854f
C3591 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.Ien 0.04854f
C3592 XA.XIR[11].XIC[9].icell.PUM VPWR 0.01015f
C3593 XA.XIR[2].XIC[11].icell.Ien Vbias 0.19161f
C3594 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.PDM 0.02104f
C3595 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR 0.39108f
C3596 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PDM 0.04035f
C3597 XA.XIR[1].XIC[13].icell.Ien Vbias 0.19173f
C3598 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3599 XA.XIR[9].XIC[13].icell.Ien Iout 0.06821f
C3600 XThR.Tn[9] XA.XIR[9].XIC[13].icell.Ien 0.15202f
C3601 XA.XIR[0].XIC[10].icell.Ien VPWR 0.19726f
C3602 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.Ien 0.04854f
C3603 XThC.Tn[3] XThR.Tn[13] 0.29362f
C3604 bias[1] Vbias 0.05009f
C3605 XA.XIR[0].XIC[6].icell.Ien Iout 0.06775f
C3606 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PDM 0.04035f
C3607 XThC.Tn[5] XA.XIR[13].XIC[5].icell.Ien 0.03605f
C3608 XA.XIR[12].XIC[0].icell.Ien Vbias 0.19149f
C3609 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PDM 0.04035f
C3610 XThC.Tn[6] Iout 0.8414f
C3611 XA.XIR[2].XIC[13].icell.PUM VPWR 0.01015f
C3612 XA.XIR[7].XIC[13].icell.Ien VPWR 0.1979f
C3613 XThC.Tn[6] XThR.Tn[9] 0.29362f
C3614 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PDM 0.02765f
C3615 XThR.Tn[11] Vbias 1.4483f
C3616 XThC.Tn[2] XThR.Tn[8] 0.29362f
C3617 XThR.Tn[13] XA.XIR[13].XIC[3].icell.Ien 0.15202f
C3618 XA.XIR[7].XIC[9].icell.PDM Vbias 0.03922f
C3619 XA.XIR[7].XIC[9].icell.Ien Iout 0.06821f
C3620 XA.XIR[1].XIC_15.icell.PUM VPWR 0.01655f
C3621 XThC.Tn[4] XA.XIR[8].XIC[4].icell.Ien 0.03605f
C3622 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.Ien 0.04854f
C3623 XA.XIR[15].XIC[7].icell.PDM Vbias 0.03922f
C3624 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.Ien 0.04854f
C3625 XA.XIR[13].XIC[0].icell.Ien VPWR 0.1979f
C3626 XThC.XTBN.Y a_2979_9615# 0.0607f
C3627 XA.XIR[12].XIC[2].icell.PUM VPWR 0.01015f
C3628 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.Ien 0.04854f
C3629 XThR.XTB7.Y XThR.XTBN.A 1.11559f
C3630 XThR.XTBN.A data[4] 0.02581f
C3631 XThR.Tn[11] XA.XIR[11].XIC[9].icell.Ien 0.15202f
C3632 XA.XIR[9].XIC[5].icell.PDM Vbias 0.03922f
C3633 XA.XIR[2].XIC[0].icell.Ien Iout 0.06814f
C3634 data[2] data[3] 0.04128f
C3635 XThR.XTB5.A XThR.XTB7.A 0.07862f
C3636 XThR.XTB7.Y XThR.Tn[6] 0.21438f
C3637 XA.XIR[5].XIC[3].icell.PUM VPWR 0.01015f
C3638 a_9827_9569# XThC.Tn[12] 0.19481f
C3639 XThC.XTB6.A data[0] 0.48493f
C3640 XThC.Tn[7] XA.XIR[6].XIC[7].icell.Ien 0.03605f
C3641 XThC.Tn[0] XThC.Tn[1] 0.53527f
C3642 XThR.Tn[0] XA.XIR[0].XIC[14].icell.Ien 0.15202f
C3643 XA.XIR[10].XIC[1].icell.Ien Iout 0.06821f
C3644 XThC.Tn[13] XA.XIR[3].XIC[13].icell.Ien 0.03605f
C3645 XThR.Tn[6] XA.XIR[6].XIC[8].icell.Ien 0.15202f
C3646 a_n1049_7787# VPWR 0.72173f
C3647 XA.XIR[1].XIC[10].icell.PDM Vbias 0.03922f
C3648 XA.XIR[6].XIC[13].icell.Ien Vbias 0.19161f
C3649 XThR.Tn[7] XA.XIR[7].XIC_15.icell.Ien 0.13564f
C3650 XA.XIR[10].XIC[14].icell.Ien Vbias 0.19161f
C3651 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PDM 0.02765f
C3652 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.Ien 0.04854f
C3653 XA.XIR[4].XIC[10].icell.PDM Vbias 0.03922f
C3654 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.Ien 0.04854f
C3655 XThC.Tn[0] XA.XIR[6].XIC[0].icell.Ien 0.03605f
C3656 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PDM 0.02765f
C3657 XThC.Tn[14] XThR.Tn[7] 0.29368f
C3658 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.Ien 0.04854f
C3659 XThC.XTB5.A a_7331_10587# 0.01243f
C3660 XA.XIR[14].XIC[7].icell.Ien Vbias 0.19161f
C3661 XThR.XTB7.A data[5] 0.06538f
C3662 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.Ien 0.04854f
C3663 XA.XIR[13].XIC[9].icell.Ien Vbias 0.19161f
C3664 XThR.XTBN.Y XThR.Tn[5] 0.59912f
C3665 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PDM 0.04035f
C3666 XA.XIR[11].XIC[13].icell.Ien Iout 0.06821f
C3667 XThC.Tn[11] Vbias 1.15701f
C3668 XA.XIR[3].XIC[10].icell.Ien VPWR 0.1979f
C3669 XA.XIR[1].XIC[14].icell.PDM VPWR 0.01002f
C3670 XA.XIR[6].XIC_15.icell.PUM VPWR 0.01655f
C3671 XA.XIR[10].XIC[14].icell.PDM VPWR 0.01002f
C3672 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout 0.06446f
C3673 XA.XIR[3].XIC[6].icell.Ien Iout 0.06821f
C3674 XThR.XTBN.A a_n997_2667# 0.01679f
C3675 XThR.Tn[3] XThR.Tn[4] 0.10564f
C3676 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PDM 0.02765f
C3677 XA.XIR[2].XIC[3].icell.Ien VPWR 0.1979f
C3678 XA.XIR[4].XIC[14].icell.PDM VPWR 0.01002f
C3679 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR 0.01493f
C3680 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PDM 0.04035f
C3681 XA.XIR[13].XIC_15.icell.PDM VPWR 0.07527f
C3682 XA.XIR[1].XIC[5].icell.Ien VPWR 0.1979f
C3683 XA.XIR[14].XIC[9].icell.PUM VPWR 0.01015f
C3684 XA.XIR[4].XIC_15.icell.Ien Iout 0.0694f
C3685 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PDM 0.0404f
C3686 XA.XIR[8].XIC[13].icell.Ien VPWR 0.1979f
C3687 XThC.Tn[13] XThR.Tn[3] 0.29363f
C3688 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.Ien 0.04854f
C3689 XThC.XTB7.A XThC.XTBN.A 0.197f
C3690 XA.XIR[8].XIC[9].icell.Ien Iout 0.06821f
C3691 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PDM 0.02765f
C3692 XThC.XTB1.Y a_7651_9569# 0.06353f
C3693 XThC.Tn[1] VPWR 6.5068f
C3694 XA.XIR[1].XIC[0].icell.PUM VPWR 0.01015f
C3695 XA.XIR[5].XIC[1].icell.Ien Vbias 0.19161f
C3696 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PDM 0.02765f
C3697 XThR.XTB6.Y XThR.XTB7.Y 2.05133f
C3698 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PDM 0.04035f
C3699 XA.XIR[4].XIC[0].icell.PUM VPWR 0.01015f
C3700 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PDM 0.02765f
C3701 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.Ien 0.04854f
C3702 XThR.Tn[14] Vbias 1.44835f
C3703 XThR.XTBN.A XThR.Tn[11] 0.11968f
C3704 XThC.Tn[9] XThR.Tn[5] 0.29362f
C3705 XA.XIR[11].XIC[0].icell.PDM Vbias 0.03915f
C3706 XA.XIR[0].XIC_15.icell.Ien VPWR 0.26622f
C3707 XThC.Tn[14] XA.XIR[5].XIC[14].icell.Ien 0.03605f
C3708 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.04035f
C3709 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PDM 0.02838f
C3710 XA.XIR[10].XIC[4].icell.PDM Vbias 0.03922f
C3711 XThR.Tn[14] XA.XIR[14].XIC[4].icell.Ien 0.15202f
C3712 XA.XIR[0].XIC[11].icell.Ien Iout 0.06775f
C3713 XThR.Tn[1] XA.XIR[1].XIC[4].icell.Ien 0.15202f
C3714 XThR.Tn[11] XA.XIR[11].XIC[14].icell.Ien 0.15202f
C3715 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PDM 0.02765f
C3716 XA.XIR[4].XIC_dummy_right.icell.Iout Iout 0.01732f
C3717 XA.XIR[10].XIC[12].icell.Ien Vbias 0.19161f
C3718 XA.XIR[4].XIC_dummy_right.icell.Iout XA.XIR[5].XIC_dummy_right.icell.Iout 0.04047f
C3719 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout 0.06446f
C3720 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PDM 0.04035f
C3721 XA.XIR[6].XIC[0].icell.Ien VPWR 0.1979f
C3722 XThC.Tn[8] data[0] 0.01643f
C3723 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.Ien 0.04854f
C3724 XThR.XTB5.A XThR.XTB7.B 0.30355f
C3725 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PDM 0.02765f
C3726 XA.XIR[15].XIC_dummy_left.icell.Iout VPWR 0.25759f
C3727 XThR.Tn[13] XA.XIR[13].XIC[8].icell.Ien 0.15202f
C3728 XThC.Tn[10] XA.XIR[7].XIC[10].icell.Ien 0.03605f
C3729 XA.XIR[7].XIC[14].icell.Ien Iout 0.06821f
C3730 a_6243_9615# XThC.Tn[6] 0.26142f
C3731 XA.XIR[5].XIC[6].icell.Ien Vbias 0.19161f
C3732 XA.XIR[11].XIC[11].icell.Ien Iout 0.06821f
C3733 XA.XIR[0].XIC_dummy_right.icell.Iout VPWR 0.12361f
C3734 XA.XIR[11].XIC_dummy_right.icell.Iout XA.XIR[12].XIC_dummy_right.icell.Iout 0.04047f
C3735 XA.XIR[13].XIC[1].icell.Ien Iout 0.06821f
C3736 XThR.XTB6.A XThR.XTB5.Y 0.01866f
C3737 XA.XIR[6].XIC[5].icell.Ien VPWR 0.1979f
C3738 XA.XIR[0].XIC[12].icell.PDM Vbias 0.03943f
C3739 XA.XIR[5].XIC[8].icell.PUM VPWR 0.01015f
C3740 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PDM 0.02765f
C3741 XA.XIR[13].XIC[14].icell.Ien Vbias 0.19161f
C3742 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PDM 0.02765f
C3743 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PDM 0.02765f
C3744 XThC.Tn[12] XA.XIR[9].XIC[12].icell.Ien 0.03605f
C3745 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PDM 0.02765f
C3746 XThR.Tn[6] XA.XIR[6].XIC[13].icell.Ien 0.15202f
C3747 XThC.XTB5.A XThC.XTBN.A 0.06305f
C3748 XThC.XTB7.A XThC.XTB3.Y 0.57441f
C3749 XThC.Tn[2] XA.XIR[11].XIC[2].icell.Ien 0.03605f
C3750 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR 0.01669f
C3751 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PDM 0.02765f
C3752 XThC.XTB7.A XThC.Tn[2] 0.12602f
C3753 XA.XIR[12].XIC[3].icell.PUM VPWR 0.01015f
C3754 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.Ien 0.04854f
C3755 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR 0.08055f
C3756 XA.XIR[14].XIC[13].icell.Ien Iout 0.06821f
C3757 XA.XIR[11].XIC[4].icell.Ien VPWR 0.1979f
C3758 XThC.Tn[13] XA.XIR[1].XIC[13].icell.Ien 0.03605f
C3759 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PDM 0.04042f
C3760 XA.XIR[13].XIC[14].icell.PDM VPWR 0.01002f
C3761 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PDM 0.02765f
C3762 XA.XIR[10].XIC[6].icell.Ien VPWR 0.1979f
C3763 XThC.Tn[11] XThR.Tn[6] 0.29362f
C3764 XThR.Tn[11] XA.XIR[11].XIC[12].icell.Ien 0.15202f
C3765 XA.XIR[10].XIC[10].icell.Ien Vbias 0.19161f
C3766 XA.XIR[1].XIC[1].icell.Ien Iout 0.06821f
C3767 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.Ien 0.04854f
C3768 XA.XIR[10].XIC[2].icell.Ien Iout 0.06821f
C3769 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.Ien 0.04854f
C3770 XThR.XTB6.Y XThR.Tn[11] 0.02465f
C3771 XA.XIR[3].XIC_15.icell.Ien VPWR 0.26829f
C3772 XThC.Tn[13] XThR.Tn[11] 0.29363f
C3773 XThR.XTB1.Y XThR.XTB6.A 0.01609f
C3774 XA.XIR[3].XIC[11].icell.Ien Iout 0.06821f
C3775 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR 0.39039f
C3776 XA.XIR[2].XIC[8].icell.Ien VPWR 0.1979f
C3777 XThC.Tn[3] XThR.Tn[7] 0.29362f
C3778 XA.XIR[1].XIC[10].icell.Ien VPWR 0.1979f
C3779 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Iout 0.01758f
C3780 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR 0.38913f
C3781 XA.XIR[2].XIC[4].icell.Ien Iout 0.06821f
C3782 XThR.Tn[8] XA.XIR[8].XIC[5].icell.Ien 0.15202f
C3783 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PDM 0.04035f
C3784 XThC.Tn[0] Vbias 0.3936f
C3785 XA.XIR[1].XIC[6].icell.Ien Iout 0.06821f
C3786 XThC.XTB6.Y XThC.Tn[9] 0.0246f
C3787 XA.XIR[6].XIC[3].icell.PDM Vbias 0.03922f
C3788 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PDM 0.02765f
C3789 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.PDM 0.02104f
C3790 XThR.XTB1.Y XThR.Tn[0] 0.1837f
C3791 XA.XIR[5].XIC[10].icell.PDM Vbias 0.03922f
C3792 XA.XIR[14].XIC[0].icell.PDM Vbias 0.03915f
C3793 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PDM 0.02812f
C3794 XThC.Tn[10] XA.XIR[8].XIC[10].icell.Ien 0.03605f
C3795 XA.XIR[8].XIC[14].icell.Ien Iout 0.06821f
C3796 XThC.Tn[14] XA.XIR[12].XIC[14].icell.Ien 0.03605f
C3797 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PDM 0.02765f
C3798 XA.XIR[13].XIC[4].icell.PDM Vbias 0.03922f
C3799 XA.XIR[3].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3800 XA.XIR[13].XIC[12].icell.Ien Vbias 0.19161f
C3801 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.Ien 0.04854f
C3802 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.04035f
C3803 XThR.Tn[5] XA.XIR[5].XIC[4].icell.Ien 0.15202f
C3804 XA.XIR[12].XIC[9].icell.PDM Vbias 0.03922f
C3805 XThR.XTB7.B XThR.Tn[9] 0.0565f
C3806 XThC.XTB5.A XThC.XTB3.Y 0.01156f
C3807 XThC.XTB1.Y XThC.XTB7.A 0.48957f
C3808 XA.XIR[9].XIC[2].icell.Ien Vbias 0.19161f
C3809 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PDM 0.02765f
C3810 XThC.Tn[2] XThR.Tn[3] 0.29362f
C3811 XThR.Tn[14] XA.XIR[14].XIC[9].icell.Ien 0.15202f
C3812 XThC.XTBN.Y XThC.Tn[14] 0.50214f
C3813 XThR.Tn[1] XA.XIR[1].XIC[9].icell.Ien 0.15202f
C3814 XA.XIR[5].XIC[14].icell.PDM VPWR 0.01002f
C3815 XThC.Tn[13] XA.XIR[6].XIC[13].icell.Ien 0.03605f
C3816 XThC.Tn[11] XThR.Tn[4] 0.29362f
C3817 XThC.Tn[4] XA.XIR[2].XIC[4].icell.Ien 0.03605f
C3818 XA.XIR[14].XIC[11].icell.Ien Iout 0.06821f
C3819 XThR.XTB5.A XThR.XTB4.Y 0.02767f
C3820 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.PDM 0.02104f
C3821 XThC.XTB4.Y XThC.Tn[9] 0.01318f
C3822 XThC.Tn[1] XA.XIR[15].XIC[1].icell.Ien 0.03184f
C3823 XThC.XTB7.Y a_10051_9569# 0.013f
C3824 XA.XIR[6].XIC[1].icell.Ien Iout 0.06821f
C3825 XThR.Tn[11] XA.XIR[11].XIC[10].icell.Ien 0.15202f
C3826 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.PDM 0.02104f
C3827 XA.XIR[5].XIC[11].icell.Ien Vbias 0.19161f
C3828 XThC.Tn[5] XThR.Tn[0] 0.29368f
C3829 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8] 0.15202f
C3830 XThC.Tn[7] XThR.Tn[5] 0.29362f
C3831 XA.XIR[9].XIC[4].icell.PUM VPWR 0.01015f
C3832 XA.XIR[3].XIC[5].icell.PDM Vbias 0.03922f
C3833 XThR.Tn[2] Iout 1.19576f
C3834 XA.XIR[8].XIC[7].icell.PDM Vbias 0.03922f
C3835 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3836 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.Ien 0.04854f
C3837 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PDM 0.02765f
C3838 XA.XIR[2].XIC[11].icell.PDM Vbias 0.03922f
C3839 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PDM 0.02765f
C3840 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.Ien 0.04854f
C3841 XThC.Tn[2] XA.XIR[14].XIC[2].icell.Ien 0.03605f
C3842 XA.XIR[12].XIC[6].icell.Ien Vbias 0.19161f
C3843 XA.XIR[6].XIC[10].icell.Ien VPWR 0.1979f
C3844 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11] 0.15202f
C3845 XA.XIR[10].XIC_15.icell.Ien Vbias 0.19195f
C3846 VPWR Vbias 98.298f
C3847 XA.XIR[6].XIC[6].icell.Ien Iout 0.06821f
C3848 XA.XIR[5].XIC[13].icell.PUM VPWR 0.01015f
C3849 XA.XIR[14].XIC[4].icell.Ien VPWR 0.19845f
C3850 XThR.XTB5.Y XThR.Tn[12] 0.32095f
C3851 XA.XIR[2].XIC_15.icell.PDM VPWR 0.07527f
C3852 XThC.XTBN.A a_8739_9569# 0.01719f
C3853 XA.XIR[13].XIC[6].icell.Ien VPWR 0.1979f
C3854 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PDM 0.0404f
C3855 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PDM 0.04035f
C3856 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.PDM 0.02104f
C3857 XA.XIR[0].XIC_dummy_left.icell.Iout Iout 0.0353f
C3858 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout 0.06446f
C3859 XA.XIR[13].XIC[10].icell.Ien Vbias 0.19161f
C3860 XA.XIR[11].XIC_15.icell.PUM VPWR 0.01655f
C3861 XA.XIR[13].XIC[2].icell.Ien Iout 0.06821f
C3862 XA.XIR[12].XIC[8].icell.PUM VPWR 0.01015f
C3863 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR 0.01604f
C3864 XThC.Tn[4] XThR.Tn[2] 0.29362f
C3865 XThC.XTB5.A XThC.XTB1.Y 0.1098f
C3866 XA.XIR[11].XIC[9].icell.Ien VPWR 0.1979f
C3867 XThC.Tn[13] XThR.Tn[14] 0.29363f
C3868 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR 0.01604f
C3869 XA.XIR[11].XIC[5].icell.Ien Iout 0.06821f
C3870 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.PDM 0.02104f
C3871 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.PDM 0.02104f
C3872 XThR.XTB3.Y XThR.XTBN.A 0.03907f
C3873 a_7875_9569# XThC.Tn[9] 0.19329f
C3874 XA.XIR[10].XIC[7].icell.Ien Iout 0.06821f
C3875 XThC.XTB2.Y XThC.Tn[9] 0.292f
C3876 XA.XIR[2].XIC[0].icell.PUM VPWR 0.01015f
C3877 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Iout 0.01728f
C3878 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.PDM 0.02104f
C3879 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PDM 0.0404f
C3880 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PDM 0.04035f
C3881 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.Ien 0.04854f
C3882 XA.XIR[2].XIC[13].icell.Ien VPWR 0.1979f
C3883 XThR.XTBN.Y XThR.Tn[9] 0.48067f
C3884 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PDM 0.02765f
C3885 XThC.Tn[0] XThR.Tn[6] 0.29365f
C3886 XA.XIR[1].XIC[1].icell.PUM VPWR 0.01015f
C3887 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3888 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.PDM 0.02104f
C3889 XA.XIR[2].XIC[9].icell.Ien Iout 0.06821f
C3890 XA.XIR[1].XIC_15.icell.Ien VPWR 0.26829f
C3891 XA.XIR[7].XIC[11].icell.PDM Vbias 0.03922f
C3892 XThR.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.15202f
C3893 XThC.XTBN.A XThC.Tn[11] 0.12129f
C3894 XThR.Tn[8] XA.XIR[8].XIC[10].icell.Ien 0.15202f
C3895 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.Ien 0.04854f
C3896 XA.XIR[4].XIC[1].icell.PUM VPWR 0.01015f
C3897 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PDM 0.02778f
C3898 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.PDM 0.02104f
C3899 XA.XIR[1].XIC[11].icell.Ien Iout 0.06821f
C3900 XA.XIR[15].XIC[9].icell.PDM Vbias 0.03922f
C3901 XA.XIR[4].XIC[4].icell.Ien Vbias 0.19161f
C3902 XThC.Tn[2] XThR.Tn[11] 0.29362f
C3903 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR 0.35555f
C3904 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PDM 0.02765f
C3905 XThC.XTBN.Y a_4067_9615# 0.08456f
C3906 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.PDM 0.02104f
C3907 XThR.Tn[11] XA.XIR[11].XIC_15.icell.Ien 0.13564f
C3908 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.Ien 0.04854f
C3909 XThR.Tn[5] XA.XIR[5].XIC[9].icell.Ien 0.15202f
C3910 XA.XIR[9].XIC[7].icell.PDM Vbias 0.03922f
C3911 XThR.XTB4.Y XThR.Tn[9] 0.01318f
C3912 XA.XIR[15].XIC[3].icell.PUM VPWR 0.01015f
C3913 XA.XIR[5].XIC[3].icell.Ien VPWR 0.1979f
C3914 XA.XIR[7].XIC_15.icell.PDM VPWR 0.07527f
C3915 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.Ien 0.04854f
C3916 XThC.XTB3.Y a_8739_9569# 0.07285f
C3917 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PDM 0.02765f
C3918 XThC.XTB6.Y XThC.Tn[7] 0.01462f
C3919 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.Ien 0.04854f
C3920 XA.XIR[9].XIC[7].icell.Ien Vbias 0.19161f
C3921 XThR.Tn[10] Iout 1.1957f
C3922 XA.XIR[4].XIC[6].icell.PUM VPWR 0.01015f
C3923 XThR.Tn[9] XThR.Tn[10] 0.114f
C3924 XA.XIR[1].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3925 XA.XIR[11].XIC[13].icell.PUM VPWR 0.01015f
C3926 XThC.Tn[3] XA.XIR[0].XIC[3].icell.Ien 0.03715f
C3927 XThR.Tn[1] XA.XIR[1].XIC[14].icell.Ien 0.15202f
C3928 XThC.Tn[5] XThR.Tn[1] 0.29364f
C3929 XThC.Tn[9] Iout 0.84042f
C3930 XThC.Tn[9] XThR.Tn[9] 0.29362f
C3931 XA.XIR[1].XIC[12].icell.PDM Vbias 0.03922f
C3932 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.Ien 0.04854f
C3933 XThC.Tn[8] XA.XIR[11].XIC[8].icell.Ien 0.03605f
C3934 XThC.Tn[14] XThR.Tn[8] 0.29368f
C3935 XThC.Tn[5] XThR.Tn[12] 0.29362f
C3936 XA.XIR[7].XIC[3].icell.Ien Vbias 0.19161f
C3937 XA.XIR[4].XIC[12].icell.PDM Vbias 0.03922f
C3938 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.Ien 0.04854f
C3939 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.Ien 0.04854f
C3940 XThC.XTB6.Y a_5949_10571# 0.01283f
C3941 XThR.XTB3.Y a_n1049_7493# 0.23056f
C3942 XA.XIR[9].XIC[9].icell.PUM VPWR 0.01015f
C3943 XThC.XTB7.B Vbias 0.09218f
C3944 XThC.XTBN.Y XThC.Tn[3] 0.62681f
C3945 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.Ien 0.04854f
C3946 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.Ien 0.04854f
C3947 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.PDM 0.02104f
C3948 XA.XIR[13].XIC_15.icell.Ien Vbias 0.19195f
C3949 XThC.Tn[0] XThR.Tn[4] 0.29369f
C3950 XThR.XTBN.A VPWR 0.90694f
C3951 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.02765f
C3952 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.PDM 0.02104f
C3953 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PDM 0.02765f
C3954 XThC.XTBN.A data[1] 0.01444f
C3955 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12] 0.15202f
C3956 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.PDM 0.02104f
C3957 XThC.Tn[5] XA.XIR[4].XIC[5].icell.Ien 0.03605f
C3958 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PDM 0.04035f
C3959 XThR.XTB5.Y a_n1049_6405# 0.24821f
C3960 XA.XIR[11].XIC[14].icell.Ien VPWR 0.19796f
C3961 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PDM 0.04042f
C3962 XThR.Tn[6] VPWR 8.22274f
C3963 XThR.XTB3.Y XThR.XTB6.Y 0.04428f
C3964 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3965 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.PDM 0.02104f
C3966 XThC.XTB4.Y XThC.Tn[7] 0.01797f
C3967 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PDM 0.02765f
C3968 XThC.Tn[4] XThR.Tn[10] 0.29362f
C3969 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Ien 0.01721f
C3970 XA.XIR[6].XIC_15.icell.Ien VPWR 0.26829f
C3971 data[7] VGND 0.49949f
C3972 data[6] VGND 0.47974f
C3973 data[4] VGND 0.59317f
C3974 data[5] VGND 1.17814f
C3975 Iout VGND 0.32002p
C3976 bias[2] VGND 0.8011f
C3977 bias[0] VGND 2.64942f
C3978 Vbias VGND 0.16815p
C3979 bias[1] VGND 0.72457f
C3980 data[3] VGND 0.49912f
C3981 data[2] VGND 0.48064f
C3982 data[0] VGND 0.59421f
C3983 data[1] VGND 1.17844f
C3984 VPWR VGND 0.34898p
C3985 a_n997_715# VGND 0.5638f
C3986 XA.XIR[15].XIC_dummy_right.icell.Iout VGND 0.7524f
C3987 XA.XIR[15].XIC_dummy_right.icell.SM VGND 0.01013f
C3988 XA.XIR[15].XIC_dummy_right.icell.Ien VGND 0.64532f
C3989 XA.XIR[15].XIC_15.icell.Ien VGND 0.44493f
C3990 XA.XIR[15].XIC[14].icell.Ien VGND 0.44523f
C3991 XA.XIR[15].XIC[13].icell.Ien VGND 0.44523f
C3992 XA.XIR[15].XIC[12].icell.Ien VGND 0.44523f
C3993 XA.XIR[15].XIC[11].icell.Ien VGND 0.44523f
C3994 XA.XIR[15].XIC[10].icell.Ien VGND 0.44523f
C3995 XA.XIR[15].XIC[9].icell.Ien VGND 0.44523f
C3996 XA.XIR[15].XIC[8].icell.Ien VGND 0.44523f
C3997 XA.XIR[15].XIC[7].icell.Ien VGND 0.44523f
C3998 XA.XIR[15].XIC[6].icell.Ien VGND 0.44523f
C3999 XA.XIR[15].XIC[5].icell.Ien VGND 0.44523f
C4000 XA.XIR[15].XIC[4].icell.Ien VGND 0.44523f
C4001 XA.XIR[15].XIC[3].icell.Ien VGND 0.44523f
C4002 XA.XIR[15].XIC[2].icell.Ien VGND 0.44523f
C4003 XA.XIR[15].XIC_dummy_left.icell.Iout VGND 0.70718f
C4004 XA.XIR[15].XIC[1].icell.Ien VGND 0.44523f
C4005 XA.XIR[15].XIC[0].icell.Ien VGND 0.44537f
C4006 XA.XIR[15].XIC_dummy_left.icell.SM VGND 0.01044f
C4007 XA.XIR[15].XIC_dummy_left.icell.Ien VGND 0.61163f
C4008 XA.XIR[15].XIC_dummy_right.icell.PDM VGND 0.23278f
C4009 XA.XIR[15].XIC_15.icell.PDM VGND 0.18786f
C4010 XA.XIR[15].XIC[14].icell.PDM VGND 0.18741f
C4011 XA.XIR[15].XIC[13].icell.PDM VGND 0.18741f
C4012 XA.XIR[15].XIC[12].icell.PDM VGND 0.18741f
C4013 XA.XIR[15].XIC[11].icell.PDM VGND 0.18741f
C4014 XA.XIR[15].XIC[10].icell.PDM VGND 0.18741f
C4015 XA.XIR[15].XIC[9].icell.PDM VGND 0.18741f
C4016 XA.XIR[15].XIC[8].icell.PDM VGND 0.18741f
C4017 XA.XIR[15].XIC[7].icell.PDM VGND 0.18741f
C4018 XA.XIR[15].XIC[6].icell.PDM VGND 0.18741f
C4019 XA.XIR[15].XIC[5].icell.PDM VGND 0.18741f
C4020 XA.XIR[15].XIC[4].icell.PDM VGND 0.18741f
C4021 XA.XIR[15].XIC[3].icell.PDM VGND 0.18741f
C4022 XA.XIR[15].XIC[2].icell.PDM VGND 0.18741f
C4023 XA.XIR[15].XIC[1].icell.PDM VGND 0.18741f
C4024 XA.XIR[15].XIC[0].icell.PDM VGND 0.18748f
C4025 XA.XIR[15].XIC_dummy_left.icell.PDM VGND 0.22703f
C4026 XA.XIR[14].XIC_dummy_right.icell.Iout VGND 0.85788f
C4027 XA.XIR[14].XIC_dummy_right.icell.SM VGND 0.01013f
C4028 XA.XIR[14].XIC_dummy_right.icell.Ien VGND 0.60818f
C4029 XA.XIR[14].XIC_15.icell.Ien VGND 0.37264f
C4030 XA.XIR[14].XIC[14].icell.Ien VGND 0.37345f
C4031 XA.XIR[14].XIC[13].icell.Ien VGND 0.37345f
C4032 XA.XIR[14].XIC[12].icell.Ien VGND 0.37345f
C4033 XA.XIR[14].XIC[11].icell.Ien VGND 0.37345f
C4034 XA.XIR[14].XIC[10].icell.Ien VGND 0.37345f
C4035 XA.XIR[14].XIC[9].icell.Ien VGND 0.37345f
C4036 XA.XIR[14].XIC[8].icell.Ien VGND 0.37345f
C4037 XA.XIR[14].XIC[7].icell.Ien VGND 0.37345f
C4038 XA.XIR[14].XIC[6].icell.Ien VGND 0.37345f
C4039 XA.XIR[14].XIC[5].icell.Ien VGND 0.37345f
C4040 XA.XIR[14].XIC[4].icell.Ien VGND 0.37345f
C4041 XA.XIR[14].XIC[3].icell.Ien VGND 0.37345f
C4042 XA.XIR[14].XIC[2].icell.Ien VGND 0.37345f
C4043 XA.XIR[14].XIC_dummy_left.icell.Iout VGND 0.80696f
C4044 XThR.Tn[14] VGND 13.42928f
C4045 XA.XIR[14].XIC[1].icell.Ien VGND 0.37345f
C4046 a_n997_1579# VGND 0.54776f
C4047 XA.XIR[14].XIC[0].icell.Ien VGND 0.37359f
C4048 XA.XIR[14].XIC_dummy_left.icell.SM VGND 0.01044f
C4049 XA.XIR[14].XIC_dummy_left.icell.Ien VGND 0.57579f
C4050 a_n997_1803# VGND 0.53619f
C4051 XA.XIR[14].XIC_dummy_right.icell.PDM VGND 0.23384f
C4052 XA.XIR[14].XIC_15.icell.PDM VGND 0.18862f
C4053 XA.XIR[14].XIC[14].icell.PDM VGND 0.18817f
C4054 XA.XIR[14].XIC[13].icell.PDM VGND 0.18817f
C4055 XA.XIR[14].XIC[12].icell.PDM VGND 0.18817f
C4056 XA.XIR[14].XIC[11].icell.PDM VGND 0.18817f
C4057 XA.XIR[14].XIC[10].icell.PDM VGND 0.18817f
C4058 XA.XIR[14].XIC[9].icell.PDM VGND 0.18817f
C4059 XA.XIR[14].XIC[8].icell.PDM VGND 0.18817f
C4060 XA.XIR[14].XIC[7].icell.PDM VGND 0.18817f
C4061 XA.XIR[14].XIC[6].icell.PDM VGND 0.18817f
C4062 XA.XIR[14].XIC[5].icell.PDM VGND 0.18817f
C4063 XA.XIR[14].XIC[4].icell.PDM VGND 0.18817f
C4064 XA.XIR[14].XIC[3].icell.PDM VGND 0.18817f
C4065 XA.XIR[14].XIC[2].icell.PDM VGND 0.18817f
C4066 XA.XIR[14].XIC[1].icell.PDM VGND 0.18817f
C4067 XA.XIR[14].XIC[0].icell.PDM VGND 0.18824f
C4068 XA.XIR[14].XIC_dummy_left.icell.PDM VGND 0.22809f
C4069 XA.XIR[13].XIC_dummy_right.icell.Iout VGND 0.85788f
C4070 XA.XIR[13].XIC_dummy_right.icell.SM VGND 0.01013f
C4071 XA.XIR[13].XIC_dummy_right.icell.Ien VGND 0.60818f
C4072 XA.XIR[13].XIC_15.icell.Ien VGND 0.37264f
C4073 XA.XIR[13].XIC[14].icell.Ien VGND 0.37345f
C4074 XA.XIR[13].XIC[13].icell.Ien VGND 0.37345f
C4075 XA.XIR[13].XIC[12].icell.Ien VGND 0.37345f
C4076 XA.XIR[13].XIC[11].icell.Ien VGND 0.37345f
C4077 XA.XIR[13].XIC[10].icell.Ien VGND 0.37345f
C4078 XA.XIR[13].XIC[9].icell.Ien VGND 0.37345f
C4079 XA.XIR[13].XIC[8].icell.Ien VGND 0.37345f
C4080 XA.XIR[13].XIC[7].icell.Ien VGND 0.37345f
C4081 XA.XIR[13].XIC[6].icell.Ien VGND 0.37345f
C4082 XA.XIR[13].XIC[5].icell.Ien VGND 0.37345f
C4083 XA.XIR[13].XIC[4].icell.Ien VGND 0.37345f
C4084 XA.XIR[13].XIC[3].icell.Ien VGND 0.37345f
C4085 XA.XIR[13].XIC[2].icell.Ien VGND 0.37345f
C4086 XA.XIR[13].XIC_dummy_left.icell.Iout VGND 0.807f
C4087 XThR.Tn[13] VGND 13.31119f
C4088 XA.XIR[13].XIC[1].icell.Ien VGND 0.37345f
C4089 XA.XIR[13].XIC[0].icell.Ien VGND 0.37359f
C4090 XA.XIR[13].XIC_dummy_left.icell.SM VGND 0.01044f
C4091 XA.XIR[13].XIC_dummy_left.icell.Ien VGND 0.57425f
C4092 XA.XIR[13].XIC_dummy_right.icell.PDM VGND 0.23384f
C4093 XA.XIR[13].XIC_15.icell.PDM VGND 0.18862f
C4094 XA.XIR[13].XIC[14].icell.PDM VGND 0.18817f
C4095 XA.XIR[13].XIC[13].icell.PDM VGND 0.18817f
C4096 XA.XIR[13].XIC[12].icell.PDM VGND 0.18817f
C4097 XA.XIR[13].XIC[11].icell.PDM VGND 0.18817f
C4098 XA.XIR[13].XIC[10].icell.PDM VGND 0.18817f
C4099 XA.XIR[13].XIC[9].icell.PDM VGND 0.18817f
C4100 XA.XIR[13].XIC[8].icell.PDM VGND 0.18817f
C4101 XA.XIR[13].XIC[7].icell.PDM VGND 0.18817f
C4102 XA.XIR[13].XIC[6].icell.PDM VGND 0.18817f
C4103 XA.XIR[13].XIC[5].icell.PDM VGND 0.18817f
C4104 XA.XIR[13].XIC[4].icell.PDM VGND 0.18817f
C4105 XA.XIR[13].XIC[3].icell.PDM VGND 0.18817f
C4106 XA.XIR[13].XIC[2].icell.PDM VGND 0.18817f
C4107 XA.XIR[13].XIC[1].icell.PDM VGND 0.18817f
C4108 XA.XIR[13].XIC[0].icell.PDM VGND 0.18824f
C4109 XA.XIR[13].XIC_dummy_left.icell.PDM VGND 0.22809f
C4110 XA.XIR[12].XIC_dummy_right.icell.Iout VGND 0.85788f
C4111 XA.XIR[12].XIC_dummy_right.icell.SM VGND 0.01013f
C4112 XA.XIR[12].XIC_dummy_right.icell.Ien VGND 0.60818f
C4113 XA.XIR[12].XIC_15.icell.Ien VGND 0.37264f
C4114 XA.XIR[12].XIC[14].icell.Ien VGND 0.37345f
C4115 XA.XIR[12].XIC[13].icell.Ien VGND 0.37345f
C4116 XA.XIR[12].XIC[12].icell.Ien VGND 0.37345f
C4117 XA.XIR[12].XIC[11].icell.Ien VGND 0.37345f
C4118 XA.XIR[12].XIC[10].icell.Ien VGND 0.37345f
C4119 XA.XIR[12].XIC[9].icell.Ien VGND 0.37345f
C4120 XA.XIR[12].XIC[8].icell.Ien VGND 0.37345f
C4121 XA.XIR[12].XIC[7].icell.Ien VGND 0.37345f
C4122 XA.XIR[12].XIC[6].icell.Ien VGND 0.37345f
C4123 XA.XIR[12].XIC[5].icell.Ien VGND 0.37345f
C4124 XA.XIR[12].XIC[4].icell.Ien VGND 0.37345f
C4125 XA.XIR[12].XIC[3].icell.Ien VGND 0.37345f
C4126 XA.XIR[12].XIC[2].icell.Ien VGND 0.37345f
C4127 XA.XIR[12].XIC_dummy_left.icell.Iout VGND 0.80565f
C4128 XThR.Tn[12] VGND 13.163f
C4129 XA.XIR[12].XIC[1].icell.Ien VGND 0.37345f
C4130 XA.XIR[12].XIC[0].icell.Ien VGND 0.37359f
C4131 XA.XIR[12].XIC_dummy_left.icell.SM VGND 0.01044f
C4132 XA.XIR[12].XIC_dummy_left.icell.Ien VGND 0.57283f
C4133 a_n997_2667# VGND 0.5457f
C4134 XA.XIR[12].XIC_dummy_right.icell.PDM VGND 0.23384f
C4135 XA.XIR[12].XIC_15.icell.PDM VGND 0.18862f
C4136 XA.XIR[12].XIC[14].icell.PDM VGND 0.18817f
C4137 XA.XIR[12].XIC[13].icell.PDM VGND 0.18817f
C4138 XA.XIR[12].XIC[12].icell.PDM VGND 0.18817f
C4139 XA.XIR[12].XIC[11].icell.PDM VGND 0.18817f
C4140 XA.XIR[12].XIC[10].icell.PDM VGND 0.18817f
C4141 XA.XIR[12].XIC[9].icell.PDM VGND 0.18817f
C4142 XA.XIR[12].XIC[8].icell.PDM VGND 0.18817f
C4143 XA.XIR[12].XIC[7].icell.PDM VGND 0.18817f
C4144 XA.XIR[12].XIC[6].icell.PDM VGND 0.18817f
C4145 XA.XIR[12].XIC[5].icell.PDM VGND 0.18817f
C4146 XA.XIR[12].XIC[4].icell.PDM VGND 0.18817f
C4147 XA.XIR[12].XIC[3].icell.PDM VGND 0.18817f
C4148 XA.XIR[12].XIC[2].icell.PDM VGND 0.18817f
C4149 XA.XIR[12].XIC[1].icell.PDM VGND 0.18817f
C4150 XA.XIR[12].XIC[0].icell.PDM VGND 0.18824f
C4151 XA.XIR[12].XIC_dummy_left.icell.PDM VGND 0.22809f
C4152 XA.XIR[11].XIC_dummy_right.icell.Iout VGND 0.85788f
C4153 XA.XIR[11].XIC_dummy_right.icell.SM VGND 0.01013f
C4154 XA.XIR[11].XIC_dummy_right.icell.Ien VGND 0.60818f
C4155 XA.XIR[11].XIC_15.icell.Ien VGND 0.37264f
C4156 XA.XIR[11].XIC[14].icell.Ien VGND 0.37345f
C4157 XA.XIR[11].XIC[13].icell.Ien VGND 0.37345f
C4158 XA.XIR[11].XIC[12].icell.Ien VGND 0.37345f
C4159 XA.XIR[11].XIC[11].icell.Ien VGND 0.37345f
C4160 XA.XIR[11].XIC[10].icell.Ien VGND 0.37345f
C4161 XA.XIR[11].XIC[9].icell.Ien VGND 0.37345f
C4162 XA.XIR[11].XIC[8].icell.Ien VGND 0.37345f
C4163 XA.XIR[11].XIC[7].icell.Ien VGND 0.37345f
C4164 XA.XIR[11].XIC[6].icell.Ien VGND 0.37345f
C4165 XA.XIR[11].XIC[5].icell.Ien VGND 0.37345f
C4166 XA.XIR[11].XIC[4].icell.Ien VGND 0.37345f
C4167 XA.XIR[11].XIC[3].icell.Ien VGND 0.37345f
C4168 XA.XIR[11].XIC[2].icell.Ien VGND 0.37345f
C4169 XA.XIR[11].XIC_dummy_left.icell.Iout VGND 0.808f
C4170 XThR.Tn[11] VGND 13.22524f
C4171 XA.XIR[11].XIC[1].icell.Ien VGND 0.37345f
C4172 a_n997_2891# VGND 0.54795f
C4173 XA.XIR[11].XIC[0].icell.Ien VGND 0.37359f
C4174 XA.XIR[11].XIC_dummy_left.icell.SM VGND 0.01044f
C4175 XA.XIR[11].XIC_dummy_left.icell.Ien VGND 0.57297f
C4176 XA.XIR[11].XIC_dummy_right.icell.PDM VGND 0.23384f
C4177 XA.XIR[11].XIC_15.icell.PDM VGND 0.18862f
C4178 XA.XIR[11].XIC[14].icell.PDM VGND 0.18817f
C4179 XA.XIR[11].XIC[13].icell.PDM VGND 0.18817f
C4180 XA.XIR[11].XIC[12].icell.PDM VGND 0.18817f
C4181 XA.XIR[11].XIC[11].icell.PDM VGND 0.18817f
C4182 XA.XIR[11].XIC[10].icell.PDM VGND 0.18817f
C4183 XA.XIR[11].XIC[9].icell.PDM VGND 0.18817f
C4184 XA.XIR[11].XIC[8].icell.PDM VGND 0.18817f
C4185 XA.XIR[11].XIC[7].icell.PDM VGND 0.18817f
C4186 XA.XIR[11].XIC[6].icell.PDM VGND 0.18817f
C4187 XA.XIR[11].XIC[5].icell.PDM VGND 0.18817f
C4188 XA.XIR[11].XIC[4].icell.PDM VGND 0.18817f
C4189 XA.XIR[11].XIC[3].icell.PDM VGND 0.18817f
C4190 XA.XIR[11].XIC[2].icell.PDM VGND 0.18817f
C4191 XA.XIR[11].XIC[1].icell.PDM VGND 0.18817f
C4192 XA.XIR[11].XIC[0].icell.PDM VGND 0.18824f
C4193 XA.XIR[11].XIC_dummy_left.icell.PDM VGND 0.22809f
C4194 XA.XIR[10].XIC_dummy_right.icell.Iout VGND 0.85788f
C4195 XA.XIR[10].XIC_dummy_right.icell.SM VGND 0.01013f
C4196 XA.XIR[10].XIC_dummy_right.icell.Ien VGND 0.60818f
C4197 XA.XIR[10].XIC_15.icell.Ien VGND 0.37264f
C4198 XA.XIR[10].XIC[14].icell.Ien VGND 0.37345f
C4199 XA.XIR[10].XIC[13].icell.Ien VGND 0.37345f
C4200 XA.XIR[10].XIC[12].icell.Ien VGND 0.37345f
C4201 XA.XIR[10].XIC[11].icell.Ien VGND 0.37345f
C4202 XA.XIR[10].XIC[10].icell.Ien VGND 0.37345f
C4203 XA.XIR[10].XIC[9].icell.Ien VGND 0.37345f
C4204 XA.XIR[10].XIC[8].icell.Ien VGND 0.37345f
C4205 XA.XIR[10].XIC[7].icell.Ien VGND 0.37345f
C4206 XA.XIR[10].XIC[6].icell.Ien VGND 0.37345f
C4207 XA.XIR[10].XIC[5].icell.Ien VGND 0.37345f
C4208 XA.XIR[10].XIC[4].icell.Ien VGND 0.37345f
C4209 XA.XIR[10].XIC[3].icell.Ien VGND 0.37345f
C4210 XA.XIR[10].XIC[2].icell.Ien VGND 0.37345f
C4211 XA.XIR[10].XIC_dummy_left.icell.Iout VGND 0.80684f
C4212 XThR.Tn[10] VGND 13.20071f
C4213 XA.XIR[10].XIC[1].icell.Ien VGND 0.37345f
C4214 XA.XIR[10].XIC[0].icell.Ien VGND 0.37359f
C4215 XA.XIR[10].XIC_dummy_left.icell.SM VGND 0.01044f
C4216 XA.XIR[10].XIC_dummy_left.icell.Ien VGND 0.57425f
C4217 XA.XIR[10].XIC_dummy_right.icell.PDM VGND 0.23384f
C4218 XA.XIR[10].XIC_15.icell.PDM VGND 0.18862f
C4219 XA.XIR[10].XIC[14].icell.PDM VGND 0.18817f
C4220 XA.XIR[10].XIC[13].icell.PDM VGND 0.18817f
C4221 XA.XIR[10].XIC[12].icell.PDM VGND 0.18817f
C4222 XA.XIR[10].XIC[11].icell.PDM VGND 0.18817f
C4223 XA.XIR[10].XIC[10].icell.PDM VGND 0.18817f
C4224 XA.XIR[10].XIC[9].icell.PDM VGND 0.18817f
C4225 XA.XIR[10].XIC[8].icell.PDM VGND 0.18817f
C4226 XA.XIR[10].XIC[7].icell.PDM VGND 0.18817f
C4227 XA.XIR[10].XIC[6].icell.PDM VGND 0.18817f
C4228 XA.XIR[10].XIC[5].icell.PDM VGND 0.18817f
C4229 XA.XIR[10].XIC[4].icell.PDM VGND 0.18817f
C4230 XA.XIR[10].XIC[3].icell.PDM VGND 0.18817f
C4231 XA.XIR[10].XIC[2].icell.PDM VGND 0.18817f
C4232 XA.XIR[10].XIC[1].icell.PDM VGND 0.18817f
C4233 XA.XIR[10].XIC[0].icell.PDM VGND 0.18824f
C4234 XA.XIR[10].XIC_dummy_left.icell.PDM VGND 0.22809f
C4235 XA.XIR[9].XIC_dummy_right.icell.Iout VGND 0.85788f
C4236 XA.XIR[9].XIC_dummy_right.icell.SM VGND 0.01013f
C4237 XA.XIR[9].XIC_dummy_right.icell.Ien VGND 0.60818f
C4238 XA.XIR[9].XIC_15.icell.Ien VGND 0.37264f
C4239 XA.XIR[9].XIC[14].icell.Ien VGND 0.37345f
C4240 XA.XIR[9].XIC[13].icell.Ien VGND 0.37345f
C4241 XA.XIR[9].XIC[12].icell.Ien VGND 0.37345f
C4242 XA.XIR[9].XIC[11].icell.Ien VGND 0.37345f
C4243 XA.XIR[9].XIC[10].icell.Ien VGND 0.37345f
C4244 XA.XIR[9].XIC[9].icell.Ien VGND 0.37345f
C4245 XA.XIR[9].XIC[8].icell.Ien VGND 0.37345f
C4246 XA.XIR[9].XIC[7].icell.Ien VGND 0.37345f
C4247 XA.XIR[9].XIC[6].icell.Ien VGND 0.37345f
C4248 XA.XIR[9].XIC[5].icell.Ien VGND 0.37345f
C4249 XA.XIR[9].XIC[4].icell.Ien VGND 0.37345f
C4250 XA.XIR[9].XIC[3].icell.Ien VGND 0.37345f
C4251 XA.XIR[9].XIC[2].icell.Ien VGND 0.37345f
C4252 XA.XIR[9].XIC_dummy_left.icell.Iout VGND 0.8087f
C4253 XA.XIR[9].XIC[1].icell.Ien VGND 0.37345f
C4254 XThR.Tn[9] VGND 13.20833f
C4255 a_n997_3755# VGND 0.54861f
C4256 XA.XIR[9].XIC[0].icell.Ien VGND 0.37359f
C4257 XA.XIR[9].XIC_dummy_left.icell.SM VGND 0.01044f
C4258 XA.XIR[9].XIC_dummy_left.icell.Ien VGND 0.57323f
C4259 a_n997_3979# VGND 0.54721f
C4260 XA.XIR[9].XIC_dummy_right.icell.PDM VGND 0.23384f
C4261 XA.XIR[9].XIC_15.icell.PDM VGND 0.18862f
C4262 XA.XIR[9].XIC[14].icell.PDM VGND 0.18817f
C4263 XA.XIR[9].XIC[13].icell.PDM VGND 0.18817f
C4264 XA.XIR[9].XIC[12].icell.PDM VGND 0.18817f
C4265 XA.XIR[9].XIC[11].icell.PDM VGND 0.18817f
C4266 XA.XIR[9].XIC[10].icell.PDM VGND 0.18817f
C4267 XA.XIR[9].XIC[9].icell.PDM VGND 0.18817f
C4268 XA.XIR[9].XIC[8].icell.PDM VGND 0.18817f
C4269 XA.XIR[9].XIC[7].icell.PDM VGND 0.18817f
C4270 XA.XIR[9].XIC[6].icell.PDM VGND 0.18817f
C4271 XA.XIR[9].XIC[5].icell.PDM VGND 0.18817f
C4272 XA.XIR[9].XIC[4].icell.PDM VGND 0.18817f
C4273 XA.XIR[9].XIC[3].icell.PDM VGND 0.18817f
C4274 XA.XIR[9].XIC[2].icell.PDM VGND 0.18817f
C4275 XA.XIR[9].XIC[1].icell.PDM VGND 0.18817f
C4276 XA.XIR[9].XIC[0].icell.PDM VGND 0.18824f
C4277 XA.XIR[9].XIC_dummy_left.icell.PDM VGND 0.22809f
C4278 XA.XIR[8].XIC_dummy_right.icell.Iout VGND 0.85788f
C4279 XA.XIR[8].XIC_dummy_right.icell.SM VGND 0.01013f
C4280 XA.XIR[8].XIC_dummy_right.icell.Ien VGND 0.60818f
C4281 XA.XIR[8].XIC_15.icell.Ien VGND 0.37264f
C4282 XA.XIR[8].XIC[14].icell.Ien VGND 0.37345f
C4283 XA.XIR[8].XIC[13].icell.Ien VGND 0.37345f
C4284 XA.XIR[8].XIC[12].icell.Ien VGND 0.37345f
C4285 XA.XIR[8].XIC[11].icell.Ien VGND 0.37345f
C4286 XA.XIR[8].XIC[10].icell.Ien VGND 0.37345f
C4287 XA.XIR[8].XIC[9].icell.Ien VGND 0.37345f
C4288 XA.XIR[8].XIC[8].icell.Ien VGND 0.37345f
C4289 XA.XIR[8].XIC[7].icell.Ien VGND 0.37345f
C4290 XA.XIR[8].XIC[6].icell.Ien VGND 0.37345f
C4291 XA.XIR[8].XIC[5].icell.Ien VGND 0.37345f
C4292 XA.XIR[8].XIC[4].icell.Ien VGND 0.37345f
C4293 XA.XIR[8].XIC[3].icell.Ien VGND 0.37345f
C4294 XA.XIR[8].XIC[2].icell.Ien VGND 0.37345f
C4295 XA.XIR[8].XIC_dummy_left.icell.Iout VGND 0.80602f
C4296 XA.XIR[8].XIC[1].icell.Ien VGND 0.37345f
C4297 XThR.Tn[8] VGND 13.18672f
C4298 XA.XIR[8].XIC[0].icell.Ien VGND 0.37359f
C4299 XA.XIR[8].XIC_dummy_left.icell.SM VGND 0.01044f
C4300 XA.XIR[8].XIC_dummy_left.icell.Ien VGND 0.57311f
C4301 XA.XIR[8].XIC_dummy_right.icell.PDM VGND 0.23384f
C4302 XA.XIR[8].XIC_15.icell.PDM VGND 0.18862f
C4303 XA.XIR[8].XIC[14].icell.PDM VGND 0.18817f
C4304 XA.XIR[8].XIC[13].icell.PDM VGND 0.18817f
C4305 XA.XIR[8].XIC[12].icell.PDM VGND 0.18817f
C4306 XA.XIR[8].XIC[11].icell.PDM VGND 0.18817f
C4307 XA.XIR[8].XIC[10].icell.PDM VGND 0.18817f
C4308 XA.XIR[8].XIC[9].icell.PDM VGND 0.18817f
C4309 XA.XIR[8].XIC[8].icell.PDM VGND 0.18817f
C4310 XA.XIR[8].XIC[7].icell.PDM VGND 0.18817f
C4311 XA.XIR[8].XIC[6].icell.PDM VGND 0.18817f
C4312 XA.XIR[8].XIC[5].icell.PDM VGND 0.18817f
C4313 XA.XIR[8].XIC[4].icell.PDM VGND 0.18817f
C4314 XA.XIR[8].XIC[3].icell.PDM VGND 0.18817f
C4315 XA.XIR[8].XIC[2].icell.PDM VGND 0.18817f
C4316 XA.XIR[8].XIC[1].icell.PDM VGND 0.18817f
C4317 XA.XIR[8].XIC[0].icell.PDM VGND 0.18824f
C4318 XA.XIR[8].XIC_dummy_left.icell.PDM VGND 0.22809f
C4319 XA.XIR[7].XIC_dummy_right.icell.Iout VGND 0.85788f
C4320 XA.XIR[7].XIC_dummy_right.icell.SM VGND 0.01013f
C4321 XA.XIR[7].XIC_dummy_right.icell.Ien VGND 0.60818f
C4322 XA.XIR[7].XIC_15.icell.Ien VGND 0.37264f
C4323 XA.XIR[7].XIC[14].icell.Ien VGND 0.37345f
C4324 XA.XIR[7].XIC[13].icell.Ien VGND 0.37345f
C4325 XA.XIR[7].XIC[12].icell.Ien VGND 0.37345f
C4326 XA.XIR[7].XIC[11].icell.Ien VGND 0.37345f
C4327 XA.XIR[7].XIC[10].icell.Ien VGND 0.37345f
C4328 XA.XIR[7].XIC[9].icell.Ien VGND 0.37345f
C4329 XA.XIR[7].XIC[8].icell.Ien VGND 0.37345f
C4330 XA.XIR[7].XIC[7].icell.Ien VGND 0.37345f
C4331 XA.XIR[7].XIC[6].icell.Ien VGND 0.37345f
C4332 XA.XIR[7].XIC[5].icell.Ien VGND 0.37345f
C4333 XA.XIR[7].XIC[4].icell.Ien VGND 0.37345f
C4334 XA.XIR[7].XIC[3].icell.Ien VGND 0.37345f
C4335 XA.XIR[7].XIC[2].icell.Ien VGND 0.37345f
C4336 XA.XIR[7].XIC_dummy_left.icell.Iout VGND 0.80634f
C4337 XA.XIR[7].XIC[1].icell.Ien VGND 0.37345f
C4338 XA.XIR[7].XIC[0].icell.Ien VGND 0.37359f
C4339 XA.XIR[7].XIC_dummy_left.icell.SM VGND 0.01044f
C4340 XThR.Tn[7] VGND 13.59514f
C4341 XThR.XTBN.A VGND 1.22814f
C4342 XA.XIR[7].XIC_dummy_left.icell.Ien VGND 0.57579f
C4343 XA.XIR[7].XIC_dummy_right.icell.PDM VGND 0.23384f
C4344 XA.XIR[7].XIC_15.icell.PDM VGND 0.18862f
C4345 XA.XIR[7].XIC[14].icell.PDM VGND 0.18817f
C4346 XA.XIR[7].XIC[13].icell.PDM VGND 0.18817f
C4347 XA.XIR[7].XIC[12].icell.PDM VGND 0.18817f
C4348 XA.XIR[7].XIC[11].icell.PDM VGND 0.18817f
C4349 XA.XIR[7].XIC[10].icell.PDM VGND 0.18817f
C4350 XA.XIR[7].XIC[9].icell.PDM VGND 0.18817f
C4351 XA.XIR[7].XIC[8].icell.PDM VGND 0.18817f
C4352 XA.XIR[7].XIC[7].icell.PDM VGND 0.18817f
C4353 XA.XIR[7].XIC[6].icell.PDM VGND 0.18817f
C4354 XA.XIR[7].XIC[5].icell.PDM VGND 0.18817f
C4355 XA.XIR[7].XIC[4].icell.PDM VGND 0.18817f
C4356 XA.XIR[7].XIC[3].icell.PDM VGND 0.18817f
C4357 XA.XIR[7].XIC[2].icell.PDM VGND 0.18817f
C4358 XA.XIR[7].XIC[1].icell.PDM VGND 0.18817f
C4359 XA.XIR[7].XIC[0].icell.PDM VGND 0.18824f
C4360 XA.XIR[7].XIC_dummy_left.icell.PDM VGND 0.22809f
C4361 XA.XIR[6].XIC_dummy_right.icell.Iout VGND 0.85788f
C4362 XA.XIR[6].XIC_dummy_right.icell.SM VGND 0.01013f
C4363 XA.XIR[6].XIC_dummy_right.icell.Ien VGND 0.60818f
C4364 XA.XIR[6].XIC_15.icell.Ien VGND 0.37264f
C4365 XA.XIR[6].XIC[14].icell.Ien VGND 0.37345f
C4366 XA.XIR[6].XIC[13].icell.Ien VGND 0.37345f
C4367 XA.XIR[6].XIC[12].icell.Ien VGND 0.37345f
C4368 XA.XIR[6].XIC[11].icell.Ien VGND 0.37345f
C4369 XA.XIR[6].XIC[10].icell.Ien VGND 0.37345f
C4370 XA.XIR[6].XIC[9].icell.Ien VGND 0.37345f
C4371 XA.XIR[6].XIC[8].icell.Ien VGND 0.37345f
C4372 XA.XIR[6].XIC[7].icell.Ien VGND 0.37345f
C4373 XA.XIR[6].XIC[6].icell.Ien VGND 0.37345f
C4374 XA.XIR[6].XIC[5].icell.Ien VGND 0.37345f
C4375 XA.XIR[6].XIC[4].icell.Ien VGND 0.37345f
C4376 XA.XIR[6].XIC[3].icell.Ien VGND 0.37345f
C4377 XA.XIR[6].XIC[2].icell.Ien VGND 0.37345f
C4378 XA.XIR[6].XIC_dummy_left.icell.Iout VGND 0.80729f
C4379 XA.XIR[6].XIC[1].icell.Ien VGND 0.37345f
C4380 XA.XIR[6].XIC[0].icell.Ien VGND 0.37359f
C4381 XA.XIR[6].XIC_dummy_left.icell.SM VGND 0.01044f
C4382 XA.XIR[6].XIC_dummy_left.icell.Ien VGND 0.57425f
C4383 XThR.Tn[6] VGND 13.26097f
C4384 a_n1049_5317# VGND 0.02283f
C4385 XThR.XTB7.Y VGND 1.36132f
C4386 XA.XIR[6].XIC_dummy_right.icell.PDM VGND 0.23384f
C4387 XA.XIR[6].XIC_15.icell.PDM VGND 0.18862f
C4388 XA.XIR[6].XIC[14].icell.PDM VGND 0.18817f
C4389 XA.XIR[6].XIC[13].icell.PDM VGND 0.18817f
C4390 XA.XIR[6].XIC[12].icell.PDM VGND 0.18817f
C4391 XA.XIR[6].XIC[11].icell.PDM VGND 0.18817f
C4392 XA.XIR[6].XIC[10].icell.PDM VGND 0.18817f
C4393 XA.XIR[6].XIC[9].icell.PDM VGND 0.18817f
C4394 XA.XIR[6].XIC[8].icell.PDM VGND 0.18817f
C4395 XA.XIR[6].XIC[7].icell.PDM VGND 0.18817f
C4396 XA.XIR[6].XIC[6].icell.PDM VGND 0.18817f
C4397 XA.XIR[6].XIC[5].icell.PDM VGND 0.18817f
C4398 XA.XIR[6].XIC[4].icell.PDM VGND 0.18817f
C4399 XA.XIR[6].XIC[3].icell.PDM VGND 0.18817f
C4400 XA.XIR[6].XIC[2].icell.PDM VGND 0.18817f
C4401 XA.XIR[6].XIC[1].icell.PDM VGND 0.18817f
C4402 XA.XIR[6].XIC[0].icell.PDM VGND 0.18824f
C4403 XA.XIR[6].XIC_dummy_left.icell.PDM VGND 0.22809f
C4404 XA.XIR[5].XIC_dummy_right.icell.Iout VGND 0.85788f
C4405 XA.XIR[5].XIC_dummy_right.icell.SM VGND 0.01013f
C4406 XA.XIR[5].XIC_dummy_right.icell.Ien VGND 0.60818f
C4407 XA.XIR[5].XIC_15.icell.Ien VGND 0.37264f
C4408 XA.XIR[5].XIC[14].icell.Ien VGND 0.37345f
C4409 XA.XIR[5].XIC[13].icell.Ien VGND 0.37345f
C4410 XA.XIR[5].XIC[12].icell.Ien VGND 0.37345f
C4411 XA.XIR[5].XIC[11].icell.Ien VGND 0.37345f
C4412 XA.XIR[5].XIC[10].icell.Ien VGND 0.37345f
C4413 XA.XIR[5].XIC[9].icell.Ien VGND 0.37345f
C4414 XA.XIR[5].XIC[8].icell.Ien VGND 0.37345f
C4415 XA.XIR[5].XIC[7].icell.Ien VGND 0.37345f
C4416 XA.XIR[5].XIC[6].icell.Ien VGND 0.37345f
C4417 XA.XIR[5].XIC[5].icell.Ien VGND 0.37345f
C4418 XA.XIR[5].XIC[4].icell.Ien VGND 0.37345f
C4419 XA.XIR[5].XIC[3].icell.Ien VGND 0.37345f
C4420 XA.XIR[5].XIC[2].icell.Ien VGND 0.37345f
C4421 XA.XIR[5].XIC_dummy_left.icell.Iout VGND 0.80598f
C4422 XA.XIR[5].XIC[1].icell.Ien VGND 0.37345f
C4423 a_n1049_5611# VGND 0.02888f
C4424 XA.XIR[5].XIC[0].icell.Ien VGND 0.37359f
C4425 XA.XIR[5].XIC_dummy_left.icell.SM VGND 0.01044f
C4426 XA.XIR[5].XIC_dummy_left.icell.Ien VGND 0.57291f
C4427 XThR.Tn[5] VGND 13.28746f
C4428 XThR.XTB6.Y VGND 1.38212f
C4429 XA.XIR[5].XIC_dummy_right.icell.PDM VGND 0.23384f
C4430 XA.XIR[5].XIC_15.icell.PDM VGND 0.18862f
C4431 XA.XIR[5].XIC[14].icell.PDM VGND 0.18817f
C4432 XA.XIR[5].XIC[13].icell.PDM VGND 0.18817f
C4433 XA.XIR[5].XIC[12].icell.PDM VGND 0.18817f
C4434 XA.XIR[5].XIC[11].icell.PDM VGND 0.18817f
C4435 XA.XIR[5].XIC[10].icell.PDM VGND 0.18817f
C4436 XA.XIR[5].XIC[9].icell.PDM VGND 0.18817f
C4437 XA.XIR[5].XIC[8].icell.PDM VGND 0.18817f
C4438 XA.XIR[5].XIC[7].icell.PDM VGND 0.18817f
C4439 XA.XIR[5].XIC[6].icell.PDM VGND 0.18817f
C4440 XA.XIR[5].XIC[5].icell.PDM VGND 0.18817f
C4441 XA.XIR[5].XIC[4].icell.PDM VGND 0.18817f
C4442 XA.XIR[5].XIC[3].icell.PDM VGND 0.18817f
C4443 XA.XIR[5].XIC[2].icell.PDM VGND 0.18817f
C4444 XA.XIR[5].XIC[1].icell.PDM VGND 0.18817f
C4445 XA.XIR[5].XIC[0].icell.PDM VGND 0.18824f
C4446 XA.XIR[5].XIC_dummy_left.icell.PDM VGND 0.22809f
C4447 XA.XIR[4].XIC_dummy_right.icell.Iout VGND 0.85788f
C4448 XA.XIR[4].XIC_dummy_right.icell.SM VGND 0.01013f
C4449 XA.XIR[4].XIC_dummy_right.icell.Ien VGND 0.60818f
C4450 XA.XIR[4].XIC_15.icell.Ien VGND 0.37264f
C4451 XA.XIR[4].XIC[14].icell.Ien VGND 0.37345f
C4452 XA.XIR[4].XIC[13].icell.Ien VGND 0.37345f
C4453 XA.XIR[4].XIC[12].icell.Ien VGND 0.37345f
C4454 XA.XIR[4].XIC[11].icell.Ien VGND 0.37345f
C4455 XA.XIR[4].XIC[10].icell.Ien VGND 0.37345f
C4456 XA.XIR[4].XIC[9].icell.Ien VGND 0.37345f
C4457 XA.XIR[4].XIC[8].icell.Ien VGND 0.37345f
C4458 XA.XIR[4].XIC[7].icell.Ien VGND 0.37345f
C4459 XA.XIR[4].XIC[6].icell.Ien VGND 0.37345f
C4460 XA.XIR[4].XIC[5].icell.Ien VGND 0.37345f
C4461 XA.XIR[4].XIC[4].icell.Ien VGND 0.37345f
C4462 XA.XIR[4].XIC[3].icell.Ien VGND 0.37345f
C4463 XA.XIR[4].XIC[2].icell.Ien VGND 0.37345f
C4464 XA.XIR[4].XIC_dummy_left.icell.Iout VGND 0.8077f
C4465 XA.XIR[4].XIC[1].icell.Ien VGND 0.37345f
C4466 XA.XIR[4].XIC[0].icell.Ien VGND 0.37359f
C4467 XA.XIR[4].XIC_dummy_left.icell.SM VGND 0.01044f
C4468 XA.XIR[4].XIC_dummy_left.icell.Ien VGND 0.57336f
C4469 XA.XIR[4].XIC_dummy_right.icell.PDM VGND 0.23384f
C4470 XA.XIR[4].XIC_15.icell.PDM VGND 0.18862f
C4471 XA.XIR[4].XIC[14].icell.PDM VGND 0.18817f
C4472 XA.XIR[4].XIC[13].icell.PDM VGND 0.18817f
C4473 XA.XIR[4].XIC[12].icell.PDM VGND 0.18817f
C4474 XA.XIR[4].XIC[11].icell.PDM VGND 0.18817f
C4475 XA.XIR[4].XIC[10].icell.PDM VGND 0.18817f
C4476 XA.XIR[4].XIC[9].icell.PDM VGND 0.18817f
C4477 XA.XIR[4].XIC[8].icell.PDM VGND 0.18817f
C4478 XA.XIR[4].XIC[7].icell.PDM VGND 0.18817f
C4479 XA.XIR[4].XIC[6].icell.PDM VGND 0.18817f
C4480 XA.XIR[4].XIC[5].icell.PDM VGND 0.18817f
C4481 XA.XIR[4].XIC[4].icell.PDM VGND 0.18817f
C4482 XA.XIR[4].XIC[3].icell.PDM VGND 0.18817f
C4483 XA.XIR[4].XIC[2].icell.PDM VGND 0.18817f
C4484 XA.XIR[4].XIC[1].icell.PDM VGND 0.18817f
C4485 XA.XIR[4].XIC[0].icell.PDM VGND 0.18824f
C4486 XA.XIR[4].XIC_dummy_left.icell.PDM VGND 0.22809f
C4487 XThR.Tn[4] VGND 13.34854f
C4488 a_n1049_6405# VGND 0.02935f
C4489 XA.XIR[3].XIC_dummy_right.icell.Iout VGND 0.85788f
C4490 XA.XIR[3].XIC_dummy_right.icell.SM VGND 0.01013f
C4491 XA.XIR[3].XIC_dummy_right.icell.Ien VGND 0.60818f
C4492 XA.XIR[3].XIC_15.icell.Ien VGND 0.37264f
C4493 XA.XIR[3].XIC[14].icell.Ien VGND 0.37345f
C4494 XA.XIR[3].XIC[13].icell.Ien VGND 0.37345f
C4495 XA.XIR[3].XIC[12].icell.Ien VGND 0.37345f
C4496 XA.XIR[3].XIC[11].icell.Ien VGND 0.37345f
C4497 XA.XIR[3].XIC[10].icell.Ien VGND 0.37345f
C4498 XA.XIR[3].XIC[9].icell.Ien VGND 0.37345f
C4499 XA.XIR[3].XIC[8].icell.Ien VGND 0.37345f
C4500 XA.XIR[3].XIC[7].icell.Ien VGND 0.37345f
C4501 XA.XIR[3].XIC[6].icell.Ien VGND 0.37345f
C4502 XA.XIR[3].XIC[5].icell.Ien VGND 0.37345f
C4503 XA.XIR[3].XIC[4].icell.Ien VGND 0.37345f
C4504 XA.XIR[3].XIC[3].icell.Ien VGND 0.37345f
C4505 XA.XIR[3].XIC[2].icell.Ien VGND 0.37345f
C4506 XThR.XTB5.Y VGND 1.32753f
C4507 XA.XIR[3].XIC_dummy_left.icell.Iout VGND 0.80611f
C4508 XA.XIR[3].XIC[1].icell.Ien VGND 0.37345f
C4509 XA.XIR[3].XIC[0].icell.Ien VGND 0.37359f
C4510 XA.XIR[3].XIC_dummy_left.icell.SM VGND 0.01044f
C4511 XA.XIR[3].XIC_dummy_left.icell.Ien VGND 0.57425f
C4512 a_n1049_6699# VGND 0.02979f
C4513 XA.XIR[3].XIC_dummy_right.icell.PDM VGND 0.23384f
C4514 XA.XIR[3].XIC_15.icell.PDM VGND 0.18862f
C4515 XA.XIR[3].XIC[14].icell.PDM VGND 0.18817f
C4516 XA.XIR[3].XIC[13].icell.PDM VGND 0.18817f
C4517 XA.XIR[3].XIC[12].icell.PDM VGND 0.18817f
C4518 XA.XIR[3].XIC[11].icell.PDM VGND 0.18817f
C4519 XA.XIR[3].XIC[10].icell.PDM VGND 0.18817f
C4520 XA.XIR[3].XIC[9].icell.PDM VGND 0.18817f
C4521 XA.XIR[3].XIC[8].icell.PDM VGND 0.18817f
C4522 XA.XIR[3].XIC[7].icell.PDM VGND 0.18817f
C4523 XA.XIR[3].XIC[6].icell.PDM VGND 0.18817f
C4524 XA.XIR[3].XIC[5].icell.PDM VGND 0.18817f
C4525 XA.XIR[3].XIC[4].icell.PDM VGND 0.18817f
C4526 XA.XIR[3].XIC[3].icell.PDM VGND 0.18817f
C4527 XA.XIR[3].XIC[2].icell.PDM VGND 0.18817f
C4528 XA.XIR[3].XIC[1].icell.PDM VGND 0.18817f
C4529 XA.XIR[3].XIC[0].icell.PDM VGND 0.18824f
C4530 XA.XIR[3].XIC_dummy_left.icell.PDM VGND 0.22809f
C4531 XA.XIR[2].XIC_dummy_right.icell.Iout VGND 0.85788f
C4532 XA.XIR[2].XIC_dummy_right.icell.SM VGND 0.01013f
C4533 XA.XIR[2].XIC_dummy_right.icell.Ien VGND 0.60818f
C4534 XA.XIR[2].XIC_15.icell.Ien VGND 0.37264f
C4535 XA.XIR[2].XIC[14].icell.Ien VGND 0.37345f
C4536 XA.XIR[2].XIC[13].icell.Ien VGND 0.37345f
C4537 XA.XIR[2].XIC[12].icell.Ien VGND 0.37345f
C4538 XA.XIR[2].XIC[11].icell.Ien VGND 0.37345f
C4539 XA.XIR[2].XIC[10].icell.Ien VGND 0.37345f
C4540 XA.XIR[2].XIC[9].icell.Ien VGND 0.37345f
C4541 XA.XIR[2].XIC[8].icell.Ien VGND 0.37345f
C4542 XA.XIR[2].XIC[7].icell.Ien VGND 0.37345f
C4543 XA.XIR[2].XIC[6].icell.Ien VGND 0.37345f
C4544 XA.XIR[2].XIC[5].icell.Ien VGND 0.37345f
C4545 XA.XIR[2].XIC[4].icell.Ien VGND 0.37345f
C4546 XA.XIR[2].XIC[3].icell.Ien VGND 0.37345f
C4547 XA.XIR[2].XIC[2].icell.Ien VGND 0.37345f
C4548 XA.XIR[2].XIC_dummy_left.icell.Iout VGND 0.80825f
C4549 XA.XIR[2].XIC[1].icell.Ien VGND 0.37345f
C4550 XThR.Tn[3] VGND 13.30321f
C4551 XThR.XTB4.Y VGND 1.76953f
C4552 XA.XIR[2].XIC[0].icell.Ien VGND 0.37359f
C4553 XA.XIR[2].XIC_dummy_left.icell.SM VGND 0.01044f
C4554 XA.XIR[2].XIC_dummy_left.icell.Ien VGND 0.57559f
C4555 XA.XIR[2].XIC_dummy_right.icell.PDM VGND 0.23384f
C4556 XA.XIR[2].XIC_15.icell.PDM VGND 0.18862f
C4557 XA.XIR[2].XIC[14].icell.PDM VGND 0.18817f
C4558 XA.XIR[2].XIC[13].icell.PDM VGND 0.18817f
C4559 XA.XIR[2].XIC[12].icell.PDM VGND 0.18817f
C4560 XA.XIR[2].XIC[11].icell.PDM VGND 0.18817f
C4561 XA.XIR[2].XIC[10].icell.PDM VGND 0.18817f
C4562 XA.XIR[2].XIC[9].icell.PDM VGND 0.18817f
C4563 XA.XIR[2].XIC[8].icell.PDM VGND 0.18817f
C4564 XA.XIR[2].XIC[7].icell.PDM VGND 0.18817f
C4565 XA.XIR[2].XIC[6].icell.PDM VGND 0.18817f
C4566 XA.XIR[2].XIC[5].icell.PDM VGND 0.18817f
C4567 XA.XIR[2].XIC[4].icell.PDM VGND 0.18817f
C4568 XA.XIR[2].XIC[3].icell.PDM VGND 0.18817f
C4569 XA.XIR[2].XIC[2].icell.PDM VGND 0.18817f
C4570 XA.XIR[2].XIC[1].icell.PDM VGND 0.18817f
C4571 XA.XIR[2].XIC[0].icell.PDM VGND 0.18824f
C4572 XA.XIR[2].XIC_dummy_left.icell.PDM VGND 0.22809f
C4573 XA.XIR[1].XIC_dummy_right.icell.Iout VGND 0.85788f
C4574 XA.XIR[1].XIC_dummy_right.icell.SM VGND 0.01013f
C4575 XA.XIR[1].XIC_dummy_right.icell.Ien VGND 0.60818f
C4576 XA.XIR[1].XIC_15.icell.Ien VGND 0.37264f
C4577 XA.XIR[1].XIC[14].icell.Ien VGND 0.37345f
C4578 XA.XIR[1].XIC[13].icell.Ien VGND 0.37345f
C4579 XA.XIR[1].XIC[12].icell.Ien VGND 0.37345f
C4580 XA.XIR[1].XIC[11].icell.Ien VGND 0.37345f
C4581 XA.XIR[1].XIC[10].icell.Ien VGND 0.37345f
C4582 XA.XIR[1].XIC[9].icell.Ien VGND 0.37345f
C4583 XA.XIR[1].XIC[8].icell.Ien VGND 0.37345f
C4584 XA.XIR[1].XIC[7].icell.Ien VGND 0.37345f
C4585 XA.XIR[1].XIC[6].icell.Ien VGND 0.37345f
C4586 XA.XIR[1].XIC[5].icell.Ien VGND 0.37345f
C4587 XA.XIR[1].XIC[4].icell.Ien VGND 0.37345f
C4588 XA.XIR[1].XIC[3].icell.Ien VGND 0.37345f
C4589 XA.XIR[1].XIC[2].icell.Ien VGND 0.37345f
C4590 XA.XIR[1].XIC_dummy_left.icell.Iout VGND 0.80611f
C4591 XA.XIR[1].XIC[1].icell.Ien VGND 0.37345f
C4592 XThR.Tn[2] VGND 13.34591f
C4593 a_n1049_7493# VGND 0.02484f
C4594 XThR.XTB3.Y VGND 2.09162f
C4595 XThR.XTB7.A VGND 1.95537f
C4596 XA.XIR[1].XIC[0].icell.Ien VGND 0.37359f
C4597 XA.XIR[1].XIC_dummy_left.icell.SM VGND 0.01044f
C4598 XA.XIR[1].XIC_dummy_left.icell.Ien VGND 0.57379f
C4599 XA.XIR[1].XIC_dummy_right.icell.PDM VGND 0.23384f
C4600 XA.XIR[1].XIC_15.icell.PDM VGND 0.18862f
C4601 XA.XIR[1].XIC[14].icell.PDM VGND 0.18817f
C4602 XA.XIR[1].XIC[13].icell.PDM VGND 0.18817f
C4603 XA.XIR[1].XIC[12].icell.PDM VGND 0.18817f
C4604 XA.XIR[1].XIC[11].icell.PDM VGND 0.18817f
C4605 XA.XIR[1].XIC[10].icell.PDM VGND 0.18817f
C4606 XA.XIR[1].XIC[9].icell.PDM VGND 0.18817f
C4607 XA.XIR[1].XIC[8].icell.PDM VGND 0.18817f
C4608 XA.XIR[1].XIC[7].icell.PDM VGND 0.18817f
C4609 XA.XIR[1].XIC[6].icell.PDM VGND 0.18817f
C4610 XA.XIR[1].XIC[5].icell.PDM VGND 0.18817f
C4611 XA.XIR[1].XIC[4].icell.PDM VGND 0.18817f
C4612 XA.XIR[1].XIC[3].icell.PDM VGND 0.18817f
C4613 XA.XIR[1].XIC[2].icell.PDM VGND 0.18817f
C4614 XA.XIR[1].XIC[1].icell.PDM VGND 0.18817f
C4615 XA.XIR[1].XIC[0].icell.PDM VGND 0.18824f
C4616 XA.XIR[1].XIC_dummy_left.icell.PDM VGND 0.22809f
C4617 a_n1049_7787# VGND 0.03397f
C4618 XA.XIR[0].XIC_dummy_right.icell.Iout VGND 0.87403f
C4619 XA.XIR[0].XIC_dummy_right.icell.SM VGND 0.01013f
C4620 XA.XIR[0].XIC_dummy_right.icell.Ien VGND 0.61797f
C4621 XA.XIR[0].XIC_15.icell.Ien VGND 0.37874f
C4622 XA.XIR[0].XIC[14].icell.Ien VGND 0.39188f
C4623 XA.XIR[0].XIC[13].icell.Ien VGND 0.39193f
C4624 XA.XIR[0].XIC[12].icell.Ien VGND 0.38856f
C4625 XA.XIR[0].XIC[11].icell.Ien VGND 0.38923f
C4626 XA.XIR[0].XIC[10].icell.Ien VGND 0.39057f
C4627 XA.XIR[0].XIC[9].icell.Ien VGND 0.38884f
C4628 XA.XIR[0].XIC[8].icell.Ien VGND 0.38932f
C4629 XA.XIR[0].XIC[7].icell.Ien VGND 0.38956f
C4630 XA.XIR[0].XIC[6].icell.Ien VGND 0.38948f
C4631 XA.XIR[0].XIC[5].icell.Ien VGND 0.38847f
C4632 XA.XIR[0].XIC[4].icell.Ien VGND 0.38861f
C4633 XA.XIR[0].XIC[3].icell.Ien VGND 0.38986f
C4634 XA.XIR[0].XIC[2].icell.Ien VGND 0.39188f
C4635 XA.XIR[0].XIC_dummy_left.icell.Iout VGND 0.83227f
C4636 XA.XIR[0].XIC[1].icell.Ien VGND 0.39188f
C4637 XA.XIR[0].XIC[0].icell.Ien VGND 0.39129f
C4638 XA.XIR[0].XIC_dummy_left.icell.SM VGND 0.01044f
C4639 XThR.Tn[1] VGND 13.34734f
C4640 XThR.XTB2.Y VGND 1.47619f
C4641 XThR.XTB6.A VGND 0.95635f
C4642 XA.XIR[0].XIC_dummy_left.icell.Ien VGND 0.58434f
C4643 XA.XIR[0].XIC_dummy_right.icell.PDM VGND 0.251f
C4644 XA.XIR[0].XIC_15.icell.PDM VGND 0.20773f
C4645 XA.XIR[0].XIC[14].icell.PDM VGND 0.24611f
C4646 XA.XIR[0].XIC[13].icell.PDM VGND 0.24595f
C4647 XA.XIR[0].XIC[12].icell.PDM VGND 0.24156f
C4648 XA.XIR[0].XIC[11].icell.PDM VGND 0.24193f
C4649 XA.XIR[0].XIC[10].icell.PDM VGND 0.24184f
C4650 XA.XIR[0].XIC[9].icell.PDM VGND 0.24156f
C4651 XA.XIR[0].XIC[8].icell.PDM VGND 0.24156f
C4652 XA.XIR[0].XIC[7].icell.PDM VGND 0.244f
C4653 XA.XIR[0].XIC[6].icell.PDM VGND 0.2412f
C4654 XA.XIR[0].XIC[5].icell.PDM VGND 0.24309f
C4655 XA.XIR[0].XIC[4].icell.PDM VGND 0.24168f
C4656 XA.XIR[0].XIC[3].icell.PDM VGND 0.24467f
C4657 XA.XIR[0].XIC[2].icell.PDM VGND 0.2459f
C4658 XA.XIR[0].XIC[1].icell.PDM VGND 0.2459f
C4659 XA.XIR[0].XIC[0].icell.PDM VGND 0.24468f
C4660 XA.XIR[0].XIC_dummy_left.icell.PDM VGND 0.24577f
C4661 XThR.Tn[0] VGND 13.64913f
C4662 a_n1049_8581# VGND 0.04333f
C4663 XThR.XTBN.Y VGND 7.54415f
C4664 XThR.XTB1.Y VGND 1.80911f
C4665 XThR.XTB7.B VGND 2.61063f
C4666 XThR.XTB5.A VGND 1.75777f
C4667 XThC.Tn[14] VGND 9.53729f
C4668 XThC.Tn[13] VGND 9.34297f
C4669 XThC.Tn[12] VGND 9.16726f
C4670 XThC.Tn[11] VGND 9.0184f
C4671 XThC.Tn[10] VGND 8.90983f
C4672 XThC.Tn[9] VGND 8.91295f
C4673 XThC.Tn[8] VGND 8.89302f
C4674 a_10915_9569# VGND 0.55837f
C4675 a_10051_9569# VGND 0.55761f
C4676 a_9827_9569# VGND 0.54461f
C4677 a_8963_9569# VGND 0.55448f
C4678 a_8739_9569# VGND 0.55288f
C4679 a_7875_9569# VGND 0.55432f
C4680 a_7651_9569# VGND 0.55717f
C4681 XThC.Tn[7] VGND 10.0223f
C4682 XThC.Tn[6] VGND 9.91412f
C4683 XThC.Tn[5] VGND 10.12609f
C4684 XThC.Tn[4] VGND 10.07042f
C4685 XThC.Tn[3] VGND 9.50738f
C4686 XThC.Tn[2] VGND 9.91895f
C4687 XThC.Tn[1] VGND 10.12244f
C4688 XThC.Tn[0] VGND 10.70185f
C4689 a_6243_9615# VGND 0.0299f
C4690 a_5949_9615# VGND 0.03432f
C4691 a_5155_9615# VGND 0.03615f
C4692 a_4861_9615# VGND 0.03632f
C4693 a_4067_9615# VGND 0.03071f
C4694 a_3773_9615# VGND 0.03867f
C4695 a_2979_9615# VGND 0.04044f
C4696 XThC.XTBN.Y VGND 7.90366f
C4697 XThC.XTB7.Y VGND 1.36247f
C4698 XThC.XTB6.Y VGND 1.3829f
C4699 XThC.XTB7.B VGND 2.73055f
C4700 XThC.XTB5.Y VGND 1.32591f
C4701 XThC.XTBN.A VGND 1.23171f
C4702 XThC.XTB4.Y VGND 1.69875f
C4703 XThC.XTB3.Y VGND 1.96765f
C4704 XThC.XTB7.A VGND 1.96056f
C4705 XThC.XTB6.A VGND 0.95757f
C4706 XThC.XTB2.Y VGND 1.47589f
C4707 XThC.XTB1.Y VGND 1.77676f
C4708 XThC.XTB5.A VGND 1.75974f
C4709 bias[0].t0 VGND 0.94587f
C4710 XThR.XTB3.Y.t1 VGND 0.06176f
C4711 XThR.XTB3.Y.n0 VGND 0.01521f
C4712 XThR.XTB3.Y.t8 VGND 0.04903f
C4713 XThR.XTB3.Y.t15 VGND 0.02889f
C4714 XThR.XTB3.Y.t13 VGND 0.04903f
C4715 XThR.XTB3.Y.t6 VGND 0.02889f
C4716 XThR.XTB3.Y.t9 VGND 0.04903f
C4717 XThR.XTB3.Y.t17 VGND 0.02889f
C4718 XThR.XTB3.Y.n1 VGND 0.08226f
C4719 XThR.XTB3.Y.n2 VGND 0.08688f
C4720 XThR.XTB3.Y.n3 VGND 0.03573f
C4721 XThR.XTB3.Y.n4 VGND 0.0707f
C4722 XThR.XTB3.Y.t12 VGND 0.04903f
C4723 XThR.XTB3.Y.t4 VGND 0.02889f
C4724 XThR.XTB3.Y.n5 VGND 0.06608f
C4725 XThR.XTB3.Y.n6 VGND 0.03236f
C4726 XThR.XTB3.Y.n7 VGND 0.02685f
C4727 XThR.XTB3.Y.t18 VGND 0.04903f
C4728 XThR.XTB3.Y.t5 VGND 0.02889f
C4729 XThR.XTB3.Y.n8 VGND 0.03005f
C4730 XThR.XTB3.Y.t7 VGND 0.04903f
C4731 XThR.XTB3.Y.t10 VGND 0.02889f
C4732 XThR.XTB3.Y.n9 VGND 0.05992f
C4733 XThR.XTB3.Y.t11 VGND 0.04903f
C4734 XThR.XTB3.Y.t16 VGND 0.02889f
C4735 XThR.XTB3.Y.n10 VGND 0.06454f
C4736 XThR.XTB3.Y.n11 VGND 0.03645f
C4737 XThR.XTB3.Y.n12 VGND 0.06034f
C4738 XThR.XTB3.Y.n13 VGND 0.03128f
C4739 XThR.XTB3.Y.n14 VGND 0.02851f
C4740 XThR.XTB3.Y.n15 VGND 0.06454f
C4741 XThR.XTB3.Y.t14 VGND 0.04903f
C4742 XThR.XTB3.Y.t3 VGND 0.02889f
C4743 XThR.XTB3.Y.n16 VGND 0.05838f
C4744 XThR.XTB3.Y.n17 VGND 0.03236f
C4745 XThR.XTB3.Y.n18 VGND 0.04707f
C4746 XThR.XTB3.Y.n19 VGND 1.31347f
C4747 XThR.XTB3.Y.t2 VGND 0.03152f
C4748 XThR.XTB3.Y.t0 VGND 0.03152f
C4749 XThR.XTB3.Y.n20 VGND 0.06766f
C4750 XThR.XTB3.Y.n21 VGND 0.157f
C4751 XThR.XTB3.Y.n22 VGND 0.03296f
C4752 XThR.XTB1.Y.t1 VGND 0.03165f
C4753 XThR.XTB1.Y.t8 VGND 0.02512f
C4754 XThR.XTB1.Y.t15 VGND 0.0148f
C4755 XThR.XTB1.Y.t14 VGND 0.02512f
C4756 XThR.XTB1.Y.t7 VGND 0.0148f
C4757 XThR.XTB1.Y.t10 VGND 0.02512f
C4758 XThR.XTB1.Y.t18 VGND 0.0148f
C4759 XThR.XTB1.Y.n1 VGND 0.04215f
C4760 XThR.XTB1.Y.n2 VGND 0.04452f
C4761 XThR.XTB1.Y.n3 VGND 0.01831f
C4762 XThR.XTB1.Y.n4 VGND 0.03623f
C4763 XThR.XTB1.Y.t13 VGND 0.02512f
C4764 XThR.XTB1.Y.t4 VGND 0.0148f
C4765 XThR.XTB1.Y.n5 VGND 0.03386f
C4766 XThR.XTB1.Y.n6 VGND 0.01658f
C4767 XThR.XTB1.Y.n7 VGND 0.01376f
C4768 XThR.XTB1.Y.t6 VGND 0.02512f
C4769 XThR.XTB1.Y.t11 VGND 0.0148f
C4770 XThR.XTB1.Y.n8 VGND 0.0154f
C4771 XThR.XTB1.Y.t12 VGND 0.02512f
C4772 XThR.XTB1.Y.t16 VGND 0.0148f
C4773 XThR.XTB1.Y.n9 VGND 0.0307f
C4774 XThR.XTB1.Y.t17 VGND 0.02512f
C4775 XThR.XTB1.Y.t5 VGND 0.0148f
C4776 XThR.XTB1.Y.n10 VGND 0.03307f
C4777 XThR.XTB1.Y.n11 VGND 0.01868f
C4778 XThR.XTB1.Y.n12 VGND 0.03092f
C4779 XThR.XTB1.Y.n13 VGND 0.01603f
C4780 XThR.XTB1.Y.n14 VGND 0.01461f
C4781 XThR.XTB1.Y.n15 VGND 0.03307f
C4782 XThR.XTB1.Y.t3 VGND 0.02512f
C4783 XThR.XTB1.Y.t9 VGND 0.0148f
C4784 XThR.XTB1.Y.n16 VGND 0.02991f
C4785 XThR.XTB1.Y.n17 VGND 0.01658f
C4786 XThR.XTB1.Y.n18 VGND 0.02412f
C4787 XThR.XTB1.Y.n19 VGND 0.75219f
C4788 XThR.XTB1.Y.t2 VGND 0.01615f
C4789 XThR.XTB1.Y.t0 VGND 0.01615f
C4790 XThR.XTB1.Y.n20 VGND 0.03467f
C4791 XThR.XTB1.Y.n21 VGND 0.08068f
C4792 XThR.XTB1.Y.n22 VGND 0.01689f
C4793 XThR.XTB4.Y.t8 VGND 0.02956f
C4794 XThR.XTB4.Y.t15 VGND 0.05016f
C4795 XThR.XTB4.Y.t16 VGND 0.02956f
C4796 XThR.XTB4.Y.t5 VGND 0.05016f
C4797 XThR.XTB4.Y.t10 VGND 0.02956f
C4798 XThR.XTB4.Y.t17 VGND 0.05016f
C4799 XThR.XTB4.Y.n0 VGND 0.08416f
C4800 XThR.XTB4.Y.n1 VGND 0.08889f
C4801 XThR.XTB4.Y.n2 VGND 0.03656f
C4802 XThR.XTB4.Y.n3 VGND 0.07234f
C4803 XThR.XTB4.Y.t13 VGND 0.02956f
C4804 XThR.XTB4.Y.t4 VGND 0.05016f
C4805 XThR.XTB4.Y.n4 VGND 0.06761f
C4806 XThR.XTB4.Y.n5 VGND 0.0331f
C4807 XThR.XTB4.Y.n6 VGND 0.01685f
C4808 XThR.XTB4.Y.n7 VGND 0.05355f
C4809 XThR.XTB4.Y.n8 VGND 0.64921f
C4810 XThR.XTB4.Y.t14 VGND 0.02956f
C4811 XThR.XTB4.Y.t7 VGND 0.05016f
C4812 XThR.XTB4.Y.n9 VGND 0.03074f
C4813 XThR.XTB4.Y.t3 VGND 0.02956f
C4814 XThR.XTB4.Y.t12 VGND 0.05016f
C4815 XThR.XTB4.Y.n10 VGND 0.0613f
C4816 XThR.XTB4.Y.t9 VGND 0.02956f
C4817 XThR.XTB4.Y.t2 VGND 0.05016f
C4818 XThR.XTB4.Y.n11 VGND 0.06603f
C4819 XThR.XTB4.Y.n12 VGND 0.03729f
C4820 XThR.XTB4.Y.n13 VGND 0.06174f
C4821 XThR.XTB4.Y.n14 VGND 0.03201f
C4822 XThR.XTB4.Y.n15 VGND 0.02916f
C4823 XThR.XTB4.Y.n16 VGND 0.06603f
C4824 XThR.XTB4.Y.t11 VGND 0.02956f
C4825 XThR.XTB4.Y.t6 VGND 0.05016f
C4826 XThR.XTB4.Y.n17 VGND 0.05972f
C4827 XThR.XTB4.Y.n18 VGND 0.0331f
C4828 XThR.XTB4.Y.n19 VGND 0.05647f
C4829 XThR.XTB4.Y.n20 VGND 1.3092f
C4830 XThR.XTB4.Y.t1 VGND 0.06491f
C4831 XThR.XTB4.Y.n21 VGND 0.12281f
C4832 XThR.XTB4.Y.n22 VGND 0.02892f
C4833 XThR.XTB4.Y.t0 VGND 0.11919f
C4834 XThR.Tn[13].t9 VGND 0.01972f
C4835 XThR.Tn[13].t11 VGND 0.01972f
C4836 XThR.Tn[13].n0 VGND 0.05989f
C4837 XThR.Tn[13].t10 VGND 0.01972f
C4838 XThR.Tn[13].t8 VGND 0.01972f
C4839 XThR.Tn[13].n1 VGND 0.04385f
C4840 XThR.Tn[13].n2 VGND 0.19937f
C4841 XThR.Tn[13].t7 VGND 0.01282f
C4842 XThR.Tn[13].t5 VGND 0.01282f
C4843 XThR.Tn[13].n3 VGND 0.03198f
C4844 XThR.Tn[13].t6 VGND 0.01282f
C4845 XThR.Tn[13].t4 VGND 0.01282f
C4846 XThR.Tn[13].n4 VGND 0.02564f
C4847 XThR.Tn[13].n5 VGND 0.0645f
C4848 XThR.Tn[13].t72 VGND 0.01542f
C4849 XThR.Tn[13].t64 VGND 0.01688f
C4850 XThR.Tn[13].n6 VGND 0.04122f
C4851 XThR.Tn[13].n7 VGND 0.07918f
C4852 XThR.Tn[13].t28 VGND 0.01542f
C4853 XThR.Tn[13].t21 VGND 0.01688f
C4854 XThR.Tn[13].n8 VGND 0.04122f
C4855 XThR.Tn[13].t44 VGND 0.01536f
C4856 XThR.Tn[13].t12 VGND 0.01683f
C4857 XThR.Tn[13].n9 VGND 0.04289f
C4858 XThR.Tn[13].n10 VGND 0.03013f
C4859 XThR.Tn[13].n12 VGND 0.09669f
C4860 XThR.Tn[13].t65 VGND 0.01542f
C4861 XThR.Tn[13].t57 VGND 0.01688f
C4862 XThR.Tn[13].n13 VGND 0.04122f
C4863 XThR.Tn[13].t19 VGND 0.01536f
C4864 XThR.Tn[13].t52 VGND 0.01683f
C4865 XThR.Tn[13].n14 VGND 0.04289f
C4866 XThR.Tn[13].n15 VGND 0.03013f
C4867 XThR.Tn[13].n17 VGND 0.09669f
C4868 XThR.Tn[13].t22 VGND 0.01542f
C4869 XThR.Tn[13].t14 VGND 0.01688f
C4870 XThR.Tn[13].n18 VGND 0.04122f
C4871 XThR.Tn[13].t34 VGND 0.01536f
C4872 XThR.Tn[13].t70 VGND 0.01683f
C4873 XThR.Tn[13].n19 VGND 0.04289f
C4874 XThR.Tn[13].n20 VGND 0.03013f
C4875 XThR.Tn[13].n22 VGND 0.09669f
C4876 XThR.Tn[13].t49 VGND 0.01542f
C4877 XThR.Tn[13].t39 VGND 0.01688f
C4878 XThR.Tn[13].n23 VGND 0.04122f
C4879 XThR.Tn[13].t66 VGND 0.01536f
C4880 XThR.Tn[13].t35 VGND 0.01683f
C4881 XThR.Tn[13].n24 VGND 0.04289f
C4882 XThR.Tn[13].n25 VGND 0.03013f
C4883 XThR.Tn[13].n27 VGND 0.09669f
C4884 XThR.Tn[13].t24 VGND 0.01542f
C4885 XThR.Tn[13].t16 VGND 0.01688f
C4886 XThR.Tn[13].n28 VGND 0.04122f
C4887 XThR.Tn[13].t37 VGND 0.01536f
C4888 XThR.Tn[13].t71 VGND 0.01683f
C4889 XThR.Tn[13].n29 VGND 0.04289f
C4890 XThR.Tn[13].n30 VGND 0.03013f
C4891 XThR.Tn[13].n32 VGND 0.09669f
C4892 XThR.Tn[13].t60 VGND 0.01542f
C4893 XThR.Tn[13].t30 VGND 0.01688f
C4894 XThR.Tn[13].n33 VGND 0.04122f
C4895 XThR.Tn[13].t13 VGND 0.01536f
C4896 XThR.Tn[13].t26 VGND 0.01683f
C4897 XThR.Tn[13].n34 VGND 0.04289f
C4898 XThR.Tn[13].n35 VGND 0.03013f
C4899 XThR.Tn[13].n37 VGND 0.09669f
C4900 XThR.Tn[13].t29 VGND 0.01542f
C4901 XThR.Tn[13].t25 VGND 0.01688f
C4902 XThR.Tn[13].n38 VGND 0.04122f
C4903 XThR.Tn[13].t43 VGND 0.01536f
C4904 XThR.Tn[13].t18 VGND 0.01683f
C4905 XThR.Tn[13].n39 VGND 0.04289f
C4906 XThR.Tn[13].n40 VGND 0.03013f
C4907 XThR.Tn[13].n42 VGND 0.09669f
C4908 XThR.Tn[13].t32 VGND 0.01542f
C4909 XThR.Tn[13].t38 VGND 0.01688f
C4910 XThR.Tn[13].n43 VGND 0.04122f
C4911 XThR.Tn[13].t48 VGND 0.01536f
C4912 XThR.Tn[13].t33 VGND 0.01683f
C4913 XThR.Tn[13].n44 VGND 0.04289f
C4914 XThR.Tn[13].n45 VGND 0.03013f
C4915 XThR.Tn[13].n47 VGND 0.09669f
C4916 XThR.Tn[13].t51 VGND 0.01542f
C4917 XThR.Tn[13].t59 VGND 0.01688f
C4918 XThR.Tn[13].n48 VGND 0.04122f
C4919 XThR.Tn[13].t68 VGND 0.01536f
C4920 XThR.Tn[13].t53 VGND 0.01683f
C4921 XThR.Tn[13].n49 VGND 0.04289f
C4922 XThR.Tn[13].n50 VGND 0.03013f
C4923 XThR.Tn[13].n52 VGND 0.09669f
C4924 XThR.Tn[13].t41 VGND 0.01542f
C4925 XThR.Tn[13].t17 VGND 0.01688f
C4926 XThR.Tn[13].n53 VGND 0.04122f
C4927 XThR.Tn[13].t58 VGND 0.01536f
C4928 XThR.Tn[13].t73 VGND 0.01683f
C4929 XThR.Tn[13].n54 VGND 0.04289f
C4930 XThR.Tn[13].n55 VGND 0.03013f
C4931 XThR.Tn[13].n57 VGND 0.09669f
C4932 XThR.Tn[13].t63 VGND 0.01542f
C4933 XThR.Tn[13].t55 VGND 0.01688f
C4934 XThR.Tn[13].n58 VGND 0.04122f
C4935 XThR.Tn[13].t15 VGND 0.01536f
C4936 XThR.Tn[13].t45 VGND 0.01683f
C4937 XThR.Tn[13].n59 VGND 0.04289f
C4938 XThR.Tn[13].n60 VGND 0.03013f
C4939 XThR.Tn[13].n62 VGND 0.09669f
C4940 XThR.Tn[13].t31 VGND 0.01542f
C4941 XThR.Tn[13].t27 VGND 0.01688f
C4942 XThR.Tn[13].n63 VGND 0.04122f
C4943 XThR.Tn[13].t46 VGND 0.01536f
C4944 XThR.Tn[13].t20 VGND 0.01683f
C4945 XThR.Tn[13].n64 VGND 0.04289f
C4946 XThR.Tn[13].n65 VGND 0.03013f
C4947 XThR.Tn[13].n67 VGND 0.09669f
C4948 XThR.Tn[13].t50 VGND 0.01542f
C4949 XThR.Tn[13].t40 VGND 0.01688f
C4950 XThR.Tn[13].n68 VGND 0.04122f
C4951 XThR.Tn[13].t67 VGND 0.01536f
C4952 XThR.Tn[13].t36 VGND 0.01683f
C4953 XThR.Tn[13].n69 VGND 0.04289f
C4954 XThR.Tn[13].n70 VGND 0.03013f
C4955 XThR.Tn[13].n72 VGND 0.09669f
C4956 XThR.Tn[13].t69 VGND 0.01542f
C4957 XThR.Tn[13].t62 VGND 0.01688f
C4958 XThR.Tn[13].n73 VGND 0.04122f
C4959 XThR.Tn[13].t23 VGND 0.01536f
C4960 XThR.Tn[13].t54 VGND 0.01683f
C4961 XThR.Tn[13].n74 VGND 0.04289f
C4962 XThR.Tn[13].n75 VGND 0.03013f
C4963 XThR.Tn[13].n77 VGND 0.09669f
C4964 XThR.Tn[13].t42 VGND 0.01542f
C4965 XThR.Tn[13].t56 VGND 0.01688f
C4966 XThR.Tn[13].n78 VGND 0.04122f
C4967 XThR.Tn[13].t61 VGND 0.01536f
C4968 XThR.Tn[13].t47 VGND 0.01683f
C4969 XThR.Tn[13].n79 VGND 0.04289f
C4970 XThR.Tn[13].n80 VGND 0.03013f
C4971 XThR.Tn[13].n82 VGND 0.09669f
C4972 XThR.Tn[13].n83 VGND 0.08787f
C4973 XThR.Tn[13].n84 VGND 0.34449f
C4974 XThR.Tn[13].t2 VGND 0.01972f
C4975 XThR.Tn[13].t0 VGND 0.01972f
C4976 XThR.Tn[13].n85 VGND 0.04262f
C4977 XThR.Tn[13].t3 VGND 0.01972f
C4978 XThR.Tn[13].t1 VGND 0.01972f
C4979 XThR.Tn[13].n86 VGND 0.06486f
C4980 XThR.Tn[13].n87 VGND 0.1801f
C4981 XThR.Tn[13].n88 VGND 0.02411f
C4982 XThC.XTB3.Y.t1 VGND 0.06296f
C4983 XThC.XTB3.Y.n0 VGND 0.04069f
C4984 XThC.XTB3.Y.n1 VGND 0.05192f
C4985 XThC.XTB3.Y.t0 VGND 0.03159f
C4986 XThC.XTB3.Y.t2 VGND 0.03159f
C4987 XThC.XTB3.Y.n2 VGND 0.06782f
C4988 XThC.XTB3.Y.t10 VGND 0.04914f
C4989 XThC.XTB3.Y.t17 VGND 0.02896f
C4990 XThC.XTB3.Y.n3 VGND 0.05852f
C4991 XThC.XTB3.Y.t14 VGND 0.04914f
C4992 XThC.XTB3.Y.t5 VGND 0.02896f
C4993 XThC.XTB3.Y.n4 VGND 0.03012f
C4994 XThC.XTB3.Y.t15 VGND 0.04914f
C4995 XThC.XTB3.Y.t6 VGND 0.02896f
C4996 XThC.XTB3.Y.n5 VGND 0.06469f
C4997 XThC.XTB3.Y.t3 VGND 0.04914f
C4998 XThC.XTB3.Y.t9 VGND 0.02896f
C4999 XThC.XTB3.Y.n6 VGND 0.06006f
C5000 XThC.XTB3.Y.n7 VGND 0.03654f
C5001 XThC.XTB3.Y.n8 VGND 0.06049f
C5002 XThC.XTB3.Y.n9 VGND 0.0234f
C5003 XThC.XTB3.Y.n10 VGND 0.02857f
C5004 XThC.XTB3.Y.n11 VGND 0.06469f
C5005 XThC.XTB3.Y.n12 VGND 0.03243f
C5006 XThC.XTB3.Y.n13 VGND 0.05514f
C5007 XThC.XTB3.Y.t16 VGND 0.04914f
C5008 XThC.XTB3.Y.t7 VGND 0.02896f
C5009 XThC.XTB3.Y.n14 VGND 0.06624f
C5010 XThC.XTB3.Y.t4 VGND 0.04914f
C5011 XThC.XTB3.Y.t13 VGND 0.02896f
C5012 XThC.XTB3.Y.t12 VGND 0.04914f
C5013 XThC.XTB3.Y.t18 VGND 0.02896f
C5014 XThC.XTB3.Y.t11 VGND 0.04914f
C5015 XThC.XTB3.Y.t8 VGND 0.02896f
C5016 XThC.XTB3.Y.n15 VGND 0.08245f
C5017 XThC.XTB3.Y.n16 VGND 0.08709f
C5018 XThC.XTB3.Y.n17 VGND 0.03356f
C5019 XThC.XTB3.Y.n18 VGND 0.07087f
C5020 XThC.XTB3.Y.n19 VGND 0.03243f
C5021 XThC.XTB3.Y.n20 VGND 0.02691f
C5022 XThC.XTB3.Y.n21 VGND 1.39635f
C5023 XThC.XTB3.Y.n22 VGND 0.14933f
C5024 XThR.Tn[8].t7 VGND 0.01984f
C5025 XThR.Tn[8].t5 VGND 0.01984f
C5026 XThR.Tn[8].n0 VGND 0.06024f
C5027 XThR.Tn[8].t8 VGND 0.01984f
C5028 XThR.Tn[8].t6 VGND 0.01984f
C5029 XThR.Tn[8].n1 VGND 0.04411f
C5030 XThR.Tn[8].n2 VGND 0.20055f
C5031 XThR.Tn[8].t1 VGND 0.0129f
C5032 XThR.Tn[8].t3 VGND 0.0129f
C5033 XThR.Tn[8].n3 VGND 0.03217f
C5034 XThR.Tn[8].t2 VGND 0.0129f
C5035 XThR.Tn[8].t4 VGND 0.0129f
C5036 XThR.Tn[8].n4 VGND 0.02579f
C5037 XThR.Tn[8].n5 VGND 0.05948f
C5038 XThR.Tn[8].t39 VGND 0.01551f
C5039 XThR.Tn[8].t33 VGND 0.01698f
C5040 XThR.Tn[8].n6 VGND 0.04146f
C5041 XThR.Tn[8].n7 VGND 0.07965f
C5042 XThR.Tn[8].t59 VGND 0.01551f
C5043 XThR.Tn[8].t49 VGND 0.01698f
C5044 XThR.Tn[8].n8 VGND 0.04146f
C5045 XThR.Tn[8].t13 VGND 0.01546f
C5046 XThR.Tn[8].t45 VGND 0.01693f
C5047 XThR.Tn[8].n9 VGND 0.04314f
C5048 XThR.Tn[8].n10 VGND 0.03031f
C5049 XThR.Tn[8].n12 VGND 0.09726f
C5050 XThR.Tn[8].t34 VGND 0.01551f
C5051 XThR.Tn[8].t26 VGND 0.01698f
C5052 XThR.Tn[8].n13 VGND 0.04146f
C5053 XThR.Tn[8].t53 VGND 0.01546f
C5054 XThR.Tn[8].t22 VGND 0.01693f
C5055 XThR.Tn[8].n14 VGND 0.04314f
C5056 XThR.Tn[8].n15 VGND 0.03031f
C5057 XThR.Tn[8].n17 VGND 0.09726f
C5058 XThR.Tn[8].t50 VGND 0.01551f
C5059 XThR.Tn[8].t43 VGND 0.01698f
C5060 XThR.Tn[8].n18 VGND 0.04146f
C5061 XThR.Tn[8].t65 VGND 0.01546f
C5062 XThR.Tn[8].t40 VGND 0.01693f
C5063 XThR.Tn[8].n19 VGND 0.04314f
C5064 XThR.Tn[8].n20 VGND 0.03031f
C5065 XThR.Tn[8].n22 VGND 0.09726f
C5066 XThR.Tn[8].t12 VGND 0.01551f
C5067 XThR.Tn[8].t70 VGND 0.01698f
C5068 XThR.Tn[8].n23 VGND 0.04146f
C5069 XThR.Tn[8].t36 VGND 0.01546f
C5070 XThR.Tn[8].t66 VGND 0.01693f
C5071 XThR.Tn[8].n24 VGND 0.04314f
C5072 XThR.Tn[8].n25 VGND 0.03031f
C5073 XThR.Tn[8].n27 VGND 0.09726f
C5074 XThR.Tn[8].t52 VGND 0.01551f
C5075 XThR.Tn[8].t44 VGND 0.01698f
C5076 XThR.Tn[8].n28 VGND 0.04146f
C5077 XThR.Tn[8].t68 VGND 0.01546f
C5078 XThR.Tn[8].t41 VGND 0.01693f
C5079 XThR.Tn[8].n29 VGND 0.04314f
C5080 XThR.Tn[8].n30 VGND 0.03031f
C5081 XThR.Tn[8].n32 VGND 0.09726f
C5082 XThR.Tn[8].t28 VGND 0.01551f
C5083 XThR.Tn[8].t61 VGND 0.01698f
C5084 XThR.Tn[8].n33 VGND 0.04146f
C5085 XThR.Tn[8].t47 VGND 0.01546f
C5086 XThR.Tn[8].t58 VGND 0.01693f
C5087 XThR.Tn[8].n34 VGND 0.04314f
C5088 XThR.Tn[8].n35 VGND 0.03031f
C5089 XThR.Tn[8].n37 VGND 0.09726f
C5090 XThR.Tn[8].t60 VGND 0.01551f
C5091 XThR.Tn[8].t56 VGND 0.01698f
C5092 XThR.Tn[8].n38 VGND 0.04146f
C5093 XThR.Tn[8].t14 VGND 0.01546f
C5094 XThR.Tn[8].t51 VGND 0.01693f
C5095 XThR.Tn[8].n39 VGND 0.04314f
C5096 XThR.Tn[8].n40 VGND 0.03031f
C5097 XThR.Tn[8].n42 VGND 0.09726f
C5098 XThR.Tn[8].t63 VGND 0.01551f
C5099 XThR.Tn[8].t69 VGND 0.01698f
C5100 XThR.Tn[8].n43 VGND 0.04146f
C5101 XThR.Tn[8].t20 VGND 0.01546f
C5102 XThR.Tn[8].t64 VGND 0.01693f
C5103 XThR.Tn[8].n44 VGND 0.04314f
C5104 XThR.Tn[8].n45 VGND 0.03031f
C5105 XThR.Tn[8].n47 VGND 0.09726f
C5106 XThR.Tn[8].t17 VGND 0.01551f
C5107 XThR.Tn[8].t27 VGND 0.01698f
C5108 XThR.Tn[8].n48 VGND 0.04146f
C5109 XThR.Tn[8].t38 VGND 0.01546f
C5110 XThR.Tn[8].t24 VGND 0.01693f
C5111 XThR.Tn[8].n49 VGND 0.04314f
C5112 XThR.Tn[8].n50 VGND 0.03031f
C5113 XThR.Tn[8].n52 VGND 0.09726f
C5114 XThR.Tn[8].t72 VGND 0.01551f
C5115 XThR.Tn[8].t46 VGND 0.01698f
C5116 XThR.Tn[8].n53 VGND 0.04146f
C5117 XThR.Tn[8].t31 VGND 0.01546f
C5118 XThR.Tn[8].t42 VGND 0.01693f
C5119 XThR.Tn[8].n54 VGND 0.04314f
C5120 XThR.Tn[8].n55 VGND 0.03031f
C5121 XThR.Tn[8].n57 VGND 0.09726f
C5122 XThR.Tn[8].t30 VGND 0.01551f
C5123 XThR.Tn[8].t21 VGND 0.01698f
C5124 XThR.Tn[8].n58 VGND 0.04146f
C5125 XThR.Tn[8].t48 VGND 0.01546f
C5126 XThR.Tn[8].t16 VGND 0.01693f
C5127 XThR.Tn[8].n59 VGND 0.04314f
C5128 XThR.Tn[8].n60 VGND 0.03031f
C5129 XThR.Tn[8].n62 VGND 0.09726f
C5130 XThR.Tn[8].t62 VGND 0.01551f
C5131 XThR.Tn[8].t57 VGND 0.01698f
C5132 XThR.Tn[8].n63 VGND 0.04146f
C5133 XThR.Tn[8].t18 VGND 0.01546f
C5134 XThR.Tn[8].t54 VGND 0.01693f
C5135 XThR.Tn[8].n64 VGND 0.04314f
C5136 XThR.Tn[8].n65 VGND 0.03031f
C5137 XThR.Tn[8].n67 VGND 0.09726f
C5138 XThR.Tn[8].t15 VGND 0.01551f
C5139 XThR.Tn[8].t71 VGND 0.01698f
C5140 XThR.Tn[8].n68 VGND 0.04146f
C5141 XThR.Tn[8].t37 VGND 0.01546f
C5142 XThR.Tn[8].t67 VGND 0.01693f
C5143 XThR.Tn[8].n69 VGND 0.04314f
C5144 XThR.Tn[8].n70 VGND 0.03031f
C5145 XThR.Tn[8].n72 VGND 0.09726f
C5146 XThR.Tn[8].t35 VGND 0.01551f
C5147 XThR.Tn[8].t29 VGND 0.01698f
C5148 XThR.Tn[8].n73 VGND 0.04146f
C5149 XThR.Tn[8].t55 VGND 0.01546f
C5150 XThR.Tn[8].t25 VGND 0.01693f
C5151 XThR.Tn[8].n74 VGND 0.04314f
C5152 XThR.Tn[8].n75 VGND 0.03031f
C5153 XThR.Tn[8].n77 VGND 0.09726f
C5154 XThR.Tn[8].t73 VGND 0.01551f
C5155 XThR.Tn[8].t23 VGND 0.01698f
C5156 XThR.Tn[8].n78 VGND 0.04146f
C5157 XThR.Tn[8].t32 VGND 0.01546f
C5158 XThR.Tn[8].t19 VGND 0.01693f
C5159 XThR.Tn[8].n79 VGND 0.04314f
C5160 XThR.Tn[8].n80 VGND 0.03031f
C5161 XThR.Tn[8].n82 VGND 0.09726f
C5162 XThR.Tn[8].n83 VGND 0.08839f
C5163 XThR.Tn[8].n84 VGND 0.27084f
C5164 XThR.Tn[8].t9 VGND 0.01984f
C5165 XThR.Tn[8].t11 VGND 0.01984f
C5166 XThR.Tn[8].n85 VGND 0.04287f
C5167 XThR.Tn[8].t0 VGND 0.01984f
C5168 XThR.Tn[8].t10 VGND 0.01984f
C5169 XThR.Tn[8].n86 VGND 0.06525f
C5170 XThR.Tn[8].n87 VGND 0.18117f
C5171 XThR.Tn[0].t4 VGND 0.01813f
C5172 XThR.Tn[0].t5 VGND 0.01813f
C5173 XThR.Tn[0].n0 VGND 0.03659f
C5174 XThR.Tn[0].t3 VGND 0.01813f
C5175 XThR.Tn[0].t2 VGND 0.01813f
C5176 XThR.Tn[0].n1 VGND 0.04281f
C5177 XThR.Tn[0].n2 VGND 0.12841f
C5178 XThR.Tn[0].t7 VGND 0.01178f
C5179 XThR.Tn[0].t8 VGND 0.01178f
C5180 XThR.Tn[0].n3 VGND 0.02683f
C5181 XThR.Tn[0].t6 VGND 0.01178f
C5182 XThR.Tn[0].t9 VGND 0.01178f
C5183 XThR.Tn[0].n4 VGND 0.02683f
C5184 XThR.Tn[0].t11 VGND 0.01178f
C5185 XThR.Tn[0].t10 VGND 0.01178f
C5186 XThR.Tn[0].n5 VGND 0.0447f
C5187 XThR.Tn[0].t1 VGND 0.01178f
C5188 XThR.Tn[0].t0 VGND 0.01178f
C5189 XThR.Tn[0].n6 VGND 0.02683f
C5190 XThR.Tn[0].n7 VGND 0.12777f
C5191 XThR.Tn[0].n8 VGND 0.07899f
C5192 XThR.Tn[0].n9 VGND 0.08914f
C5193 XThR.Tn[0].t48 VGND 0.01417f
C5194 XThR.Tn[0].t40 VGND 0.01551f
C5195 XThR.Tn[0].n10 VGND 0.03788f
C5196 XThR.Tn[0].n11 VGND 0.07277f
C5197 XThR.Tn[0].t67 VGND 0.01417f
C5198 XThR.Tn[0].t58 VGND 0.01551f
C5199 XThR.Tn[0].n12 VGND 0.03788f
C5200 XThR.Tn[0].t24 VGND 0.01412f
C5201 XThR.Tn[0].t50 VGND 0.01546f
C5202 XThR.Tn[0].n13 VGND 0.03941f
C5203 XThR.Tn[0].n14 VGND 0.02769f
C5204 XThR.Tn[0].n16 VGND 0.08885f
C5205 XThR.Tn[0].t41 VGND 0.01417f
C5206 XThR.Tn[0].t33 VGND 0.01551f
C5207 XThR.Tn[0].n17 VGND 0.03788f
C5208 XThR.Tn[0].t61 VGND 0.01412f
C5209 XThR.Tn[0].t26 VGND 0.01546f
C5210 XThR.Tn[0].n18 VGND 0.03941f
C5211 XThR.Tn[0].n19 VGND 0.02769f
C5212 XThR.Tn[0].n21 VGND 0.08885f
C5213 XThR.Tn[0].t59 VGND 0.01417f
C5214 XThR.Tn[0].t51 VGND 0.01551f
C5215 XThR.Tn[0].n22 VGND 0.03788f
C5216 XThR.Tn[0].t12 VGND 0.01412f
C5217 XThR.Tn[0].t44 VGND 0.01546f
C5218 XThR.Tn[0].n23 VGND 0.03941f
C5219 XThR.Tn[0].n24 VGND 0.02769f
C5220 XThR.Tn[0].n26 VGND 0.08885f
C5221 XThR.Tn[0].t21 VGND 0.01417f
C5222 XThR.Tn[0].t15 VGND 0.01551f
C5223 XThR.Tn[0].n27 VGND 0.03788f
C5224 XThR.Tn[0].t43 VGND 0.01412f
C5225 XThR.Tn[0].t72 VGND 0.01546f
C5226 XThR.Tn[0].n28 VGND 0.03941f
C5227 XThR.Tn[0].n29 VGND 0.02769f
C5228 XThR.Tn[0].n31 VGND 0.08885f
C5229 XThR.Tn[0].t60 VGND 0.01417f
C5230 XThR.Tn[0].t52 VGND 0.01551f
C5231 XThR.Tn[0].n32 VGND 0.03788f
C5232 XThR.Tn[0].t13 VGND 0.01412f
C5233 XThR.Tn[0].t46 VGND 0.01546f
C5234 XThR.Tn[0].n33 VGND 0.03941f
C5235 XThR.Tn[0].n34 VGND 0.02769f
C5236 XThR.Tn[0].n36 VGND 0.08885f
C5237 XThR.Tn[0].t35 VGND 0.01417f
C5238 XThR.Tn[0].t68 VGND 0.01551f
C5239 XThR.Tn[0].n37 VGND 0.03788f
C5240 XThR.Tn[0].t54 VGND 0.01412f
C5241 XThR.Tn[0].t64 VGND 0.01546f
C5242 XThR.Tn[0].n38 VGND 0.03941f
C5243 XThR.Tn[0].n39 VGND 0.02769f
C5244 XThR.Tn[0].n41 VGND 0.08885f
C5245 XThR.Tn[0].t66 VGND 0.01417f
C5246 XThR.Tn[0].t63 VGND 0.01551f
C5247 XThR.Tn[0].n42 VGND 0.03788f
C5248 XThR.Tn[0].t23 VGND 0.01412f
C5249 XThR.Tn[0].t55 VGND 0.01546f
C5250 XThR.Tn[0].n43 VGND 0.03941f
C5251 XThR.Tn[0].n44 VGND 0.02769f
C5252 XThR.Tn[0].n46 VGND 0.08885f
C5253 XThR.Tn[0].t70 VGND 0.01417f
C5254 XThR.Tn[0].t14 VGND 0.01551f
C5255 XThR.Tn[0].n47 VGND 0.03788f
C5256 XThR.Tn[0].t28 VGND 0.01412f
C5257 XThR.Tn[0].t71 VGND 0.01546f
C5258 XThR.Tn[0].n48 VGND 0.03941f
C5259 XThR.Tn[0].n49 VGND 0.02769f
C5260 XThR.Tn[0].n51 VGND 0.08885f
C5261 XThR.Tn[0].t25 VGND 0.01417f
C5262 XThR.Tn[0].t34 VGND 0.01551f
C5263 XThR.Tn[0].n52 VGND 0.03788f
C5264 XThR.Tn[0].t47 VGND 0.01412f
C5265 XThR.Tn[0].t29 VGND 0.01546f
C5266 XThR.Tn[0].n53 VGND 0.03941f
C5267 XThR.Tn[0].n54 VGND 0.02769f
C5268 XThR.Tn[0].n56 VGND 0.08885f
C5269 XThR.Tn[0].t17 VGND 0.01417f
C5270 XThR.Tn[0].t53 VGND 0.01551f
C5271 XThR.Tn[0].n57 VGND 0.03788f
C5272 XThR.Tn[0].t38 VGND 0.01412f
C5273 XThR.Tn[0].t49 VGND 0.01546f
C5274 XThR.Tn[0].n58 VGND 0.03941f
C5275 XThR.Tn[0].n59 VGND 0.02769f
C5276 XThR.Tn[0].n61 VGND 0.08885f
C5277 XThR.Tn[0].t37 VGND 0.01417f
C5278 XThR.Tn[0].t31 VGND 0.01551f
C5279 XThR.Tn[0].n62 VGND 0.03788f
C5280 XThR.Tn[0].t56 VGND 0.01412f
C5281 XThR.Tn[0].t19 VGND 0.01546f
C5282 XThR.Tn[0].n63 VGND 0.03941f
C5283 XThR.Tn[0].n64 VGND 0.02769f
C5284 XThR.Tn[0].n66 VGND 0.08885f
C5285 XThR.Tn[0].t69 VGND 0.01417f
C5286 XThR.Tn[0].t65 VGND 0.01551f
C5287 XThR.Tn[0].n67 VGND 0.03788f
C5288 XThR.Tn[0].t27 VGND 0.01412f
C5289 XThR.Tn[0].t57 VGND 0.01546f
C5290 XThR.Tn[0].n68 VGND 0.03941f
C5291 XThR.Tn[0].n69 VGND 0.02769f
C5292 XThR.Tn[0].n71 VGND 0.08885f
C5293 XThR.Tn[0].t22 VGND 0.01417f
C5294 XThR.Tn[0].t16 VGND 0.01551f
C5295 XThR.Tn[0].n72 VGND 0.03788f
C5296 XThR.Tn[0].t45 VGND 0.01412f
C5297 XThR.Tn[0].t73 VGND 0.01546f
C5298 XThR.Tn[0].n73 VGND 0.03941f
C5299 XThR.Tn[0].n74 VGND 0.02769f
C5300 XThR.Tn[0].n76 VGND 0.08885f
C5301 XThR.Tn[0].t42 VGND 0.01417f
C5302 XThR.Tn[0].t36 VGND 0.01551f
C5303 XThR.Tn[0].n77 VGND 0.03788f
C5304 XThR.Tn[0].t62 VGND 0.01412f
C5305 XThR.Tn[0].t30 VGND 0.01546f
C5306 XThR.Tn[0].n78 VGND 0.03941f
C5307 XThR.Tn[0].n79 VGND 0.02769f
C5308 XThR.Tn[0].n81 VGND 0.08885f
C5309 XThR.Tn[0].t18 VGND 0.01417f
C5310 XThR.Tn[0].t32 VGND 0.01551f
C5311 XThR.Tn[0].n82 VGND 0.03788f
C5312 XThR.Tn[0].t39 VGND 0.01412f
C5313 XThR.Tn[0].t20 VGND 0.01546f
C5314 XThR.Tn[0].n83 VGND 0.03941f
C5315 XThR.Tn[0].n84 VGND 0.02769f
C5316 XThR.Tn[0].n86 VGND 0.08885f
C5317 XThR.Tn[0].n87 VGND 0.08075f
C5318 XThR.Tn[0].n88 VGND 0.2312f
C5319 XThR.Tn[7].t7 VGND 0.01208f
C5320 XThR.Tn[7].t4 VGND 0.01208f
C5321 XThR.Tn[7].n0 VGND 0.03728f
C5322 XThR.Tn[7].t6 VGND 0.01208f
C5323 XThR.Tn[7].t5 VGND 0.01208f
C5324 XThR.Tn[7].n1 VGND 0.02668f
C5325 XThR.Tn[7].n2 VGND 0.13681f
C5326 XThR.Tn[7].t2 VGND 0.01858f
C5327 XThR.Tn[7].t3 VGND 0.01858f
C5328 XThR.Tn[7].n3 VGND 0.05658f
C5329 XThR.Tn[7].t1 VGND 0.01858f
C5330 XThR.Tn[7].t0 VGND 0.01858f
C5331 XThR.Tn[7].n4 VGND 0.04117f
C5332 XThR.Tn[7].n5 VGND 0.18115f
C5333 XThR.Tn[7].n6 VGND 0.02257f
C5334 XThR.Tn[7].t53 VGND 0.01452f
C5335 XThR.Tn[7].t45 VGND 0.0159f
C5336 XThR.Tn[7].n7 VGND 0.03883f
C5337 XThR.Tn[7].n8 VGND 0.0746f
C5338 XThR.Tn[7].t8 VGND 0.01452f
C5339 XThR.Tn[7].t60 VGND 0.0159f
C5340 XThR.Tn[7].n9 VGND 0.03883f
C5341 XThR.Tn[7].t26 VGND 0.01448f
C5342 XThR.Tn[7].t38 VGND 0.01585f
C5343 XThR.Tn[7].n10 VGND 0.04041f
C5344 XThR.Tn[7].n11 VGND 0.02839f
C5345 XThR.Tn[7].n13 VGND 0.09109f
C5346 XThR.Tn[7].t47 VGND 0.01452f
C5347 XThR.Tn[7].t37 VGND 0.0159f
C5348 XThR.Tn[7].n14 VGND 0.03883f
C5349 XThR.Tn[7].t66 VGND 0.01448f
C5350 XThR.Tn[7].t15 VGND 0.01585f
C5351 XThR.Tn[7].n15 VGND 0.04041f
C5352 XThR.Tn[7].n16 VGND 0.02839f
C5353 XThR.Tn[7].n18 VGND 0.09109f
C5354 XThR.Tn[7].t62 VGND 0.01452f
C5355 XThR.Tn[7].t55 VGND 0.0159f
C5356 XThR.Tn[7].n19 VGND 0.03883f
C5357 XThR.Tn[7].t18 VGND 0.01448f
C5358 XThR.Tn[7].t32 VGND 0.01585f
C5359 XThR.Tn[7].n20 VGND 0.04041f
C5360 XThR.Tn[7].n21 VGND 0.02839f
C5361 XThR.Tn[7].n23 VGND 0.09109f
C5362 XThR.Tn[7].t25 VGND 0.01452f
C5363 XThR.Tn[7].t21 VGND 0.0159f
C5364 XThR.Tn[7].n24 VGND 0.03883f
C5365 XThR.Tn[7].t50 VGND 0.01448f
C5366 XThR.Tn[7].t63 VGND 0.01585f
C5367 XThR.Tn[7].n25 VGND 0.04041f
C5368 XThR.Tn[7].n26 VGND 0.02839f
C5369 XThR.Tn[7].n28 VGND 0.09109f
C5370 XThR.Tn[7].t65 VGND 0.01452f
C5371 XThR.Tn[7].t56 VGND 0.0159f
C5372 XThR.Tn[7].n29 VGND 0.03883f
C5373 XThR.Tn[7].t19 VGND 0.01448f
C5374 XThR.Tn[7].t34 VGND 0.01585f
C5375 XThR.Tn[7].n30 VGND 0.04041f
C5376 XThR.Tn[7].n31 VGND 0.02839f
C5377 XThR.Tn[7].n33 VGND 0.09109f
C5378 XThR.Tn[7].t40 VGND 0.01452f
C5379 XThR.Tn[7].t11 VGND 0.0159f
C5380 XThR.Tn[7].n34 VGND 0.03883f
C5381 XThR.Tn[7].t58 VGND 0.01448f
C5382 XThR.Tn[7].t54 VGND 0.01585f
C5383 XThR.Tn[7].n35 VGND 0.04041f
C5384 XThR.Tn[7].n36 VGND 0.02839f
C5385 XThR.Tn[7].n38 VGND 0.09109f
C5386 XThR.Tn[7].t9 VGND 0.01452f
C5387 XThR.Tn[7].t68 VGND 0.0159f
C5388 XThR.Tn[7].n39 VGND 0.03883f
C5389 XThR.Tn[7].t27 VGND 0.01448f
C5390 XThR.Tn[7].t46 VGND 0.01585f
C5391 XThR.Tn[7].n40 VGND 0.04041f
C5392 XThR.Tn[7].n41 VGND 0.02839f
C5393 XThR.Tn[7].n43 VGND 0.09109f
C5394 XThR.Tn[7].t14 VGND 0.01452f
C5395 XThR.Tn[7].t20 VGND 0.0159f
C5396 XThR.Tn[7].n44 VGND 0.03883f
C5397 XThR.Tn[7].t31 VGND 0.01448f
C5398 XThR.Tn[7].t61 VGND 0.01585f
C5399 XThR.Tn[7].n45 VGND 0.04041f
C5400 XThR.Tn[7].n46 VGND 0.02839f
C5401 XThR.Tn[7].n48 VGND 0.09109f
C5402 XThR.Tn[7].t29 VGND 0.01452f
C5403 XThR.Tn[7].t39 VGND 0.0159f
C5404 XThR.Tn[7].n49 VGND 0.03883f
C5405 XThR.Tn[7].t52 VGND 0.01448f
C5406 XThR.Tn[7].t16 VGND 0.01585f
C5407 XThR.Tn[7].n50 VGND 0.04041f
C5408 XThR.Tn[7].n51 VGND 0.02839f
C5409 XThR.Tn[7].n53 VGND 0.09109f
C5410 XThR.Tn[7].t23 VGND 0.01452f
C5411 XThR.Tn[7].t57 VGND 0.0159f
C5412 XThR.Tn[7].n54 VGND 0.03883f
C5413 XThR.Tn[7].t43 VGND 0.01448f
C5414 XThR.Tn[7].t36 VGND 0.01585f
C5415 XThR.Tn[7].n55 VGND 0.04041f
C5416 XThR.Tn[7].n56 VGND 0.02839f
C5417 XThR.Tn[7].n58 VGND 0.09109f
C5418 XThR.Tn[7].t42 VGND 0.01452f
C5419 XThR.Tn[7].t33 VGND 0.0159f
C5420 XThR.Tn[7].n59 VGND 0.03883f
C5421 XThR.Tn[7].t59 VGND 0.01448f
C5422 XThR.Tn[7].t10 VGND 0.01585f
C5423 XThR.Tn[7].n60 VGND 0.04041f
C5424 XThR.Tn[7].n61 VGND 0.02839f
C5425 XThR.Tn[7].n63 VGND 0.09109f
C5426 XThR.Tn[7].t12 VGND 0.01452f
C5427 XThR.Tn[7].t69 VGND 0.0159f
C5428 XThR.Tn[7].n64 VGND 0.03883f
C5429 XThR.Tn[7].t30 VGND 0.01448f
C5430 XThR.Tn[7].t48 VGND 0.01585f
C5431 XThR.Tn[7].n65 VGND 0.04041f
C5432 XThR.Tn[7].n66 VGND 0.02839f
C5433 XThR.Tn[7].n68 VGND 0.09109f
C5434 XThR.Tn[7].t28 VGND 0.01452f
C5435 XThR.Tn[7].t22 VGND 0.0159f
C5436 XThR.Tn[7].n69 VGND 0.03883f
C5437 XThR.Tn[7].t51 VGND 0.01448f
C5438 XThR.Tn[7].t64 VGND 0.01585f
C5439 XThR.Tn[7].n70 VGND 0.04041f
C5440 XThR.Tn[7].n71 VGND 0.02839f
C5441 XThR.Tn[7].n73 VGND 0.09109f
C5442 XThR.Tn[7].t49 VGND 0.01452f
C5443 XThR.Tn[7].t41 VGND 0.0159f
C5444 XThR.Tn[7].n74 VGND 0.03883f
C5445 XThR.Tn[7].t67 VGND 0.01448f
C5446 XThR.Tn[7].t17 VGND 0.01585f
C5447 XThR.Tn[7].n75 VGND 0.04041f
C5448 XThR.Tn[7].n76 VGND 0.02839f
C5449 XThR.Tn[7].n78 VGND 0.09109f
C5450 XThR.Tn[7].t24 VGND 0.01452f
C5451 XThR.Tn[7].t35 VGND 0.0159f
C5452 XThR.Tn[7].n79 VGND 0.03883f
C5453 XThR.Tn[7].t44 VGND 0.01448f
C5454 XThR.Tn[7].t13 VGND 0.01585f
C5455 XThR.Tn[7].n80 VGND 0.04041f
C5456 XThR.Tn[7].n81 VGND 0.02839f
C5457 XThR.Tn[7].n83 VGND 0.09109f
C5458 XThR.Tn[7].n84 VGND 0.08278f
C5459 XThR.Tn[7].n85 VGND 0.33606f
C5460 XThR.Tn[11].t11 VGND 0.01276f
C5461 XThR.Tn[11].t2 VGND 0.01276f
C5462 XThR.Tn[11].n0 VGND 0.02551f
C5463 XThR.Tn[11].t10 VGND 0.01276f
C5464 XThR.Tn[11].t0 VGND 0.01276f
C5465 XThR.Tn[11].n1 VGND 0.03182f
C5466 XThR.Tn[11].n2 VGND 0.06418f
C5467 XThR.Tn[11].t4 VGND 0.01963f
C5468 XThR.Tn[11].t6 VGND 0.01963f
C5469 XThR.Tn[11].n3 VGND 0.05959f
C5470 XThR.Tn[11].t5 VGND 0.01963f
C5471 XThR.Tn[11].t7 VGND 0.01963f
C5472 XThR.Tn[11].n4 VGND 0.04363f
C5473 XThR.Tn[11].n5 VGND 0.19837f
C5474 XThR.Tn[11].t3 VGND 0.01963f
C5475 XThR.Tn[11].t9 VGND 0.01963f
C5476 XThR.Tn[11].n6 VGND 0.0424f
C5477 XThR.Tn[11].t1 VGND 0.01963f
C5478 XThR.Tn[11].t8 VGND 0.01963f
C5479 XThR.Tn[11].n7 VGND 0.06454f
C5480 XThR.Tn[11].n8 VGND 0.1792f
C5481 XThR.Tn[11].n9 VGND 0.02399f
C5482 XThR.Tn[11].t56 VGND 0.01534f
C5483 XThR.Tn[11].t48 VGND 0.0168f
C5484 XThR.Tn[11].n10 VGND 0.04101f
C5485 XThR.Tn[11].n11 VGND 0.07879f
C5486 XThR.Tn[11].t12 VGND 0.01534f
C5487 XThR.Tn[11].t67 VGND 0.0168f
C5488 XThR.Tn[11].n12 VGND 0.04101f
C5489 XThR.Tn[11].t27 VGND 0.01529f
C5490 XThR.Tn[11].t58 VGND 0.01674f
C5491 XThR.Tn[11].n13 VGND 0.04267f
C5492 XThR.Tn[11].n14 VGND 0.02998f
C5493 XThR.Tn[11].n16 VGND 0.0962f
C5494 XThR.Tn[11].t49 VGND 0.01534f
C5495 XThR.Tn[11].t41 VGND 0.0168f
C5496 XThR.Tn[11].n17 VGND 0.04101f
C5497 XThR.Tn[11].t65 VGND 0.01529f
C5498 XThR.Tn[11].t36 VGND 0.01674f
C5499 XThR.Tn[11].n18 VGND 0.04267f
C5500 XThR.Tn[11].n19 VGND 0.02998f
C5501 XThR.Tn[11].n21 VGND 0.0962f
C5502 XThR.Tn[11].t68 VGND 0.01534f
C5503 XThR.Tn[11].t60 VGND 0.0168f
C5504 XThR.Tn[11].n22 VGND 0.04101f
C5505 XThR.Tn[11].t18 VGND 0.01529f
C5506 XThR.Tn[11].t54 VGND 0.01674f
C5507 XThR.Tn[11].n23 VGND 0.04267f
C5508 XThR.Tn[11].n24 VGND 0.02998f
C5509 XThR.Tn[11].n26 VGND 0.0962f
C5510 XThR.Tn[11].t33 VGND 0.01534f
C5511 XThR.Tn[11].t23 VGND 0.0168f
C5512 XThR.Tn[11].n27 VGND 0.04101f
C5513 XThR.Tn[11].t50 VGND 0.01529f
C5514 XThR.Tn[11].t19 VGND 0.01674f
C5515 XThR.Tn[11].n28 VGND 0.04267f
C5516 XThR.Tn[11].n29 VGND 0.02998f
C5517 XThR.Tn[11].n31 VGND 0.0962f
C5518 XThR.Tn[11].t70 VGND 0.01534f
C5519 XThR.Tn[11].t62 VGND 0.0168f
C5520 XThR.Tn[11].n32 VGND 0.04101f
C5521 XThR.Tn[11].t21 VGND 0.01529f
C5522 XThR.Tn[11].t55 VGND 0.01674f
C5523 XThR.Tn[11].n33 VGND 0.04267f
C5524 XThR.Tn[11].n34 VGND 0.02998f
C5525 XThR.Tn[11].n36 VGND 0.0962f
C5526 XThR.Tn[11].t44 VGND 0.01534f
C5527 XThR.Tn[11].t14 VGND 0.0168f
C5528 XThR.Tn[11].n37 VGND 0.04101f
C5529 XThR.Tn[11].t59 VGND 0.01529f
C5530 XThR.Tn[11].t72 VGND 0.01674f
C5531 XThR.Tn[11].n38 VGND 0.04267f
C5532 XThR.Tn[11].n39 VGND 0.02998f
C5533 XThR.Tn[11].n41 VGND 0.0962f
C5534 XThR.Tn[11].t13 VGND 0.01534f
C5535 XThR.Tn[11].t71 VGND 0.0168f
C5536 XThR.Tn[11].n42 VGND 0.04101f
C5537 XThR.Tn[11].t28 VGND 0.01529f
C5538 XThR.Tn[11].t64 VGND 0.01674f
C5539 XThR.Tn[11].n43 VGND 0.04267f
C5540 XThR.Tn[11].n44 VGND 0.02998f
C5541 XThR.Tn[11].n46 VGND 0.0962f
C5542 XThR.Tn[11].t16 VGND 0.01534f
C5543 XThR.Tn[11].t22 VGND 0.0168f
C5544 XThR.Tn[11].n47 VGND 0.04101f
C5545 XThR.Tn[11].t32 VGND 0.01529f
C5546 XThR.Tn[11].t17 VGND 0.01674f
C5547 XThR.Tn[11].n48 VGND 0.04267f
C5548 XThR.Tn[11].n49 VGND 0.02998f
C5549 XThR.Tn[11].n51 VGND 0.0962f
C5550 XThR.Tn[11].t35 VGND 0.01534f
C5551 XThR.Tn[11].t43 VGND 0.0168f
C5552 XThR.Tn[11].n52 VGND 0.04101f
C5553 XThR.Tn[11].t52 VGND 0.01529f
C5554 XThR.Tn[11].t37 VGND 0.01674f
C5555 XThR.Tn[11].n53 VGND 0.04267f
C5556 XThR.Tn[11].n54 VGND 0.02998f
C5557 XThR.Tn[11].n56 VGND 0.0962f
C5558 XThR.Tn[11].t25 VGND 0.01534f
C5559 XThR.Tn[11].t63 VGND 0.0168f
C5560 XThR.Tn[11].n57 VGND 0.04101f
C5561 XThR.Tn[11].t42 VGND 0.01529f
C5562 XThR.Tn[11].t57 VGND 0.01674f
C5563 XThR.Tn[11].n58 VGND 0.04267f
C5564 XThR.Tn[11].n59 VGND 0.02998f
C5565 XThR.Tn[11].n61 VGND 0.0962f
C5566 XThR.Tn[11].t47 VGND 0.01534f
C5567 XThR.Tn[11].t39 VGND 0.0168f
C5568 XThR.Tn[11].n62 VGND 0.04101f
C5569 XThR.Tn[11].t61 VGND 0.01529f
C5570 XThR.Tn[11].t29 VGND 0.01674f
C5571 XThR.Tn[11].n63 VGND 0.04267f
C5572 XThR.Tn[11].n64 VGND 0.02998f
C5573 XThR.Tn[11].n66 VGND 0.0962f
C5574 XThR.Tn[11].t15 VGND 0.01534f
C5575 XThR.Tn[11].t73 VGND 0.0168f
C5576 XThR.Tn[11].n67 VGND 0.04101f
C5577 XThR.Tn[11].t30 VGND 0.01529f
C5578 XThR.Tn[11].t66 VGND 0.01674f
C5579 XThR.Tn[11].n68 VGND 0.04267f
C5580 XThR.Tn[11].n69 VGND 0.02998f
C5581 XThR.Tn[11].n71 VGND 0.0962f
C5582 XThR.Tn[11].t34 VGND 0.01534f
C5583 XThR.Tn[11].t24 VGND 0.0168f
C5584 XThR.Tn[11].n72 VGND 0.04101f
C5585 XThR.Tn[11].t51 VGND 0.01529f
C5586 XThR.Tn[11].t20 VGND 0.01674f
C5587 XThR.Tn[11].n73 VGND 0.04267f
C5588 XThR.Tn[11].n74 VGND 0.02998f
C5589 XThR.Tn[11].n76 VGND 0.0962f
C5590 XThR.Tn[11].t53 VGND 0.01534f
C5591 XThR.Tn[11].t46 VGND 0.0168f
C5592 XThR.Tn[11].n77 VGND 0.04101f
C5593 XThR.Tn[11].t69 VGND 0.01529f
C5594 XThR.Tn[11].t38 VGND 0.01674f
C5595 XThR.Tn[11].n78 VGND 0.04267f
C5596 XThR.Tn[11].n79 VGND 0.02998f
C5597 XThR.Tn[11].n81 VGND 0.0962f
C5598 XThR.Tn[11].t26 VGND 0.01534f
C5599 XThR.Tn[11].t40 VGND 0.0168f
C5600 XThR.Tn[11].n82 VGND 0.04101f
C5601 XThR.Tn[11].t45 VGND 0.01529f
C5602 XThR.Tn[11].t31 VGND 0.01674f
C5603 XThR.Tn[11].n83 VGND 0.04267f
C5604 XThR.Tn[11].n84 VGND 0.02998f
C5605 XThR.Tn[11].n86 VGND 0.0962f
C5606 XThR.Tn[11].n87 VGND 0.08743f
C5607 XThR.Tn[11].n88 VGND 0.31334f
C5608 XThR.Tn[4].t5 VGND 0.01874f
C5609 XThR.Tn[4].t6 VGND 0.01874f
C5610 XThR.Tn[4].n0 VGND 0.03782f
C5611 XThR.Tn[4].t4 VGND 0.01874f
C5612 XThR.Tn[4].t7 VGND 0.01874f
C5613 XThR.Tn[4].n1 VGND 0.04425f
C5614 XThR.Tn[4].n2 VGND 0.13273f
C5615 XThR.Tn[4].t11 VGND 0.01218f
C5616 XThR.Tn[4].t8 VGND 0.01218f
C5617 XThR.Tn[4].n3 VGND 0.02773f
C5618 XThR.Tn[4].t10 VGND 0.01218f
C5619 XThR.Tn[4].t9 VGND 0.01218f
C5620 XThR.Tn[4].n4 VGND 0.02773f
C5621 XThR.Tn[4].t0 VGND 0.01218f
C5622 XThR.Tn[4].t1 VGND 0.01218f
C5623 XThR.Tn[4].n5 VGND 0.04621f
C5624 XThR.Tn[4].t3 VGND 0.01218f
C5625 XThR.Tn[4].t2 VGND 0.01218f
C5626 XThR.Tn[4].n6 VGND 0.02773f
C5627 XThR.Tn[4].n7 VGND 0.13207f
C5628 XThR.Tn[4].n8 VGND 0.08165f
C5629 XThR.Tn[4].n9 VGND 0.09214f
C5630 XThR.Tn[4].t44 VGND 0.01464f
C5631 XThR.Tn[4].t38 VGND 0.01603f
C5632 XThR.Tn[4].n10 VGND 0.03916f
C5633 XThR.Tn[4].n11 VGND 0.07522f
C5634 XThR.Tn[4].t65 VGND 0.01464f
C5635 XThR.Tn[4].t54 VGND 0.01603f
C5636 XThR.Tn[4].n12 VGND 0.03916f
C5637 XThR.Tn[4].t19 VGND 0.0146f
C5638 XThR.Tn[4].t50 VGND 0.01598f
C5639 XThR.Tn[4].n13 VGND 0.04074f
C5640 XThR.Tn[4].n14 VGND 0.02862f
C5641 XThR.Tn[4].n16 VGND 0.09185f
C5642 XThR.Tn[4].t39 VGND 0.01464f
C5643 XThR.Tn[4].t31 VGND 0.01603f
C5644 XThR.Tn[4].n17 VGND 0.03916f
C5645 XThR.Tn[4].t58 VGND 0.0146f
C5646 XThR.Tn[4].t27 VGND 0.01598f
C5647 XThR.Tn[4].n18 VGND 0.04074f
C5648 XThR.Tn[4].n19 VGND 0.02862f
C5649 XThR.Tn[4].n21 VGND 0.09185f
C5650 XThR.Tn[4].t55 VGND 0.01464f
C5651 XThR.Tn[4].t48 VGND 0.01603f
C5652 XThR.Tn[4].n22 VGND 0.03916f
C5653 XThR.Tn[4].t70 VGND 0.0146f
C5654 XThR.Tn[4].t45 VGND 0.01598f
C5655 XThR.Tn[4].n23 VGND 0.04074f
C5656 XThR.Tn[4].n24 VGND 0.02862f
C5657 XThR.Tn[4].n26 VGND 0.09185f
C5658 XThR.Tn[4].t17 VGND 0.01464f
C5659 XThR.Tn[4].t13 VGND 0.01603f
C5660 XThR.Tn[4].n27 VGND 0.03916f
C5661 XThR.Tn[4].t41 VGND 0.0146f
C5662 XThR.Tn[4].t71 VGND 0.01598f
C5663 XThR.Tn[4].n28 VGND 0.04074f
C5664 XThR.Tn[4].n29 VGND 0.02862f
C5665 XThR.Tn[4].n31 VGND 0.09185f
C5666 XThR.Tn[4].t57 VGND 0.01464f
C5667 XThR.Tn[4].t49 VGND 0.01603f
C5668 XThR.Tn[4].n32 VGND 0.03916f
C5669 XThR.Tn[4].t73 VGND 0.0146f
C5670 XThR.Tn[4].t46 VGND 0.01598f
C5671 XThR.Tn[4].n33 VGND 0.04074f
C5672 XThR.Tn[4].n34 VGND 0.02862f
C5673 XThR.Tn[4].n36 VGND 0.09185f
C5674 XThR.Tn[4].t33 VGND 0.01464f
C5675 XThR.Tn[4].t66 VGND 0.01603f
C5676 XThR.Tn[4].n37 VGND 0.03916f
C5677 XThR.Tn[4].t52 VGND 0.0146f
C5678 XThR.Tn[4].t63 VGND 0.01598f
C5679 XThR.Tn[4].n38 VGND 0.04074f
C5680 XThR.Tn[4].n39 VGND 0.02862f
C5681 XThR.Tn[4].n41 VGND 0.09185f
C5682 XThR.Tn[4].t64 VGND 0.01464f
C5683 XThR.Tn[4].t61 VGND 0.01603f
C5684 XThR.Tn[4].n42 VGND 0.03916f
C5685 XThR.Tn[4].t18 VGND 0.0146f
C5686 XThR.Tn[4].t56 VGND 0.01598f
C5687 XThR.Tn[4].n43 VGND 0.04074f
C5688 XThR.Tn[4].n44 VGND 0.02862f
C5689 XThR.Tn[4].n46 VGND 0.09185f
C5690 XThR.Tn[4].t68 VGND 0.01464f
C5691 XThR.Tn[4].t12 VGND 0.01603f
C5692 XThR.Tn[4].n47 VGND 0.03916f
C5693 XThR.Tn[4].t25 VGND 0.0146f
C5694 XThR.Tn[4].t69 VGND 0.01598f
C5695 XThR.Tn[4].n48 VGND 0.04074f
C5696 XThR.Tn[4].n49 VGND 0.02862f
C5697 XThR.Tn[4].n51 VGND 0.09185f
C5698 XThR.Tn[4].t22 VGND 0.01464f
C5699 XThR.Tn[4].t32 VGND 0.01603f
C5700 XThR.Tn[4].n52 VGND 0.03916f
C5701 XThR.Tn[4].t43 VGND 0.0146f
C5702 XThR.Tn[4].t29 VGND 0.01598f
C5703 XThR.Tn[4].n53 VGND 0.04074f
C5704 XThR.Tn[4].n54 VGND 0.02862f
C5705 XThR.Tn[4].n56 VGND 0.09185f
C5706 XThR.Tn[4].t15 VGND 0.01464f
C5707 XThR.Tn[4].t51 VGND 0.01603f
C5708 XThR.Tn[4].n57 VGND 0.03916f
C5709 XThR.Tn[4].t36 VGND 0.0146f
C5710 XThR.Tn[4].t47 VGND 0.01598f
C5711 XThR.Tn[4].n58 VGND 0.04074f
C5712 XThR.Tn[4].n59 VGND 0.02862f
C5713 XThR.Tn[4].n61 VGND 0.09185f
C5714 XThR.Tn[4].t35 VGND 0.01464f
C5715 XThR.Tn[4].t26 VGND 0.01603f
C5716 XThR.Tn[4].n62 VGND 0.03916f
C5717 XThR.Tn[4].t53 VGND 0.0146f
C5718 XThR.Tn[4].t21 VGND 0.01598f
C5719 XThR.Tn[4].n63 VGND 0.04074f
C5720 XThR.Tn[4].n64 VGND 0.02862f
C5721 XThR.Tn[4].n66 VGND 0.09185f
C5722 XThR.Tn[4].t67 VGND 0.01464f
C5723 XThR.Tn[4].t62 VGND 0.01603f
C5724 XThR.Tn[4].n67 VGND 0.03916f
C5725 XThR.Tn[4].t23 VGND 0.0146f
C5726 XThR.Tn[4].t59 VGND 0.01598f
C5727 XThR.Tn[4].n68 VGND 0.04074f
C5728 XThR.Tn[4].n69 VGND 0.02862f
C5729 XThR.Tn[4].n71 VGND 0.09185f
C5730 XThR.Tn[4].t20 VGND 0.01464f
C5731 XThR.Tn[4].t14 VGND 0.01603f
C5732 XThR.Tn[4].n72 VGND 0.03916f
C5733 XThR.Tn[4].t42 VGND 0.0146f
C5734 XThR.Tn[4].t72 VGND 0.01598f
C5735 XThR.Tn[4].n73 VGND 0.04074f
C5736 XThR.Tn[4].n74 VGND 0.02862f
C5737 XThR.Tn[4].n76 VGND 0.09185f
C5738 XThR.Tn[4].t40 VGND 0.01464f
C5739 XThR.Tn[4].t34 VGND 0.01603f
C5740 XThR.Tn[4].n77 VGND 0.03916f
C5741 XThR.Tn[4].t60 VGND 0.0146f
C5742 XThR.Tn[4].t30 VGND 0.01598f
C5743 XThR.Tn[4].n78 VGND 0.04074f
C5744 XThR.Tn[4].n79 VGND 0.02862f
C5745 XThR.Tn[4].n81 VGND 0.09185f
C5746 XThR.Tn[4].t16 VGND 0.01464f
C5747 XThR.Tn[4].t28 VGND 0.01603f
C5748 XThR.Tn[4].n82 VGND 0.03916f
C5749 XThR.Tn[4].t37 VGND 0.0146f
C5750 XThR.Tn[4].t24 VGND 0.01598f
C5751 XThR.Tn[4].n83 VGND 0.04074f
C5752 XThR.Tn[4].n84 VGND 0.02862f
C5753 XThR.Tn[4].n86 VGND 0.09185f
C5754 XThR.Tn[4].n87 VGND 0.08347f
C5755 XThR.Tn[4].n88 VGND 0.15769f
C5756 XThC.Tn[7].n0 VGND 0.02998f
C5757 XThC.Tn[7].n1 VGND 0.02145f
C5758 XThC.Tn[7].n2 VGND 0.1061f
C5759 XThC.Tn[7].t0 VGND 0.01494f
C5760 XThC.Tn[7].t3 VGND 0.01494f
C5761 XThC.Tn[7].n3 VGND 0.03218f
C5762 XThC.Tn[7].t2 VGND 0.01494f
C5763 XThC.Tn[7].t1 VGND 0.01494f
C5764 XThC.Tn[7].n4 VGND 0.04886f
C5765 XThC.Tn[7].n5 VGND 0.14364f
C5766 XThC.Tn[7].t8 VGND 0.01184f
C5767 XThC.Tn[7].t11 VGND 0.01294f
C5768 XThC.Tn[7].n6 VGND 0.02888f
C5769 XThC.Tn[7].n7 VGND 0.01978f
C5770 XThC.Tn[7].n8 VGND 0.06494f
C5771 XThC.Tn[7].t25 VGND 0.01184f
C5772 XThC.Tn[7].t30 VGND 0.01294f
C5773 XThC.Tn[7].n9 VGND 0.02888f
C5774 XThC.Tn[7].n10 VGND 0.01978f
C5775 XThC.Tn[7].n11 VGND 0.06512f
C5776 XThC.Tn[7].n12 VGND 0.10732f
C5777 XThC.Tn[7].t27 VGND 0.01184f
C5778 XThC.Tn[7].t34 VGND 0.01294f
C5779 XThC.Tn[7].n13 VGND 0.02888f
C5780 XThC.Tn[7].n14 VGND 0.01978f
C5781 XThC.Tn[7].n15 VGND 0.06512f
C5782 XThC.Tn[7].n16 VGND 0.10732f
C5783 XThC.Tn[7].t29 VGND 0.01184f
C5784 XThC.Tn[7].t35 VGND 0.01294f
C5785 XThC.Tn[7].n17 VGND 0.02888f
C5786 XThC.Tn[7].n18 VGND 0.01978f
C5787 XThC.Tn[7].n19 VGND 0.06512f
C5788 XThC.Tn[7].n20 VGND 0.10732f
C5789 XThC.Tn[7].t18 VGND 0.01184f
C5790 XThC.Tn[7].t22 VGND 0.01294f
C5791 XThC.Tn[7].n21 VGND 0.02888f
C5792 XThC.Tn[7].n22 VGND 0.01978f
C5793 XThC.Tn[7].n23 VGND 0.06512f
C5794 XThC.Tn[7].n24 VGND 0.10732f
C5795 XThC.Tn[7].t20 VGND 0.01184f
C5796 XThC.Tn[7].t23 VGND 0.01294f
C5797 XThC.Tn[7].n25 VGND 0.02888f
C5798 XThC.Tn[7].n26 VGND 0.01978f
C5799 XThC.Tn[7].n27 VGND 0.06512f
C5800 XThC.Tn[7].n28 VGND 0.10732f
C5801 XThC.Tn[7].t33 VGND 0.01184f
C5802 XThC.Tn[7].t39 VGND 0.01294f
C5803 XThC.Tn[7].n29 VGND 0.02888f
C5804 XThC.Tn[7].n30 VGND 0.01978f
C5805 XThC.Tn[7].n31 VGND 0.06512f
C5806 XThC.Tn[7].n32 VGND 0.10732f
C5807 XThC.Tn[7].t10 VGND 0.01184f
C5808 XThC.Tn[7].t14 VGND 0.01294f
C5809 XThC.Tn[7].n33 VGND 0.02888f
C5810 XThC.Tn[7].n34 VGND 0.01978f
C5811 XThC.Tn[7].n35 VGND 0.06512f
C5812 XThC.Tn[7].n36 VGND 0.10732f
C5813 XThC.Tn[7].t12 VGND 0.01184f
C5814 XThC.Tn[7].t16 VGND 0.01294f
C5815 XThC.Tn[7].n37 VGND 0.02888f
C5816 XThC.Tn[7].n38 VGND 0.01978f
C5817 XThC.Tn[7].n39 VGND 0.06512f
C5818 XThC.Tn[7].n40 VGND 0.10732f
C5819 XThC.Tn[7].t31 VGND 0.01184f
C5820 XThC.Tn[7].t36 VGND 0.01294f
C5821 XThC.Tn[7].n41 VGND 0.02888f
C5822 XThC.Tn[7].n42 VGND 0.01978f
C5823 XThC.Tn[7].n43 VGND 0.06512f
C5824 XThC.Tn[7].n44 VGND 0.10732f
C5825 XThC.Tn[7].t32 VGND 0.01184f
C5826 XThC.Tn[7].t38 VGND 0.01294f
C5827 XThC.Tn[7].n45 VGND 0.02888f
C5828 XThC.Tn[7].n46 VGND 0.01978f
C5829 XThC.Tn[7].n47 VGND 0.06512f
C5830 XThC.Tn[7].n48 VGND 0.10732f
C5831 XThC.Tn[7].t13 VGND 0.01184f
C5832 XThC.Tn[7].t17 VGND 0.01294f
C5833 XThC.Tn[7].n49 VGND 0.02888f
C5834 XThC.Tn[7].n50 VGND 0.01978f
C5835 XThC.Tn[7].n51 VGND 0.06512f
C5836 XThC.Tn[7].n52 VGND 0.10732f
C5837 XThC.Tn[7].t21 VGND 0.01184f
C5838 XThC.Tn[7].t26 VGND 0.01294f
C5839 XThC.Tn[7].n53 VGND 0.02888f
C5840 XThC.Tn[7].n54 VGND 0.01978f
C5841 XThC.Tn[7].n55 VGND 0.06512f
C5842 XThC.Tn[7].n56 VGND 0.10732f
C5843 XThC.Tn[7].t24 VGND 0.01184f
C5844 XThC.Tn[7].t28 VGND 0.01294f
C5845 XThC.Tn[7].n57 VGND 0.02888f
C5846 XThC.Tn[7].n58 VGND 0.01978f
C5847 XThC.Tn[7].n59 VGND 0.06512f
C5848 XThC.Tn[7].n60 VGND 0.10732f
C5849 XThC.Tn[7].t37 VGND 0.01184f
C5850 XThC.Tn[7].t9 VGND 0.01294f
C5851 XThC.Tn[7].n61 VGND 0.02888f
C5852 XThC.Tn[7].n62 VGND 0.01978f
C5853 XThC.Tn[7].n63 VGND 0.06512f
C5854 XThC.Tn[7].n64 VGND 0.10732f
C5855 XThC.Tn[7].t15 VGND 0.01184f
C5856 XThC.Tn[7].t19 VGND 0.01294f
C5857 XThC.Tn[7].n65 VGND 0.02888f
C5858 XThC.Tn[7].n66 VGND 0.01978f
C5859 XThC.Tn[7].n67 VGND 0.06512f
C5860 XThC.Tn[7].n68 VGND 0.10732f
C5861 XThC.Tn[7].n69 VGND 0.26952f
C5862 XThC.Tn[7].n70 VGND 0.01788f
C5863 XThR.Tn[1].t4 VGND 0.01839f
C5864 XThR.Tn[1].t5 VGND 0.01839f
C5865 XThR.Tn[1].n0 VGND 0.03711f
C5866 XThR.Tn[1].t7 VGND 0.01839f
C5867 XThR.Tn[1].t6 VGND 0.01839f
C5868 XThR.Tn[1].n1 VGND 0.04342f
C5869 XThR.Tn[1].n2 VGND 0.12156f
C5870 XThR.Tn[1].t11 VGND 0.01195f
C5871 XThR.Tn[1].t8 VGND 0.01195f
C5872 XThR.Tn[1].n3 VGND 0.02721f
C5873 XThR.Tn[1].t10 VGND 0.01195f
C5874 XThR.Tn[1].t9 VGND 0.01195f
C5875 XThR.Tn[1].n4 VGND 0.02721f
C5876 XThR.Tn[1].t2 VGND 0.01195f
C5877 XThR.Tn[1].t1 VGND 0.01195f
C5878 XThR.Tn[1].n5 VGND 0.02721f
C5879 XThR.Tn[1].t3 VGND 0.01195f
C5880 XThR.Tn[1].t0 VGND 0.01195f
C5881 XThR.Tn[1].n6 VGND 0.04535f
C5882 XThR.Tn[1].n7 VGND 0.1296f
C5883 XThR.Tn[1].n8 VGND 0.08012f
C5884 XThR.Tn[1].n9 VGND 0.09042f
C5885 XThR.Tn[1].t24 VGND 0.01437f
C5886 XThR.Tn[1].t18 VGND 0.01573f
C5887 XThR.Tn[1].n10 VGND 0.03842f
C5888 XThR.Tn[1].n11 VGND 0.07381f
C5889 XThR.Tn[1].t44 VGND 0.01437f
C5890 XThR.Tn[1].t34 VGND 0.01573f
C5891 XThR.Tn[1].n12 VGND 0.03842f
C5892 XThR.Tn[1].t61 VGND 0.01432f
C5893 XThR.Tn[1].t30 VGND 0.01568f
C5894 XThR.Tn[1].n13 VGND 0.03998f
C5895 XThR.Tn[1].n14 VGND 0.02809f
C5896 XThR.Tn[1].n16 VGND 0.09013f
C5897 XThR.Tn[1].t19 VGND 0.01437f
C5898 XThR.Tn[1].t73 VGND 0.01573f
C5899 XThR.Tn[1].n17 VGND 0.03842f
C5900 XThR.Tn[1].t38 VGND 0.01432f
C5901 XThR.Tn[1].t69 VGND 0.01568f
C5902 XThR.Tn[1].n18 VGND 0.03998f
C5903 XThR.Tn[1].n19 VGND 0.02809f
C5904 XThR.Tn[1].n21 VGND 0.09013f
C5905 XThR.Tn[1].t35 VGND 0.01437f
C5906 XThR.Tn[1].t28 VGND 0.01573f
C5907 XThR.Tn[1].n22 VGND 0.03842f
C5908 XThR.Tn[1].t50 VGND 0.01432f
C5909 XThR.Tn[1].t25 VGND 0.01568f
C5910 XThR.Tn[1].n23 VGND 0.03998f
C5911 XThR.Tn[1].n24 VGND 0.02809f
C5912 XThR.Tn[1].n26 VGND 0.09013f
C5913 XThR.Tn[1].t59 VGND 0.01437f
C5914 XThR.Tn[1].t55 VGND 0.01573f
C5915 XThR.Tn[1].n27 VGND 0.03842f
C5916 XThR.Tn[1].t21 VGND 0.01432f
C5917 XThR.Tn[1].t51 VGND 0.01568f
C5918 XThR.Tn[1].n28 VGND 0.03998f
C5919 XThR.Tn[1].n29 VGND 0.02809f
C5920 XThR.Tn[1].n31 VGND 0.09013f
C5921 XThR.Tn[1].t37 VGND 0.01437f
C5922 XThR.Tn[1].t29 VGND 0.01573f
C5923 XThR.Tn[1].n32 VGND 0.03842f
C5924 XThR.Tn[1].t53 VGND 0.01432f
C5925 XThR.Tn[1].t26 VGND 0.01568f
C5926 XThR.Tn[1].n33 VGND 0.03998f
C5927 XThR.Tn[1].n34 VGND 0.02809f
C5928 XThR.Tn[1].n36 VGND 0.09013f
C5929 XThR.Tn[1].t13 VGND 0.01437f
C5930 XThR.Tn[1].t46 VGND 0.01573f
C5931 XThR.Tn[1].n37 VGND 0.03842f
C5932 XThR.Tn[1].t32 VGND 0.01432f
C5933 XThR.Tn[1].t43 VGND 0.01568f
C5934 XThR.Tn[1].n38 VGND 0.03998f
C5935 XThR.Tn[1].n39 VGND 0.02809f
C5936 XThR.Tn[1].n41 VGND 0.09013f
C5937 XThR.Tn[1].t45 VGND 0.01437f
C5938 XThR.Tn[1].t41 VGND 0.01573f
C5939 XThR.Tn[1].n42 VGND 0.03842f
C5940 XThR.Tn[1].t60 VGND 0.01432f
C5941 XThR.Tn[1].t36 VGND 0.01568f
C5942 XThR.Tn[1].n43 VGND 0.03998f
C5943 XThR.Tn[1].n44 VGND 0.02809f
C5944 XThR.Tn[1].n46 VGND 0.09013f
C5945 XThR.Tn[1].t48 VGND 0.01437f
C5946 XThR.Tn[1].t54 VGND 0.01573f
C5947 XThR.Tn[1].n47 VGND 0.03842f
C5948 XThR.Tn[1].t67 VGND 0.01432f
C5949 XThR.Tn[1].t49 VGND 0.01568f
C5950 XThR.Tn[1].n48 VGND 0.03998f
C5951 XThR.Tn[1].n49 VGND 0.02809f
C5952 XThR.Tn[1].n51 VGND 0.09013f
C5953 XThR.Tn[1].t64 VGND 0.01437f
C5954 XThR.Tn[1].t12 VGND 0.01573f
C5955 XThR.Tn[1].n52 VGND 0.03842f
C5956 XThR.Tn[1].t23 VGND 0.01432f
C5957 XThR.Tn[1].t71 VGND 0.01568f
C5958 XThR.Tn[1].n53 VGND 0.03998f
C5959 XThR.Tn[1].n54 VGND 0.02809f
C5960 XThR.Tn[1].n56 VGND 0.09013f
C5961 XThR.Tn[1].t57 VGND 0.01437f
C5962 XThR.Tn[1].t31 VGND 0.01573f
C5963 XThR.Tn[1].n57 VGND 0.03842f
C5964 XThR.Tn[1].t16 VGND 0.01432f
C5965 XThR.Tn[1].t27 VGND 0.01568f
C5966 XThR.Tn[1].n58 VGND 0.03998f
C5967 XThR.Tn[1].n59 VGND 0.02809f
C5968 XThR.Tn[1].n61 VGND 0.09013f
C5969 XThR.Tn[1].t15 VGND 0.01437f
C5970 XThR.Tn[1].t68 VGND 0.01573f
C5971 XThR.Tn[1].n62 VGND 0.03842f
C5972 XThR.Tn[1].t33 VGND 0.01432f
C5973 XThR.Tn[1].t63 VGND 0.01568f
C5974 XThR.Tn[1].n63 VGND 0.03998f
C5975 XThR.Tn[1].n64 VGND 0.02809f
C5976 XThR.Tn[1].n66 VGND 0.09013f
C5977 XThR.Tn[1].t47 VGND 0.01437f
C5978 XThR.Tn[1].t42 VGND 0.01573f
C5979 XThR.Tn[1].n67 VGND 0.03842f
C5980 XThR.Tn[1].t65 VGND 0.01432f
C5981 XThR.Tn[1].t39 VGND 0.01568f
C5982 XThR.Tn[1].n68 VGND 0.03998f
C5983 XThR.Tn[1].n69 VGND 0.02809f
C5984 XThR.Tn[1].n71 VGND 0.09013f
C5985 XThR.Tn[1].t62 VGND 0.01437f
C5986 XThR.Tn[1].t56 VGND 0.01573f
C5987 XThR.Tn[1].n72 VGND 0.03842f
C5988 XThR.Tn[1].t22 VGND 0.01432f
C5989 XThR.Tn[1].t52 VGND 0.01568f
C5990 XThR.Tn[1].n73 VGND 0.03998f
C5991 XThR.Tn[1].n74 VGND 0.02809f
C5992 XThR.Tn[1].n76 VGND 0.09013f
C5993 XThR.Tn[1].t20 VGND 0.01437f
C5994 XThR.Tn[1].t14 VGND 0.01573f
C5995 XThR.Tn[1].n77 VGND 0.03842f
C5996 XThR.Tn[1].t40 VGND 0.01432f
C5997 XThR.Tn[1].t72 VGND 0.01568f
C5998 XThR.Tn[1].n78 VGND 0.03998f
C5999 XThR.Tn[1].n79 VGND 0.02809f
C6000 XThR.Tn[1].n81 VGND 0.09013f
C6001 XThR.Tn[1].t58 VGND 0.01437f
C6002 XThR.Tn[1].t70 VGND 0.01573f
C6003 XThR.Tn[1].n82 VGND 0.03842f
C6004 XThR.Tn[1].t17 VGND 0.01432f
C6005 XThR.Tn[1].t66 VGND 0.01568f
C6006 XThR.Tn[1].n83 VGND 0.03998f
C6007 XThR.Tn[1].n84 VGND 0.02809f
C6008 XThR.Tn[1].n86 VGND 0.09013f
C6009 XThR.Tn[1].n87 VGND 0.0819f
C6010 XThR.Tn[1].n88 VGND 0.23576f
C6011 XThR.Tn[1].n89 VGND 0.03847f
C6012 XThC.Tn[8].t9 VGND 0.01061f
C6013 XThC.Tn[8].t8 VGND 0.01061f
C6014 XThC.Tn[8].n0 VGND 0.02645f
C6015 XThC.Tn[8].t11 VGND 0.01061f
C6016 XThC.Tn[8].t10 VGND 0.01061f
C6017 XThC.Tn[8].n1 VGND 0.02121f
C6018 XThC.Tn[8].n2 VGND 0.05336f
C6019 XThC.Tn[8].n3 VGND 0.01995f
C6020 XThC.Tn[8].t43 VGND 0.01293f
C6021 XThC.Tn[8].t41 VGND 0.01413f
C6022 XThC.Tn[8].n4 VGND 0.03153f
C6023 XThC.Tn[8].n5 VGND 0.0216f
C6024 XThC.Tn[8].n6 VGND 0.07091f
C6025 XThC.Tn[8].t29 VGND 0.01293f
C6026 XThC.Tn[8].t26 VGND 0.01413f
C6027 XThC.Tn[8].n7 VGND 0.03153f
C6028 XThC.Tn[8].n8 VGND 0.0216f
C6029 XThC.Tn[8].n9 VGND 0.0711f
C6030 XThC.Tn[8].n10 VGND 0.11718f
C6031 XThC.Tn[8].t34 VGND 0.01293f
C6032 XThC.Tn[8].t28 VGND 0.01413f
C6033 XThC.Tn[8].n11 VGND 0.03153f
C6034 XThC.Tn[8].n12 VGND 0.0216f
C6035 XThC.Tn[8].n13 VGND 0.0711f
C6036 XThC.Tn[8].n14 VGND 0.11718f
C6037 XThC.Tn[8].t35 VGND 0.01293f
C6038 XThC.Tn[8].t30 VGND 0.01413f
C6039 XThC.Tn[8].n15 VGND 0.03153f
C6040 XThC.Tn[8].n16 VGND 0.0216f
C6041 XThC.Tn[8].n17 VGND 0.0711f
C6042 XThC.Tn[8].n18 VGND 0.11718f
C6043 XThC.Tn[8].t22 VGND 0.01293f
C6044 XThC.Tn[8].t19 VGND 0.01413f
C6045 XThC.Tn[8].n19 VGND 0.03153f
C6046 XThC.Tn[8].n20 VGND 0.0216f
C6047 XThC.Tn[8].n21 VGND 0.0711f
C6048 XThC.Tn[8].n22 VGND 0.11718f
C6049 XThC.Tn[8].t23 VGND 0.01293f
C6050 XThC.Tn[8].t20 VGND 0.01413f
C6051 XThC.Tn[8].n23 VGND 0.03153f
C6052 XThC.Tn[8].n24 VGND 0.0216f
C6053 XThC.Tn[8].n25 VGND 0.0711f
C6054 XThC.Tn[8].n26 VGND 0.11718f
C6055 XThC.Tn[8].t39 VGND 0.01293f
C6056 XThC.Tn[8].t33 VGND 0.01413f
C6057 XThC.Tn[8].n27 VGND 0.03153f
C6058 XThC.Tn[8].n28 VGND 0.0216f
C6059 XThC.Tn[8].n29 VGND 0.0711f
C6060 XThC.Tn[8].n30 VGND 0.11718f
C6061 XThC.Tn[8].t14 VGND 0.01293f
C6062 XThC.Tn[8].t42 VGND 0.01413f
C6063 XThC.Tn[8].n31 VGND 0.03153f
C6064 XThC.Tn[8].n32 VGND 0.0216f
C6065 XThC.Tn[8].n33 VGND 0.0711f
C6066 XThC.Tn[8].n34 VGND 0.11718f
C6067 XThC.Tn[8].t16 VGND 0.01293f
C6068 XThC.Tn[8].t12 VGND 0.01413f
C6069 XThC.Tn[8].n35 VGND 0.03153f
C6070 XThC.Tn[8].n36 VGND 0.0216f
C6071 XThC.Tn[8].n37 VGND 0.0711f
C6072 XThC.Tn[8].n38 VGND 0.11718f
C6073 XThC.Tn[8].t36 VGND 0.01293f
C6074 XThC.Tn[8].t31 VGND 0.01413f
C6075 XThC.Tn[8].n39 VGND 0.03153f
C6076 XThC.Tn[8].n40 VGND 0.0216f
C6077 XThC.Tn[8].n41 VGND 0.0711f
C6078 XThC.Tn[8].n42 VGND 0.11718f
C6079 XThC.Tn[8].t38 VGND 0.01293f
C6080 XThC.Tn[8].t32 VGND 0.01413f
C6081 XThC.Tn[8].n43 VGND 0.03153f
C6082 XThC.Tn[8].n44 VGND 0.0216f
C6083 XThC.Tn[8].n45 VGND 0.0711f
C6084 XThC.Tn[8].n46 VGND 0.11718f
C6085 XThC.Tn[8].t17 VGND 0.01293f
C6086 XThC.Tn[8].t13 VGND 0.01413f
C6087 XThC.Tn[8].n47 VGND 0.03153f
C6088 XThC.Tn[8].n48 VGND 0.0216f
C6089 XThC.Tn[8].n49 VGND 0.0711f
C6090 XThC.Tn[8].n50 VGND 0.11718f
C6091 XThC.Tn[8].t25 VGND 0.01293f
C6092 XThC.Tn[8].t21 VGND 0.01413f
C6093 XThC.Tn[8].n51 VGND 0.03153f
C6094 XThC.Tn[8].n52 VGND 0.0216f
C6095 XThC.Tn[8].n53 VGND 0.0711f
C6096 XThC.Tn[8].n54 VGND 0.11718f
C6097 XThC.Tn[8].t27 VGND 0.01293f
C6098 XThC.Tn[8].t24 VGND 0.01413f
C6099 XThC.Tn[8].n55 VGND 0.03153f
C6100 XThC.Tn[8].n56 VGND 0.0216f
C6101 XThC.Tn[8].n57 VGND 0.0711f
C6102 XThC.Tn[8].n58 VGND 0.11718f
C6103 XThC.Tn[8].t40 VGND 0.01293f
C6104 XThC.Tn[8].t37 VGND 0.01413f
C6105 XThC.Tn[8].n59 VGND 0.03153f
C6106 XThC.Tn[8].n60 VGND 0.0216f
C6107 XThC.Tn[8].n61 VGND 0.0711f
C6108 XThC.Tn[8].n62 VGND 0.11718f
C6109 XThC.Tn[8].t18 VGND 0.01293f
C6110 XThC.Tn[8].t15 VGND 0.01413f
C6111 XThC.Tn[8].n63 VGND 0.03153f
C6112 XThC.Tn[8].n64 VGND 0.0216f
C6113 XThC.Tn[8].n65 VGND 0.0711f
C6114 XThC.Tn[8].n66 VGND 0.11718f
C6115 XThC.Tn[8].n67 VGND 0.49072f
C6116 XThC.Tn[8].n68 VGND 0.19206f
C6117 XThC.Tn[8].t5 VGND 0.01632f
C6118 XThC.Tn[8].t6 VGND 0.01632f
C6119 XThC.Tn[8].n69 VGND 0.03525f
C6120 XThC.Tn[8].t4 VGND 0.01632f
C6121 XThC.Tn[8].t7 VGND 0.01632f
C6122 XThC.Tn[8].n70 VGND 0.05365f
C6123 XThC.Tn[8].n71 VGND 0.14908f
C6124 XThC.Tn[8].n72 VGND 0.02344f
C6125 XThC.Tn[8].t2 VGND 0.01632f
C6126 XThC.Tn[8].t1 VGND 0.01632f
C6127 XThC.Tn[8].n73 VGND 0.03627f
C6128 XThC.Tn[8].t0 VGND 0.01632f
C6129 XThC.Tn[8].t3 VGND 0.01632f
C6130 XThC.Tn[8].n74 VGND 0.04954f
C6131 XThC.Tn[8].n75 VGND 0.16142f
C6132 XThC.XTB1.Y.t2 VGND 0.03224f
C6133 XThC.XTB1.Y.n0 VGND 0.02084f
C6134 XThC.XTB1.Y.n1 VGND 0.02659f
C6135 XThC.XTB1.Y.t1 VGND 0.01618f
C6136 XThC.XTB1.Y.t0 VGND 0.01618f
C6137 XThC.XTB1.Y.n2 VGND 0.03473f
C6138 XThC.XTB1.Y.t17 VGND 0.02517f
C6139 XThC.XTB1.Y.t5 VGND 0.01483f
C6140 XThC.XTB1.Y.n3 VGND 0.02997f
C6141 XThC.XTB1.Y.t6 VGND 0.02517f
C6142 XThC.XTB1.Y.t12 VGND 0.01483f
C6143 XThC.XTB1.Y.n4 VGND 0.01542f
C6144 XThC.XTB1.Y.t8 VGND 0.02517f
C6145 XThC.XTB1.Y.t13 VGND 0.01483f
C6146 XThC.XTB1.Y.n5 VGND 0.03313f
C6147 XThC.XTB1.Y.t11 VGND 0.02517f
C6148 XThC.XTB1.Y.t16 VGND 0.01483f
C6149 XThC.XTB1.Y.n6 VGND 0.03076f
C6150 XThC.XTB1.Y.n7 VGND 0.01871f
C6151 XThC.XTB1.Y.n8 VGND 0.03098f
C6152 XThC.XTB1.Y.n9 VGND 0.01198f
C6153 XThC.XTB1.Y.n10 VGND 0.01463f
C6154 XThC.XTB1.Y.n11 VGND 0.03313f
C6155 XThC.XTB1.Y.n12 VGND 0.01661f
C6156 XThC.XTB1.Y.n13 VGND 0.02824f
C6157 XThC.XTB1.Y.t18 VGND 0.02517f
C6158 XThC.XTB1.Y.t9 VGND 0.01483f
C6159 XThC.XTB1.Y.n14 VGND 0.03392f
C6160 XThC.XTB1.Y.t7 VGND 0.02517f
C6161 XThC.XTB1.Y.t15 VGND 0.01483f
C6162 XThC.XTB1.Y.t14 VGND 0.02517f
C6163 XThC.XTB1.Y.t3 VGND 0.01483f
C6164 XThC.XTB1.Y.t10 VGND 0.02517f
C6165 XThC.XTB1.Y.t4 VGND 0.01483f
C6166 XThC.XTB1.Y.n15 VGND 0.04223f
C6167 XThC.XTB1.Y.n16 VGND 0.0446f
C6168 XThC.XTB1.Y.n17 VGND 0.01719f
C6169 XThC.XTB1.Y.n18 VGND 0.0363f
C6170 XThC.XTB1.Y.n19 VGND 0.01661f
C6171 XThC.XTB1.Y.n20 VGND 0.01378f
C6172 XThC.XTB1.Y.n21 VGND 0.77148f
C6173 XThC.XTB1.Y.n22 VGND 0.07634f
C6174 XThC.Tn[14].n0 VGND 0.02478f
C6175 XThC.Tn[14].n1 VGND 0.01987f
C6176 XThC.Tn[14].n2 VGND 0.04998f
C6177 XThC.Tn[14].t43 VGND 0.01211f
C6178 XThC.Tn[14].t38 VGND 0.01323f
C6179 XThC.Tn[14].n3 VGND 0.02954f
C6180 XThC.Tn[14].n4 VGND 0.02024f
C6181 XThC.Tn[14].n5 VGND 0.06643f
C6182 XThC.Tn[14].t29 VGND 0.01211f
C6183 XThC.Tn[14].t22 VGND 0.01323f
C6184 XThC.Tn[14].n6 VGND 0.02954f
C6185 XThC.Tn[14].n7 VGND 0.02024f
C6186 XThC.Tn[14].n8 VGND 0.06661f
C6187 XThC.Tn[14].n9 VGND 0.10978f
C6188 XThC.Tn[14].t32 VGND 0.01211f
C6189 XThC.Tn[14].t25 VGND 0.01323f
C6190 XThC.Tn[14].n10 VGND 0.02954f
C6191 XThC.Tn[14].n11 VGND 0.02024f
C6192 XThC.Tn[14].n12 VGND 0.06661f
C6193 XThC.Tn[14].n13 VGND 0.10978f
C6194 XThC.Tn[14].t34 VGND 0.01211f
C6195 XThC.Tn[14].t26 VGND 0.01323f
C6196 XThC.Tn[14].n14 VGND 0.02954f
C6197 XThC.Tn[14].n15 VGND 0.02024f
C6198 XThC.Tn[14].n16 VGND 0.06661f
C6199 XThC.Tn[14].n17 VGND 0.10978f
C6200 XThC.Tn[14].t20 VGND 0.01211f
C6201 XThC.Tn[14].t14 VGND 0.01323f
C6202 XThC.Tn[14].n18 VGND 0.02954f
C6203 XThC.Tn[14].n19 VGND 0.02024f
C6204 XThC.Tn[14].n20 VGND 0.06661f
C6205 XThC.Tn[14].n21 VGND 0.10978f
C6206 XThC.Tn[14].t23 VGND 0.01211f
C6207 XThC.Tn[14].t17 VGND 0.01323f
C6208 XThC.Tn[14].n22 VGND 0.02954f
C6209 XThC.Tn[14].n23 VGND 0.02024f
C6210 XThC.Tn[14].n24 VGND 0.06661f
C6211 XThC.Tn[14].n25 VGND 0.10978f
C6212 XThC.Tn[14].t37 VGND 0.01211f
C6213 XThC.Tn[14].t31 VGND 0.01323f
C6214 XThC.Tn[14].n26 VGND 0.02954f
C6215 XThC.Tn[14].n27 VGND 0.02024f
C6216 XThC.Tn[14].n28 VGND 0.06661f
C6217 XThC.Tn[14].n29 VGND 0.10978f
C6218 XThC.Tn[14].t13 VGND 0.01211f
C6219 XThC.Tn[14].t39 VGND 0.01323f
C6220 XThC.Tn[14].n30 VGND 0.02954f
C6221 XThC.Tn[14].n31 VGND 0.02024f
C6222 XThC.Tn[14].n32 VGND 0.06661f
C6223 XThC.Tn[14].n33 VGND 0.10978f
C6224 XThC.Tn[14].t15 VGND 0.01211f
C6225 XThC.Tn[14].t41 VGND 0.01323f
C6226 XThC.Tn[14].n34 VGND 0.02954f
C6227 XThC.Tn[14].n35 VGND 0.02024f
C6228 XThC.Tn[14].n36 VGND 0.06661f
C6229 XThC.Tn[14].n37 VGND 0.10978f
C6230 XThC.Tn[14].t35 VGND 0.01211f
C6231 XThC.Tn[14].t27 VGND 0.01323f
C6232 XThC.Tn[14].n38 VGND 0.02954f
C6233 XThC.Tn[14].n39 VGND 0.02024f
C6234 XThC.Tn[14].n40 VGND 0.06661f
C6235 XThC.Tn[14].n41 VGND 0.10978f
C6236 XThC.Tn[14].t36 VGND 0.01211f
C6237 XThC.Tn[14].t30 VGND 0.01323f
C6238 XThC.Tn[14].n42 VGND 0.02954f
C6239 XThC.Tn[14].n43 VGND 0.02024f
C6240 XThC.Tn[14].n44 VGND 0.06661f
C6241 XThC.Tn[14].n45 VGND 0.10978f
C6242 XThC.Tn[14].t16 VGND 0.01211f
C6243 XThC.Tn[14].t42 VGND 0.01323f
C6244 XThC.Tn[14].n46 VGND 0.02954f
C6245 XThC.Tn[14].n47 VGND 0.02024f
C6246 XThC.Tn[14].n48 VGND 0.06661f
C6247 XThC.Tn[14].n49 VGND 0.10978f
C6248 XThC.Tn[14].t24 VGND 0.01211f
C6249 XThC.Tn[14].t19 VGND 0.01323f
C6250 XThC.Tn[14].n50 VGND 0.02954f
C6251 XThC.Tn[14].n51 VGND 0.02024f
C6252 XThC.Tn[14].n52 VGND 0.06661f
C6253 XThC.Tn[14].n53 VGND 0.10978f
C6254 XThC.Tn[14].t28 VGND 0.01211f
C6255 XThC.Tn[14].t21 VGND 0.01323f
C6256 XThC.Tn[14].n54 VGND 0.02954f
C6257 XThC.Tn[14].n55 VGND 0.02024f
C6258 XThC.Tn[14].n56 VGND 0.06661f
C6259 XThC.Tn[14].n57 VGND 0.10978f
C6260 XThC.Tn[14].t40 VGND 0.01211f
C6261 XThC.Tn[14].t33 VGND 0.01323f
C6262 XThC.Tn[14].n58 VGND 0.02954f
C6263 XThC.Tn[14].n59 VGND 0.02024f
C6264 XThC.Tn[14].n60 VGND 0.06661f
C6265 XThC.Tn[14].n61 VGND 0.10978f
C6266 XThC.Tn[14].t18 VGND 0.01211f
C6267 XThC.Tn[14].t12 VGND 0.01323f
C6268 XThC.Tn[14].n62 VGND 0.02954f
C6269 XThC.Tn[14].n63 VGND 0.02024f
C6270 XThC.Tn[14].n64 VGND 0.06661f
C6271 XThC.Tn[14].n65 VGND 0.10978f
C6272 XThC.Tn[14].n66 VGND 0.72002f
C6273 XThC.Tn[14].n67 VGND 0.21181f
C6274 XThC.Tn[14].t4 VGND 0.01528f
C6275 XThC.Tn[14].t5 VGND 0.01528f
C6276 XThC.Tn[14].n68 VGND 0.03302f
C6277 XThC.Tn[14].t7 VGND 0.01528f
C6278 XThC.Tn[14].t6 VGND 0.01528f
C6279 XThC.Tn[14].n69 VGND 0.05026f
C6280 XThC.Tn[14].n70 VGND 0.13966f
C6281 XThC.Tn[14].n71 VGND 0.02196f
C6282 XThC.Tn[14].t1 VGND 0.01528f
C6283 XThC.Tn[14].t0 VGND 0.01528f
C6284 XThC.Tn[14].n72 VGND 0.03398f
C6285 XThC.Tn[14].t3 VGND 0.01528f
C6286 XThC.Tn[14].t2 VGND 0.01528f
C6287 XThC.Tn[14].n73 VGND 0.04641f
C6288 XThC.Tn[14].n74 VGND 0.15122f
C6289 XThR.Tn[10].t10 VGND 0.01984f
C6290 XThR.Tn[10].t8 VGND 0.01984f
C6291 XThR.Tn[10].n0 VGND 0.06023f
C6292 XThR.Tn[10].t11 VGND 0.01984f
C6293 XThR.Tn[10].t9 VGND 0.01984f
C6294 XThR.Tn[10].n1 VGND 0.0441f
C6295 XThR.Tn[10].n2 VGND 0.20051f
C6296 XThR.Tn[10].t7 VGND 0.01289f
C6297 XThR.Tn[10].t6 VGND 0.01289f
C6298 XThR.Tn[10].n3 VGND 0.03216f
C6299 XThR.Tn[10].t2 VGND 0.01289f
C6300 XThR.Tn[10].t3 VGND 0.01289f
C6301 XThR.Tn[10].n4 VGND 0.02579f
C6302 XThR.Tn[10].n5 VGND 0.05947f
C6303 XThR.Tn[10].t54 VGND 0.0155f
C6304 XThR.Tn[10].t47 VGND 0.01698f
C6305 XThR.Tn[10].n6 VGND 0.04146f
C6306 XThR.Tn[10].n7 VGND 0.07964f
C6307 XThR.Tn[10].t13 VGND 0.0155f
C6308 XThR.Tn[10].t63 VGND 0.01698f
C6309 XThR.Tn[10].n8 VGND 0.04146f
C6310 XThR.Tn[10].t50 VGND 0.01545f
C6311 XThR.Tn[10].t60 VGND 0.01692f
C6312 XThR.Tn[10].n9 VGND 0.04313f
C6313 XThR.Tn[10].n10 VGND 0.0303f
C6314 XThR.Tn[10].n12 VGND 0.09724f
C6315 XThR.Tn[10].t48 VGND 0.0155f
C6316 XThR.Tn[10].t41 VGND 0.01698f
C6317 XThR.Tn[10].n13 VGND 0.04146f
C6318 XThR.Tn[10].t23 VGND 0.01545f
C6319 XThR.Tn[10].t36 VGND 0.01692f
C6320 XThR.Tn[10].n14 VGND 0.04313f
C6321 XThR.Tn[10].n15 VGND 0.0303f
C6322 XThR.Tn[10].n17 VGND 0.09724f
C6323 XThR.Tn[10].t65 VGND 0.0155f
C6324 XThR.Tn[10].t58 VGND 0.01698f
C6325 XThR.Tn[10].n18 VGND 0.04146f
C6326 XThR.Tn[10].t40 VGND 0.01545f
C6327 XThR.Tn[10].t55 VGND 0.01692f
C6328 XThR.Tn[10].n19 VGND 0.04313f
C6329 XThR.Tn[10].n20 VGND 0.0303f
C6330 XThR.Tn[10].n22 VGND 0.09724f
C6331 XThR.Tn[10].t30 VGND 0.0155f
C6332 XThR.Tn[10].t26 VGND 0.01698f
C6333 XThR.Tn[10].n23 VGND 0.04146f
C6334 XThR.Tn[10].t70 VGND 0.01545f
C6335 XThR.Tn[10].t21 VGND 0.01692f
C6336 XThR.Tn[10].n24 VGND 0.04313f
C6337 XThR.Tn[10].n25 VGND 0.0303f
C6338 XThR.Tn[10].n27 VGND 0.09724f
C6339 XThR.Tn[10].t67 VGND 0.0155f
C6340 XThR.Tn[10].t59 VGND 0.01698f
C6341 XThR.Tn[10].n28 VGND 0.04146f
C6342 XThR.Tn[10].t42 VGND 0.01545f
C6343 XThR.Tn[10].t56 VGND 0.01692f
C6344 XThR.Tn[10].n29 VGND 0.04313f
C6345 XThR.Tn[10].n30 VGND 0.0303f
C6346 XThR.Tn[10].n32 VGND 0.09724f
C6347 XThR.Tn[10].t44 VGND 0.0155f
C6348 XThR.Tn[10].t15 VGND 0.01698f
C6349 XThR.Tn[10].n33 VGND 0.04146f
C6350 XThR.Tn[10].t18 VGND 0.01545f
C6351 XThR.Tn[10].t12 VGND 0.01692f
C6352 XThR.Tn[10].n34 VGND 0.04313f
C6353 XThR.Tn[10].n35 VGND 0.0303f
C6354 XThR.Tn[10].n37 VGND 0.09724f
C6355 XThR.Tn[10].t14 VGND 0.0155f
C6356 XThR.Tn[10].t69 VGND 0.01698f
C6357 XThR.Tn[10].n38 VGND 0.04146f
C6358 XThR.Tn[10].t51 VGND 0.01545f
C6359 XThR.Tn[10].t66 VGND 0.01692f
C6360 XThR.Tn[10].n39 VGND 0.04313f
C6361 XThR.Tn[10].n40 VGND 0.0303f
C6362 XThR.Tn[10].n42 VGND 0.09724f
C6363 XThR.Tn[10].t17 VGND 0.0155f
C6364 XThR.Tn[10].t24 VGND 0.01698f
C6365 XThR.Tn[10].n43 VGND 0.04146f
C6366 XThR.Tn[10].t53 VGND 0.01545f
C6367 XThR.Tn[10].t20 VGND 0.01692f
C6368 XThR.Tn[10].n44 VGND 0.04313f
C6369 XThR.Tn[10].n45 VGND 0.0303f
C6370 XThR.Tn[10].n47 VGND 0.09724f
C6371 XThR.Tn[10].t33 VGND 0.0155f
C6372 XThR.Tn[10].t43 VGND 0.01698f
C6373 XThR.Tn[10].n48 VGND 0.04146f
C6374 XThR.Tn[10].t73 VGND 0.01545f
C6375 XThR.Tn[10].t38 VGND 0.01692f
C6376 XThR.Tn[10].n49 VGND 0.04313f
C6377 XThR.Tn[10].n50 VGND 0.0303f
C6378 XThR.Tn[10].n52 VGND 0.09724f
C6379 XThR.Tn[10].t28 VGND 0.0155f
C6380 XThR.Tn[10].t61 VGND 0.01698f
C6381 XThR.Tn[10].n53 VGND 0.04146f
C6382 XThR.Tn[10].t62 VGND 0.01545f
C6383 XThR.Tn[10].t57 VGND 0.01692f
C6384 XThR.Tn[10].n54 VGND 0.04313f
C6385 XThR.Tn[10].n55 VGND 0.0303f
C6386 XThR.Tn[10].n57 VGND 0.09724f
C6387 XThR.Tn[10].t46 VGND 0.0155f
C6388 XThR.Tn[10].t35 VGND 0.01698f
C6389 XThR.Tn[10].n58 VGND 0.04146f
C6390 XThR.Tn[10].t19 VGND 0.01545f
C6391 XThR.Tn[10].t32 VGND 0.01692f
C6392 XThR.Tn[10].n59 VGND 0.04313f
C6393 XThR.Tn[10].n60 VGND 0.0303f
C6394 XThR.Tn[10].n62 VGND 0.09724f
C6395 XThR.Tn[10].t16 VGND 0.0155f
C6396 XThR.Tn[10].t72 VGND 0.01698f
C6397 XThR.Tn[10].n63 VGND 0.04146f
C6398 XThR.Tn[10].t52 VGND 0.01545f
C6399 XThR.Tn[10].t68 VGND 0.01692f
C6400 XThR.Tn[10].n64 VGND 0.04313f
C6401 XThR.Tn[10].n65 VGND 0.0303f
C6402 XThR.Tn[10].n67 VGND 0.09724f
C6403 XThR.Tn[10].t31 VGND 0.0155f
C6404 XThR.Tn[10].t27 VGND 0.01698f
C6405 XThR.Tn[10].n68 VGND 0.04146f
C6406 XThR.Tn[10].t71 VGND 0.01545f
C6407 XThR.Tn[10].t22 VGND 0.01692f
C6408 XThR.Tn[10].n69 VGND 0.04313f
C6409 XThR.Tn[10].n70 VGND 0.0303f
C6410 XThR.Tn[10].n72 VGND 0.09724f
C6411 XThR.Tn[10].t49 VGND 0.0155f
C6412 XThR.Tn[10].t45 VGND 0.01698f
C6413 XThR.Tn[10].n73 VGND 0.04146f
C6414 XThR.Tn[10].t25 VGND 0.01545f
C6415 XThR.Tn[10].t39 VGND 0.01692f
C6416 XThR.Tn[10].n74 VGND 0.04313f
C6417 XThR.Tn[10].n75 VGND 0.0303f
C6418 XThR.Tn[10].n77 VGND 0.09724f
C6419 XThR.Tn[10].t29 VGND 0.0155f
C6420 XThR.Tn[10].t37 VGND 0.01698f
C6421 XThR.Tn[10].n78 VGND 0.04146f
C6422 XThR.Tn[10].t64 VGND 0.01545f
C6423 XThR.Tn[10].t34 VGND 0.01692f
C6424 XThR.Tn[10].n79 VGND 0.04313f
C6425 XThR.Tn[10].n80 VGND 0.0303f
C6426 XThR.Tn[10].n82 VGND 0.09724f
C6427 XThR.Tn[10].n83 VGND 0.08837f
C6428 XThR.Tn[10].n84 VGND 0.27206f
C6429 XThR.Tn[10].t4 VGND 0.01984f
C6430 XThR.Tn[10].t5 VGND 0.01984f
C6431 XThR.Tn[10].n85 VGND 0.04286f
C6432 XThR.Tn[10].t1 VGND 0.01984f
C6433 XThR.Tn[10].t0 VGND 0.01984f
C6434 XThR.Tn[10].n86 VGND 0.06524f
C6435 XThR.Tn[10].n87 VGND 0.18114f
C6436 XThC.Tn[3].t5 VGND 0.01413f
C6437 XThC.Tn[3].t4 VGND 0.01413f
C6438 XThC.Tn[3].n0 VGND 0.02852f
C6439 XThC.Tn[3].t7 VGND 0.01413f
C6440 XThC.Tn[3].t6 VGND 0.01413f
C6441 XThC.Tn[3].n1 VGND 0.03337f
C6442 XThC.Tn[3].n2 VGND 0.10009f
C6443 XThC.Tn[3].n3 VGND 0.02091f
C6444 XThC.Tn[3].n4 VGND 0.03484f
C6445 XThC.Tn[3].n5 VGND 0.02091f
C6446 XThC.Tn[3].n6 VGND 0.09959f
C6447 XThC.Tn[3].n7 VGND 0.02091f
C6448 XThC.Tn[3].n8 VGND 0.06156f
C6449 XThC.Tn[3].n9 VGND 0.06948f
C6450 XThC.Tn[3].t12 VGND 0.0112f
C6451 XThC.Tn[3].t42 VGND 0.01223f
C6452 XThC.Tn[3].n10 VGND 0.0273f
C6453 XThC.Tn[3].n11 VGND 0.01871f
C6454 XThC.Tn[3].n12 VGND 0.0614f
C6455 XThC.Tn[3].t30 VGND 0.0112f
C6456 XThC.Tn[3].t27 VGND 0.01223f
C6457 XThC.Tn[3].n13 VGND 0.0273f
C6458 XThC.Tn[3].n14 VGND 0.01871f
C6459 XThC.Tn[3].n15 VGND 0.06157f
C6460 XThC.Tn[3].n16 VGND 0.10147f
C6461 XThC.Tn[3].t35 VGND 0.0112f
C6462 XThC.Tn[3].t29 VGND 0.01223f
C6463 XThC.Tn[3].n17 VGND 0.0273f
C6464 XThC.Tn[3].n18 VGND 0.01871f
C6465 XThC.Tn[3].n19 VGND 0.06157f
C6466 XThC.Tn[3].n20 VGND 0.10147f
C6467 XThC.Tn[3].t36 VGND 0.0112f
C6468 XThC.Tn[3].t31 VGND 0.01223f
C6469 XThC.Tn[3].n21 VGND 0.0273f
C6470 XThC.Tn[3].n22 VGND 0.01871f
C6471 XThC.Tn[3].n23 VGND 0.06157f
C6472 XThC.Tn[3].n24 VGND 0.10147f
C6473 XThC.Tn[3].t23 VGND 0.0112f
C6474 XThC.Tn[3].t20 VGND 0.01223f
C6475 XThC.Tn[3].n25 VGND 0.0273f
C6476 XThC.Tn[3].n26 VGND 0.01871f
C6477 XThC.Tn[3].n27 VGND 0.06157f
C6478 XThC.Tn[3].n28 VGND 0.10147f
C6479 XThC.Tn[3].t24 VGND 0.0112f
C6480 XThC.Tn[3].t21 VGND 0.01223f
C6481 XThC.Tn[3].n29 VGND 0.0273f
C6482 XThC.Tn[3].n30 VGND 0.01871f
C6483 XThC.Tn[3].n31 VGND 0.06157f
C6484 XThC.Tn[3].n32 VGND 0.10147f
C6485 XThC.Tn[3].t40 VGND 0.0112f
C6486 XThC.Tn[3].t34 VGND 0.01223f
C6487 XThC.Tn[3].n33 VGND 0.0273f
C6488 XThC.Tn[3].n34 VGND 0.01871f
C6489 XThC.Tn[3].n35 VGND 0.06157f
C6490 XThC.Tn[3].n36 VGND 0.10147f
C6491 XThC.Tn[3].t15 VGND 0.0112f
C6492 XThC.Tn[3].t43 VGND 0.01223f
C6493 XThC.Tn[3].n37 VGND 0.0273f
C6494 XThC.Tn[3].n38 VGND 0.01871f
C6495 XThC.Tn[3].n39 VGND 0.06157f
C6496 XThC.Tn[3].n40 VGND 0.10147f
C6497 XThC.Tn[3].t17 VGND 0.0112f
C6498 XThC.Tn[3].t13 VGND 0.01223f
C6499 XThC.Tn[3].n41 VGND 0.0273f
C6500 XThC.Tn[3].n42 VGND 0.01871f
C6501 XThC.Tn[3].n43 VGND 0.06157f
C6502 XThC.Tn[3].n44 VGND 0.10147f
C6503 XThC.Tn[3].t37 VGND 0.0112f
C6504 XThC.Tn[3].t32 VGND 0.01223f
C6505 XThC.Tn[3].n45 VGND 0.0273f
C6506 XThC.Tn[3].n46 VGND 0.01871f
C6507 XThC.Tn[3].n47 VGND 0.06157f
C6508 XThC.Tn[3].n48 VGND 0.10147f
C6509 XThC.Tn[3].t39 VGND 0.0112f
C6510 XThC.Tn[3].t33 VGND 0.01223f
C6511 XThC.Tn[3].n49 VGND 0.0273f
C6512 XThC.Tn[3].n50 VGND 0.01871f
C6513 XThC.Tn[3].n51 VGND 0.06157f
C6514 XThC.Tn[3].n52 VGND 0.10147f
C6515 XThC.Tn[3].t18 VGND 0.0112f
C6516 XThC.Tn[3].t14 VGND 0.01223f
C6517 XThC.Tn[3].n53 VGND 0.0273f
C6518 XThC.Tn[3].n54 VGND 0.01871f
C6519 XThC.Tn[3].n55 VGND 0.06157f
C6520 XThC.Tn[3].n56 VGND 0.10147f
C6521 XThC.Tn[3].t26 VGND 0.0112f
C6522 XThC.Tn[3].t22 VGND 0.01223f
C6523 XThC.Tn[3].n57 VGND 0.0273f
C6524 XThC.Tn[3].n58 VGND 0.01871f
C6525 XThC.Tn[3].n59 VGND 0.06157f
C6526 XThC.Tn[3].n60 VGND 0.10147f
C6527 XThC.Tn[3].t28 VGND 0.0112f
C6528 XThC.Tn[3].t25 VGND 0.01223f
C6529 XThC.Tn[3].n61 VGND 0.0273f
C6530 XThC.Tn[3].n62 VGND 0.01871f
C6531 XThC.Tn[3].n63 VGND 0.06157f
C6532 XThC.Tn[3].n64 VGND 0.10147f
C6533 XThC.Tn[3].t41 VGND 0.0112f
C6534 XThC.Tn[3].t38 VGND 0.01223f
C6535 XThC.Tn[3].n65 VGND 0.0273f
C6536 XThC.Tn[3].n66 VGND 0.01871f
C6537 XThC.Tn[3].n67 VGND 0.06157f
C6538 XThC.Tn[3].n68 VGND 0.10147f
C6539 XThC.Tn[3].t19 VGND 0.0112f
C6540 XThC.Tn[3].t16 VGND 0.01223f
C6541 XThC.Tn[3].n69 VGND 0.0273f
C6542 XThC.Tn[3].n70 VGND 0.01871f
C6543 XThC.Tn[3].n71 VGND 0.06157f
C6544 XThC.Tn[3].n72 VGND 0.10147f
C6545 XThC.Tn[3].n73 VGND 0.59675f
C6546 XThC.Tn[3].n74 VGND 0.08605f
C6547 XThC.Tn[1].t3 VGND 0.01343f
C6548 XThC.Tn[1].t2 VGND 0.01343f
C6549 XThC.Tn[1].n0 VGND 0.02712f
C6550 XThC.Tn[1].t1 VGND 0.01343f
C6551 XThC.Tn[1].t0 VGND 0.01343f
C6552 XThC.Tn[1].n1 VGND 0.03173f
C6553 XThC.Tn[1].n2 VGND 0.09517f
C6554 XThC.Tn[1].n3 VGND 0.03313f
C6555 XThC.Tn[1].n4 VGND 0.01988f
C6556 XThC.Tn[1].n5 VGND 0.09469f
C6557 XThC.Tn[1].n6 VGND 0.01988f
C6558 XThC.Tn[1].n7 VGND 0.05854f
C6559 XThC.Tn[1].n8 VGND 0.01988f
C6560 XThC.Tn[1].n9 VGND 0.06606f
C6561 XThC.Tn[1].t31 VGND 0.01065f
C6562 XThC.Tn[1].t29 VGND 0.01163f
C6563 XThC.Tn[1].n10 VGND 0.02596f
C6564 XThC.Tn[1].n11 VGND 0.01779f
C6565 XThC.Tn[1].n12 VGND 0.05838f
C6566 XThC.Tn[1].t17 VGND 0.01065f
C6567 XThC.Tn[1].t14 VGND 0.01163f
C6568 XThC.Tn[1].n13 VGND 0.02596f
C6569 XThC.Tn[1].n14 VGND 0.01779f
C6570 XThC.Tn[1].n15 VGND 0.05854f
C6571 XThC.Tn[1].n16 VGND 0.09648f
C6572 XThC.Tn[1].t22 VGND 0.01065f
C6573 XThC.Tn[1].t16 VGND 0.01163f
C6574 XThC.Tn[1].n17 VGND 0.02596f
C6575 XThC.Tn[1].n18 VGND 0.01779f
C6576 XThC.Tn[1].n19 VGND 0.05854f
C6577 XThC.Tn[1].n20 VGND 0.09648f
C6578 XThC.Tn[1].t23 VGND 0.01065f
C6579 XThC.Tn[1].t18 VGND 0.01163f
C6580 XThC.Tn[1].n21 VGND 0.02596f
C6581 XThC.Tn[1].n22 VGND 0.01779f
C6582 XThC.Tn[1].n23 VGND 0.05854f
C6583 XThC.Tn[1].n24 VGND 0.09648f
C6584 XThC.Tn[1].t42 VGND 0.01065f
C6585 XThC.Tn[1].t39 VGND 0.01163f
C6586 XThC.Tn[1].n25 VGND 0.02596f
C6587 XThC.Tn[1].n26 VGND 0.01779f
C6588 XThC.Tn[1].n27 VGND 0.05854f
C6589 XThC.Tn[1].n28 VGND 0.09648f
C6590 XThC.Tn[1].t43 VGND 0.01065f
C6591 XThC.Tn[1].t40 VGND 0.01163f
C6592 XThC.Tn[1].n29 VGND 0.02596f
C6593 XThC.Tn[1].n30 VGND 0.01779f
C6594 XThC.Tn[1].n31 VGND 0.05854f
C6595 XThC.Tn[1].n32 VGND 0.09648f
C6596 XThC.Tn[1].t27 VGND 0.01065f
C6597 XThC.Tn[1].t21 VGND 0.01163f
C6598 XThC.Tn[1].n33 VGND 0.02596f
C6599 XThC.Tn[1].n34 VGND 0.01779f
C6600 XThC.Tn[1].n35 VGND 0.05854f
C6601 XThC.Tn[1].n36 VGND 0.09648f
C6602 XThC.Tn[1].t34 VGND 0.01065f
C6603 XThC.Tn[1].t30 VGND 0.01163f
C6604 XThC.Tn[1].n37 VGND 0.02596f
C6605 XThC.Tn[1].n38 VGND 0.01779f
C6606 XThC.Tn[1].n39 VGND 0.05854f
C6607 XThC.Tn[1].n40 VGND 0.09648f
C6608 XThC.Tn[1].t36 VGND 0.01065f
C6609 XThC.Tn[1].t32 VGND 0.01163f
C6610 XThC.Tn[1].n41 VGND 0.02596f
C6611 XThC.Tn[1].n42 VGND 0.01779f
C6612 XThC.Tn[1].n43 VGND 0.05854f
C6613 XThC.Tn[1].n44 VGND 0.09648f
C6614 XThC.Tn[1].t24 VGND 0.01065f
C6615 XThC.Tn[1].t19 VGND 0.01163f
C6616 XThC.Tn[1].n45 VGND 0.02596f
C6617 XThC.Tn[1].n46 VGND 0.01779f
C6618 XThC.Tn[1].n47 VGND 0.05854f
C6619 XThC.Tn[1].n48 VGND 0.09648f
C6620 XThC.Tn[1].t26 VGND 0.01065f
C6621 XThC.Tn[1].t20 VGND 0.01163f
C6622 XThC.Tn[1].n49 VGND 0.02596f
C6623 XThC.Tn[1].n50 VGND 0.01779f
C6624 XThC.Tn[1].n51 VGND 0.05854f
C6625 XThC.Tn[1].n52 VGND 0.09648f
C6626 XThC.Tn[1].t37 VGND 0.01065f
C6627 XThC.Tn[1].t33 VGND 0.01163f
C6628 XThC.Tn[1].n53 VGND 0.02596f
C6629 XThC.Tn[1].n54 VGND 0.01779f
C6630 XThC.Tn[1].n55 VGND 0.05854f
C6631 XThC.Tn[1].n56 VGND 0.09648f
C6632 XThC.Tn[1].t13 VGND 0.01065f
C6633 XThC.Tn[1].t41 VGND 0.01163f
C6634 XThC.Tn[1].n57 VGND 0.02596f
C6635 XThC.Tn[1].n58 VGND 0.01779f
C6636 XThC.Tn[1].n59 VGND 0.05854f
C6637 XThC.Tn[1].n60 VGND 0.09648f
C6638 XThC.Tn[1].t15 VGND 0.01065f
C6639 XThC.Tn[1].t12 VGND 0.01163f
C6640 XThC.Tn[1].n61 VGND 0.02596f
C6641 XThC.Tn[1].n62 VGND 0.01779f
C6642 XThC.Tn[1].n63 VGND 0.05854f
C6643 XThC.Tn[1].n64 VGND 0.09648f
C6644 XThC.Tn[1].t28 VGND 0.01065f
C6645 XThC.Tn[1].t25 VGND 0.01163f
C6646 XThC.Tn[1].n65 VGND 0.02596f
C6647 XThC.Tn[1].n66 VGND 0.01779f
C6648 XThC.Tn[1].n67 VGND 0.05854f
C6649 XThC.Tn[1].n68 VGND 0.09648f
C6650 XThC.Tn[1].t38 VGND 0.01065f
C6651 XThC.Tn[1].t35 VGND 0.01163f
C6652 XThC.Tn[1].n69 VGND 0.02596f
C6653 XThC.Tn[1].n70 VGND 0.01779f
C6654 XThC.Tn[1].n71 VGND 0.05854f
C6655 XThC.Tn[1].n72 VGND 0.09648f
C6656 XThC.Tn[1].n73 VGND 0.49027f
C6657 XThC.Tn[1].n74 VGND 0.09316f
C6658 Vbias.t260 VGND 0.17892f
C6659 Vbias.n0 VGND 0.19478f
C6660 Vbias.t79 VGND 0.17892f
C6661 Vbias.n1 VGND 0.19512f
C6662 Vbias.n2 VGND 0.1294f
C6663 Vbias.t174 VGND 0.17892f
C6664 Vbias.n3 VGND 0.19512f
C6665 Vbias.n4 VGND 0.1294f
C6666 Vbias.t182 VGND 0.17892f
C6667 Vbias.n5 VGND 0.19512f
C6668 Vbias.n6 VGND 0.1294f
C6669 Vbias.t15 VGND 0.17892f
C6670 Vbias.n7 VGND 0.19512f
C6671 Vbias.n8 VGND 0.1294f
C6672 Vbias.t101 VGND 0.17892f
C6673 Vbias.n9 VGND 0.19512f
C6674 Vbias.n10 VGND 0.1294f
C6675 Vbias.t184 VGND 0.17892f
C6676 Vbias.n11 VGND 0.19512f
C6677 Vbias.n12 VGND 0.1294f
C6678 Vbias.t19 VGND 0.17892f
C6679 Vbias.n13 VGND 0.19512f
C6680 Vbias.n14 VGND 0.1294f
C6681 Vbias.t39 VGND 0.17892f
C6682 Vbias.n15 VGND 0.19512f
C6683 Vbias.n16 VGND 0.1294f
C6684 Vbias.t111 VGND 0.17892f
C6685 Vbias.n17 VGND 0.19512f
C6686 Vbias.n18 VGND 0.1294f
C6687 Vbias.t202 VGND 0.17892f
C6688 Vbias.n19 VGND 0.19512f
C6689 Vbias.n20 VGND 0.1294f
C6690 Vbias.t223 VGND 0.17892f
C6691 Vbias.n21 VGND 0.19512f
C6692 Vbias.n22 VGND 0.1294f
C6693 Vbias.t114 VGND 0.17892f
C6694 Vbias.n23 VGND 0.19512f
C6695 Vbias.n24 VGND 0.1294f
C6696 Vbias.t142 VGND 0.17892f
C6697 Vbias.n25 VGND 0.19512f
C6698 Vbias.n26 VGND 0.1294f
C6699 Vbias.t151 VGND 0.17892f
C6700 Vbias.n27 VGND 0.19512f
C6701 Vbias.n28 VGND 0.1294f
C6702 Vbias.t61 VGND 0.17892f
C6703 Vbias.n29 VGND 0.19512f
C6704 Vbias.n30 VGND 0.1294f
C6705 Vbias.n31 VGND 0.54301f
C6706 Vbias.t140 VGND 0.17892f
C6707 Vbias.n32 VGND 0.19478f
C6708 Vbias.t216 VGND 0.17892f
C6709 Vbias.n33 VGND 0.19512f
C6710 Vbias.n34 VGND 0.1294f
C6711 Vbias.t59 VGND 0.17892f
C6712 Vbias.n35 VGND 0.19512f
C6713 Vbias.n36 VGND 0.1294f
C6714 Vbias.t67 VGND 0.17892f
C6715 Vbias.n37 VGND 0.19512f
C6716 Vbias.n38 VGND 0.1294f
C6717 Vbias.t152 VGND 0.17892f
C6718 Vbias.n39 VGND 0.19512f
C6719 Vbias.n40 VGND 0.1294f
C6720 Vbias.t245 VGND 0.17892f
C6721 Vbias.n41 VGND 0.19512f
C6722 Vbias.n42 VGND 0.1294f
C6723 Vbias.t72 VGND 0.17892f
C6724 Vbias.n43 VGND 0.19512f
C6725 Vbias.n44 VGND 0.1294f
C6726 Vbias.t158 VGND 0.17892f
C6727 Vbias.n45 VGND 0.19512f
C6728 Vbias.n46 VGND 0.1294f
C6729 Vbias.t178 VGND 0.17892f
C6730 Vbias.n47 VGND 0.19512f
C6731 Vbias.n48 VGND 0.1294f
C6732 Vbias.t254 VGND 0.17892f
C6733 Vbias.n49 VGND 0.19512f
C6734 Vbias.n50 VGND 0.1294f
C6735 Vbias.t84 VGND 0.17892f
C6736 Vbias.n51 VGND 0.19512f
C6737 Vbias.n52 VGND 0.1294f
C6738 Vbias.t106 VGND 0.17892f
C6739 Vbias.n53 VGND 0.19512f
C6740 Vbias.n54 VGND 0.1294f
C6741 Vbias.t259 VGND 0.17892f
C6742 Vbias.n55 VGND 0.19512f
C6743 Vbias.n56 VGND 0.1294f
C6744 Vbias.t26 VGND 0.17892f
C6745 Vbias.n57 VGND 0.19512f
C6746 Vbias.n58 VGND 0.1294f
C6747 Vbias.t35 VGND 0.17892f
C6748 Vbias.n59 VGND 0.19512f
C6749 Vbias.n60 VGND 0.1294f
C6750 Vbias.t194 VGND 0.17892f
C6751 Vbias.n61 VGND 0.19512f
C6752 Vbias.n62 VGND 0.1294f
C6753 Vbias.n63 VGND 0.55864f
C6754 Vbias.t215 VGND 0.17892f
C6755 Vbias.n64 VGND 0.19478f
C6756 Vbias.t31 VGND 0.17892f
C6757 Vbias.n65 VGND 0.19512f
C6758 Vbias.n66 VGND 0.1294f
C6759 Vbias.t132 VGND 0.17892f
C6760 Vbias.n67 VGND 0.19512f
C6761 Vbias.n68 VGND 0.1294f
C6762 Vbias.t139 VGND 0.17892f
C6763 Vbias.n69 VGND 0.19512f
C6764 Vbias.n70 VGND 0.1294f
C6765 Vbias.t224 VGND 0.17892f
C6766 Vbias.n71 VGND 0.19512f
C6767 Vbias.n72 VGND 0.1294f
C6768 Vbias.t58 VGND 0.17892f
C6769 Vbias.n73 VGND 0.19512f
C6770 Vbias.n74 VGND 0.1294f
C6771 Vbias.t145 VGND 0.17892f
C6772 Vbias.n75 VGND 0.19512f
C6773 Vbias.n76 VGND 0.1294f
C6774 Vbias.t230 VGND 0.17892f
C6775 Vbias.n77 VGND 0.19512f
C6776 Vbias.n78 VGND 0.1294f
C6777 Vbias.t253 VGND 0.17892f
C6778 Vbias.n79 VGND 0.19512f
C6779 Vbias.n80 VGND 0.1294f
C6780 Vbias.t71 VGND 0.17892f
C6781 Vbias.n81 VGND 0.19512f
C6782 Vbias.n82 VGND 0.1294f
C6783 Vbias.t157 VGND 0.17892f
C6784 Vbias.n83 VGND 0.19512f
C6785 Vbias.n84 VGND 0.1294f
C6786 Vbias.t177 VGND 0.17892f
C6787 Vbias.n85 VGND 0.19512f
C6788 Vbias.n86 VGND 0.1294f
C6789 Vbias.t77 VGND 0.17892f
C6790 Vbias.n87 VGND 0.19512f
C6791 Vbias.n88 VGND 0.1294f
C6792 Vbias.t97 VGND 0.17892f
C6793 Vbias.n89 VGND 0.19512f
C6794 Vbias.n90 VGND 0.1294f
C6795 Vbias.t104 VGND 0.17892f
C6796 Vbias.n91 VGND 0.19512f
C6797 Vbias.n92 VGND 0.1294f
C6798 Vbias.t13 VGND 0.17892f
C6799 Vbias.n93 VGND 0.19512f
C6800 Vbias.n94 VGND 0.1294f
C6801 Vbias.n95 VGND 0.55864f
C6802 Vbias.t30 VGND 0.17892f
C6803 Vbias.n96 VGND 0.19478f
C6804 Vbias.t100 VGND 0.17892f
C6805 Vbias.n97 VGND 0.19512f
C6806 Vbias.n98 VGND 0.1294f
C6807 Vbias.t203 VGND 0.17892f
C6808 Vbias.n99 VGND 0.19512f
C6809 Vbias.n100 VGND 0.1294f
C6810 Vbias.t214 VGND 0.17892f
C6811 Vbias.n101 VGND 0.19512f
C6812 Vbias.n102 VGND 0.1294f
C6813 Vbias.t38 VGND 0.17892f
C6814 Vbias.n103 VGND 0.19512f
C6815 Vbias.n104 VGND 0.1294f
C6816 Vbias.t131 VGND 0.17892f
C6817 Vbias.n105 VGND 0.19512f
C6818 Vbias.n106 VGND 0.1294f
C6819 Vbias.t218 VGND 0.17892f
C6820 Vbias.n107 VGND 0.19512f
C6821 Vbias.n108 VGND 0.1294f
C6822 Vbias.t42 VGND 0.17892f
C6823 Vbias.n109 VGND 0.19512f
C6824 Vbias.n110 VGND 0.1294f
C6825 Vbias.t70 VGND 0.17892f
C6826 Vbias.n111 VGND 0.19512f
C6827 Vbias.n112 VGND 0.1294f
C6828 Vbias.t143 VGND 0.17892f
C6829 Vbias.n113 VGND 0.19512f
C6830 Vbias.n114 VGND 0.1294f
C6831 Vbias.t228 VGND 0.17892f
C6832 Vbias.n115 VGND 0.19512f
C6833 Vbias.n116 VGND 0.1294f
C6834 Vbias.t252 VGND 0.17892f
C6835 Vbias.n117 VGND 0.19512f
C6836 Vbias.n118 VGND 0.1294f
C6837 Vbias.t148 VGND 0.17892f
C6838 Vbias.n119 VGND 0.19512f
C6839 Vbias.n120 VGND 0.1294f
C6840 Vbias.t170 VGND 0.17892f
C6841 Vbias.n121 VGND 0.19512f
C6842 Vbias.n122 VGND 0.1294f
C6843 Vbias.t175 VGND 0.17892f
C6844 Vbias.n123 VGND 0.19512f
C6845 Vbias.n124 VGND 0.1294f
C6846 Vbias.t86 VGND 0.17892f
C6847 Vbias.n125 VGND 0.19512f
C6848 Vbias.n126 VGND 0.1294f
C6849 Vbias.n127 VGND 0.55864f
C6850 Vbias.t186 VGND 0.17892f
C6851 Vbias.n128 VGND 0.19478f
C6852 Vbias.t6 VGND 0.17892f
C6853 Vbias.n129 VGND 0.19512f
C6854 Vbias.n130 VGND 0.1294f
C6855 Vbias.t103 VGND 0.17892f
C6856 Vbias.n131 VGND 0.19512f
C6857 Vbias.n132 VGND 0.1294f
C6858 Vbias.t115 VGND 0.17892f
C6859 Vbias.n133 VGND 0.19512f
C6860 Vbias.n134 VGND 0.1294f
C6861 Vbias.t206 VGND 0.17892f
C6862 Vbias.n135 VGND 0.19512f
C6863 Vbias.n136 VGND 0.1294f
C6864 Vbias.t34 VGND 0.17892f
C6865 Vbias.n137 VGND 0.19512f
C6866 Vbias.n138 VGND 0.1294f
C6867 Vbias.t116 VGND 0.17892f
C6868 Vbias.n139 VGND 0.19512f
C6869 Vbias.n140 VGND 0.1294f
C6870 Vbias.t209 VGND 0.17892f
C6871 Vbias.n141 VGND 0.19512f
C6872 Vbias.n142 VGND 0.1294f
C6873 Vbias.t231 VGND 0.17892f
C6874 Vbias.n143 VGND 0.19512f
C6875 Vbias.n144 VGND 0.1294f
C6876 Vbias.t43 VGND 0.17892f
C6877 Vbias.n145 VGND 0.19512f
C6878 Vbias.n146 VGND 0.1294f
C6879 Vbias.t134 VGND 0.17892f
C6880 Vbias.n147 VGND 0.19512f
C6881 Vbias.n148 VGND 0.1294f
C6882 Vbias.t159 VGND 0.17892f
C6883 Vbias.n149 VGND 0.19512f
C6884 Vbias.n150 VGND 0.1294f
C6885 Vbias.t47 VGND 0.17892f
C6886 Vbias.n151 VGND 0.19512f
C6887 Vbias.n152 VGND 0.1294f
C6888 Vbias.t78 VGND 0.17892f
C6889 Vbias.n153 VGND 0.19512f
C6890 Vbias.n154 VGND 0.1294f
C6891 Vbias.t85 VGND 0.17892f
C6892 Vbias.n155 VGND 0.19512f
C6893 Vbias.n156 VGND 0.1294f
C6894 Vbias.t249 VGND 0.17892f
C6895 Vbias.n157 VGND 0.19512f
C6896 Vbias.n158 VGND 0.1294f
C6897 Vbias.n159 VGND 0.55864f
C6898 Vbias.t55 VGND 0.17892f
C6899 Vbias.n160 VGND 0.19478f
C6900 Vbias.t128 VGND 0.17892f
C6901 Vbias.n161 VGND 0.19512f
C6902 Vbias.n162 VGND 0.1294f
C6903 Vbias.t226 VGND 0.17892f
C6904 Vbias.n163 VGND 0.19512f
C6905 Vbias.n164 VGND 0.1294f
C6906 Vbias.t241 VGND 0.17892f
C6907 Vbias.n165 VGND 0.19512f
C6908 Vbias.n166 VGND 0.1294f
C6909 Vbias.t66 VGND 0.17892f
C6910 Vbias.n167 VGND 0.19512f
C6911 Vbias.n168 VGND 0.1294f
C6912 Vbias.t155 VGND 0.17892f
C6913 Vbias.n169 VGND 0.19512f
C6914 Vbias.n170 VGND 0.1294f
C6915 Vbias.t244 VGND 0.17892f
C6916 Vbias.n171 VGND 0.19512f
C6917 Vbias.n172 VGND 0.1294f
C6918 Vbias.t74 VGND 0.17892f
C6919 Vbias.n173 VGND 0.19512f
C6920 Vbias.n174 VGND 0.1294f
C6921 Vbias.t94 VGND 0.17892f
C6922 Vbias.n175 VGND 0.19512f
C6923 Vbias.n176 VGND 0.1294f
C6924 Vbias.t167 VGND 0.17892f
C6925 Vbias.n177 VGND 0.19512f
C6926 Vbias.n178 VGND 0.1294f
C6927 Vbias.t256 VGND 0.17892f
C6928 Vbias.n179 VGND 0.19512f
C6929 Vbias.n180 VGND 0.1294f
C6930 Vbias.t22 VGND 0.17892f
C6931 Vbias.n181 VGND 0.19512f
C6932 Vbias.n182 VGND 0.1294f
C6933 Vbias.t172 VGND 0.17892f
C6934 Vbias.n183 VGND 0.19512f
C6935 Vbias.n184 VGND 0.1294f
C6936 Vbias.t191 VGND 0.17892f
C6937 Vbias.n185 VGND 0.19512f
C6938 Vbias.n186 VGND 0.1294f
C6939 Vbias.t207 VGND 0.17892f
C6940 Vbias.n187 VGND 0.19512f
C6941 Vbias.n188 VGND 0.1294f
C6942 Vbias.t109 VGND 0.17892f
C6943 Vbias.n189 VGND 0.19512f
C6944 Vbias.n190 VGND 0.1294f
C6945 Vbias.n191 VGND 0.55864f
C6946 Vbias.t189 VGND 0.17892f
C6947 Vbias.n192 VGND 0.19478f
C6948 Vbias.t10 VGND 0.17892f
C6949 Vbias.n193 VGND 0.19512f
C6950 Vbias.n194 VGND 0.1294f
C6951 Vbias.t108 VGND 0.17892f
C6952 Vbias.n195 VGND 0.19512f
C6953 Vbias.n196 VGND 0.1294f
C6954 Vbias.t117 VGND 0.17892f
C6955 Vbias.n197 VGND 0.19512f
C6956 Vbias.n198 VGND 0.1294f
C6957 Vbias.t208 VGND 0.17892f
C6958 Vbias.n199 VGND 0.19512f
C6959 Vbias.n200 VGND 0.1294f
C6960 Vbias.t36 VGND 0.17892f
C6961 Vbias.n201 VGND 0.19512f
C6962 Vbias.n202 VGND 0.1294f
C6963 Vbias.t120 VGND 0.17892f
C6964 Vbias.n203 VGND 0.19512f
C6965 Vbias.n204 VGND 0.1294f
C6966 Vbias.t212 VGND 0.17892f
C6967 Vbias.n205 VGND 0.19512f
C6968 Vbias.n206 VGND 0.1294f
C6969 Vbias.t234 VGND 0.17892f
C6970 Vbias.n207 VGND 0.19512f
C6971 Vbias.n208 VGND 0.1294f
C6972 Vbias.t46 VGND 0.17892f
C6973 Vbias.n209 VGND 0.19512f
C6974 Vbias.n210 VGND 0.1294f
C6975 Vbias.t136 VGND 0.17892f
C6976 Vbias.n211 VGND 0.19512f
C6977 Vbias.n212 VGND 0.1294f
C6978 Vbias.t162 VGND 0.17892f
C6979 Vbias.n213 VGND 0.19512f
C6980 Vbias.n214 VGND 0.1294f
C6981 Vbias.t51 VGND 0.17892f
C6982 Vbias.n215 VGND 0.19512f
C6983 Vbias.n216 VGND 0.1294f
C6984 Vbias.t80 VGND 0.17892f
C6985 Vbias.n217 VGND 0.19512f
C6986 Vbias.n218 VGND 0.1294f
C6987 Vbias.t89 VGND 0.17892f
C6988 Vbias.n219 VGND 0.19512f
C6989 Vbias.n220 VGND 0.1294f
C6990 Vbias.t250 VGND 0.17892f
C6991 Vbias.n221 VGND 0.19512f
C6992 Vbias.n222 VGND 0.1294f
C6993 Vbias.n223 VGND 0.55864f
C6994 Vbias.t9 VGND 0.17892f
C6995 Vbias.n224 VGND 0.19478f
C6996 Vbias.t83 VGND 0.17892f
C6997 Vbias.n225 VGND 0.19512f
C6998 Vbias.n226 VGND 0.1294f
C6999 Vbias.t180 VGND 0.17892f
C7000 Vbias.n227 VGND 0.19512f
C7001 Vbias.n228 VGND 0.1294f
C7002 Vbias.t188 VGND 0.17892f
C7003 Vbias.n229 VGND 0.19512f
C7004 Vbias.n230 VGND 0.1294f
C7005 Vbias.t23 VGND 0.17892f
C7006 Vbias.n231 VGND 0.19512f
C7007 Vbias.n232 VGND 0.1294f
C7008 Vbias.t107 VGND 0.17892f
C7009 Vbias.n233 VGND 0.19512f
C7010 Vbias.n234 VGND 0.1294f
C7011 Vbias.t192 VGND 0.17892f
C7012 Vbias.n235 VGND 0.19512f
C7013 Vbias.n236 VGND 0.1294f
C7014 Vbias.t28 VGND 0.17892f
C7015 Vbias.n237 VGND 0.19512f
C7016 Vbias.n238 VGND 0.1294f
C7017 Vbias.t45 VGND 0.17892f
C7018 Vbias.n239 VGND 0.19512f
C7019 Vbias.n240 VGND 0.1294f
C7020 Vbias.t119 VGND 0.17892f
C7021 Vbias.n241 VGND 0.19512f
C7022 Vbias.n242 VGND 0.1294f
C7023 Vbias.t211 VGND 0.17892f
C7024 Vbias.n243 VGND 0.19512f
C7025 Vbias.n244 VGND 0.1294f
C7026 Vbias.t233 VGND 0.17892f
C7027 Vbias.n245 VGND 0.19512f
C7028 Vbias.n246 VGND 0.1294f
C7029 Vbias.t123 VGND 0.17892f
C7030 Vbias.n247 VGND 0.19512f
C7031 Vbias.n248 VGND 0.1294f
C7032 Vbias.t149 VGND 0.17892f
C7033 Vbias.n249 VGND 0.19512f
C7034 Vbias.n250 VGND 0.1294f
C7035 Vbias.t161 VGND 0.17892f
C7036 Vbias.n251 VGND 0.19512f
C7037 Vbias.n252 VGND 0.1294f
C7038 Vbias.t64 VGND 0.17892f
C7039 Vbias.n253 VGND 0.19512f
C7040 Vbias.n254 VGND 0.1294f
C7041 Vbias.n255 VGND 0.55864f
C7042 Vbias.t82 VGND 0.17892f
C7043 Vbias.n256 VGND 0.19478f
C7044 Vbias.t154 VGND 0.17892f
C7045 Vbias.n257 VGND 0.19512f
C7046 Vbias.n258 VGND 0.1294f
C7047 Vbias.t257 VGND 0.17892f
C7048 Vbias.n259 VGND 0.19512f
C7049 Vbias.n260 VGND 0.1294f
C7050 Vbias.t8 VGND 0.17892f
C7051 Vbias.n261 VGND 0.19512f
C7052 Vbias.n262 VGND 0.1294f
C7053 Vbias.t93 VGND 0.17892f
C7054 Vbias.n263 VGND 0.19512f
C7055 Vbias.n264 VGND 0.1294f
C7056 Vbias.t179 VGND 0.17892f
C7057 Vbias.n265 VGND 0.19512f
C7058 Vbias.n266 VGND 0.1294f
C7059 Vbias.t11 VGND 0.17892f
C7060 Vbias.n267 VGND 0.19512f
C7061 Vbias.n268 VGND 0.1294f
C7062 Vbias.t98 VGND 0.17892f
C7063 Vbias.n269 VGND 0.19512f
C7064 Vbias.n270 VGND 0.1294f
C7065 Vbias.t118 VGND 0.17892f
C7066 Vbias.n271 VGND 0.19512f
C7067 Vbias.n272 VGND 0.1294f
C7068 Vbias.t190 VGND 0.17892f
C7069 Vbias.n273 VGND 0.19512f
C7070 Vbias.n274 VGND 0.1294f
C7071 Vbias.t27 VGND 0.17892f
C7072 Vbias.n275 VGND 0.19512f
C7073 Vbias.n276 VGND 0.1294f
C7074 Vbias.t44 VGND 0.17892f
C7075 Vbias.n277 VGND 0.19512f
C7076 Vbias.n278 VGND 0.1294f
C7077 Vbias.t197 VGND 0.17892f
C7078 Vbias.n279 VGND 0.19512f
C7079 Vbias.n280 VGND 0.1294f
C7080 Vbias.t220 VGND 0.17892f
C7081 Vbias.n281 VGND 0.19512f
C7082 Vbias.n282 VGND 0.1294f
C7083 Vbias.t232 VGND 0.17892f
C7084 Vbias.n283 VGND 0.19512f
C7085 Vbias.n284 VGND 0.1294f
C7086 Vbias.t137 VGND 0.17892f
C7087 Vbias.n285 VGND 0.19512f
C7088 Vbias.n286 VGND 0.1294f
C7089 Vbias.n287 VGND 0.55864f
C7090 Vbias.t49 VGND 0.17892f
C7091 Vbias.n288 VGND 0.19478f
C7092 Vbias.t122 VGND 0.17892f
C7093 Vbias.n289 VGND 0.19512f
C7094 Vbias.n290 VGND 0.1294f
C7095 Vbias.t222 VGND 0.17892f
C7096 Vbias.n291 VGND 0.19512f
C7097 Vbias.n292 VGND 0.1294f
C7098 Vbias.t235 VGND 0.17892f
C7099 Vbias.n293 VGND 0.19512f
C7100 Vbias.n294 VGND 0.1294f
C7101 Vbias.t63 VGND 0.17892f
C7102 Vbias.n295 VGND 0.19512f
C7103 Vbias.n296 VGND 0.1294f
C7104 Vbias.t150 VGND 0.17892f
C7105 Vbias.n297 VGND 0.19512f
C7106 Vbias.n298 VGND 0.1294f
C7107 Vbias.t237 VGND 0.17892f
C7108 Vbias.n299 VGND 0.19512f
C7109 Vbias.n300 VGND 0.1294f
C7110 Vbias.t68 VGND 0.17892f
C7111 Vbias.n301 VGND 0.19512f
C7112 Vbias.n302 VGND 0.1294f
C7113 Vbias.t91 VGND 0.17892f
C7114 Vbias.n303 VGND 0.19512f
C7115 Vbias.n304 VGND 0.1294f
C7116 Vbias.t164 VGND 0.17892f
C7117 Vbias.n305 VGND 0.19512f
C7118 Vbias.n306 VGND 0.1294f
C7119 Vbias.t251 VGND 0.17892f
C7120 Vbias.n307 VGND 0.19512f
C7121 Vbias.n308 VGND 0.1294f
C7122 Vbias.t21 VGND 0.17892f
C7123 Vbias.n309 VGND 0.19512f
C7124 Vbias.n310 VGND 0.1294f
C7125 Vbias.t168 VGND 0.17892f
C7126 Vbias.n311 VGND 0.19512f
C7127 Vbias.n312 VGND 0.1294f
C7128 Vbias.t187 VGND 0.17892f
C7129 Vbias.n313 VGND 0.19512f
C7130 Vbias.n314 VGND 0.1294f
C7131 Vbias.t204 VGND 0.17892f
C7132 Vbias.n315 VGND 0.19512f
C7133 Vbias.n316 VGND 0.1294f
C7134 Vbias.t105 VGND 0.17892f
C7135 Vbias.n317 VGND 0.19512f
C7136 Vbias.n318 VGND 0.1294f
C7137 Vbias.n319 VGND 0.55864f
C7138 Vbias.t121 VGND 0.17892f
C7139 Vbias.n320 VGND 0.19478f
C7140 Vbias.t195 VGND 0.17892f
C7141 Vbias.n321 VGND 0.19512f
C7142 Vbias.n322 VGND 0.1294f
C7143 Vbias.t37 VGND 0.17892f
C7144 Vbias.n323 VGND 0.19512f
C7145 Vbias.n324 VGND 0.1294f
C7146 Vbias.t48 VGND 0.17892f
C7147 Vbias.n325 VGND 0.19512f
C7148 Vbias.n326 VGND 0.1294f
C7149 Vbias.t135 VGND 0.17892f
C7150 Vbias.n327 VGND 0.19512f
C7151 Vbias.n328 VGND 0.1294f
C7152 Vbias.t221 VGND 0.17892f
C7153 Vbias.n329 VGND 0.19512f
C7154 Vbias.n330 VGND 0.1294f
C7155 Vbias.t50 VGND 0.17892f
C7156 Vbias.n331 VGND 0.19512f
C7157 Vbias.n332 VGND 0.1294f
C7158 Vbias.t138 VGND 0.17892f
C7159 Vbias.n333 VGND 0.19512f
C7160 Vbias.n334 VGND 0.1294f
C7161 Vbias.t163 VGND 0.17892f
C7162 Vbias.n335 VGND 0.19512f
C7163 Vbias.n336 VGND 0.1294f
C7164 Vbias.t236 VGND 0.17892f
C7165 Vbias.n337 VGND 0.19512f
C7166 Vbias.n338 VGND 0.1294f
C7167 Vbias.t65 VGND 0.17892f
C7168 Vbias.n339 VGND 0.19512f
C7169 Vbias.n340 VGND 0.1294f
C7170 Vbias.t90 VGND 0.17892f
C7171 Vbias.n341 VGND 0.19512f
C7172 Vbias.n342 VGND 0.1294f
C7173 Vbias.t243 VGND 0.17892f
C7174 Vbias.n343 VGND 0.19512f
C7175 Vbias.n344 VGND 0.1294f
C7176 Vbias.t7 VGND 0.17892f
C7177 Vbias.n345 VGND 0.19512f
C7178 Vbias.n346 VGND 0.1294f
C7179 Vbias.t20 VGND 0.17892f
C7180 Vbias.n347 VGND 0.19512f
C7181 Vbias.n348 VGND 0.1294f
C7182 Vbias.t176 VGND 0.17892f
C7183 Vbias.n349 VGND 0.19512f
C7184 Vbias.n350 VGND 0.1294f
C7185 Vbias.n351 VGND 0.55864f
C7186 Vbias.t198 VGND 0.17892f
C7187 Vbias.n352 VGND 0.19478f
C7188 Vbias.t17 VGND 0.17892f
C7189 Vbias.n353 VGND 0.19512f
C7190 Vbias.n354 VGND 0.1294f
C7191 Vbias.t113 VGND 0.17892f
C7192 Vbias.n355 VGND 0.19512f
C7193 Vbias.n356 VGND 0.1294f
C7194 Vbias.t124 VGND 0.17892f
C7195 Vbias.n357 VGND 0.19512f
C7196 Vbias.n358 VGND 0.1294f
C7197 Vbias.t213 VGND 0.17892f
C7198 Vbias.n359 VGND 0.19512f
C7199 Vbias.n360 VGND 0.1294f
C7200 Vbias.t40 VGND 0.17892f
C7201 Vbias.n361 VGND 0.19512f
C7202 Vbias.n362 VGND 0.1294f
C7203 Vbias.t127 VGND 0.17892f
C7204 Vbias.n363 VGND 0.19512f
C7205 Vbias.n364 VGND 0.1294f
C7206 Vbias.t219 VGND 0.17892f
C7207 Vbias.n365 VGND 0.19512f
C7208 Vbias.n366 VGND 0.1294f
C7209 Vbias.t240 VGND 0.17892f
C7210 Vbias.n367 VGND 0.19512f
C7211 Vbias.n368 VGND 0.1294f
C7212 Vbias.t54 VGND 0.17892f
C7213 Vbias.n369 VGND 0.19512f
C7214 Vbias.n370 VGND 0.1294f
C7215 Vbias.t144 VGND 0.17892f
C7216 Vbias.n371 VGND 0.19512f
C7217 Vbias.n372 VGND 0.1294f
C7218 Vbias.t166 VGND 0.17892f
C7219 Vbias.n373 VGND 0.19512f
C7220 Vbias.n374 VGND 0.1294f
C7221 Vbias.t62 VGND 0.17892f
C7222 Vbias.n375 VGND 0.19512f
C7223 Vbias.n376 VGND 0.1294f
C7224 Vbias.t81 VGND 0.17892f
C7225 Vbias.n377 VGND 0.19512f
C7226 Vbias.n378 VGND 0.1294f
C7227 Vbias.t92 VGND 0.17892f
C7228 Vbias.n379 VGND 0.19512f
C7229 Vbias.n380 VGND 0.1294f
C7230 Vbias.t255 VGND 0.17892f
C7231 Vbias.n381 VGND 0.19512f
C7232 Vbias.n382 VGND 0.1294f
C7233 Vbias.n383 VGND 0.55864f
C7234 Vbias.t16 VGND 0.17892f
C7235 Vbias.n384 VGND 0.19478f
C7236 Vbias.t88 VGND 0.17892f
C7237 Vbias.n385 VGND 0.19512f
C7238 Vbias.n386 VGND 0.1294f
C7239 Vbias.t185 VGND 0.17892f
C7240 Vbias.n387 VGND 0.19512f
C7241 Vbias.n388 VGND 0.1294f
C7242 Vbias.t196 VGND 0.17892f
C7243 Vbias.n389 VGND 0.19512f
C7244 Vbias.n390 VGND 0.1294f
C7245 Vbias.t29 VGND 0.17892f
C7246 Vbias.n391 VGND 0.19512f
C7247 Vbias.n392 VGND 0.1294f
C7248 Vbias.t112 VGND 0.17892f
C7249 Vbias.n393 VGND 0.19512f
C7250 Vbias.n394 VGND 0.1294f
C7251 Vbias.t200 VGND 0.17892f
C7252 Vbias.n395 VGND 0.19512f
C7253 Vbias.n396 VGND 0.1294f
C7254 Vbias.t33 VGND 0.17892f
C7255 Vbias.n397 VGND 0.19512f
C7256 Vbias.n398 VGND 0.1294f
C7257 Vbias.t53 VGND 0.17892f
C7258 Vbias.n399 VGND 0.19512f
C7259 Vbias.n400 VGND 0.1294f
C7260 Vbias.t126 VGND 0.17892f
C7261 Vbias.n401 VGND 0.19512f
C7262 Vbias.n402 VGND 0.1294f
C7263 Vbias.t217 VGND 0.17892f
C7264 Vbias.n403 VGND 0.19512f
C7265 Vbias.n404 VGND 0.1294f
C7266 Vbias.t239 VGND 0.17892f
C7267 Vbias.n405 VGND 0.19512f
C7268 Vbias.n406 VGND 0.1294f
C7269 Vbias.t133 VGND 0.17892f
C7270 Vbias.n407 VGND 0.19512f
C7271 Vbias.n408 VGND 0.1294f
C7272 Vbias.t153 VGND 0.17892f
C7273 Vbias.n409 VGND 0.19512f
C7274 Vbias.n410 VGND 0.1294f
C7275 Vbias.t165 VGND 0.17892f
C7276 Vbias.n411 VGND 0.19512f
C7277 Vbias.n412 VGND 0.1294f
C7278 Vbias.t73 VGND 0.17892f
C7279 Vbias.n413 VGND 0.19512f
C7280 Vbias.n414 VGND 0.1294f
C7281 Vbias.n415 VGND 0.55864f
C7282 Vbias.t87 VGND 0.17892f
C7283 Vbias.n416 VGND 0.19478f
C7284 Vbias.t160 VGND 0.17892f
C7285 Vbias.n417 VGND 0.19512f
C7286 Vbias.n418 VGND 0.1294f
C7287 Vbias.t261 VGND 0.17892f
C7288 Vbias.n419 VGND 0.19512f
C7289 Vbias.n420 VGND 0.1294f
C7290 Vbias.t14 VGND 0.17892f
C7291 Vbias.n421 VGND 0.19512f
C7292 Vbias.n422 VGND 0.1294f
C7293 Vbias.t99 VGND 0.17892f
C7294 Vbias.n423 VGND 0.19512f
C7295 Vbias.n424 VGND 0.1294f
C7296 Vbias.t183 VGND 0.17892f
C7297 Vbias.n425 VGND 0.19512f
C7298 Vbias.n426 VGND 0.1294f
C7299 Vbias.t18 VGND 0.17892f
C7300 Vbias.n427 VGND 0.19512f
C7301 Vbias.n428 VGND 0.1294f
C7302 Vbias.t102 VGND 0.17892f
C7303 Vbias.n429 VGND 0.19512f
C7304 Vbias.n430 VGND 0.1294f
C7305 Vbias.t125 VGND 0.17892f
C7306 Vbias.n431 VGND 0.19512f
C7307 Vbias.n432 VGND 0.1294f
C7308 Vbias.t199 VGND 0.17892f
C7309 Vbias.n433 VGND 0.19512f
C7310 Vbias.n434 VGND 0.1294f
C7311 Vbias.t32 VGND 0.17892f
C7312 Vbias.n435 VGND 0.19512f
C7313 Vbias.n436 VGND 0.1294f
C7314 Vbias.t52 VGND 0.17892f
C7315 Vbias.n437 VGND 0.19512f
C7316 Vbias.n438 VGND 0.1294f
C7317 Vbias.t205 VGND 0.17892f
C7318 Vbias.n439 VGND 0.19512f
C7319 Vbias.n440 VGND 0.1294f
C7320 Vbias.t225 VGND 0.17892f
C7321 Vbias.n441 VGND 0.19512f
C7322 Vbias.n442 VGND 0.1294f
C7323 Vbias.t238 VGND 0.17892f
C7324 Vbias.n443 VGND 0.19512f
C7325 Vbias.n444 VGND 0.1294f
C7326 Vbias.t146 VGND 0.17892f
C7327 Vbias.n445 VGND 0.19512f
C7328 Vbias.n446 VGND 0.1294f
C7329 Vbias.n447 VGND 0.55864f
C7330 Vbias.t57 VGND 0.17892f
C7331 Vbias.n448 VGND 0.19478f
C7332 Vbias.t130 VGND 0.17892f
C7333 Vbias.n449 VGND 0.19512f
C7334 Vbias.n450 VGND 0.1294f
C7335 Vbias.t229 VGND 0.17892f
C7336 Vbias.n451 VGND 0.19512f
C7337 Vbias.n452 VGND 0.1294f
C7338 Vbias.t242 VGND 0.17892f
C7339 Vbias.n453 VGND 0.19512f
C7340 Vbias.n454 VGND 0.1294f
C7341 Vbias.t69 VGND 0.17892f
C7342 Vbias.n455 VGND 0.19512f
C7343 Vbias.n456 VGND 0.1294f
C7344 Vbias.t156 VGND 0.17892f
C7345 Vbias.n457 VGND 0.19512f
C7346 Vbias.n458 VGND 0.1294f
C7347 Vbias.t247 VGND 0.17892f
C7348 Vbias.n459 VGND 0.19512f
C7349 Vbias.n460 VGND 0.1294f
C7350 Vbias.t76 VGND 0.17892f
C7351 Vbias.n461 VGND 0.19512f
C7352 Vbias.n462 VGND 0.1294f
C7353 Vbias.t96 VGND 0.17892f
C7354 Vbias.n463 VGND 0.19512f
C7355 Vbias.n464 VGND 0.1294f
C7356 Vbias.t171 VGND 0.17892f
C7357 Vbias.n465 VGND 0.19512f
C7358 Vbias.n466 VGND 0.1294f
C7359 Vbias.t258 VGND 0.17892f
C7360 Vbias.n467 VGND 0.19512f
C7361 Vbias.n468 VGND 0.1294f
C7362 Vbias.t25 VGND 0.17892f
C7363 Vbias.n469 VGND 0.19512f
C7364 Vbias.n470 VGND 0.1294f
C7365 Vbias.t173 VGND 0.17892f
C7366 Vbias.n471 VGND 0.19512f
C7367 Vbias.n472 VGND 0.1294f
C7368 Vbias.t193 VGND 0.17892f
C7369 Vbias.n473 VGND 0.19512f
C7370 Vbias.n474 VGND 0.1294f
C7371 Vbias.t210 VGND 0.17892f
C7372 Vbias.n475 VGND 0.19512f
C7373 Vbias.n476 VGND 0.1294f
C7374 Vbias.t110 VGND 0.17892f
C7375 Vbias.n477 VGND 0.19512f
C7376 Vbias.n478 VGND 0.1294f
C7377 Vbias.n479 VGND 0.55864f
C7378 Vbias.t129 VGND 0.17892f
C7379 Vbias.n480 VGND 0.19478f
C7380 Vbias.t201 VGND 0.17892f
C7381 Vbias.n481 VGND 0.19512f
C7382 Vbias.n482 VGND 0.1294f
C7383 Vbias.t41 VGND 0.17892f
C7384 Vbias.n483 VGND 0.19512f
C7385 Vbias.n484 VGND 0.1294f
C7386 Vbias.t56 VGND 0.17892f
C7387 Vbias.n485 VGND 0.19512f
C7388 Vbias.n486 VGND 0.1294f
C7389 Vbias.t141 VGND 0.17892f
C7390 Vbias.n487 VGND 0.19512f
C7391 Vbias.n488 VGND 0.1294f
C7392 Vbias.t227 VGND 0.17892f
C7393 Vbias.n489 VGND 0.19512f
C7394 Vbias.n490 VGND 0.1294f
C7395 Vbias.t60 VGND 0.17892f
C7396 Vbias.n491 VGND 0.19512f
C7397 Vbias.n492 VGND 0.1294f
C7398 Vbias.t147 VGND 0.17892f
C7399 Vbias.n493 VGND 0.19512f
C7400 Vbias.n494 VGND 0.1294f
C7401 Vbias.t169 VGND 0.17892f
C7402 Vbias.n495 VGND 0.19512f
C7403 Vbias.n496 VGND 0.1294f
C7404 Vbias.t246 VGND 0.17892f
C7405 Vbias.n497 VGND 0.19512f
C7406 Vbias.n498 VGND 0.1294f
C7407 Vbias.t75 VGND 0.17892f
C7408 Vbias.n499 VGND 0.19512f
C7409 Vbias.n500 VGND 0.1294f
C7410 Vbias.t95 VGND 0.17892f
C7411 Vbias.n501 VGND 0.19512f
C7412 Vbias.n502 VGND 0.1294f
C7413 Vbias.t248 VGND 0.17892f
C7414 Vbias.n503 VGND 0.19512f
C7415 Vbias.n504 VGND 0.1294f
C7416 Vbias.t12 VGND 0.17892f
C7417 Vbias.n505 VGND 0.19512f
C7418 Vbias.n506 VGND 0.1294f
C7419 Vbias.t24 VGND 0.17892f
C7420 Vbias.n507 VGND 0.19512f
C7421 Vbias.n508 VGND 0.1294f
C7422 Vbias.t181 VGND 0.17892f
C7423 Vbias.n509 VGND 0.19512f
C7424 Vbias.n510 VGND 0.1294f
C7425 Vbias.n511 VGND 0.64971f
C7426 Vbias.t2 VGND 0.03656f
C7427 Vbias.t5 VGND 0.03656f
C7428 Vbias.n512 VGND 0.24632f
C7429 Vbias.t4 VGND 0.03656f
C7430 Vbias.t3 VGND 0.03656f
C7431 Vbias.n513 VGND 0.24632f
C7432 Vbias.n514 VGND 0.74347f
C7433 Vbias.t1 VGND 0.17053f
C7434 Vbias.t0 VGND 0.67054f
C7435 Vbias.n515 VGND 1.24142f
C7436 Vbias.n516 VGND 0.47748f
C7437 Vbias.n517 VGND 1.11804f
C7438 XThC.Tn[2].t5 VGND 0.01376f
C7439 XThC.Tn[2].t4 VGND 0.01376f
C7440 XThC.Tn[2].n0 VGND 0.02778f
C7441 XThC.Tn[2].t3 VGND 0.01376f
C7442 XThC.Tn[2].t2 VGND 0.01376f
C7443 XThC.Tn[2].n1 VGND 0.03251f
C7444 XThC.Tn[2].n2 VGND 0.091f
C7445 XThC.Tn[2].n3 VGND 0.02037f
C7446 XThC.Tn[2].n4 VGND 0.02037f
C7447 XThC.Tn[2].n5 VGND 0.02037f
C7448 XThC.Tn[2].n6 VGND 0.03395f
C7449 XThC.Tn[2].n7 VGND 0.09702f
C7450 XThC.Tn[2].n8 VGND 0.05998f
C7451 XThC.Tn[2].n9 VGND 0.06769f
C7452 XThC.Tn[2].t20 VGND 0.01091f
C7453 XThC.Tn[2].t18 VGND 0.01192f
C7454 XThC.Tn[2].n10 VGND 0.0266f
C7455 XThC.Tn[2].n11 VGND 0.01822f
C7456 XThC.Tn[2].n12 VGND 0.05982f
C7457 XThC.Tn[2].t38 VGND 0.01091f
C7458 XThC.Tn[2].t35 VGND 0.01192f
C7459 XThC.Tn[2].n13 VGND 0.0266f
C7460 XThC.Tn[2].n14 VGND 0.01822f
C7461 XThC.Tn[2].n15 VGND 0.05998f
C7462 XThC.Tn[2].n16 VGND 0.09886f
C7463 XThC.Tn[2].t43 VGND 0.01091f
C7464 XThC.Tn[2].t37 VGND 0.01192f
C7465 XThC.Tn[2].n17 VGND 0.0266f
C7466 XThC.Tn[2].n18 VGND 0.01822f
C7467 XThC.Tn[2].n19 VGND 0.05998f
C7468 XThC.Tn[2].n20 VGND 0.09886f
C7469 XThC.Tn[2].t12 VGND 0.01091f
C7470 XThC.Tn[2].t39 VGND 0.01192f
C7471 XThC.Tn[2].n21 VGND 0.0266f
C7472 XThC.Tn[2].n22 VGND 0.01822f
C7473 XThC.Tn[2].n23 VGND 0.05998f
C7474 XThC.Tn[2].n24 VGND 0.09886f
C7475 XThC.Tn[2].t31 VGND 0.01091f
C7476 XThC.Tn[2].t28 VGND 0.01192f
C7477 XThC.Tn[2].n25 VGND 0.0266f
C7478 XThC.Tn[2].n26 VGND 0.01822f
C7479 XThC.Tn[2].n27 VGND 0.05998f
C7480 XThC.Tn[2].n28 VGND 0.09886f
C7481 XThC.Tn[2].t32 VGND 0.01091f
C7482 XThC.Tn[2].t29 VGND 0.01192f
C7483 XThC.Tn[2].n29 VGND 0.0266f
C7484 XThC.Tn[2].n30 VGND 0.01822f
C7485 XThC.Tn[2].n31 VGND 0.05998f
C7486 XThC.Tn[2].n32 VGND 0.09886f
C7487 XThC.Tn[2].t16 VGND 0.01091f
C7488 XThC.Tn[2].t42 VGND 0.01192f
C7489 XThC.Tn[2].n33 VGND 0.0266f
C7490 XThC.Tn[2].n34 VGND 0.01822f
C7491 XThC.Tn[2].n35 VGND 0.05998f
C7492 XThC.Tn[2].n36 VGND 0.09886f
C7493 XThC.Tn[2].t23 VGND 0.01091f
C7494 XThC.Tn[2].t19 VGND 0.01192f
C7495 XThC.Tn[2].n37 VGND 0.0266f
C7496 XThC.Tn[2].n38 VGND 0.01822f
C7497 XThC.Tn[2].n39 VGND 0.05998f
C7498 XThC.Tn[2].n40 VGND 0.09886f
C7499 XThC.Tn[2].t25 VGND 0.01091f
C7500 XThC.Tn[2].t21 VGND 0.01192f
C7501 XThC.Tn[2].n41 VGND 0.0266f
C7502 XThC.Tn[2].n42 VGND 0.01822f
C7503 XThC.Tn[2].n43 VGND 0.05998f
C7504 XThC.Tn[2].n44 VGND 0.09886f
C7505 XThC.Tn[2].t13 VGND 0.01091f
C7506 XThC.Tn[2].t40 VGND 0.01192f
C7507 XThC.Tn[2].n45 VGND 0.0266f
C7508 XThC.Tn[2].n46 VGND 0.01822f
C7509 XThC.Tn[2].n47 VGND 0.05998f
C7510 XThC.Tn[2].n48 VGND 0.09886f
C7511 XThC.Tn[2].t15 VGND 0.01091f
C7512 XThC.Tn[2].t41 VGND 0.01192f
C7513 XThC.Tn[2].n49 VGND 0.0266f
C7514 XThC.Tn[2].n50 VGND 0.01822f
C7515 XThC.Tn[2].n51 VGND 0.05998f
C7516 XThC.Tn[2].n52 VGND 0.09886f
C7517 XThC.Tn[2].t26 VGND 0.01091f
C7518 XThC.Tn[2].t22 VGND 0.01192f
C7519 XThC.Tn[2].n53 VGND 0.0266f
C7520 XThC.Tn[2].n54 VGND 0.01822f
C7521 XThC.Tn[2].n55 VGND 0.05998f
C7522 XThC.Tn[2].n56 VGND 0.09886f
C7523 XThC.Tn[2].t34 VGND 0.01091f
C7524 XThC.Tn[2].t30 VGND 0.01192f
C7525 XThC.Tn[2].n57 VGND 0.0266f
C7526 XThC.Tn[2].n58 VGND 0.01822f
C7527 XThC.Tn[2].n59 VGND 0.05998f
C7528 XThC.Tn[2].n60 VGND 0.09886f
C7529 XThC.Tn[2].t36 VGND 0.01091f
C7530 XThC.Tn[2].t33 VGND 0.01192f
C7531 XThC.Tn[2].n61 VGND 0.0266f
C7532 XThC.Tn[2].n62 VGND 0.01822f
C7533 XThC.Tn[2].n63 VGND 0.05998f
C7534 XThC.Tn[2].n64 VGND 0.09886f
C7535 XThC.Tn[2].t17 VGND 0.01091f
C7536 XThC.Tn[2].t14 VGND 0.01192f
C7537 XThC.Tn[2].n65 VGND 0.0266f
C7538 XThC.Tn[2].n66 VGND 0.01822f
C7539 XThC.Tn[2].n67 VGND 0.05998f
C7540 XThC.Tn[2].n68 VGND 0.09886f
C7541 XThC.Tn[2].t27 VGND 0.01091f
C7542 XThC.Tn[2].t24 VGND 0.01192f
C7543 XThC.Tn[2].n69 VGND 0.0266f
C7544 XThC.Tn[2].n70 VGND 0.01822f
C7545 XThC.Tn[2].n71 VGND 0.05998f
C7546 XThC.Tn[2].n72 VGND 0.09886f
C7547 XThC.Tn[2].n73 VGND 0.38259f
C7548 XThC.Tn[2].n74 VGND 0.08113f
C7549 XThC.Tn[2].n75 VGND 0.0288f
C7550 XThC.Tn[4].t5 VGND 0.01387f
C7551 XThC.Tn[4].t4 VGND 0.01387f
C7552 XThC.Tn[4].n0 VGND 0.028f
C7553 XThC.Tn[4].t7 VGND 0.01387f
C7554 XThC.Tn[4].t6 VGND 0.01387f
C7555 XThC.Tn[4].n1 VGND 0.03276f
C7556 XThC.Tn[4].n2 VGND 0.09172f
C7557 XThC.Tn[4].n3 VGND 0.02053f
C7558 XThC.Tn[4].n4 VGND 0.02053f
C7559 XThC.Tn[4].n5 VGND 0.02053f
C7560 XThC.Tn[4].n6 VGND 0.03421f
C7561 XThC.Tn[4].n7 VGND 0.09778f
C7562 XThC.Tn[4].n8 VGND 0.06045f
C7563 XThC.Tn[4].n9 VGND 0.06822f
C7564 XThC.Tn[4].t28 VGND 0.01099f
C7565 XThC.Tn[4].t26 VGND 0.01201f
C7566 XThC.Tn[4].n10 VGND 0.02681f
C7567 XThC.Tn[4].n11 VGND 0.01837f
C7568 XThC.Tn[4].n12 VGND 0.06029f
C7569 XThC.Tn[4].t14 VGND 0.01099f
C7570 XThC.Tn[4].t43 VGND 0.01201f
C7571 XThC.Tn[4].n13 VGND 0.02681f
C7572 XThC.Tn[4].n14 VGND 0.01837f
C7573 XThC.Tn[4].n15 VGND 0.06045f
C7574 XThC.Tn[4].n16 VGND 0.09963f
C7575 XThC.Tn[4].t19 VGND 0.01099f
C7576 XThC.Tn[4].t13 VGND 0.01201f
C7577 XThC.Tn[4].n17 VGND 0.02681f
C7578 XThC.Tn[4].n18 VGND 0.01837f
C7579 XThC.Tn[4].n19 VGND 0.06045f
C7580 XThC.Tn[4].n20 VGND 0.09963f
C7581 XThC.Tn[4].t20 VGND 0.01099f
C7582 XThC.Tn[4].t15 VGND 0.01201f
C7583 XThC.Tn[4].n21 VGND 0.02681f
C7584 XThC.Tn[4].n22 VGND 0.01837f
C7585 XThC.Tn[4].n23 VGND 0.06045f
C7586 XThC.Tn[4].n24 VGND 0.09963f
C7587 XThC.Tn[4].t39 VGND 0.01099f
C7588 XThC.Tn[4].t36 VGND 0.01201f
C7589 XThC.Tn[4].n25 VGND 0.02681f
C7590 XThC.Tn[4].n26 VGND 0.01837f
C7591 XThC.Tn[4].n27 VGND 0.06045f
C7592 XThC.Tn[4].n28 VGND 0.09963f
C7593 XThC.Tn[4].t40 VGND 0.01099f
C7594 XThC.Tn[4].t37 VGND 0.01201f
C7595 XThC.Tn[4].n29 VGND 0.02681f
C7596 XThC.Tn[4].n30 VGND 0.01837f
C7597 XThC.Tn[4].n31 VGND 0.06045f
C7598 XThC.Tn[4].n32 VGND 0.09963f
C7599 XThC.Tn[4].t24 VGND 0.01099f
C7600 XThC.Tn[4].t18 VGND 0.01201f
C7601 XThC.Tn[4].n33 VGND 0.02681f
C7602 XThC.Tn[4].n34 VGND 0.01837f
C7603 XThC.Tn[4].n35 VGND 0.06045f
C7604 XThC.Tn[4].n36 VGND 0.09963f
C7605 XThC.Tn[4].t31 VGND 0.01099f
C7606 XThC.Tn[4].t27 VGND 0.01201f
C7607 XThC.Tn[4].n37 VGND 0.02681f
C7608 XThC.Tn[4].n38 VGND 0.01837f
C7609 XThC.Tn[4].n39 VGND 0.06045f
C7610 XThC.Tn[4].n40 VGND 0.09963f
C7611 XThC.Tn[4].t33 VGND 0.01099f
C7612 XThC.Tn[4].t29 VGND 0.01201f
C7613 XThC.Tn[4].n41 VGND 0.02681f
C7614 XThC.Tn[4].n42 VGND 0.01837f
C7615 XThC.Tn[4].n43 VGND 0.06045f
C7616 XThC.Tn[4].n44 VGND 0.09963f
C7617 XThC.Tn[4].t21 VGND 0.01099f
C7618 XThC.Tn[4].t16 VGND 0.01201f
C7619 XThC.Tn[4].n45 VGND 0.02681f
C7620 XThC.Tn[4].n46 VGND 0.01837f
C7621 XThC.Tn[4].n47 VGND 0.06045f
C7622 XThC.Tn[4].n48 VGND 0.09963f
C7623 XThC.Tn[4].t23 VGND 0.01099f
C7624 XThC.Tn[4].t17 VGND 0.01201f
C7625 XThC.Tn[4].n49 VGND 0.02681f
C7626 XThC.Tn[4].n50 VGND 0.01837f
C7627 XThC.Tn[4].n51 VGND 0.06045f
C7628 XThC.Tn[4].n52 VGND 0.09963f
C7629 XThC.Tn[4].t34 VGND 0.01099f
C7630 XThC.Tn[4].t30 VGND 0.01201f
C7631 XThC.Tn[4].n53 VGND 0.02681f
C7632 XThC.Tn[4].n54 VGND 0.01837f
C7633 XThC.Tn[4].n55 VGND 0.06045f
C7634 XThC.Tn[4].n56 VGND 0.09963f
C7635 XThC.Tn[4].t42 VGND 0.01099f
C7636 XThC.Tn[4].t38 VGND 0.01201f
C7637 XThC.Tn[4].n57 VGND 0.02681f
C7638 XThC.Tn[4].n58 VGND 0.01837f
C7639 XThC.Tn[4].n59 VGND 0.06045f
C7640 XThC.Tn[4].n60 VGND 0.09963f
C7641 XThC.Tn[4].t12 VGND 0.01099f
C7642 XThC.Tn[4].t41 VGND 0.01201f
C7643 XThC.Tn[4].n61 VGND 0.02681f
C7644 XThC.Tn[4].n62 VGND 0.01837f
C7645 XThC.Tn[4].n63 VGND 0.06045f
C7646 XThC.Tn[4].n64 VGND 0.09963f
C7647 XThC.Tn[4].t25 VGND 0.01099f
C7648 XThC.Tn[4].t22 VGND 0.01201f
C7649 XThC.Tn[4].n65 VGND 0.02681f
C7650 XThC.Tn[4].n66 VGND 0.01837f
C7651 XThC.Tn[4].n67 VGND 0.06045f
C7652 XThC.Tn[4].n68 VGND 0.09963f
C7653 XThC.Tn[4].t35 VGND 0.01099f
C7654 XThC.Tn[4].t32 VGND 0.01201f
C7655 XThC.Tn[4].n69 VGND 0.02681f
C7656 XThC.Tn[4].n70 VGND 0.01837f
C7657 XThC.Tn[4].n71 VGND 0.06045f
C7658 XThC.Tn[4].n72 VGND 0.09963f
C7659 XThC.Tn[4].n73 VGND 0.12212f
C7660 XThC.Tn[4].n74 VGND 0.02903f
C7661 XThR.Tn[5].t10 VGND 0.01876f
C7662 XThR.Tn[5].t11 VGND 0.01876f
C7663 XThR.Tn[5].n0 VGND 0.03786f
C7664 XThR.Tn[5].t9 VGND 0.01876f
C7665 XThR.Tn[5].t8 VGND 0.01876f
C7666 XThR.Tn[5].n1 VGND 0.0443f
C7667 XThR.Tn[5].n2 VGND 0.124f
C7668 XThR.Tn[5].t7 VGND 0.01219f
C7669 XThR.Tn[5].t4 VGND 0.01219f
C7670 XThR.Tn[5].n3 VGND 0.02776f
C7671 XThR.Tn[5].t6 VGND 0.01219f
C7672 XThR.Tn[5].t5 VGND 0.01219f
C7673 XThR.Tn[5].n4 VGND 0.02776f
C7674 XThR.Tn[5].t0 VGND 0.01219f
C7675 XThR.Tn[5].t1 VGND 0.01219f
C7676 XThR.Tn[5].n5 VGND 0.04626f
C7677 XThR.Tn[5].t3 VGND 0.01219f
C7678 XThR.Tn[5].t2 VGND 0.01219f
C7679 XThR.Tn[5].n6 VGND 0.02776f
C7680 XThR.Tn[5].n7 VGND 0.13221f
C7681 XThR.Tn[5].n8 VGND 0.08173f
C7682 XThR.Tn[5].n9 VGND 0.09224f
C7683 XThR.Tn[5].t17 VGND 0.01466f
C7684 XThR.Tn[5].t72 VGND 0.01605f
C7685 XThR.Tn[5].n10 VGND 0.03919f
C7686 XThR.Tn[5].n11 VGND 0.07529f
C7687 XThR.Tn[5].t39 VGND 0.01466f
C7688 XThR.Tn[5].t26 VGND 0.01605f
C7689 XThR.Tn[5].n12 VGND 0.03919f
C7690 XThR.Tn[5].t13 VGND 0.01461f
C7691 XThR.Tn[5].t23 VGND 0.016f
C7692 XThR.Tn[5].n13 VGND 0.04078f
C7693 XThR.Tn[5].n14 VGND 0.02865f
C7694 XThR.Tn[5].n16 VGND 0.09194f
C7695 XThR.Tn[5].t73 VGND 0.01466f
C7696 XThR.Tn[5].t66 VGND 0.01605f
C7697 XThR.Tn[5].n17 VGND 0.03919f
C7698 XThR.Tn[5].t48 VGND 0.01461f
C7699 XThR.Tn[5].t61 VGND 0.016f
C7700 XThR.Tn[5].n18 VGND 0.04078f
C7701 XThR.Tn[5].n19 VGND 0.02865f
C7702 XThR.Tn[5].n21 VGND 0.09194f
C7703 XThR.Tn[5].t28 VGND 0.01466f
C7704 XThR.Tn[5].t21 VGND 0.01605f
C7705 XThR.Tn[5].n22 VGND 0.03919f
C7706 XThR.Tn[5].t65 VGND 0.01461f
C7707 XThR.Tn[5].t18 VGND 0.016f
C7708 XThR.Tn[5].n23 VGND 0.04078f
C7709 XThR.Tn[5].n24 VGND 0.02865f
C7710 XThR.Tn[5].n26 VGND 0.09194f
C7711 XThR.Tn[5].t55 VGND 0.01466f
C7712 XThR.Tn[5].t51 VGND 0.01605f
C7713 XThR.Tn[5].n27 VGND 0.03919f
C7714 XThR.Tn[5].t33 VGND 0.01461f
C7715 XThR.Tn[5].t46 VGND 0.016f
C7716 XThR.Tn[5].n28 VGND 0.04078f
C7717 XThR.Tn[5].n29 VGND 0.02865f
C7718 XThR.Tn[5].n31 VGND 0.09194f
C7719 XThR.Tn[5].t30 VGND 0.01466f
C7720 XThR.Tn[5].t22 VGND 0.01605f
C7721 XThR.Tn[5].n32 VGND 0.03919f
C7722 XThR.Tn[5].t67 VGND 0.01461f
C7723 XThR.Tn[5].t19 VGND 0.016f
C7724 XThR.Tn[5].n33 VGND 0.04078f
C7725 XThR.Tn[5].n34 VGND 0.02865f
C7726 XThR.Tn[5].n36 VGND 0.09194f
C7727 XThR.Tn[5].t69 VGND 0.01466f
C7728 XThR.Tn[5].t40 VGND 0.01605f
C7729 XThR.Tn[5].n37 VGND 0.03919f
C7730 XThR.Tn[5].t43 VGND 0.01461f
C7731 XThR.Tn[5].t37 VGND 0.016f
C7732 XThR.Tn[5].n38 VGND 0.04078f
C7733 XThR.Tn[5].n39 VGND 0.02865f
C7734 XThR.Tn[5].n41 VGND 0.09194f
C7735 XThR.Tn[5].t38 VGND 0.01466f
C7736 XThR.Tn[5].t32 VGND 0.01605f
C7737 XThR.Tn[5].n42 VGND 0.03919f
C7738 XThR.Tn[5].t14 VGND 0.01461f
C7739 XThR.Tn[5].t29 VGND 0.016f
C7740 XThR.Tn[5].n43 VGND 0.04078f
C7741 XThR.Tn[5].n44 VGND 0.02865f
C7742 XThR.Tn[5].n46 VGND 0.09194f
C7743 XThR.Tn[5].t42 VGND 0.01466f
C7744 XThR.Tn[5].t49 VGND 0.01605f
C7745 XThR.Tn[5].n47 VGND 0.03919f
C7746 XThR.Tn[5].t16 VGND 0.01461f
C7747 XThR.Tn[5].t45 VGND 0.016f
C7748 XThR.Tn[5].n48 VGND 0.04078f
C7749 XThR.Tn[5].n49 VGND 0.02865f
C7750 XThR.Tn[5].n51 VGND 0.09194f
C7751 XThR.Tn[5].t58 VGND 0.01466f
C7752 XThR.Tn[5].t68 VGND 0.01605f
C7753 XThR.Tn[5].n52 VGND 0.03919f
C7754 XThR.Tn[5].t36 VGND 0.01461f
C7755 XThR.Tn[5].t63 VGND 0.016f
C7756 XThR.Tn[5].n53 VGND 0.04078f
C7757 XThR.Tn[5].n54 VGND 0.02865f
C7758 XThR.Tn[5].n56 VGND 0.09194f
C7759 XThR.Tn[5].t53 VGND 0.01466f
C7760 XThR.Tn[5].t24 VGND 0.01605f
C7761 XThR.Tn[5].n57 VGND 0.03919f
C7762 XThR.Tn[5].t25 VGND 0.01461f
C7763 XThR.Tn[5].t20 VGND 0.016f
C7764 XThR.Tn[5].n58 VGND 0.04078f
C7765 XThR.Tn[5].n59 VGND 0.02865f
C7766 XThR.Tn[5].n61 VGND 0.09194f
C7767 XThR.Tn[5].t71 VGND 0.01466f
C7768 XThR.Tn[5].t60 VGND 0.01605f
C7769 XThR.Tn[5].n62 VGND 0.03919f
C7770 XThR.Tn[5].t44 VGND 0.01461f
C7771 XThR.Tn[5].t57 VGND 0.016f
C7772 XThR.Tn[5].n63 VGND 0.04078f
C7773 XThR.Tn[5].n64 VGND 0.02865f
C7774 XThR.Tn[5].n66 VGND 0.09194f
C7775 XThR.Tn[5].t41 VGND 0.01466f
C7776 XThR.Tn[5].t35 VGND 0.01605f
C7777 XThR.Tn[5].n67 VGND 0.03919f
C7778 XThR.Tn[5].t15 VGND 0.01461f
C7779 XThR.Tn[5].t31 VGND 0.016f
C7780 XThR.Tn[5].n68 VGND 0.04078f
C7781 XThR.Tn[5].n69 VGND 0.02865f
C7782 XThR.Tn[5].n71 VGND 0.09194f
C7783 XThR.Tn[5].t56 VGND 0.01466f
C7784 XThR.Tn[5].t52 VGND 0.01605f
C7785 XThR.Tn[5].n72 VGND 0.03919f
C7786 XThR.Tn[5].t34 VGND 0.01461f
C7787 XThR.Tn[5].t47 VGND 0.016f
C7788 XThR.Tn[5].n73 VGND 0.04078f
C7789 XThR.Tn[5].n74 VGND 0.02865f
C7790 XThR.Tn[5].n76 VGND 0.09194f
C7791 XThR.Tn[5].t12 VGND 0.01466f
C7792 XThR.Tn[5].t70 VGND 0.01605f
C7793 XThR.Tn[5].n77 VGND 0.03919f
C7794 XThR.Tn[5].t50 VGND 0.01461f
C7795 XThR.Tn[5].t64 VGND 0.016f
C7796 XThR.Tn[5].n78 VGND 0.04078f
C7797 XThR.Tn[5].n79 VGND 0.02865f
C7798 XThR.Tn[5].n81 VGND 0.09194f
C7799 XThR.Tn[5].t54 VGND 0.01466f
C7800 XThR.Tn[5].t62 VGND 0.01605f
C7801 XThR.Tn[5].n82 VGND 0.03919f
C7802 XThR.Tn[5].t27 VGND 0.01461f
C7803 XThR.Tn[5].t59 VGND 0.016f
C7804 XThR.Tn[5].n83 VGND 0.04078f
C7805 XThR.Tn[5].n84 VGND 0.02865f
C7806 XThR.Tn[5].n86 VGND 0.09194f
C7807 XThR.Tn[5].n87 VGND 0.08355f
C7808 XThR.Tn[5].n88 VGND 0.16182f
C7809 XThR.Tn[5].n89 VGND 0.03925f
C7810 XThR.Tn[3].t2 VGND 0.01866f
C7811 XThR.Tn[3].t3 VGND 0.01866f
C7812 XThR.Tn[3].n0 VGND 0.03766f
C7813 XThR.Tn[3].t1 VGND 0.01866f
C7814 XThR.Tn[3].t4 VGND 0.01866f
C7815 XThR.Tn[3].n1 VGND 0.04406f
C7816 XThR.Tn[3].n2 VGND 0.12334f
C7817 XThR.Tn[3].t8 VGND 0.01213f
C7818 XThR.Tn[3].t5 VGND 0.01213f
C7819 XThR.Tn[3].n3 VGND 0.02761f
C7820 XThR.Tn[3].t7 VGND 0.01213f
C7821 XThR.Tn[3].t6 VGND 0.01213f
C7822 XThR.Tn[3].n4 VGND 0.02761f
C7823 XThR.Tn[3].t9 VGND 0.01213f
C7824 XThR.Tn[3].t10 VGND 0.01213f
C7825 XThR.Tn[3].n5 VGND 0.02761f
C7826 XThR.Tn[3].t0 VGND 0.01213f
C7827 XThR.Tn[3].t11 VGND 0.01213f
C7828 XThR.Tn[3].n6 VGND 0.04601f
C7829 XThR.Tn[3].n7 VGND 0.1315f
C7830 XThR.Tn[3].n8 VGND 0.08129f
C7831 XThR.Tn[3].n9 VGND 0.09175f
C7832 XThR.Tn[3].t64 VGND 0.01458f
C7833 XThR.Tn[3].t57 VGND 0.01597f
C7834 XThR.Tn[3].n10 VGND 0.03899f
C7835 XThR.Tn[3].n11 VGND 0.07489f
C7836 XThR.Tn[3].t18 VGND 0.01458f
C7837 XThR.Tn[3].t70 VGND 0.01597f
C7838 XThR.Tn[3].n12 VGND 0.03899f
C7839 XThR.Tn[3].t24 VGND 0.01453f
C7840 XThR.Tn[3].t55 VGND 0.01591f
C7841 XThR.Tn[3].n13 VGND 0.04056f
C7842 XThR.Tn[3].n14 VGND 0.0285f
C7843 XThR.Tn[3].n16 VGND 0.09145f
C7844 XThR.Tn[3].t59 VGND 0.01458f
C7845 XThR.Tn[3].t49 VGND 0.01597f
C7846 XThR.Tn[3].n17 VGND 0.03899f
C7847 XThR.Tn[3].t62 VGND 0.01453f
C7848 XThR.Tn[3].t29 VGND 0.01591f
C7849 XThR.Tn[3].n18 VGND 0.04056f
C7850 XThR.Tn[3].n19 VGND 0.0285f
C7851 XThR.Tn[3].n21 VGND 0.09145f
C7852 XThR.Tn[3].t71 VGND 0.01458f
C7853 XThR.Tn[3].t67 VGND 0.01597f
C7854 XThR.Tn[3].n22 VGND 0.03899f
C7855 XThR.Tn[3].t12 VGND 0.01453f
C7856 XThR.Tn[3].t47 VGND 0.01591f
C7857 XThR.Tn[3].n23 VGND 0.04056f
C7858 XThR.Tn[3].n24 VGND 0.0285f
C7859 XThR.Tn[3].n26 VGND 0.09145f
C7860 XThR.Tn[3].t39 VGND 0.01458f
C7861 XThR.Tn[3].t33 VGND 0.01597f
C7862 XThR.Tn[3].n27 VGND 0.03899f
C7863 XThR.Tn[3].t42 VGND 0.01453f
C7864 XThR.Tn[3].t13 VGND 0.01591f
C7865 XThR.Tn[3].n28 VGND 0.04056f
C7866 XThR.Tn[3].n29 VGND 0.0285f
C7867 XThR.Tn[3].n31 VGND 0.09145f
C7868 XThR.Tn[3].t72 VGND 0.01458f
C7869 XThR.Tn[3].t68 VGND 0.01597f
C7870 XThR.Tn[3].n32 VGND 0.03899f
C7871 XThR.Tn[3].t16 VGND 0.01453f
C7872 XThR.Tn[3].t48 VGND 0.01591f
C7873 XThR.Tn[3].n33 VGND 0.04056f
C7874 XThR.Tn[3].n34 VGND 0.0285f
C7875 XThR.Tn[3].n36 VGND 0.09145f
C7876 XThR.Tn[3].t52 VGND 0.01458f
C7877 XThR.Tn[3].t20 VGND 0.01597f
C7878 XThR.Tn[3].n37 VGND 0.03899f
C7879 XThR.Tn[3].t56 VGND 0.01453f
C7880 XThR.Tn[3].t66 VGND 0.01591f
C7881 XThR.Tn[3].n38 VGND 0.04056f
C7882 XThR.Tn[3].n39 VGND 0.0285f
C7883 XThR.Tn[3].n41 VGND 0.09145f
C7884 XThR.Tn[3].t19 VGND 0.01458f
C7885 XThR.Tn[3].t14 VGND 0.01597f
C7886 XThR.Tn[3].n42 VGND 0.03899f
C7887 XThR.Tn[3].t23 VGND 0.01453f
C7888 XThR.Tn[3].t61 VGND 0.01591f
C7889 XThR.Tn[3].n43 VGND 0.04056f
C7890 XThR.Tn[3].n44 VGND 0.0285f
C7891 XThR.Tn[3].n46 VGND 0.09145f
C7892 XThR.Tn[3].t22 VGND 0.01458f
C7893 XThR.Tn[3].t31 VGND 0.01597f
C7894 XThR.Tn[3].n47 VGND 0.03899f
C7895 XThR.Tn[3].t28 VGND 0.01453f
C7896 XThR.Tn[3].t73 VGND 0.01591f
C7897 XThR.Tn[3].n48 VGND 0.04056f
C7898 XThR.Tn[3].n49 VGND 0.0285f
C7899 XThR.Tn[3].n51 VGND 0.09145f
C7900 XThR.Tn[3].t41 VGND 0.01458f
C7901 XThR.Tn[3].t51 VGND 0.01597f
C7902 XThR.Tn[3].n52 VGND 0.03899f
C7903 XThR.Tn[3].t45 VGND 0.01453f
C7904 XThR.Tn[3].t30 VGND 0.01591f
C7905 XThR.Tn[3].n53 VGND 0.04056f
C7906 XThR.Tn[3].n54 VGND 0.0285f
C7907 XThR.Tn[3].n56 VGND 0.09145f
C7908 XThR.Tn[3].t35 VGND 0.01458f
C7909 XThR.Tn[3].t69 VGND 0.01597f
C7910 XThR.Tn[3].n57 VGND 0.03899f
C7911 XThR.Tn[3].t37 VGND 0.01453f
C7912 XThR.Tn[3].t50 VGND 0.01591f
C7913 XThR.Tn[3].n58 VGND 0.04056f
C7914 XThR.Tn[3].n59 VGND 0.0285f
C7915 XThR.Tn[3].n61 VGND 0.09145f
C7916 XThR.Tn[3].t54 VGND 0.01458f
C7917 XThR.Tn[3].t44 VGND 0.01597f
C7918 XThR.Tn[3].n62 VGND 0.03899f
C7919 XThR.Tn[3].t58 VGND 0.01453f
C7920 XThR.Tn[3].t25 VGND 0.01591f
C7921 XThR.Tn[3].n63 VGND 0.04056f
C7922 XThR.Tn[3].n64 VGND 0.0285f
C7923 XThR.Tn[3].n66 VGND 0.09145f
C7924 XThR.Tn[3].t21 VGND 0.01458f
C7925 XThR.Tn[3].t17 VGND 0.01597f
C7926 XThR.Tn[3].n67 VGND 0.03899f
C7927 XThR.Tn[3].t26 VGND 0.01453f
C7928 XThR.Tn[3].t63 VGND 0.01591f
C7929 XThR.Tn[3].n68 VGND 0.04056f
C7930 XThR.Tn[3].n69 VGND 0.0285f
C7931 XThR.Tn[3].n71 VGND 0.09145f
C7932 XThR.Tn[3].t40 VGND 0.01458f
C7933 XThR.Tn[3].t34 VGND 0.01597f
C7934 XThR.Tn[3].n72 VGND 0.03899f
C7935 XThR.Tn[3].t43 VGND 0.01453f
C7936 XThR.Tn[3].t15 VGND 0.01591f
C7937 XThR.Tn[3].n73 VGND 0.04056f
C7938 XThR.Tn[3].n74 VGND 0.0285f
C7939 XThR.Tn[3].n76 VGND 0.09145f
C7940 XThR.Tn[3].t60 VGND 0.01458f
C7941 XThR.Tn[3].t53 VGND 0.01597f
C7942 XThR.Tn[3].n77 VGND 0.03899f
C7943 XThR.Tn[3].t65 VGND 0.01453f
C7944 XThR.Tn[3].t32 VGND 0.01591f
C7945 XThR.Tn[3].n78 VGND 0.04056f
C7946 XThR.Tn[3].n79 VGND 0.0285f
C7947 XThR.Tn[3].n81 VGND 0.09145f
C7948 XThR.Tn[3].t36 VGND 0.01458f
C7949 XThR.Tn[3].t46 VGND 0.01597f
C7950 XThR.Tn[3].n82 VGND 0.03899f
C7951 XThR.Tn[3].t38 VGND 0.01453f
C7952 XThR.Tn[3].t27 VGND 0.01591f
C7953 XThR.Tn[3].n83 VGND 0.04056f
C7954 XThR.Tn[3].n84 VGND 0.0285f
C7955 XThR.Tn[3].n86 VGND 0.09145f
C7956 XThR.Tn[3].n87 VGND 0.08311f
C7957 XThR.Tn[3].n88 VGND 0.18407f
C7958 XThR.Tn[3].n89 VGND 0.03904f
C7959 XThC.XTB4.Y.t4 VGND 0.02956f
C7960 XThC.XTB4.Y.t13 VGND 0.05016f
C7961 XThC.XTB4.Y.n0 VGND 0.05972f
C7962 XThC.XTB4.Y.t7 VGND 0.02956f
C7963 XThC.XTB4.Y.t17 VGND 0.05016f
C7964 XThC.XTB4.Y.n1 VGND 0.03074f
C7965 XThC.XTB4.Y.t10 VGND 0.02956f
C7966 XThC.XTB4.Y.t2 VGND 0.05016f
C7967 XThC.XTB4.Y.n2 VGND 0.06603f
C7968 XThC.XTB4.Y.t14 VGND 0.02956f
C7969 XThC.XTB4.Y.t3 VGND 0.05016f
C7970 XThC.XTB4.Y.n3 VGND 0.0613f
C7971 XThC.XTB4.Y.n4 VGND 0.03729f
C7972 XThC.XTB4.Y.n5 VGND 0.06174f
C7973 XThC.XTB4.Y.n6 VGND 0.02389f
C7974 XThC.XTB4.Y.n7 VGND 0.02916f
C7975 XThC.XTB4.Y.n8 VGND 0.06603f
C7976 XThC.XTB4.Y.n9 VGND 0.0331f
C7977 XThC.XTB4.Y.n10 VGND 0.06459f
C7978 XThC.XTB4.Y.t5 VGND 0.02956f
C7979 XThC.XTB4.Y.t16 VGND 0.05016f
C7980 XThC.XTB4.Y.n11 VGND 0.06761f
C7981 XThC.XTB4.Y.t9 VGND 0.02956f
C7982 XThC.XTB4.Y.t6 VGND 0.05016f
C7983 XThC.XTB4.Y.t15 VGND 0.02956f
C7984 XThC.XTB4.Y.t12 VGND 0.05016f
C7985 XThC.XTB4.Y.t11 VGND 0.02956f
C7986 XThC.XTB4.Y.t8 VGND 0.05016f
C7987 XThC.XTB4.Y.n12 VGND 0.08416f
C7988 XThC.XTB4.Y.n13 VGND 0.08889f
C7989 XThC.XTB4.Y.n14 VGND 0.03426f
C7990 XThC.XTB4.Y.n15 VGND 0.07234f
C7991 XThC.XTB4.Y.n16 VGND 0.0331f
C7992 XThC.XTB4.Y.n17 VGND 0.02701f
C7993 XThC.XTB4.Y.n18 VGND 0.63971f
C7994 XThC.XTB4.Y.n19 VGND 1.30917f
C7995 XThC.XTB4.Y.t1 VGND 0.06491f
C7996 XThC.XTB4.Y.n20 VGND 0.11223f
C7997 XThC.XTB4.Y.t0 VGND 0.12238f
C7998 XThC.XTB4.Y.n21 VGND 0.16166f
C7999 XThC.Tn[0].t8 VGND 0.01406f
C8000 XThC.Tn[0].t7 VGND 0.01406f
C8001 XThC.Tn[0].n0 VGND 0.02837f
C8002 XThC.Tn[0].t10 VGND 0.01406f
C8003 XThC.Tn[0].t9 VGND 0.01406f
C8004 XThC.Tn[0].n1 VGND 0.0332f
C8005 XThC.Tn[0].n2 VGND 0.09293f
C8006 XThC.Tn[0].n3 VGND 0.02081f
C8007 XThC.Tn[0].n4 VGND 0.02081f
C8008 XThC.Tn[0].n5 VGND 0.02081f
C8009 XThC.Tn[0].n6 VGND 0.03467f
C8010 XThC.Tn[0].n7 VGND 0.09908f
C8011 XThC.Tn[0].n8 VGND 0.06125f
C8012 XThC.Tn[0].n9 VGND 0.06913f
C8013 XThC.Tn[0].t18 VGND 0.01114f
C8014 XThC.Tn[0].t22 VGND 0.01217f
C8015 XThC.Tn[0].n10 VGND 0.02717f
C8016 XThC.Tn[0].n11 VGND 0.01861f
C8017 XThC.Tn[0].n12 VGND 0.06109f
C8018 XThC.Tn[0].t35 VGND 0.01114f
C8019 XThC.Tn[0].t41 VGND 0.01217f
C8020 XThC.Tn[0].n13 VGND 0.02717f
C8021 XThC.Tn[0].n14 VGND 0.01861f
C8022 XThC.Tn[0].n15 VGND 0.06126f
C8023 XThC.Tn[0].n16 VGND 0.10096f
C8024 XThC.Tn[0].t37 VGND 0.01114f
C8025 XThC.Tn[0].t12 VGND 0.01217f
C8026 XThC.Tn[0].n17 VGND 0.02717f
C8027 XThC.Tn[0].n18 VGND 0.01861f
C8028 XThC.Tn[0].n19 VGND 0.06126f
C8029 XThC.Tn[0].n20 VGND 0.10096f
C8030 XThC.Tn[0].t39 VGND 0.01114f
C8031 XThC.Tn[0].t13 VGND 0.01217f
C8032 XThC.Tn[0].n21 VGND 0.02717f
C8033 XThC.Tn[0].n22 VGND 0.01861f
C8034 XThC.Tn[0].n23 VGND 0.06126f
C8035 XThC.Tn[0].n24 VGND 0.10096f
C8036 XThC.Tn[0].t28 VGND 0.01114f
C8037 XThC.Tn[0].t32 VGND 0.01217f
C8038 XThC.Tn[0].n25 VGND 0.02717f
C8039 XThC.Tn[0].n26 VGND 0.01861f
C8040 XThC.Tn[0].n27 VGND 0.06126f
C8041 XThC.Tn[0].n28 VGND 0.10096f
C8042 XThC.Tn[0].t30 VGND 0.01114f
C8043 XThC.Tn[0].t34 VGND 0.01217f
C8044 XThC.Tn[0].n29 VGND 0.02717f
C8045 XThC.Tn[0].n30 VGND 0.01861f
C8046 XThC.Tn[0].n31 VGND 0.06126f
C8047 XThC.Tn[0].n32 VGND 0.10096f
C8048 XThC.Tn[0].t43 VGND 0.01114f
C8049 XThC.Tn[0].t17 VGND 0.01217f
C8050 XThC.Tn[0].n33 VGND 0.02717f
C8051 XThC.Tn[0].n34 VGND 0.01861f
C8052 XThC.Tn[0].n35 VGND 0.06126f
C8053 XThC.Tn[0].n36 VGND 0.10096f
C8054 XThC.Tn[0].t20 VGND 0.01114f
C8055 XThC.Tn[0].t25 VGND 0.01217f
C8056 XThC.Tn[0].n37 VGND 0.02717f
C8057 XThC.Tn[0].n38 VGND 0.01861f
C8058 XThC.Tn[0].n39 VGND 0.06126f
C8059 XThC.Tn[0].n40 VGND 0.10096f
C8060 XThC.Tn[0].t21 VGND 0.01114f
C8061 XThC.Tn[0].t26 VGND 0.01217f
C8062 XThC.Tn[0].n41 VGND 0.02717f
C8063 XThC.Tn[0].n42 VGND 0.01861f
C8064 XThC.Tn[0].n43 VGND 0.06126f
C8065 XThC.Tn[0].n44 VGND 0.10096f
C8066 XThC.Tn[0].t40 VGND 0.01114f
C8067 XThC.Tn[0].t15 VGND 0.01217f
C8068 XThC.Tn[0].n45 VGND 0.02717f
C8069 XThC.Tn[0].n46 VGND 0.01861f
C8070 XThC.Tn[0].n47 VGND 0.06126f
C8071 XThC.Tn[0].n48 VGND 0.10096f
C8072 XThC.Tn[0].t42 VGND 0.01114f
C8073 XThC.Tn[0].t16 VGND 0.01217f
C8074 XThC.Tn[0].n49 VGND 0.02717f
C8075 XThC.Tn[0].n50 VGND 0.01861f
C8076 XThC.Tn[0].n51 VGND 0.06126f
C8077 XThC.Tn[0].n52 VGND 0.10096f
C8078 XThC.Tn[0].t23 VGND 0.01114f
C8079 XThC.Tn[0].t27 VGND 0.01217f
C8080 XThC.Tn[0].n53 VGND 0.02717f
C8081 XThC.Tn[0].n54 VGND 0.01861f
C8082 XThC.Tn[0].n55 VGND 0.06126f
C8083 XThC.Tn[0].n56 VGND 0.10096f
C8084 XThC.Tn[0].t31 VGND 0.01114f
C8085 XThC.Tn[0].t36 VGND 0.01217f
C8086 XThC.Tn[0].n57 VGND 0.02717f
C8087 XThC.Tn[0].n58 VGND 0.01861f
C8088 XThC.Tn[0].n59 VGND 0.06126f
C8089 XThC.Tn[0].n60 VGND 0.10096f
C8090 XThC.Tn[0].t33 VGND 0.01114f
C8091 XThC.Tn[0].t38 VGND 0.01217f
C8092 XThC.Tn[0].n61 VGND 0.02717f
C8093 XThC.Tn[0].n62 VGND 0.01861f
C8094 XThC.Tn[0].n63 VGND 0.06126f
C8095 XThC.Tn[0].n64 VGND 0.10096f
C8096 XThC.Tn[0].t14 VGND 0.01114f
C8097 XThC.Tn[0].t19 VGND 0.01217f
C8098 XThC.Tn[0].n65 VGND 0.02717f
C8099 XThC.Tn[0].n66 VGND 0.01861f
C8100 XThC.Tn[0].n67 VGND 0.06126f
C8101 XThC.Tn[0].n68 VGND 0.10096f
C8102 XThC.Tn[0].t24 VGND 0.01114f
C8103 XThC.Tn[0].t29 VGND 0.01217f
C8104 XThC.Tn[0].n69 VGND 0.02717f
C8105 XThC.Tn[0].n70 VGND 0.01861f
C8106 XThC.Tn[0].n71 VGND 0.06126f
C8107 XThC.Tn[0].n72 VGND 0.10096f
C8108 XThC.Tn[0].n73 VGND 0.70587f
C8109 XThC.Tn[0].n74 VGND 0.07565f
C8110 XThC.Tn[0].n75 VGND 0.02941f
C8111 XThC.Tn[13].t11 VGND 0.01009f
C8112 XThC.Tn[13].t9 VGND 0.01009f
C8113 XThC.Tn[13].n0 VGND 0.02515f
C8114 XThC.Tn[13].t8 VGND 0.01009f
C8115 XThC.Tn[13].t10 VGND 0.01009f
C8116 XThC.Tn[13].n1 VGND 0.02017f
C8117 XThC.Tn[13].n2 VGND 0.04651f
C8118 XThC.Tn[13].t29 VGND 0.0123f
C8119 XThC.Tn[13].t27 VGND 0.01343f
C8120 XThC.Tn[13].n3 VGND 0.02999f
C8121 XThC.Tn[13].n4 VGND 0.02054f
C8122 XThC.Tn[13].n5 VGND 0.06743f
C8123 XThC.Tn[13].t15 VGND 0.0123f
C8124 XThC.Tn[13].t12 VGND 0.01343f
C8125 XThC.Tn[13].n6 VGND 0.02999f
C8126 XThC.Tn[13].n7 VGND 0.02054f
C8127 XThC.Tn[13].n8 VGND 0.06762f
C8128 XThC.Tn[13].n9 VGND 0.11144f
C8129 XThC.Tn[13].t20 VGND 0.0123f
C8130 XThC.Tn[13].t14 VGND 0.01343f
C8131 XThC.Tn[13].n10 VGND 0.02999f
C8132 XThC.Tn[13].n11 VGND 0.02054f
C8133 XThC.Tn[13].n12 VGND 0.06762f
C8134 XThC.Tn[13].n13 VGND 0.11144f
C8135 XThC.Tn[13].t21 VGND 0.0123f
C8136 XThC.Tn[13].t16 VGND 0.01343f
C8137 XThC.Tn[13].n14 VGND 0.02999f
C8138 XThC.Tn[13].n15 VGND 0.02054f
C8139 XThC.Tn[13].n16 VGND 0.06762f
C8140 XThC.Tn[13].n17 VGND 0.11144f
C8141 XThC.Tn[13].t40 VGND 0.0123f
C8142 XThC.Tn[13].t37 VGND 0.01343f
C8143 XThC.Tn[13].n18 VGND 0.02999f
C8144 XThC.Tn[13].n19 VGND 0.02054f
C8145 XThC.Tn[13].n20 VGND 0.06762f
C8146 XThC.Tn[13].n21 VGND 0.11144f
C8147 XThC.Tn[13].t41 VGND 0.0123f
C8148 XThC.Tn[13].t38 VGND 0.01343f
C8149 XThC.Tn[13].n22 VGND 0.02999f
C8150 XThC.Tn[13].n23 VGND 0.02054f
C8151 XThC.Tn[13].n24 VGND 0.06762f
C8152 XThC.Tn[13].n25 VGND 0.11144f
C8153 XThC.Tn[13].t25 VGND 0.0123f
C8154 XThC.Tn[13].t19 VGND 0.01343f
C8155 XThC.Tn[13].n26 VGND 0.02999f
C8156 XThC.Tn[13].n27 VGND 0.02054f
C8157 XThC.Tn[13].n28 VGND 0.06762f
C8158 XThC.Tn[13].n29 VGND 0.11144f
C8159 XThC.Tn[13].t32 VGND 0.0123f
C8160 XThC.Tn[13].t28 VGND 0.01343f
C8161 XThC.Tn[13].n30 VGND 0.02999f
C8162 XThC.Tn[13].n31 VGND 0.02054f
C8163 XThC.Tn[13].n32 VGND 0.06762f
C8164 XThC.Tn[13].n33 VGND 0.11144f
C8165 XThC.Tn[13].t34 VGND 0.0123f
C8166 XThC.Tn[13].t30 VGND 0.01343f
C8167 XThC.Tn[13].n34 VGND 0.02999f
C8168 XThC.Tn[13].n35 VGND 0.02054f
C8169 XThC.Tn[13].n36 VGND 0.06762f
C8170 XThC.Tn[13].n37 VGND 0.11144f
C8171 XThC.Tn[13].t22 VGND 0.0123f
C8172 XThC.Tn[13].t17 VGND 0.01343f
C8173 XThC.Tn[13].n38 VGND 0.02999f
C8174 XThC.Tn[13].n39 VGND 0.02054f
C8175 XThC.Tn[13].n40 VGND 0.06762f
C8176 XThC.Tn[13].n41 VGND 0.11144f
C8177 XThC.Tn[13].t24 VGND 0.0123f
C8178 XThC.Tn[13].t18 VGND 0.01343f
C8179 XThC.Tn[13].n42 VGND 0.02999f
C8180 XThC.Tn[13].n43 VGND 0.02054f
C8181 XThC.Tn[13].n44 VGND 0.06762f
C8182 XThC.Tn[13].n45 VGND 0.11144f
C8183 XThC.Tn[13].t35 VGND 0.0123f
C8184 XThC.Tn[13].t31 VGND 0.01343f
C8185 XThC.Tn[13].n46 VGND 0.02999f
C8186 XThC.Tn[13].n47 VGND 0.02054f
C8187 XThC.Tn[13].n48 VGND 0.06762f
C8188 XThC.Tn[13].n49 VGND 0.11144f
C8189 XThC.Tn[13].t43 VGND 0.0123f
C8190 XThC.Tn[13].t39 VGND 0.01343f
C8191 XThC.Tn[13].n50 VGND 0.02999f
C8192 XThC.Tn[13].n51 VGND 0.02054f
C8193 XThC.Tn[13].n52 VGND 0.06762f
C8194 XThC.Tn[13].n53 VGND 0.11144f
C8195 XThC.Tn[13].t13 VGND 0.0123f
C8196 XThC.Tn[13].t42 VGND 0.01343f
C8197 XThC.Tn[13].n54 VGND 0.02999f
C8198 XThC.Tn[13].n55 VGND 0.02054f
C8199 XThC.Tn[13].n56 VGND 0.06762f
C8200 XThC.Tn[13].n57 VGND 0.11144f
C8201 XThC.Tn[13].t26 VGND 0.0123f
C8202 XThC.Tn[13].t23 VGND 0.01343f
C8203 XThC.Tn[13].n58 VGND 0.02999f
C8204 XThC.Tn[13].n59 VGND 0.02054f
C8205 XThC.Tn[13].n60 VGND 0.06762f
C8206 XThC.Tn[13].n61 VGND 0.11144f
C8207 XThC.Tn[13].t36 VGND 0.0123f
C8208 XThC.Tn[13].t33 VGND 0.01343f
C8209 XThC.Tn[13].n62 VGND 0.02999f
C8210 XThC.Tn[13].n63 VGND 0.02054f
C8211 XThC.Tn[13].n64 VGND 0.06762f
C8212 XThC.Tn[13].n65 VGND 0.11144f
C8213 XThC.Tn[13].n66 VGND 0.57793f
C8214 XThC.Tn[13].n67 VGND 0.20323f
C8215 XThC.Tn[13].t6 VGND 0.01552f
C8216 XThC.Tn[13].t5 VGND 0.01552f
C8217 XThC.Tn[13].n68 VGND 0.03352f
C8218 XThC.Tn[13].t4 VGND 0.01552f
C8219 XThC.Tn[13].t7 VGND 0.01552f
C8220 XThC.Tn[13].n69 VGND 0.05284f
C8221 XThC.Tn[13].n70 VGND 0.13995f
C8222 XThC.Tn[13].n71 VGND 0.0103f
C8223 XThC.Tn[13].t1 VGND 0.01552f
C8224 XThC.Tn[13].t0 VGND 0.01552f
C8225 XThC.Tn[13].n72 VGND 0.04711f
C8226 XThC.Tn[13].t3 VGND 0.01552f
C8227 XThC.Tn[13].t2 VGND 0.01552f
C8228 XThC.Tn[13].n73 VGND 0.03449f
C8229 XThC.Tn[13].n74 VGND 0.15351f
C8230 XThC.Tn[12].t7 VGND 0.01022f
C8231 XThC.Tn[12].t6 VGND 0.01022f
C8232 XThC.Tn[12].n0 VGND 0.02548f
C8233 XThC.Tn[12].t5 VGND 0.01022f
C8234 XThC.Tn[12].t4 VGND 0.01022f
C8235 XThC.Tn[12].n1 VGND 0.02043f
C8236 XThC.Tn[12].n2 VGND 0.0514f
C8237 XThC.Tn[12].t37 VGND 0.01246f
C8238 XThC.Tn[12].t35 VGND 0.01361f
C8239 XThC.Tn[12].n3 VGND 0.03037f
C8240 XThC.Tn[12].n4 VGND 0.02081f
C8241 XThC.Tn[12].n5 VGND 0.0683f
C8242 XThC.Tn[12].t23 VGND 0.01246f
C8243 XThC.Tn[12].t20 VGND 0.01361f
C8244 XThC.Tn[12].n6 VGND 0.03037f
C8245 XThC.Tn[12].n7 VGND 0.02081f
C8246 XThC.Tn[12].n8 VGND 0.06849f
C8247 XThC.Tn[12].n9 VGND 0.11288f
C8248 XThC.Tn[12].t28 VGND 0.01246f
C8249 XThC.Tn[12].t22 VGND 0.01361f
C8250 XThC.Tn[12].n10 VGND 0.03037f
C8251 XThC.Tn[12].n11 VGND 0.02081f
C8252 XThC.Tn[12].n12 VGND 0.06849f
C8253 XThC.Tn[12].n13 VGND 0.11288f
C8254 XThC.Tn[12].t29 VGND 0.01246f
C8255 XThC.Tn[12].t24 VGND 0.01361f
C8256 XThC.Tn[12].n14 VGND 0.03037f
C8257 XThC.Tn[12].n15 VGND 0.02081f
C8258 XThC.Tn[12].n16 VGND 0.06849f
C8259 XThC.Tn[12].n17 VGND 0.11288f
C8260 XThC.Tn[12].t16 VGND 0.01246f
C8261 XThC.Tn[12].t13 VGND 0.01361f
C8262 XThC.Tn[12].n18 VGND 0.03037f
C8263 XThC.Tn[12].n19 VGND 0.02081f
C8264 XThC.Tn[12].n20 VGND 0.06849f
C8265 XThC.Tn[12].n21 VGND 0.11288f
C8266 XThC.Tn[12].t17 VGND 0.01246f
C8267 XThC.Tn[12].t14 VGND 0.01361f
C8268 XThC.Tn[12].n22 VGND 0.03037f
C8269 XThC.Tn[12].n23 VGND 0.02081f
C8270 XThC.Tn[12].n24 VGND 0.06849f
C8271 XThC.Tn[12].n25 VGND 0.11288f
C8272 XThC.Tn[12].t33 VGND 0.01246f
C8273 XThC.Tn[12].t27 VGND 0.01361f
C8274 XThC.Tn[12].n26 VGND 0.03037f
C8275 XThC.Tn[12].n27 VGND 0.02081f
C8276 XThC.Tn[12].n28 VGND 0.06849f
C8277 XThC.Tn[12].n29 VGND 0.11288f
C8278 XThC.Tn[12].t40 VGND 0.01246f
C8279 XThC.Tn[12].t36 VGND 0.01361f
C8280 XThC.Tn[12].n30 VGND 0.03037f
C8281 XThC.Tn[12].n31 VGND 0.02081f
C8282 XThC.Tn[12].n32 VGND 0.06849f
C8283 XThC.Tn[12].n33 VGND 0.11288f
C8284 XThC.Tn[12].t42 VGND 0.01246f
C8285 XThC.Tn[12].t38 VGND 0.01361f
C8286 XThC.Tn[12].n34 VGND 0.03037f
C8287 XThC.Tn[12].n35 VGND 0.02081f
C8288 XThC.Tn[12].n36 VGND 0.06849f
C8289 XThC.Tn[12].n37 VGND 0.11288f
C8290 XThC.Tn[12].t30 VGND 0.01246f
C8291 XThC.Tn[12].t25 VGND 0.01361f
C8292 XThC.Tn[12].n38 VGND 0.03037f
C8293 XThC.Tn[12].n39 VGND 0.02081f
C8294 XThC.Tn[12].n40 VGND 0.06849f
C8295 XThC.Tn[12].n41 VGND 0.11288f
C8296 XThC.Tn[12].t32 VGND 0.01246f
C8297 XThC.Tn[12].t26 VGND 0.01361f
C8298 XThC.Tn[12].n42 VGND 0.03037f
C8299 XThC.Tn[12].n43 VGND 0.02081f
C8300 XThC.Tn[12].n44 VGND 0.06849f
C8301 XThC.Tn[12].n45 VGND 0.11288f
C8302 XThC.Tn[12].t43 VGND 0.01246f
C8303 XThC.Tn[12].t39 VGND 0.01361f
C8304 XThC.Tn[12].n46 VGND 0.03037f
C8305 XThC.Tn[12].n47 VGND 0.02081f
C8306 XThC.Tn[12].n48 VGND 0.06849f
C8307 XThC.Tn[12].n49 VGND 0.11288f
C8308 XThC.Tn[12].t19 VGND 0.01246f
C8309 XThC.Tn[12].t15 VGND 0.01361f
C8310 XThC.Tn[12].n50 VGND 0.03037f
C8311 XThC.Tn[12].n51 VGND 0.02081f
C8312 XThC.Tn[12].n52 VGND 0.06849f
C8313 XThC.Tn[12].n53 VGND 0.11288f
C8314 XThC.Tn[12].t21 VGND 0.01246f
C8315 XThC.Tn[12].t18 VGND 0.01361f
C8316 XThC.Tn[12].n54 VGND 0.03037f
C8317 XThC.Tn[12].n55 VGND 0.02081f
C8318 XThC.Tn[12].n56 VGND 0.06849f
C8319 XThC.Tn[12].n57 VGND 0.11288f
C8320 XThC.Tn[12].t34 VGND 0.01246f
C8321 XThC.Tn[12].t31 VGND 0.01361f
C8322 XThC.Tn[12].n58 VGND 0.03037f
C8323 XThC.Tn[12].n59 VGND 0.02081f
C8324 XThC.Tn[12].n60 VGND 0.06849f
C8325 XThC.Tn[12].n61 VGND 0.11288f
C8326 XThC.Tn[12].t12 VGND 0.01246f
C8327 XThC.Tn[12].t41 VGND 0.01361f
C8328 XThC.Tn[12].n62 VGND 0.03037f
C8329 XThC.Tn[12].n63 VGND 0.02081f
C8330 XThC.Tn[12].n64 VGND 0.06849f
C8331 XThC.Tn[12].n65 VGND 0.11288f
C8332 XThC.Tn[12].n66 VGND 0.53677f
C8333 XThC.Tn[12].n67 VGND 0.19068f
C8334 XThC.Tn[12].t1 VGND 0.01572f
C8335 XThC.Tn[12].t2 VGND 0.01572f
C8336 XThC.Tn[12].n68 VGND 0.03396f
C8337 XThC.Tn[12].t0 VGND 0.01572f
C8338 XThC.Tn[12].t3 VGND 0.01572f
C8339 XThC.Tn[12].n69 VGND 0.05168f
C8340 XThC.Tn[12].n70 VGND 0.1436f
C8341 XThC.Tn[12].n71 VGND 0.02258f
C8342 XThC.Tn[12].t9 VGND 0.01572f
C8343 XThC.Tn[12].t8 VGND 0.01572f
C8344 XThC.Tn[12].n72 VGND 0.04772f
C8345 XThC.Tn[12].t11 VGND 0.01572f
C8346 XThC.Tn[12].t10 VGND 0.01572f
C8347 XThC.Tn[12].n73 VGND 0.03494f
C8348 XThC.Tn[12].n74 VGND 0.15549f
C8349 XThC.Tn[11].t8 VGND 0.01038f
C8350 XThC.Tn[11].t11 VGND 0.01038f
C8351 XThC.Tn[11].n0 VGND 0.0259f
C8352 XThC.Tn[11].t7 VGND 0.01038f
C8353 XThC.Tn[11].t5 VGND 0.01038f
C8354 XThC.Tn[11].n1 VGND 0.02077f
C8355 XThC.Tn[11].n2 VGND 0.04789f
C8356 XThC.Tn[11].t20 VGND 0.01266f
C8357 XThC.Tn[11].t18 VGND 0.01383f
C8358 XThC.Tn[11].n3 VGND 0.03087f
C8359 XThC.Tn[11].n4 VGND 0.02115f
C8360 XThC.Tn[11].n5 VGND 0.06943f
C8361 XThC.Tn[11].t38 VGND 0.01266f
C8362 XThC.Tn[11].t35 VGND 0.01383f
C8363 XThC.Tn[11].n6 VGND 0.03087f
C8364 XThC.Tn[11].n7 VGND 0.02115f
C8365 XThC.Tn[11].n8 VGND 0.06962f
C8366 XThC.Tn[11].n9 VGND 0.11473f
C8367 XThC.Tn[11].t43 VGND 0.01266f
C8368 XThC.Tn[11].t37 VGND 0.01383f
C8369 XThC.Tn[11].n10 VGND 0.03087f
C8370 XThC.Tn[11].n11 VGND 0.02115f
C8371 XThC.Tn[11].n12 VGND 0.06962f
C8372 XThC.Tn[11].n13 VGND 0.11473f
C8373 XThC.Tn[11].t12 VGND 0.01266f
C8374 XThC.Tn[11].t39 VGND 0.01383f
C8375 XThC.Tn[11].n14 VGND 0.03087f
C8376 XThC.Tn[11].n15 VGND 0.02115f
C8377 XThC.Tn[11].n16 VGND 0.06962f
C8378 XThC.Tn[11].n17 VGND 0.11473f
C8379 XThC.Tn[11].t31 VGND 0.01266f
C8380 XThC.Tn[11].t28 VGND 0.01383f
C8381 XThC.Tn[11].n18 VGND 0.03087f
C8382 XThC.Tn[11].n19 VGND 0.02115f
C8383 XThC.Tn[11].n20 VGND 0.06962f
C8384 XThC.Tn[11].n21 VGND 0.11473f
C8385 XThC.Tn[11].t32 VGND 0.01266f
C8386 XThC.Tn[11].t29 VGND 0.01383f
C8387 XThC.Tn[11].n22 VGND 0.03087f
C8388 XThC.Tn[11].n23 VGND 0.02115f
C8389 XThC.Tn[11].n24 VGND 0.06962f
C8390 XThC.Tn[11].n25 VGND 0.11473f
C8391 XThC.Tn[11].t16 VGND 0.01266f
C8392 XThC.Tn[11].t42 VGND 0.01383f
C8393 XThC.Tn[11].n26 VGND 0.03087f
C8394 XThC.Tn[11].n27 VGND 0.02115f
C8395 XThC.Tn[11].n28 VGND 0.06962f
C8396 XThC.Tn[11].n29 VGND 0.11473f
C8397 XThC.Tn[11].t23 VGND 0.01266f
C8398 XThC.Tn[11].t19 VGND 0.01383f
C8399 XThC.Tn[11].n30 VGND 0.03087f
C8400 XThC.Tn[11].n31 VGND 0.02115f
C8401 XThC.Tn[11].n32 VGND 0.06962f
C8402 XThC.Tn[11].n33 VGND 0.11473f
C8403 XThC.Tn[11].t25 VGND 0.01266f
C8404 XThC.Tn[11].t21 VGND 0.01383f
C8405 XThC.Tn[11].n34 VGND 0.03087f
C8406 XThC.Tn[11].n35 VGND 0.02115f
C8407 XThC.Tn[11].n36 VGND 0.06962f
C8408 XThC.Tn[11].n37 VGND 0.11473f
C8409 XThC.Tn[11].t13 VGND 0.01266f
C8410 XThC.Tn[11].t40 VGND 0.01383f
C8411 XThC.Tn[11].n38 VGND 0.03087f
C8412 XThC.Tn[11].n39 VGND 0.02115f
C8413 XThC.Tn[11].n40 VGND 0.06962f
C8414 XThC.Tn[11].n41 VGND 0.11473f
C8415 XThC.Tn[11].t15 VGND 0.01266f
C8416 XThC.Tn[11].t41 VGND 0.01383f
C8417 XThC.Tn[11].n42 VGND 0.03087f
C8418 XThC.Tn[11].n43 VGND 0.02115f
C8419 XThC.Tn[11].n44 VGND 0.06962f
C8420 XThC.Tn[11].n45 VGND 0.11473f
C8421 XThC.Tn[11].t26 VGND 0.01266f
C8422 XThC.Tn[11].t22 VGND 0.01383f
C8423 XThC.Tn[11].n46 VGND 0.03087f
C8424 XThC.Tn[11].n47 VGND 0.02115f
C8425 XThC.Tn[11].n48 VGND 0.06962f
C8426 XThC.Tn[11].n49 VGND 0.11473f
C8427 XThC.Tn[11].t34 VGND 0.01266f
C8428 XThC.Tn[11].t30 VGND 0.01383f
C8429 XThC.Tn[11].n50 VGND 0.03087f
C8430 XThC.Tn[11].n51 VGND 0.02115f
C8431 XThC.Tn[11].n52 VGND 0.06962f
C8432 XThC.Tn[11].n53 VGND 0.11473f
C8433 XThC.Tn[11].t36 VGND 0.01266f
C8434 XThC.Tn[11].t33 VGND 0.01383f
C8435 XThC.Tn[11].n54 VGND 0.03087f
C8436 XThC.Tn[11].n55 VGND 0.02115f
C8437 XThC.Tn[11].n56 VGND 0.06962f
C8438 XThC.Tn[11].n57 VGND 0.11473f
C8439 XThC.Tn[11].t17 VGND 0.01266f
C8440 XThC.Tn[11].t14 VGND 0.01383f
C8441 XThC.Tn[11].n58 VGND 0.03087f
C8442 XThC.Tn[11].n59 VGND 0.02115f
C8443 XThC.Tn[11].n60 VGND 0.06962f
C8444 XThC.Tn[11].n61 VGND 0.11473f
C8445 XThC.Tn[11].t27 VGND 0.01266f
C8446 XThC.Tn[11].t24 VGND 0.01383f
C8447 XThC.Tn[11].n62 VGND 0.03087f
C8448 XThC.Tn[11].n63 VGND 0.02115f
C8449 XThC.Tn[11].n64 VGND 0.06962f
C8450 XThC.Tn[11].n65 VGND 0.11473f
C8451 XThC.Tn[11].n66 VGND 0.53249f
C8452 XThC.Tn[11].n67 VGND 0.20859f
C8453 XThC.Tn[11].t6 VGND 0.01597f
C8454 XThC.Tn[11].t10 VGND 0.01597f
C8455 XThC.Tn[11].n68 VGND 0.03451f
C8456 XThC.Tn[11].t4 VGND 0.01597f
C8457 XThC.Tn[11].t9 VGND 0.01597f
C8458 XThC.Tn[11].n69 VGND 0.05441f
C8459 XThC.Tn[11].n70 VGND 0.14409f
C8460 XThC.Tn[11].n71 VGND 0.01061f
C8461 XThC.Tn[11].t2 VGND 0.01597f
C8462 XThC.Tn[11].t1 VGND 0.01597f
C8463 XThC.Tn[11].n72 VGND 0.03551f
C8464 XThC.Tn[11].t0 VGND 0.01597f
C8465 XThC.Tn[11].t3 VGND 0.01597f
C8466 XThC.Tn[11].n73 VGND 0.0485f
C8467 XThC.Tn[11].n74 VGND 0.15805f
C8468 XThC.Tn[9].t9 VGND 0.01057f
C8469 XThC.Tn[9].t8 VGND 0.01057f
C8470 XThC.Tn[9].n0 VGND 0.02637f
C8471 XThC.Tn[9].t10 VGND 0.01057f
C8472 XThC.Tn[9].t11 VGND 0.01057f
C8473 XThC.Tn[9].n1 VGND 0.02114f
C8474 XThC.Tn[9].n2 VGND 0.04875f
C8475 XThC.Tn[9].t26 VGND 0.01289f
C8476 XThC.Tn[9].t12 VGND 0.01408f
C8477 XThC.Tn[9].n3 VGND 0.03143f
C8478 XThC.Tn[9].n4 VGND 0.02153f
C8479 XThC.Tn[9].n5 VGND 0.07068f
C8480 XThC.Tn[9].t13 VGND 0.01289f
C8481 XThC.Tn[9].t30 VGND 0.01408f
C8482 XThC.Tn[9].n6 VGND 0.03143f
C8483 XThC.Tn[9].n7 VGND 0.02153f
C8484 XThC.Tn[9].n8 VGND 0.07088f
C8485 XThC.Tn[9].n9 VGND 0.11681f
C8486 XThC.Tn[9].t15 VGND 0.01289f
C8487 XThC.Tn[9].t34 VGND 0.01408f
C8488 XThC.Tn[9].n10 VGND 0.03143f
C8489 XThC.Tn[9].n11 VGND 0.02153f
C8490 XThC.Tn[9].n12 VGND 0.07088f
C8491 XThC.Tn[9].n13 VGND 0.11681f
C8492 XThC.Tn[9].t17 VGND 0.01289f
C8493 XThC.Tn[9].t35 VGND 0.01408f
C8494 XThC.Tn[9].n14 VGND 0.03143f
C8495 XThC.Tn[9].n15 VGND 0.02153f
C8496 XThC.Tn[9].n16 VGND 0.07088f
C8497 XThC.Tn[9].n17 VGND 0.11681f
C8498 XThC.Tn[9].t39 VGND 0.01289f
C8499 XThC.Tn[9].t24 VGND 0.01408f
C8500 XThC.Tn[9].n18 VGND 0.03143f
C8501 XThC.Tn[9].n19 VGND 0.02153f
C8502 XThC.Tn[9].n20 VGND 0.07088f
C8503 XThC.Tn[9].n21 VGND 0.11681f
C8504 XThC.Tn[9].t40 VGND 0.01289f
C8505 XThC.Tn[9].t25 VGND 0.01408f
C8506 XThC.Tn[9].n22 VGND 0.03143f
C8507 XThC.Tn[9].n23 VGND 0.02153f
C8508 XThC.Tn[9].n24 VGND 0.07088f
C8509 XThC.Tn[9].n25 VGND 0.11681f
C8510 XThC.Tn[9].t22 VGND 0.01289f
C8511 XThC.Tn[9].t38 VGND 0.01408f
C8512 XThC.Tn[9].n26 VGND 0.03143f
C8513 XThC.Tn[9].n27 VGND 0.02153f
C8514 XThC.Tn[9].n28 VGND 0.07088f
C8515 XThC.Tn[9].n29 VGND 0.11681f
C8516 XThC.Tn[9].t28 VGND 0.01289f
C8517 XThC.Tn[9].t14 VGND 0.01408f
C8518 XThC.Tn[9].n30 VGND 0.03143f
C8519 XThC.Tn[9].n31 VGND 0.02153f
C8520 XThC.Tn[9].n32 VGND 0.07088f
C8521 XThC.Tn[9].n33 VGND 0.11681f
C8522 XThC.Tn[9].t31 VGND 0.01289f
C8523 XThC.Tn[9].t16 VGND 0.01408f
C8524 XThC.Tn[9].n34 VGND 0.03143f
C8525 XThC.Tn[9].n35 VGND 0.02153f
C8526 XThC.Tn[9].n36 VGND 0.07088f
C8527 XThC.Tn[9].n37 VGND 0.11681f
C8528 XThC.Tn[9].t19 VGND 0.01289f
C8529 XThC.Tn[9].t36 VGND 0.01408f
C8530 XThC.Tn[9].n38 VGND 0.03143f
C8531 XThC.Tn[9].n39 VGND 0.02153f
C8532 XThC.Tn[9].n40 VGND 0.07088f
C8533 XThC.Tn[9].n41 VGND 0.11681f
C8534 XThC.Tn[9].t21 VGND 0.01289f
C8535 XThC.Tn[9].t37 VGND 0.01408f
C8536 XThC.Tn[9].n42 VGND 0.03143f
C8537 XThC.Tn[9].n43 VGND 0.02153f
C8538 XThC.Tn[9].n44 VGND 0.07088f
C8539 XThC.Tn[9].n45 VGND 0.11681f
C8540 XThC.Tn[9].t32 VGND 0.01289f
C8541 XThC.Tn[9].t18 VGND 0.01408f
C8542 XThC.Tn[9].n46 VGND 0.03143f
C8543 XThC.Tn[9].n47 VGND 0.02153f
C8544 XThC.Tn[9].n48 VGND 0.07088f
C8545 XThC.Tn[9].n49 VGND 0.11681f
C8546 XThC.Tn[9].t42 VGND 0.01289f
C8547 XThC.Tn[9].t27 VGND 0.01408f
C8548 XThC.Tn[9].n50 VGND 0.03143f
C8549 XThC.Tn[9].n51 VGND 0.02153f
C8550 XThC.Tn[9].n52 VGND 0.07088f
C8551 XThC.Tn[9].n53 VGND 0.11681f
C8552 XThC.Tn[9].t43 VGND 0.01289f
C8553 XThC.Tn[9].t29 VGND 0.01408f
C8554 XThC.Tn[9].n54 VGND 0.03143f
C8555 XThC.Tn[9].n55 VGND 0.02153f
C8556 XThC.Tn[9].n56 VGND 0.07088f
C8557 XThC.Tn[9].n57 VGND 0.11681f
C8558 XThC.Tn[9].t23 VGND 0.01289f
C8559 XThC.Tn[9].t41 VGND 0.01408f
C8560 XThC.Tn[9].n58 VGND 0.03143f
C8561 XThC.Tn[9].n59 VGND 0.02153f
C8562 XThC.Tn[9].n60 VGND 0.07088f
C8563 XThC.Tn[9].n61 VGND 0.11681f
C8564 XThC.Tn[9].t33 VGND 0.01289f
C8565 XThC.Tn[9].t20 VGND 0.01408f
C8566 XThC.Tn[9].n62 VGND 0.03143f
C8567 XThC.Tn[9].n63 VGND 0.02153f
C8568 XThC.Tn[9].n64 VGND 0.07088f
C8569 XThC.Tn[9].n65 VGND 0.11681f
C8570 XThC.Tn[9].n66 VGND 0.50212f
C8571 XThC.Tn[9].n67 VGND 0.21237f
C8572 XThC.Tn[9].t4 VGND 0.01626f
C8573 XThC.Tn[9].t7 VGND 0.01626f
C8574 XThC.Tn[9].n68 VGND 0.03514f
C8575 XThC.Tn[9].t6 VGND 0.01626f
C8576 XThC.Tn[9].t5 VGND 0.01626f
C8577 XThC.Tn[9].n69 VGND 0.05539f
C8578 XThC.Tn[9].n70 VGND 0.1467f
C8579 XThC.Tn[9].n71 VGND 0.0108f
C8580 XThC.Tn[9].t1 VGND 0.01626f
C8581 XThC.Tn[9].t0 VGND 0.01626f
C8582 XThC.Tn[9].n72 VGND 0.04938f
C8583 XThC.Tn[9].t3 VGND 0.01626f
C8584 XThC.Tn[9].t2 VGND 0.01626f
C8585 XThC.Tn[9].n73 VGND 0.03615f
C8586 XThC.Tn[9].n74 VGND 0.16091f
C8587 XThC.Tn[5].t7 VGND 0.01432f
C8588 XThC.Tn[5].t6 VGND 0.01432f
C8589 XThC.Tn[5].n0 VGND 0.02891f
C8590 XThC.Tn[5].t5 VGND 0.01432f
C8591 XThC.Tn[5].t4 VGND 0.01432f
C8592 XThC.Tn[5].n1 VGND 0.03382f
C8593 XThC.Tn[5].n2 VGND 0.10145f
C8594 XThC.Tn[5].n3 VGND 0.0212f
C8595 XThC.Tn[5].n4 VGND 0.03532f
C8596 XThC.Tn[5].n5 VGND 0.0212f
C8597 XThC.Tn[5].n6 VGND 0.10095f
C8598 XThC.Tn[5].n7 VGND 0.0212f
C8599 XThC.Tn[5].n8 VGND 0.06241f
C8600 XThC.Tn[5].n9 VGND 0.07043f
C8601 XThC.Tn[5].t15 VGND 0.01135f
C8602 XThC.Tn[5].t33 VGND 0.0124f
C8603 XThC.Tn[5].n10 VGND 0.02768f
C8604 XThC.Tn[5].n11 VGND 0.01896f
C8605 XThC.Tn[5].n12 VGND 0.06224f
C8606 XThC.Tn[5].t34 VGND 0.01135f
C8607 XThC.Tn[5].t19 VGND 0.0124f
C8608 XThC.Tn[5].n13 VGND 0.02768f
C8609 XThC.Tn[5].n14 VGND 0.01896f
C8610 XThC.Tn[5].n15 VGND 0.06241f
C8611 XThC.Tn[5].n16 VGND 0.10286f
C8612 XThC.Tn[5].t36 VGND 0.01135f
C8613 XThC.Tn[5].t23 VGND 0.0124f
C8614 XThC.Tn[5].n17 VGND 0.02768f
C8615 XThC.Tn[5].n18 VGND 0.01896f
C8616 XThC.Tn[5].n19 VGND 0.06241f
C8617 XThC.Tn[5].n20 VGND 0.10286f
C8618 XThC.Tn[5].t38 VGND 0.01135f
C8619 XThC.Tn[5].t24 VGND 0.0124f
C8620 XThC.Tn[5].n21 VGND 0.02768f
C8621 XThC.Tn[5].n22 VGND 0.01896f
C8622 XThC.Tn[5].n23 VGND 0.06241f
C8623 XThC.Tn[5].n24 VGND 0.10286f
C8624 XThC.Tn[5].t28 VGND 0.01135f
C8625 XThC.Tn[5].t13 VGND 0.0124f
C8626 XThC.Tn[5].n25 VGND 0.02768f
C8627 XThC.Tn[5].n26 VGND 0.01896f
C8628 XThC.Tn[5].n27 VGND 0.06241f
C8629 XThC.Tn[5].n28 VGND 0.10286f
C8630 XThC.Tn[5].t29 VGND 0.01135f
C8631 XThC.Tn[5].t14 VGND 0.0124f
C8632 XThC.Tn[5].n29 VGND 0.02768f
C8633 XThC.Tn[5].n30 VGND 0.01896f
C8634 XThC.Tn[5].n31 VGND 0.06241f
C8635 XThC.Tn[5].n32 VGND 0.10286f
C8636 XThC.Tn[5].t43 VGND 0.01135f
C8637 XThC.Tn[5].t27 VGND 0.0124f
C8638 XThC.Tn[5].n33 VGND 0.02768f
C8639 XThC.Tn[5].n34 VGND 0.01896f
C8640 XThC.Tn[5].n35 VGND 0.06241f
C8641 XThC.Tn[5].n36 VGND 0.10286f
C8642 XThC.Tn[5].t17 VGND 0.01135f
C8643 XThC.Tn[5].t35 VGND 0.0124f
C8644 XThC.Tn[5].n37 VGND 0.02768f
C8645 XThC.Tn[5].n38 VGND 0.01896f
C8646 XThC.Tn[5].n39 VGND 0.06241f
C8647 XThC.Tn[5].n40 VGND 0.10286f
C8648 XThC.Tn[5].t20 VGND 0.01135f
C8649 XThC.Tn[5].t37 VGND 0.0124f
C8650 XThC.Tn[5].n41 VGND 0.02768f
C8651 XThC.Tn[5].n42 VGND 0.01896f
C8652 XThC.Tn[5].n43 VGND 0.06241f
C8653 XThC.Tn[5].n44 VGND 0.10286f
C8654 XThC.Tn[5].t40 VGND 0.01135f
C8655 XThC.Tn[5].t25 VGND 0.0124f
C8656 XThC.Tn[5].n45 VGND 0.02768f
C8657 XThC.Tn[5].n46 VGND 0.01896f
C8658 XThC.Tn[5].n47 VGND 0.06241f
C8659 XThC.Tn[5].n48 VGND 0.10286f
C8660 XThC.Tn[5].t42 VGND 0.01135f
C8661 XThC.Tn[5].t26 VGND 0.0124f
C8662 XThC.Tn[5].n49 VGND 0.02768f
C8663 XThC.Tn[5].n50 VGND 0.01896f
C8664 XThC.Tn[5].n51 VGND 0.06241f
C8665 XThC.Tn[5].n52 VGND 0.10286f
C8666 XThC.Tn[5].t21 VGND 0.01135f
C8667 XThC.Tn[5].t39 VGND 0.0124f
C8668 XThC.Tn[5].n53 VGND 0.02768f
C8669 XThC.Tn[5].n54 VGND 0.01896f
C8670 XThC.Tn[5].n55 VGND 0.06241f
C8671 XThC.Tn[5].n56 VGND 0.10286f
C8672 XThC.Tn[5].t31 VGND 0.01135f
C8673 XThC.Tn[5].t16 VGND 0.0124f
C8674 XThC.Tn[5].n57 VGND 0.02768f
C8675 XThC.Tn[5].n58 VGND 0.01896f
C8676 XThC.Tn[5].n59 VGND 0.06241f
C8677 XThC.Tn[5].n60 VGND 0.10286f
C8678 XThC.Tn[5].t32 VGND 0.01135f
C8679 XThC.Tn[5].t18 VGND 0.0124f
C8680 XThC.Tn[5].n61 VGND 0.02768f
C8681 XThC.Tn[5].n62 VGND 0.01896f
C8682 XThC.Tn[5].n63 VGND 0.06241f
C8683 XThC.Tn[5].n64 VGND 0.10286f
C8684 XThC.Tn[5].t12 VGND 0.01135f
C8685 XThC.Tn[5].t30 VGND 0.0124f
C8686 XThC.Tn[5].n65 VGND 0.02768f
C8687 XThC.Tn[5].n66 VGND 0.01896f
C8688 XThC.Tn[5].n67 VGND 0.06241f
C8689 XThC.Tn[5].n68 VGND 0.10286f
C8690 XThC.Tn[5].t22 VGND 0.01135f
C8691 XThC.Tn[5].t41 VGND 0.0124f
C8692 XThC.Tn[5].n69 VGND 0.02768f
C8693 XThC.Tn[5].n70 VGND 0.01896f
C8694 XThC.Tn[5].n71 VGND 0.06241f
C8695 XThC.Tn[5].n72 VGND 0.10286f
C8696 XThC.Tn[5].n73 VGND 0.11705f
C8697 XThR.Tn[9].t10 VGND 0.01974f
C8698 XThR.Tn[9].t8 VGND 0.01974f
C8699 XThR.Tn[9].n0 VGND 0.05994f
C8700 XThR.Tn[9].t11 VGND 0.01974f
C8701 XThR.Tn[9].t9 VGND 0.01974f
C8702 XThR.Tn[9].n1 VGND 0.04388f
C8703 XThR.Tn[9].n2 VGND 0.19953f
C8704 XThR.Tn[9].t5 VGND 0.01283f
C8705 XThR.Tn[9].t7 VGND 0.01283f
C8706 XThR.Tn[9].n3 VGND 0.032f
C8707 XThR.Tn[9].t4 VGND 0.01283f
C8708 XThR.Tn[9].t6 VGND 0.01283f
C8709 XThR.Tn[9].n4 VGND 0.02566f
C8710 XThR.Tn[9].n5 VGND 0.06456f
C8711 XThR.Tn[9].t17 VGND 0.01543f
C8712 XThR.Tn[9].t71 VGND 0.01689f
C8713 XThR.Tn[9].n6 VGND 0.04125f
C8714 XThR.Tn[9].n7 VGND 0.07925f
C8715 XThR.Tn[9].t35 VGND 0.01543f
C8716 XThR.Tn[9].t28 VGND 0.01689f
C8717 XThR.Tn[9].n8 VGND 0.04125f
C8718 XThR.Tn[9].t50 VGND 0.01538f
C8719 XThR.Tn[9].t19 VGND 0.01684f
C8720 XThR.Tn[9].n9 VGND 0.04292f
C8721 XThR.Tn[9].n10 VGND 0.03015f
C8722 XThR.Tn[9].n12 VGND 0.09677f
C8723 XThR.Tn[9].t72 VGND 0.01543f
C8724 XThR.Tn[9].t64 VGND 0.01689f
C8725 XThR.Tn[9].n13 VGND 0.04125f
C8726 XThR.Tn[9].t26 VGND 0.01538f
C8727 XThR.Tn[9].t59 VGND 0.01684f
C8728 XThR.Tn[9].n14 VGND 0.04292f
C8729 XThR.Tn[9].n15 VGND 0.03015f
C8730 XThR.Tn[9].n17 VGND 0.09677f
C8731 XThR.Tn[9].t29 VGND 0.01543f
C8732 XThR.Tn[9].t21 VGND 0.01689f
C8733 XThR.Tn[9].n18 VGND 0.04125f
C8734 XThR.Tn[9].t41 VGND 0.01538f
C8735 XThR.Tn[9].t15 VGND 0.01684f
C8736 XThR.Tn[9].n19 VGND 0.04292f
C8737 XThR.Tn[9].n20 VGND 0.03015f
C8738 XThR.Tn[9].n22 VGND 0.09677f
C8739 XThR.Tn[9].t56 VGND 0.01543f
C8740 XThR.Tn[9].t46 VGND 0.01689f
C8741 XThR.Tn[9].n23 VGND 0.04125f
C8742 XThR.Tn[9].t73 VGND 0.01538f
C8743 XThR.Tn[9].t42 VGND 0.01684f
C8744 XThR.Tn[9].n24 VGND 0.04292f
C8745 XThR.Tn[9].n25 VGND 0.03015f
C8746 XThR.Tn[9].n27 VGND 0.09677f
C8747 XThR.Tn[9].t31 VGND 0.01543f
C8748 XThR.Tn[9].t23 VGND 0.01689f
C8749 XThR.Tn[9].n28 VGND 0.04125f
C8750 XThR.Tn[9].t44 VGND 0.01538f
C8751 XThR.Tn[9].t16 VGND 0.01684f
C8752 XThR.Tn[9].n29 VGND 0.04292f
C8753 XThR.Tn[9].n30 VGND 0.03015f
C8754 XThR.Tn[9].n32 VGND 0.09677f
C8755 XThR.Tn[9].t67 VGND 0.01543f
C8756 XThR.Tn[9].t37 VGND 0.01689f
C8757 XThR.Tn[9].n33 VGND 0.04125f
C8758 XThR.Tn[9].t20 VGND 0.01538f
C8759 XThR.Tn[9].t33 VGND 0.01684f
C8760 XThR.Tn[9].n34 VGND 0.04292f
C8761 XThR.Tn[9].n35 VGND 0.03015f
C8762 XThR.Tn[9].n37 VGND 0.09677f
C8763 XThR.Tn[9].t36 VGND 0.01543f
C8764 XThR.Tn[9].t32 VGND 0.01689f
C8765 XThR.Tn[9].n38 VGND 0.04125f
C8766 XThR.Tn[9].t51 VGND 0.01538f
C8767 XThR.Tn[9].t25 VGND 0.01684f
C8768 XThR.Tn[9].n39 VGND 0.04292f
C8769 XThR.Tn[9].n40 VGND 0.03015f
C8770 XThR.Tn[9].n42 VGND 0.09677f
C8771 XThR.Tn[9].t39 VGND 0.01543f
C8772 XThR.Tn[9].t45 VGND 0.01689f
C8773 XThR.Tn[9].n43 VGND 0.04125f
C8774 XThR.Tn[9].t55 VGND 0.01538f
C8775 XThR.Tn[9].t40 VGND 0.01684f
C8776 XThR.Tn[9].n44 VGND 0.04292f
C8777 XThR.Tn[9].n45 VGND 0.03015f
C8778 XThR.Tn[9].n47 VGND 0.09677f
C8779 XThR.Tn[9].t58 VGND 0.01543f
C8780 XThR.Tn[9].t66 VGND 0.01689f
C8781 XThR.Tn[9].n48 VGND 0.04125f
C8782 XThR.Tn[9].t13 VGND 0.01538f
C8783 XThR.Tn[9].t60 VGND 0.01684f
C8784 XThR.Tn[9].n49 VGND 0.04292f
C8785 XThR.Tn[9].n50 VGND 0.03015f
C8786 XThR.Tn[9].n52 VGND 0.09677f
C8787 XThR.Tn[9].t48 VGND 0.01543f
C8788 XThR.Tn[9].t24 VGND 0.01689f
C8789 XThR.Tn[9].n53 VGND 0.04125f
C8790 XThR.Tn[9].t65 VGND 0.01538f
C8791 XThR.Tn[9].t18 VGND 0.01684f
C8792 XThR.Tn[9].n54 VGND 0.04292f
C8793 XThR.Tn[9].n55 VGND 0.03015f
C8794 XThR.Tn[9].n57 VGND 0.09677f
C8795 XThR.Tn[9].t70 VGND 0.01543f
C8796 XThR.Tn[9].t62 VGND 0.01689f
C8797 XThR.Tn[9].n58 VGND 0.04125f
C8798 XThR.Tn[9].t22 VGND 0.01538f
C8799 XThR.Tn[9].t52 VGND 0.01684f
C8800 XThR.Tn[9].n59 VGND 0.04292f
C8801 XThR.Tn[9].n60 VGND 0.03015f
C8802 XThR.Tn[9].n62 VGND 0.09677f
C8803 XThR.Tn[9].t38 VGND 0.01543f
C8804 XThR.Tn[9].t34 VGND 0.01689f
C8805 XThR.Tn[9].n63 VGND 0.04125f
C8806 XThR.Tn[9].t53 VGND 0.01538f
C8807 XThR.Tn[9].t27 VGND 0.01684f
C8808 XThR.Tn[9].n64 VGND 0.04292f
C8809 XThR.Tn[9].n65 VGND 0.03015f
C8810 XThR.Tn[9].n67 VGND 0.09677f
C8811 XThR.Tn[9].t57 VGND 0.01543f
C8812 XThR.Tn[9].t47 VGND 0.01689f
C8813 XThR.Tn[9].n68 VGND 0.04125f
C8814 XThR.Tn[9].t12 VGND 0.01538f
C8815 XThR.Tn[9].t43 VGND 0.01684f
C8816 XThR.Tn[9].n69 VGND 0.04292f
C8817 XThR.Tn[9].n70 VGND 0.03015f
C8818 XThR.Tn[9].n72 VGND 0.09677f
C8819 XThR.Tn[9].t14 VGND 0.01543f
C8820 XThR.Tn[9].t69 VGND 0.01689f
C8821 XThR.Tn[9].n73 VGND 0.04125f
C8822 XThR.Tn[9].t30 VGND 0.01538f
C8823 XThR.Tn[9].t61 VGND 0.01684f
C8824 XThR.Tn[9].n74 VGND 0.04292f
C8825 XThR.Tn[9].n75 VGND 0.03015f
C8826 XThR.Tn[9].n77 VGND 0.09677f
C8827 XThR.Tn[9].t49 VGND 0.01543f
C8828 XThR.Tn[9].t63 VGND 0.01689f
C8829 XThR.Tn[9].n78 VGND 0.04125f
C8830 XThR.Tn[9].t68 VGND 0.01538f
C8831 XThR.Tn[9].t54 VGND 0.01684f
C8832 XThR.Tn[9].n79 VGND 0.04292f
C8833 XThR.Tn[9].n80 VGND 0.03015f
C8834 XThR.Tn[9].n82 VGND 0.09677f
C8835 XThR.Tn[9].n83 VGND 0.08794f
C8836 XThR.Tn[9].n84 VGND 0.28527f
C8837 XThR.Tn[9].t2 VGND 0.01974f
C8838 XThR.Tn[9].t0 VGND 0.01974f
C8839 XThR.Tn[9].n85 VGND 0.04265f
C8840 XThR.Tn[9].t3 VGND 0.01974f
C8841 XThR.Tn[9].t1 VGND 0.01974f
C8842 XThR.Tn[9].n86 VGND 0.06492f
C8843 XThR.Tn[9].n87 VGND 0.18025f
C8844 XThR.Tn[9].n88 VGND 0.02413f
C8845 XThC.Tn[6].t7 VGND 0.0146f
C8846 XThC.Tn[6].t6 VGND 0.0146f
C8847 XThC.Tn[6].n0 VGND 0.02948f
C8848 XThC.Tn[6].t5 VGND 0.0146f
C8849 XThC.Tn[6].t4 VGND 0.0146f
C8850 XThC.Tn[6].n1 VGND 0.03449f
C8851 XThC.Tn[6].n2 VGND 0.09656f
C8852 XThC.Tn[6].n3 VGND 0.03602f
C8853 XThC.Tn[6].n4 VGND 0.02162f
C8854 XThC.Tn[6].n5 VGND 0.10295f
C8855 XThC.Tn[6].n6 VGND 0.02162f
C8856 XThC.Tn[6].n7 VGND 0.06364f
C8857 XThC.Tn[6].n8 VGND 0.02162f
C8858 XThC.Tn[6].n9 VGND 0.07182f
C8859 XThC.Tn[6].t23 VGND 0.01158f
C8860 XThC.Tn[6].t26 VGND 0.01264f
C8861 XThC.Tn[6].n10 VGND 0.02823f
C8862 XThC.Tn[6].n11 VGND 0.01934f
C8863 XThC.Tn[6].n12 VGND 0.06347f
C8864 XThC.Tn[6].t40 VGND 0.01158f
C8865 XThC.Tn[6].t13 VGND 0.01264f
C8866 XThC.Tn[6].n13 VGND 0.02823f
C8867 XThC.Tn[6].n14 VGND 0.01934f
C8868 XThC.Tn[6].n15 VGND 0.06365f
C8869 XThC.Tn[6].n16 VGND 0.1049f
C8870 XThC.Tn[6].t42 VGND 0.01158f
C8871 XThC.Tn[6].t17 VGND 0.01264f
C8872 XThC.Tn[6].n17 VGND 0.02823f
C8873 XThC.Tn[6].n18 VGND 0.01934f
C8874 XThC.Tn[6].n19 VGND 0.06365f
C8875 XThC.Tn[6].n20 VGND 0.1049f
C8876 XThC.Tn[6].t12 VGND 0.01158f
C8877 XThC.Tn[6].t18 VGND 0.01264f
C8878 XThC.Tn[6].n21 VGND 0.02823f
C8879 XThC.Tn[6].n22 VGND 0.01934f
C8880 XThC.Tn[6].n23 VGND 0.06365f
C8881 XThC.Tn[6].n24 VGND 0.1049f
C8882 XThC.Tn[6].t33 VGND 0.01158f
C8883 XThC.Tn[6].t37 VGND 0.01264f
C8884 XThC.Tn[6].n25 VGND 0.02823f
C8885 XThC.Tn[6].n26 VGND 0.01934f
C8886 XThC.Tn[6].n27 VGND 0.06365f
C8887 XThC.Tn[6].n28 VGND 0.1049f
C8888 XThC.Tn[6].t35 VGND 0.01158f
C8889 XThC.Tn[6].t38 VGND 0.01264f
C8890 XThC.Tn[6].n29 VGND 0.02823f
C8891 XThC.Tn[6].n30 VGND 0.01934f
C8892 XThC.Tn[6].n31 VGND 0.06365f
C8893 XThC.Tn[6].n32 VGND 0.1049f
C8894 XThC.Tn[6].t16 VGND 0.01158f
C8895 XThC.Tn[6].t22 VGND 0.01264f
C8896 XThC.Tn[6].n33 VGND 0.02823f
C8897 XThC.Tn[6].n34 VGND 0.01934f
C8898 XThC.Tn[6].n35 VGND 0.06365f
C8899 XThC.Tn[6].n36 VGND 0.1049f
C8900 XThC.Tn[6].t25 VGND 0.01158f
C8901 XThC.Tn[6].t29 VGND 0.01264f
C8902 XThC.Tn[6].n37 VGND 0.02823f
C8903 XThC.Tn[6].n38 VGND 0.01934f
C8904 XThC.Tn[6].n39 VGND 0.06365f
C8905 XThC.Tn[6].n40 VGND 0.1049f
C8906 XThC.Tn[6].t27 VGND 0.01158f
C8907 XThC.Tn[6].t31 VGND 0.01264f
C8908 XThC.Tn[6].n41 VGND 0.02823f
C8909 XThC.Tn[6].n42 VGND 0.01934f
C8910 XThC.Tn[6].n43 VGND 0.06365f
C8911 XThC.Tn[6].n44 VGND 0.1049f
C8912 XThC.Tn[6].t14 VGND 0.01158f
C8913 XThC.Tn[6].t19 VGND 0.01264f
C8914 XThC.Tn[6].n45 VGND 0.02823f
C8915 XThC.Tn[6].n46 VGND 0.01934f
C8916 XThC.Tn[6].n47 VGND 0.06365f
C8917 XThC.Tn[6].n48 VGND 0.1049f
C8918 XThC.Tn[6].t15 VGND 0.01158f
C8919 XThC.Tn[6].t21 VGND 0.01264f
C8920 XThC.Tn[6].n49 VGND 0.02823f
C8921 XThC.Tn[6].n50 VGND 0.01934f
C8922 XThC.Tn[6].n51 VGND 0.06365f
C8923 XThC.Tn[6].n52 VGND 0.1049f
C8924 XThC.Tn[6].t28 VGND 0.01158f
C8925 XThC.Tn[6].t32 VGND 0.01264f
C8926 XThC.Tn[6].n53 VGND 0.02823f
C8927 XThC.Tn[6].n54 VGND 0.01934f
C8928 XThC.Tn[6].n55 VGND 0.06365f
C8929 XThC.Tn[6].n56 VGND 0.1049f
C8930 XThC.Tn[6].t36 VGND 0.01158f
C8931 XThC.Tn[6].t41 VGND 0.01264f
C8932 XThC.Tn[6].n57 VGND 0.02823f
C8933 XThC.Tn[6].n58 VGND 0.01934f
C8934 XThC.Tn[6].n59 VGND 0.06365f
C8935 XThC.Tn[6].n60 VGND 0.1049f
C8936 XThC.Tn[6].t39 VGND 0.01158f
C8937 XThC.Tn[6].t43 VGND 0.01264f
C8938 XThC.Tn[6].n61 VGND 0.02823f
C8939 XThC.Tn[6].n62 VGND 0.01934f
C8940 XThC.Tn[6].n63 VGND 0.06365f
C8941 XThC.Tn[6].n64 VGND 0.1049f
C8942 XThC.Tn[6].t20 VGND 0.01158f
C8943 XThC.Tn[6].t24 VGND 0.01264f
C8944 XThC.Tn[6].n65 VGND 0.02823f
C8945 XThC.Tn[6].n66 VGND 0.01934f
C8946 XThC.Tn[6].n67 VGND 0.06365f
C8947 XThC.Tn[6].n68 VGND 0.1049f
C8948 XThC.Tn[6].t30 VGND 0.01158f
C8949 XThC.Tn[6].t34 VGND 0.01264f
C8950 XThC.Tn[6].n69 VGND 0.02823f
C8951 XThC.Tn[6].n70 VGND 0.01934f
C8952 XThC.Tn[6].n71 VGND 0.06365f
C8953 XThC.Tn[6].n72 VGND 0.1049f
C8954 XThC.Tn[6].n73 VGND 0.11666f
C8955 XThC.Tn[6].n74 VGND 0.03056f
C8956 XThC.XTBN.Y.n0 VGND 0.01531f
C8957 XThC.XTBN.Y.t50 VGND 0.01024f
C8958 XThC.XTBN.Y.t18 VGND 0.01024f
C8959 XThC.XTBN.Y.n1 VGND 0.01477f
C8960 XThC.XTBN.Y.t120 VGND 0.01024f
C8961 XThC.XTBN.Y.t114 VGND 0.01024f
C8962 XThC.XTBN.Y.n3 VGND 0.0138f
C8963 XThC.XTBN.Y.n5 VGND 0.01477f
C8964 XThC.XTBN.Y.n10 VGND 0.02164f
C8965 XThC.XTBN.Y.t79 VGND 0.01024f
C8966 XThC.XTBN.Y.t36 VGND 0.01024f
C8967 XThC.XTBN.Y.n13 VGND 0.01477f
C8968 XThC.XTBN.Y.t26 VGND 0.01024f
C8969 XThC.XTBN.Y.t21 VGND 0.01024f
C8970 XThC.XTBN.Y.n15 VGND 0.0138f
C8971 XThC.XTBN.Y.n17 VGND 0.01477f
C8972 XThC.XTBN.Y.n22 VGND 0.02164f
C8973 XThC.XTBN.Y.n25 VGND 0.11789f
C8974 XThC.XTBN.Y.t106 VGND 0.01024f
C8975 XThC.XTBN.Y.t70 VGND 0.01024f
C8976 XThC.XTBN.Y.n26 VGND 0.01477f
C8977 XThC.XTBN.Y.t56 VGND 0.01024f
C8978 XThC.XTBN.Y.t48 VGND 0.01024f
C8979 XThC.XTBN.Y.n28 VGND 0.0138f
C8980 XThC.XTBN.Y.n30 VGND 0.01477f
C8981 XThC.XTBN.Y.n35 VGND 0.02164f
C8982 XThC.XTBN.Y.n38 VGND 0.07443f
C8983 XThC.XTBN.Y.t39 VGND 0.01024f
C8984 XThC.XTBN.Y.t122 VGND 0.01024f
C8985 XThC.XTBN.Y.n39 VGND 0.01477f
C8986 XThC.XTBN.Y.t109 VGND 0.01024f
C8987 XThC.XTBN.Y.t102 VGND 0.01024f
C8988 XThC.XTBN.Y.n41 VGND 0.0138f
C8989 XThC.XTBN.Y.n43 VGND 0.01477f
C8990 XThC.XTBN.Y.n48 VGND 0.02164f
C8991 XThC.XTBN.Y.n51 VGND 0.07443f
C8992 XThC.XTBN.Y.t47 VGND 0.01024f
C8993 XThC.XTBN.Y.t17 VGND 0.01024f
C8994 XThC.XTBN.Y.n52 VGND 0.01477f
C8995 XThC.XTBN.Y.t116 VGND 0.01024f
C8996 XThC.XTBN.Y.t111 VGND 0.01024f
C8997 XThC.XTBN.Y.n54 VGND 0.0138f
C8998 XThC.XTBN.Y.n56 VGND 0.01477f
C8999 XThC.XTBN.Y.n61 VGND 0.02164f
C9000 XThC.XTBN.Y.n64 VGND 0.07443f
C9001 XThC.XTBN.Y.t101 VGND 0.01024f
C9002 XThC.XTBN.Y.t63 VGND 0.01024f
C9003 XThC.XTBN.Y.n65 VGND 0.01477f
C9004 XThC.XTBN.Y.t52 VGND 0.01024f
C9005 XThC.XTBN.Y.t44 VGND 0.01024f
C9006 XThC.XTBN.Y.n67 VGND 0.0138f
C9007 XThC.XTBN.Y.n69 VGND 0.01477f
C9008 XThC.XTBN.Y.n74 VGND 0.02164f
C9009 XThC.XTBN.Y.n77 VGND 0.07443f
C9010 XThC.XTBN.Y.t25 VGND 0.01024f
C9011 XThC.XTBN.Y.t100 VGND 0.01024f
C9012 XThC.XTBN.Y.n78 VGND 0.01477f
C9013 XThC.XTBN.Y.t93 VGND 0.01024f
C9014 XThC.XTBN.Y.t90 VGND 0.01024f
C9015 XThC.XTBN.Y.n80 VGND 0.0138f
C9016 XThC.XTBN.Y.n82 VGND 0.01477f
C9017 XThC.XTBN.Y.n87 VGND 0.02164f
C9018 XThC.XTBN.Y.n90 VGND 0.06646f
C9019 XThC.XTBN.Y.t46 VGND 0.01024f
C9020 XThC.XTBN.Y.t6 VGND 0.01024f
C9021 XThC.XTBN.Y.n92 VGND 0.01243f
C9022 XThC.XTBN.Y.t12 VGND 0.01024f
C9023 XThC.XTBN.Y.n93 VGND 0.01348f
C9024 XThC.XTBN.Y.n95 VGND 0.01252f
C9025 XThC.XTBN.Y.n98 VGND 0.01348f
C9026 XThC.XTBN.Y.t54 VGND 0.01024f
C9027 XThC.XTBN.Y.n99 VGND 0.01227f
C9028 XThC.XTBN.Y.n101 VGND 0.01009f
C9029 XThC.XTBN.Y.t38 VGND 0.01024f
C9030 XThC.XTBN.Y.t113 VGND 0.01024f
C9031 XThC.XTBN.Y.n103 VGND 0.01243f
C9032 XThC.XTBN.Y.t119 VGND 0.01024f
C9033 XThC.XTBN.Y.n104 VGND 0.01348f
C9034 XThC.XTBN.Y.n106 VGND 0.01252f
C9035 XThC.XTBN.Y.n109 VGND 0.01348f
C9036 XThC.XTBN.Y.t42 VGND 0.01024f
C9037 XThC.XTBN.Y.n110 VGND 0.01227f
C9038 XThC.XTBN.Y.n113 VGND 0.11256f
C9039 XThC.XTBN.Y.t30 VGND 0.01024f
C9040 XThC.XTBN.Y.t98 VGND 0.01024f
C9041 XThC.XTBN.Y.n115 VGND 0.01243f
C9042 XThC.XTBN.Y.t103 VGND 0.01024f
C9043 XThC.XTBN.Y.n116 VGND 0.01348f
C9044 XThC.XTBN.Y.n118 VGND 0.01252f
C9045 XThC.XTBN.Y.n121 VGND 0.01348f
C9046 XThC.XTBN.Y.t34 VGND 0.01024f
C9047 XThC.XTBN.Y.n122 VGND 0.01227f
C9048 XThC.XTBN.Y.n125 VGND 0.07521f
C9049 XThC.XTBN.Y.t96 VGND 0.01024f
C9050 XThC.XTBN.Y.t51 VGND 0.01024f
C9051 XThC.XTBN.Y.n127 VGND 0.01243f
C9052 XThC.XTBN.Y.t58 VGND 0.01024f
C9053 XThC.XTBN.Y.n128 VGND 0.01348f
C9054 XThC.XTBN.Y.n130 VGND 0.01252f
C9055 XThC.XTBN.Y.n133 VGND 0.01348f
C9056 XThC.XTBN.Y.t99 VGND 0.01024f
C9057 XThC.XTBN.Y.n134 VGND 0.01227f
C9058 XThC.XTBN.Y.n137 VGND 0.07521f
C9059 XThC.XTBN.Y.t88 VGND 0.01024f
C9060 XThC.XTBN.Y.t37 VGND 0.01024f
C9061 XThC.XTBN.Y.n139 VGND 0.01243f
C9062 XThC.XTBN.Y.t40 VGND 0.01024f
C9063 XThC.XTBN.Y.n140 VGND 0.01348f
C9064 XThC.XTBN.Y.n142 VGND 0.01252f
C9065 XThC.XTBN.Y.n145 VGND 0.01348f
C9066 XThC.XTBN.Y.t91 VGND 0.01024f
C9067 XThC.XTBN.Y.n146 VGND 0.01227f
C9068 XThC.XTBN.Y.n149 VGND 0.07534f
C9069 XThC.XTBN.Y.t7 VGND 0.01024f
C9070 XThC.XTBN.Y.t81 VGND 0.01024f
C9071 XThC.XTBN.Y.n151 VGND 0.01243f
C9072 XThC.XTBN.Y.t86 VGND 0.01024f
C9073 XThC.XTBN.Y.n152 VGND 0.01348f
C9074 XThC.XTBN.Y.n154 VGND 0.01252f
C9075 XThC.XTBN.Y.n157 VGND 0.01348f
C9076 XThC.XTBN.Y.t13 VGND 0.01024f
C9077 XThC.XTBN.Y.n158 VGND 0.01227f
C9078 XThC.XTBN.Y.n161 VGND 0.07521f
C9079 XThC.XTBN.Y.t23 VGND 0.01024f
C9080 XThC.XTBN.Y.t95 VGND 0.01024f
C9081 XThC.XTBN.Y.n163 VGND 0.01243f
C9082 XThC.XTBN.Y.t97 VGND 0.01024f
C9083 XThC.XTBN.Y.n164 VGND 0.01348f
C9084 XThC.XTBN.Y.n166 VGND 0.01252f
C9085 XThC.XTBN.Y.n169 VGND 0.01348f
C9086 XThC.XTBN.Y.t28 VGND 0.01024f
C9087 XThC.XTBN.Y.n170 VGND 0.01227f
C9088 XThC.XTBN.Y.n173 VGND 0.08751f
C9089 XThC.XTBN.Y.n174 VGND 0.11019f
C9090 XThC.XTBN.Y.t75 VGND 0.01024f
C9091 XThC.XTBN.Y.t33 VGND 0.01024f
C9092 XThC.XTBN.Y.n175 VGND 0.01477f
C9093 XThC.XTBN.Y.t27 VGND 0.01024f
C9094 XThC.XTBN.Y.n176 VGND 0.02293f
C9095 XThC.XTBN.Y.n181 VGND 0.01477f
C9096 XThC.XTBN.Y.t9 VGND 0.01024f
C9097 XThC.XTBN.Y.n182 VGND 0.0138f
C9098 XThC.XTBN.Y.n186 VGND 0.11129f
C9099 XThC.XTBN.Y.n187 VGND 0.02169f
C9100 XThC.XTBN.Y.n191 VGND 0.01513f
C9101 XThC.XTBN.Y.n192 VGND 0.0307f
C9102 XThR.Tn[12].t11 VGND 0.01974f
C9103 XThR.Tn[12].t9 VGND 0.01974f
C9104 XThR.Tn[12].n0 VGND 0.05994f
C9105 XThR.Tn[12].t8 VGND 0.01974f
C9106 XThR.Tn[12].t10 VGND 0.01974f
C9107 XThR.Tn[12].n1 VGND 0.04388f
C9108 XThR.Tn[12].n2 VGND 0.19954f
C9109 XThR.Tn[12].t7 VGND 0.01283f
C9110 XThR.Tn[12].t5 VGND 0.01283f
C9111 XThR.Tn[12].n3 VGND 0.032f
C9112 XThR.Tn[12].t6 VGND 0.01283f
C9113 XThR.Tn[12].t4 VGND 0.01283f
C9114 XThR.Tn[12].n4 VGND 0.02566f
C9115 XThR.Tn[12].n5 VGND 0.05917f
C9116 XThR.Tn[12].t36 VGND 0.01543f
C9117 XThR.Tn[12].t28 VGND 0.01689f
C9118 XThR.Tn[12].n6 VGND 0.04125f
C9119 XThR.Tn[12].n7 VGND 0.07925f
C9120 XThR.Tn[12].t53 VGND 0.01543f
C9121 XThR.Tn[12].t43 VGND 0.01689f
C9122 XThR.Tn[12].n8 VGND 0.04125f
C9123 XThR.Tn[12].t71 VGND 0.01538f
C9124 XThR.Tn[12].t21 VGND 0.01684f
C9125 XThR.Tn[12].n9 VGND 0.04292f
C9126 XThR.Tn[12].n10 VGND 0.03016f
C9127 XThR.Tn[12].n12 VGND 0.09677f
C9128 XThR.Tn[12].t30 VGND 0.01543f
C9129 XThR.Tn[12].t20 VGND 0.01689f
C9130 XThR.Tn[12].n13 VGND 0.04125f
C9131 XThR.Tn[12].t49 VGND 0.01538f
C9132 XThR.Tn[12].t60 VGND 0.01684f
C9133 XThR.Tn[12].n14 VGND 0.04292f
C9134 XThR.Tn[12].n15 VGND 0.03016f
C9135 XThR.Tn[12].n17 VGND 0.09677f
C9136 XThR.Tn[12].t45 VGND 0.01543f
C9137 XThR.Tn[12].t38 VGND 0.01689f
C9138 XThR.Tn[12].n18 VGND 0.04125f
C9139 XThR.Tn[12].t63 VGND 0.01538f
C9140 XThR.Tn[12].t15 VGND 0.01684f
C9141 XThR.Tn[12].n19 VGND 0.04292f
C9142 XThR.Tn[12].n20 VGND 0.03016f
C9143 XThR.Tn[12].n22 VGND 0.09677f
C9144 XThR.Tn[12].t70 VGND 0.01543f
C9145 XThR.Tn[12].t66 VGND 0.01689f
C9146 XThR.Tn[12].n23 VGND 0.04125f
C9147 XThR.Tn[12].t33 VGND 0.01538f
C9148 XThR.Tn[12].t46 VGND 0.01684f
C9149 XThR.Tn[12].n24 VGND 0.04292f
C9150 XThR.Tn[12].n25 VGND 0.03016f
C9151 XThR.Tn[12].n27 VGND 0.09677f
C9152 XThR.Tn[12].t48 VGND 0.01543f
C9153 XThR.Tn[12].t39 VGND 0.01689f
C9154 XThR.Tn[12].n28 VGND 0.04125f
C9155 XThR.Tn[12].t64 VGND 0.01538f
C9156 XThR.Tn[12].t17 VGND 0.01684f
C9157 XThR.Tn[12].n29 VGND 0.04292f
C9158 XThR.Tn[12].n30 VGND 0.03016f
C9159 XThR.Tn[12].n32 VGND 0.09677f
C9160 XThR.Tn[12].t23 VGND 0.01543f
C9161 XThR.Tn[12].t56 VGND 0.01689f
C9162 XThR.Tn[12].n33 VGND 0.04125f
C9163 XThR.Tn[12].t41 VGND 0.01538f
C9164 XThR.Tn[12].t37 VGND 0.01684f
C9165 XThR.Tn[12].n34 VGND 0.04292f
C9166 XThR.Tn[12].n35 VGND 0.03016f
C9167 XThR.Tn[12].n37 VGND 0.09677f
C9168 XThR.Tn[12].t54 VGND 0.01543f
C9169 XThR.Tn[12].t51 VGND 0.01689f
C9170 XThR.Tn[12].n38 VGND 0.04125f
C9171 XThR.Tn[12].t72 VGND 0.01538f
C9172 XThR.Tn[12].t29 VGND 0.01684f
C9173 XThR.Tn[12].n39 VGND 0.04292f
C9174 XThR.Tn[12].n40 VGND 0.03016f
C9175 XThR.Tn[12].n42 VGND 0.09677f
C9176 XThR.Tn[12].t59 VGND 0.01543f
C9177 XThR.Tn[12].t65 VGND 0.01689f
C9178 XThR.Tn[12].n43 VGND 0.04125f
C9179 XThR.Tn[12].t14 VGND 0.01538f
C9180 XThR.Tn[12].t44 VGND 0.01684f
C9181 XThR.Tn[12].n44 VGND 0.04292f
C9182 XThR.Tn[12].n45 VGND 0.03016f
C9183 XThR.Tn[12].n47 VGND 0.09677f
C9184 XThR.Tn[12].t12 VGND 0.01543f
C9185 XThR.Tn[12].t22 VGND 0.01689f
C9186 XThR.Tn[12].n48 VGND 0.04125f
C9187 XThR.Tn[12].t35 VGND 0.01538f
C9188 XThR.Tn[12].t61 VGND 0.01684f
C9189 XThR.Tn[12].n49 VGND 0.04292f
C9190 XThR.Tn[12].n50 VGND 0.03016f
C9191 XThR.Tn[12].n52 VGND 0.09677f
C9192 XThR.Tn[12].t68 VGND 0.01543f
C9193 XThR.Tn[12].t40 VGND 0.01689f
C9194 XThR.Tn[12].n53 VGND 0.04125f
C9195 XThR.Tn[12].t26 VGND 0.01538f
C9196 XThR.Tn[12].t19 VGND 0.01684f
C9197 XThR.Tn[12].n54 VGND 0.04292f
C9198 XThR.Tn[12].n55 VGND 0.03016f
C9199 XThR.Tn[12].n57 VGND 0.09677f
C9200 XThR.Tn[12].t25 VGND 0.01543f
C9201 XThR.Tn[12].t16 VGND 0.01689f
C9202 XThR.Tn[12].n58 VGND 0.04125f
C9203 XThR.Tn[12].t42 VGND 0.01538f
C9204 XThR.Tn[12].t55 VGND 0.01684f
C9205 XThR.Tn[12].n59 VGND 0.04292f
C9206 XThR.Tn[12].n60 VGND 0.03016f
C9207 XThR.Tn[12].n62 VGND 0.09677f
C9208 XThR.Tn[12].t57 VGND 0.01543f
C9209 XThR.Tn[12].t52 VGND 0.01689f
C9210 XThR.Tn[12].n63 VGND 0.04125f
C9211 XThR.Tn[12].t13 VGND 0.01538f
C9212 XThR.Tn[12].t31 VGND 0.01684f
C9213 XThR.Tn[12].n64 VGND 0.04292f
C9214 XThR.Tn[12].n65 VGND 0.03016f
C9215 XThR.Tn[12].n67 VGND 0.09677f
C9216 XThR.Tn[12].t73 VGND 0.01543f
C9217 XThR.Tn[12].t67 VGND 0.01689f
C9218 XThR.Tn[12].n68 VGND 0.04125f
C9219 XThR.Tn[12].t34 VGND 0.01538f
C9220 XThR.Tn[12].t47 VGND 0.01684f
C9221 XThR.Tn[12].n69 VGND 0.04292f
C9222 XThR.Tn[12].n70 VGND 0.03016f
C9223 XThR.Tn[12].n72 VGND 0.09677f
C9224 XThR.Tn[12].t32 VGND 0.01543f
C9225 XThR.Tn[12].t24 VGND 0.01689f
C9226 XThR.Tn[12].n73 VGND 0.04125f
C9227 XThR.Tn[12].t50 VGND 0.01538f
C9228 XThR.Tn[12].t62 VGND 0.01684f
C9229 XThR.Tn[12].n74 VGND 0.04292f
C9230 XThR.Tn[12].n75 VGND 0.03016f
C9231 XThR.Tn[12].n77 VGND 0.09677f
C9232 XThR.Tn[12].t69 VGND 0.01543f
C9233 XThR.Tn[12].t18 VGND 0.01689f
C9234 XThR.Tn[12].n78 VGND 0.04125f
C9235 XThR.Tn[12].t27 VGND 0.01538f
C9236 XThR.Tn[12].t58 VGND 0.01684f
C9237 XThR.Tn[12].n79 VGND 0.04292f
C9238 XThR.Tn[12].n80 VGND 0.03016f
C9239 XThR.Tn[12].n82 VGND 0.09677f
C9240 XThR.Tn[12].n83 VGND 0.08794f
C9241 XThR.Tn[12].n84 VGND 0.29993f
C9242 XThR.Tn[12].t2 VGND 0.01974f
C9243 XThR.Tn[12].t0 VGND 0.01974f
C9244 XThR.Tn[12].n85 VGND 0.04265f
C9245 XThR.Tn[12].t3 VGND 0.01974f
C9246 XThR.Tn[12].t1 VGND 0.01974f
C9247 XThR.Tn[12].n86 VGND 0.06492f
C9248 XThR.Tn[12].n87 VGND 0.18025f
C9249 XThR.Tn[14].t8 VGND 0.02012f
C9250 XThR.Tn[14].t9 VGND 0.02012f
C9251 XThR.Tn[14].n0 VGND 0.06109f
C9252 XThR.Tn[14].t10 VGND 0.02012f
C9253 XThR.Tn[14].t11 VGND 0.02012f
C9254 XThR.Tn[14].n1 VGND 0.04473f
C9255 XThR.Tn[14].n2 VGND 0.20337f
C9256 XThR.Tn[14].t6 VGND 0.01308f
C9257 XThR.Tn[14].t7 VGND 0.01308f
C9258 XThR.Tn[14].n3 VGND 0.03262f
C9259 XThR.Tn[14].t4 VGND 0.01308f
C9260 XThR.Tn[14].t5 VGND 0.01308f
C9261 XThR.Tn[14].n4 VGND 0.02616f
C9262 XThR.Tn[14].n5 VGND 0.06031f
C9263 XThR.Tn[14].t69 VGND 0.01572f
C9264 XThR.Tn[14].t62 VGND 0.01722f
C9265 XThR.Tn[14].n6 VGND 0.04205f
C9266 XThR.Tn[14].n7 VGND 0.08077f
C9267 XThR.Tn[14].t24 VGND 0.01572f
C9268 XThR.Tn[14].t13 VGND 0.01722f
C9269 XThR.Tn[14].n8 VGND 0.04205f
C9270 XThR.Tn[14].t28 VGND 0.01567f
C9271 XThR.Tn[14].t60 VGND 0.01716f
C9272 XThR.Tn[14].n9 VGND 0.04375f
C9273 XThR.Tn[14].n10 VGND 0.03073f
C9274 XThR.Tn[14].n12 VGND 0.09863f
C9275 XThR.Tn[14].t64 VGND 0.01572f
C9276 XThR.Tn[14].t54 VGND 0.01722f
C9277 XThR.Tn[14].n13 VGND 0.04205f
C9278 XThR.Tn[14].t67 VGND 0.01567f
C9279 XThR.Tn[14].t34 VGND 0.01716f
C9280 XThR.Tn[14].n14 VGND 0.04375f
C9281 XThR.Tn[14].n15 VGND 0.03073f
C9282 XThR.Tn[14].n17 VGND 0.09863f
C9283 XThR.Tn[14].t14 VGND 0.01572f
C9284 XThR.Tn[14].t72 VGND 0.01722f
C9285 XThR.Tn[14].n18 VGND 0.04205f
C9286 XThR.Tn[14].t17 VGND 0.01567f
C9287 XThR.Tn[14].t52 VGND 0.01716f
C9288 XThR.Tn[14].n19 VGND 0.04375f
C9289 XThR.Tn[14].n20 VGND 0.03073f
C9290 XThR.Tn[14].n22 VGND 0.09863f
C9291 XThR.Tn[14].t44 VGND 0.01572f
C9292 XThR.Tn[14].t38 VGND 0.01722f
C9293 XThR.Tn[14].n23 VGND 0.04205f
C9294 XThR.Tn[14].t47 VGND 0.01567f
C9295 XThR.Tn[14].t18 VGND 0.01716f
C9296 XThR.Tn[14].n24 VGND 0.04375f
C9297 XThR.Tn[14].n25 VGND 0.03073f
C9298 XThR.Tn[14].n27 VGND 0.09863f
C9299 XThR.Tn[14].t15 VGND 0.01572f
C9300 XThR.Tn[14].t73 VGND 0.01722f
C9301 XThR.Tn[14].n28 VGND 0.04205f
C9302 XThR.Tn[14].t21 VGND 0.01567f
C9303 XThR.Tn[14].t53 VGND 0.01716f
C9304 XThR.Tn[14].n29 VGND 0.04375f
C9305 XThR.Tn[14].n30 VGND 0.03073f
C9306 XThR.Tn[14].n32 VGND 0.09863f
C9307 XThR.Tn[14].t57 VGND 0.01572f
C9308 XThR.Tn[14].t25 VGND 0.01722f
C9309 XThR.Tn[14].n33 VGND 0.04205f
C9310 XThR.Tn[14].t61 VGND 0.01567f
C9311 XThR.Tn[14].t71 VGND 0.01716f
C9312 XThR.Tn[14].n34 VGND 0.04375f
C9313 XThR.Tn[14].n35 VGND 0.03073f
C9314 XThR.Tn[14].n37 VGND 0.09863f
C9315 XThR.Tn[14].t23 VGND 0.01572f
C9316 XThR.Tn[14].t19 VGND 0.01722f
C9317 XThR.Tn[14].n38 VGND 0.04205f
C9318 XThR.Tn[14].t29 VGND 0.01567f
C9319 XThR.Tn[14].t66 VGND 0.01716f
C9320 XThR.Tn[14].n39 VGND 0.04375f
C9321 XThR.Tn[14].n40 VGND 0.03073f
C9322 XThR.Tn[14].n42 VGND 0.09863f
C9323 XThR.Tn[14].t27 VGND 0.01572f
C9324 XThR.Tn[14].t36 VGND 0.01722f
C9325 XThR.Tn[14].n43 VGND 0.04205f
C9326 XThR.Tn[14].t33 VGND 0.01567f
C9327 XThR.Tn[14].t16 VGND 0.01716f
C9328 XThR.Tn[14].n44 VGND 0.04375f
C9329 XThR.Tn[14].n45 VGND 0.03073f
C9330 XThR.Tn[14].n47 VGND 0.09863f
C9331 XThR.Tn[14].t46 VGND 0.01572f
C9332 XThR.Tn[14].t56 VGND 0.01722f
C9333 XThR.Tn[14].n48 VGND 0.04205f
C9334 XThR.Tn[14].t50 VGND 0.01567f
C9335 XThR.Tn[14].t35 VGND 0.01716f
C9336 XThR.Tn[14].n49 VGND 0.04375f
C9337 XThR.Tn[14].n50 VGND 0.03073f
C9338 XThR.Tn[14].n52 VGND 0.09863f
C9339 XThR.Tn[14].t40 VGND 0.01572f
C9340 XThR.Tn[14].t12 VGND 0.01722f
C9341 XThR.Tn[14].n53 VGND 0.04205f
C9342 XThR.Tn[14].t42 VGND 0.01567f
C9343 XThR.Tn[14].t55 VGND 0.01716f
C9344 XThR.Tn[14].n54 VGND 0.04375f
C9345 XThR.Tn[14].n55 VGND 0.03073f
C9346 XThR.Tn[14].n57 VGND 0.09863f
C9347 XThR.Tn[14].t59 VGND 0.01572f
C9348 XThR.Tn[14].t49 VGND 0.01722f
C9349 XThR.Tn[14].n58 VGND 0.04205f
C9350 XThR.Tn[14].t63 VGND 0.01567f
C9351 XThR.Tn[14].t30 VGND 0.01716f
C9352 XThR.Tn[14].n59 VGND 0.04375f
C9353 XThR.Tn[14].n60 VGND 0.03073f
C9354 XThR.Tn[14].n62 VGND 0.09863f
C9355 XThR.Tn[14].t26 VGND 0.01572f
C9356 XThR.Tn[14].t22 VGND 0.01722f
C9357 XThR.Tn[14].n63 VGND 0.04205f
C9358 XThR.Tn[14].t31 VGND 0.01567f
C9359 XThR.Tn[14].t68 VGND 0.01716f
C9360 XThR.Tn[14].n64 VGND 0.04375f
C9361 XThR.Tn[14].n65 VGND 0.03073f
C9362 XThR.Tn[14].n67 VGND 0.09863f
C9363 XThR.Tn[14].t45 VGND 0.01572f
C9364 XThR.Tn[14].t39 VGND 0.01722f
C9365 XThR.Tn[14].n68 VGND 0.04205f
C9366 XThR.Tn[14].t48 VGND 0.01567f
C9367 XThR.Tn[14].t20 VGND 0.01716f
C9368 XThR.Tn[14].n69 VGND 0.04375f
C9369 XThR.Tn[14].n70 VGND 0.03073f
C9370 XThR.Tn[14].n72 VGND 0.09863f
C9371 XThR.Tn[14].t65 VGND 0.01572f
C9372 XThR.Tn[14].t58 VGND 0.01722f
C9373 XThR.Tn[14].n73 VGND 0.04205f
C9374 XThR.Tn[14].t70 VGND 0.01567f
C9375 XThR.Tn[14].t37 VGND 0.01716f
C9376 XThR.Tn[14].n74 VGND 0.04375f
C9377 XThR.Tn[14].n75 VGND 0.03073f
C9378 XThR.Tn[14].n77 VGND 0.09863f
C9379 XThR.Tn[14].t41 VGND 0.01572f
C9380 XThR.Tn[14].t51 VGND 0.01722f
C9381 XThR.Tn[14].n78 VGND 0.04205f
C9382 XThR.Tn[14].t43 VGND 0.01567f
C9383 XThR.Tn[14].t32 VGND 0.01716f
C9384 XThR.Tn[14].n79 VGND 0.04375f
C9385 XThR.Tn[14].n80 VGND 0.03073f
C9386 XThR.Tn[14].n82 VGND 0.09863f
C9387 XThR.Tn[14].n83 VGND 0.08963f
C9388 XThR.Tn[14].n84 VGND 0.36005f
C9389 XThR.Tn[14].t2 VGND 0.02012f
C9390 XThR.Tn[14].t3 VGND 0.02012f
C9391 XThR.Tn[14].n85 VGND 0.04347f
C9392 XThR.Tn[14].t0 VGND 0.02012f
C9393 XThR.Tn[14].t1 VGND 0.02012f
C9394 XThR.Tn[14].n86 VGND 0.06616f
C9395 XThR.Tn[14].n87 VGND 0.18371f
C9396 XThR.Tn[6].t7 VGND 0.01859f
C9397 XThR.Tn[6].t4 VGND 0.01859f
C9398 XThR.Tn[6].n0 VGND 0.03751f
C9399 XThR.Tn[6].t6 VGND 0.01859f
C9400 XThR.Tn[6].t5 VGND 0.01859f
C9401 XThR.Tn[6].n1 VGND 0.04389f
C9402 XThR.Tn[6].n2 VGND 0.13166f
C9403 XThR.Tn[6].t8 VGND 0.01208f
C9404 XThR.Tn[6].t9 VGND 0.01208f
C9405 XThR.Tn[6].n3 VGND 0.02751f
C9406 XThR.Tn[6].t11 VGND 0.01208f
C9407 XThR.Tn[6].t10 VGND 0.01208f
C9408 XThR.Tn[6].n4 VGND 0.02751f
C9409 XThR.Tn[6].t0 VGND 0.01208f
C9410 XThR.Tn[6].t1 VGND 0.01208f
C9411 XThR.Tn[6].n5 VGND 0.04584f
C9412 XThR.Tn[6].t3 VGND 0.01208f
C9413 XThR.Tn[6].t2 VGND 0.01208f
C9414 XThR.Tn[6].n6 VGND 0.02751f
C9415 XThR.Tn[6].n7 VGND 0.13101f
C9416 XThR.Tn[6].n8 VGND 0.08099f
C9417 XThR.Tn[6].n9 VGND 0.0914f
C9418 XThR.Tn[6].t62 VGND 0.01453f
C9419 XThR.Tn[6].t56 VGND 0.01591f
C9420 XThR.Tn[6].n10 VGND 0.03884f
C9421 XThR.Tn[6].n11 VGND 0.07461f
C9422 XThR.Tn[6].t20 VGND 0.01453f
C9423 XThR.Tn[6].t72 VGND 0.01591f
C9424 XThR.Tn[6].n12 VGND 0.03884f
C9425 XThR.Tn[6].t36 VGND 0.01448f
C9426 XThR.Tn[6].t68 VGND 0.01585f
C9427 XThR.Tn[6].n13 VGND 0.04041f
C9428 XThR.Tn[6].n14 VGND 0.02839f
C9429 XThR.Tn[6].n16 VGND 0.09111f
C9430 XThR.Tn[6].t57 VGND 0.01453f
C9431 XThR.Tn[6].t49 VGND 0.01591f
C9432 XThR.Tn[6].n17 VGND 0.03884f
C9433 XThR.Tn[6].t14 VGND 0.01448f
C9434 XThR.Tn[6].t45 VGND 0.01585f
C9435 XThR.Tn[6].n18 VGND 0.04041f
C9436 XThR.Tn[6].n19 VGND 0.02839f
C9437 XThR.Tn[6].n21 VGND 0.09111f
C9438 XThR.Tn[6].t73 VGND 0.01453f
C9439 XThR.Tn[6].t66 VGND 0.01591f
C9440 XThR.Tn[6].n22 VGND 0.03884f
C9441 XThR.Tn[6].t26 VGND 0.01448f
C9442 XThR.Tn[6].t63 VGND 0.01585f
C9443 XThR.Tn[6].n23 VGND 0.04041f
C9444 XThR.Tn[6].n24 VGND 0.02839f
C9445 XThR.Tn[6].n26 VGND 0.09111f
C9446 XThR.Tn[6].t35 VGND 0.01453f
C9447 XThR.Tn[6].t31 VGND 0.01591f
C9448 XThR.Tn[6].n27 VGND 0.03884f
C9449 XThR.Tn[6].t59 VGND 0.01448f
C9450 XThR.Tn[6].t27 VGND 0.01585f
C9451 XThR.Tn[6].n28 VGND 0.04041f
C9452 XThR.Tn[6].n29 VGND 0.02839f
C9453 XThR.Tn[6].n31 VGND 0.09111f
C9454 XThR.Tn[6].t13 VGND 0.01453f
C9455 XThR.Tn[6].t67 VGND 0.01591f
C9456 XThR.Tn[6].n32 VGND 0.03884f
C9457 XThR.Tn[6].t29 VGND 0.01448f
C9458 XThR.Tn[6].t64 VGND 0.01585f
C9459 XThR.Tn[6].n33 VGND 0.04041f
C9460 XThR.Tn[6].n34 VGND 0.02839f
C9461 XThR.Tn[6].n36 VGND 0.09111f
C9462 XThR.Tn[6].t51 VGND 0.01453f
C9463 XThR.Tn[6].t22 VGND 0.01591f
C9464 XThR.Tn[6].n37 VGND 0.03884f
C9465 XThR.Tn[6].t70 VGND 0.01448f
C9466 XThR.Tn[6].t19 VGND 0.01585f
C9467 XThR.Tn[6].n38 VGND 0.04041f
C9468 XThR.Tn[6].n39 VGND 0.02839f
C9469 XThR.Tn[6].n41 VGND 0.09111f
C9470 XThR.Tn[6].t21 VGND 0.01453f
C9471 XThR.Tn[6].t17 VGND 0.01591f
C9472 XThR.Tn[6].n42 VGND 0.03884f
C9473 XThR.Tn[6].t37 VGND 0.01448f
C9474 XThR.Tn[6].t12 VGND 0.01585f
C9475 XThR.Tn[6].n43 VGND 0.04041f
C9476 XThR.Tn[6].n44 VGND 0.02839f
C9477 XThR.Tn[6].n46 VGND 0.09111f
C9478 XThR.Tn[6].t24 VGND 0.01453f
C9479 XThR.Tn[6].t30 VGND 0.01591f
C9480 XThR.Tn[6].n47 VGND 0.03884f
C9481 XThR.Tn[6].t43 VGND 0.01448f
C9482 XThR.Tn[6].t25 VGND 0.01585f
C9483 XThR.Tn[6].n48 VGND 0.04041f
C9484 XThR.Tn[6].n49 VGND 0.02839f
C9485 XThR.Tn[6].n51 VGND 0.09111f
C9486 XThR.Tn[6].t40 VGND 0.01453f
C9487 XThR.Tn[6].t50 VGND 0.01591f
C9488 XThR.Tn[6].n52 VGND 0.03884f
C9489 XThR.Tn[6].t61 VGND 0.01448f
C9490 XThR.Tn[6].t47 VGND 0.01585f
C9491 XThR.Tn[6].n53 VGND 0.04041f
C9492 XThR.Tn[6].n54 VGND 0.02839f
C9493 XThR.Tn[6].n56 VGND 0.09111f
C9494 XThR.Tn[6].t33 VGND 0.01453f
C9495 XThR.Tn[6].t69 VGND 0.01591f
C9496 XThR.Tn[6].n57 VGND 0.03884f
C9497 XThR.Tn[6].t54 VGND 0.01448f
C9498 XThR.Tn[6].t65 VGND 0.01585f
C9499 XThR.Tn[6].n58 VGND 0.04041f
C9500 XThR.Tn[6].n59 VGND 0.02839f
C9501 XThR.Tn[6].n61 VGND 0.09111f
C9502 XThR.Tn[6].t53 VGND 0.01453f
C9503 XThR.Tn[6].t44 VGND 0.01591f
C9504 XThR.Tn[6].n62 VGND 0.03884f
C9505 XThR.Tn[6].t71 VGND 0.01448f
C9506 XThR.Tn[6].t39 VGND 0.01585f
C9507 XThR.Tn[6].n63 VGND 0.04041f
C9508 XThR.Tn[6].n64 VGND 0.02839f
C9509 XThR.Tn[6].n66 VGND 0.09111f
C9510 XThR.Tn[6].t23 VGND 0.01453f
C9511 XThR.Tn[6].t18 VGND 0.01591f
C9512 XThR.Tn[6].n67 VGND 0.03884f
C9513 XThR.Tn[6].t41 VGND 0.01448f
C9514 XThR.Tn[6].t15 VGND 0.01585f
C9515 XThR.Tn[6].n68 VGND 0.04041f
C9516 XThR.Tn[6].n69 VGND 0.02839f
C9517 XThR.Tn[6].n71 VGND 0.09111f
C9518 XThR.Tn[6].t38 VGND 0.01453f
C9519 XThR.Tn[6].t32 VGND 0.01591f
C9520 XThR.Tn[6].n72 VGND 0.03884f
C9521 XThR.Tn[6].t60 VGND 0.01448f
C9522 XThR.Tn[6].t28 VGND 0.01585f
C9523 XThR.Tn[6].n73 VGND 0.04041f
C9524 XThR.Tn[6].n74 VGND 0.02839f
C9525 XThR.Tn[6].n76 VGND 0.09111f
C9526 XThR.Tn[6].t58 VGND 0.01453f
C9527 XThR.Tn[6].t52 VGND 0.01591f
C9528 XThR.Tn[6].n77 VGND 0.03884f
C9529 XThR.Tn[6].t16 VGND 0.01448f
C9530 XThR.Tn[6].t48 VGND 0.01585f
C9531 XThR.Tn[6].n78 VGND 0.04041f
C9532 XThR.Tn[6].n79 VGND 0.02839f
C9533 XThR.Tn[6].n81 VGND 0.09111f
C9534 XThR.Tn[6].t34 VGND 0.01453f
C9535 XThR.Tn[6].t46 VGND 0.01591f
C9536 XThR.Tn[6].n82 VGND 0.03884f
C9537 XThR.Tn[6].t55 VGND 0.01448f
C9538 XThR.Tn[6].t42 VGND 0.01585f
C9539 XThR.Tn[6].n83 VGND 0.04041f
C9540 XThR.Tn[6].n84 VGND 0.02839f
C9541 XThR.Tn[6].n86 VGND 0.09111f
C9542 XThR.Tn[6].n87 VGND 0.08279f
C9543 XThR.Tn[6].n88 VGND 0.13782f
C9544 XThC.Tn[10].t2 VGND 0.01051f
C9545 XThC.Tn[10].t7 VGND 0.01051f
C9546 XThC.Tn[10].n0 VGND 0.02621f
C9547 XThC.Tn[10].t11 VGND 0.01051f
C9548 XThC.Tn[10].t3 VGND 0.01051f
C9549 XThC.Tn[10].n1 VGND 0.02101f
C9550 XThC.Tn[10].n2 VGND 0.05286f
C9551 XThC.Tn[10].n3 VGND 0.02293f
C9552 XThC.Tn[10].t38 VGND 0.01281f
C9553 XThC.Tn[10].t36 VGND 0.014f
C9554 XThC.Tn[10].n4 VGND 0.03124f
C9555 XThC.Tn[10].n5 VGND 0.0214f
C9556 XThC.Tn[10].n6 VGND 0.07025f
C9557 XThC.Tn[10].t24 VGND 0.01281f
C9558 XThC.Tn[10].t21 VGND 0.014f
C9559 XThC.Tn[10].n7 VGND 0.03124f
C9560 XThC.Tn[10].n8 VGND 0.0214f
C9561 XThC.Tn[10].n9 VGND 0.07045f
C9562 XThC.Tn[10].n10 VGND 0.1161f
C9563 XThC.Tn[10].t29 VGND 0.01281f
C9564 XThC.Tn[10].t23 VGND 0.014f
C9565 XThC.Tn[10].n11 VGND 0.03124f
C9566 XThC.Tn[10].n12 VGND 0.0214f
C9567 XThC.Tn[10].n13 VGND 0.07045f
C9568 XThC.Tn[10].n14 VGND 0.1161f
C9569 XThC.Tn[10].t30 VGND 0.01281f
C9570 XThC.Tn[10].t25 VGND 0.014f
C9571 XThC.Tn[10].n15 VGND 0.03124f
C9572 XThC.Tn[10].n16 VGND 0.0214f
C9573 XThC.Tn[10].n17 VGND 0.07045f
C9574 XThC.Tn[10].n18 VGND 0.1161f
C9575 XThC.Tn[10].t17 VGND 0.01281f
C9576 XThC.Tn[10].t14 VGND 0.014f
C9577 XThC.Tn[10].n19 VGND 0.03124f
C9578 XThC.Tn[10].n20 VGND 0.0214f
C9579 XThC.Tn[10].n21 VGND 0.07045f
C9580 XThC.Tn[10].n22 VGND 0.1161f
C9581 XThC.Tn[10].t18 VGND 0.01281f
C9582 XThC.Tn[10].t15 VGND 0.014f
C9583 XThC.Tn[10].n23 VGND 0.03124f
C9584 XThC.Tn[10].n24 VGND 0.0214f
C9585 XThC.Tn[10].n25 VGND 0.07045f
C9586 XThC.Tn[10].n26 VGND 0.1161f
C9587 XThC.Tn[10].t34 VGND 0.01281f
C9588 XThC.Tn[10].t28 VGND 0.014f
C9589 XThC.Tn[10].n27 VGND 0.03124f
C9590 XThC.Tn[10].n28 VGND 0.0214f
C9591 XThC.Tn[10].n29 VGND 0.07045f
C9592 XThC.Tn[10].n30 VGND 0.1161f
C9593 XThC.Tn[10].t41 VGND 0.01281f
C9594 XThC.Tn[10].t37 VGND 0.014f
C9595 XThC.Tn[10].n31 VGND 0.03124f
C9596 XThC.Tn[10].n32 VGND 0.0214f
C9597 XThC.Tn[10].n33 VGND 0.07045f
C9598 XThC.Tn[10].n34 VGND 0.1161f
C9599 XThC.Tn[10].t43 VGND 0.01281f
C9600 XThC.Tn[10].t39 VGND 0.014f
C9601 XThC.Tn[10].n35 VGND 0.03124f
C9602 XThC.Tn[10].n36 VGND 0.0214f
C9603 XThC.Tn[10].n37 VGND 0.07045f
C9604 XThC.Tn[10].n38 VGND 0.1161f
C9605 XThC.Tn[10].t31 VGND 0.01281f
C9606 XThC.Tn[10].t26 VGND 0.014f
C9607 XThC.Tn[10].n39 VGND 0.03124f
C9608 XThC.Tn[10].n40 VGND 0.0214f
C9609 XThC.Tn[10].n41 VGND 0.07045f
C9610 XThC.Tn[10].n42 VGND 0.1161f
C9611 XThC.Tn[10].t33 VGND 0.01281f
C9612 XThC.Tn[10].t27 VGND 0.014f
C9613 XThC.Tn[10].n43 VGND 0.03124f
C9614 XThC.Tn[10].n44 VGND 0.0214f
C9615 XThC.Tn[10].n45 VGND 0.07045f
C9616 XThC.Tn[10].n46 VGND 0.1161f
C9617 XThC.Tn[10].t12 VGND 0.01281f
C9618 XThC.Tn[10].t40 VGND 0.014f
C9619 XThC.Tn[10].n47 VGND 0.03124f
C9620 XThC.Tn[10].n48 VGND 0.0214f
C9621 XThC.Tn[10].n49 VGND 0.07045f
C9622 XThC.Tn[10].n50 VGND 0.1161f
C9623 XThC.Tn[10].t20 VGND 0.01281f
C9624 XThC.Tn[10].t16 VGND 0.014f
C9625 XThC.Tn[10].n51 VGND 0.03124f
C9626 XThC.Tn[10].n52 VGND 0.0214f
C9627 XThC.Tn[10].n53 VGND 0.07045f
C9628 XThC.Tn[10].n54 VGND 0.1161f
C9629 XThC.Tn[10].t22 VGND 0.01281f
C9630 XThC.Tn[10].t19 VGND 0.014f
C9631 XThC.Tn[10].n55 VGND 0.03124f
C9632 XThC.Tn[10].n56 VGND 0.0214f
C9633 XThC.Tn[10].n57 VGND 0.07045f
C9634 XThC.Tn[10].n58 VGND 0.1161f
C9635 XThC.Tn[10].t35 VGND 0.01281f
C9636 XThC.Tn[10].t32 VGND 0.014f
C9637 XThC.Tn[10].n59 VGND 0.03124f
C9638 XThC.Tn[10].n60 VGND 0.0214f
C9639 XThC.Tn[10].n61 VGND 0.07045f
C9640 XThC.Tn[10].n62 VGND 0.1161f
C9641 XThC.Tn[10].t13 VGND 0.01281f
C9642 XThC.Tn[10].t42 VGND 0.014f
C9643 XThC.Tn[10].n63 VGND 0.03124f
C9644 XThC.Tn[10].n64 VGND 0.0214f
C9645 XThC.Tn[10].n65 VGND 0.07045f
C9646 XThC.Tn[10].n66 VGND 0.1161f
C9647 XThC.Tn[10].n67 VGND 0.49806f
C9648 XThC.Tn[10].n68 VGND 0.18958f
C9649 XThC.Tn[10].t6 VGND 0.01617f
C9650 XThC.Tn[10].t5 VGND 0.01617f
C9651 XThC.Tn[10].n69 VGND 0.03493f
C9652 XThC.Tn[10].t10 VGND 0.01617f
C9653 XThC.Tn[10].t1 VGND 0.01617f
C9654 XThC.Tn[10].n70 VGND 0.05316f
C9655 XThC.Tn[10].n71 VGND 0.1477f
C9656 XThC.Tn[10].n72 VGND 0.02322f
C9657 XThC.Tn[10].t4 VGND 0.01617f
C9658 XThC.Tn[10].t8 VGND 0.01617f
C9659 XThC.Tn[10].n73 VGND 0.03593f
C9660 XThC.Tn[10].t0 VGND 0.01617f
C9661 XThC.Tn[10].t9 VGND 0.01617f
C9662 XThC.Tn[10].n74 VGND 0.04908f
C9663 XThC.Tn[10].n75 VGND 0.15993f
C9664 Iout.n0 VGND 0.22693f
C9665 Iout.n1 VGND 1.18657f
C9666 Iout.n2 VGND 0.22693f
C9667 Iout.n3 VGND 0.22693f
C9668 Iout.t21 VGND 0.02185f
C9669 Iout.n4 VGND 0.04859f
C9670 Iout.n5 VGND 0.19196f
C9671 Iout.n6 VGND 0.22693f
C9672 Iout.n7 VGND 1.18657f
C9673 Iout.n8 VGND 0.22693f
C9674 Iout.t31 VGND 0.02185f
C9675 Iout.n9 VGND 0.04859f
C9676 Iout.n10 VGND 0.19196f
C9677 Iout.n11 VGND 0.22693f
C9678 Iout.n12 VGND 1.18657f
C9679 Iout.n13 VGND 0.22693f
C9680 Iout.t157 VGND 0.02185f
C9681 Iout.n14 VGND 0.04859f
C9682 Iout.n15 VGND 0.19196f
C9683 Iout.n16 VGND 0.22693f
C9684 Iout.n17 VGND 1.18657f
C9685 Iout.n18 VGND 0.22693f
C9686 Iout.t50 VGND 0.02185f
C9687 Iout.n19 VGND 0.04859f
C9688 Iout.n20 VGND 0.19196f
C9689 Iout.n21 VGND 0.47048f
C9690 Iout.t57 VGND 0.02185f
C9691 Iout.n22 VGND 0.04859f
C9692 Iout.n23 VGND 0.28309f
C9693 Iout.n24 VGND 0.22693f
C9694 Iout.n25 VGND 0.22693f
C9695 Iout.n26 VGND 0.22693f
C9696 Iout.n27 VGND 0.22693f
C9697 Iout.n28 VGND 0.22693f
C9698 Iout.n29 VGND 0.22693f
C9699 Iout.n30 VGND 0.22693f
C9700 Iout.n31 VGND 0.22693f
C9701 Iout.n32 VGND 0.22693f
C9702 Iout.n33 VGND 0.22693f
C9703 Iout.n34 VGND 0.22693f
C9704 Iout.n35 VGND 0.22693f
C9705 Iout.n36 VGND 0.22693f
C9706 Iout.n37 VGND 0.22693f
C9707 Iout.t103 VGND 0.02185f
C9708 Iout.n38 VGND 0.04859f
C9709 Iout.n39 VGND 0.02471f
C9710 Iout.n40 VGND 0.22693f
C9711 Iout.n41 VGND 0.04528f
C9712 Iout.t244 VGND 0.02185f
C9713 Iout.n42 VGND 0.04859f
C9714 Iout.n43 VGND 0.02471f
C9715 Iout.t67 VGND 0.02185f
C9716 Iout.n44 VGND 0.04859f
C9717 Iout.n45 VGND 0.02471f
C9718 Iout.n46 VGND 0.22693f
C9719 Iout.t199 VGND 0.02185f
C9720 Iout.n47 VGND 0.04859f
C9721 Iout.n48 VGND 0.02471f
C9722 Iout.n49 VGND 0.22693f
C9723 Iout.t218 VGND 0.02185f
C9724 Iout.n50 VGND 0.04859f
C9725 Iout.n51 VGND 0.02471f
C9726 Iout.n52 VGND 0.22693f
C9727 Iout.t123 VGND 0.02185f
C9728 Iout.n53 VGND 0.04859f
C9729 Iout.n54 VGND 0.02471f
C9730 Iout.n55 VGND 0.22693f
C9731 Iout.t159 VGND 0.02185f
C9732 Iout.n56 VGND 0.04859f
C9733 Iout.n57 VGND 0.02471f
C9734 Iout.n58 VGND 0.22693f
C9735 Iout.t170 VGND 0.02185f
C9736 Iout.n59 VGND 0.04859f
C9737 Iout.n60 VGND 0.02471f
C9738 Iout.n61 VGND 0.22693f
C9739 Iout.t198 VGND 0.02185f
C9740 Iout.n62 VGND 0.04859f
C9741 Iout.n63 VGND 0.02471f
C9742 Iout.n64 VGND 0.22693f
C9743 Iout.t65 VGND 0.02185f
C9744 Iout.n65 VGND 0.04859f
C9745 Iout.n66 VGND 0.02471f
C9746 Iout.n67 VGND 0.22693f
C9747 Iout.t37 VGND 0.02185f
C9748 Iout.n68 VGND 0.04859f
C9749 Iout.n69 VGND 0.02471f
C9750 Iout.n70 VGND 0.22693f
C9751 Iout.t211 VGND 0.02185f
C9752 Iout.n71 VGND 0.04859f
C9753 Iout.n72 VGND 0.02471f
C9754 Iout.n73 VGND 0.22693f
C9755 Iout.t105 VGND 0.02185f
C9756 Iout.n74 VGND 0.04859f
C9757 Iout.n75 VGND 0.02471f
C9758 Iout.n76 VGND 0.22693f
C9759 Iout.t132 VGND 0.02185f
C9760 Iout.n77 VGND 0.04859f
C9761 Iout.n78 VGND 0.02471f
C9762 Iout.n79 VGND 0.22693f
C9763 Iout.n80 VGND 0.22693f
C9764 Iout.t187 VGND 0.02185f
C9765 Iout.n81 VGND 0.04859f
C9766 Iout.n82 VGND 0.02471f
C9767 Iout.n83 VGND 0.22693f
C9768 Iout.n84 VGND 0.04528f
C9769 Iout.t77 VGND 0.02185f
C9770 Iout.n85 VGND 0.04859f
C9771 Iout.n86 VGND 0.02471f
C9772 Iout.t192 VGND 0.02185f
C9773 Iout.n87 VGND 0.04859f
C9774 Iout.n88 VGND 0.02471f
C9775 Iout.n89 VGND 0.22693f
C9776 Iout.t52 VGND 0.02185f
C9777 Iout.n90 VGND 0.04859f
C9778 Iout.n91 VGND 0.02471f
C9779 Iout.n92 VGND 0.22693f
C9780 Iout.t79 VGND 0.02185f
C9781 Iout.n93 VGND 0.04859f
C9782 Iout.n94 VGND 0.02471f
C9783 Iout.n95 VGND 0.22693f
C9784 Iout.t238 VGND 0.02185f
C9785 Iout.n96 VGND 0.04859f
C9786 Iout.n97 VGND 0.02471f
C9787 Iout.n98 VGND 0.22693f
C9788 Iout.t48 VGND 0.02185f
C9789 Iout.n99 VGND 0.04859f
C9790 Iout.n100 VGND 0.02471f
C9791 Iout.n101 VGND 0.22693f
C9792 Iout.t188 VGND 0.02185f
C9793 Iout.n102 VGND 0.04859f
C9794 Iout.n103 VGND 0.02471f
C9795 Iout.n104 VGND 0.22693f
C9796 Iout.t138 VGND 0.02185f
C9797 Iout.n105 VGND 0.04859f
C9798 Iout.n106 VGND 0.02471f
C9799 Iout.n107 VGND 0.22693f
C9800 Iout.t239 VGND 0.02185f
C9801 Iout.n108 VGND 0.04859f
C9802 Iout.n109 VGND 0.02471f
C9803 Iout.n110 VGND 0.22693f
C9804 Iout.t84 VGND 0.02185f
C9805 Iout.n111 VGND 0.04859f
C9806 Iout.n112 VGND 0.02471f
C9807 Iout.n113 VGND 0.22693f
C9808 Iout.t161 VGND 0.02185f
C9809 Iout.n114 VGND 0.04859f
C9810 Iout.n115 VGND 0.02471f
C9811 Iout.n116 VGND 0.22693f
C9812 Iout.t34 VGND 0.02185f
C9813 Iout.n117 VGND 0.04859f
C9814 Iout.n118 VGND 0.02471f
C9815 Iout.n119 VGND 0.22693f
C9816 Iout.t240 VGND 0.02185f
C9817 Iout.n120 VGND 0.04859f
C9818 Iout.n121 VGND 0.02471f
C9819 Iout.n122 VGND 0.04528f
C9820 Iout.t148 VGND 0.02185f
C9821 Iout.n123 VGND 0.04859f
C9822 Iout.n124 VGND 0.02471f
C9823 Iout.n125 VGND 0.22693f
C9824 Iout.n126 VGND 0.22693f
C9825 Iout.t78 VGND 0.02185f
C9826 Iout.n127 VGND 0.04859f
C9827 Iout.n128 VGND 0.02471f
C9828 Iout.n129 VGND 0.04528f
C9829 Iout.t232 VGND 0.02185f
C9830 Iout.n130 VGND 0.04859f
C9831 Iout.n131 VGND 0.02471f
C9832 Iout.n132 VGND 0.22693f
C9833 Iout.t220 VGND 0.02185f
C9834 Iout.n133 VGND 0.04859f
C9835 Iout.n134 VGND 0.02471f
C9836 Iout.n135 VGND 0.04528f
C9837 Iout.t55 VGND 0.02185f
C9838 Iout.n136 VGND 0.04859f
C9839 Iout.n137 VGND 0.02471f
C9840 Iout.n138 VGND 0.22693f
C9841 Iout.n139 VGND 0.22693f
C9842 Iout.t135 VGND 0.02185f
C9843 Iout.n140 VGND 0.04859f
C9844 Iout.n141 VGND 0.02471f
C9845 Iout.n142 VGND 0.04528f
C9846 Iout.t91 VGND 0.02185f
C9847 Iout.n143 VGND 0.04859f
C9848 Iout.n144 VGND 0.02471f
C9849 Iout.n145 VGND 0.13396f
C9850 Iout.t145 VGND 0.02185f
C9851 Iout.n146 VGND 0.04859f
C9852 Iout.n147 VGND 0.02471f
C9853 Iout.n148 VGND 0.04528f
C9854 Iout.t153 VGND 0.02185f
C9855 Iout.n149 VGND 0.04859f
C9856 Iout.n150 VGND 0.02471f
C9857 Iout.n151 VGND 0.22693f
C9858 Iout.n152 VGND 0.13396f
C9859 Iout.n153 VGND 0.22693f
C9860 Iout.n154 VGND 0.22693f
C9861 Iout.n155 VGND 0.22693f
C9862 Iout.t108 VGND 0.02185f
C9863 Iout.n156 VGND 0.04859f
C9864 Iout.n157 VGND 0.02471f
C9865 Iout.n158 VGND 0.22693f
C9866 Iout.n159 VGND 0.22693f
C9867 Iout.n160 VGND 0.22693f
C9868 Iout.n161 VGND 0.22693f
C9869 Iout.n162 VGND 0.22693f
C9870 Iout.n163 VGND 0.22693f
C9871 Iout.n164 VGND 0.22693f
C9872 Iout.n165 VGND 0.22693f
C9873 Iout.n166 VGND 0.22693f
C9874 Iout.n167 VGND 0.22693f
C9875 Iout.t80 VGND 0.02185f
C9876 Iout.n168 VGND 0.04859f
C9877 Iout.n169 VGND 0.02471f
C9878 Iout.n170 VGND 0.22693f
C9879 Iout.n171 VGND 0.04528f
C9880 Iout.t134 VGND 0.02185f
C9881 Iout.n172 VGND 0.04859f
C9882 Iout.n173 VGND 0.02471f
C9883 Iout.t76 VGND 0.02185f
C9884 Iout.n174 VGND 0.04859f
C9885 Iout.n175 VGND 0.02471f
C9886 Iout.n176 VGND 0.22693f
C9887 Iout.t255 VGND 0.02185f
C9888 Iout.n177 VGND 0.04859f
C9889 Iout.n178 VGND 0.02471f
C9890 Iout.n179 VGND 0.22693f
C9891 Iout.t245 VGND 0.02185f
C9892 Iout.n180 VGND 0.04859f
C9893 Iout.n181 VGND 0.02471f
C9894 Iout.n182 VGND 0.22693f
C9895 Iout.t5 VGND 0.02185f
C9896 Iout.n183 VGND 0.04859f
C9897 Iout.n184 VGND 0.02471f
C9898 Iout.n185 VGND 0.22693f
C9899 Iout.t182 VGND 0.02185f
C9900 Iout.n186 VGND 0.04859f
C9901 Iout.n187 VGND 0.02471f
C9902 Iout.n188 VGND 0.22693f
C9903 Iout.t248 VGND 0.02185f
C9904 Iout.n189 VGND 0.04859f
C9905 Iout.n190 VGND 0.02471f
C9906 Iout.n191 VGND 0.13396f
C9907 Iout.t234 VGND 0.02185f
C9908 Iout.n192 VGND 0.04859f
C9909 Iout.n193 VGND 0.02471f
C9910 Iout.n194 VGND 0.04528f
C9911 Iout.t133 VGND 0.02185f
C9912 Iout.n195 VGND 0.04859f
C9913 Iout.n196 VGND 0.02471f
C9914 Iout.n197 VGND 0.13396f
C9915 Iout.n198 VGND 0.04528f
C9916 Iout.t20 VGND 0.02185f
C9917 Iout.n199 VGND 0.04859f
C9918 Iout.n200 VGND 0.02471f
C9919 Iout.n201 VGND 0.04528f
C9920 Iout.t35 VGND 0.02185f
C9921 Iout.n202 VGND 0.04859f
C9922 Iout.n203 VGND 0.02471f
C9923 Iout.n204 VGND 0.13396f
C9924 Iout.n205 VGND 0.04528f
C9925 Iout.t61 VGND 0.02185f
C9926 Iout.n206 VGND 0.04859f
C9927 Iout.n207 VGND 0.02471f
C9928 Iout.n208 VGND 0.13396f
C9929 Iout.n209 VGND 0.04528f
C9930 Iout.t205 VGND 0.02185f
C9931 Iout.n210 VGND 0.04859f
C9932 Iout.n211 VGND 0.02471f
C9933 Iout.n212 VGND 0.13396f
C9934 Iout.n213 VGND 0.04528f
C9935 Iout.t62 VGND 0.02185f
C9936 Iout.n214 VGND 0.04859f
C9937 Iout.n215 VGND 0.02471f
C9938 Iout.n216 VGND 0.13396f
C9939 Iout.n217 VGND 0.04528f
C9940 Iout.t160 VGND 0.02185f
C9941 Iout.n218 VGND 0.04859f
C9942 Iout.n219 VGND 0.02471f
C9943 Iout.n220 VGND 0.13396f
C9944 Iout.n221 VGND 0.04528f
C9945 Iout.t139 VGND 0.02185f
C9946 Iout.n222 VGND 0.04859f
C9947 Iout.n223 VGND 0.02471f
C9948 Iout.n224 VGND 0.13396f
C9949 Iout.n225 VGND 0.04528f
C9950 Iout.t75 VGND 0.02185f
C9951 Iout.n226 VGND 0.04859f
C9952 Iout.n227 VGND 0.02471f
C9953 Iout.n228 VGND 0.04528f
C9954 Iout.n229 VGND 0.13396f
C9955 Iout.n230 VGND 0.22693f
C9956 Iout.n231 VGND 0.04528f
C9957 Iout.t117 VGND 0.02185f
C9958 Iout.n232 VGND 0.04859f
C9959 Iout.n233 VGND 0.02471f
C9960 Iout.n234 VGND 0.04528f
C9961 Iout.t72 VGND 0.02185f
C9962 Iout.n235 VGND 0.04859f
C9963 Iout.n236 VGND 0.02471f
C9964 Iout.n237 VGND 0.04528f
C9965 Iout.t3 VGND 0.02185f
C9966 Iout.n238 VGND 0.04859f
C9967 Iout.n239 VGND 0.02471f
C9968 Iout.n240 VGND 0.04528f
C9969 Iout.t118 VGND 0.02185f
C9970 Iout.n241 VGND 0.04859f
C9971 Iout.n242 VGND 0.02471f
C9972 Iout.n243 VGND 0.04528f
C9973 Iout.t216 VGND 0.02185f
C9974 Iout.n244 VGND 0.04859f
C9975 Iout.n245 VGND 0.02471f
C9976 Iout.n246 VGND 0.04528f
C9977 Iout.t42 VGND 0.02185f
C9978 Iout.n247 VGND 0.04859f
C9979 Iout.n248 VGND 0.02471f
C9980 Iout.n249 VGND 0.04528f
C9981 Iout.t178 VGND 0.02185f
C9982 Iout.n250 VGND 0.04859f
C9983 Iout.n251 VGND 0.02471f
C9984 Iout.t121 VGND 0.02185f
C9985 Iout.n252 VGND 0.04859f
C9986 Iout.n253 VGND 0.02471f
C9987 Iout.n254 VGND 0.04528f
C9988 Iout.t110 VGND 0.02185f
C9989 Iout.n255 VGND 0.04859f
C9990 Iout.n256 VGND 0.02471f
C9991 Iout.n257 VGND 0.04528f
C9992 Iout.n258 VGND 0.22693f
C9993 Iout.t13 VGND 0.02185f
C9994 Iout.n259 VGND 0.04859f
C9995 Iout.n260 VGND 0.02471f
C9996 Iout.n261 VGND 0.04528f
C9997 Iout.n262 VGND 0.22693f
C9998 Iout.n263 VGND 0.22693f
C9999 Iout.n264 VGND 0.04528f
C10000 Iout.t210 VGND 0.02185f
C10001 Iout.n265 VGND 0.04859f
C10002 Iout.n266 VGND 0.02471f
C10003 Iout.n267 VGND 0.04528f
C10004 Iout.n268 VGND 0.22693f
C10005 Iout.n269 VGND 0.22693f
C10006 Iout.n270 VGND 0.04528f
C10007 Iout.t243 VGND 0.02185f
C10008 Iout.n271 VGND 0.04859f
C10009 Iout.n272 VGND 0.02471f
C10010 Iout.n273 VGND 0.04528f
C10011 Iout.n274 VGND 0.22693f
C10012 Iout.n275 VGND 0.22693f
C10013 Iout.n276 VGND 0.04528f
C10014 Iout.t179 VGND 0.02185f
C10015 Iout.n277 VGND 0.04859f
C10016 Iout.n278 VGND 0.02471f
C10017 Iout.n279 VGND 0.04528f
C10018 Iout.n280 VGND 0.22693f
C10019 Iout.n281 VGND 0.22693f
C10020 Iout.n282 VGND 0.04528f
C10021 Iout.t114 VGND 0.02185f
C10022 Iout.n283 VGND 0.04859f
C10023 Iout.n284 VGND 0.02471f
C10024 Iout.n285 VGND 0.04528f
C10025 Iout.n286 VGND 0.22693f
C10026 Iout.n287 VGND 0.22693f
C10027 Iout.n288 VGND 0.04528f
C10028 Iout.t226 VGND 0.02185f
C10029 Iout.n289 VGND 0.04859f
C10030 Iout.n290 VGND 0.02471f
C10031 Iout.n291 VGND 0.04528f
C10032 Iout.n292 VGND 0.22693f
C10033 Iout.n293 VGND 0.22693f
C10034 Iout.n294 VGND 0.04528f
C10035 Iout.t181 VGND 0.02185f
C10036 Iout.n295 VGND 0.04859f
C10037 Iout.n296 VGND 0.02471f
C10038 Iout.n297 VGND 0.04528f
C10039 Iout.n298 VGND 0.22693f
C10040 Iout.n299 VGND 0.22693f
C10041 Iout.n300 VGND 0.04528f
C10042 Iout.t2 VGND 0.02185f
C10043 Iout.n301 VGND 0.04859f
C10044 Iout.n302 VGND 0.02471f
C10045 Iout.n303 VGND 0.04528f
C10046 Iout.n304 VGND 0.22693f
C10047 Iout.t183 VGND 0.02185f
C10048 Iout.n305 VGND 0.04859f
C10049 Iout.n306 VGND 0.02471f
C10050 Iout.n307 VGND 0.04528f
C10051 Iout.t194 VGND 0.02185f
C10052 Iout.n308 VGND 0.04859f
C10053 Iout.n309 VGND 0.02471f
C10054 Iout.n310 VGND 0.04528f
C10055 Iout.t18 VGND 0.02185f
C10056 Iout.n311 VGND 0.04859f
C10057 Iout.n312 VGND 0.02471f
C10058 Iout.n313 VGND 0.04528f
C10059 Iout.t165 VGND 0.02185f
C10060 Iout.n314 VGND 0.04859f
C10061 Iout.n315 VGND 0.02471f
C10062 Iout.n316 VGND 0.04528f
C10063 Iout.t191 VGND 0.02185f
C10064 Iout.n317 VGND 0.04859f
C10065 Iout.n318 VGND 0.02471f
C10066 Iout.n319 VGND 0.04528f
C10067 Iout.t176 VGND 0.02185f
C10068 Iout.n320 VGND 0.04859f
C10069 Iout.n321 VGND 0.02471f
C10070 Iout.n322 VGND 0.04528f
C10071 Iout.t186 VGND 0.02185f
C10072 Iout.n323 VGND 0.04859f
C10073 Iout.n324 VGND 0.02471f
C10074 Iout.n325 VGND 0.04528f
C10075 Iout.t171 VGND 0.02185f
C10076 Iout.n326 VGND 0.04859f
C10077 Iout.n327 VGND 0.02471f
C10078 Iout.n328 VGND 0.04528f
C10079 Iout.t128 VGND 0.02185f
C10080 Iout.n329 VGND 0.04859f
C10081 Iout.n330 VGND 0.02471f
C10082 Iout.n331 VGND 0.04528f
C10083 Iout.n332 VGND 0.22693f
C10084 Iout.t180 VGND 0.02185f
C10085 Iout.n333 VGND 0.04859f
C10086 Iout.n334 VGND 0.02471f
C10087 Iout.n335 VGND 0.04528f
C10088 Iout.t83 VGND 0.02185f
C10089 Iout.n336 VGND 0.04859f
C10090 Iout.n337 VGND 0.02471f
C10091 Iout.n338 VGND 0.04528f
C10092 Iout.t28 VGND 0.02185f
C10093 Iout.n339 VGND 0.04859f
C10094 Iout.n340 VGND 0.02471f
C10095 Iout.n341 VGND 0.04528f
C10096 Iout.t115 VGND 0.02185f
C10097 Iout.n342 VGND 0.04859f
C10098 Iout.n343 VGND 0.02471f
C10099 Iout.n344 VGND 0.04528f
C10100 Iout.t40 VGND 0.02185f
C10101 Iout.n345 VGND 0.04859f
C10102 Iout.n346 VGND 0.02471f
C10103 Iout.n347 VGND 0.04528f
C10104 Iout.t107 VGND 0.02185f
C10105 Iout.n348 VGND 0.04859f
C10106 Iout.n349 VGND 0.02471f
C10107 Iout.n350 VGND 0.04528f
C10108 Iout.t96 VGND 0.02185f
C10109 Iout.n351 VGND 0.04859f
C10110 Iout.n352 VGND 0.02471f
C10111 Iout.n353 VGND 0.04528f
C10112 Iout.t222 VGND 0.02185f
C10113 Iout.n354 VGND 0.04859f
C10114 Iout.n355 VGND 0.02471f
C10115 Iout.n356 VGND 0.04528f
C10116 Iout.t204 VGND 0.02185f
C10117 Iout.n357 VGND 0.04859f
C10118 Iout.n358 VGND 0.02471f
C10119 Iout.n359 VGND 0.04528f
C10120 Iout.t212 VGND 0.02185f
C10121 Iout.n360 VGND 0.04859f
C10122 Iout.n361 VGND 0.02471f
C10123 Iout.n362 VGND 0.04528f
C10124 Iout.t102 VGND 0.02185f
C10125 Iout.n363 VGND 0.04859f
C10126 Iout.n364 VGND 0.02471f
C10127 Iout.n365 VGND 0.04528f
C10128 Iout.t81 VGND 0.02185f
C10129 Iout.n366 VGND 0.04859f
C10130 Iout.n367 VGND 0.02471f
C10131 Iout.n368 VGND 0.04528f
C10132 Iout.n369 VGND 0.22693f
C10133 Iout.t223 VGND 0.02185f
C10134 Iout.n370 VGND 0.04859f
C10135 Iout.n371 VGND 0.02471f
C10136 Iout.n372 VGND 0.04528f
C10137 Iout.n373 VGND 0.22693f
C10138 Iout.n374 VGND 0.22693f
C10139 Iout.n375 VGND 0.04528f
C10140 Iout.t25 VGND 0.02185f
C10141 Iout.n376 VGND 0.04859f
C10142 Iout.n377 VGND 0.02471f
C10143 Iout.t237 VGND 0.02185f
C10144 Iout.n378 VGND 0.04859f
C10145 Iout.n379 VGND 0.02471f
C10146 Iout.n380 VGND 0.04528f
C10147 Iout.n381 VGND 0.22693f
C10148 Iout.n382 VGND 0.22693f
C10149 Iout.n383 VGND 0.04528f
C10150 Iout.t97 VGND 0.02185f
C10151 Iout.n384 VGND 0.04859f
C10152 Iout.n385 VGND 0.02471f
C10153 Iout.t113 VGND 0.02185f
C10154 Iout.n386 VGND 0.04859f
C10155 Iout.n387 VGND 0.02471f
C10156 Iout.n388 VGND 0.04528f
C10157 Iout.n389 VGND 0.22693f
C10158 Iout.n390 VGND 0.22693f
C10159 Iout.n391 VGND 0.04528f
C10160 Iout.t30 VGND 0.02185f
C10161 Iout.n392 VGND 0.04859f
C10162 Iout.n393 VGND 0.02471f
C10163 Iout.t7 VGND 0.02185f
C10164 Iout.n394 VGND 0.04859f
C10165 Iout.n395 VGND 0.02471f
C10166 Iout.n396 VGND 0.04528f
C10167 Iout.n397 VGND 0.22693f
C10168 Iout.n398 VGND 0.22693f
C10169 Iout.n399 VGND 0.04528f
C10170 Iout.t140 VGND 0.02185f
C10171 Iout.n400 VGND 0.04859f
C10172 Iout.n401 VGND 0.02471f
C10173 Iout.t6 VGND 0.02185f
C10174 Iout.n402 VGND 0.04859f
C10175 Iout.n403 VGND 0.02471f
C10176 Iout.n404 VGND 0.04528f
C10177 Iout.n405 VGND 0.22693f
C10178 Iout.n406 VGND 0.22693f
C10179 Iout.n407 VGND 0.04528f
C10180 Iout.t14 VGND 0.02185f
C10181 Iout.n408 VGND 0.04859f
C10182 Iout.n409 VGND 0.02471f
C10183 Iout.t154 VGND 0.02185f
C10184 Iout.n410 VGND 0.04859f
C10185 Iout.n411 VGND 0.02471f
C10186 Iout.n412 VGND 0.04528f
C10187 Iout.n413 VGND 0.22693f
C10188 Iout.n414 VGND 0.22693f
C10189 Iout.n415 VGND 0.04528f
C10190 Iout.t206 VGND 0.02185f
C10191 Iout.n416 VGND 0.04859f
C10192 Iout.n417 VGND 0.02471f
C10193 Iout.t111 VGND 0.02185f
C10194 Iout.n418 VGND 0.04859f
C10195 Iout.n419 VGND 0.02471f
C10196 Iout.n420 VGND 0.04528f
C10197 Iout.n421 VGND 0.22693f
C10198 Iout.n422 VGND 0.22693f
C10199 Iout.n423 VGND 0.04528f
C10200 Iout.t185 VGND 0.02185f
C10201 Iout.n424 VGND 0.04859f
C10202 Iout.n425 VGND 0.02471f
C10203 Iout.t207 VGND 0.02185f
C10204 Iout.n426 VGND 0.04859f
C10205 Iout.n427 VGND 0.02471f
C10206 Iout.n428 VGND 0.04528f
C10207 Iout.n429 VGND 0.22693f
C10208 Iout.n430 VGND 0.22693f
C10209 Iout.n431 VGND 0.04528f
C10210 Iout.t15 VGND 0.02185f
C10211 Iout.n432 VGND 0.04859f
C10212 Iout.n433 VGND 0.02471f
C10213 Iout.t112 VGND 0.02185f
C10214 Iout.n434 VGND 0.04859f
C10215 Iout.n435 VGND 0.02471f
C10216 Iout.n436 VGND 0.22693f
C10217 Iout.n437 VGND 0.04528f
C10218 Iout.t247 VGND 0.02185f
C10219 Iout.n438 VGND 0.04859f
C10220 Iout.n439 VGND 0.02471f
C10221 Iout.n440 VGND 0.04528f
C10222 Iout.t126 VGND 0.02185f
C10223 Iout.n441 VGND 0.04859f
C10224 Iout.n442 VGND 0.02471f
C10225 Iout.n443 VGND 0.04528f
C10226 Iout.n444 VGND 0.22693f
C10227 Iout.n445 VGND 0.22693f
C10228 Iout.n446 VGND 0.04528f
C10229 Iout.t190 VGND 0.02185f
C10230 Iout.n447 VGND 0.04859f
C10231 Iout.n448 VGND 0.02471f
C10232 Iout.t45 VGND 0.02185f
C10233 Iout.n449 VGND 0.04859f
C10234 Iout.n450 VGND 0.02471f
C10235 Iout.n451 VGND 0.04528f
C10236 Iout.t152 VGND 0.02185f
C10237 Iout.n452 VGND 0.04859f
C10238 Iout.n453 VGND 0.02471f
C10239 Iout.n454 VGND 0.04528f
C10240 Iout.n455 VGND 0.22693f
C10241 Iout.n456 VGND 0.22693f
C10242 Iout.n457 VGND 0.04528f
C10243 Iout.t73 VGND 0.02185f
C10244 Iout.n458 VGND 0.04859f
C10245 Iout.n459 VGND 0.02471f
C10246 Iout.t136 VGND 0.02185f
C10247 Iout.n460 VGND 0.04859f
C10248 Iout.n461 VGND 0.02471f
C10249 Iout.n462 VGND 0.04528f
C10250 Iout.t173 VGND 0.02185f
C10251 Iout.n463 VGND 0.04859f
C10252 Iout.n464 VGND 0.02471f
C10253 Iout.n465 VGND 0.04528f
C10254 Iout.n466 VGND 0.22693f
C10255 Iout.n467 VGND 0.22693f
C10256 Iout.n468 VGND 0.04528f
C10257 Iout.t74 VGND 0.02185f
C10258 Iout.n469 VGND 0.04859f
C10259 Iout.n470 VGND 0.02471f
C10260 Iout.n471 VGND 0.04528f
C10261 Iout.t19 VGND 0.02185f
C10262 Iout.n472 VGND 0.04859f
C10263 Iout.n473 VGND 0.02471f
C10264 Iout.n474 VGND 0.04528f
C10265 Iout.n475 VGND 0.22693f
C10266 Iout.n476 VGND 0.22693f
C10267 Iout.n477 VGND 0.04528f
C10268 Iout.t168 VGND 0.02185f
C10269 Iout.n478 VGND 0.04859f
C10270 Iout.n479 VGND 0.02471f
C10271 Iout.t143 VGND 0.02185f
C10272 Iout.n480 VGND 0.04859f
C10273 Iout.n481 VGND 0.02471f
C10274 Iout.n482 VGND 0.04528f
C10275 Iout.t26 VGND 0.02185f
C10276 Iout.n483 VGND 0.04859f
C10277 Iout.n484 VGND 0.02471f
C10278 Iout.n485 VGND 0.04528f
C10279 Iout.n486 VGND 0.22693f
C10280 Iout.n487 VGND 0.22693f
C10281 Iout.n488 VGND 0.04528f
C10282 Iout.t124 VGND 0.02185f
C10283 Iout.n489 VGND 0.04859f
C10284 Iout.n490 VGND 0.02471f
C10285 Iout.t203 VGND 0.02185f
C10286 Iout.n491 VGND 0.04859f
C10287 Iout.n492 VGND 0.02471f
C10288 Iout.n493 VGND 0.04528f
C10289 Iout.t93 VGND 0.02185f
C10290 Iout.n494 VGND 0.04859f
C10291 Iout.n495 VGND 0.02471f
C10292 Iout.n496 VGND 0.04528f
C10293 Iout.n497 VGND 0.22693f
C10294 Iout.n498 VGND 0.13396f
C10295 Iout.n499 VGND 0.04528f
C10296 Iout.t249 VGND 0.02185f
C10297 Iout.n500 VGND 0.04859f
C10298 Iout.n501 VGND 0.02471f
C10299 Iout.n502 VGND 0.13396f
C10300 Iout.n503 VGND 0.04528f
C10301 Iout.t39 VGND 0.02185f
C10302 Iout.n504 VGND 0.04859f
C10303 Iout.n505 VGND 0.02471f
C10304 Iout.n506 VGND 0.04528f
C10305 Iout.t86 VGND 0.02185f
C10306 Iout.n507 VGND 0.04859f
C10307 Iout.n508 VGND 0.02471f
C10308 Iout.t33 VGND 0.02185f
C10309 Iout.n509 VGND 0.04859f
C10310 Iout.n510 VGND 0.02471f
C10311 Iout.n511 VGND 0.13396f
C10312 Iout.n512 VGND 0.04528f
C10313 Iout.t9 VGND 0.02185f
C10314 Iout.n513 VGND 0.04859f
C10315 Iout.n514 VGND 0.02471f
C10316 Iout.n515 VGND 0.04528f
C10317 Iout.n516 VGND 0.13396f
C10318 Iout.n517 VGND 0.22693f
C10319 Iout.n518 VGND 0.04528f
C10320 Iout.t95 VGND 0.02185f
C10321 Iout.n519 VGND 0.04859f
C10322 Iout.n520 VGND 0.02471f
C10323 Iout.n521 VGND 0.04528f
C10324 Iout.n522 VGND 0.22693f
C10325 Iout.n523 VGND 0.22693f
C10326 Iout.n524 VGND 0.04528f
C10327 Iout.t214 VGND 0.02185f
C10328 Iout.n525 VGND 0.04859f
C10329 Iout.n526 VGND 0.02471f
C10330 Iout.n527 VGND 0.04528f
C10331 Iout.n528 VGND 0.22693f
C10332 Iout.n529 VGND 0.22693f
C10333 Iout.n530 VGND 0.04528f
C10334 Iout.t125 VGND 0.02185f
C10335 Iout.n531 VGND 0.04859f
C10336 Iout.n532 VGND 0.02471f
C10337 Iout.n533 VGND 0.04528f
C10338 Iout.t69 VGND 0.02185f
C10339 Iout.n534 VGND 0.04859f
C10340 Iout.n535 VGND 0.02471f
C10341 Iout.t58 VGND 0.02185f
C10342 Iout.n536 VGND 0.04859f
C10343 Iout.n537 VGND 0.02471f
C10344 Iout.n538 VGND 0.04528f
C10345 Iout.n539 VGND 0.22693f
C10346 Iout.n540 VGND 0.22693f
C10347 Iout.n541 VGND 0.04528f
C10348 Iout.t16 VGND 0.02185f
C10349 Iout.n542 VGND 0.04859f
C10350 Iout.n543 VGND 0.02471f
C10351 Iout.n544 VGND 0.04528f
C10352 Iout.n545 VGND 0.22693f
C10353 Iout.n546 VGND 0.22693f
C10354 Iout.n547 VGND 0.04528f
C10355 Iout.t89 VGND 0.02185f
C10356 Iout.n548 VGND 0.04859f
C10357 Iout.n549 VGND 0.02471f
C10358 Iout.n550 VGND 0.04528f
C10359 Iout.n551 VGND 0.22693f
C10360 Iout.n552 VGND 0.22693f
C10361 Iout.n553 VGND 0.04528f
C10362 Iout.t184 VGND 0.02185f
C10363 Iout.n554 VGND 0.04859f
C10364 Iout.n555 VGND 0.02471f
C10365 Iout.n556 VGND 0.04528f
C10366 Iout.t166 VGND 0.02185f
C10367 Iout.n557 VGND 0.04859f
C10368 Iout.n558 VGND 0.02471f
C10369 Iout.t49 VGND 0.02185f
C10370 Iout.n559 VGND 0.04859f
C10371 Iout.n560 VGND 0.02471f
C10372 Iout.n561 VGND 0.04528f
C10373 Iout.n562 VGND 0.22693f
C10374 Iout.t44 VGND 0.02185f
C10375 Iout.n563 VGND 0.04859f
C10376 Iout.n564 VGND 0.02471f
C10377 Iout.n565 VGND 0.04528f
C10378 Iout.n566 VGND 0.22693f
C10379 Iout.n567 VGND 0.22693f
C10380 Iout.n568 VGND 0.04528f
C10381 Iout.t24 VGND 0.02185f
C10382 Iout.n569 VGND 0.04859f
C10383 Iout.n570 VGND 0.02471f
C10384 Iout.n571 VGND 0.04528f
C10385 Iout.n572 VGND 0.22693f
C10386 Iout.t162 VGND 0.02185f
C10387 Iout.n573 VGND 0.04859f
C10388 Iout.n574 VGND 0.02471f
C10389 Iout.n575 VGND 0.04528f
C10390 Iout.t167 VGND 0.02185f
C10391 Iout.n576 VGND 0.04859f
C10392 Iout.n577 VGND 0.02471f
C10393 Iout.n578 VGND 0.04528f
C10394 Iout.n579 VGND 0.22693f
C10395 Iout.n580 VGND 0.22693f
C10396 Iout.n581 VGND 0.04528f
C10397 Iout.t169 VGND 0.02185f
C10398 Iout.n582 VGND 0.04859f
C10399 Iout.n583 VGND 0.02471f
C10400 Iout.n584 VGND 0.04528f
C10401 Iout.n585 VGND 0.22693f
C10402 Iout.n586 VGND 0.22693f
C10403 Iout.n587 VGND 0.04528f
C10404 Iout.t66 VGND 0.02185f
C10405 Iout.n588 VGND 0.04859f
C10406 Iout.n589 VGND 0.02471f
C10407 Iout.n590 VGND 0.04528f
C10408 Iout.n591 VGND 0.22693f
C10409 Iout.n592 VGND 0.22693f
C10410 Iout.n593 VGND 0.04528f
C10411 Iout.t219 VGND 0.02185f
C10412 Iout.n594 VGND 0.04859f
C10413 Iout.n595 VGND 0.02471f
C10414 Iout.n596 VGND 0.04528f
C10415 Iout.n597 VGND 0.22693f
C10416 Iout.n598 VGND 0.22693f
C10417 Iout.n599 VGND 0.04528f
C10418 Iout.t32 VGND 0.02185f
C10419 Iout.n600 VGND 0.04859f
C10420 Iout.n601 VGND 0.02471f
C10421 Iout.n602 VGND 0.04528f
C10422 Iout.n603 VGND 0.22693f
C10423 Iout.n604 VGND 0.22693f
C10424 Iout.n605 VGND 0.04528f
C10425 Iout.t99 VGND 0.02185f
C10426 Iout.n606 VGND 0.04859f
C10427 Iout.n607 VGND 0.02471f
C10428 Iout.n608 VGND 0.04528f
C10429 Iout.n609 VGND 0.22693f
C10430 Iout.n610 VGND 0.22693f
C10431 Iout.n611 VGND 0.04528f
C10432 Iout.t11 VGND 0.02185f
C10433 Iout.n612 VGND 0.04859f
C10434 Iout.n613 VGND 0.02471f
C10435 Iout.n614 VGND 0.04528f
C10436 Iout.n615 VGND 0.22693f
C10437 Iout.n616 VGND 0.22693f
C10438 Iout.n617 VGND 0.04528f
C10439 Iout.t177 VGND 0.02185f
C10440 Iout.n618 VGND 0.04859f
C10441 Iout.n619 VGND 0.02471f
C10442 Iout.n620 VGND 0.04528f
C10443 Iout.n621 VGND 0.22693f
C10444 Iout.n622 VGND 0.22693f
C10445 Iout.n623 VGND 0.04528f
C10446 Iout.t17 VGND 0.02185f
C10447 Iout.n624 VGND 0.04859f
C10448 Iout.n625 VGND 0.02471f
C10449 Iout.n626 VGND 0.04528f
C10450 Iout.n627 VGND 0.22693f
C10451 Iout.n628 VGND 0.22693f
C10452 Iout.n629 VGND 0.04528f
C10453 Iout.t129 VGND 0.02185f
C10454 Iout.n630 VGND 0.04859f
C10455 Iout.n631 VGND 0.02471f
C10456 Iout.n632 VGND 0.04528f
C10457 Iout.n633 VGND 0.22693f
C10458 Iout.n634 VGND 0.22693f
C10459 Iout.n635 VGND 0.04528f
C10460 Iout.t29 VGND 0.02185f
C10461 Iout.n636 VGND 0.04859f
C10462 Iout.n637 VGND 0.02471f
C10463 Iout.n638 VGND 0.04528f
C10464 Iout.n639 VGND 0.22693f
C10465 Iout.n640 VGND 0.22693f
C10466 Iout.n641 VGND 0.04528f
C10467 Iout.t144 VGND 0.02185f
C10468 Iout.n642 VGND 0.04859f
C10469 Iout.n643 VGND 0.02471f
C10470 Iout.n644 VGND 0.04528f
C10471 Iout.n645 VGND 0.22693f
C10472 Iout.n646 VGND 0.22693f
C10473 Iout.n647 VGND 0.04528f
C10474 Iout.t164 VGND 0.02185f
C10475 Iout.n648 VGND 0.04859f
C10476 Iout.n649 VGND 0.02471f
C10477 Iout.n650 VGND 0.04528f
C10478 Iout.n651 VGND 0.22693f
C10479 Iout.n652 VGND 0.22693f
C10480 Iout.n653 VGND 0.04528f
C10481 Iout.t235 VGND 0.02185f
C10482 Iout.n654 VGND 0.04859f
C10483 Iout.n655 VGND 0.02471f
C10484 Iout.n656 VGND 0.04528f
C10485 Iout.t208 VGND 0.02185f
C10486 Iout.n657 VGND 0.04859f
C10487 Iout.n658 VGND 0.02471f
C10488 Iout.n659 VGND 0.04528f
C10489 Iout.t109 VGND 0.02185f
C10490 Iout.n660 VGND 0.04859f
C10491 Iout.n661 VGND 0.02471f
C10492 Iout.n662 VGND 0.04528f
C10493 Iout.t12 VGND 0.02185f
C10494 Iout.n663 VGND 0.04859f
C10495 Iout.n664 VGND 0.02471f
C10496 Iout.n665 VGND 0.04528f
C10497 Iout.t71 VGND 0.02185f
C10498 Iout.n666 VGND 0.04859f
C10499 Iout.n667 VGND 0.02471f
C10500 Iout.n668 VGND 0.04528f
C10501 Iout.t104 VGND 0.02185f
C10502 Iout.n669 VGND 0.04859f
C10503 Iout.n670 VGND 0.02471f
C10504 Iout.n671 VGND 0.04528f
C10505 Iout.t224 VGND 0.02185f
C10506 Iout.n672 VGND 0.04859f
C10507 Iout.n673 VGND 0.02471f
C10508 Iout.n674 VGND 0.04528f
C10509 Iout.t56 VGND 0.02185f
C10510 Iout.n675 VGND 0.04859f
C10511 Iout.n676 VGND 0.02471f
C10512 Iout.n677 VGND 0.04528f
C10513 Iout.t156 VGND 0.02185f
C10514 Iout.n678 VGND 0.04859f
C10515 Iout.n679 VGND 0.02471f
C10516 Iout.n680 VGND 0.04528f
C10517 Iout.t85 VGND 0.02185f
C10518 Iout.n681 VGND 0.04859f
C10519 Iout.n682 VGND 0.02471f
C10520 Iout.n683 VGND 0.04528f
C10521 Iout.t225 VGND 0.02185f
C10522 Iout.n684 VGND 0.04859f
C10523 Iout.n685 VGND 0.02471f
C10524 Iout.n686 VGND 0.04528f
C10525 Iout.t151 VGND 0.02185f
C10526 Iout.n687 VGND 0.04859f
C10527 Iout.n688 VGND 0.02471f
C10528 Iout.n689 VGND 0.04528f
C10529 Iout.t229 VGND 0.02185f
C10530 Iout.n690 VGND 0.04859f
C10531 Iout.n691 VGND 0.02471f
C10532 Iout.t193 VGND 0.02185f
C10533 Iout.n692 VGND 0.04859f
C10534 Iout.n693 VGND 0.02471f
C10535 Iout.n694 VGND 0.04528f
C10536 Iout.t59 VGND 0.02185f
C10537 Iout.n695 VGND 0.04859f
C10538 Iout.n696 VGND 0.02471f
C10539 Iout.n697 VGND 0.04528f
C10540 Iout.n698 VGND 0.22693f
C10541 Iout.t101 VGND 0.02185f
C10542 Iout.n699 VGND 0.04859f
C10543 Iout.n700 VGND 0.02471f
C10544 Iout.n701 VGND 0.04528f
C10545 Iout.n702 VGND 0.22693f
C10546 Iout.n703 VGND 0.22693f
C10547 Iout.n704 VGND 0.04528f
C10548 Iout.t23 VGND 0.02185f
C10549 Iout.n705 VGND 0.04859f
C10550 Iout.n706 VGND 0.02471f
C10551 Iout.n707 VGND 0.04528f
C10552 Iout.n708 VGND 0.22693f
C10553 Iout.n709 VGND 0.22693f
C10554 Iout.n710 VGND 0.04528f
C10555 Iout.t98 VGND 0.02185f
C10556 Iout.n711 VGND 0.04859f
C10557 Iout.n712 VGND 0.02471f
C10558 Iout.n713 VGND 0.04528f
C10559 Iout.n714 VGND 0.22693f
C10560 Iout.n715 VGND 0.22693f
C10561 Iout.n716 VGND 0.04528f
C10562 Iout.t46 VGND 0.02185f
C10563 Iout.n717 VGND 0.04859f
C10564 Iout.n718 VGND 0.02471f
C10565 Iout.n719 VGND 0.04528f
C10566 Iout.n720 VGND 0.22693f
C10567 Iout.n721 VGND 0.22693f
C10568 Iout.n722 VGND 0.04528f
C10569 Iout.t242 VGND 0.02185f
C10570 Iout.n723 VGND 0.04859f
C10571 Iout.n724 VGND 0.02471f
C10572 Iout.n725 VGND 0.04528f
C10573 Iout.n726 VGND 0.22693f
C10574 Iout.n727 VGND 0.22693f
C10575 Iout.n728 VGND 0.04528f
C10576 Iout.t231 VGND 0.02185f
C10577 Iout.n729 VGND 0.04859f
C10578 Iout.n730 VGND 0.02471f
C10579 Iout.n731 VGND 0.04528f
C10580 Iout.n732 VGND 0.22693f
C10581 Iout.n733 VGND 0.22693f
C10582 Iout.n734 VGND 0.04528f
C10583 Iout.t202 VGND 0.02185f
C10584 Iout.n735 VGND 0.04859f
C10585 Iout.n736 VGND 0.02471f
C10586 Iout.n737 VGND 0.04528f
C10587 Iout.n738 VGND 0.22693f
C10588 Iout.n739 VGND 0.22693f
C10589 Iout.n740 VGND 0.04528f
C10590 Iout.t137 VGND 0.02185f
C10591 Iout.n741 VGND 0.04859f
C10592 Iout.n742 VGND 0.02471f
C10593 Iout.n743 VGND 0.04528f
C10594 Iout.n744 VGND 0.22693f
C10595 Iout.n745 VGND 0.22693f
C10596 Iout.n746 VGND 0.04528f
C10597 Iout.t130 VGND 0.02185f
C10598 Iout.n747 VGND 0.04859f
C10599 Iout.n748 VGND 0.02471f
C10600 Iout.n749 VGND 0.04528f
C10601 Iout.n750 VGND 0.22693f
C10602 Iout.n751 VGND 0.22693f
C10603 Iout.n752 VGND 0.04528f
C10604 Iout.t88 VGND 0.02185f
C10605 Iout.n753 VGND 0.04859f
C10606 Iout.n754 VGND 0.02471f
C10607 Iout.n755 VGND 0.04528f
C10608 Iout.n756 VGND 0.22693f
C10609 Iout.n757 VGND 0.22693f
C10610 Iout.n758 VGND 0.04528f
C10611 Iout.t106 VGND 0.02185f
C10612 Iout.n759 VGND 0.04859f
C10613 Iout.n760 VGND 0.02471f
C10614 Iout.n761 VGND 0.04528f
C10615 Iout.n762 VGND 0.22693f
C10616 Iout.n763 VGND 0.22693f
C10617 Iout.n764 VGND 0.04528f
C10618 Iout.t100 VGND 0.02185f
C10619 Iout.n765 VGND 0.04859f
C10620 Iout.n766 VGND 0.02471f
C10621 Iout.n767 VGND 0.04528f
C10622 Iout.n768 VGND 0.22693f
C10623 Iout.n769 VGND 0.22693f
C10624 Iout.n770 VGND 0.04528f
C10625 Iout.t41 VGND 0.02185f
C10626 Iout.n771 VGND 0.04859f
C10627 Iout.n772 VGND 0.02471f
C10628 Iout.n773 VGND 0.04528f
C10629 Iout.n774 VGND 0.22693f
C10630 Iout.n775 VGND 0.22693f
C10631 Iout.n776 VGND 0.04528f
C10632 Iout.t51 VGND 0.02185f
C10633 Iout.n777 VGND 0.04859f
C10634 Iout.n778 VGND 0.02471f
C10635 Iout.n779 VGND 0.04528f
C10636 Iout.n780 VGND 0.22693f
C10637 Iout.t53 VGND 0.02185f
C10638 Iout.n781 VGND 0.04859f
C10639 Iout.n782 VGND 0.02471f
C10640 Iout.n783 VGND 0.04528f
C10641 Iout.t147 VGND 0.02185f
C10642 Iout.n784 VGND 0.04859f
C10643 Iout.n785 VGND 0.02471f
C10644 Iout.n786 VGND 0.04528f
C10645 Iout.t197 VGND 0.02185f
C10646 Iout.n787 VGND 0.04859f
C10647 Iout.n788 VGND 0.02471f
C10648 Iout.n789 VGND 0.04528f
C10649 Iout.t27 VGND 0.02185f
C10650 Iout.n790 VGND 0.04859f
C10651 Iout.n791 VGND 0.02471f
C10652 Iout.n792 VGND 0.04528f
C10653 Iout.t22 VGND 0.02185f
C10654 Iout.n793 VGND 0.04859f
C10655 Iout.n794 VGND 0.02471f
C10656 Iout.n795 VGND 0.04528f
C10657 Iout.t174 VGND 0.02185f
C10658 Iout.n796 VGND 0.04859f
C10659 Iout.n797 VGND 0.02471f
C10660 Iout.n798 VGND 0.04528f
C10661 Iout.t131 VGND 0.02185f
C10662 Iout.n799 VGND 0.04859f
C10663 Iout.n800 VGND 0.02471f
C10664 Iout.n801 VGND 0.04528f
C10665 Iout.t230 VGND 0.02185f
C10666 Iout.n802 VGND 0.04859f
C10667 Iout.n803 VGND 0.02471f
C10668 Iout.n804 VGND 0.04528f
C10669 Iout.t122 VGND 0.02185f
C10670 Iout.n805 VGND 0.04859f
C10671 Iout.n806 VGND 0.02471f
C10672 Iout.n807 VGND 0.04528f
C10673 Iout.t189 VGND 0.02185f
C10674 Iout.n808 VGND 0.04859f
C10675 Iout.n809 VGND 0.02471f
C10676 Iout.n810 VGND 0.04528f
C10677 Iout.t228 VGND 0.02185f
C10678 Iout.n811 VGND 0.04859f
C10679 Iout.n812 VGND 0.02471f
C10680 Iout.n813 VGND 0.04528f
C10681 Iout.t47 VGND 0.02185f
C10682 Iout.n814 VGND 0.04859f
C10683 Iout.n815 VGND 0.02471f
C10684 Iout.n816 VGND 0.04528f
C10685 Iout.t92 VGND 0.02185f
C10686 Iout.n817 VGND 0.04859f
C10687 Iout.n818 VGND 0.02471f
C10688 Iout.n819 VGND 0.04528f
C10689 Iout.t252 VGND 0.02185f
C10690 Iout.n820 VGND 0.04859f
C10691 Iout.n821 VGND 0.02471f
C10692 Iout.n822 VGND 0.04528f
C10693 Iout.t233 VGND 0.02185f
C10694 Iout.n823 VGND 0.04859f
C10695 Iout.n824 VGND 0.02471f
C10696 Iout.n825 VGND 0.04528f
C10697 Iout.n826 VGND 0.22693f
C10698 Iout.t163 VGND 0.02185f
C10699 Iout.n827 VGND 0.04859f
C10700 Iout.n828 VGND 0.02471f
C10701 Iout.n829 VGND 0.07746f
C10702 Iout.n830 VGND 0.47048f
C10703 Iout.n831 VGND 0.04528f
C10704 Iout.t116 VGND 0.02185f
C10705 Iout.n832 VGND 0.04859f
C10706 Iout.n833 VGND 0.02471f
C10707 Iout.t141 VGND 0.02185f
C10708 Iout.n834 VGND 0.04859f
C10709 Iout.n835 VGND 0.02471f
C10710 Iout.n836 VGND 0.04528f
C10711 Iout.n837 VGND 0.47048f
C10712 Iout.n838 VGND 0.07746f
C10713 Iout.t254 VGND 0.02185f
C10714 Iout.n839 VGND 0.04859f
C10715 Iout.n840 VGND 0.02471f
C10716 Iout.t158 VGND 0.02185f
C10717 Iout.n841 VGND 0.04859f
C10718 Iout.n842 VGND 0.02471f
C10719 Iout.n843 VGND 0.07746f
C10720 Iout.n844 VGND 0.47048f
C10721 Iout.n845 VGND 0.04528f
C10722 Iout.t70 VGND 0.02185f
C10723 Iout.n846 VGND 0.04859f
C10724 Iout.n847 VGND 0.02471f
C10725 Iout.t217 VGND 0.02185f
C10726 Iout.n848 VGND 0.04859f
C10727 Iout.n849 VGND 0.02471f
C10728 Iout.n850 VGND 0.04528f
C10729 Iout.n851 VGND 0.47048f
C10730 Iout.n852 VGND 0.07746f
C10731 Iout.t87 VGND 0.02185f
C10732 Iout.n853 VGND 0.04859f
C10733 Iout.n854 VGND 0.02471f
C10734 Iout.t43 VGND 0.02185f
C10735 Iout.n855 VGND 0.04859f
C10736 Iout.n856 VGND 0.02471f
C10737 Iout.n857 VGND 0.07746f
C10738 Iout.n858 VGND 0.47048f
C10739 Iout.n859 VGND 0.04528f
C10740 Iout.t149 VGND 0.02185f
C10741 Iout.n860 VGND 0.04859f
C10742 Iout.n861 VGND 0.02471f
C10743 Iout.t119 VGND 0.02185f
C10744 Iout.n862 VGND 0.04859f
C10745 Iout.n863 VGND 0.02471f
C10746 Iout.n864 VGND 0.04528f
C10747 Iout.n865 VGND 0.47048f
C10748 Iout.n866 VGND 0.07746f
C10749 Iout.t146 VGND 0.02185f
C10750 Iout.n867 VGND 0.04859f
C10751 Iout.n868 VGND 0.02471f
C10752 Iout.t253 VGND 0.02185f
C10753 Iout.n869 VGND 0.04859f
C10754 Iout.n870 VGND 0.02471f
C10755 Iout.n871 VGND 0.07746f
C10756 Iout.n872 VGND 0.47048f
C10757 Iout.n873 VGND 0.04528f
C10758 Iout.t241 VGND 0.02185f
C10759 Iout.n874 VGND 0.04859f
C10760 Iout.n875 VGND 0.02471f
C10761 Iout.t175 VGND 0.02185f
C10762 Iout.n876 VGND 0.04859f
C10763 Iout.n877 VGND 0.02471f
C10764 Iout.n878 VGND 0.04528f
C10765 Iout.n879 VGND 0.47048f
C10766 Iout.n880 VGND 0.07746f
C10767 Iout.t82 VGND 0.02185f
C10768 Iout.n881 VGND 0.04859f
C10769 Iout.n882 VGND 0.02471f
C10770 Iout.t68 VGND 0.02185f
C10771 Iout.n883 VGND 0.04859f
C10772 Iout.n884 VGND 0.02471f
C10773 Iout.n885 VGND 0.07746f
C10774 Iout.n886 VGND 0.47048f
C10775 Iout.n887 VGND 0.04528f
C10776 Iout.t60 VGND 0.02185f
C10777 Iout.n888 VGND 0.04859f
C10778 Iout.n889 VGND 0.02471f
C10779 Iout.t94 VGND 0.02185f
C10780 Iout.n890 VGND 0.04859f
C10781 Iout.n891 VGND 0.02471f
C10782 Iout.n892 VGND 0.04528f
C10783 Iout.n893 VGND 0.47048f
C10784 Iout.n894 VGND 0.07746f
C10785 Iout.t150 VGND 0.02185f
C10786 Iout.n895 VGND 0.04859f
C10787 Iout.n896 VGND 0.02471f
C10788 Iout.t246 VGND 0.02185f
C10789 Iout.n897 VGND 0.04859f
C10790 Iout.n898 VGND 0.02471f
C10791 Iout.n899 VGND 0.07746f
C10792 Iout.n900 VGND 0.47048f
C10793 Iout.n901 VGND 0.04528f
C10794 Iout.t38 VGND 0.02185f
C10795 Iout.n902 VGND 0.04859f
C10796 Iout.n903 VGND 0.02471f
C10797 Iout.t127 VGND 0.02185f
C10798 Iout.n904 VGND 0.04859f
C10799 Iout.n905 VGND 0.02471f
C10800 Iout.n906 VGND 0.04528f
C10801 Iout.n907 VGND 0.47048f
C10802 Iout.n908 VGND 0.07746f
C10803 Iout.t120 VGND 0.02185f
C10804 Iout.n909 VGND 0.04859f
C10805 Iout.n910 VGND 0.02471f
C10806 Iout.t251 VGND 0.02185f
C10807 Iout.n911 VGND 0.04859f
C10808 Iout.n912 VGND 0.02471f
C10809 Iout.n913 VGND 0.07746f
C10810 Iout.n914 VGND 0.47048f
C10811 Iout.n915 VGND 0.04528f
C10812 Iout.t215 VGND 0.02185f
C10813 Iout.n916 VGND 0.04859f
C10814 Iout.n917 VGND 0.02471f
C10815 Iout.t209 VGND 0.02185f
C10816 Iout.n918 VGND 0.04859f
C10817 Iout.n919 VGND 0.02471f
C10818 Iout.n920 VGND 0.04528f
C10819 Iout.n921 VGND 0.47048f
C10820 Iout.n922 VGND 0.07746f
C10821 Iout.t0 VGND 0.02185f
C10822 Iout.n923 VGND 0.04859f
C10823 Iout.n924 VGND 0.02471f
C10824 Iout.n925 VGND 0.07746f
C10825 Iout.t90 VGND 0.02185f
C10826 Iout.n926 VGND 0.04859f
C10827 Iout.n927 VGND 0.02471f
C10828 Iout.n928 VGND 0.07746f
C10829 Iout.n929 VGND 0.47048f
C10830 Iout.n930 VGND 0.04528f
C10831 Iout.t4 VGND 0.02185f
C10832 Iout.n931 VGND 0.04859f
C10833 Iout.n932 VGND 0.02471f
C10834 Iout.n933 VGND 0.04528f
C10835 Iout.t1 VGND 0.02185f
C10836 Iout.n934 VGND 0.04859f
C10837 Iout.n935 VGND 0.19196f
C10838 Iout.n936 VGND 2.51438f
C10839 Iout.n937 VGND 1.18657f
C10840 Iout.t221 VGND 0.02185f
C10841 Iout.n938 VGND 0.04859f
C10842 Iout.n939 VGND 0.19196f
C10843 Iout.n940 VGND 0.04528f
C10844 Iout.n941 VGND 0.22693f
C10845 Iout.n942 VGND 0.22693f
C10846 Iout.n943 VGND 0.04528f
C10847 Iout.t155 VGND 0.02185f
C10848 Iout.n944 VGND 0.04859f
C10849 Iout.n945 VGND 0.02471f
C10850 Iout.n946 VGND 0.04528f
C10851 Iout.n947 VGND 0.22693f
C10852 Iout.n948 VGND 0.22693f
C10853 Iout.n949 VGND 0.04528f
C10854 Iout.t196 VGND 0.02185f
C10855 Iout.n950 VGND 0.04859f
C10856 Iout.n951 VGND 0.02471f
C10857 Iout.n952 VGND 0.04528f
C10858 Iout.t227 VGND 0.02185f
C10859 Iout.n953 VGND 0.04859f
C10860 Iout.n954 VGND 0.19196f
C10861 Iout.n955 VGND 1.18657f
C10862 Iout.n956 VGND 1.18657f
C10863 Iout.t36 VGND 0.02185f
C10864 Iout.n957 VGND 0.04859f
C10865 Iout.n958 VGND 0.19196f
C10866 Iout.n959 VGND 0.04528f
C10867 Iout.n960 VGND 0.22693f
C10868 Iout.n961 VGND 0.22693f
C10869 Iout.n962 VGND 0.04528f
C10870 Iout.t142 VGND 0.02185f
C10871 Iout.n963 VGND 0.04859f
C10872 Iout.n964 VGND 0.02471f
C10873 Iout.n965 VGND 0.04528f
C10874 Iout.n966 VGND 0.22693f
C10875 Iout.n967 VGND 0.22693f
C10876 Iout.n968 VGND 0.04528f
C10877 Iout.t10 VGND 0.02185f
C10878 Iout.n969 VGND 0.04859f
C10879 Iout.n970 VGND 0.02471f
C10880 Iout.n971 VGND 0.04528f
C10881 Iout.t172 VGND 0.02185f
C10882 Iout.n972 VGND 0.04859f
C10883 Iout.n973 VGND 0.19196f
C10884 Iout.n974 VGND 1.18657f
C10885 Iout.n975 VGND 1.18657f
C10886 Iout.t201 VGND 0.02185f
C10887 Iout.n976 VGND 0.04859f
C10888 Iout.n977 VGND 0.19196f
C10889 Iout.n978 VGND 0.04528f
C10890 Iout.n979 VGND 0.22693f
C10891 Iout.n980 VGND 0.22693f
C10892 Iout.n981 VGND 0.04528f
C10893 Iout.t195 VGND 0.02185f
C10894 Iout.n982 VGND 0.04859f
C10895 Iout.n983 VGND 0.02471f
C10896 Iout.n984 VGND 0.04528f
C10897 Iout.n985 VGND 0.22693f
C10898 Iout.n986 VGND 0.22693f
C10899 Iout.n987 VGND 0.04528f
C10900 Iout.t250 VGND 0.02185f
C10901 Iout.n988 VGND 0.04859f
C10902 Iout.n989 VGND 0.02471f
C10903 Iout.n990 VGND 0.04528f
C10904 Iout.t8 VGND 0.02185f
C10905 Iout.n991 VGND 0.04859f
C10906 Iout.n992 VGND 0.19196f
C10907 Iout.n993 VGND 1.18657f
C10908 Iout.n994 VGND 1.18657f
C10909 Iout.t236 VGND 0.02185f
C10910 Iout.n995 VGND 0.04859f
C10911 Iout.n996 VGND 0.19196f
C10912 Iout.n997 VGND 0.04528f
C10913 Iout.n998 VGND 0.22693f
C10914 Iout.n999 VGND 0.22693f
C10915 Iout.n1000 VGND 0.04528f
C10916 Iout.t213 VGND 0.02185f
C10917 Iout.n1001 VGND 0.04859f
C10918 Iout.n1002 VGND 0.02471f
C10919 Iout.n1003 VGND 0.04528f
C10920 Iout.n1004 VGND 0.22693f
C10921 Iout.n1005 VGND 0.22693f
C10922 Iout.n1006 VGND 0.04528f
C10923 Iout.t63 VGND 0.02185f
C10924 Iout.n1007 VGND 0.04859f
C10925 Iout.n1008 VGND 0.02471f
C10926 Iout.n1009 VGND 0.04528f
C10927 Iout.t200 VGND 0.02185f
C10928 Iout.n1010 VGND 0.04859f
C10929 Iout.n1011 VGND 0.19196f
C10930 Iout.n1012 VGND 1.18657f
C10931 Iout.n1013 VGND 1.06545f
C10932 Iout.t54 VGND 0.02185f
C10933 Iout.n1014 VGND 0.04859f
C10934 Iout.n1015 VGND 0.19196f
C10935 Iout.n1016 VGND 0.04528f
C10936 Iout.n1017 VGND 0.22693f
C10937 Iout.n1018 VGND 0.13396f
C10938 Iout.n1019 VGND 0.04528f
C10939 Iout.t64 VGND 0.02185f
C10940 Iout.n1020 VGND 0.04859f
C10941 Iout.n1021 VGND 0.19196f
C10942 Iout.n1022 VGND 0.22043f
C10943 VPWR.n0 VGND 0.03902f
C10944 VPWR.t1414 VGND 0.24677f
C10945 VPWR.t1213 VGND 0.1092f
C10946 VPWR.t1417 VGND 0.31484f
C10947 VPWR.t1523 VGND 0.11913f
C10948 VPWR.t424 VGND 0.11913f
C10949 VPWR.t420 VGND 0.11913f
C10950 VPWR.t443 VGND 0.11913f
C10951 VPWR.t439 VGND 0.11913f
C10952 VPWR.t435 VGND 0.11913f
C10953 VPWR.t616 VGND 0.08368f
C10954 VPWR.n1 VGND 0.15203f
C10955 VPWR.n2 VGND 0.08044f
C10956 VPWR.t1214 VGND 0.04759f
C10957 VPWR.t617 VGND 0.01193f
C10958 VPWR.t436 VGND 0.01193f
C10959 VPWR.n4 VGND 0.02619f
C10960 VPWR.t440 VGND 0.01193f
C10961 VPWR.t444 VGND 0.01193f
C10962 VPWR.n5 VGND 0.02615f
C10963 VPWR.n6 VGND 0.0537f
C10964 VPWR.n7 VGND 0.15138f
C10965 VPWR.n8 VGND 0.04793f
C10966 VPWR.n9 VGND 0.0352f
C10967 VPWR.n10 VGND 0.0631f
C10968 VPWR.n12 VGND 0.01357f
C10969 VPWR.n13 VGND 0.01591f
C10970 VPWR.n14 VGND 0.02333f
C10971 VPWR.n15 VGND 0.07062f
C10972 VPWR.n16 VGND 0.01006f
C10973 VPWR.t1415 VGND 0.04758f
C10974 VPWR.n17 VGND 0.06119f
C10975 VPWR.n18 VGND 0.27944f
C10976 VPWR.n19 VGND 0.81484f
C10977 VPWR.n20 VGND 0.26524f
C10978 VPWR.n21 VGND 0.84572f
C10979 VPWR.n22 VGND 0.11562f
C10980 VPWR.t298 VGND 0.01021f
C10981 VPWR.n23 VGND 0.02493f
C10982 VPWR.n24 VGND 0.06622f
C10983 VPWR.t187 VGND 0.01021f
C10984 VPWR.n25 VGND 0.02493f
C10985 VPWR.n26 VGND 0.13327f
C10986 VPWR.t335 VGND 0.01021f
C10987 VPWR.n27 VGND 0.02493f
C10988 VPWR.n28 VGND 0.10618f
C10989 VPWR.t227 VGND 0.01021f
C10990 VPWR.n29 VGND 0.02493f
C10991 VPWR.n30 VGND 0.10618f
C10992 VPWR.t43 VGND 0.01021f
C10993 VPWR.n31 VGND 0.02493f
C10994 VPWR.n32 VGND 0.10618f
C10995 VPWR.t220 VGND 0.01021f
C10996 VPWR.n33 VGND 0.02493f
C10997 VPWR.n34 VGND 0.10618f
C10998 VPWR.t115 VGND 0.01021f
C10999 VPWR.n35 VGND 0.02493f
C11000 VPWR.n36 VGND 0.10618f
C11001 VPWR.t155 VGND 0.01021f
C11002 VPWR.n37 VGND 0.02493f
C11003 VPWR.n38 VGND 0.10618f
C11004 VPWR.t48 VGND 0.01021f
C11005 VPWR.n39 VGND 0.02493f
C11006 VPWR.n40 VGND 0.10618f
C11007 VPWR.t322 VGND 0.01021f
C11008 VPWR.n41 VGND 0.02493f
C11009 VPWR.n42 VGND 0.10618f
C11010 VPWR.t214 VGND 0.01021f
C11011 VPWR.n43 VGND 0.02493f
C11012 VPWR.n44 VGND 0.10618f
C11013 VPWR.t365 VGND 0.01021f
C11014 VPWR.n45 VGND 0.02493f
C11015 VPWR.n46 VGND 0.10618f
C11016 VPWR.t147 VGND 0.01021f
C11017 VPWR.n47 VGND 0.02493f
C11018 VPWR.n48 VGND 0.10618f
C11019 VPWR.t35 VGND 0.01021f
C11020 VPWR.n49 VGND 0.02493f
C11021 VPWR.n50 VGND 0.10618f
C11022 VPWR.t314 VGND 0.01021f
C11023 VPWR.n51 VGND 0.02493f
C11024 VPWR.n52 VGND 0.10618f
C11025 VPWR.t357 VGND 0.01021f
C11026 VPWR.n53 VGND 0.02493f
C11027 VPWR.n54 VGND 0.11497f
C11028 VPWR.n55 VGND 0.09598f
C11029 VPWR.t146 VGND 0.02774f
C11030 VPWR.t251 VGND 0.02465f
C11031 VPWR.n56 VGND 0.0762f
C11032 VPWR.t7 VGND 0.07675f
C11033 VPWR.t21 VGND 0.02774f
C11034 VPWR.t8 VGND 0.02465f
C11035 VPWR.n57 VGND 0.0762f
C11036 VPWR.n58 VGND 0.02861f
C11037 VPWR.n59 VGND 0.11584f
C11038 VPWR.n60 VGND 0.11584f
C11039 VPWR.n61 VGND 0.02861f
C11040 VPWR.t2 VGND 0.02774f
C11041 VPWR.t375 VGND 0.02465f
C11042 VPWR.n62 VGND 0.0762f
C11043 VPWR.t241 VGND 0.07675f
C11044 VPWR.t152 VGND 0.02774f
C11045 VPWR.t242 VGND 0.02465f
C11046 VPWR.n63 VGND 0.0762f
C11047 VPWR.n64 VGND 0.02861f
C11048 VPWR.n65 VGND 0.11584f
C11049 VPWR.n66 VGND 0.11584f
C11050 VPWR.n67 VGND 0.02861f
C11051 VPWR.t122 VGND 0.02774f
C11052 VPWR.t114 VGND 0.02465f
C11053 VPWR.n68 VGND 0.0762f
C11054 VPWR.t95 VGND 0.07675f
C11055 VPWR.t378 VGND 0.02774f
C11056 VPWR.t96 VGND 0.02465f
C11057 VPWR.n69 VGND 0.0762f
C11058 VPWR.n70 VGND 0.02861f
C11059 VPWR.n71 VGND 0.11584f
C11060 VPWR.n72 VGND 0.11584f
C11061 VPWR.n73 VGND 0.02861f
C11062 VPWR.t248 VGND 0.02774f
C11063 VPWR.t329 VGND 0.02465f
C11064 VPWR.n74 VGND 0.0762f
C11065 VPWR.t218 VGND 0.07675f
C11066 VPWR.t232 VGND 0.02774f
C11067 VPWR.t219 VGND 0.02465f
C11068 VPWR.n75 VGND 0.0762f
C11069 VPWR.n76 VGND 0.02861f
C11070 VPWR.n77 VGND 0.11584f
C11071 VPWR.n78 VGND 0.11584f
C11072 VPWR.n79 VGND 0.02861f
C11073 VPWR.t72 VGND 0.02774f
C11074 VPWR.t91 VGND 0.02465f
C11075 VPWR.n80 VGND 0.0762f
C11076 VPWR.t55 VGND 0.07675f
C11077 VPWR.t351 VGND 0.02774f
C11078 VPWR.t56 VGND 0.02465f
C11079 VPWR.n81 VGND 0.0762f
C11080 VPWR.n82 VGND 0.02861f
C11081 VPWR.n83 VGND 0.11584f
C11082 VPWR.n84 VGND 0.11584f
C11083 VPWR.n85 VGND 0.02861f
C11084 VPWR.t195 VGND 0.02774f
C11085 VPWR.t332 VGND 0.02465f
C11086 VPWR.n86 VGND 0.0762f
C11087 VPWR.t176 VGND 0.07675f
C11088 VPWR.t186 VGND 0.02774f
C11089 VPWR.t177 VGND 0.02465f
C11090 VPWR.n87 VGND 0.0762f
C11091 VPWR.n88 VGND 0.02861f
C11092 VPWR.n89 VGND 0.11584f
C11093 VPWR.n90 VGND 0.11584f
C11094 VPWR.n91 VGND 0.02861f
C11095 VPWR.t75 VGND 0.02774f
C11096 VPWR.t69 VGND 0.02465f
C11097 VPWR.n92 VGND 0.0762f
C11098 VPWR.t306 VGND 0.07675f
C11099 VPWR.t310 VGND 0.02774f
C11100 VPWR.t307 VGND 0.02465f
C11101 VPWR.n93 VGND 0.0762f
C11102 VPWR.n94 VGND 0.02861f
C11103 VPWR.n95 VGND 0.11584f
C11104 VPWR.n96 VGND 0.11584f
C11105 VPWR.n97 VGND 0.02861f
C11106 VPWR.t198 VGND 0.02774f
C11107 VPWR.t289 VGND 0.02465f
C11108 VPWR.n98 VGND 0.0762f
C11109 VPWR.t52 VGND 0.12083f
C11110 VPWR.t28 VGND 0.06535f
C11111 VPWR.t159 VGND 0.07675f
C11112 VPWR.t53 VGND 0.02774f
C11113 VPWR.t160 VGND 0.02465f
C11114 VPWR.n99 VGND 0.0762f
C11115 VPWR.t287 VGND 0.01021f
C11116 VPWR.n100 VGND 0.02492f
C11117 VPWR.n101 VGND 0.02734f
C11118 VPWR.n103 VGND 0.01517f
C11119 VPWR.t158 VGND 0.01021f
C11120 VPWR.n104 VGND 0.02492f
C11121 VPWR.n105 VGND 0.02734f
C11122 VPWR.t51 VGND 0.01018f
C11123 VPWR.n106 VGND 0.02594f
C11124 VPWR.n107 VGND 0.01639f
C11125 VPWR.t27 VGND 0.01033f
C11126 VPWR.n108 VGND 0.02304f
C11127 VPWR.n109 VGND 0.02346f
C11128 VPWR.n110 VGND 0.01479f
C11129 VPWR.n112 VGND 0.01517f
C11130 VPWR.n113 VGND 0.0221f
C11131 VPWR.t249 VGND 0.01021f
C11132 VPWR.n114 VGND 0.02492f
C11133 VPWR.n115 VGND 0.02734f
C11134 VPWR.t144 VGND 0.01018f
C11135 VPWR.n116 VGND 0.02594f
C11136 VPWR.n117 VGND 0.03075f
C11137 VPWR.t128 VGND 0.01033f
C11138 VPWR.n119 VGND 0.02304f
C11139 VPWR.n120 VGND 0.02346f
C11140 VPWR.n121 VGND 0.01479f
C11141 VPWR.n123 VGND 0.01517f
C11142 VPWR.n124 VGND 0.02116f
C11143 VPWR.t6 VGND 0.01021f
C11144 VPWR.n125 VGND 0.02492f
C11145 VPWR.n126 VGND 0.02734f
C11146 VPWR.t19 VGND 0.01018f
C11147 VPWR.n127 VGND 0.02594f
C11148 VPWR.n128 VGND 0.03075f
C11149 VPWR.t277 VGND 0.01033f
C11150 VPWR.n130 VGND 0.02304f
C11151 VPWR.n131 VGND 0.02346f
C11152 VPWR.n132 VGND 0.01479f
C11153 VPWR.n134 VGND 0.01517f
C11154 VPWR.n135 VGND 0.01985f
C11155 VPWR.n136 VGND 0.1762f
C11156 VPWR.t373 VGND 0.01021f
C11157 VPWR.n137 VGND 0.02492f
C11158 VPWR.n138 VGND 0.02734f
C11159 VPWR.t0 VGND 0.01018f
C11160 VPWR.n139 VGND 0.02594f
C11161 VPWR.n140 VGND 0.03075f
C11162 VPWR.t252 VGND 0.01033f
C11163 VPWR.n142 VGND 0.02304f
C11164 VPWR.n143 VGND 0.02346f
C11165 VPWR.n144 VGND 0.01479f
C11166 VPWR.n146 VGND 0.01517f
C11167 VPWR.n147 VGND 0.01985f
C11168 VPWR.n148 VGND 0.14641f
C11169 VPWR.t240 VGND 0.01021f
C11170 VPWR.n149 VGND 0.02492f
C11171 VPWR.n150 VGND 0.02734f
C11172 VPWR.t150 VGND 0.01018f
C11173 VPWR.n151 VGND 0.02594f
C11174 VPWR.n152 VGND 0.03075f
C11175 VPWR.t233 VGND 0.01033f
C11176 VPWR.n154 VGND 0.02304f
C11177 VPWR.n155 VGND 0.02346f
C11178 VPWR.n156 VGND 0.01479f
C11179 VPWR.n158 VGND 0.01517f
C11180 VPWR.n159 VGND 0.01985f
C11181 VPWR.n160 VGND 0.14641f
C11182 VPWR.t112 VGND 0.01021f
C11183 VPWR.n161 VGND 0.02492f
C11184 VPWR.n162 VGND 0.02734f
C11185 VPWR.t120 VGND 0.01018f
C11186 VPWR.n163 VGND 0.02594f
C11187 VPWR.n164 VGND 0.03075f
C11188 VPWR.t379 VGND 0.01033f
C11189 VPWR.n166 VGND 0.02304f
C11190 VPWR.n167 VGND 0.02346f
C11191 VPWR.n168 VGND 0.01479f
C11192 VPWR.n170 VGND 0.01517f
C11193 VPWR.n171 VGND 0.01985f
C11194 VPWR.n172 VGND 0.14641f
C11195 VPWR.t94 VGND 0.01021f
C11196 VPWR.n173 VGND 0.02492f
C11197 VPWR.n174 VGND 0.02734f
C11198 VPWR.t376 VGND 0.01018f
C11199 VPWR.n175 VGND 0.02594f
C11200 VPWR.n176 VGND 0.03075f
C11201 VPWR.t360 VGND 0.01033f
C11202 VPWR.n178 VGND 0.02304f
C11203 VPWR.n179 VGND 0.02346f
C11204 VPWR.n180 VGND 0.01479f
C11205 VPWR.n182 VGND 0.01517f
C11206 VPWR.n183 VGND 0.01985f
C11207 VPWR.n184 VGND 0.14641f
C11208 VPWR.t327 VGND 0.01021f
C11209 VPWR.n185 VGND 0.02492f
C11210 VPWR.n186 VGND 0.02734f
C11211 VPWR.t246 VGND 0.01018f
C11212 VPWR.n187 VGND 0.02594f
C11213 VPWR.n188 VGND 0.03075f
C11214 VPWR.t199 VGND 0.01033f
C11215 VPWR.n190 VGND 0.02304f
C11216 VPWR.n191 VGND 0.02346f
C11217 VPWR.n192 VGND 0.01479f
C11218 VPWR.n194 VGND 0.01517f
C11219 VPWR.n195 VGND 0.01985f
C11220 VPWR.n196 VGND 0.14641f
C11221 VPWR.t217 VGND 0.01021f
C11222 VPWR.n197 VGND 0.02492f
C11223 VPWR.n198 VGND 0.02734f
C11224 VPWR.t230 VGND 0.01018f
C11225 VPWR.n199 VGND 0.02594f
C11226 VPWR.n200 VGND 0.03075f
C11227 VPWR.t97 VGND 0.01033f
C11228 VPWR.n202 VGND 0.02304f
C11229 VPWR.n203 VGND 0.02346f
C11230 VPWR.n204 VGND 0.01479f
C11231 VPWR.n206 VGND 0.01517f
C11232 VPWR.n207 VGND 0.01985f
C11233 VPWR.n208 VGND 0.14641f
C11234 VPWR.t89 VGND 0.01021f
C11235 VPWR.n209 VGND 0.02492f
C11236 VPWR.n210 VGND 0.02734f
C11237 VPWR.t70 VGND 0.01018f
C11238 VPWR.n211 VGND 0.02594f
C11239 VPWR.n212 VGND 0.03075f
C11240 VPWR.t62 VGND 0.01033f
C11241 VPWR.n214 VGND 0.02304f
C11242 VPWR.n215 VGND 0.02346f
C11243 VPWR.n216 VGND 0.01479f
C11244 VPWR.n218 VGND 0.01517f
C11245 VPWR.n219 VGND 0.01985f
C11246 VPWR.n220 VGND 0.14641f
C11247 VPWR.t54 VGND 0.01021f
C11248 VPWR.n221 VGND 0.02492f
C11249 VPWR.n222 VGND 0.02734f
C11250 VPWR.t349 VGND 0.01018f
C11251 VPWR.n223 VGND 0.02594f
C11252 VPWR.n224 VGND 0.03075f
C11253 VPWR.t225 VGND 0.01033f
C11254 VPWR.n226 VGND 0.02304f
C11255 VPWR.n227 VGND 0.02346f
C11256 VPWR.n228 VGND 0.01479f
C11257 VPWR.n230 VGND 0.01517f
C11258 VPWR.n231 VGND 0.01985f
C11259 VPWR.n232 VGND 0.14641f
C11260 VPWR.t330 VGND 0.01021f
C11261 VPWR.n233 VGND 0.02492f
C11262 VPWR.n234 VGND 0.02734f
C11263 VPWR.t193 VGND 0.01018f
C11264 VPWR.n235 VGND 0.02594f
C11265 VPWR.n236 VGND 0.03075f
C11266 VPWR.t201 VGND 0.01033f
C11267 VPWR.n238 VGND 0.02304f
C11268 VPWR.n239 VGND 0.02346f
C11269 VPWR.n240 VGND 0.01479f
C11270 VPWR.n242 VGND 0.01517f
C11271 VPWR.n243 VGND 0.01985f
C11272 VPWR.n244 VGND 0.14641f
C11273 VPWR.t175 VGND 0.01021f
C11274 VPWR.n245 VGND 0.02492f
C11275 VPWR.n246 VGND 0.02734f
C11276 VPWR.t184 VGND 0.01018f
C11277 VPWR.n247 VGND 0.02594f
C11278 VPWR.n248 VGND 0.03075f
C11279 VPWR.t57 VGND 0.01033f
C11280 VPWR.n250 VGND 0.02304f
C11281 VPWR.n251 VGND 0.02346f
C11282 VPWR.n252 VGND 0.01479f
C11283 VPWR.n254 VGND 0.01517f
C11284 VPWR.n255 VGND 0.01985f
C11285 VPWR.n256 VGND 0.14641f
C11286 VPWR.t67 VGND 0.01021f
C11287 VPWR.n257 VGND 0.02492f
C11288 VPWR.n258 VGND 0.02734f
C11289 VPWR.t73 VGND 0.01018f
C11290 VPWR.n259 VGND 0.02594f
C11291 VPWR.n260 VGND 0.03075f
C11292 VPWR.t333 VGND 0.01033f
C11293 VPWR.n262 VGND 0.02304f
C11294 VPWR.n263 VGND 0.02346f
C11295 VPWR.n264 VGND 0.01479f
C11296 VPWR.n266 VGND 0.01517f
C11297 VPWR.n267 VGND 0.01985f
C11298 VPWR.n268 VGND 0.14641f
C11299 VPWR.t305 VGND 0.01021f
C11300 VPWR.n269 VGND 0.02492f
C11301 VPWR.n270 VGND 0.02734f
C11302 VPWR.t308 VGND 0.01018f
C11303 VPWR.n271 VGND 0.02594f
C11304 VPWR.n272 VGND 0.03075f
C11305 VPWR.t293 VGND 0.01033f
C11306 VPWR.n274 VGND 0.02304f
C11307 VPWR.n275 VGND 0.02346f
C11308 VPWR.n276 VGND 0.01479f
C11309 VPWR.n278 VGND 0.01517f
C11310 VPWR.n279 VGND 0.01985f
C11311 VPWR.n280 VGND 0.14641f
C11312 VPWR.n281 VGND 0.19753f
C11313 VPWR.n282 VGND 0.01985f
C11314 VPWR.n283 VGND 0.01479f
C11315 VPWR.t163 VGND 0.01033f
C11316 VPWR.n284 VGND 0.02304f
C11317 VPWR.n285 VGND 0.02346f
C11318 VPWR.t196 VGND 0.01018f
C11319 VPWR.n287 VGND 0.02594f
C11320 VPWR.n288 VGND 0.03075f
C11321 VPWR.n289 VGND 0.02861f
C11322 VPWR.t1118 VGND 0.02774f
C11323 VPWR.t1025 VGND 0.02465f
C11324 VPWR.n290 VGND 0.0762f
C11325 VPWR.t1117 VGND 0.12083f
C11326 VPWR.t1389 VGND 0.06535f
C11327 VPWR.t1024 VGND 0.07675f
C11328 VPWR.t601 VGND 0.02774f
C11329 VPWR.t359 VGND 0.02465f
C11330 VPWR.n291 VGND 0.0762f
C11331 VPWR.n292 VGND 0.01496f
C11332 VPWR.n293 VGND 0.06343f
C11333 VPWR.t358 VGND 0.11101f
C11334 VPWR.t1385 VGND 0.06535f
C11335 VPWR.t600 VGND 0.09955f
C11336 VPWR.t1361 VGND 0.02774f
C11337 VPWR.t773 VGND 0.02465f
C11338 VPWR.n294 VGND 0.0762f
C11339 VPWR.n295 VGND 0.01496f
C11340 VPWR.n297 VGND 0.0901f
C11341 VPWR.t772 VGND 0.07675f
C11342 VPWR.t1887 VGND 0.06535f
C11343 VPWR.t1360 VGND 0.09955f
C11344 VPWR.t1712 VGND 0.02774f
C11345 VPWR.t742 VGND 0.02465f
C11346 VPWR.n298 VGND 0.0762f
C11347 VPWR.n299 VGND 0.01496f
C11348 VPWR.n301 VGND 0.0901f
C11349 VPWR.t741 VGND 0.07675f
C11350 VPWR.t987 VGND 0.06535f
C11351 VPWR.t1711 VGND 0.09955f
C11352 VPWR.t1261 VGND 0.02774f
C11353 VPWR.t1915 VGND 0.02465f
C11354 VPWR.n302 VGND 0.0762f
C11355 VPWR.n303 VGND 0.01496f
C11356 VPWR.n305 VGND 0.0901f
C11357 VPWR.t1914 VGND 0.07675f
C11358 VPWR.t988 VGND 0.06535f
C11359 VPWR.t1260 VGND 0.09955f
C11360 VPWR.t1313 VGND 0.02774f
C11361 VPWR.t1255 VGND 0.02465f
C11362 VPWR.n306 VGND 0.0762f
C11363 VPWR.n307 VGND 0.01496f
C11364 VPWR.n309 VGND 0.0901f
C11365 VPWR.t1254 VGND 0.07675f
C11366 VPWR.t1883 VGND 0.06535f
C11367 VPWR.t1312 VGND 0.09955f
C11368 VPWR.t1231 VGND 0.02774f
C11369 VPWR.t1319 VGND 0.02465f
C11370 VPWR.n310 VGND 0.0762f
C11371 VPWR.n311 VGND 0.01496f
C11372 VPWR.n313 VGND 0.0901f
C11373 VPWR.t1318 VGND 0.07675f
C11374 VPWR.t1884 VGND 0.06535f
C11375 VPWR.t1230 VGND 0.09955f
C11376 VPWR.t842 VGND 0.02774f
C11377 VPWR.t1241 VGND 0.02465f
C11378 VPWR.n314 VGND 0.0762f
C11379 VPWR.n315 VGND 0.01496f
C11380 VPWR.n317 VGND 0.0901f
C11381 VPWR.t1240 VGND 0.07675f
C11382 VPWR.t991 VGND 0.06535f
C11383 VPWR.t841 VGND 0.09955f
C11384 VPWR.t836 VGND 0.02774f
C11385 VPWR.t944 VGND 0.02465f
C11386 VPWR.n318 VGND 0.0762f
C11387 VPWR.n319 VGND 0.01496f
C11388 VPWR.n321 VGND 0.0901f
C11389 VPWR.t943 VGND 0.07675f
C11390 VPWR.t1386 VGND 0.06535f
C11391 VPWR.t835 VGND 0.09955f
C11392 VPWR.t803 VGND 0.02774f
C11393 VPWR.t651 VGND 0.02465f
C11394 VPWR.n322 VGND 0.0762f
C11395 VPWR.n323 VGND 0.01496f
C11396 VPWR.n325 VGND 0.0901f
C11397 VPWR.t650 VGND 0.07675f
C11398 VPWR.t1387 VGND 0.06535f
C11399 VPWR.t802 VGND 0.09955f
C11400 VPWR.t1148 VGND 0.02774f
C11401 VPWR.t809 VGND 0.02465f
C11402 VPWR.n326 VGND 0.0762f
C11403 VPWR.n327 VGND 0.01496f
C11404 VPWR.n329 VGND 0.0901f
C11405 VPWR.t808 VGND 0.07675f
C11406 VPWR.t989 VGND 0.06535f
C11407 VPWR.t1147 VGND 0.09955f
C11408 VPWR.t1338 VGND 0.02774f
C11409 VPWR.t1154 VGND 0.02465f
C11410 VPWR.n330 VGND 0.0762f
C11411 VPWR.n331 VGND 0.01496f
C11412 VPWR.n333 VGND 0.0901f
C11413 VPWR.t1153 VGND 0.07675f
C11414 VPWR.t990 VGND 0.06535f
C11415 VPWR.t1337 VGND 0.09955f
C11416 VPWR.t393 VGND 0.02774f
C11417 VPWR.t1544 VGND 0.02465f
C11418 VPWR.n334 VGND 0.0762f
C11419 VPWR.n335 VGND 0.01496f
C11420 VPWR.n337 VGND 0.0901f
C11421 VPWR.t1543 VGND 0.07675f
C11422 VPWR.t1388 VGND 0.06535f
C11423 VPWR.t392 VGND 0.09955f
C11424 VPWR.t1467 VGND 0.02774f
C11425 VPWR.t1267 VGND 0.02465f
C11426 VPWR.n338 VGND 0.0762f
C11427 VPWR.n339 VGND 0.01496f
C11428 VPWR.n341 VGND 0.0901f
C11429 VPWR.t1266 VGND 0.07675f
C11430 VPWR.t1885 VGND 0.06535f
C11431 VPWR.t1466 VGND 0.09955f
C11432 VPWR.t1677 VGND 0.02774f
C11433 VPWR.t1443 VGND 0.02465f
C11434 VPWR.n342 VGND 0.0762f
C11435 VPWR.n343 VGND 0.01496f
C11436 VPWR.n345 VGND 0.0901f
C11437 VPWR.t1442 VGND 0.07675f
C11438 VPWR.t1886 VGND 0.06535f
C11439 VPWR.t1676 VGND 0.09955f
C11440 VPWR.t1204 VGND 0.02774f
C11441 VPWR.t470 VGND 0.02465f
C11442 VPWR.n346 VGND 0.0762f
C11443 VPWR.n347 VGND 0.01496f
C11444 VPWR.n349 VGND 0.0901f
C11445 VPWR.t469 VGND 0.07675f
C11446 VPWR.t1384 VGND 0.06535f
C11447 VPWR.t1203 VGND 0.09955f
C11448 VPWR.n350 VGND 0.0901f
C11449 VPWR.n352 VGND 0.01496f
C11450 VPWR.n353 VGND 0.11584f
C11451 VPWR.n354 VGND 0.84042f
C11452 VPWR.n355 VGND 0.11584f
C11453 VPWR.t1112 VGND 0.02774f
C11454 VPWR.t1200 VGND 0.02465f
C11455 VPWR.n356 VGND 0.0762f
C11456 VPWR.t1111 VGND 0.12083f
C11457 VPWR.t1169 VGND 0.06535f
C11458 VPWR.t1199 VGND 0.07675f
C11459 VPWR.t473 VGND 0.09955f
C11460 VPWR.t1021 VGND 0.02774f
C11461 VPWR.t1562 VGND 0.02465f
C11462 VPWR.n357 VGND 0.0762f
C11463 VPWR.n358 VGND 0.11584f
C11464 VPWR.n359 VGND 0.11584f
C11465 VPWR.t474 VGND 0.02774f
C11466 VPWR.t1435 VGND 0.02465f
C11467 VPWR.n360 VGND 0.0762f
C11468 VPWR.t763 VGND 0.06535f
C11469 VPWR.t1434 VGND 0.07675f
C11470 VPWR.t1514 VGND 0.09955f
C11471 VPWR.t1459 VGND 0.02774f
C11472 VPWR.t1279 VGND 0.02465f
C11473 VPWR.n361 VGND 0.0762f
C11474 VPWR.n362 VGND 0.11584f
C11475 VPWR.n363 VGND 0.11584f
C11476 VPWR.t1515 VGND 0.02774f
C11477 VPWR.t589 VGND 0.02465f
C11478 VPWR.n364 VGND 0.0762f
C11479 VPWR.t1168 VGND 0.06535f
C11480 VPWR.t588 VGND 0.07675f
C11481 VPWR.t1134 VGND 0.09955f
C11482 VPWR.t1548 VGND 0.02774f
C11483 VPWR.t1141 VGND 0.02465f
C11484 VPWR.n365 VGND 0.0762f
C11485 VPWR.n366 VGND 0.11584f
C11486 VPWR.n367 VGND 0.11584f
C11487 VPWR.t1135 VGND 0.02774f
C11488 VPWR.t819 VGND 0.02465f
C11489 VPWR.n368 VGND 0.0762f
C11490 VPWR.t1218 VGND 0.06535f
C11491 VPWR.t818 VGND 0.07675f
C11492 VPWR.t934 VGND 0.09955f
C11493 VPWR.t813 VGND 0.02774f
C11494 VPWR.t895 VGND 0.02465f
C11495 VPWR.n369 VGND 0.0762f
C11496 VPWR.n370 VGND 0.11584f
C11497 VPWR.n371 VGND 0.11584f
C11498 VPWR.t935 VGND 0.02774f
C11499 VPWR.t555 VGND 0.02465f
C11500 VPWR.n372 VGND 0.0762f
C11501 VPWR.t1166 VGND 0.06535f
C11502 VPWR.t554 VGND 0.07675f
C11503 VPWR.t1236 VGND 0.09955f
C11504 VPWR.t948 VGND 0.02774f
C11505 VPWR.t1871 VGND 0.02465f
C11506 VPWR.n373 VGND 0.0762f
C11507 VPWR.n374 VGND 0.11584f
C11508 VPWR.n375 VGND 0.11584f
C11509 VPWR.t1237 VGND 0.02774f
C11510 VPWR.t1344 VGND 0.02465f
C11511 VPWR.n376 VGND 0.0762f
C11512 VPWR.t920 VGND 0.06535f
C11513 VPWR.t1343 VGND 0.07675f
C11514 VPWR.t1250 VGND 0.09955f
C11515 VPWR.t1323 VGND 0.02774f
C11516 VPWR.t1841 VGND 0.02465f
C11517 VPWR.n377 VGND 0.0762f
C11518 VPWR.n378 VGND 0.11584f
C11519 VPWR.n379 VGND 0.11584f
C11520 VPWR.t1251 VGND 0.02774f
C11521 VPWR.t1925 VGND 0.02465f
C11522 VPWR.n380 VGND 0.0762f
C11523 VPWR.t766 VGND 0.06535f
C11524 VPWR.t1924 VGND 0.07675f
C11525 VPWR.t737 VGND 0.09955f
C11526 VPWR.t1718 VGND 0.02774f
C11527 VPWR.t762 VGND 0.02465f
C11528 VPWR.n381 VGND 0.0762f
C11529 VPWR.n382 VGND 0.11584f
C11530 VPWR.n383 VGND 0.11584f
C11531 VPWR.t738 VGND 0.02774f
C11532 VPWR.t785 VGND 0.02465f
C11533 VPWR.n384 VGND 0.0762f
C11534 VPWR.t764 VGND 0.06535f
C11535 VPWR.t784 VGND 0.07675f
C11536 VPWR.t609 VGND 0.02774f
C11537 VPWR.t316 VGND 0.02465f
C11538 VPWR.n385 VGND 0.0762f
C11539 VPWR.t529 VGND 0.02774f
C11540 VPWR.t37 VGND 0.02465f
C11541 VPWR.n386 VGND 0.0762f
C11542 VPWR.t1121 VGND 0.12083f
C11543 VPWR.t1433 VGND 0.06535f
C11544 VPWR.t973 VGND 0.07675f
C11545 VPWR.t1122 VGND 0.02774f
C11546 VPWR.t974 VGND 0.02465f
C11547 VPWR.n387 VGND 0.0762f
C11548 VPWR.n388 VGND 0.01496f
C11549 VPWR.n390 VGND 0.0901f
C11550 VPWR.t828 VGND 0.09955f
C11551 VPWR.t1347 VGND 0.06535f
C11552 VPWR.t837 VGND 0.07675f
C11553 VPWR.t829 VGND 0.02774f
C11554 VPWR.t838 VGND 0.02465f
C11555 VPWR.n391 VGND 0.0762f
C11556 VPWR.n392 VGND 0.01496f
C11557 VPWR.n394 VGND 0.0901f
C11558 VPWR.t1555 VGND 0.09955f
C11559 VPWR.t1650 VGND 0.06535f
C11560 VPWR.t1452 VGND 0.07675f
C11561 VPWR.t1556 VGND 0.02774f
C11562 VPWR.t1453 VGND 0.02465f
C11563 VPWR.n395 VGND 0.0762f
C11564 VPWR.n396 VGND 0.01496f
C11565 VPWR.n398 VGND 0.0901f
C11566 VPWR.t1478 VGND 0.09955f
C11567 VPWR.t1649 VGND 0.06535f
C11568 VPWR.t1518 VGND 0.07675f
C11569 VPWR.t1479 VGND 0.02774f
C11570 VPWR.t1519 VGND 0.02465f
C11571 VPWR.n399 VGND 0.0762f
C11572 VPWR.n400 VGND 0.01496f
C11573 VPWR.n402 VGND 0.0901f
C11574 VPWR.t1394 VGND 0.09955f
C11575 VPWR.t1432 VGND 0.06535f
C11576 VPWR.t1639 VGND 0.07675f
C11577 VPWR.t1395 VGND 0.02774f
C11578 VPWR.t1640 VGND 0.02465f
C11579 VPWR.n403 VGND 0.0762f
C11580 VPWR.n404 VGND 0.01496f
C11581 VPWR.n406 VGND 0.0901f
C11582 VPWR.t1333 VGND 0.09955f
C11583 VPWR.t1655 VGND 0.06535f
C11584 VPWR.t630 VGND 0.07675f
C11585 VPWR.t1334 VGND 0.02774f
C11586 VPWR.t631 VGND 0.02465f
C11587 VPWR.n407 VGND 0.0762f
C11588 VPWR.n408 VGND 0.01496f
C11589 VPWR.n410 VGND 0.0901f
C11590 VPWR.t624 VGND 0.09955f
C11591 VPWR.t1654 VGND 0.06535f
C11592 VPWR.t798 VGND 0.07675f
C11593 VPWR.t625 VGND 0.02774f
C11594 VPWR.t799 VGND 0.02465f
C11595 VPWR.n411 VGND 0.0762f
C11596 VPWR.n412 VGND 0.01496f
C11597 VPWR.n414 VGND 0.0901f
C11598 VPWR.t792 VGND 0.09955f
C11599 VPWR.t1431 VGND 0.06535f
C11600 VPWR.t400 VGND 0.07675f
C11601 VPWR.t793 VGND 0.02774f
C11602 VPWR.t401 VGND 0.02465f
C11603 VPWR.n415 VGND 0.0762f
C11604 VPWR.n416 VGND 0.01496f
C11605 VPWR.n418 VGND 0.0901f
C11606 VPWR.t658 VGND 0.09955f
C11607 VPWR.t1430 VGND 0.06535f
C11608 VPWR.t699 VGND 0.07675f
C11609 VPWR.t659 VGND 0.02774f
C11610 VPWR.t700 VGND 0.02465f
C11611 VPWR.n419 VGND 0.0762f
C11612 VPWR.n420 VGND 0.01496f
C11613 VPWR.n422 VGND 0.0901f
C11614 VPWR.t548 VGND 0.09955f
C11615 VPWR.t1656 VGND 0.06535f
C11616 VPWR.t516 VGND 0.07675f
C11617 VPWR.t549 VGND 0.02774f
C11618 VPWR.t517 VGND 0.02465f
C11619 VPWR.n423 VGND 0.0762f
C11620 VPWR.n424 VGND 0.01496f
C11621 VPWR.n426 VGND 0.0901f
C11622 VPWR.t510 VGND 0.09955f
C11623 VPWR.t1648 VGND 0.06535f
C11624 VPWR.t926 VGND 0.07675f
C11625 VPWR.t511 VGND 0.02774f
C11626 VPWR.t927 VGND 0.02465f
C11627 VPWR.n427 VGND 0.0762f
C11628 VPWR.n428 VGND 0.01496f
C11629 VPWR.n430 VGND 0.0901f
C11630 VPWR.t1668 VGND 0.09955f
C11631 VPWR.t1647 VGND 0.06535f
C11632 VPWR.t1356 VGND 0.07675f
C11633 VPWR.t1669 VGND 0.02774f
C11634 VPWR.t1357 VGND 0.02465f
C11635 VPWR.n431 VGND 0.0762f
C11636 VPWR.n432 VGND 0.01496f
C11637 VPWR.n434 VGND 0.0901f
C11638 VPWR.t1286 VGND 0.09955f
C11639 VPWR.t1653 VGND 0.06535f
C11640 VPWR.t1723 VGND 0.07675f
C11641 VPWR.t1287 VGND 0.02774f
C11642 VPWR.t1724 VGND 0.02465f
C11643 VPWR.n435 VGND 0.0762f
C11644 VPWR.n436 VGND 0.01496f
C11645 VPWR.n438 VGND 0.0901f
C11646 VPWR.t1300 VGND 0.09955f
C11647 VPWR.t1652 VGND 0.06535f
C11648 VPWR.t1372 VGND 0.07675f
C11649 VPWR.t1301 VGND 0.02774f
C11650 VPWR.t1373 VGND 0.02465f
C11651 VPWR.n439 VGND 0.0762f
C11652 VPWR.n440 VGND 0.01496f
C11653 VPWR.n442 VGND 0.0901f
C11654 VPWR.t1500 VGND 0.09955f
C11655 VPWR.t1651 VGND 0.06535f
C11656 VPWR.t612 VGND 0.07675f
C11657 VPWR.t1501 VGND 0.02774f
C11658 VPWR.t613 VGND 0.02465f
C11659 VPWR.n443 VGND 0.0762f
C11660 VPWR.n444 VGND 0.01496f
C11661 VPWR.n446 VGND 0.0901f
C11662 VPWR.t528 VGND 0.09955f
C11663 VPWR.t1429 VGND 0.06535f
C11664 VPWR.t36 VGND 0.11101f
C11665 VPWR.n447 VGND 0.06343f
C11666 VPWR.n448 VGND 0.01496f
C11667 VPWR.n449 VGND 0.11584f
C11668 VPWR.n450 VGND 0.84572f
C11669 VPWR.n451 VGND 0.11584f
C11670 VPWR.t1847 VGND 0.02774f
C11671 VPWR.t149 VGND 0.02465f
C11672 VPWR.n452 VGND 0.0762f
C11673 VPWR.t530 VGND 0.07675f
C11674 VPWR.t413 VGND 0.02774f
C11675 VPWR.t531 VGND 0.02465f
C11676 VPWR.n453 VGND 0.0762f
C11677 VPWR.n454 VGND 0.11584f
C11678 VPWR.n455 VGND 0.11584f
C11679 VPWR.t1078 VGND 0.02774f
C11680 VPWR.t1880 VGND 0.02465f
C11681 VPWR.n456 VGND 0.0762f
C11682 VPWR.t1304 VGND 0.07675f
C11683 VPWR.t1574 VGND 0.02774f
C11684 VPWR.t1305 VGND 0.02465f
C11685 VPWR.n457 VGND 0.0762f
C11686 VPWR.n458 VGND 0.11584f
C11687 VPWR.n459 VGND 0.11584f
C11688 VPWR.t1606 VGND 0.02774f
C11689 VPWR.t1570 VGND 0.02465f
C11690 VPWR.n460 VGND 0.0762f
C11691 VPWR.t1609 VGND 0.07675f
C11692 VPWR.t746 VGND 0.02774f
C11693 VPWR.t1610 VGND 0.02465f
C11694 VPWR.n461 VGND 0.0762f
C11695 VPWR.n462 VGND 0.11584f
C11696 VPWR.n463 VGND 0.11584f
C11697 VPWR.t1685 VGND 0.02774f
C11698 VPWR.t754 VGND 0.02465f
C11699 VPWR.n464 VGND 0.0762f
C11700 VPWR.t1032 VGND 0.07675f
C11701 VPWR.t901 VGND 0.02774f
C11702 VPWR.t1033 VGND 0.02465f
C11703 VPWR.n465 VGND 0.0762f
C11704 VPWR.n466 VGND 0.11584f
C11705 VPWR.n467 VGND 0.11584f
C11706 VPWR.t1580 VGND 0.02774f
C11707 VPWR.t663 VGND 0.02465f
C11708 VPWR.n468 VGND 0.0762f
C11709 VPWR.t1583 VGND 0.07675f
C11710 VPWR.t960 VGND 0.02774f
C11711 VPWR.t1584 VGND 0.02465f
C11712 VPWR.n469 VGND 0.0762f
C11713 VPWR.n470 VGND 0.11584f
C11714 VPWR.n471 VGND 0.11584f
C11715 VPWR.t1596 VGND 0.02774f
C11716 VPWR.t653 VGND 0.02465f
C11717 VPWR.n472 VGND 0.0762f
C11718 VPWR.t1623 VGND 0.07675f
C11719 VPWR.t1509 VGND 0.02774f
C11720 VPWR.t1624 VGND 0.02465f
C11721 VPWR.n473 VGND 0.0762f
C11722 VPWR.n474 VGND 0.11584f
C11723 VPWR.n475 VGND 0.11584f
C11724 VPWR.t1493 VGND 0.02774f
C11725 VPWR.t1397 VGND 0.02465f
C11726 VPWR.n476 VGND 0.0762f
C11727 VPWR.t1472 VGND 0.07675f
C11728 VPWR.t690 VGND 0.02774f
C11729 VPWR.t1473 VGND 0.02465f
C11730 VPWR.n477 VGND 0.0762f
C11731 VPWR.n478 VGND 0.11584f
C11732 VPWR.n479 VGND 0.11584f
C11733 VPWR.t1192 VGND 0.02774f
C11734 VPWR.t1027 VGND 0.02465f
C11735 VPWR.n480 VGND 0.0762f
C11736 VPWR.t1130 VGND 0.12083f
C11737 VPWR.t769 VGND 0.06535f
C11738 VPWR.t1014 VGND 0.07675f
C11739 VPWR.t1131 VGND 0.02774f
C11740 VPWR.t1015 VGND 0.02465f
C11741 VPWR.n481 VGND 0.0762f
C11742 VPWR.t1120 VGND 0.02774f
C11743 VPWR.t1023 VGND 0.02465f
C11744 VPWR.n482 VGND 0.0762f
C11745 VPWR.t1119 VGND 0.12083f
C11746 VPWR.t1867 VGND 0.06535f
C11747 VPWR.t1022 VGND 0.07675f
C11748 VPWR.t599 VGND 0.02774f
C11749 VPWR.t367 VGND 0.02465f
C11750 VPWR.n483 VGND 0.0762f
C11751 VPWR.n484 VGND 0.01496f
C11752 VPWR.n485 VGND 0.06343f
C11753 VPWR.t366 VGND 0.11101f
C11754 VPWR.t978 VGND 0.06535f
C11755 VPWR.t598 VGND 0.09955f
C11756 VPWR.t1359 VGND 0.02774f
C11757 VPWR.t771 VGND 0.02465f
C11758 VPWR.n486 VGND 0.0762f
C11759 VPWR.n487 VGND 0.01496f
C11760 VPWR.n489 VGND 0.0901f
C11761 VPWR.t770 VGND 0.07675f
C11762 VPWR.t1378 VGND 0.06535f
C11763 VPWR.t1358 VGND 0.09955f
C11764 VPWR.t1307 VGND 0.02774f
C11765 VPWR.t740 VGND 0.02465f
C11766 VPWR.n490 VGND 0.0762f
C11767 VPWR.n491 VGND 0.01496f
C11768 VPWR.n493 VGND 0.0901f
C11769 VPWR.t739 VGND 0.07675f
C11770 VPWR.t1657 VGND 0.06535f
C11771 VPWR.t1306 VGND 0.09955f
C11772 VPWR.t1259 VGND 0.02774f
C11773 VPWR.t1911 VGND 0.02465f
C11774 VPWR.n494 VGND 0.0762f
C11775 VPWR.n495 VGND 0.01496f
C11776 VPWR.n497 VGND 0.0901f
C11777 VPWR.t1910 VGND 0.07675f
C11778 VPWR.t1658 VGND 0.06535f
C11779 VPWR.t1258 VGND 0.09955f
C11780 VPWR.t1311 VGND 0.02774f
C11781 VPWR.t1253 VGND 0.02465f
C11782 VPWR.n498 VGND 0.0762f
C11783 VPWR.n499 VGND 0.01496f
C11784 VPWR.n501 VGND 0.0901f
C11785 VPWR.t1252 VGND 0.07675f
C11786 VPWR.t1868 VGND 0.06535f
C11787 VPWR.t1310 VGND 0.09955f
C11788 VPWR.t519 VGND 0.02774f
C11789 VPWR.t1315 VGND 0.02465f
C11790 VPWR.n502 VGND 0.0762f
C11791 VPWR.n503 VGND 0.01496f
C11792 VPWR.n505 VGND 0.0901f
C11793 VPWR.t1314 VGND 0.07675f
C11794 VPWR.t1375 VGND 0.06535f
C11795 VPWR.t518 VGND 0.09955f
C11796 VPWR.t840 VGND 0.02774f
C11797 VPWR.t1239 VGND 0.02465f
C11798 VPWR.n506 VGND 0.0762f
C11799 VPWR.n507 VGND 0.01496f
C11800 VPWR.n509 VGND 0.0901f
C11801 VPWR.t1238 VGND 0.07675f
C11802 VPWR.t1661 VGND 0.06535f
C11803 VPWR.t839 VGND 0.09955f
C11804 VPWR.t832 VGND 0.02774f
C11805 VPWR.t844 VGND 0.02465f
C11806 VPWR.n510 VGND 0.0762f
C11807 VPWR.n511 VGND 0.01496f
C11808 VPWR.n513 VGND 0.0901f
C11809 VPWR.t843 VGND 0.07675f
C11810 VPWR.t979 VGND 0.06535f
C11811 VPWR.t831 VGND 0.09955f
C11812 VPWR.t801 VGND 0.02774f
C11813 VPWR.t647 VGND 0.02465f
C11814 VPWR.n514 VGND 0.0762f
C11815 VPWR.n515 VGND 0.01496f
C11816 VPWR.n517 VGND 0.0901f
C11817 VPWR.t646 VGND 0.07675f
C11818 VPWR.t1865 VGND 0.06535f
C11819 VPWR.t800 VGND 0.09955f
C11820 VPWR.t1146 VGND 0.02774f
C11821 VPWR.t805 VGND 0.02465f
C11822 VPWR.n518 VGND 0.0762f
C11823 VPWR.n519 VGND 0.01496f
C11824 VPWR.n521 VGND 0.0901f
C11825 VPWR.t804 VGND 0.07675f
C11826 VPWR.t1659 VGND 0.06535f
C11827 VPWR.t1145 VGND 0.09955f
C11828 VPWR.t1336 VGND 0.02774f
C11829 VPWR.t1150 VGND 0.02465f
C11830 VPWR.n522 VGND 0.0762f
C11831 VPWR.n523 VGND 0.01496f
C11832 VPWR.n525 VGND 0.0901f
C11833 VPWR.t1149 VGND 0.07675f
C11834 VPWR.t1660 VGND 0.06535f
C11835 VPWR.t1335 VGND 0.09955f
C11836 VPWR.t391 VGND 0.02774f
C11837 VPWR.t1540 VGND 0.02465f
C11838 VPWR.n526 VGND 0.0762f
C11839 VPWR.n527 VGND 0.01496f
C11840 VPWR.n529 VGND 0.0901f
C11841 VPWR.t1539 VGND 0.07675f
C11842 VPWR.t1866 VGND 0.06535f
C11843 VPWR.t390 VGND 0.09955f
C11844 VPWR.t1471 VGND 0.02774f
C11845 VPWR.t1265 VGND 0.02465f
C11846 VPWR.n530 VGND 0.0762f
C11847 VPWR.n531 VGND 0.01496f
C11848 VPWR.n533 VGND 0.0901f
C11849 VPWR.t1264 VGND 0.07675f
C11850 VPWR.t1376 VGND 0.06535f
C11851 VPWR.t1470 VGND 0.09955f
C11852 VPWR.t1675 VGND 0.02774f
C11853 VPWR.t1445 VGND 0.02465f
C11854 VPWR.n534 VGND 0.0762f
C11855 VPWR.n535 VGND 0.01496f
C11856 VPWR.n537 VGND 0.0901f
C11857 VPWR.t1444 VGND 0.07675f
C11858 VPWR.t1377 VGND 0.06535f
C11859 VPWR.t1674 VGND 0.09955f
C11860 VPWR.t1202 VGND 0.02774f
C11861 VPWR.t1679 VGND 0.02465f
C11862 VPWR.n538 VGND 0.0762f
C11863 VPWR.n539 VGND 0.01496f
C11864 VPWR.n541 VGND 0.0901f
C11865 VPWR.t1678 VGND 0.07675f
C11866 VPWR.t977 VGND 0.06535f
C11867 VPWR.t1201 VGND 0.09955f
C11868 VPWR.n542 VGND 0.0901f
C11869 VPWR.n544 VGND 0.01496f
C11870 VPWR.n545 VGND 0.11584f
C11871 VPWR.n546 VGND 0.84042f
C11872 VPWR.n547 VGND 0.11584f
C11873 VPWR.t1106 VGND 0.02774f
C11874 VPWR.t861 VGND 0.02465f
C11875 VPWR.n548 VGND 0.0762f
C11876 VPWR.t1105 VGND 0.12083f
C11877 VPWR.t1263 VGND 0.06535f
C11878 VPWR.t860 VGND 0.07675f
C11879 VPWR.t1709 VGND 0.09955f
C11880 VPWR.t853 VGND 0.02774f
C11881 VPWR.t1903 VGND 0.02465f
C11882 VPWR.n549 VGND 0.0762f
C11883 VPWR.n550 VGND 0.11584f
C11884 VPWR.n551 VGND 0.11584f
C11885 VPWR.t1710 VGND 0.02774f
C11886 VPWR.t1485 VGND 0.02465f
C11887 VPWR.n552 VGND 0.0762f
C11888 VPWR.t1644 VGND 0.06535f
C11889 VPWR.t1484 VGND 0.07675f
C11890 VPWR.t1274 VGND 0.09955f
C11891 VPWR.t1447 VGND 0.02774f
C11892 VPWR.t995 VGND 0.02465f
C11893 VPWR.n553 VGND 0.0762f
C11894 VPWR.n554 VGND 0.11584f
C11895 VPWR.n555 VGND 0.11584f
C11896 VPWR.t1275 VGND 0.02774f
C11897 VPWR.t1704 VGND 0.02465f
C11898 VPWR.n556 VGND 0.0762f
C11899 VPWR.t1262 VGND 0.06535f
C11900 VPWR.t1703 VGND 0.07675f
C11901 VPWR.t911 VGND 0.09955f
C11902 VPWR.t1696 VGND 0.02774f
C11903 VPWR.t954 VGND 0.02465f
C11904 VPWR.n557 VGND 0.0762f
C11905 VPWR.n558 VGND 0.11584f
C11906 VPWR.n559 VGND 0.11584f
C11907 VPWR.t912 VGND 0.02774f
C11908 VPWR.t491 VGND 0.02465f
C11909 VPWR.n560 VGND 0.0762f
C11910 VPWR.t1050 VGND 0.06535f
C11911 VPWR.t490 VGND 0.07675f
C11912 VPWR.t886 VGND 0.09955f
C11913 VPWR.t483 VGND 0.02774f
C11914 VPWR.t868 VGND 0.02465f
C11915 VPWR.n561 VGND 0.0762f
C11916 VPWR.n562 VGND 0.11584f
C11917 VPWR.n563 VGND 0.11584f
C11918 VPWR.t887 VGND 0.02774f
C11919 VPWR.t1186 VGND 0.02465f
C11920 VPWR.n564 VGND 0.0762f
C11921 VPWR.t1055 VGND 0.06535f
C11922 VPWR.t1185 VGND 0.07675f
C11923 VPWR.t723 VGND 0.09955f
C11924 VPWR.t885 VGND 0.02774f
C11925 VPWR.t732 VGND 0.02465f
C11926 VPWR.n565 VGND 0.0762f
C11927 VPWR.n566 VGND 0.11584f
C11928 VPWR.n567 VGND 0.11584f
C11929 VPWR.t724 VGND 0.02774f
C11930 VPWR.t1616 VGND 0.02465f
C11931 VPWR.n568 VGND 0.0762f
C11932 VPWR.t1642 VGND 0.06535f
C11933 VPWR.t1615 VGND 0.07675f
C11934 VPWR.t1828 VGND 0.09955f
C11935 VPWR.t1175 VGND 0.02774f
C11936 VPWR.t1837 VGND 0.02465f
C11937 VPWR.n569 VGND 0.0762f
C11938 VPWR.n570 VGND 0.11584f
C11939 VPWR.n571 VGND 0.11584f
C11940 VPWR.t1829 VGND 0.02774f
C11941 VPWR.t1086 VGND 0.02465f
C11942 VPWR.n572 VGND 0.0762f
C11943 VPWR.t1049 VGND 0.06535f
C11944 VPWR.t1085 VGND 0.07675f
C11945 VPWR.t564 VGND 0.09955f
C11946 VPWR.t1917 VGND 0.02774f
C11947 VPWR.t409 VGND 0.02465f
C11948 VPWR.n573 VGND 0.0762f
C11949 VPWR.n574 VGND 0.11584f
C11950 VPWR.n575 VGND 0.11584f
C11951 VPWR.t565 VGND 0.02774f
C11952 VPWR.t505 VGND 0.02465f
C11953 VPWR.n576 VGND 0.0762f
C11954 VPWR.t1645 VGND 0.06535f
C11955 VPWR.t504 VGND 0.07675f
C11956 VPWR.t781 VGND 0.02774f
C11957 VPWR.t216 VGND 0.02465f
C11958 VPWR.n577 VGND 0.0762f
C11959 VPWR.t605 VGND 0.02774f
C11960 VPWR.t324 VGND 0.02465f
C11961 VPWR.n578 VGND 0.0762f
C11962 VPWR.t1113 VGND 0.12083f
C11963 VPWR.t1428 VGND 0.06535f
C11964 VPWR.t1197 VGND 0.07675f
C11965 VPWR.t1114 VGND 0.02774f
C11966 VPWR.t1198 VGND 0.02465f
C11967 VPWR.n579 VGND 0.0762f
C11968 VPWR.n580 VGND 0.01496f
C11969 VPWR.n582 VGND 0.0901f
C11970 VPWR.t1018 VGND 0.09955f
C11971 VPWR.t1423 VGND 0.06535f
C11972 VPWR.t1597 VGND 0.07675f
C11973 VPWR.t1019 VGND 0.02774f
C11974 VPWR.t1598 VGND 0.02465f
C11975 VPWR.n583 VGND 0.0762f
C11976 VPWR.n584 VGND 0.01496f
C11977 VPWR.n586 VGND 0.0901f
C11978 VPWR.t471 VGND 0.09955f
C11979 VPWR.t698 VGND 0.06535f
C11980 VPWR.t1436 VGND 0.07675f
C11981 VPWR.t472 VGND 0.02774f
C11982 VPWR.t1437 VGND 0.02465f
C11983 VPWR.n587 VGND 0.0762f
C11984 VPWR.n588 VGND 0.01496f
C11985 VPWR.n590 VGND 0.0901f
C11986 VPWR.t1460 VGND 0.09955f
C11987 VPWR.t697 VGND 0.06535f
C11988 VPWR.t1276 VGND 0.07675f
C11989 VPWR.t1461 VGND 0.02774f
C11990 VPWR.t1277 VGND 0.02465f
C11991 VPWR.n591 VGND 0.0762f
C11992 VPWR.n592 VGND 0.01496f
C11993 VPWR.n594 VGND 0.0901f
C11994 VPWR.t396 VGND 0.09955f
C11995 VPWR.t1427 VGND 0.06535f
C11996 VPWR.t586 VGND 0.07675f
C11997 VPWR.t397 VGND 0.02774f
C11998 VPWR.t587 VGND 0.02465f
C11999 VPWR.n595 VGND 0.0762f
C12000 VPWR.n596 VGND 0.01496f
C12001 VPWR.n598 VGND 0.0901f
C12002 VPWR.t1545 VGND 0.09955f
C12003 VPWR.t1878 VGND 0.06535f
C12004 VPWR.t1138 VGND 0.07675f
C12005 VPWR.t1546 VGND 0.02774f
C12006 VPWR.t1139 VGND 0.02465f
C12007 VPWR.n599 VGND 0.0762f
C12008 VPWR.n600 VGND 0.01496f
C12009 VPWR.n602 VGND 0.0901f
C12010 VPWR.t1155 VGND 0.09955f
C12011 VPWR.t1877 VGND 0.06535f
C12012 VPWR.t816 VGND 0.07675f
C12013 VPWR.t1156 VGND 0.02774f
C12014 VPWR.t817 VGND 0.02465f
C12015 VPWR.n603 VGND 0.0762f
C12016 VPWR.n604 VGND 0.01496f
C12017 VPWR.n606 VGND 0.0901f
C12018 VPWR.t810 VGND 0.09955f
C12019 VPWR.t1426 VGND 0.06535f
C12020 VPWR.t892 VGND 0.07675f
C12021 VPWR.t811 VGND 0.02774f
C12022 VPWR.t893 VGND 0.02465f
C12023 VPWR.n607 VGND 0.0762f
C12024 VPWR.n608 VGND 0.01496f
C12025 VPWR.n610 VGND 0.0901f
C12026 VPWR.t932 VGND 0.09955f
C12027 VPWR.t1425 VGND 0.06535f
C12028 VPWR.t951 VGND 0.07675f
C12029 VPWR.t933 VGND 0.02774f
C12030 VPWR.t952 VGND 0.02465f
C12031 VPWR.n611 VGND 0.0762f
C12032 VPWR.n612 VGND 0.01496f
C12033 VPWR.n614 VGND 0.0901f
C12034 VPWR.t945 VGND 0.09955f
C12035 VPWR.t1422 VGND 0.06535f
C12036 VPWR.t1244 VGND 0.07675f
C12037 VPWR.t946 VGND 0.02774f
C12038 VPWR.t1245 VGND 0.02465f
C12039 VPWR.n615 VGND 0.0762f
C12040 VPWR.n616 VGND 0.01496f
C12041 VPWR.n618 VGND 0.0901f
C12042 VPWR.t1234 VGND 0.09955f
C12043 VPWR.t696 VGND 0.06535f
C12044 VPWR.t1341 VGND 0.07675f
C12045 VPWR.t1235 VGND 0.02774f
C12046 VPWR.t1342 VGND 0.02465f
C12047 VPWR.n619 VGND 0.0762f
C12048 VPWR.n620 VGND 0.01496f
C12049 VPWR.n622 VGND 0.0901f
C12050 VPWR.t1320 VGND 0.09955f
C12051 VPWR.t695 VGND 0.06535f
C12052 VPWR.t1838 VGND 0.07675f
C12053 VPWR.t1321 VGND 0.02774f
C12054 VPWR.t1839 VGND 0.02465f
C12055 VPWR.n623 VGND 0.0762f
C12056 VPWR.n624 VGND 0.01496f
C12057 VPWR.n626 VGND 0.0901f
C12058 VPWR.t1248 VGND 0.09955f
C12059 VPWR.t1876 VGND 0.06535f
C12060 VPWR.t1922 VGND 0.07675f
C12061 VPWR.t1249 VGND 0.02774f
C12062 VPWR.t1923 VGND 0.02465f
C12063 VPWR.n627 VGND 0.0762f
C12064 VPWR.n628 VGND 0.01496f
C12065 VPWR.n630 VGND 0.0901f
C12066 VPWR.t1715 VGND 0.09955f
C12067 VPWR.t1875 VGND 0.06535f
C12068 VPWR.t759 VGND 0.07675f
C12069 VPWR.t1716 VGND 0.02774f
C12070 VPWR.t760 VGND 0.02465f
C12071 VPWR.n631 VGND 0.0762f
C12072 VPWR.n632 VGND 0.01496f
C12073 VPWR.n634 VGND 0.0901f
C12074 VPWR.t735 VGND 0.09955f
C12075 VPWR.t1874 VGND 0.06535f
C12076 VPWR.t782 VGND 0.07675f
C12077 VPWR.t736 VGND 0.02774f
C12078 VPWR.t783 VGND 0.02465f
C12079 VPWR.n635 VGND 0.0762f
C12080 VPWR.n636 VGND 0.01496f
C12081 VPWR.n638 VGND 0.0901f
C12082 VPWR.t604 VGND 0.09955f
C12083 VPWR.t1424 VGND 0.06535f
C12084 VPWR.t323 VGND 0.11101f
C12085 VPWR.n639 VGND 0.06343f
C12086 VPWR.n640 VGND 0.01496f
C12087 VPWR.n641 VGND 0.11584f
C12088 VPWR.n642 VGND 0.84572f
C12089 VPWR.n643 VGND 0.11584f
C12090 VPWR.t523 VGND 0.02774f
C12091 VPWR.t50 VGND 0.02465f
C12092 VPWR.n644 VGND 0.0762f
C12093 VPWR.t606 VGND 0.07675f
C12094 VPWR.t1497 VGND 0.02774f
C12095 VPWR.t607 VGND 0.02465f
C12096 VPWR.n645 VGND 0.0762f
C12097 VPWR.n646 VGND 0.11584f
C12098 VPWR.n647 VGND 0.11584f
C12099 VPWR.t1297 VGND 0.02774f
C12100 VPWR.t1503 VGND 0.02465f
C12101 VPWR.n648 VGND 0.0762f
C12102 VPWR.t1719 VGND 0.07675f
C12103 VPWR.t1283 VGND 0.02774f
C12104 VPWR.t1720 VGND 0.02465f
C12105 VPWR.n649 VGND 0.0762f
C12106 VPWR.n650 VGND 0.11584f
C12107 VPWR.n651 VGND 0.11584f
C12108 VPWR.t1665 VGND 0.02774f
C12109 VPWR.t1353 VGND 0.02465f
C12110 VPWR.n652 VGND 0.0762f
C12111 VPWR.t922 VGND 0.07675f
C12112 VPWR.t507 VGND 0.02774f
C12113 VPWR.t923 VGND 0.02465f
C12114 VPWR.n653 VGND 0.0762f
C12115 VPWR.n654 VGND 0.11584f
C12116 VPWR.n655 VGND 0.11584f
C12117 VPWR.t545 VGND 0.02774f
C12118 VPWR.t513 VGND 0.02465f
C12119 VPWR.n656 VGND 0.0762f
C12120 VPWR.t550 VGND 0.07675f
C12121 VPWR.t872 VGND 0.02774f
C12122 VPWR.t551 VGND 0.02465f
C12123 VPWR.n657 VGND 0.0762f
C12124 VPWR.n658 VGND 0.11584f
C12125 VPWR.n659 VGND 0.11584f
C12126 VPWR.t1590 VGND 0.02774f
C12127 VPWR.t937 VGND 0.02465f
C12128 VPWR.n660 VGND 0.0762f
C12129 VPWR.t794 VGND 0.07675f
C12130 VPWR.t621 VGND 0.02774f
C12131 VPWR.t795 VGND 0.02465f
C12132 VPWR.n661 VGND 0.0762f
C12133 VPWR.n662 VGND 0.11584f
C12134 VPWR.n663 VGND 0.11584f
C12135 VPWR.t1330 VGND 0.02774f
C12136 VPWR.t627 VGND 0.02465f
C12137 VPWR.n664 VGND 0.0762f
C12138 VPWR.t1635 VGND 0.07675f
C12139 VPWR.t999 VGND 0.02774f
C12140 VPWR.t1636 VGND 0.02465f
C12141 VPWR.n665 VGND 0.0762f
C12142 VPWR.n666 VGND 0.11584f
C12143 VPWR.n667 VGND 0.11584f
C12144 VPWR.t1483 VGND 0.02774f
C12145 VPWR.t399 VGND 0.02465f
C12146 VPWR.n668 VGND 0.0762f
C12147 VPWR.t1456 VGND 0.07675f
C12148 VPWR.t1552 VGND 0.02774f
C12149 VPWR.t1457 VGND 0.02465f
C12150 VPWR.n669 VGND 0.0762f
C12151 VPWR.n670 VGND 0.11584f
C12152 VPWR.n671 VGND 0.11584f
C12153 VPWR.t825 VGND 0.02774f
C12154 VPWR.t1558 VGND 0.02465f
C12155 VPWR.n672 VGND 0.0762f
C12156 VPWR.t1125 VGND 0.12083f
C12157 VPWR.t1061 VGND 0.06535f
C12158 VPWR.t969 VGND 0.07675f
C12159 VPWR.t1126 VGND 0.02774f
C12160 VPWR.t970 VGND 0.02465f
C12161 VPWR.n673 VGND 0.0762f
C12162 VPWR.t1133 VGND 0.02774f
C12163 VPWR.t1011 VGND 0.02465f
C12164 VPWR.n674 VGND 0.0762f
C12165 VPWR.t1132 VGND 0.12083f
C12166 VPWR.t633 VGND 0.06535f
C12167 VPWR.t1010 VGND 0.07675f
C12168 VPWR.t1845 VGND 0.02774f
C12169 VPWR.t157 VGND 0.02465f
C12170 VPWR.n675 VGND 0.0762f
C12171 VPWR.n676 VGND 0.01496f
C12172 VPWR.n677 VGND 0.06343f
C12173 VPWR.t156 VGND 0.11101f
C12174 VPWR.t1822 VGND 0.06535f
C12175 VPWR.t1844 VGND 0.09955f
C12176 VPWR.t411 VGND 0.02774f
C12177 VPWR.t527 VGND 0.02465f
C12178 VPWR.n678 VGND 0.0762f
C12179 VPWR.n679 VGND 0.01496f
C12180 VPWR.n681 VGND 0.0901f
C12181 VPWR.t526 VGND 0.07675f
C12182 VPWR.t1351 VGND 0.06535f
C12183 VPWR.t410 VGND 0.09955f
C12184 VPWR.t1076 VGND 0.02774f
C12185 VPWR.t417 VGND 0.02465f
C12186 VPWR.n682 VGND 0.0762f
C12187 VPWR.n683 VGND 0.01496f
C12188 VPWR.n685 VGND 0.0901f
C12189 VPWR.t416 VGND 0.07675f
C12190 VPWR.t1064 VGND 0.06535f
C12191 VPWR.t1075 VGND 0.09955f
C12192 VPWR.t1572 VGND 0.02774f
C12193 VPWR.t1303 VGND 0.02465f
C12194 VPWR.n686 VGND 0.0762f
C12195 VPWR.n687 VGND 0.01496f
C12196 VPWR.n689 VGND 0.0901f
C12197 VPWR.t1302 VGND 0.07675f
C12198 VPWR.t1065 VGND 0.06535f
C12199 VPWR.t1571 VGND 0.09955f
C12200 VPWR.t1620 VGND 0.02774f
C12201 VPWR.t1566 VGND 0.02465f
C12202 VPWR.n690 VGND 0.0762f
C12203 VPWR.n691 VGND 0.01496f
C12204 VPWR.n693 VGND 0.0901f
C12205 VPWR.t1565 VGND 0.07675f
C12206 VPWR.t634 VGND 0.06535f
C12207 VPWR.t1619 VGND 0.09955f
C12208 VPWR.t744 VGND 0.02774f
C12209 VPWR.t1608 VGND 0.02465f
C12210 VPWR.n694 VGND 0.0762f
C12211 VPWR.n695 VGND 0.01496f
C12212 VPWR.n697 VGND 0.0901f
C12213 VPWR.t1607 VGND 0.07675f
C12214 VPWR.t1348 VGND 0.06535f
C12215 VPWR.t743 VGND 0.09955f
C12216 VPWR.t1683 VGND 0.02774f
C12217 VPWR.t750 VGND 0.02465f
C12218 VPWR.n698 VGND 0.0762f
C12219 VPWR.n699 VGND 0.01496f
C12220 VPWR.n701 VGND 0.0901f
C12221 VPWR.t749 VGND 0.07675f
C12222 VPWR.t1068 VGND 0.06535f
C12223 VPWR.t1682 VGND 0.09955f
C12224 VPWR.t899 VGND 0.02774f
C12225 VPWR.t1687 VGND 0.02465f
C12226 VPWR.n702 VGND 0.0762f
C12227 VPWR.n703 VGND 0.01496f
C12228 VPWR.n705 VGND 0.0901f
C12229 VPWR.t1686 VGND 0.07675f
C12230 VPWR.t1823 VGND 0.06535f
C12231 VPWR.t898 VGND 0.09955f
C12232 VPWR.t1578 VGND 0.02774f
C12233 VPWR.t661 VGND 0.02465f
C12234 VPWR.n706 VGND 0.0762f
C12235 VPWR.n707 VGND 0.01496f
C12236 VPWR.n709 VGND 0.0901f
C12237 VPWR.t660 VGND 0.07675f
C12238 VPWR.t1144 VGND 0.06535f
C12239 VPWR.t1577 VGND 0.09955f
C12240 VPWR.t958 VGND 0.02774f
C12241 VPWR.t1582 VGND 0.02465f
C12242 VPWR.n710 VGND 0.0762f
C12243 VPWR.n711 VGND 0.01496f
C12244 VPWR.n713 VGND 0.0901f
C12245 VPWR.t1581 VGND 0.07675f
C12246 VPWR.t1066 VGND 0.06535f
C12247 VPWR.t957 VGND 0.09955f
C12248 VPWR.t1594 VGND 0.02774f
C12249 VPWR.t962 VGND 0.02465f
C12250 VPWR.n714 VGND 0.0762f
C12251 VPWR.n715 VGND 0.01496f
C12252 VPWR.n717 VGND 0.0901f
C12253 VPWR.t961 VGND 0.07675f
C12254 VPWR.t1067 VGND 0.06535f
C12255 VPWR.t1593 VGND 0.09955f
C12256 VPWR.t1507 VGND 0.02774f
C12257 VPWR.t1622 VGND 0.02465f
C12258 VPWR.n718 VGND 0.0762f
C12259 VPWR.n719 VGND 0.01496f
C12260 VPWR.n721 VGND 0.0901f
C12261 VPWR.t1621 VGND 0.07675f
C12262 VPWR.t632 VGND 0.06535f
C12263 VPWR.t1506 VGND 0.09955f
C12264 VPWR.t1495 VGND 0.02774f
C12265 VPWR.t1393 VGND 0.02465f
C12266 VPWR.n722 VGND 0.0762f
C12267 VPWR.n723 VGND 0.01496f
C12268 VPWR.n725 VGND 0.0901f
C12269 VPWR.t1392 VGND 0.07675f
C12270 VPWR.t1349 VGND 0.06535f
C12271 VPWR.t1494 VGND 0.09955f
C12272 VPWR.t688 VGND 0.02774f
C12273 VPWR.t1475 VGND 0.02465f
C12274 VPWR.n726 VGND 0.0762f
C12275 VPWR.n727 VGND 0.01496f
C12276 VPWR.n729 VGND 0.0901f
C12277 VPWR.t1474 VGND 0.07675f
C12278 VPWR.t1350 VGND 0.06535f
C12279 VPWR.t687 VGND 0.09955f
C12280 VPWR.t1190 VGND 0.02774f
C12281 VPWR.t692 VGND 0.02465f
C12282 VPWR.n730 VGND 0.0762f
C12283 VPWR.n731 VGND 0.01496f
C12284 VPWR.n733 VGND 0.0901f
C12285 VPWR.t691 VGND 0.07675f
C12286 VPWR.t1821 VGND 0.06535f
C12287 VPWR.t1189 VGND 0.09955f
C12288 VPWR.n734 VGND 0.0901f
C12289 VPWR.n736 VGND 0.01496f
C12290 VPWR.n737 VGND 0.11584f
C12291 VPWR.n738 VGND 0.84042f
C12292 VPWR.n739 VGND 0.11584f
C12293 VPWR.t1129 VGND 0.02774f
C12294 VPWR.t823 VGND 0.02465f
C12295 VPWR.n740 VGND 0.0762f
C12296 VPWR.t1128 VGND 0.12083f
C12297 VPWR.t1629 VGND 0.06535f
C12298 VPWR.t822 VGND 0.07675f
C12299 VPWR.t1028 VGND 0.09955f
C12300 VPWR.t1013 VGND 0.02774f
C12301 VPWR.t1031 VGND 0.02465f
C12302 VPWR.n741 VGND 0.0762f
C12303 VPWR.n742 VGND 0.11584f
C12304 VPWR.n743 VGND 0.11584f
C12305 VPWR.t1029 VGND 0.02774f
C12306 VPWR.t1465 VGND 0.02465f
C12307 VPWR.n744 VGND 0.0762f
C12308 VPWR.t1633 VGND 0.06535f
C12309 VPWR.t1464 VGND 0.07675f
C12310 VPWR.t1510 VGND 0.09955f
C12311 VPWR.t1489 VGND 0.02774f
C12312 VPWR.t389 VGND 0.02465f
C12313 VPWR.n745 VGND 0.0762f
C12314 VPWR.n746 VGND 0.11584f
C12315 VPWR.n747 VGND 0.11584f
C12316 VPWR.t1511 VGND 0.02774f
C12317 VPWR.t1628 VGND 0.02465f
C12318 VPWR.n748 VGND 0.0762f
C12319 VPWR.t468 VGND 0.06535f
C12320 VPWR.t1627 VGND 0.07675f
C12321 VPWR.t654 VGND 0.09955f
C12322 VPWR.t1626 VGND 0.02774f
C12323 VPWR.t657 VGND 0.02465f
C12324 VPWR.n749 VGND 0.0762f
C12325 VPWR.n750 VGND 0.11584f
C12326 VPWR.n751 VGND 0.11584f
C12327 VPWR.t655 VGND 0.02774f
C12328 VPWR.t1588 VGND 0.02465f
C12329 VPWR.n752 VGND 0.0762f
C12330 VPWR.t1601 VGND 0.06535f
C12331 VPWR.t1587 VGND 0.07675f
C12332 VPWR.t664 VGND 0.09955f
C12333 VPWR.t1586 VGND 0.02774f
C12334 VPWR.t834 VGND 0.02465f
C12335 VPWR.n753 VGND 0.0762f
C12336 VPWR.n754 VGND 0.11584f
C12337 VPWR.n755 VGND 0.11584f
C12338 VPWR.t665 VGND 0.02774f
C12339 VPWR.t1037 VGND 0.02465f
C12340 VPWR.n756 VGND 0.0762f
C12341 VPWR.t466 VGND 0.06535f
C12342 VPWR.t1036 VGND 0.07675f
C12343 VPWR.t751 VGND 0.09955f
C12344 VPWR.t1035 VGND 0.02774f
C12345 VPWR.t756 VGND 0.02465f
C12346 VPWR.n757 VGND 0.0762f
C12347 VPWR.n758 VGND 0.11584f
C12348 VPWR.n759 VGND 0.11584f
C12349 VPWR.t752 VGND 0.02774f
C12350 VPWR.t1663 VGND 0.02465f
C12351 VPWR.n760 VGND 0.0762f
C12352 VPWR.t1631 VGND 0.06535f
C12353 VPWR.t1662 VGND 0.07675f
C12354 VPWR.t1567 VGND 0.09955f
C12355 VPWR.t879 VGND 0.02774f
C12356 VPWR.t1533 VGND 0.02465f
C12357 VPWR.n761 VGND 0.0762f
C12358 VPWR.n762 VGND 0.11584f
C12359 VPWR.n763 VGND 0.11584f
C12360 VPWR.t1568 VGND 0.02774f
C12361 VPWR.t1309 VGND 0.02465f
C12362 VPWR.n764 VGND 0.0762f
C12363 VPWR.t1600 VGND 0.06535f
C12364 VPWR.t1308 VGND 0.07675f
C12365 VPWR.t418 VGND 0.09955f
C12366 VPWR.t1080 VGND 0.02774f
C12367 VPWR.t1882 VGND 0.02465f
C12368 VPWR.n765 VGND 0.0762f
C12369 VPWR.n766 VGND 0.11584f
C12370 VPWR.n767 VGND 0.11584f
C12371 VPWR.t419 VGND 0.02774f
C12372 VPWR.t533 VGND 0.02465f
C12373 VPWR.n768 VGND 0.0762f
C12374 VPWR.t1634 VGND 0.06535f
C12375 VPWR.t532 VGND 0.07675f
C12376 VPWR.t1849 VGND 0.02774f
C12377 VPWR.t117 VGND 0.02465f
C12378 VPWR.n769 VGND 0.0762f
C12379 VPWR.t777 VGND 0.02774f
C12380 VPWR.t222 VGND 0.02465f
C12381 VPWR.n770 VGND 0.0762f
C12382 VPWR.t1107 VGND 0.12083f
C12383 VPWR.t707 VGND 0.06535f
C12384 VPWR.t858 VGND 0.07675f
C12385 VPWR.t1108 VGND 0.02774f
C12386 VPWR.t859 VGND 0.02465f
C12387 VPWR.n771 VGND 0.0762f
C12388 VPWR.n772 VGND 0.01496f
C12389 VPWR.n774 VGND 0.0901f
C12390 VPWR.t433 VGND 0.09955f
C12391 VPWR.t702 VGND 0.06535f
C12392 VPWR.t1898 VGND 0.07675f
C12393 VPWR.t434 VGND 0.02774f
C12394 VPWR.t1899 VGND 0.02465f
C12395 VPWR.n775 VGND 0.0762f
C12396 VPWR.n776 VGND 0.01496f
C12397 VPWR.n778 VGND 0.0901f
C12398 VPWR.t1707 VGND 0.09955f
C12399 VPWR.t1004 VGND 0.06535f
C12400 VPWR.t1468 VGND 0.07675f
C12401 VPWR.t1708 VGND 0.02774f
C12402 VPWR.t1469 VGND 0.02465f
C12403 VPWR.n779 VGND 0.0762f
C12404 VPWR.n780 VGND 0.01496f
C12405 VPWR.n782 VGND 0.0901f
C12406 VPWR.t1448 VGND 0.09955f
C12407 VPWR.t1003 VGND 0.06535f
C12408 VPWR.t992 VGND 0.07675f
C12409 VPWR.t1449 VGND 0.02774f
C12410 VPWR.t993 VGND 0.02465f
C12411 VPWR.n783 VGND 0.0762f
C12412 VPWR.n784 VGND 0.01496f
C12413 VPWR.n786 VGND 0.0901f
C12414 VPWR.t1270 VGND 0.09955f
C12415 VPWR.t706 VGND 0.06535f
C12416 VPWR.t1699 VGND 0.07675f
C12417 VPWR.t1271 VGND 0.02774f
C12418 VPWR.t1700 VGND 0.02465f
C12419 VPWR.n787 VGND 0.0762f
C12420 VPWR.n788 VGND 0.01496f
C12421 VPWR.n790 VGND 0.0901f
C12422 VPWR.t1693 VGND 0.09955f
C12423 VPWR.t1009 VGND 0.06535f
C12424 VPWR.t915 VGND 0.07675f
C12425 VPWR.t1694 VGND 0.02774f
C12426 VPWR.t916 VGND 0.02465f
C12427 VPWR.n791 VGND 0.0762f
C12428 VPWR.n792 VGND 0.01496f
C12429 VPWR.n794 VGND 0.0901f
C12430 VPWR.t909 VGND 0.09955f
C12431 VPWR.t1008 VGND 0.06535f
C12432 VPWR.t486 VGND 0.07675f
C12433 VPWR.t910 VGND 0.02774f
C12434 VPWR.t487 VGND 0.02465f
C12435 VPWR.n795 VGND 0.0762f
C12436 VPWR.n796 VGND 0.01496f
C12437 VPWR.n798 VGND 0.0901f
C12438 VPWR.t480 VGND 0.09955f
C12439 VPWR.t705 VGND 0.06535f
C12440 VPWR.t668 VGND 0.07675f
C12441 VPWR.t481 VGND 0.02774f
C12442 VPWR.t669 VGND 0.02465f
C12443 VPWR.n799 VGND 0.0762f
C12444 VPWR.n800 VGND 0.01496f
C12445 VPWR.n802 VGND 0.0901f
C12446 VPWR.t648 VGND 0.09955f
C12447 VPWR.t704 VGND 0.06535f
C12448 VPWR.t1181 VGND 0.07675f
C12449 VPWR.t649 VGND 0.02774f
C12450 VPWR.t1182 VGND 0.02465f
C12451 VPWR.n803 VGND 0.0762f
C12452 VPWR.n804 VGND 0.01496f
C12453 VPWR.n806 VGND 0.0901f
C12454 VPWR.t882 VGND 0.09955f
C12455 VPWR.t701 VGND 0.06535f
C12456 VPWR.t729 VGND 0.07675f
C12457 VPWR.t883 VGND 0.02774f
C12458 VPWR.t730 VGND 0.02465f
C12459 VPWR.n807 VGND 0.0762f
C12460 VPWR.n808 VGND 0.01496f
C12461 VPWR.n810 VGND 0.0901f
C12462 VPWR.t721 VGND 0.09955f
C12463 VPWR.t1002 VGND 0.06535f
C12464 VPWR.t1611 VGND 0.07675f
C12465 VPWR.t722 VGND 0.02774f
C12466 VPWR.t1612 VGND 0.02465f
C12467 VPWR.n811 VGND 0.0762f
C12468 VPWR.n812 VGND 0.01496f
C12469 VPWR.n814 VGND 0.0901f
C12470 VPWR.t1172 VGND 0.09955f
C12471 VPWR.t1001 VGND 0.06535f
C12472 VPWR.t1834 VGND 0.07675f
C12473 VPWR.t1173 VGND 0.02774f
C12474 VPWR.t1835 VGND 0.02465f
C12475 VPWR.n815 VGND 0.0762f
C12476 VPWR.n816 VGND 0.01496f
C12477 VPWR.n818 VGND 0.0901f
C12478 VPWR.t536 VGND 0.09955f
C12479 VPWR.t1007 VGND 0.06535f
C12480 VPWR.t1083 VGND 0.07675f
C12481 VPWR.t537 VGND 0.02774f
C12482 VPWR.t1084 VGND 0.02465f
C12483 VPWR.n819 VGND 0.0762f
C12484 VPWR.n820 VGND 0.01496f
C12485 VPWR.n822 VGND 0.0901f
C12486 VPWR.t1912 VGND 0.09955f
C12487 VPWR.t1006 VGND 0.06535f
C12488 VPWR.t406 VGND 0.07675f
C12489 VPWR.t1913 VGND 0.02774f
C12490 VPWR.t407 VGND 0.02465f
C12491 VPWR.n823 VGND 0.0762f
C12492 VPWR.n824 VGND 0.01496f
C12493 VPWR.n826 VGND 0.0901f
C12494 VPWR.t562 VGND 0.09955f
C12495 VPWR.t1005 VGND 0.06535f
C12496 VPWR.t1852 VGND 0.07675f
C12497 VPWR.t563 VGND 0.02774f
C12498 VPWR.t1853 VGND 0.02465f
C12499 VPWR.n827 VGND 0.0762f
C12500 VPWR.n828 VGND 0.01496f
C12501 VPWR.n830 VGND 0.0901f
C12502 VPWR.t776 VGND 0.09955f
C12503 VPWR.t703 VGND 0.06535f
C12504 VPWR.t221 VGND 0.11101f
C12505 VPWR.n831 VGND 0.06343f
C12506 VPWR.n832 VGND 0.01496f
C12507 VPWR.n833 VGND 0.11584f
C12508 VPWR.n834 VGND 0.84572f
C12509 VPWR.n835 VGND 0.11584f
C12510 VPWR.t525 VGND 0.02774f
C12511 VPWR.t45 VGND 0.02465f
C12512 VPWR.n836 VGND 0.0762f
C12513 VPWR.t610 VGND 0.07675f
C12514 VPWR.t1499 VGND 0.02774f
C12515 VPWR.t611 VGND 0.02465f
C12516 VPWR.n837 VGND 0.0762f
C12517 VPWR.n838 VGND 0.11584f
C12518 VPWR.n839 VGND 0.11584f
C12519 VPWR.t1299 VGND 0.02774f
C12520 VPWR.t1371 VGND 0.02465f
C12521 VPWR.n840 VGND 0.0762f
C12522 VPWR.t1721 VGND 0.07675f
C12523 VPWR.t1285 VGND 0.02774f
C12524 VPWR.t1722 VGND 0.02465f
C12525 VPWR.n841 VGND 0.0762f
C12526 VPWR.n842 VGND 0.11584f
C12527 VPWR.n843 VGND 0.11584f
C12528 VPWR.t1667 VGND 0.02774f
C12529 VPWR.t1355 VGND 0.02465f
C12530 VPWR.n844 VGND 0.0762f
C12531 VPWR.t924 VGND 0.07675f
C12532 VPWR.t509 VGND 0.02774f
C12533 VPWR.t925 VGND 0.02465f
C12534 VPWR.n845 VGND 0.0762f
C12535 VPWR.n846 VGND 0.11584f
C12536 VPWR.n847 VGND 0.11584f
C12537 VPWR.t547 VGND 0.02774f
C12538 VPWR.t515 VGND 0.02465f
C12539 VPWR.n848 VGND 0.0762f
C12540 VPWR.t552 VGND 0.07675f
C12541 VPWR.t874 VGND 0.02774f
C12542 VPWR.t553 VGND 0.02465f
C12543 VPWR.n849 VGND 0.0762f
C12544 VPWR.n850 VGND 0.11584f
C12545 VPWR.n851 VGND 0.11584f
C12546 VPWR.t791 VGND 0.02774f
C12547 VPWR.t939 VGND 0.02465f
C12548 VPWR.n852 VGND 0.0762f
C12549 VPWR.t796 VGND 0.07675f
C12550 VPWR.t623 VGND 0.02774f
C12551 VPWR.t797 VGND 0.02465f
C12552 VPWR.n853 VGND 0.0762f
C12553 VPWR.n854 VGND 0.11584f
C12554 VPWR.n855 VGND 0.11584f
C12555 VPWR.t1332 VGND 0.02774f
C12556 VPWR.t629 VGND 0.02465f
C12557 VPWR.n856 VGND 0.0762f
C12558 VPWR.t1637 VGND 0.07675f
C12559 VPWR.t1391 VGND 0.02774f
C12560 VPWR.t1638 VGND 0.02465f
C12561 VPWR.n857 VGND 0.0762f
C12562 VPWR.n858 VGND 0.11584f
C12563 VPWR.n859 VGND 0.11584f
C12564 VPWR.t1481 VGND 0.02774f
C12565 VPWR.t1517 VGND 0.02465f
C12566 VPWR.n860 VGND 0.0762f
C12567 VPWR.t1454 VGND 0.07675f
C12568 VPWR.t1554 VGND 0.02774f
C12569 VPWR.t1455 VGND 0.02465f
C12570 VPWR.n861 VGND 0.0762f
C12571 VPWR.n862 VGND 0.11584f
C12572 VPWR.n863 VGND 0.11584f
C12573 VPWR.t827 VGND 0.02774f
C12574 VPWR.t1560 VGND 0.02465f
C12575 VPWR.n864 VGND 0.0762f
C12576 VPWR.t1123 VGND 0.12083f
C12577 VPWR.t713 VGND 0.06535f
C12578 VPWR.t971 VGND 0.07675f
C12579 VPWR.t1124 VGND 0.02774f
C12580 VPWR.t972 VGND 0.02465f
C12581 VPWR.n865 VGND 0.0762f
C12582 VPWR.t1110 VGND 0.02774f
C12583 VPWR.t857 VGND 0.02465f
C12584 VPWR.n866 VGND 0.0762f
C12585 VPWR.t1109 VGND 0.12083f
C12586 VPWR.t968 VGND 0.06535f
C12587 VPWR.t856 VGND 0.07675f
C12588 VPWR.t775 VGND 0.02774f
C12589 VPWR.t229 VGND 0.02465f
C12590 VPWR.n867 VGND 0.0762f
C12591 VPWR.n868 VGND 0.01496f
C12592 VPWR.n869 VGND 0.06343f
C12593 VPWR.t228 VGND 0.11101f
C12594 VPWR.t964 VGND 0.06535f
C12595 VPWR.t774 VGND 0.09955f
C12596 VPWR.t561 VGND 0.02774f
C12597 VPWR.t1851 VGND 0.02465f
C12598 VPWR.n870 VGND 0.0762f
C12599 VPWR.n871 VGND 0.01496f
C12600 VPWR.n873 VGND 0.0901f
C12601 VPWR.t1850 VGND 0.07675f
C12602 VPWR.t846 VGND 0.06535f
C12603 VPWR.t560 VGND 0.09955f
C12604 VPWR.t1909 VGND 0.02774f
C12605 VPWR.t405 VGND 0.02465f
C12606 VPWR.n874 VGND 0.0762f
C12607 VPWR.n875 VGND 0.01496f
C12608 VPWR.n877 VGND 0.0901f
C12609 VPWR.t404 VGND 0.07675f
C12610 VPWR.t847 VGND 0.06535f
C12611 VPWR.t1908 VGND 0.09955f
C12612 VPWR.t535 VGND 0.02774f
C12613 VPWR.t1082 VGND 0.02465f
C12614 VPWR.n878 VGND 0.0762f
C12615 VPWR.n879 VGND 0.01496f
C12616 VPWR.n881 VGND 0.0901f
C12617 VPWR.t1081 VGND 0.07675f
C12618 VPWR.t848 VGND 0.06535f
C12619 VPWR.t534 VGND 0.09955f
C12620 VPWR.t1171 VGND 0.02774f
C12621 VPWR.t1833 VGND 0.02465f
C12622 VPWR.n882 VGND 0.0762f
C12623 VPWR.n883 VGND 0.01496f
C12624 VPWR.n885 VGND 0.0901f
C12625 VPWR.t1832 VGND 0.07675f
C12626 VPWR.t1859 VGND 0.06535f
C12627 VPWR.t1170 VGND 0.09955f
C12628 VPWR.t720 VGND 0.02774f
C12629 VPWR.t1177 VGND 0.02465f
C12630 VPWR.n886 VGND 0.0762f
C12631 VPWR.n887 VGND 0.01496f
C12632 VPWR.n889 VGND 0.0901f
C12633 VPWR.t1176 VGND 0.07675f
C12634 VPWR.t1860 VGND 0.06535f
C12635 VPWR.t719 VGND 0.09955f
C12636 VPWR.t881 VGND 0.02774f
C12637 VPWR.t728 VGND 0.02465f
C12638 VPWR.n890 VGND 0.0762f
C12639 VPWR.n891 VGND 0.01496f
C12640 VPWR.n893 VGND 0.0901f
C12641 VPWR.t727 VGND 0.07675f
C12642 VPWR.t851 VGND 0.06535f
C12643 VPWR.t880 VGND 0.09955f
C12644 VPWR.t645 VGND 0.02774f
C12645 VPWR.t1180 VGND 0.02465f
C12646 VPWR.n894 VGND 0.0762f
C12647 VPWR.n895 VGND 0.01496f
C12648 VPWR.n897 VGND 0.0901f
C12649 VPWR.t1179 VGND 0.07675f
C12650 VPWR.t965 VGND 0.06535f
C12651 VPWR.t644 VGND 0.09955f
C12652 VPWR.t479 VGND 0.02774f
C12653 VPWR.t667 VGND 0.02465f
C12654 VPWR.n898 VGND 0.0762f
C12655 VPWR.n899 VGND 0.01496f
C12656 VPWR.n901 VGND 0.0901f
C12657 VPWR.t666 VGND 0.07675f
C12658 VPWR.t966 VGND 0.06535f
C12659 VPWR.t478 VGND 0.09955f
C12660 VPWR.t908 VGND 0.02774f
C12661 VPWR.t485 VGND 0.02465f
C12662 VPWR.n902 VGND 0.0762f
C12663 VPWR.n903 VGND 0.01496f
C12664 VPWR.n905 VGND 0.0901f
C12665 VPWR.t484 VGND 0.07675f
C12666 VPWR.t849 VGND 0.06535f
C12667 VPWR.t907 VGND 0.09955f
C12668 VPWR.t1673 VGND 0.02774f
C12669 VPWR.t914 VGND 0.02465f
C12670 VPWR.n906 VGND 0.0762f
C12671 VPWR.n907 VGND 0.01496f
C12672 VPWR.n909 VGND 0.0901f
C12673 VPWR.t913 VGND 0.07675f
C12674 VPWR.t850 VGND 0.06535f
C12675 VPWR.t1672 VGND 0.09955f
C12676 VPWR.t1269 VGND 0.02774f
C12677 VPWR.t1698 VGND 0.02465f
C12678 VPWR.n910 VGND 0.0762f
C12679 VPWR.n911 VGND 0.01496f
C12680 VPWR.n913 VGND 0.0901f
C12681 VPWR.t1697 VGND 0.07675f
C12682 VPWR.t967 VGND 0.06535f
C12683 VPWR.t1268 VGND 0.09955f
C12684 VPWR.t1451 VGND 0.02774f
C12685 VPWR.t1513 VGND 0.02465f
C12686 VPWR.n914 VGND 0.0762f
C12687 VPWR.n915 VGND 0.01496f
C12688 VPWR.n917 VGND 0.0901f
C12689 VPWR.t1512 VGND 0.07675f
C12690 VPWR.t1861 VGND 0.06535f
C12691 VPWR.t1450 VGND 0.09955f
C12692 VPWR.t1706 VGND 0.02774f
C12693 VPWR.t1487 VGND 0.02465f
C12694 VPWR.n918 VGND 0.0762f
C12695 VPWR.n919 VGND 0.01496f
C12696 VPWR.n921 VGND 0.0901f
C12697 VPWR.t1486 VGND 0.07675f
C12698 VPWR.t845 VGND 0.06535f
C12699 VPWR.t1705 VGND 0.09955f
C12700 VPWR.t432 VGND 0.02774f
C12701 VPWR.t1897 VGND 0.02465f
C12702 VPWR.n922 VGND 0.0762f
C12703 VPWR.n923 VGND 0.01496f
C12704 VPWR.n925 VGND 0.0901f
C12705 VPWR.t1896 VGND 0.07675f
C12706 VPWR.t963 VGND 0.06535f
C12707 VPWR.t431 VGND 0.09955f
C12708 VPWR.n926 VGND 0.0901f
C12709 VPWR.n928 VGND 0.01496f
C12710 VPWR.n929 VGND 0.11584f
C12711 VPWR.n930 VGND 0.84042f
C12712 VPWR.n931 VGND 0.11584f
C12713 VPWR.t1116 VGND 0.02774f
C12714 VPWR.t1196 VGND 0.02465f
C12715 VPWR.n932 VGND 0.0762f
C12716 VPWR.t1115 VGND 0.12083f
C12717 VPWR.t539 VGND 0.06535f
C12718 VPWR.t1195 VGND 0.07675f
C12719 VPWR.t1680 VGND 0.09955f
C12720 VPWR.t1017 VGND 0.02774f
C12721 VPWR.t476 VGND 0.02465f
C12722 VPWR.n933 VGND 0.0762f
C12723 VPWR.n934 VGND 0.11584f
C12724 VPWR.n935 VGND 0.11584f
C12725 VPWR.t1681 VGND 0.02774f
C12726 VPWR.t1439 VGND 0.02465f
C12727 VPWR.n936 VGND 0.0762f
C12728 VPWR.t543 VGND 0.06535f
C12729 VPWR.t1438 VGND 0.07675f
C12730 VPWR.t394 VGND 0.09955f
C12731 VPWR.t1463 VGND 0.02774f
C12732 VPWR.t1273 VGND 0.02465f
C12733 VPWR.n937 VGND 0.0762f
C12734 VPWR.n938 VGND 0.11584f
C12735 VPWR.n939 VGND 0.11584f
C12736 VPWR.t395 VGND 0.02774f
C12737 VPWR.t1550 VGND 0.02465f
C12738 VPWR.n940 VGND 0.0762f
C12739 VPWR.t538 VGND 0.06535f
C12740 VPWR.t1549 VGND 0.07675f
C12741 VPWR.t1151 VGND 0.09955f
C12742 VPWR.t1542 VGND 0.02774f
C12743 VPWR.t1137 VGND 0.02465f
C12744 VPWR.n941 VGND 0.0762f
C12745 VPWR.n942 VGND 0.11584f
C12746 VPWR.n943 VGND 0.11584f
C12747 VPWR.t1152 VGND 0.02774f
C12748 VPWR.t815 VGND 0.02465f
C12749 VPWR.n944 VGND 0.0762f
C12750 VPWR.t905 VGND 0.06535f
C12751 VPWR.t814 VGND 0.07675f
C12752 VPWR.t930 VGND 0.09955f
C12753 VPWR.t807 VGND 0.02774f
C12754 VPWR.t889 VGND 0.02465f
C12755 VPWR.n945 VGND 0.0762f
C12756 VPWR.n946 VGND 0.11584f
C12757 VPWR.n947 VGND 0.11584f
C12758 VPWR.t931 VGND 0.02774f
C12759 VPWR.t950 VGND 0.02465f
C12760 VPWR.n948 VGND 0.0762f
C12761 VPWR.t1857 VGND 0.06535f
C12762 VPWR.t949 VGND 0.07675f
C12763 VPWR.t1232 VGND 0.09955f
C12764 VPWR.t942 VGND 0.02774f
C12765 VPWR.t1243 VGND 0.02465f
C12766 VPWR.n949 VGND 0.0762f
C12767 VPWR.n950 VGND 0.11584f
C12768 VPWR.n951 VGND 0.11584f
C12769 VPWR.t1233 VGND 0.02774f
C12770 VPWR.t1340 VGND 0.02465f
C12771 VPWR.n952 VGND 0.0762f
C12772 VPWR.t541 VGND 0.06535f
C12773 VPWR.t1339 VGND 0.07675f
C12774 VPWR.t1246 VGND 0.09955f
C12775 VPWR.t1317 VGND 0.02774f
C12776 VPWR.t1257 VGND 0.02465f
C12777 VPWR.n953 VGND 0.0762f
C12778 VPWR.n954 VGND 0.11584f
C12779 VPWR.n955 VGND 0.11584f
C12780 VPWR.t1247 VGND 0.02774f
C12781 VPWR.t1919 VGND 0.02465f
C12782 VPWR.n956 VGND 0.0762f
C12783 VPWR.t904 VGND 0.06535f
C12784 VPWR.t1918 VGND 0.07675f
C12785 VPWR.t733 VGND 0.09955f
C12786 VPWR.t1714 VGND 0.02774f
C12787 VPWR.t758 VGND 0.02465f
C12788 VPWR.n957 VGND 0.0762f
C12789 VPWR.n958 VGND 0.11584f
C12790 VPWR.n959 VGND 0.11584f
C12791 VPWR.t734 VGND 0.02774f
C12792 VPWR.t779 VGND 0.02465f
C12793 VPWR.n960 VGND 0.0762f
C12794 VPWR.t902 VGND 0.06535f
C12795 VPWR.t778 VGND 0.07675f
C12796 VPWR.t603 VGND 0.02774f
C12797 VPWR.t337 VGND 0.02465f
C12798 VPWR.n961 VGND 0.0762f
C12799 VPWR.t787 VGND 0.02774f
C12800 VPWR.t189 VGND 0.02465f
C12801 VPWR.n962 VGND 0.0762f
C12802 VPWR.t1103 VGND 0.12083f
C12803 VPWR.t1038 VGND 0.06535f
C12804 VPWR.t1193 VGND 0.07675f
C12805 VPWR.t1104 VGND 0.02774f
C12806 VPWR.t1194 VGND 0.02465f
C12807 VPWR.n963 VGND 0.0762f
C12808 VPWR.n964 VGND 0.01496f
C12809 VPWR.n966 VGND 0.0901f
C12810 VPWR.t854 VGND 0.09955f
C12811 VPWR.t1383 VGND 0.06535f
C12812 VPWR.t1904 VGND 0.07675f
C12813 VPWR.t855 VGND 0.02774f
C12814 VPWR.t1905 VGND 0.02465f
C12815 VPWR.n967 VGND 0.0762f
C12816 VPWR.n968 VGND 0.01496f
C12817 VPWR.n970 VGND 0.0901f
C12818 VPWR.t1900 VGND 0.09955f
C12819 VPWR.t1044 VGND 0.06535f
C12820 VPWR.t1476 VGND 0.07675f
C12821 VPWR.t1901 VGND 0.02774f
C12822 VPWR.t1477 VGND 0.02465f
C12823 VPWR.n971 VGND 0.0762f
C12824 VPWR.n972 VGND 0.01496f
C12825 VPWR.n974 VGND 0.0901f
C12826 VPWR.t1440 VGND 0.09955f
C12827 VPWR.t1043 VGND 0.06535f
C12828 VPWR.t996 VGND 0.07675f
C12829 VPWR.t1441 VGND 0.02774f
C12830 VPWR.t997 VGND 0.02465f
C12831 VPWR.n975 VGND 0.0762f
C12832 VPWR.n976 VGND 0.01496f
C12833 VPWR.n978 VGND 0.0901f
C12834 VPWR.t1280 VGND 0.09955f
C12835 VPWR.t940 VGND 0.06535f
C12836 VPWR.t1591 VGND 0.07675f
C12837 VPWR.t1281 VGND 0.02774f
C12838 VPWR.t1592 VGND 0.02465f
C12839 VPWR.n979 VGND 0.0762f
C12840 VPWR.n980 VGND 0.01496f
C12841 VPWR.n982 VGND 0.0901f
C12842 VPWR.t1701 VGND 0.09955f
C12843 VPWR.t1381 VGND 0.06535f
C12844 VPWR.t955 VGND 0.07675f
C12845 VPWR.t1702 VGND 0.02774f
C12846 VPWR.t956 VGND 0.02465f
C12847 VPWR.n983 VGND 0.0762f
C12848 VPWR.n984 VGND 0.01496f
C12849 VPWR.n986 VGND 0.0901f
C12850 VPWR.t917 VGND 0.09955f
C12851 VPWR.t1380 VGND 0.06535f
C12852 VPWR.t492 VGND 0.07675f
C12853 VPWR.t918 VGND 0.02774f
C12854 VPWR.t493 VGND 0.02465f
C12855 VPWR.n987 VGND 0.0762f
C12856 VPWR.n988 VGND 0.01496f
C12857 VPWR.n990 VGND 0.0901f
C12858 VPWR.t488 VGND 0.09955f
C12859 VPWR.t594 VGND 0.06535f
C12860 VPWR.t869 VGND 0.07675f
C12861 VPWR.t489 VGND 0.02774f
C12862 VPWR.t870 VGND 0.02465f
C12863 VPWR.n991 VGND 0.0762f
C12864 VPWR.n992 VGND 0.01496f
C12865 VPWR.n994 VGND 0.0901f
C12866 VPWR.t890 VGND 0.09955f
C12867 VPWR.t593 VGND 0.06535f
C12868 VPWR.t1187 VGND 0.07675f
C12869 VPWR.t891 VGND 0.02774f
C12870 VPWR.t1188 VGND 0.02465f
C12871 VPWR.n995 VGND 0.0762f
C12872 VPWR.n996 VGND 0.01496f
C12873 VPWR.n998 VGND 0.0901f
C12874 VPWR.t1183 VGND 0.09955f
C12875 VPWR.t1382 VGND 0.06535f
C12876 VPWR.t747 VGND 0.07675f
C12877 VPWR.t1184 VGND 0.02774f
C12878 VPWR.t748 VGND 0.02465f
C12879 VPWR.n999 VGND 0.0762f
C12880 VPWR.n1000 VGND 0.01496f
C12881 VPWR.n1002 VGND 0.0901f
C12882 VPWR.t725 VGND 0.09955f
C12883 VPWR.t1040 VGND 0.06535f
C12884 VPWR.t1617 VGND 0.07675f
C12885 VPWR.t726 VGND 0.02774f
C12886 VPWR.t1618 VGND 0.02465f
C12887 VPWR.n1003 VGND 0.0762f
C12888 VPWR.n1004 VGND 0.01496f
C12889 VPWR.n1006 VGND 0.0901f
C12890 VPWR.t1613 VGND 0.09955f
C12891 VPWR.t1039 VGND 0.06535f
C12892 VPWR.t1575 VGND 0.07675f
C12893 VPWR.t1614 VGND 0.02774f
C12894 VPWR.t1576 VGND 0.02465f
C12895 VPWR.n1007 VGND 0.0762f
C12896 VPWR.n1008 VGND 0.01496f
C12897 VPWR.n1010 VGND 0.0901f
C12898 VPWR.t1830 VGND 0.09955f
C12899 VPWR.t1379 VGND 0.06535f
C12900 VPWR.t1294 VGND 0.07675f
C12901 VPWR.t1831 VGND 0.02774f
C12902 VPWR.t1295 VGND 0.02465f
C12903 VPWR.n1011 VGND 0.0762f
C12904 VPWR.n1012 VGND 0.01496f
C12905 VPWR.n1014 VGND 0.0901f
C12906 VPWR.t1920 VGND 0.09955f
C12907 VPWR.t1046 VGND 0.06535f
C12908 VPWR.t414 VGND 0.07675f
C12909 VPWR.t1921 VGND 0.02774f
C12910 VPWR.t415 VGND 0.02465f
C12911 VPWR.n1015 VGND 0.0762f
C12912 VPWR.n1016 VGND 0.01496f
C12913 VPWR.n1018 VGND 0.0901f
C12914 VPWR.t402 VGND 0.09955f
C12915 VPWR.t1045 VGND 0.06535f
C12916 VPWR.t520 VGND 0.07675f
C12917 VPWR.t403 VGND 0.02774f
C12918 VPWR.t521 VGND 0.02465f
C12919 VPWR.n1019 VGND 0.0762f
C12920 VPWR.n1020 VGND 0.01496f
C12921 VPWR.n1022 VGND 0.0901f
C12922 VPWR.t786 VGND 0.09955f
C12923 VPWR.t592 VGND 0.06535f
C12924 VPWR.t188 VGND 0.11101f
C12925 VPWR.n1023 VGND 0.06343f
C12926 VPWR.n1024 VGND 0.01496f
C12927 VPWR.n1025 VGND 0.11584f
C12928 VPWR.n1026 VGND 4.86825f
C12929 VPWR.n1027 VGND 0.05468f
C12930 VPWR.n1028 VGND -0.01553f
C12931 VPWR.t190 VGND 0.01018f
C12932 VPWR.n1029 VGND 0.02533f
C12933 VPWR.t192 VGND 0.02231f
C12934 VPWR.n1031 VGND 0.04766f
C12935 VPWR.t300 VGND 0.02465f
C12936 VPWR.n1032 VGND 0.03907f
C12937 VPWR.t788 VGND 0.07675f
C12938 VPWR.t82 VGND 0.01018f
C12939 VPWR.n1033 VGND 0.02533f
C12940 VPWR.t84 VGND 0.02231f
C12941 VPWR.n1035 VGND 0.04766f
C12942 VPWR.t789 VGND 0.02465f
C12943 VPWR.n1036 VGND 0.03907f
C12944 VPWR.n1037 VGND -0.01553f
C12945 VPWR.n1038 VGND 0.05468f
C12946 VPWR.t41 VGND 0.01033f
C12947 VPWR.n1039 VGND 0.02305f
C12948 VPWR.n1040 VGND 0.01579f
C12949 VPWR.n1041 VGND 0.05199f
C12950 VPWR.n1042 VGND 0.08114f
C12951 VPWR.n1043 VGND 0.0453f
C12952 VPWR.n1044 VGND 0.05468f
C12953 VPWR.n1045 VGND -0.01553f
C12954 VPWR.t168 VGND 0.01018f
C12955 VPWR.n1046 VGND 0.02533f
C12956 VPWR.t170 VGND 0.02231f
C12957 VPWR.n1048 VGND 0.04766f
C12958 VPWR.t1843 VGND 0.02465f
C12959 VPWR.n1049 VGND 0.03907f
C12960 VPWR.t1842 VGND 0.07675f
C12961 VPWR.t33 VGND 0.09955f
C12962 VPWR.t209 VGND 0.01018f
C12963 VPWR.n1050 VGND 0.02533f
C12964 VPWR.t211 VGND 0.02231f
C12965 VPWR.n1052 VGND 0.04766f
C12966 VPWR.t1074 VGND 0.02465f
C12967 VPWR.n1053 VGND 0.03907f
C12968 VPWR.n1055 VGND 0.16128f
C12969 VPWR.n1056 VGND 0.06953f
C12970 VPWR.n1057 VGND 0.02861f
C12971 VPWR.t264 VGND 0.02774f
C12972 VPWR.t256 VGND 0.02465f
C12973 VPWR.n1058 VGND 0.0762f
C12974 VPWR.t255 VGND 0.07675f
C12975 VPWR.t10 VGND 0.09955f
C12976 VPWR.t292 VGND 0.02774f
C12977 VPWR.t284 VGND 0.02465f
C12978 VPWR.n1059 VGND 0.0762f
C12979 VPWR.t11 VGND 0.02774f
C12980 VPWR.t135 VGND 0.02465f
C12981 VPWR.n1061 VGND 0.0762f
C12982 VPWR.t13 VGND 0.06535f
C12983 VPWR.t134 VGND 0.11101f
C12984 VPWR.n1062 VGND 0.0634f
C12985 VPWR.n1063 VGND 0.01414f
C12986 VPWR.t133 VGND 0.01021f
C12987 VPWR.n1064 VGND 0.02492f
C12988 VPWR.n1065 VGND 0.02734f
C12989 VPWR.n1067 VGND 0.01517f
C12990 VPWR.n1068 VGND 0.14641f
C12991 VPWR.t254 VGND 0.01021f
C12992 VPWR.n1069 VGND 0.02492f
C12993 VPWR.n1070 VGND 0.02734f
C12994 VPWR.n1071 VGND 0.01427f
C12995 VPWR.n1074 VGND 0.01427f
C12996 VPWR.t260 VGND 0.01033f
C12997 VPWR.n1076 VGND 0.02304f
C12998 VPWR.n1077 VGND 0.02346f
C12999 VPWR.n1078 VGND 0.01517f
C13000 VPWR.n1079 VGND 0.14641f
C13001 VPWR.t362 VGND 0.01021f
C13002 VPWR.n1080 VGND 0.02492f
C13003 VPWR.n1081 VGND 0.02734f
C13004 VPWR.n1082 VGND 0.01427f
C13005 VPWR.n1084 VGND 0.01427f
C13006 VPWR.t368 VGND 0.01033f
C13007 VPWR.n1086 VGND 0.02304f
C13008 VPWR.n1087 VGND 0.02346f
C13009 VPWR.n1088 VGND 0.01517f
C13010 VPWR.n1089 VGND 0.14641f
C13011 VPWR.t354 VGND 0.01021f
C13012 VPWR.n1090 VGND 0.02492f
C13013 VPWR.n1091 VGND 0.02734f
C13014 VPWR.n1092 VGND 0.01427f
C13015 VPWR.n1094 VGND 0.01427f
C13016 VPWR.t87 VGND 0.01033f
C13017 VPWR.n1096 VGND 0.02304f
C13018 VPWR.n1097 VGND 0.02346f
C13019 VPWR.n1098 VGND 0.01517f
C13020 VPWR.n1099 VGND 0.14641f
C13021 VPWR.t59 VGND 0.01021f
C13022 VPWR.n1100 VGND 0.02492f
C13023 VPWR.n1101 VGND 0.02734f
C13024 VPWR.n1102 VGND 0.01427f
C13025 VPWR.n1104 VGND 0.01427f
C13026 VPWR.t171 VGND 0.01033f
C13027 VPWR.n1106 VGND 0.02304f
C13028 VPWR.n1107 VGND 0.02346f
C13029 VPWR.n1108 VGND 0.01517f
C13030 VPWR.n1109 VGND 0.0221f
C13031 VPWR.t165 VGND 0.01021f
C13032 VPWR.n1110 VGND 0.02492f
C13033 VPWR.n1111 VGND 0.02734f
C13034 VPWR.n1112 VGND 0.01517f
C13035 VPWR.t311 VGND 0.01018f
C13036 VPWR.n1114 VGND 0.02594f
C13037 VPWR.n1115 VGND 0.01639f
C13038 VPWR.t301 VGND 0.01033f
C13039 VPWR.n1116 VGND 0.02304f
C13040 VPWR.n1117 VGND 0.02346f
C13041 VPWR.n1118 VGND 0.01479f
C13042 VPWR.t29 VGND 0.01021f
C13043 VPWR.n1119 VGND 0.02492f
C13044 VPWR.n1120 VGND 0.02734f
C13045 VPWR.t313 VGND 0.02774f
C13046 VPWR.t31 VGND 0.02465f
C13047 VPWR.n1122 VGND 0.0762f
C13048 VPWR.t312 VGND 0.12083f
C13049 VPWR.t302 VGND 0.06535f
C13050 VPWR.t30 VGND 0.07675f
C13051 VPWR.t182 VGND 0.09955f
C13052 VPWR.t81 VGND 0.02774f
C13053 VPWR.t167 VGND 0.02465f
C13054 VPWR.n1123 VGND 0.0762f
C13055 VPWR.t181 VGND 0.01018f
C13056 VPWR.n1125 VGND 0.02594f
C13057 VPWR.n1126 VGND 0.03075f
C13058 VPWR.n1127 VGND 0.02861f
C13059 VPWR.n1128 VGND 0.11584f
C13060 VPWR.n1130 VGND 0.01496f
C13061 VPWR.n1131 VGND 0.05468f
C13062 VPWR.n1132 VGND 0.0453f
C13063 VPWR.t352 VGND 0.01033f
C13064 VPWR.n1133 VGND 0.02305f
C13065 VPWR.n1134 VGND 0.01579f
C13066 VPWR.n1135 VGND 0.05199f
C13067 VPWR.n1136 VGND 0.08114f
C13068 VPWR.n1137 VGND 0.05468f
C13069 VPWR.n1138 VGND 0.05468f
C13070 VPWR.n1139 VGND 0.05468f
C13071 VPWR.n1140 VGND 0.05468f
C13072 VPWR.n1141 VGND 0.05468f
C13073 VPWR.n1142 VGND 0.05468f
C13074 VPWR.n1143 VGND 0.0453f
C13075 VPWR.n1145 VGND -0.01553f
C13076 VPWR.t295 VGND 0.01018f
C13077 VPWR.n1146 VGND 0.02533f
C13078 VPWR.t297 VGND 0.02231f
C13079 VPWR.n1148 VGND 0.04766f
C13080 VPWR.t1873 VGND 0.02465f
C13081 VPWR.n1149 VGND 0.03907f
C13082 VPWR.t1872 VGND 0.07675f
C13083 VPWR.t42 VGND 0.06535f
C13084 VPWR.t169 VGND 0.09955f
C13085 VPWR.t38 VGND 0.01018f
C13086 VPWR.n1150 VGND 0.02533f
C13087 VPWR.t40 VGND 0.02231f
C13088 VPWR.n1152 VGND 0.04766f
C13089 VPWR.t1346 VGND 0.02465f
C13090 VPWR.n1153 VGND 0.03907f
C13091 VPWR.t279 VGND 0.01018f
C13092 VPWR.n1156 VGND 0.02533f
C13093 VPWR.t281 VGND 0.02231f
C13094 VPWR.n1158 VGND 0.04766f
C13095 VPWR.t557 VGND 0.02465f
C13096 VPWR.n1159 VGND 0.03907f
C13097 VPWR.t896 VGND 0.07675f
C13098 VPWR.t138 VGND 0.01018f
C13099 VPWR.n1160 VGND 0.02533f
C13100 VPWR.t140 VGND 0.02231f
C13101 VPWR.n1162 VGND 0.04766f
C13102 VPWR.t897 VGND 0.02465f
C13103 VPWR.n1163 VGND 0.03907f
C13104 VPWR.t16 VGND 0.01018f
C13105 VPWR.n1166 VGND 0.02533f
C13106 VPWR.t18 VGND 0.02231f
C13107 VPWR.n1168 VGND 0.04766f
C13108 VPWR.t821 VGND 0.02465f
C13109 VPWR.n1169 VGND 0.03907f
C13110 VPWR.t1142 VGND 0.07675f
C13111 VPWR.t265 VGND 0.01018f
C13112 VPWR.n1170 VGND 0.02533f
C13113 VPWR.t267 VGND 0.02231f
C13114 VPWR.n1172 VGND 0.04766f
C13115 VPWR.t1143 VGND 0.02465f
C13116 VPWR.n1173 VGND 0.03907f
C13117 VPWR.t76 VGND 0.01018f
C13118 VPWR.n1176 VGND 0.02594f
C13119 VPWR.n1177 VGND 0.03075f
C13120 VPWR.n1178 VGND 0.02861f
C13121 VPWR.t66 VGND 0.02774f
C13122 VPWR.t61 VGND 0.02465f
C13123 VPWR.n1179 VGND 0.0762f
C13124 VPWR.t172 VGND 0.06535f
C13125 VPWR.t179 VGND 0.07675f
C13126 VPWR.t183 VGND 0.02774f
C13127 VPWR.t180 VGND 0.02465f
C13128 VPWR.n1180 VGND 0.0762f
C13129 VPWR.n1182 VGND 0.0901f
C13130 VPWR.t347 VGND 0.09955f
C13131 VPWR.t213 VGND 0.06535f
C13132 VPWR.t339 VGND 0.07675f
C13133 VPWR.t348 VGND 0.02774f
C13134 VPWR.t340 VGND 0.02465f
C13135 VPWR.n1183 VGND 0.0762f
C13136 VPWR.n1185 VGND 0.0901f
C13137 VPWR.t65 VGND 0.09955f
C13138 VPWR.t321 VGND 0.06535f
C13139 VPWR.t60 VGND 0.07675f
C13140 VPWR.t137 VGND 0.06535f
C13141 VPWR.t263 VGND 0.09955f
C13142 VPWR.t26 VGND 0.02774f
C13143 VPWR.t127 VGND 0.02465f
C13144 VPWR.n1186 VGND 0.0762f
C13145 VPWR.n1188 VGND 0.0901f
C13146 VPWR.t126 VGND 0.07675f
C13147 VPWR.t111 VGND 0.06535f
C13148 VPWR.t25 VGND 0.09955f
C13149 VPWR.t5 VGND 0.02774f
C13150 VPWR.t383 VGND 0.02465f
C13151 VPWR.n1189 VGND 0.0762f
C13152 VPWR.n1191 VGND 0.0901f
C13153 VPWR.t382 VGND 0.07675f
C13154 VPWR.t261 VGND 0.06535f
C13155 VPWR.t4 VGND 0.09955f
C13156 VPWR.t259 VGND 0.02774f
C13157 VPWR.t364 VGND 0.02465f
C13158 VPWR.n1192 VGND 0.0762f
C13159 VPWR.t3 VGND 0.01018f
C13160 VPWR.n1194 VGND 0.02594f
C13161 VPWR.n1195 VGND 0.03075f
C13162 VPWR.n1196 VGND 0.02861f
C13163 VPWR.n1197 VGND 0.01427f
C13164 VPWR.n1199 VGND 0.0901f
C13165 VPWR.t363 VGND 0.07675f
C13166 VPWR.t239 VGND 0.06535f
C13167 VPWR.t258 VGND 0.09955f
C13168 VPWR.t132 VGND 0.02774f
C13169 VPWR.t205 VGND 0.02465f
C13170 VPWR.n1200 VGND 0.0762f
C13171 VPWR.n1202 VGND 0.0901f
C13172 VPWR.t204 VGND 0.07675f
C13173 VPWR.t86 VGND 0.06535f
C13174 VPWR.t131 VGND 0.09955f
C13175 VPWR.t106 VGND 0.02774f
C13176 VPWR.t101 VGND 0.02465f
C13177 VPWR.n1203 VGND 0.0762f
C13178 VPWR.n1205 VGND 0.0901f
C13179 VPWR.t100 VGND 0.07675f
C13180 VPWR.t369 VGND 0.06535f
C13181 VPWR.t105 VGND 0.09955f
C13182 VPWR.t345 VGND 0.02774f
C13183 VPWR.t356 VGND 0.02465f
C13184 VPWR.n1206 VGND 0.0762f
C13185 VPWR.t104 VGND 0.01018f
C13186 VPWR.n1208 VGND 0.02594f
C13187 VPWR.n1209 VGND 0.03075f
C13188 VPWR.n1210 VGND 0.02861f
C13189 VPWR.n1211 VGND 0.01427f
C13190 VPWR.n1213 VGND 0.0901f
C13191 VPWR.t355 VGND 0.07675f
C13192 VPWR.t326 VGND 0.06535f
C13193 VPWR.t344 VGND 0.09955f
C13194 VPWR.t237 VGND 0.02774f
C13195 VPWR.t319 VGND 0.02465f
C13196 VPWR.n1214 VGND 0.0762f
C13197 VPWR.n1216 VGND 0.0901f
C13198 VPWR.t318 VGND 0.07675f
C13199 VPWR.t103 VGND 0.06535f
C13200 VPWR.t236 VGND 0.09955f
C13201 VPWR.t78 VGND 0.02774f
C13202 VPWR.t208 VGND 0.02465f
C13203 VPWR.n1217 VGND 0.0762f
C13204 VPWR.n1219 VGND 0.0901f
C13205 VPWR.t207 VGND 0.07675f
C13206 VPWR.t88 VGND 0.06535f
C13207 VPWR.t77 VGND 0.09955f
C13208 VPWR.n1220 VGND 0.0901f
C13209 VPWR.n1222 VGND 0.01427f
C13210 VPWR.t243 VGND 0.01018f
C13211 VPWR.n1224 VGND 0.02533f
C13212 VPWR.t245 VGND 0.02231f
C13213 VPWR.n1226 VGND 0.04766f
C13214 VPWR.t591 VGND 0.02465f
C13215 VPWR.n1227 VGND 0.03907f
C13216 VPWR.t108 VGND 0.12083f
C13217 VPWR.t93 VGND 0.06535f
C13218 VPWR.t429 VGND 0.07675f
C13219 VPWR.t107 VGND 0.01018f
C13220 VPWR.n1228 VGND 0.02533f
C13221 VPWR.t109 VGND 0.02231f
C13222 VPWR.n1230 VGND 0.04766f
C13223 VPWR.t430 VGND 0.02465f
C13224 VPWR.n1231 VGND 0.03907f
C13225 VPWR.n1232 VGND -0.01553f
C13226 VPWR.n1233 VGND 0.03902f
C13227 VPWR.t580 VGND 0.81233f
C13228 VPWR.n1234 VGND 0.44305f
C13229 VPWR.t566 VGND 0.81233f
C13230 VPWR.n1235 VGND 0.34456f
C13231 VPWR.n1236 VGND 0.24212f
C13232 VPWR.t1216 VGND 0.04759f
C13233 VPWR.t1057 VGND 0.01193f
C13234 VPWR.t1060 VGND 0.01193f
C13235 VPWR.n1238 VGND 0.02619f
C13236 VPWR.t1742 VGND 0.01193f
C13237 VPWR.t581 VGND 0.01193f
C13238 VPWR.n1239 VGND 0.02615f
C13239 VPWR.t1738 VGND 0.01193f
C13240 VPWR.t1737 VGND 0.01193f
C13241 VPWR.n1240 VGND 0.02615f
C13242 VPWR.n1241 VGND 0.08676f
C13243 VPWR.n1242 VGND 0.15138f
C13244 VPWR.n1243 VGND 0.04793f
C13245 VPWR.n1244 VGND 0.0352f
C13246 VPWR.t1734 VGND 0.01193f
C13247 VPWR.t1739 VGND 0.01193f
C13248 VPWR.n1245 VGND 0.02619f
C13249 VPWR.n1246 VGND 0.10742f
C13250 VPWR.n1248 VGND 0.01357f
C13251 VPWR.n1249 VGND 0.01591f
C13252 VPWR.n1250 VGND 0.02333f
C13253 VPWR.t1215 VGND 0.04759f
C13254 VPWR.n1251 VGND 0.12538f
C13255 VPWR.n1252 VGND 0.01006f
C13256 VPWR.t583 VGND 0.04758f
C13257 VPWR.t567 VGND 0.04758f
C13258 VPWR.n1253 VGND 0.11195f
C13259 VPWR.n1254 VGND 0.27944f
C13260 VPWR.n1255 VGND 1.36622f
C13261 VPWR.n1256 VGND 0.03902f
C13262 VPWR.t494 VGND 0.81233f
C13263 VPWR.n1257 VGND 0.44305f
C13264 VPWR.t637 VGND 0.81233f
C13265 VPWR.n1258 VGND 0.34456f
C13266 VPWR.n1259 VGND 0.2443f
C13267 VPWR.t501 VGND 0.01193f
C13268 VPWR.t499 VGND 0.01193f
C13269 VPWR.n1261 VGND 0.02619f
C13270 VPWR.t498 VGND 0.01193f
C13271 VPWR.t495 VGND 0.01193f
C13272 VPWR.n1262 VGND 0.02615f
C13273 VPWR.t980 VGND 0.01193f
C13274 VPWR.t981 VGND 0.01193f
C13275 VPWR.n1263 VGND 0.02615f
C13276 VPWR.n1264 VGND 0.08676f
C13277 VPWR.n1265 VGND 0.15138f
C13278 VPWR.n1266 VGND 0.04793f
C13279 VPWR.n1267 VGND 0.0352f
C13280 VPWR.t1538 VGND 0.01193f
C13281 VPWR.t1289 VGND 0.01193f
C13282 VPWR.n1268 VGND 0.02619f
C13283 VPWR.n1269 VGND 0.10742f
C13284 VPWR.n1271 VGND 0.01357f
C13285 VPWR.n1272 VGND 0.01591f
C13286 VPWR.n1273 VGND 0.0229f
C13287 VPWR.t1217 VGND 0.04752f
C13288 VPWR.n1275 VGND 0.0508f
C13289 VPWR.t1413 VGND 0.04762f
C13290 VPWR.n1277 VGND 0.07585f
C13291 VPWR.n1278 VGND 0.27944f
C13292 VPWR.n1279 VGND 1.36622f
C13293 VPWR.n1280 VGND 0.03902f
C13294 VPWR.t584 VGND 0.81233f
C13295 VPWR.n1281 VGND 0.44305f
C13296 VPWR.t421 VGND 0.81233f
C13297 VPWR.n1282 VGND 0.34456f
C13298 VPWR.n1283 VGND 0.2443f
C13299 VPWR.t1212 VGND 0.01193f
C13300 VPWR.t1210 VGND 0.01193f
C13301 VPWR.n1285 VGND 0.02619f
C13302 VPWR.t1209 VGND 0.01193f
C13303 VPWR.t1208 VGND 0.01193f
C13304 VPWR.n1286 VGND 0.02615f
C13305 VPWR.t1405 VGND 0.01193f
C13306 VPWR.t1412 VGND 0.01193f
C13307 VPWR.n1287 VGND 0.02615f
C13308 VPWR.n1288 VGND 0.08676f
C13309 VPWR.n1289 VGND 0.15138f
C13310 VPWR.n1290 VGND 0.04793f
C13311 VPWR.n1291 VGND 0.0352f
C13312 VPWR.t1409 VGND 0.01193f
C13313 VPWR.t1406 VGND 0.01193f
C13314 VPWR.n1292 VGND 0.02619f
C13315 VPWR.n1293 VGND 0.10742f
C13316 VPWR.n1295 VGND 0.01357f
C13317 VPWR.n1296 VGND 0.01591f
C13318 VPWR.n1297 VGND 0.0229f
C13319 VPWR.n1298 VGND 0.01164f
C13320 VPWR.n1299 VGND 0.01089f
C13321 VPWR.t585 VGND 0.04762f
C13322 VPWR.t568 VGND 0.04762f
C13323 VPWR.n1300 VGND 0.14066f
C13324 VPWR.n1301 VGND 0.27944f
C13325 VPWR.n1302 VGND 1.36622f
C13326 VPWR.t1728 VGND 0.04755f
C13327 VPWR.t1070 VGND 0.04762f
C13328 VPWR.t1730 VGND 0.04722f
C13329 VPWR.n1303 VGND 0.12244f
C13330 VPWR.t1227 VGND 0.04668f
C13331 VPWR.n1304 VGND 0.05641f
C13332 VPWR.n1305 VGND 0.03902f
C13333 VPWR.t619 VGND 0.04494f
C13334 VPWR.n1306 VGND 0.04274f
C13335 VPWR.t442 VGND 0.01193f
C13336 VPWR.t1421 VGND 0.01193f
C13337 VPWR.n1307 VGND 0.02607f
C13338 VPWR.t423 VGND 0.04175f
C13339 VPWR.n1308 VGND 0.06262f
C13340 VPWR.n1309 VGND 0.03902f
C13341 VPWR.t1224 VGND 0.04757f
C13342 VPWR.n1310 VGND 0.05989f
C13343 VPWR.n1311 VGND 0.0229f
C13344 VPWR.n1312 VGND 0.03902f
C13345 VPWR.n1313 VGND 0.01006f
C13346 VPWR.t636 VGND 0.01193f
C13347 VPWR.t639 VGND 0.01193f
C13348 VPWR.n1314 VGND 0.02607f
C13349 VPWR.n1315 VGND 0.0382f
C13350 VPWR.n1316 VGND 0.01006f
C13351 VPWR.n1317 VGND 0.02927f
C13352 VPWR.n1318 VGND 0.02927f
C13353 VPWR.n1319 VGND 0.03902f
C13354 VPWR.t438 VGND 0.01193f
C13355 VPWR.t615 VGND 0.01193f
C13356 VPWR.n1321 VGND 0.02607f
C13357 VPWR.n1322 VGND 0.03001f
C13358 VPWR.t1229 VGND 0.01193f
C13359 VPWR.t864 VGND 0.01193f
C13360 VPWR.n1323 VGND 0.02607f
C13361 VPWR.n1324 VGND 0.03317f
C13362 VPWR.n1326 VGND 0.03542f
C13363 VPWR.n1327 VGND 0.01336f
C13364 VPWR.t1047 VGND 0.04001f
C13365 VPWR.t1727 VGND 0.09002f
C13366 VPWR.t1069 VGND 0.10503f
C13367 VPWR.t1729 VGND 0.19505f
C13368 VPWR.t1223 VGND 0.10495f
C13369 VPWR.t638 VGND 0.11913f
C13370 VPWR.t635 VGND 0.11582f
C13371 VPWR.t1420 VGND 0.18523f
C13372 VPWR.t441 VGND 0.15754f
C13373 VPWR.t422 VGND 0.10503f
C13374 VPWR.t614 VGND 0.10503f
C13375 VPWR.t863 VGND 0.10503f
C13376 VPWR.t437 VGND 0.10503f
C13377 VPWR.t1228 VGND 0.10503f
C13378 VPWR.t618 VGND 0.10503f
C13379 VPWR.t1226 VGND 0.10378f
C13380 VPWR.n1329 VGND 0.35694f
C13381 VPWR.n1330 VGND 0.14503f
C13382 VPWR.n1331 VGND 0.01591f
C13383 VPWR.n1332 VGND 0.02927f
C13384 VPWR.n1333 VGND 0.0352f
C13385 VPWR.n1335 VGND 0.05293f
C13386 VPWR.n1336 VGND 0.26353f
C13387 VPWR.n1337 VGND 1.36622f
C13388 VPWR.t569 VGND 0.04678f
C13389 VPWR.t984 VGND 0.04665f
C13390 VPWR.t1374 VGND 0.04758f
C13391 VPWR.n1338 VGND 0.0663f
C13392 VPWR.t1743 VGND 0.04542f
C13393 VPWR.t1740 VGND 0.04542f
C13394 VPWR.n1339 VGND 0.08241f
C13395 VPWR.n1340 VGND 0.03902f
C13396 VPWR.n1342 VGND 0.03902f
C13397 VPWR.t1058 VGND 0.01193f
C13398 VPWR.t710 VGND 0.01193f
C13399 VPWR.n1343 VGND 0.02607f
C13400 VPWR.t1741 VGND 0.01193f
C13401 VPWR.t1522 VGND 0.01193f
C13402 VPWR.n1344 VGND 0.02607f
C13403 VPWR.n1345 VGND 0.05311f
C13404 VPWR.t1524 VGND 0.04757f
C13405 VPWR.t641 VGND 0.04757f
C13406 VPWR.n1346 VGND 0.10964f
C13407 VPWR.n1347 VGND 0.0229f
C13408 VPWR.n1348 VGND 0.03902f
C13409 VPWR.n1349 VGND 0.01006f
C13410 VPWR.t1398 VGND 0.01193f
C13411 VPWR.t426 VGND 0.01193f
C13412 VPWR.n1350 VGND 0.02607f
C13413 VPWR.t1416 VGND 0.01193f
C13414 VPWR.t1419 VGND 0.01193f
C13415 VPWR.n1351 VGND 0.02607f
C13416 VPWR.n1352 VGND 0.06002f
C13417 VPWR.n1353 VGND 0.01006f
C13418 VPWR.n1354 VGND 0.03902f
C13419 VPWR.n1355 VGND 0.03902f
C13420 VPWR.n1356 VGND 0.03902f
C13421 VPWR.t582 VGND 0.01193f
C13422 VPWR.t1059 VGND 0.01193f
C13423 VPWR.n1358 VGND 0.02607f
C13424 VPWR.t1736 VGND 0.01193f
C13425 VPWR.t1735 VGND 0.01193f
C13426 VPWR.n1359 VGND 0.02607f
C13427 VPWR.n1360 VGND 0.05311f
C13428 VPWR.n1363 VGND 0.03902f
C13429 VPWR.n1364 VGND 0.02927f
C13430 VPWR.t425 VGND 0.81233f
C13431 VPWR.n1366 VGND 0.44305f
C13432 VPWR.t640 VGND 0.81233f
C13433 VPWR.n1367 VGND 0.34456f
C13434 VPWR.n1368 VGND 0.24212f
C13435 VPWR.n1369 VGND 0.01591f
C13436 VPWR.n1370 VGND 0.02927f
C13437 VPWR.n1371 VGND 0.03542f
C13438 VPWR.n1373 VGND 0.04852f
C13439 VPWR.n1374 VGND 0.06572f
C13440 VPWR.n1375 VGND 0.26332f
C13441 VPWR.n1376 VGND 1.36622f
C13442 VPWR.t1071 VGND 0.04752f
C13443 VPWR.t1072 VGND 0.04752f
C13444 VPWR.n1377 VGND 0.01164f
C13445 VPWR.t497 VGND 0.04542f
C13446 VPWR.t1288 VGND 0.04542f
C13447 VPWR.n1378 VGND 0.08241f
C13448 VPWR.n1379 VGND 0.03902f
C13449 VPWR.n1381 VGND 0.03902f
C13450 VPWR.t502 VGND 0.01193f
C13451 VPWR.t1525 VGND 0.01193f
C13452 VPWR.n1382 VGND 0.02607f
C13453 VPWR.t1726 VGND 0.01193f
C13454 VPWR.t643 VGND 0.01193f
C13455 VPWR.n1383 VGND 0.02607f
C13456 VPWR.n1384 VGND 0.05311f
C13457 VPWR.t708 VGND 0.04757f
C13458 VPWR.t1521 VGND 0.04757f
C13459 VPWR.n1385 VGND 0.10964f
C13460 VPWR.n1386 VGND 0.0229f
C13461 VPWR.n1387 VGND 0.03902f
C13462 VPWR.n1388 VGND 0.01006f
C13463 VPWR.t1418 VGND 0.01193f
C13464 VPWR.t862 VGND 0.01193f
C13465 VPWR.n1389 VGND 0.02607f
C13466 VPWR.t709 VGND 0.01193f
C13467 VPWR.t1400 VGND 0.01193f
C13468 VPWR.n1390 VGND 0.02607f
C13469 VPWR.n1391 VGND 0.06002f
C13470 VPWR.n1392 VGND 0.01006f
C13471 VPWR.n1393 VGND 0.03902f
C13472 VPWR.n1394 VGND 0.03902f
C13473 VPWR.n1395 VGND 0.03902f
C13474 VPWR.t503 VGND 0.01193f
C13475 VPWR.t500 VGND 0.01193f
C13476 VPWR.n1397 VGND 0.02607f
C13477 VPWR.t1725 VGND 0.01193f
C13478 VPWR.t1537 VGND 0.01193f
C13479 VPWR.n1398 VGND 0.02607f
C13480 VPWR.n1399 VGND 0.05311f
C13481 VPWR.n1402 VGND 0.03902f
C13482 VPWR.n1403 VGND 0.02927f
C13483 VPWR.t496 VGND 0.81233f
C13484 VPWR.n1405 VGND 0.44305f
C13485 VPWR.t642 VGND 0.81233f
C13486 VPWR.n1406 VGND 0.34456f
C13487 VPWR.n1407 VGND 0.2443f
C13488 VPWR.n1408 VGND 0.01591f
C13489 VPWR.n1409 VGND 0.02927f
C13490 VPWR.n1410 VGND 0.03542f
C13491 VPWR.n1412 VGND 0.09606f
C13492 VPWR.n1413 VGND 0.26757f
C13493 VPWR.n1414 VGND 1.36622f
C13494 VPWR.t1211 VGND 0.04542f
C13495 VPWR.t1407 VGND 0.04542f
C13496 VPWR.n1415 VGND 0.08241f
C13497 VPWR.n1416 VGND 0.03902f
C13498 VPWR.n1418 VGND 0.03902f
C13499 VPWR.t1206 VGND 0.01193f
C13500 VPWR.t711 VGND 0.01193f
C13501 VPWR.n1419 VGND 0.02607f
C13502 VPWR.t1408 VGND 0.01193f
C13503 VPWR.t1222 VGND 0.01193f
C13504 VPWR.n1420 VGND 0.02607f
C13505 VPWR.n1421 VGND 0.05311f
C13506 VPWR.t1526 VGND 0.04757f
C13507 VPWR.t866 VGND 0.04757f
C13508 VPWR.n1422 VGND 0.10964f
C13509 VPWR.n1423 VGND 0.0229f
C13510 VPWR.n1424 VGND 0.03902f
C13511 VPWR.n1425 VGND 0.01006f
C13512 VPWR.t1399 VGND 0.01193f
C13513 VPWR.t428 VGND 0.01193f
C13514 VPWR.n1426 VGND 0.02607f
C13515 VPWR.t1225 VGND 0.01193f
C13516 VPWR.t1520 VGND 0.01193f
C13517 VPWR.n1427 VGND 0.02607f
C13518 VPWR.n1428 VGND 0.06002f
C13519 VPWR.n1429 VGND 0.01006f
C13520 VPWR.n1430 VGND 0.03902f
C13521 VPWR.n1431 VGND 0.03902f
C13522 VPWR.n1432 VGND 0.03902f
C13523 VPWR.t1207 VGND 0.01193f
C13524 VPWR.t1205 VGND 0.01193f
C13525 VPWR.n1434 VGND 0.02607f
C13526 VPWR.t1411 VGND 0.01193f
C13527 VPWR.t1410 VGND 0.01193f
C13528 VPWR.n1435 VGND 0.02607f
C13529 VPWR.n1436 VGND 0.05311f
C13530 VPWR.n1439 VGND 0.03902f
C13531 VPWR.n1440 VGND 0.02927f
C13532 VPWR.t427 VGND 0.62314f
C13533 VPWR.n1442 VGND 0.35652f
C13534 VPWR.t865 VGND 0.62314f
C13535 VPWR.n1443 VGND 0.27936f
C13536 VPWR.n1444 VGND 0.2342f
C13537 VPWR.n1445 VGND 0.35804f
C13538 VPWR.n1446 VGND 5.20598f
C13539 VPWR.n1447 VGND 7.62137f
C13540 VPWR.n1448 VGND 0.06953f
C13541 VPWR.n1449 VGND 0.91576f
C13542 VPWR.n1450 VGND 0.84042f
C13543 VPWR.n1451 VGND 0.05397f
C13544 VPWR.n1452 VGND 0.0453f
C13545 VPWR.t92 VGND 0.01033f
C13546 VPWR.n1453 VGND 0.02305f
C13547 VPWR.n1454 VGND 0.01579f
C13548 VPWR.n1455 VGND 0.05199f
C13549 VPWR.n1456 VGND 0.06463f
C13550 VPWR.n1457 VGND 0.07639f
C13551 VPWR.t223 VGND 0.01033f
C13552 VPWR.n1458 VGND 0.02305f
C13553 VPWR.n1459 VGND 0.01579f
C13554 VPWR.n1460 VGND 0.05199f
C13555 VPWR.n1461 VGND 0.08114f
C13556 VPWR.n1462 VGND 0.07639f
C13557 VPWR.n1463 VGND 0.05468f
C13558 VPWR.n1464 VGND 0.0453f
C13559 VPWR.n1465 VGND 0.11584f
C13560 VPWR.n1466 VGND 0.01496f
C13561 VPWR.n1468 VGND 0.0901f
C13562 VPWR.t269 VGND 0.09955f
C13563 VPWR.t224 VGND 0.06535f
C13564 VPWR.t1563 VGND 0.07675f
C13565 VPWR.t268 VGND 0.01018f
C13566 VPWR.n1469 VGND 0.02533f
C13567 VPWR.t270 VGND 0.02231f
C13568 VPWR.n1471 VGND 0.04766f
C13569 VPWR.t1564 VGND 0.02465f
C13570 VPWR.n1472 VGND 0.03907f
C13571 VPWR.n1473 VGND 0.01496f
C13572 VPWR.n1475 VGND 0.0901f
C13573 VPWR.t371 VGND 0.09955f
C13574 VPWR.t353 VGND 0.06535f
C13575 VPWR.t1490 VGND 0.07675f
C13576 VPWR.t370 VGND 0.01018f
C13577 VPWR.n1476 VGND 0.02533f
C13578 VPWR.t372 VGND 0.02231f
C13579 VPWR.n1478 VGND 0.04766f
C13580 VPWR.t1491 VGND 0.02465f
C13581 VPWR.n1479 VGND 0.03907f
C13582 VPWR.n1481 VGND 0.0901f
C13583 VPWR.t142 VGND 0.09955f
C13584 VPWR.t15 VGND 0.06535f
C13585 VPWR.t1504 VGND 0.07675f
C13586 VPWR.t141 VGND 0.01018f
C13587 VPWR.n1482 VGND 0.02533f
C13588 VPWR.t143 VGND 0.02231f
C13589 VPWR.n1484 VGND 0.04766f
C13590 VPWR.t1505 VGND 0.02465f
C13591 VPWR.n1485 VGND 0.03907f
C13592 VPWR.n1487 VGND 0.06953f
C13593 VPWR.n1488 VGND -0.01553f
C13594 VPWR.n1489 VGND 0.11584f
C13595 VPWR.n1490 VGND 0.01496f
C13596 VPWR.n1492 VGND 0.0901f
C13597 VPWR.t244 VGND 0.09955f
C13598 VPWR.t119 VGND 0.06535f
C13599 VPWR.t590 VGND 0.07675f
C13600 VPWR.t274 VGND 0.06535f
C13601 VPWR.t266 VGND 0.09955f
C13602 VPWR.n1493 VGND 0.0901f
C13603 VPWR.n1495 VGND 0.01496f
C13604 VPWR.n1496 VGND 0.0453f
C13605 VPWR.n1497 VGND 0.11584f
C13606 VPWR.n1498 VGND -0.01553f
C13607 VPWR.n1499 VGND 0.06953f
C13608 VPWR.n1500 VGND 0.06953f
C13609 VPWR.n1501 VGND -0.01553f
C13610 VPWR.n1502 VGND 0.0453f
C13611 VPWR.n1503 VGND 0.11584f
C13612 VPWR.n1504 VGND 0.01496f
C13613 VPWR.n1506 VGND 0.0901f
C13614 VPWR.t17 VGND 0.09955f
C13615 VPWR.t276 VGND 0.06535f
C13616 VPWR.t820 VGND 0.07675f
C13617 VPWR.t124 VGND 0.06535f
C13618 VPWR.t139 VGND 0.09955f
C13619 VPWR.n1507 VGND 0.0901f
C13620 VPWR.n1509 VGND 0.01496f
C13621 VPWR.n1510 VGND 0.0453f
C13622 VPWR.n1511 VGND 0.11584f
C13623 VPWR.n1512 VGND -0.01553f
C13624 VPWR.n1513 VGND 0.06953f
C13625 VPWR.n1514 VGND 0.06953f
C13626 VPWR.n1515 VGND -0.01553f
C13627 VPWR.n1516 VGND 0.0453f
C13628 VPWR.n1517 VGND 0.11584f
C13629 VPWR.n1518 VGND 0.01496f
C13630 VPWR.n1520 VGND 0.0901f
C13631 VPWR.t280 VGND 0.09955f
C13632 VPWR.t154 VGND 0.06535f
C13633 VPWR.t556 VGND 0.07675f
C13634 VPWR.t272 VGND 0.06535f
C13635 VPWR.t296 VGND 0.09955f
C13636 VPWR.n1521 VGND 0.0901f
C13637 VPWR.n1523 VGND 0.01496f
C13638 VPWR.n1524 VGND 0.0453f
C13639 VPWR.n1525 VGND 0.11584f
C13640 VPWR.n1526 VGND -0.01553f
C13641 VPWR.n1527 VGND 0.06953f
C13642 VPWR.n1528 VGND 0.06953f
C13643 VPWR.n1529 VGND 0.06953f
C13644 VPWR.n1530 VGND 0.06953f
C13645 VPWR.n1531 VGND -0.01553f
C13646 VPWR.n1532 VGND 0.11584f
C13647 VPWR.n1533 VGND 0.01496f
C13648 VPWR.n1535 VGND 0.0901f
C13649 VPWR.t1345 VGND 0.07675f
C13650 VPWR.t23 VGND 0.06535f
C13651 VPWR.t39 VGND 0.09955f
C13652 VPWR.n1536 VGND 0.0901f
C13653 VPWR.n1538 VGND 0.01496f
C13654 VPWR.n1539 VGND 0.11584f
C13655 VPWR.n1540 VGND 0.0453f
C13656 VPWR.n1541 VGND 0.05468f
C13657 VPWR.n1542 VGND 0.07639f
C13658 VPWR.t22 VGND 0.01033f
C13659 VPWR.n1543 VGND 0.02305f
C13660 VPWR.n1544 VGND 0.01579f
C13661 VPWR.n1545 VGND 0.05199f
C13662 VPWR.n1546 VGND 0.08114f
C13663 VPWR.n1547 VGND 0.07639f
C13664 VPWR.t271 VGND 0.01033f
C13665 VPWR.n1548 VGND 0.02305f
C13666 VPWR.n1549 VGND 0.01579f
C13667 VPWR.n1550 VGND 0.05199f
C13668 VPWR.n1551 VGND 0.08114f
C13669 VPWR.n1552 VGND 0.07639f
C13670 VPWR.t153 VGND 0.01033f
C13671 VPWR.n1553 VGND 0.02305f
C13672 VPWR.n1554 VGND 0.01579f
C13673 VPWR.n1555 VGND 0.05199f
C13674 VPWR.n1556 VGND 0.08114f
C13675 VPWR.n1557 VGND 0.07639f
C13676 VPWR.t123 VGND 0.01033f
C13677 VPWR.n1558 VGND 0.02305f
C13678 VPWR.n1559 VGND 0.01579f
C13679 VPWR.n1560 VGND 0.05199f
C13680 VPWR.n1561 VGND 0.08114f
C13681 VPWR.n1562 VGND 0.07639f
C13682 VPWR.t275 VGND 0.01033f
C13683 VPWR.n1563 VGND 0.02305f
C13684 VPWR.n1564 VGND 0.01579f
C13685 VPWR.n1565 VGND 0.05199f
C13686 VPWR.n1566 VGND 0.08114f
C13687 VPWR.n1567 VGND 0.07639f
C13688 VPWR.t273 VGND 0.01033f
C13689 VPWR.n1568 VGND 0.02305f
C13690 VPWR.n1569 VGND 0.01579f
C13691 VPWR.n1570 VGND 0.05199f
C13692 VPWR.n1571 VGND 0.08114f
C13693 VPWR.n1572 VGND 0.07639f
C13694 VPWR.t118 VGND 0.01033f
C13695 VPWR.n1573 VGND 0.02305f
C13696 VPWR.n1574 VGND 0.01579f
C13697 VPWR.n1575 VGND 0.05199f
C13698 VPWR.n1576 VGND 0.08114f
C13699 VPWR.n1577 VGND 0.07639f
C13700 VPWR.t14 VGND 0.01033f
C13701 VPWR.n1578 VGND 0.02305f
C13702 VPWR.n1579 VGND 0.01579f
C13703 VPWR.n1580 VGND 0.05199f
C13704 VPWR.n1581 VGND 0.08114f
C13705 VPWR.n1582 VGND 0.07639f
C13706 VPWR.n1583 VGND 0.05468f
C13707 VPWR.n1584 VGND 0.0453f
C13708 VPWR.n1585 VGND 0.11584f
C13709 VPWR.n1586 VGND -0.01553f
C13710 VPWR.n1587 VGND 0.06953f
C13711 VPWR.n1588 VGND 0.06953f
C13712 VPWR.n1589 VGND -0.01553f
C13713 VPWR.n1591 VGND 0.01427f
C13714 VPWR.n1593 VGND 0.0901f
C13715 VPWR.t166 VGND 0.07675f
C13716 VPWR.t47 VGND 0.06535f
C13717 VPWR.t80 VGND 0.09955f
C13718 VPWR.n1594 VGND 0.0901f
C13719 VPWR.n1596 VGND 0.01427f
C13720 VPWR.n1597 VGND 0.02861f
C13721 VPWR.t79 VGND 0.01018f
C13722 VPWR.n1598 VGND 0.02594f
C13723 VPWR.n1599 VGND 0.03075f
C13724 VPWR.t46 VGND 0.01033f
C13725 VPWR.n1601 VGND 0.02304f
C13726 VPWR.n1602 VGND 0.02346f
C13727 VPWR.n1603 VGND 0.01479f
C13728 VPWR.n1605 VGND 0.01517f
C13729 VPWR.n1606 VGND 0.01985f
C13730 VPWR.n1607 VGND 0.19753f
C13731 VPWR.n1608 VGND 0.14641f
C13732 VPWR.n1609 VGND 0.01985f
C13733 VPWR.n1610 VGND 0.01479f
C13734 VPWR.t178 VGND 0.01021f
C13735 VPWR.n1611 VGND 0.02492f
C13736 VPWR.n1612 VGND 0.02734f
C13737 VPWR.n1613 VGND 0.02861f
C13738 VPWR.t346 VGND 0.01018f
C13739 VPWR.n1614 VGND 0.02594f
C13740 VPWR.n1615 VGND 0.03075f
C13741 VPWR.t212 VGND 0.01033f
C13742 VPWR.n1617 VGND 0.02304f
C13743 VPWR.n1618 VGND 0.02346f
C13744 VPWR.n1619 VGND 0.01517f
C13745 VPWR.n1620 VGND 0.01985f
C13746 VPWR.n1621 VGND 0.01479f
C13747 VPWR.t338 VGND 0.01021f
C13748 VPWR.n1622 VGND 0.02492f
C13749 VPWR.n1623 VGND 0.02734f
C13750 VPWR.n1624 VGND 0.02861f
C13751 VPWR.t64 VGND 0.01018f
C13752 VPWR.n1625 VGND 0.02594f
C13753 VPWR.n1626 VGND 0.03075f
C13754 VPWR.t320 VGND 0.01033f
C13755 VPWR.n1628 VGND 0.02304f
C13756 VPWR.n1629 VGND 0.02346f
C13757 VPWR.n1630 VGND 0.01479f
C13758 VPWR.n1632 VGND 0.01517f
C13759 VPWR.n1633 VGND 0.01985f
C13760 VPWR.n1634 VGND 0.14641f
C13761 VPWR.n1635 VGND 0.14641f
C13762 VPWR.n1636 VGND 0.01985f
C13763 VPWR.n1637 VGND 0.01479f
C13764 VPWR.t206 VGND 0.01021f
C13765 VPWR.n1638 VGND 0.02492f
C13766 VPWR.n1639 VGND 0.02734f
C13767 VPWR.n1640 VGND 0.02861f
C13768 VPWR.t235 VGND 0.01018f
C13769 VPWR.n1641 VGND 0.02594f
C13770 VPWR.n1642 VGND 0.03075f
C13771 VPWR.t102 VGND 0.01033f
C13772 VPWR.n1644 VGND 0.02304f
C13773 VPWR.n1645 VGND 0.02346f
C13774 VPWR.n1646 VGND 0.01517f
C13775 VPWR.n1647 VGND 0.01985f
C13776 VPWR.n1648 VGND 0.01479f
C13777 VPWR.t317 VGND 0.01021f
C13778 VPWR.n1649 VGND 0.02492f
C13779 VPWR.n1650 VGND 0.02734f
C13780 VPWR.n1651 VGND 0.02861f
C13781 VPWR.t343 VGND 0.01018f
C13782 VPWR.n1652 VGND 0.02594f
C13783 VPWR.n1653 VGND 0.03075f
C13784 VPWR.t325 VGND 0.01033f
C13785 VPWR.n1655 VGND 0.02304f
C13786 VPWR.n1656 VGND 0.02346f
C13787 VPWR.n1657 VGND 0.01479f
C13788 VPWR.n1659 VGND 0.01517f
C13789 VPWR.n1660 VGND 0.01985f
C13790 VPWR.n1661 VGND 0.14641f
C13791 VPWR.n1662 VGND 0.14641f
C13792 VPWR.n1663 VGND 0.01985f
C13793 VPWR.n1664 VGND 0.01479f
C13794 VPWR.t99 VGND 0.01021f
C13795 VPWR.n1665 VGND 0.02492f
C13796 VPWR.n1666 VGND 0.02734f
C13797 VPWR.n1667 VGND 0.02861f
C13798 VPWR.t130 VGND 0.01018f
C13799 VPWR.n1668 VGND 0.02594f
C13800 VPWR.n1669 VGND 0.03075f
C13801 VPWR.t85 VGND 0.01033f
C13802 VPWR.n1671 VGND 0.02304f
C13803 VPWR.n1672 VGND 0.02346f
C13804 VPWR.n1673 VGND 0.01517f
C13805 VPWR.n1674 VGND 0.01985f
C13806 VPWR.n1675 VGND 0.01479f
C13807 VPWR.t203 VGND 0.01021f
C13808 VPWR.n1676 VGND 0.02492f
C13809 VPWR.n1677 VGND 0.02734f
C13810 VPWR.n1678 VGND 0.02861f
C13811 VPWR.t257 VGND 0.01018f
C13812 VPWR.n1679 VGND 0.02594f
C13813 VPWR.n1680 VGND 0.03075f
C13814 VPWR.t238 VGND 0.01033f
C13815 VPWR.n1682 VGND 0.02304f
C13816 VPWR.n1683 VGND 0.02346f
C13817 VPWR.n1684 VGND 0.01479f
C13818 VPWR.n1686 VGND 0.01517f
C13819 VPWR.n1687 VGND 0.01985f
C13820 VPWR.n1688 VGND 0.14641f
C13821 VPWR.n1689 VGND 0.14641f
C13822 VPWR.n1690 VGND 0.01985f
C13823 VPWR.n1691 VGND 0.01479f
C13824 VPWR.t381 VGND 0.01021f
C13825 VPWR.n1692 VGND 0.02492f
C13826 VPWR.n1693 VGND 0.02734f
C13827 VPWR.n1694 VGND 0.02861f
C13828 VPWR.t24 VGND 0.01018f
C13829 VPWR.n1695 VGND 0.02594f
C13830 VPWR.n1696 VGND 0.03075f
C13831 VPWR.t110 VGND 0.01033f
C13832 VPWR.n1698 VGND 0.02304f
C13833 VPWR.n1699 VGND 0.02346f
C13834 VPWR.n1700 VGND 0.01517f
C13835 VPWR.n1701 VGND 0.01985f
C13836 VPWR.n1702 VGND 0.01479f
C13837 VPWR.t125 VGND 0.01021f
C13838 VPWR.n1703 VGND 0.02492f
C13839 VPWR.n1704 VGND 0.02734f
C13840 VPWR.n1705 VGND 0.02861f
C13841 VPWR.t262 VGND 0.01018f
C13842 VPWR.n1706 VGND 0.02594f
C13843 VPWR.n1707 VGND 0.03075f
C13844 VPWR.t136 VGND 0.01033f
C13845 VPWR.n1709 VGND 0.02304f
C13846 VPWR.n1710 VGND 0.02346f
C13847 VPWR.n1711 VGND 0.01479f
C13848 VPWR.n1713 VGND 0.01517f
C13849 VPWR.n1714 VGND 0.01985f
C13850 VPWR.n1715 VGND 0.14641f
C13851 VPWR.t282 VGND 0.01021f
C13852 VPWR.n1716 VGND 0.02492f
C13853 VPWR.n1717 VGND 0.02734f
C13854 VPWR.t290 VGND 0.01018f
C13855 VPWR.n1718 VGND 0.02594f
C13856 VPWR.n1719 VGND 0.03075f
C13857 VPWR.t161 VGND 0.01033f
C13858 VPWR.n1721 VGND 0.02304f
C13859 VPWR.n1722 VGND 0.02346f
C13860 VPWR.n1723 VGND 0.01479f
C13861 VPWR.n1725 VGND 0.01517f
C13862 VPWR.n1726 VGND 0.01985f
C13863 VPWR.n1727 VGND 0.1762f
C13864 VPWR.n1728 VGND 0.02116f
C13865 VPWR.n1729 VGND 0.01479f
C13866 VPWR.t12 VGND 0.01033f
C13867 VPWR.n1730 VGND 0.02304f
C13868 VPWR.n1731 VGND 0.02346f
C13869 VPWR.t9 VGND 0.01018f
C13870 VPWR.n1733 VGND 0.02594f
C13871 VPWR.n1734 VGND 0.03075f
C13872 VPWR.n1735 VGND 0.02861f
C13873 VPWR.n1737 VGND 0.01427f
C13874 VPWR.n1739 VGND 0.0901f
C13875 VPWR.t283 VGND 0.07675f
C13876 VPWR.t162 VGND 0.06535f
C13877 VPWR.t291 VGND 0.09955f
C13878 VPWR.n1740 VGND 0.0901f
C13879 VPWR.n1742 VGND 0.01427f
C13880 VPWR.n1744 VGND 0.0453f
C13881 VPWR.t32 VGND 0.01018f
C13882 VPWR.n1745 VGND 0.02533f
C13883 VPWR.t34 VGND 0.02231f
C13884 VPWR.n1747 VGND 0.04766f
C13885 VPWR.t686 VGND 0.02465f
C13886 VPWR.n1748 VGND 0.03907f
C13887 VPWR.t304 VGND 0.06535f
C13888 VPWR.t685 VGND 0.07675f
C13889 VPWR.t342 VGND 0.06535f
C13890 VPWR.t83 VGND 0.09955f
C13891 VPWR.n1749 VGND 0.0901f
C13892 VPWR.n1751 VGND 0.01496f
C13893 VPWR.n1752 VGND 0.11584f
C13894 VPWR.n1753 VGND -0.01553f
C13895 VPWR.n1754 VGND 0.06953f
C13896 VPWR.n1755 VGND 0.06953f
C13897 VPWR.n1756 VGND -0.01553f
C13898 VPWR.n1757 VGND 0.11584f
C13899 VPWR.n1758 VGND 0.01496f
C13900 VPWR.n1760 VGND 0.0901f
C13901 VPWR.t1073 VGND 0.07675f
C13902 VPWR.t286 VGND 0.06535f
C13903 VPWR.t210 VGND 0.09955f
C13904 VPWR.n1761 VGND 0.0901f
C13905 VPWR.n1763 VGND 0.01496f
C13906 VPWR.n1764 VGND 0.11584f
C13907 VPWR.n1765 VGND 0.0453f
C13908 VPWR.n1766 VGND 0.05468f
C13909 VPWR.n1767 VGND 0.07639f
C13910 VPWR.t285 VGND 0.01033f
C13911 VPWR.n1768 VGND 0.02305f
C13912 VPWR.n1769 VGND 0.01579f
C13913 VPWR.n1770 VGND 0.05199f
C13914 VPWR.n1771 VGND 0.08114f
C13915 VPWR.n1772 VGND 0.07639f
C13916 VPWR.t303 VGND 0.01033f
C13917 VPWR.n1773 VGND 0.02305f
C13918 VPWR.n1774 VGND 0.01579f
C13919 VPWR.n1775 VGND 0.05199f
C13920 VPWR.n1776 VGND 0.08114f
C13921 VPWR.t173 VGND 0.01033f
C13922 VPWR.n1777 VGND 0.02305f
C13923 VPWR.n1778 VGND 0.01579f
C13924 VPWR.n1779 VGND 0.05197f
C13925 VPWR.n1780 VGND 0.04278f
C13926 VPWR.t341 VGND 0.01033f
C13927 VPWR.n1781 VGND 0.02305f
C13928 VPWR.n1782 VGND 0.01579f
C13929 VPWR.n1783 VGND 0.05199f
C13930 VPWR.n1784 VGND 0.08114f
C13931 VPWR.n1785 VGND 0.07639f
C13932 VPWR.n1786 VGND 0.05468f
C13933 VPWR.n1787 VGND 0.0453f
C13934 VPWR.n1788 VGND 0.11584f
C13935 VPWR.n1789 VGND 0.01496f
C13936 VPWR.n1791 VGND 0.0901f
C13937 VPWR.t191 VGND 0.09955f
C13938 VPWR.t174 VGND 0.06535f
C13939 VPWR.t299 VGND 0.11101f
C13940 VPWR.n1792 VGND 0.06343f
C13941 VPWR.n1793 VGND 0.01496f
C13942 VPWR.n1794 VGND 0.11584f
C13943 VPWR.n1795 VGND 0.13705f
C13944 VPWR.n1796 VGND 0.84572f
C13945 VPWR.n1797 VGND 0.06953f
C13946 VPWR.n1798 VGND 0.06953f
C13947 VPWR.n1799 VGND 0.06953f
C13948 VPWR.n1800 VGND 0.06953f
C13949 VPWR.n1801 VGND 0.06953f
C13950 VPWR.n1802 VGND 0.06953f
C13951 VPWR.n1803 VGND 0.06953f
C13952 VPWR.n1804 VGND 0.06953f
C13953 VPWR.n1805 VGND 0.06953f
C13954 VPWR.n1806 VGND 0.06953f
C13955 VPWR.n1807 VGND 0.06953f
C13956 VPWR.n1808 VGND 0.06953f
C13957 VPWR.n1809 VGND 0.06953f
C13958 VPWR.n1810 VGND 0.06953f
C13959 VPWR.n1811 VGND 0.06953f
C13960 VPWR.n1812 VGND 0.16128f
C13961 VPWR.n1813 VGND 0.84572f
C13962 VPWR.n1814 VGND 0.84572f
C13963 VPWR.n1815 VGND 0.16128f
C13964 VPWR.n1816 VGND 0.11584f
C13965 VPWR.n1817 VGND 0.01496f
C13966 VPWR.n1818 VGND 0.06343f
C13967 VPWR.t336 VGND 0.11101f
C13968 VPWR.t1856 VGND 0.06535f
C13969 VPWR.t602 VGND 0.09955f
C13970 VPWR.n1819 VGND 0.0901f
C13971 VPWR.n1821 VGND 0.01496f
C13972 VPWR.n1822 VGND 0.11584f
C13973 VPWR.n1823 VGND 0.06953f
C13974 VPWR.n1824 VGND 0.06953f
C13975 VPWR.n1825 VGND 0.11584f
C13976 VPWR.n1826 VGND 0.01496f
C13977 VPWR.n1828 VGND 0.0901f
C13978 VPWR.t757 VGND 0.07675f
C13979 VPWR.t903 VGND 0.06535f
C13980 VPWR.t1713 VGND 0.09955f
C13981 VPWR.n1829 VGND 0.0901f
C13982 VPWR.n1831 VGND 0.01496f
C13983 VPWR.n1832 VGND 0.11584f
C13984 VPWR.n1833 VGND 0.06953f
C13985 VPWR.n1834 VGND 0.06953f
C13986 VPWR.n1835 VGND 0.11584f
C13987 VPWR.n1836 VGND 0.01496f
C13988 VPWR.n1838 VGND 0.0901f
C13989 VPWR.t1256 VGND 0.07675f
C13990 VPWR.t540 VGND 0.06535f
C13991 VPWR.t1316 VGND 0.09955f
C13992 VPWR.n1839 VGND 0.0901f
C13993 VPWR.n1841 VGND 0.01496f
C13994 VPWR.n1842 VGND 0.11584f
C13995 VPWR.n1843 VGND 0.06953f
C13996 VPWR.n1844 VGND 0.06953f
C13997 VPWR.n1845 VGND 0.11584f
C13998 VPWR.n1846 VGND 0.01496f
C13999 VPWR.n1848 VGND 0.0901f
C14000 VPWR.t1242 VGND 0.07675f
C14001 VPWR.t1854 VGND 0.06535f
C14002 VPWR.t941 VGND 0.09955f
C14003 VPWR.n1849 VGND 0.0901f
C14004 VPWR.n1851 VGND 0.01496f
C14005 VPWR.n1852 VGND 0.11584f
C14006 VPWR.n1853 VGND 0.06953f
C14007 VPWR.n1854 VGND 0.06953f
C14008 VPWR.n1855 VGND 0.11584f
C14009 VPWR.n1856 VGND 0.01496f
C14010 VPWR.n1858 VGND 0.0901f
C14011 VPWR.t888 VGND 0.07675f
C14012 VPWR.t1858 VGND 0.06535f
C14013 VPWR.t806 VGND 0.09955f
C14014 VPWR.n1859 VGND 0.0901f
C14015 VPWR.n1861 VGND 0.01496f
C14016 VPWR.n1862 VGND 0.11584f
C14017 VPWR.n1863 VGND 0.06953f
C14018 VPWR.n1864 VGND 0.06953f
C14019 VPWR.n1865 VGND 0.11584f
C14020 VPWR.n1866 VGND 0.01496f
C14021 VPWR.n1868 VGND 0.0901f
C14022 VPWR.t1136 VGND 0.07675f
C14023 VPWR.t906 VGND 0.06535f
C14024 VPWR.t1541 VGND 0.09955f
C14025 VPWR.n1869 VGND 0.0901f
C14026 VPWR.n1871 VGND 0.01496f
C14027 VPWR.n1872 VGND 0.11584f
C14028 VPWR.n1873 VGND 0.06953f
C14029 VPWR.n1874 VGND 0.06953f
C14030 VPWR.n1875 VGND 0.11584f
C14031 VPWR.n1876 VGND 0.01496f
C14032 VPWR.n1878 VGND 0.0901f
C14033 VPWR.t1272 VGND 0.07675f
C14034 VPWR.t542 VGND 0.06535f
C14035 VPWR.t1462 VGND 0.09955f
C14036 VPWR.n1879 VGND 0.0901f
C14037 VPWR.n1881 VGND 0.01496f
C14038 VPWR.n1882 VGND 0.11584f
C14039 VPWR.n1883 VGND 0.06953f
C14040 VPWR.n1884 VGND 0.06953f
C14041 VPWR.n1885 VGND 0.11584f
C14042 VPWR.n1886 VGND 0.01496f
C14043 VPWR.n1888 VGND 0.0901f
C14044 VPWR.t475 VGND 0.07675f
C14045 VPWR.t1855 VGND 0.06535f
C14046 VPWR.t1016 VGND 0.09955f
C14047 VPWR.n1889 VGND 0.0901f
C14048 VPWR.n1891 VGND 0.01496f
C14049 VPWR.n1892 VGND 0.11584f
C14050 VPWR.n1893 VGND 0.06953f
C14051 VPWR.n1894 VGND 0.84042f
C14052 VPWR.n1895 VGND 0.16128f
C14053 VPWR.n1896 VGND 0.06953f
C14054 VPWR.n1897 VGND 0.06953f
C14055 VPWR.n1898 VGND 0.06953f
C14056 VPWR.n1899 VGND 0.06953f
C14057 VPWR.n1900 VGND 0.06953f
C14058 VPWR.n1901 VGND 0.06953f
C14059 VPWR.n1902 VGND 0.06953f
C14060 VPWR.n1903 VGND 0.06953f
C14061 VPWR.n1904 VGND 0.06953f
C14062 VPWR.n1905 VGND 0.06953f
C14063 VPWR.n1906 VGND 0.06953f
C14064 VPWR.n1907 VGND 0.06953f
C14065 VPWR.n1908 VGND 0.06953f
C14066 VPWR.n1909 VGND 0.06953f
C14067 VPWR.n1910 VGND 0.06953f
C14068 VPWR.n1911 VGND 0.84042f
C14069 VPWR.n1912 VGND 0.84042f
C14070 VPWR.n1913 VGND 0.06953f
C14071 VPWR.n1914 VGND 0.11584f
C14072 VPWR.n1915 VGND 0.01496f
C14073 VPWR.n1917 VGND 0.0901f
C14074 VPWR.t826 VGND 0.09955f
C14075 VPWR.t1824 VGND 0.06535f
C14076 VPWR.t1559 VGND 0.07675f
C14077 VPWR.t717 VGND 0.06535f
C14078 VPWR.t1553 VGND 0.09955f
C14079 VPWR.n1918 VGND 0.0901f
C14080 VPWR.n1920 VGND 0.01496f
C14081 VPWR.n1921 VGND 0.11584f
C14082 VPWR.n1922 VGND 0.06953f
C14083 VPWR.n1923 VGND 0.06953f
C14084 VPWR.n1924 VGND 0.11584f
C14085 VPWR.n1925 VGND 0.01496f
C14086 VPWR.n1927 VGND 0.0901f
C14087 VPWR.t1480 VGND 0.09955f
C14088 VPWR.t716 VGND 0.06535f
C14089 VPWR.t1516 VGND 0.07675f
C14090 VPWR.t712 VGND 0.06535f
C14091 VPWR.t1390 VGND 0.09955f
C14092 VPWR.n1928 VGND 0.0901f
C14093 VPWR.n1930 VGND 0.01496f
C14094 VPWR.n1931 VGND 0.11584f
C14095 VPWR.n1932 VGND 0.06953f
C14096 VPWR.n1933 VGND 0.06953f
C14097 VPWR.n1934 VGND 0.11584f
C14098 VPWR.n1935 VGND 0.01496f
C14099 VPWR.n1937 VGND 0.0901f
C14100 VPWR.t1331 VGND 0.09955f
C14101 VPWR.t1530 VGND 0.06535f
C14102 VPWR.t628 VGND 0.07675f
C14103 VPWR.t1529 VGND 0.06535f
C14104 VPWR.t622 VGND 0.09955f
C14105 VPWR.n1938 VGND 0.0901f
C14106 VPWR.n1940 VGND 0.01496f
C14107 VPWR.n1941 VGND 0.11584f
C14108 VPWR.n1942 VGND 0.06953f
C14109 VPWR.n1943 VGND 0.06953f
C14110 VPWR.n1944 VGND 0.11584f
C14111 VPWR.n1945 VGND 0.01496f
C14112 VPWR.n1947 VGND 0.0901f
C14113 VPWR.t790 VGND 0.09955f
C14114 VPWR.t1827 VGND 0.06535f
C14115 VPWR.t938 VGND 0.07675f
C14116 VPWR.t1826 VGND 0.06535f
C14117 VPWR.t873 VGND 0.09955f
C14118 VPWR.n1948 VGND 0.0901f
C14119 VPWR.n1950 VGND 0.01496f
C14120 VPWR.n1951 VGND 0.11584f
C14121 VPWR.n1952 VGND 0.06953f
C14122 VPWR.n1953 VGND 0.06953f
C14123 VPWR.n1954 VGND 0.11584f
C14124 VPWR.n1955 VGND 0.01496f
C14125 VPWR.n1957 VGND 0.0901f
C14126 VPWR.t546 VGND 0.09955f
C14127 VPWR.t1531 VGND 0.06535f
C14128 VPWR.t514 VGND 0.07675f
C14129 VPWR.t715 VGND 0.06535f
C14130 VPWR.t508 VGND 0.09955f
C14131 VPWR.n1958 VGND 0.0901f
C14132 VPWR.n1960 VGND 0.01496f
C14133 VPWR.n1961 VGND 0.11584f
C14134 VPWR.n1962 VGND 0.06953f
C14135 VPWR.n1963 VGND 0.06953f
C14136 VPWR.n1964 VGND 0.11584f
C14137 VPWR.n1965 VGND 0.01496f
C14138 VPWR.n1967 VGND 0.0901f
C14139 VPWR.t1666 VGND 0.09955f
C14140 VPWR.t714 VGND 0.06535f
C14141 VPWR.t1354 VGND 0.07675f
C14142 VPWR.t1528 VGND 0.06535f
C14143 VPWR.t1284 VGND 0.09955f
C14144 VPWR.n1968 VGND 0.0901f
C14145 VPWR.n1970 VGND 0.01496f
C14146 VPWR.n1971 VGND 0.11584f
C14147 VPWR.n1972 VGND 0.06953f
C14148 VPWR.n1973 VGND 0.06953f
C14149 VPWR.n1974 VGND 0.11584f
C14150 VPWR.n1975 VGND 0.01496f
C14151 VPWR.n1977 VGND 0.0901f
C14152 VPWR.t1298 VGND 0.09955f
C14153 VPWR.t1527 VGND 0.06535f
C14154 VPWR.t1370 VGND 0.07675f
C14155 VPWR.t718 VGND 0.06535f
C14156 VPWR.t1498 VGND 0.09955f
C14157 VPWR.n1978 VGND 0.0901f
C14158 VPWR.n1980 VGND 0.01496f
C14159 VPWR.n1981 VGND 0.11584f
C14160 VPWR.n1982 VGND 0.06953f
C14161 VPWR.n1983 VGND 0.06953f
C14162 VPWR.n1984 VGND 0.11584f
C14163 VPWR.n1985 VGND 0.01496f
C14164 VPWR.n1987 VGND 0.0901f
C14165 VPWR.t524 VGND 0.09955f
C14166 VPWR.t1825 VGND 0.06535f
C14167 VPWR.t44 VGND 0.11101f
C14168 VPWR.n1988 VGND 0.06343f
C14169 VPWR.n1989 VGND 0.01496f
C14170 VPWR.n1990 VGND 0.11584f
C14171 VPWR.n1991 VGND 0.16128f
C14172 VPWR.n1992 VGND 0.84572f
C14173 VPWR.n1993 VGND 0.06953f
C14174 VPWR.n1994 VGND 0.06953f
C14175 VPWR.n1995 VGND 0.06953f
C14176 VPWR.n1996 VGND 0.06953f
C14177 VPWR.n1997 VGND 0.06953f
C14178 VPWR.n1998 VGND 0.06953f
C14179 VPWR.n1999 VGND 0.06953f
C14180 VPWR.n2000 VGND 0.06953f
C14181 VPWR.n2001 VGND 0.06953f
C14182 VPWR.n2002 VGND 0.06953f
C14183 VPWR.n2003 VGND 0.06953f
C14184 VPWR.n2004 VGND 0.06953f
C14185 VPWR.n2005 VGND 0.06953f
C14186 VPWR.n2006 VGND 0.06953f
C14187 VPWR.n2007 VGND 0.06953f
C14188 VPWR.n2008 VGND 0.16128f
C14189 VPWR.n2009 VGND 0.84572f
C14190 VPWR.n2010 VGND 0.84572f
C14191 VPWR.n2011 VGND 0.16128f
C14192 VPWR.n2012 VGND 0.11584f
C14193 VPWR.n2013 VGND 0.01496f
C14194 VPWR.n2014 VGND 0.06343f
C14195 VPWR.t116 VGND 0.11101f
C14196 VPWR.t465 VGND 0.06535f
C14197 VPWR.t1848 VGND 0.09955f
C14198 VPWR.n2015 VGND 0.0901f
C14199 VPWR.n2017 VGND 0.01496f
C14200 VPWR.n2018 VGND 0.11584f
C14201 VPWR.n2019 VGND 0.06953f
C14202 VPWR.n2020 VGND 0.06953f
C14203 VPWR.n2021 VGND 0.11584f
C14204 VPWR.n2022 VGND 0.01496f
C14205 VPWR.n2024 VGND 0.0901f
C14206 VPWR.t1881 VGND 0.07675f
C14207 VPWR.t1599 VGND 0.06535f
C14208 VPWR.t1079 VGND 0.09955f
C14209 VPWR.n2025 VGND 0.0901f
C14210 VPWR.n2027 VGND 0.01496f
C14211 VPWR.n2028 VGND 0.11584f
C14212 VPWR.n2029 VGND 0.06953f
C14213 VPWR.n2030 VGND 0.06953f
C14214 VPWR.n2031 VGND 0.11584f
C14215 VPWR.n2032 VGND 0.01496f
C14216 VPWR.n2034 VGND 0.0901f
C14217 VPWR.t1532 VGND 0.07675f
C14218 VPWR.t1630 VGND 0.06535f
C14219 VPWR.t878 VGND 0.09955f
C14220 VPWR.n2035 VGND 0.0901f
C14221 VPWR.n2037 VGND 0.01496f
C14222 VPWR.n2038 VGND 0.11584f
C14223 VPWR.n2039 VGND 0.06953f
C14224 VPWR.n2040 VGND 0.06953f
C14225 VPWR.n2041 VGND 0.11584f
C14226 VPWR.n2042 VGND 0.01496f
C14227 VPWR.n2044 VGND 0.0901f
C14228 VPWR.t755 VGND 0.07675f
C14229 VPWR.t1603 VGND 0.06535f
C14230 VPWR.t1034 VGND 0.09955f
C14231 VPWR.n2045 VGND 0.0901f
C14232 VPWR.n2047 VGND 0.01496f
C14233 VPWR.n2048 VGND 0.11584f
C14234 VPWR.n2049 VGND 0.06953f
C14235 VPWR.n2050 VGND 0.06953f
C14236 VPWR.n2051 VGND 0.11584f
C14237 VPWR.n2052 VGND 0.01496f
C14238 VPWR.n2054 VGND 0.0901f
C14239 VPWR.t833 VGND 0.07675f
C14240 VPWR.t467 VGND 0.06535f
C14241 VPWR.t1585 VGND 0.09955f
C14242 VPWR.n2055 VGND 0.0901f
C14243 VPWR.n2057 VGND 0.01496f
C14244 VPWR.n2058 VGND 0.11584f
C14245 VPWR.n2059 VGND 0.06953f
C14246 VPWR.n2060 VGND 0.06953f
C14247 VPWR.n2061 VGND 0.11584f
C14248 VPWR.n2062 VGND 0.01496f
C14249 VPWR.n2064 VGND 0.0901f
C14250 VPWR.t656 VGND 0.07675f
C14251 VPWR.t1602 VGND 0.06535f
C14252 VPWR.t1625 VGND 0.09955f
C14253 VPWR.n2065 VGND 0.0901f
C14254 VPWR.n2067 VGND 0.01496f
C14255 VPWR.n2068 VGND 0.11584f
C14256 VPWR.n2069 VGND 0.06953f
C14257 VPWR.n2070 VGND 0.06953f
C14258 VPWR.n2071 VGND 0.11584f
C14259 VPWR.n2072 VGND 0.01496f
C14260 VPWR.n2074 VGND 0.0901f
C14261 VPWR.t388 VGND 0.07675f
C14262 VPWR.t1632 VGND 0.06535f
C14263 VPWR.t1488 VGND 0.09955f
C14264 VPWR.n2075 VGND 0.0901f
C14265 VPWR.n2077 VGND 0.01496f
C14266 VPWR.n2078 VGND 0.11584f
C14267 VPWR.n2079 VGND 0.06953f
C14268 VPWR.n2080 VGND 0.06953f
C14269 VPWR.n2081 VGND 0.11584f
C14270 VPWR.n2082 VGND 0.01496f
C14271 VPWR.n2084 VGND 0.0901f
C14272 VPWR.t1030 VGND 0.07675f
C14273 VPWR.t1604 VGND 0.06535f
C14274 VPWR.t1012 VGND 0.09955f
C14275 VPWR.n2085 VGND 0.0901f
C14276 VPWR.n2087 VGND 0.01496f
C14277 VPWR.n2088 VGND 0.11584f
C14278 VPWR.n2089 VGND 0.06953f
C14279 VPWR.n2090 VGND 0.84042f
C14280 VPWR.n2091 VGND 0.16128f
C14281 VPWR.n2092 VGND 0.06953f
C14282 VPWR.n2093 VGND 0.06953f
C14283 VPWR.n2094 VGND 0.06953f
C14284 VPWR.n2095 VGND 0.06953f
C14285 VPWR.n2096 VGND 0.06953f
C14286 VPWR.n2097 VGND 0.06953f
C14287 VPWR.n2098 VGND 0.06953f
C14288 VPWR.n2099 VGND 0.06953f
C14289 VPWR.n2100 VGND 0.06953f
C14290 VPWR.n2101 VGND 0.06953f
C14291 VPWR.n2102 VGND 0.06953f
C14292 VPWR.n2103 VGND 0.06953f
C14293 VPWR.n2104 VGND 0.06953f
C14294 VPWR.n2105 VGND 0.06953f
C14295 VPWR.n2106 VGND 0.06953f
C14296 VPWR.n2107 VGND 0.84042f
C14297 VPWR.n2108 VGND 0.84042f
C14298 VPWR.n2109 VGND 0.06953f
C14299 VPWR.n2110 VGND 0.11584f
C14300 VPWR.n2111 VGND 0.01496f
C14301 VPWR.n2113 VGND 0.0901f
C14302 VPWR.t824 VGND 0.09955f
C14303 VPWR.t982 VGND 0.06535f
C14304 VPWR.t1557 VGND 0.07675f
C14305 VPWR.t1158 VGND 0.06535f
C14306 VPWR.t1551 VGND 0.09955f
C14307 VPWR.n2114 VGND 0.0901f
C14308 VPWR.n2116 VGND 0.01496f
C14309 VPWR.n2117 VGND 0.11584f
C14310 VPWR.n2118 VGND 0.06953f
C14311 VPWR.n2119 VGND 0.06953f
C14312 VPWR.n2120 VGND 0.11584f
C14313 VPWR.n2121 VGND 0.01496f
C14314 VPWR.n2123 VGND 0.0901f
C14315 VPWR.t1482 VGND 0.09955f
C14316 VPWR.t1157 VGND 0.06535f
C14317 VPWR.t398 VGND 0.07675f
C14318 VPWR.t877 VGND 0.06535f
C14319 VPWR.t998 VGND 0.09955f
C14320 VPWR.n2124 VGND 0.0901f
C14321 VPWR.n2126 VGND 0.01496f
C14322 VPWR.n2127 VGND 0.11584f
C14323 VPWR.n2128 VGND 0.06953f
C14324 VPWR.n2129 VGND 0.06953f
C14325 VPWR.n2130 VGND 0.11584f
C14326 VPWR.n2131 VGND 0.01496f
C14327 VPWR.n2133 VGND 0.0901f
C14328 VPWR.t1329 VGND 0.09955f
C14329 VPWR.t1691 VGND 0.06535f
C14330 VPWR.t626 VGND 0.07675f
C14331 VPWR.t1690 VGND 0.06535f
C14332 VPWR.t620 VGND 0.09955f
C14333 VPWR.n2134 VGND 0.0901f
C14334 VPWR.n2136 VGND 0.01496f
C14335 VPWR.n2137 VGND 0.11584f
C14336 VPWR.n2138 VGND 0.06953f
C14337 VPWR.n2139 VGND 0.06953f
C14338 VPWR.n2140 VGND 0.11584f
C14339 VPWR.n2141 VGND 0.01496f
C14340 VPWR.n2143 VGND 0.0901f
C14341 VPWR.t1589 VGND 0.09955f
C14342 VPWR.t876 VGND 0.06535f
C14343 VPWR.t936 VGND 0.07675f
C14344 VPWR.t875 VGND 0.06535f
C14345 VPWR.t871 VGND 0.09955f
C14346 VPWR.n2144 VGND 0.0901f
C14347 VPWR.n2146 VGND 0.01496f
C14348 VPWR.n2147 VGND 0.11584f
C14349 VPWR.n2148 VGND 0.06953f
C14350 VPWR.n2149 VGND 0.06953f
C14351 VPWR.n2150 VGND 0.11584f
C14352 VPWR.n2151 VGND 0.01496f
C14353 VPWR.n2153 VGND 0.0901f
C14354 VPWR.t544 VGND 0.09955f
C14355 VPWR.t1692 VGND 0.06535f
C14356 VPWR.t512 VGND 0.07675f
C14357 VPWR.t1063 VGND 0.06535f
C14358 VPWR.t506 VGND 0.09955f
C14359 VPWR.n2154 VGND 0.0901f
C14360 VPWR.n2156 VGND 0.01496f
C14361 VPWR.n2157 VGND 0.11584f
C14362 VPWR.n2158 VGND 0.06953f
C14363 VPWR.n2159 VGND 0.06953f
C14364 VPWR.n2160 VGND 0.11584f
C14365 VPWR.n2161 VGND 0.01496f
C14366 VPWR.n2163 VGND 0.0901f
C14367 VPWR.t1664 VGND 0.09955f
C14368 VPWR.t1062 VGND 0.06535f
C14369 VPWR.t1352 VGND 0.07675f
C14370 VPWR.t1689 VGND 0.06535f
C14371 VPWR.t1282 VGND 0.09955f
C14372 VPWR.n2164 VGND 0.0901f
C14373 VPWR.n2166 VGND 0.01496f
C14374 VPWR.n2167 VGND 0.11584f
C14375 VPWR.n2168 VGND 0.06953f
C14376 VPWR.n2169 VGND 0.06953f
C14377 VPWR.n2170 VGND 0.11584f
C14378 VPWR.n2171 VGND 0.01496f
C14379 VPWR.n2173 VGND 0.0901f
C14380 VPWR.t1296 VGND 0.09955f
C14381 VPWR.t1688 VGND 0.06535f
C14382 VPWR.t1502 VGND 0.07675f
C14383 VPWR.t1159 VGND 0.06535f
C14384 VPWR.t1496 VGND 0.09955f
C14385 VPWR.n2174 VGND 0.0901f
C14386 VPWR.n2176 VGND 0.01496f
C14387 VPWR.n2177 VGND 0.11584f
C14388 VPWR.n2178 VGND 0.06953f
C14389 VPWR.n2179 VGND 0.06953f
C14390 VPWR.n2180 VGND 0.11584f
C14391 VPWR.n2181 VGND 0.01496f
C14392 VPWR.n2183 VGND 0.0901f
C14393 VPWR.t522 VGND 0.09955f
C14394 VPWR.t983 VGND 0.06535f
C14395 VPWR.t49 VGND 0.11101f
C14396 VPWR.n2184 VGND 0.06343f
C14397 VPWR.n2185 VGND 0.01496f
C14398 VPWR.n2186 VGND 0.11584f
C14399 VPWR.n2187 VGND 0.16128f
C14400 VPWR.n2188 VGND 0.84572f
C14401 VPWR.n2189 VGND 0.06953f
C14402 VPWR.n2190 VGND 0.06953f
C14403 VPWR.n2191 VGND 0.06953f
C14404 VPWR.n2192 VGND 0.06953f
C14405 VPWR.n2193 VGND 0.06953f
C14406 VPWR.n2194 VGND 0.06953f
C14407 VPWR.n2195 VGND 0.06953f
C14408 VPWR.n2196 VGND 0.06953f
C14409 VPWR.n2197 VGND 0.06953f
C14410 VPWR.n2198 VGND 0.06953f
C14411 VPWR.n2199 VGND 0.06953f
C14412 VPWR.n2200 VGND 0.06953f
C14413 VPWR.n2201 VGND 0.06953f
C14414 VPWR.n2202 VGND 0.06953f
C14415 VPWR.n2203 VGND 0.06953f
C14416 VPWR.n2204 VGND 0.16128f
C14417 VPWR.n2205 VGND 0.84572f
C14418 VPWR.n2206 VGND 0.84572f
C14419 VPWR.n2207 VGND 0.16128f
C14420 VPWR.n2208 VGND 0.11584f
C14421 VPWR.n2209 VGND 0.01496f
C14422 VPWR.n2210 VGND 0.06343f
C14423 VPWR.t215 VGND 0.11101f
C14424 VPWR.t1054 VGND 0.06535f
C14425 VPWR.t780 VGND 0.09955f
C14426 VPWR.n2211 VGND 0.0901f
C14427 VPWR.n2213 VGND 0.01496f
C14428 VPWR.n2214 VGND 0.11584f
C14429 VPWR.n2215 VGND 0.06953f
C14430 VPWR.n2216 VGND 0.06953f
C14431 VPWR.n2217 VGND 0.11584f
C14432 VPWR.n2218 VGND 0.01496f
C14433 VPWR.n2220 VGND 0.0901f
C14434 VPWR.t408 VGND 0.07675f
C14435 VPWR.t1646 VGND 0.06535f
C14436 VPWR.t1916 VGND 0.09955f
C14437 VPWR.n2221 VGND 0.0901f
C14438 VPWR.n2223 VGND 0.01496f
C14439 VPWR.n2224 VGND 0.11584f
C14440 VPWR.n2225 VGND 0.06953f
C14441 VPWR.n2226 VGND 0.06953f
C14442 VPWR.n2227 VGND 0.11584f
C14443 VPWR.n2228 VGND 0.01496f
C14444 VPWR.n2230 VGND 0.0901f
C14445 VPWR.t1836 VGND 0.07675f
C14446 VPWR.t1641 VGND 0.06535f
C14447 VPWR.t1174 VGND 0.09955f
C14448 VPWR.n2231 VGND 0.0901f
C14449 VPWR.n2233 VGND 0.01496f
C14450 VPWR.n2234 VGND 0.11584f
C14451 VPWR.n2235 VGND 0.06953f
C14452 VPWR.n2236 VGND 0.06953f
C14453 VPWR.n2237 VGND 0.11584f
C14454 VPWR.n2238 VGND 0.01496f
C14455 VPWR.n2240 VGND 0.0901f
C14456 VPWR.t731 VGND 0.07675f
C14457 VPWR.t1052 VGND 0.06535f
C14458 VPWR.t884 VGND 0.09955f
C14459 VPWR.n2241 VGND 0.0901f
C14460 VPWR.n2243 VGND 0.01496f
C14461 VPWR.n2244 VGND 0.11584f
C14462 VPWR.n2245 VGND 0.06953f
C14463 VPWR.n2246 VGND 0.06953f
C14464 VPWR.n2247 VGND 0.11584f
C14465 VPWR.n2248 VGND 0.01496f
C14466 VPWR.n2250 VGND 0.0901f
C14467 VPWR.t867 VGND 0.07675f
C14468 VPWR.t1056 VGND 0.06535f
C14469 VPWR.t482 VGND 0.09955f
C14470 VPWR.n2251 VGND 0.0901f
C14471 VPWR.n2253 VGND 0.01496f
C14472 VPWR.n2254 VGND 0.11584f
C14473 VPWR.n2255 VGND 0.06953f
C14474 VPWR.n2256 VGND 0.06953f
C14475 VPWR.n2257 VGND 0.11584f
C14476 VPWR.n2258 VGND 0.01496f
C14477 VPWR.n2260 VGND 0.0901f
C14478 VPWR.t953 VGND 0.07675f
C14479 VPWR.t1051 VGND 0.06535f
C14480 VPWR.t1695 VGND 0.09955f
C14481 VPWR.n2261 VGND 0.0901f
C14482 VPWR.n2263 VGND 0.01496f
C14483 VPWR.n2264 VGND 0.11584f
C14484 VPWR.n2265 VGND 0.06953f
C14485 VPWR.n2266 VGND 0.06953f
C14486 VPWR.n2267 VGND 0.11584f
C14487 VPWR.n2268 VGND 0.01496f
C14488 VPWR.n2270 VGND 0.0901f
C14489 VPWR.t994 VGND 0.07675f
C14490 VPWR.t1643 VGND 0.06535f
C14491 VPWR.t1446 VGND 0.09955f
C14492 VPWR.n2271 VGND 0.0901f
C14493 VPWR.n2273 VGND 0.01496f
C14494 VPWR.n2274 VGND 0.11584f
C14495 VPWR.n2275 VGND 0.06953f
C14496 VPWR.n2276 VGND 0.06953f
C14497 VPWR.n2277 VGND 0.11584f
C14498 VPWR.n2278 VGND 0.01496f
C14499 VPWR.n2280 VGND 0.0901f
C14500 VPWR.t1902 VGND 0.07675f
C14501 VPWR.t1053 VGND 0.06535f
C14502 VPWR.t852 VGND 0.09955f
C14503 VPWR.n2281 VGND 0.0901f
C14504 VPWR.n2283 VGND 0.01496f
C14505 VPWR.n2284 VGND 0.11584f
C14506 VPWR.n2285 VGND 0.06953f
C14507 VPWR.n2286 VGND 0.84042f
C14508 VPWR.n2287 VGND 0.16128f
C14509 VPWR.n2288 VGND 0.06953f
C14510 VPWR.n2289 VGND 0.06953f
C14511 VPWR.n2290 VGND 0.06953f
C14512 VPWR.n2291 VGND 0.06953f
C14513 VPWR.n2292 VGND 0.06953f
C14514 VPWR.n2293 VGND 0.06953f
C14515 VPWR.n2294 VGND 0.06953f
C14516 VPWR.n2295 VGND 0.06953f
C14517 VPWR.n2296 VGND 0.06953f
C14518 VPWR.n2297 VGND 0.06953f
C14519 VPWR.n2298 VGND 0.06953f
C14520 VPWR.n2299 VGND 0.06953f
C14521 VPWR.n2300 VGND 0.06953f
C14522 VPWR.n2301 VGND 0.06953f
C14523 VPWR.n2302 VGND 0.06953f
C14524 VPWR.n2303 VGND 0.84042f
C14525 VPWR.n2304 VGND 0.84042f
C14526 VPWR.n2305 VGND 0.06953f
C14527 VPWR.n2306 VGND 0.11584f
C14528 VPWR.n2307 VGND 0.01496f
C14529 VPWR.n2309 VGND 0.0901f
C14530 VPWR.t1191 VGND 0.09955f
C14531 VPWR.t1731 VGND 0.06535f
C14532 VPWR.t1026 VGND 0.07675f
C14533 VPWR.t1327 VGND 0.06535f
C14534 VPWR.t689 VGND 0.09955f
C14535 VPWR.n2310 VGND 0.0901f
C14536 VPWR.n2312 VGND 0.01496f
C14537 VPWR.n2313 VGND 0.11584f
C14538 VPWR.n2314 VGND 0.06953f
C14539 VPWR.n2315 VGND 0.06953f
C14540 VPWR.n2316 VGND 0.11584f
C14541 VPWR.n2317 VGND 0.01496f
C14542 VPWR.n2319 VGND 0.0901f
C14543 VPWR.t1492 VGND 0.09955f
C14544 VPWR.t1326 VGND 0.06535f
C14545 VPWR.t1396 VGND 0.07675f
C14546 VPWR.t768 VGND 0.06535f
C14547 VPWR.t1508 VGND 0.09955f
C14548 VPWR.n2320 VGND 0.0901f
C14549 VPWR.n2322 VGND 0.01496f
C14550 VPWR.n2323 VGND 0.11584f
C14551 VPWR.n2324 VGND 0.06953f
C14552 VPWR.n2325 VGND 0.06953f
C14553 VPWR.n2326 VGND 0.11584f
C14554 VPWR.n2327 VGND 0.01496f
C14555 VPWR.n2329 VGND 0.0901f
C14556 VPWR.t1595 VGND 0.09955f
C14557 VPWR.t1163 VGND 0.06535f
C14558 VPWR.t652 VGND 0.07675f
C14559 VPWR.t1162 VGND 0.06535f
C14560 VPWR.t959 VGND 0.09955f
C14561 VPWR.n2330 VGND 0.0901f
C14562 VPWR.n2332 VGND 0.01496f
C14563 VPWR.n2333 VGND 0.11584f
C14564 VPWR.n2334 VGND 0.06953f
C14565 VPWR.n2335 VGND 0.06953f
C14566 VPWR.n2336 VGND 0.11584f
C14567 VPWR.n2337 VGND 0.01496f
C14568 VPWR.n2339 VGND 0.0901f
C14569 VPWR.t1579 VGND 0.09955f
C14570 VPWR.t767 VGND 0.06535f
C14571 VPWR.t662 VGND 0.07675f
C14572 VPWR.t1733 VGND 0.06535f
C14573 VPWR.t900 VGND 0.09955f
C14574 VPWR.n2340 VGND 0.0901f
C14575 VPWR.n2342 VGND 0.01496f
C14576 VPWR.n2343 VGND 0.11584f
C14577 VPWR.n2344 VGND 0.06953f
C14578 VPWR.n2345 VGND 0.06953f
C14579 VPWR.n2346 VGND 0.11584f
C14580 VPWR.n2347 VGND 0.01496f
C14581 VPWR.n2349 VGND 0.0901f
C14582 VPWR.t1684 VGND 0.09955f
C14583 VPWR.t1164 VGND 0.06535f
C14584 VPWR.t753 VGND 0.07675f
C14585 VPWR.t1325 VGND 0.06535f
C14586 VPWR.t745 VGND 0.09955f
C14587 VPWR.n2350 VGND 0.0901f
C14588 VPWR.n2352 VGND 0.01496f
C14589 VPWR.n2353 VGND 0.11584f
C14590 VPWR.n2354 VGND 0.06953f
C14591 VPWR.n2355 VGND 0.06953f
C14592 VPWR.n2356 VGND 0.11584f
C14593 VPWR.n2357 VGND 0.01496f
C14594 VPWR.n2359 VGND 0.0901f
C14595 VPWR.t1605 VGND 0.09955f
C14596 VPWR.t1324 VGND 0.06535f
C14597 VPWR.t1569 VGND 0.07675f
C14598 VPWR.t1161 VGND 0.06535f
C14599 VPWR.t1573 VGND 0.09955f
C14600 VPWR.n2360 VGND 0.0901f
C14601 VPWR.n2362 VGND 0.01496f
C14602 VPWR.n2363 VGND 0.11584f
C14603 VPWR.n2364 VGND 0.06953f
C14604 VPWR.n2365 VGND 0.06953f
C14605 VPWR.n2366 VGND 0.11584f
C14606 VPWR.n2367 VGND 0.01496f
C14607 VPWR.n2369 VGND 0.0901f
C14608 VPWR.t1077 VGND 0.09955f
C14609 VPWR.t1160 VGND 0.06535f
C14610 VPWR.t1879 VGND 0.07675f
C14611 VPWR.t1328 VGND 0.06535f
C14612 VPWR.t412 VGND 0.09955f
C14613 VPWR.n2370 VGND 0.0901f
C14614 VPWR.n2372 VGND 0.01496f
C14615 VPWR.n2373 VGND 0.11584f
C14616 VPWR.n2374 VGND 0.06953f
C14617 VPWR.n2375 VGND 0.06953f
C14618 VPWR.n2376 VGND 0.11584f
C14619 VPWR.n2377 VGND 0.01496f
C14620 VPWR.n2379 VGND 0.0901f
C14621 VPWR.t1846 VGND 0.09955f
C14622 VPWR.t1732 VGND 0.06535f
C14623 VPWR.t148 VGND 0.11101f
C14624 VPWR.n2380 VGND 0.06343f
C14625 VPWR.n2381 VGND 0.01496f
C14626 VPWR.n2382 VGND 0.11584f
C14627 VPWR.n2383 VGND 0.16128f
C14628 VPWR.n2384 VGND 0.84572f
C14629 VPWR.n2385 VGND 0.06953f
C14630 VPWR.n2386 VGND 0.06953f
C14631 VPWR.n2387 VGND 0.06953f
C14632 VPWR.n2388 VGND 0.06953f
C14633 VPWR.n2389 VGND 0.06953f
C14634 VPWR.n2390 VGND 0.06953f
C14635 VPWR.n2391 VGND 0.06953f
C14636 VPWR.n2392 VGND 0.06953f
C14637 VPWR.n2393 VGND 0.06953f
C14638 VPWR.n2394 VGND 0.06953f
C14639 VPWR.n2395 VGND 0.06953f
C14640 VPWR.n2396 VGND 0.06953f
C14641 VPWR.n2397 VGND 0.06953f
C14642 VPWR.n2398 VGND 0.06953f
C14643 VPWR.n2399 VGND 0.06953f
C14644 VPWR.n2400 VGND 0.16128f
C14645 VPWR.n2401 VGND 0.84572f
C14646 VPWR.n2402 VGND 0.84572f
C14647 VPWR.n2403 VGND 0.16128f
C14648 VPWR.n2404 VGND 0.11584f
C14649 VPWR.n2405 VGND 0.01496f
C14650 VPWR.n2406 VGND 0.06343f
C14651 VPWR.t315 VGND 0.11101f
C14652 VPWR.t1165 VGND 0.06535f
C14653 VPWR.t608 VGND 0.09955f
C14654 VPWR.n2407 VGND 0.0901f
C14655 VPWR.n2409 VGND 0.01496f
C14656 VPWR.n2410 VGND 0.11584f
C14657 VPWR.n2411 VGND 0.06953f
C14658 VPWR.n2412 VGND 0.06953f
C14659 VPWR.n2413 VGND 0.11584f
C14660 VPWR.n2414 VGND 0.01496f
C14661 VPWR.n2416 VGND 0.0901f
C14662 VPWR.t761 VGND 0.07675f
C14663 VPWR.t765 VGND 0.06535f
C14664 VPWR.t1717 VGND 0.09955f
C14665 VPWR.n2417 VGND 0.0901f
C14666 VPWR.n2419 VGND 0.01496f
C14667 VPWR.n2420 VGND 0.11584f
C14668 VPWR.n2421 VGND 0.06953f
C14669 VPWR.n2422 VGND 0.06953f
C14670 VPWR.n2423 VGND 0.11584f
C14671 VPWR.n2424 VGND 0.01496f
C14672 VPWR.n2426 VGND 0.0901f
C14673 VPWR.t1840 VGND 0.07675f
C14674 VPWR.t919 VGND 0.06535f
C14675 VPWR.t1322 VGND 0.09955f
C14676 VPWR.n2427 VGND 0.0901f
C14677 VPWR.n2429 VGND 0.01496f
C14678 VPWR.n2430 VGND 0.11584f
C14679 VPWR.n2431 VGND 0.06953f
C14680 VPWR.n2432 VGND 0.06953f
C14681 VPWR.n2433 VGND 0.11584f
C14682 VPWR.n2434 VGND 0.01496f
C14683 VPWR.n2436 VGND 0.0901f
C14684 VPWR.t1870 VGND 0.07675f
C14685 VPWR.t1220 VGND 0.06535f
C14686 VPWR.t947 VGND 0.09955f
C14687 VPWR.n2437 VGND 0.0901f
C14688 VPWR.n2439 VGND 0.01496f
C14689 VPWR.n2440 VGND 0.11584f
C14690 VPWR.n2441 VGND 0.06953f
C14691 VPWR.n2442 VGND 0.06953f
C14692 VPWR.n2443 VGND 0.11584f
C14693 VPWR.n2444 VGND 0.01496f
C14694 VPWR.n2446 VGND 0.0901f
C14695 VPWR.t894 VGND 0.07675f
C14696 VPWR.t1167 VGND 0.06535f
C14697 VPWR.t812 VGND 0.09955f
C14698 VPWR.n2447 VGND 0.0901f
C14699 VPWR.n2449 VGND 0.01496f
C14700 VPWR.n2450 VGND 0.11584f
C14701 VPWR.n2451 VGND 0.06953f
C14702 VPWR.n2452 VGND 0.06953f
C14703 VPWR.n2453 VGND 0.11584f
C14704 VPWR.n2454 VGND 0.01496f
C14705 VPWR.n2456 VGND 0.0901f
C14706 VPWR.t1140 VGND 0.07675f
C14707 VPWR.t1219 VGND 0.06535f
C14708 VPWR.t1547 VGND 0.09955f
C14709 VPWR.n2457 VGND 0.0901f
C14710 VPWR.n2459 VGND 0.01496f
C14711 VPWR.n2460 VGND 0.11584f
C14712 VPWR.n2461 VGND 0.06953f
C14713 VPWR.n2462 VGND 0.06953f
C14714 VPWR.n2463 VGND 0.11584f
C14715 VPWR.n2464 VGND 0.01496f
C14716 VPWR.n2466 VGND 0.0901f
C14717 VPWR.t1278 VGND 0.07675f
C14718 VPWR.t921 VGND 0.06535f
C14719 VPWR.t1458 VGND 0.09955f
C14720 VPWR.n2467 VGND 0.0901f
C14721 VPWR.n2469 VGND 0.01496f
C14722 VPWR.n2470 VGND 0.11584f
C14723 VPWR.n2471 VGND 0.06953f
C14724 VPWR.n2472 VGND 0.06953f
C14725 VPWR.n2473 VGND 0.11584f
C14726 VPWR.n2474 VGND 0.01496f
C14727 VPWR.n2476 VGND 0.0901f
C14728 VPWR.t1561 VGND 0.07675f
C14729 VPWR.t1221 VGND 0.06535f
C14730 VPWR.t1020 VGND 0.09955f
C14731 VPWR.n2477 VGND 0.0901f
C14732 VPWR.n2479 VGND 0.01496f
C14733 VPWR.n2480 VGND 0.11584f
C14734 VPWR.n2481 VGND 0.06953f
C14735 VPWR.n2482 VGND 0.84042f
C14736 VPWR.n2483 VGND 0.16128f
C14737 VPWR.n2484 VGND 0.06953f
C14738 VPWR.n2485 VGND 0.06953f
C14739 VPWR.n2486 VGND 0.06953f
C14740 VPWR.n2487 VGND 0.06953f
C14741 VPWR.n2488 VGND 0.06953f
C14742 VPWR.n2489 VGND 0.06953f
C14743 VPWR.n2490 VGND 0.06953f
C14744 VPWR.n2491 VGND 0.06953f
C14745 VPWR.n2492 VGND 0.06953f
C14746 VPWR.n2493 VGND 0.06953f
C14747 VPWR.n2494 VGND 0.06953f
C14748 VPWR.n2495 VGND 0.06953f
C14749 VPWR.n2496 VGND 0.06953f
C14750 VPWR.n2497 VGND 0.06953f
C14751 VPWR.n2498 VGND 0.06953f
C14752 VPWR.n2499 VGND 0.84042f
C14753 VPWR.n2500 VGND 0.47566f
C14754 VPWR.n2501 VGND 0.06953f
C14755 VPWR.n2502 VGND 0.07205f
C14756 VPWR.n2504 VGND 0.01427f
C14757 VPWR.n2506 VGND 0.0901f
C14758 VPWR.t197 VGND 0.09955f
C14759 VPWR.t164 VGND 0.06535f
C14760 VPWR.t288 VGND 0.07675f
C14761 VPWR.t294 VGND 0.06535f
C14762 VPWR.t309 VGND 0.09955f
C14763 VPWR.n2507 VGND 0.0901f
C14764 VPWR.n2509 VGND 0.01427f
C14765 VPWR.n2511 VGND 0.07205f
C14766 VPWR.n2512 VGND 0.06953f
C14767 VPWR.n2513 VGND 0.06953f
C14768 VPWR.n2514 VGND 0.07205f
C14769 VPWR.n2516 VGND 0.01427f
C14770 VPWR.n2518 VGND 0.0901f
C14771 VPWR.t74 VGND 0.09955f
C14772 VPWR.t334 VGND 0.06535f
C14773 VPWR.t68 VGND 0.07675f
C14774 VPWR.t58 VGND 0.06535f
C14775 VPWR.t185 VGND 0.09955f
C14776 VPWR.n2519 VGND 0.0901f
C14777 VPWR.n2521 VGND 0.01427f
C14778 VPWR.n2523 VGND 0.07205f
C14779 VPWR.n2524 VGND 0.06953f
C14780 VPWR.n2525 VGND 0.06953f
C14781 VPWR.n2526 VGND 0.07205f
C14782 VPWR.n2528 VGND 0.01427f
C14783 VPWR.n2530 VGND 0.0901f
C14784 VPWR.t194 VGND 0.09955f
C14785 VPWR.t202 VGND 0.06535f
C14786 VPWR.t331 VGND 0.07675f
C14787 VPWR.t226 VGND 0.06535f
C14788 VPWR.t350 VGND 0.09955f
C14789 VPWR.n2531 VGND 0.0901f
C14790 VPWR.n2533 VGND 0.01427f
C14791 VPWR.n2535 VGND 0.07205f
C14792 VPWR.n2536 VGND 0.06953f
C14793 VPWR.n2537 VGND 0.06953f
C14794 VPWR.n2538 VGND 0.07205f
C14795 VPWR.n2540 VGND 0.01427f
C14796 VPWR.n2542 VGND 0.0901f
C14797 VPWR.t71 VGND 0.09955f
C14798 VPWR.t63 VGND 0.06535f
C14799 VPWR.t90 VGND 0.07675f
C14800 VPWR.t98 VGND 0.06535f
C14801 VPWR.t231 VGND 0.09955f
C14802 VPWR.n2543 VGND 0.0901f
C14803 VPWR.n2545 VGND 0.01427f
C14804 VPWR.n2547 VGND 0.07205f
C14805 VPWR.n2548 VGND 0.06953f
C14806 VPWR.n2549 VGND 0.06953f
C14807 VPWR.n2550 VGND 0.07205f
C14808 VPWR.n2552 VGND 0.01427f
C14809 VPWR.n2554 VGND 0.0901f
C14810 VPWR.t247 VGND 0.09955f
C14811 VPWR.t200 VGND 0.06535f
C14812 VPWR.t328 VGND 0.07675f
C14813 VPWR.t361 VGND 0.06535f
C14814 VPWR.t377 VGND 0.09955f
C14815 VPWR.n2555 VGND 0.0901f
C14816 VPWR.n2557 VGND 0.01427f
C14817 VPWR.n2559 VGND 0.07205f
C14818 VPWR.n2560 VGND 0.06953f
C14819 VPWR.n2561 VGND 0.06953f
C14820 VPWR.n2562 VGND 0.07205f
C14821 VPWR.n2564 VGND 0.01427f
C14822 VPWR.n2566 VGND 0.0901f
C14823 VPWR.t121 VGND 0.09955f
C14824 VPWR.t380 VGND 0.06535f
C14825 VPWR.t113 VGND 0.07675f
C14826 VPWR.t234 VGND 0.06535f
C14827 VPWR.t151 VGND 0.09955f
C14828 VPWR.n2567 VGND 0.0901f
C14829 VPWR.n2569 VGND 0.01427f
C14830 VPWR.n2571 VGND 0.07205f
C14831 VPWR.n2572 VGND 0.06953f
C14832 VPWR.n2573 VGND 0.06953f
C14833 VPWR.n2574 VGND 0.07205f
C14834 VPWR.n2576 VGND 0.01427f
C14835 VPWR.n2578 VGND 0.0901f
C14836 VPWR.t1 VGND 0.09955f
C14837 VPWR.t253 VGND 0.06535f
C14838 VPWR.t374 VGND 0.07675f
C14839 VPWR.t278 VGND 0.06535f
C14840 VPWR.t20 VGND 0.09955f
C14841 VPWR.n2579 VGND 0.0901f
C14842 VPWR.n2581 VGND 0.01427f
C14843 VPWR.n2583 VGND 0.07205f
C14844 VPWR.n2584 VGND 0.06953f
C14845 VPWR.n2585 VGND 0.06953f
C14846 VPWR.n2586 VGND 0.07205f
C14847 VPWR.n2588 VGND 0.01427f
C14848 VPWR.n2590 VGND 0.0901f
C14849 VPWR.t145 VGND 0.09955f
C14850 VPWR.t129 VGND 0.06535f
C14851 VPWR.t250 VGND 0.11101f
C14852 VPWR.n2591 VGND 0.0634f
C14853 VPWR.n2592 VGND 0.01414f
C14854 VPWR.n2594 VGND 0.09036f
C14855 VPWR.n2595 VGND 0.16128f
C14856 VPWR.n2596 VGND 2.21691f
C14857 VPWR.n2597 VGND 0.90282f
C14858 VPWR.n2598 VGND 0.37828f
C14859 VPWR.t1090 VGND 0.04542f
C14860 VPWR.t1364 VGND 0.04542f
C14861 VPWR.n2599 VGND 0.08241f
C14862 VPWR.n2600 VGND 0.03902f
C14863 VPWR.t1088 VGND 0.01193f
C14864 VPWR.t1096 VGND 0.01193f
C14865 VPWR.n2601 VGND 0.02561f
C14866 VPWR.t1369 VGND 0.01193f
C14867 VPWR.t1363 VGND 0.01193f
C14868 VPWR.n2602 VGND 0.02561f
C14869 VPWR.n2604 VGND 0.03902f
C14870 VPWR.t1813 VGND 0.01193f
C14871 VPWR.t1794 VGND 0.01193f
C14872 VPWR.n2605 VGND 0.02561f
C14873 VPWR.t1777 VGND 0.01193f
C14874 VPWR.t1783 VGND 0.01193f
C14875 VPWR.n2606 VGND 0.02561f
C14876 VPWR.t1790 VGND 0.04757f
C14877 VPWR.t1769 VGND 0.04757f
C14878 VPWR.n2607 VGND 0.1097f
C14879 VPWR.n2608 VGND 0.0352f
C14880 VPWR.n2609 VGND 0.01134f
C14881 VPWR.n2610 VGND 0.05148f
C14882 VPWR.t1771 VGND 0.01193f
C14883 VPWR.t1094 VGND 0.01193f
C14884 VPWR.n2612 VGND 0.02561f
C14885 VPWR.t1789 VGND 0.01193f
C14886 VPWR.t1367 VGND 0.01193f
C14887 VPWR.n2613 VGND 0.02561f
C14888 VPWR.n2614 VGND 0.05148f
C14889 VPWR.n2615 VGND 0.01187f
C14890 VPWR.n2616 VGND 0.03902f
C14891 VPWR.n2617 VGND 0.03902f
C14892 VPWR.n2618 VGND 0.03902f
C14893 VPWR.n2619 VGND 0.01067f
C14894 VPWR.n2620 VGND 0.05148f
C14895 VPWR.n2621 VGND 0.01006f
C14896 VPWR.n2623 VGND 0.03902f
C14897 VPWR.n2624 VGND 0.02927f
C14898 VPWR.t1768 VGND 0.14254f
C14899 VPWR.t1776 VGND 0.21006f
C14900 VPWR.t1782 VGND 0.21006f
C14901 VPWR.t1770 VGND 0.21006f
C14902 VPWR.t1093 VGND 0.21006f
C14903 VPWR.t1087 VGND 0.21006f
C14904 VPWR.t1095 VGND 0.21006f
C14905 VPWR.t1089 VGND 0.46766f
C14906 VPWR.n2626 VGND 0.51043f
C14907 VPWR.n2627 VGND 0.01484f
C14908 VPWR.n2628 VGND 0.8953f
C14909 VPWR.n2629 VGND 0.03902f
C14910 VPWR.t1766 VGND 0.14254f
C14911 VPWR.t1779 VGND 0.21006f
C14912 VPWR.t1753 VGND 0.21006f
C14913 VPWR.t1805 VGND 0.21006f
C14914 VPWR.t576 VGND 0.21006f
C14915 VPWR.t671 VGND 0.21006f
C14916 VPWR.t574 VGND 0.21006f
C14917 VPWR.t675 VGND 0.34509f
C14918 VPWR.t975 VGND 0.36635f
C14919 VPWR.n2630 VGND 0.51698f
C14920 VPWR.n2631 VGND 0.14706f
C14921 VPWR.n2632 VGND 0.03902f
C14922 VPWR.t1864 VGND 0.01193f
C14923 VPWR.t575 VGND 0.01193f
C14924 VPWR.n2633 VGND 0.02561f
C14925 VPWR.t672 VGND 0.01193f
C14926 VPWR.t682 VGND 0.01193f
C14927 VPWR.n2634 VGND 0.02561f
C14928 VPWR.n2635 VGND 0.05148f
C14929 VPWR.n2636 VGND 0.03902f
C14930 VPWR.t1816 VGND 0.01193f
C14931 VPWR.t577 VGND 0.01193f
C14932 VPWR.n2637 VGND 0.02561f
C14933 VPWR.t1806 VGND 0.01193f
C14934 VPWR.t679 VGND 0.01193f
C14935 VPWR.n2638 VGND 0.02561f
C14936 VPWR.t1767 VGND 0.04757f
C14937 VPWR.t1815 VGND 0.04757f
C14938 VPWR.n2640 VGND 0.1097f
C14939 VPWR.t1798 VGND 0.01193f
C14940 VPWR.t1773 VGND 0.01193f
C14941 VPWR.n2641 VGND 0.02561f
C14942 VPWR.t1780 VGND 0.01193f
C14943 VPWR.t1754 VGND 0.01193f
C14944 VPWR.n2642 VGND 0.02561f
C14945 VPWR.n2643 VGND 0.05148f
C14946 VPWR.n2644 VGND 0.01134f
C14947 VPWR.n2645 VGND 0.0352f
C14948 VPWR.n2646 VGND 0.03902f
C14949 VPWR.n2647 VGND 0.03902f
C14950 VPWR.n2648 VGND 0.01187f
C14951 VPWR.n2649 VGND 0.05148f
C14952 VPWR.n2651 VGND 0.01067f
C14953 VPWR.n2652 VGND 0.03902f
C14954 VPWR.n2653 VGND 0.03902f
C14955 VPWR.n2654 VGND 0.01006f
C14956 VPWR.t1863 VGND 0.04542f
C14957 VPWR.t676 VGND 0.04542f
C14958 VPWR.n2656 VGND 0.08241f
C14959 VPWR.n2658 VGND 0.02927f
C14960 VPWR.n2659 VGND 0.01484f
C14961 VPWR.n2660 VGND 0.02927f
C14962 VPWR.n2661 VGND 0.01164f
C14963 VPWR.t976 VGND 0.04752f
C14964 VPWR.t1869 VGND 0.04752f
C14965 VPWR.n2663 VGND 0.09606f
C14966 VPWR.n2664 VGND 0.02715f
C14967 VPWR.n2665 VGND 1.36261f
C14968 VPWR.n2666 VGND 0.03902f
C14969 VPWR.t597 VGND 0.04665f
C14970 VPWR.t1800 VGND 0.14254f
C14971 VPWR.t1757 VGND 0.21006f
C14972 VPWR.t1807 VGND 0.21006f
C14973 VPWR.t1784 VGND 0.21006f
C14974 VPWR.t459 VGND 0.21006f
C14975 VPWR.t453 VGND 0.21006f
C14976 VPWR.t461 VGND 0.21006f
C14977 VPWR.t455 VGND 0.34509f
C14978 VPWR.t1401 VGND 0.13254f
C14979 VPWR.t596 VGND 0.10503f
C14980 VPWR.t928 VGND 0.23381f
C14981 VPWR.n2667 VGND 0.45821f
C14982 VPWR.n2668 VGND 0.14488f
C14983 VPWR.n2669 VGND 0.03902f
C14984 VPWR.t454 VGND 0.01193f
C14985 VPWR.t462 VGND 0.01193f
C14986 VPWR.n2670 VGND 0.02561f
C14987 VPWR.t1178 VGND 0.01193f
C14988 VPWR.t595 VGND 0.01193f
C14989 VPWR.n2671 VGND 0.02561f
C14990 VPWR.n2672 VGND 0.05148f
C14991 VPWR.n2673 VGND 0.03902f
C14992 VPWR.t1802 VGND 0.01193f
C14993 VPWR.t460 VGND 0.01193f
C14994 VPWR.n2674 VGND 0.02561f
C14995 VPWR.t1785 VGND 0.01193f
C14996 VPWR.t1000 VGND 0.01193f
C14997 VPWR.n2675 VGND 0.02561f
C14998 VPWR.t1814 VGND 0.04757f
C14999 VPWR.t1801 VGND 0.04757f
C15000 VPWR.n2677 VGND 0.1097f
C15001 VPWR.t1774 VGND 0.01193f
C15002 VPWR.t1820 VGND 0.01193f
C15003 VPWR.n2678 VGND 0.02561f
C15004 VPWR.t1758 VGND 0.01193f
C15005 VPWR.t1808 VGND 0.01193f
C15006 VPWR.n2679 VGND 0.02561f
C15007 VPWR.n2680 VGND 0.05148f
C15008 VPWR.n2681 VGND 0.01134f
C15009 VPWR.n2682 VGND 0.0352f
C15010 VPWR.n2683 VGND 0.03902f
C15011 VPWR.n2684 VGND 0.03902f
C15012 VPWR.n2685 VGND 0.01187f
C15013 VPWR.n2686 VGND 0.05148f
C15014 VPWR.n2688 VGND 0.01067f
C15015 VPWR.n2689 VGND 0.03902f
C15016 VPWR.n2690 VGND 0.03902f
C15017 VPWR.n2691 VGND 0.01006f
C15018 VPWR.t456 VGND 0.04542f
C15019 VPWR.t477 VGND 0.04542f
C15020 VPWR.n2693 VGND 0.08241f
C15021 VPWR.n2695 VGND 0.02927f
C15022 VPWR.n2696 VGND 0.01484f
C15023 VPWR.n2697 VGND 0.02927f
C15024 VPWR.t929 VGND 0.04758f
C15025 VPWR.n2698 VGND 0.0663f
C15026 VPWR.n2700 VGND 0.04852f
C15027 VPWR.t1402 VGND 0.04677f
C15028 VPWR.n2701 VGND 0.06062f
C15029 VPWR.n2702 VGND 0.02312f
C15030 VPWR.n2703 VGND 1.36261f
C15031 VPWR.n2704 VGND 0.03902f
C15032 VPWR.t1803 VGND 0.08084f
C15033 VPWR.t1761 VGND 0.11913f
C15034 VPWR.t1809 VGND 0.11582f
C15035 VPWR.t1787 VGND 0.18523f
C15036 VPWR.t1888 VGND 0.15754f
C15037 VPWR.t1791 VGND 0.10503f
C15038 VPWR.t1894 VGND 0.10503f
C15039 VPWR.t1763 VGND 0.10503f
C15040 VPWR.t578 VGND 0.10503f
C15041 VPWR.t1795 VGND 0.10503f
C15042 VPWR.t1892 VGND 0.10503f
C15043 VPWR.t1818 VGND 0.14629f
C15044 VPWR.t1536 VGND 0.08252f
C15045 VPWR.t1290 VGND 0.09002f
C15046 VPWR.t1670 VGND 0.10503f
C15047 VPWR.t1292 VGND 0.19505f
C15048 VPWR.n2705 VGND 0.31443f
C15049 VPWR.n2706 VGND 0.14503f
C15050 VPWR.t1293 VGND 0.04722f
C15051 VPWR.n2707 VGND 0.03902f
C15052 VPWR.t1819 VGND 0.04668f
C15053 VPWR.t1893 VGND 0.04494f
C15054 VPWR.t1764 VGND 0.01193f
C15055 VPWR.t1796 VGND 0.01193f
C15056 VPWR.n2708 VGND 0.02561f
C15057 VPWR.t1895 VGND 0.01193f
C15058 VPWR.t579 VGND 0.01193f
C15059 VPWR.n2709 VGND 0.02561f
C15060 VPWR.n2710 VGND 0.0292f
C15061 VPWR.n2711 VGND 0.03902f
C15062 VPWR.t1788 VGND 0.01193f
C15063 VPWR.t1889 VGND 0.01193f
C15064 VPWR.n2712 VGND 0.02561f
C15065 VPWR.t1804 VGND 0.04757f
C15066 VPWR.n2714 VGND 0.05995f
C15067 VPWR.t1762 VGND 0.01193f
C15068 VPWR.t1810 VGND 0.01193f
C15069 VPWR.n2715 VGND 0.02561f
C15070 VPWR.n2716 VGND 0.0292f
C15071 VPWR.n2717 VGND 0.01134f
C15072 VPWR.n2718 VGND 0.0352f
C15073 VPWR.n2719 VGND 0.03902f
C15074 VPWR.n2720 VGND 0.03902f
C15075 VPWR.n2721 VGND 0.01187f
C15076 VPWR.n2722 VGND 0.02852f
C15077 VPWR.t1792 VGND 0.04175f
C15078 VPWR.n2723 VGND 0.03329f
C15079 VPWR.n2725 VGND 0.03902f
C15080 VPWR.n2726 VGND 0.03902f
C15081 VPWR.n2727 VGND 0.03235f
C15082 VPWR.n2728 VGND 0.01006f
C15083 VPWR.n2729 VGND 0.04282f
C15084 VPWR.n2730 VGND 0.05641f
C15085 VPWR.n2732 VGND 0.02312f
C15086 VPWR.n2733 VGND 0.01484f
C15087 VPWR.n2734 VGND 0.02927f
C15088 VPWR.t1671 VGND 0.04762f
C15089 VPWR.n2735 VGND 0.12244f
C15090 VPWR.t1291 VGND 0.04755f
C15091 VPWR.n2737 VGND 0.05293f
C15092 VPWR.n2738 VGND 0.0229f
C15093 VPWR.n2739 VGND 1.36261f
C15094 VPWR.n2740 VGND 0.0352f
C15095 VPWR.t1797 VGND 0.55515f
C15096 VPWR.t1756 VGND 0.21006f
C15097 VPWR.t1786 VGND 0.21006f
C15098 VPWR.t1760 VGND 0.21006f
C15099 VPWR.t1097 VGND 0.21006f
C15100 VPWR.t1091 VGND 0.21006f
C15101 VPWR.t1099 VGND 0.21006f
C15102 VPWR.t1101 VGND 0.19005f
C15103 VPWR.t445 VGND 0.46012f
C15104 VPWR.t1746 VGND 0.12753f
C15105 VPWR.n2741 VGND 0.27567f
C15106 VPWR.n2742 VGND 0.14706f
C15107 VPWR.t1098 VGND 0.01193f
C15108 VPWR.t1092 VGND 0.01193f
C15109 VPWR.n2743 VGND 0.02615f
C15110 VPWR.t1366 VGND 0.01193f
C15111 VPWR.t1365 VGND 0.01193f
C15112 VPWR.n2744 VGND 0.02615f
C15113 VPWR.n2745 VGND 0.09924f
C15114 VPWR.n2746 VGND 0.08046f
C15115 VPWR.t1100 VGND 0.01193f
C15116 VPWR.t1102 VGND 0.01193f
C15117 VPWR.n2747 VGND 0.02619f
C15118 VPWR.t1368 VGND 0.01193f
C15119 VPWR.t1362 VGND 0.01193f
C15120 VPWR.n2748 VGND 0.02619f
C15121 VPWR.n2749 VGND 0.10878f
C15122 VPWR.n2751 VGND 0.31423f
C15123 VPWR.n2752 VGND 0.01484f
C15124 VPWR.n2753 VGND 0.01357f
C15125 VPWR.n2754 VGND 0.01164f
C15126 VPWR.n2755 VGND 0.01089f
C15127 VPWR.t446 VGND 0.04762f
C15128 VPWR.t1535 VGND 0.04762f
C15129 VPWR.n2756 VGND 0.14066f
C15130 VPWR.n2757 VGND 0.02927f
C15131 VPWR.n2758 VGND 1.36261f
C15132 VPWR.n2759 VGND 0.0352f
C15133 VPWR.t1778 VGND 0.55515f
C15134 VPWR.t1811 VGND 0.21006f
C15135 VPWR.t1765 VGND 0.21006f
C15136 VPWR.t1812 VGND 0.21006f
C15137 VPWR.t572 VGND 0.21006f
C15138 VPWR.t680 VGND 0.21006f
C15139 VPWR.t673 VGND 0.21006f
C15140 VPWR.t677 VGND 0.19005f
C15141 VPWR.t386 VGND 0.40886f
C15142 VPWR.t1748 VGND 0.09002f
C15143 VPWR.t1752 VGND 0.08877f
C15144 VPWR.n2760 VGND 0.27442f
C15145 VPWR.n2761 VGND 0.14706f
C15146 VPWR.t573 VGND 0.01193f
C15147 VPWR.t1862 VGND 0.01193f
C15148 VPWR.n2762 VGND 0.02615f
C15149 VPWR.t670 VGND 0.01193f
C15150 VPWR.t681 VGND 0.01193f
C15151 VPWR.n2763 VGND 0.02615f
C15152 VPWR.n2764 VGND 0.09924f
C15153 VPWR.n2765 VGND 0.08046f
C15154 VPWR.t1907 VGND 0.01193f
C15155 VPWR.t1906 VGND 0.01193f
C15156 VPWR.n2766 VGND 0.02619f
C15157 VPWR.t674 VGND 0.01193f
C15158 VPWR.t678 VGND 0.01193f
C15159 VPWR.n2767 VGND 0.02619f
C15160 VPWR.n2768 VGND 0.10878f
C15161 VPWR.n2770 VGND 0.31423f
C15162 VPWR.n2771 VGND 0.01484f
C15163 VPWR.n2772 VGND 0.01336f
C15164 VPWR.t1749 VGND 0.04752f
C15165 VPWR.n2774 VGND 0.0508f
C15166 VPWR.t387 VGND 0.04762f
C15167 VPWR.n2776 VGND 0.07585f
C15168 VPWR.n2777 VGND 0.02927f
C15169 VPWR.n2778 VGND 1.36261f
C15170 VPWR.n2779 VGND 0.03563f
C15171 VPWR.t1759 VGND 0.55515f
C15172 VPWR.t1772 VGND 0.21006f
C15173 VPWR.t1799 VGND 0.21006f
C15174 VPWR.t1775 VGND 0.21006f
C15175 VPWR.t463 VGND 0.21006f
C15176 VPWR.t457 VGND 0.21006f
C15177 VPWR.t449 VGND 0.21006f
C15178 VPWR.t451 VGND 0.19005f
C15179 VPWR.t447 VGND 0.43512f
C15180 VPWR.t1744 VGND 0.15004f
C15181 VPWR.n2780 VGND 0.27316f
C15182 VPWR.n2781 VGND 0.14488f
C15183 VPWR.t1747 VGND 0.04759f
C15184 VPWR.t464 VGND 0.01193f
C15185 VPWR.t458 VGND 0.01193f
C15186 VPWR.n2782 VGND 0.02615f
C15187 VPWR.t985 VGND 0.01193f
C15188 VPWR.t1048 VGND 0.01193f
C15189 VPWR.n2783 VGND 0.02615f
C15190 VPWR.n2784 VGND 0.09924f
C15191 VPWR.n2785 VGND 0.08046f
C15192 VPWR.t450 VGND 0.01193f
C15193 VPWR.t452 VGND 0.01193f
C15194 VPWR.n2786 VGND 0.02619f
C15195 VPWR.t986 VGND 0.01193f
C15196 VPWR.t830 VGND 0.01193f
C15197 VPWR.n2787 VGND 0.02619f
C15198 VPWR.n2788 VGND 0.10878f
C15199 VPWR.n2790 VGND 0.31423f
C15200 VPWR.n2791 VGND 0.01484f
C15201 VPWR.n2792 VGND 0.01315f
C15202 VPWR.t1745 VGND 0.04759f
C15203 VPWR.n2793 VGND 0.12538f
C15204 VPWR.n2794 VGND 0.01006f
C15205 VPWR.t448 VGND 0.04758f
C15206 VPWR.t1534 VGND 0.04758f
C15207 VPWR.n2795 VGND 0.11195f
C15208 VPWR.n2796 VGND 0.02927f
C15209 VPWR.n2797 VGND 1.36261f
C15210 VPWR.n2798 VGND 0.03563f
C15211 VPWR.t385 VGND 0.04758f
C15212 VPWR.n2799 VGND 0.01315f
C15213 VPWR.t1751 VGND 0.04759f
C15214 VPWR.n2800 VGND 0.01484f
C15215 VPWR.t1793 VGND 0.31484f
C15216 VPWR.t1817 VGND 0.11913f
C15217 VPWR.t1781 VGND 0.11913f
C15218 VPWR.t1755 VGND 0.11913f
C15219 VPWR.t1890 VGND 0.11913f
C15220 VPWR.t683 VGND 0.11913f
C15221 VPWR.t693 VGND 0.11913f
C15222 VPWR.t558 VGND 0.10779f
C15223 VPWR.t384 VGND 0.24677f
C15224 VPWR.t1750 VGND 0.08509f
C15225 VPWR.n2801 VGND 0.15203f
C15226 VPWR.t694 VGND 0.01193f
C15227 VPWR.t559 VGND 0.01193f
C15228 VPWR.n2802 VGND 0.02619f
C15229 VPWR.n2803 VGND 0.06446f
C15230 VPWR.t1891 VGND 0.01193f
C15231 VPWR.t684 VGND 0.01193f
C15232 VPWR.n2804 VGND 0.02726f
C15233 VPWR.n2805 VGND 0.14554f
C15234 VPWR.n2806 VGND 0.31423f
C15235 VPWR.n2808 VGND 0.08044f
C15236 VPWR.n2809 VGND 0.07062f
C15237 VPWR.n2810 VGND 0.01006f
C15238 VPWR.n2811 VGND 0.06119f
C15239 VPWR.n2812 VGND 0.02927f
C15240 VPWR.n2813 VGND 1.98291f
C15241 VPWR.n2814 VGND 1.6059f
C15242 VPWR.t1042 VGND 0.02419f
C15243 VPWR.n2815 VGND 0.10843f
C15244 VPWR.n2816 VGND 0.23867f
C15245 VPWR.n2817 VGND 0.06294f
C15246 VPWR.n2818 VGND 0.02989f
C15247 VPWR.n2819 VGND 0.0365f
C15248 VPWR.n2820 VGND 0.07398f
C15249 VPWR.n2821 VGND 0.09644f
C15250 VPWR.n2822 VGND 0.07398f
C15251 VPWR.t570 VGND 2.32707f
C15252 VPWR.t1041 VGND 0.73498f
C15253 VPWR.n2823 VGND 0.0972f
C15254 VPWR.n2824 VGND 0.38456f
C15255 VPWR.t571 VGND 0.02418f
C15256 VPWR.n2825 VGND 0.14806f
C15257 VPWR.n2826 VGND 0.01495f
C15258 VPWR.n2827 VGND 0.08157f
C15259 VPWR.n2828 VGND 0.07323f
C15260 VPWR.n2829 VGND 0.0972f
C15261 VPWR.n2830 VGND 0.06121f
C15262 VPWR.t1127 VGND 0.02418f
C15263 VPWR.n2831 VGND 0.14806f
C15264 VPWR.n2832 VGND 0.01495f
C15265 VPWR.n2833 VGND 0.0972f
C15266 VPWR.n2834 VGND 0.06361f
C15267 VPWR.n2835 VGND 0.07255f
C15268 VPWR.n2836 VGND 1.39067f
C15269 VPWR.n2837 VGND 0.07255f
C15270 VPWR.n2838 VGND 0.06361f
C15271 VPWR.n2839 VGND 0.0972f
C15272 VPWR.n2840 VGND 0.08149f
C15273 VPWR.n2841 VGND 0.06741f
C15274 VPWR.n2842 VGND 0.83594f
C15275 VPWR.n2843 VGND 0.0526f
C15276 VPWR.n2844 VGND 0.07357f
C15277 VPWR.n2845 VGND 0.05115f
C15278 VPWR.n2846 VGND 0.01495f
C15279 VPWR.n2847 VGND 0.0526f
C15280 VPWR.n2848 VGND 0.04039f
C15281 VPWR.n2849 VGND 0.1445f
C15282 VPWR.n2850 VGND 0.05693f
C15283 VPWR.n2851 VGND 0.0365f
C15284 VPWR.t1403 VGND 0.28776f
C15285 VPWR.n2852 VGND 0.06741f
C15286 VPWR.n2853 VGND 0.08149f
C15287 VPWR.n2854 VGND 0.02989f
C15288 VPWR.n2855 VGND 1.68424f
C15289 VPWR.n2856 VGND 0.02989f
C15290 VPWR.n2857 VGND 0.02989f
C15291 VPWR.n2858 VGND 0.07428f
C15292 VPWR.n2859 VGND 0.04078f
C15293 VPWR.n2860 VGND 0.31586f
C15294 VPWR.n2861 VGND 0.25988f
C15295 VPWR.t1404 VGND 0.02417f
C15296 VPWR.n2862 VGND 0.18289f
C15297 VPWR.n2863 VGND 2.89587f
C15298 XThR.Tn[2].t11 VGND 0.01864f
C15299 XThR.Tn[2].t8 VGND 0.01864f
C15300 XThR.Tn[2].n0 VGND 0.03762f
C15301 XThR.Tn[2].t10 VGND 0.01864f
C15302 XThR.Tn[2].t9 VGND 0.01864f
C15303 XThR.Tn[2].n1 VGND 0.04402f
C15304 XThR.Tn[2].n2 VGND 0.13203f
C15305 XThR.Tn[2].t6 VGND 0.01211f
C15306 XThR.Tn[2].t7 VGND 0.01211f
C15307 XThR.Tn[2].n3 VGND 0.02759f
C15308 XThR.Tn[2].t5 VGND 0.01211f
C15309 XThR.Tn[2].t4 VGND 0.01211f
C15310 XThR.Tn[2].n4 VGND 0.02759f
C15311 XThR.Tn[2].t2 VGND 0.01211f
C15312 XThR.Tn[2].t3 VGND 0.01211f
C15313 XThR.Tn[2].n5 VGND 0.02759f
C15314 XThR.Tn[2].t0 VGND 0.01211f
C15315 XThR.Tn[2].t1 VGND 0.01211f
C15316 XThR.Tn[2].n6 VGND 0.04596f
C15317 XThR.Tn[2].n7 VGND 0.13137f
C15318 XThR.Tn[2].n8 VGND 0.08121f
C15319 XThR.Tn[2].n9 VGND 0.09165f
C15320 XThR.Tn[2].t21 VGND 0.01457f
C15321 XThR.Tn[2].t14 VGND 0.01595f
C15322 XThR.Tn[2].n10 VGND 0.03895f
C15323 XThR.Tn[2].n11 VGND 0.07482f
C15324 XThR.Tn[2].t40 VGND 0.01457f
C15325 XThR.Tn[2].t31 VGND 0.01595f
C15326 XThR.Tn[2].n12 VGND 0.03895f
C15327 XThR.Tn[2].t55 VGND 0.01452f
C15328 XThR.Tn[2].t66 VGND 0.0159f
C15329 XThR.Tn[2].n13 VGND 0.04052f
C15330 XThR.Tn[2].n14 VGND 0.02847f
C15331 XThR.Tn[2].n16 VGND 0.09136f
C15332 XThR.Tn[2].t15 VGND 0.01457f
C15333 XThR.Tn[2].t67 VGND 0.01595f
C15334 XThR.Tn[2].n17 VGND 0.03895f
C15335 XThR.Tn[2].t30 VGND 0.01452f
C15336 XThR.Tn[2].t43 VGND 0.0159f
C15337 XThR.Tn[2].n18 VGND 0.04052f
C15338 XThR.Tn[2].n19 VGND 0.02847f
C15339 XThR.Tn[2].n21 VGND 0.09136f
C15340 XThR.Tn[2].t32 VGND 0.01457f
C15341 XThR.Tn[2].t23 VGND 0.01595f
C15342 XThR.Tn[2].n22 VGND 0.03895f
C15343 XThR.Tn[2].t47 VGND 0.01452f
C15344 XThR.Tn[2].t60 VGND 0.0159f
C15345 XThR.Tn[2].n23 VGND 0.04052f
C15346 XThR.Tn[2].n24 VGND 0.02847f
C15347 XThR.Tn[2].n26 VGND 0.09136f
C15348 XThR.Tn[2].t58 VGND 0.01457f
C15349 XThR.Tn[2].t50 VGND 0.01595f
C15350 XThR.Tn[2].n27 VGND 0.03895f
C15351 XThR.Tn[2].t16 VGND 0.01452f
C15352 XThR.Tn[2].t28 VGND 0.0159f
C15353 XThR.Tn[2].n28 VGND 0.04052f
C15354 XThR.Tn[2].n29 VGND 0.02847f
C15355 XThR.Tn[2].n31 VGND 0.09136f
C15356 XThR.Tn[2].t34 VGND 0.01457f
C15357 XThR.Tn[2].t25 VGND 0.01595f
C15358 XThR.Tn[2].n32 VGND 0.03895f
C15359 XThR.Tn[2].t48 VGND 0.01452f
C15360 XThR.Tn[2].t62 VGND 0.0159f
C15361 XThR.Tn[2].n33 VGND 0.04052f
C15362 XThR.Tn[2].n34 VGND 0.02847f
C15363 XThR.Tn[2].n36 VGND 0.09136f
C15364 XThR.Tn[2].t70 VGND 0.01457f
C15365 XThR.Tn[2].t41 VGND 0.01595f
C15366 XThR.Tn[2].n37 VGND 0.03895f
C15367 XThR.Tn[2].t22 VGND 0.01452f
C15368 XThR.Tn[2].t20 VGND 0.0159f
C15369 XThR.Tn[2].n38 VGND 0.04052f
C15370 XThR.Tn[2].n39 VGND 0.02847f
C15371 XThR.Tn[2].n41 VGND 0.09136f
C15372 XThR.Tn[2].t39 VGND 0.01457f
C15373 XThR.Tn[2].t35 VGND 0.01595f
C15374 XThR.Tn[2].n42 VGND 0.03895f
C15375 XThR.Tn[2].t54 VGND 0.01452f
C15376 XThR.Tn[2].t12 VGND 0.0159f
C15377 XThR.Tn[2].n43 VGND 0.04052f
C15378 XThR.Tn[2].n44 VGND 0.02847f
C15379 XThR.Tn[2].n46 VGND 0.09136f
C15380 XThR.Tn[2].t44 VGND 0.01457f
C15381 XThR.Tn[2].t49 VGND 0.01595f
C15382 XThR.Tn[2].n47 VGND 0.03895f
C15383 XThR.Tn[2].t57 VGND 0.01452f
C15384 XThR.Tn[2].t27 VGND 0.0159f
C15385 XThR.Tn[2].n48 VGND 0.04052f
C15386 XThR.Tn[2].n49 VGND 0.02847f
C15387 XThR.Tn[2].n51 VGND 0.09136f
C15388 XThR.Tn[2].t61 VGND 0.01457f
C15389 XThR.Tn[2].t69 VGND 0.01595f
C15390 XThR.Tn[2].n52 VGND 0.03895f
C15391 XThR.Tn[2].t18 VGND 0.01452f
C15392 XThR.Tn[2].t45 VGND 0.0159f
C15393 XThR.Tn[2].n53 VGND 0.04052f
C15394 XThR.Tn[2].n54 VGND 0.02847f
C15395 XThR.Tn[2].n56 VGND 0.09136f
C15396 XThR.Tn[2].t52 VGND 0.01457f
C15397 XThR.Tn[2].t26 VGND 0.01595f
C15398 XThR.Tn[2].n57 VGND 0.03895f
C15399 XThR.Tn[2].t68 VGND 0.01452f
C15400 XThR.Tn[2].t63 VGND 0.0159f
C15401 XThR.Tn[2].n58 VGND 0.04052f
C15402 XThR.Tn[2].n59 VGND 0.02847f
C15403 XThR.Tn[2].n61 VGND 0.09136f
C15404 XThR.Tn[2].t73 VGND 0.01457f
C15405 XThR.Tn[2].t64 VGND 0.01595f
C15406 XThR.Tn[2].n62 VGND 0.03895f
C15407 XThR.Tn[2].t24 VGND 0.01452f
C15408 XThR.Tn[2].t37 VGND 0.0159f
C15409 XThR.Tn[2].n63 VGND 0.04052f
C15410 XThR.Tn[2].n64 VGND 0.02847f
C15411 XThR.Tn[2].n66 VGND 0.09136f
C15412 XThR.Tn[2].t42 VGND 0.01457f
C15413 XThR.Tn[2].t36 VGND 0.01595f
C15414 XThR.Tn[2].n67 VGND 0.03895f
C15415 XThR.Tn[2].t56 VGND 0.01452f
C15416 XThR.Tn[2].t13 VGND 0.0159f
C15417 XThR.Tn[2].n68 VGND 0.04052f
C15418 XThR.Tn[2].n69 VGND 0.02847f
C15419 XThR.Tn[2].n71 VGND 0.09136f
C15420 XThR.Tn[2].t59 VGND 0.01457f
C15421 XThR.Tn[2].t51 VGND 0.01595f
C15422 XThR.Tn[2].n72 VGND 0.03895f
C15423 XThR.Tn[2].t17 VGND 0.01452f
C15424 XThR.Tn[2].t29 VGND 0.0159f
C15425 XThR.Tn[2].n73 VGND 0.04052f
C15426 XThR.Tn[2].n74 VGND 0.02847f
C15427 XThR.Tn[2].n76 VGND 0.09136f
C15428 XThR.Tn[2].t19 VGND 0.01457f
C15429 XThR.Tn[2].t72 VGND 0.01595f
C15430 XThR.Tn[2].n77 VGND 0.03895f
C15431 XThR.Tn[2].t33 VGND 0.01452f
C15432 XThR.Tn[2].t46 VGND 0.0159f
C15433 XThR.Tn[2].n78 VGND 0.04052f
C15434 XThR.Tn[2].n79 VGND 0.02847f
C15435 XThR.Tn[2].n81 VGND 0.09136f
C15436 XThR.Tn[2].t53 VGND 0.01457f
C15437 XThR.Tn[2].t65 VGND 0.01595f
C15438 XThR.Tn[2].n82 VGND 0.03895f
C15439 XThR.Tn[2].t71 VGND 0.01452f
C15440 XThR.Tn[2].t38 VGND 0.0159f
C15441 XThR.Tn[2].n83 VGND 0.04052f
C15442 XThR.Tn[2].n84 VGND 0.02847f
C15443 XThR.Tn[2].n86 VGND 0.09136f
C15444 XThR.Tn[2].n87 VGND 0.08302f
C15445 XThR.Tn[2].n88 VGND 0.17991f
.ends

