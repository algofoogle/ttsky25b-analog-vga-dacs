magic
tech sky130A
magscale 1 2
timestamp 1762784779
<< locali >>
rect -220 404 -172 410
rect -220 370 -214 404
rect -180 370 -172 404
rect -220 362 -172 370
rect 770 390 860 396
rect -300 308 -252 312
rect -300 268 -296 308
rect -256 268 -252 308
rect -32 303 16 308
rect -32 302 106 303
rect -32 268 -26 302
rect 8 268 106 302
rect -300 264 -252 268
rect -32 263 106 268
rect -32 260 16 263
rect 770 200 776 390
rect 854 200 860 390
rect 770 194 860 200
rect -220 -66 -172 -60
rect -220 -100 -214 -66
rect -180 -100 -172 -66
rect -220 -108 -172 -100
rect 770 -104 860 -98
rect -32 -167 16 -162
rect -32 -168 106 -167
rect -32 -202 -26 -168
rect 8 -202 106 -168
rect -32 -207 106 -202
rect -32 -210 16 -207
rect 770 -294 776 -104
rect 854 -294 860 -104
rect 770 -300 860 -294
rect -220 -684 -172 -678
rect -220 -718 -214 -684
rect -180 -718 -172 -684
rect -220 -726 -172 -718
rect -310 -788 -242 -776
rect -310 -826 -292 -788
rect -132 -784 -80 -776
rect -132 -818 -122 -784
rect -88 -818 -80 -784
rect -132 -828 -80 -818
rect -32 -785 16 -780
rect -32 -786 154 -785
rect -32 -820 -26 -786
rect 8 -820 154 -786
rect -32 -825 154 -820
rect -32 -828 16 -825
rect -256 -1154 -208 -1148
rect -256 -1188 -250 -1154
rect -216 -1188 -208 -1154
rect -256 -1196 -208 -1188
rect -68 -1255 -20 -1250
rect -68 -1256 70 -1255
rect -176 -1262 -128 -1256
rect -176 -1296 -168 -1262
rect -134 -1296 -128 -1262
rect -176 -1304 -128 -1296
rect -68 -1290 -62 -1256
rect -28 -1290 70 -1256
rect -68 -1295 70 -1290
rect 170 -1295 222 -1255
rect -68 -1298 -20 -1295
rect -130 -1772 -82 -1766
rect -130 -1806 -124 -1772
rect -90 -1806 -82 -1772
rect -130 -1814 -82 -1806
rect -300 -1868 -252 -1864
rect -300 -1908 -296 -1868
rect -256 -1908 -252 -1868
rect -300 -1912 -252 -1908
rect -130 -1870 -82 -1864
rect -130 -1904 -122 -1870
rect -88 -1904 -82 -1870
rect -130 -1912 -82 -1904
rect -14 -1873 34 -1868
rect -14 -1874 124 -1873
rect -14 -1908 -8 -1874
rect 26 -1908 124 -1874
rect -14 -1913 124 -1908
rect 238 -1913 290 -1873
rect -14 -1916 34 -1913
rect -14 -2343 34 -2340
rect -130 -2350 -82 -2344
rect -130 -2384 -122 -2350
rect -88 -2384 -82 -2350
rect -130 -2392 -82 -2384
rect -14 -2348 124 -2343
rect -14 -2382 -8 -2348
rect 26 -2382 124 -2348
rect -14 -2383 124 -2382
rect -14 -2388 34 -2383
rect 306 -2385 358 -2345
rect -130 -2510 -82 -2502
rect -130 -2544 -124 -2510
rect -90 -2544 -82 -2510
rect -130 -2550 -82 -2544
rect -130 -2800 -82 -2794
rect -130 -2834 -124 -2800
rect -90 -2834 -82 -2800
rect -130 -2842 -82 -2834
rect -130 -2958 -82 -2952
rect -130 -2992 -122 -2958
rect -88 -2992 -82 -2958
rect -130 -3000 -82 -2992
rect -14 -2961 34 -2956
rect -14 -2962 124 -2961
rect -14 -2996 -8 -2962
rect 26 -2996 124 -2962
rect -14 -3001 124 -2996
rect 374 -3001 426 -2961
rect -14 -3004 34 -3001
rect 420 -3366 496 -3360
rect -312 -3440 -244 -3432
rect -312 -3474 -296 -3440
rect -262 -3474 -244 -3440
rect -312 -3480 -244 -3474
rect -208 -3436 104 -3432
rect -208 -3476 -196 -3436
rect -84 -3476 104 -3436
rect -208 -3480 -72 -3476
rect 420 -3546 426 -3366
rect 490 -3546 496 -3366
rect 420 -3552 496 -3546
rect -300 -3846 -252 -3842
rect -300 -3886 -296 -3846
rect -256 -3886 -252 -3846
rect -300 -3890 -252 -3886
rect -34 -4056 80 -4044
rect -34 -4096 -28 -4056
rect 12 -4096 80 -4056
rect -34 -4108 80 -4096
rect 34 -4516 86 -4508
rect 34 -4556 40 -4516
rect 80 -4556 86 -4516
rect 34 -4564 86 -4556
rect -166 -5498 -106 -5486
rect -166 -5708 -160 -5498
rect -112 -5708 -106 -5498
rect 162 -5610 230 -5604
rect 162 -5650 176 -5610
rect 216 -5650 230 -5610
rect 162 -5656 230 -5650
rect -166 -5720 -106 -5708
<< viali >>
rect -214 370 -180 404
rect -296 268 -256 308
rect -122 268 -88 302
rect -26 268 8 302
rect 688 264 728 300
rect 776 200 854 390
rect -214 -100 -180 -66
rect -296 -210 -260 -174
rect -122 -206 -88 -172
rect -26 -202 8 -168
rect 688 -204 728 -168
rect 776 -294 854 -104
rect -214 -718 -180 -684
rect -292 -826 -242 -788
rect -122 -818 -88 -784
rect -26 -820 8 -786
rect 688 -824 728 -788
rect 776 -888 842 -698
rect -250 -1188 -216 -1154
rect -168 -1296 -134 -1262
rect -62 -1290 -28 -1256
rect 688 -1292 728 -1256
rect 776 -1382 842 -1192
rect -124 -1806 -90 -1772
rect -296 -1908 -256 -1868
rect -122 -1904 -88 -1870
rect -8 -1908 26 -1874
rect 688 -1912 728 -1876
rect 776 -1976 842 -1786
rect -296 -2386 -260 -2350
rect -122 -2384 -88 -2350
rect -8 -2382 26 -2348
rect 688 -2382 728 -2346
rect 776 -2470 842 -2280
rect -124 -2544 -90 -2510
rect -124 -2834 -90 -2800
rect -292 -2993 -258 -2959
rect -122 -2992 -88 -2958
rect -8 -2996 26 -2962
rect 688 -3000 728 -2964
rect 776 -3064 842 -2874
rect -296 -3474 -262 -3440
rect -196 -3476 -84 -3436
rect 260 -3476 372 -3436
rect 426 -3546 490 -3366
rect -296 -3886 -256 -3846
rect -294 -4082 -260 -4048
rect -124 -4082 -90 -4048
rect -28 -4096 12 -4056
rect 388 -4084 472 -3976
rect 798 -4082 838 -4046
rect -250 -4562 -210 -4522
rect 40 -4556 80 -4516
rect 388 -4632 472 -4524
rect 798 -4562 838 -4526
rect -182 -4682 -142 -4642
rect -296 -5172 -260 -5136
rect -126 -5172 -86 -5132
rect 110 -5170 146 -5134
rect 388 -5172 472 -5064
rect 798 -5170 838 -5134
rect -209 -5265 -169 -5225
rect -250 -5648 -214 -5612
rect -160 -5708 -112 -5498
rect 176 -5650 216 -5610
rect 388 -5720 472 -5612
rect 798 -5650 838 -5614
rect -250 -6258 -214 -6222
rect -160 -6262 -124 -6154
rect 244 -6260 284 -6220
rect 388 -6260 472 -6152
rect 798 -6258 838 -6222
rect 300 -6740 340 -6700
rect 388 -6808 472 -6700
rect 798 -6738 838 -6702
rect 300 -7356 340 -7316
rect 388 -7348 472 -7240
rect 798 -7346 838 -7310
<< metal1 >>
rect -618 634 -324 640
rect -618 550 -612 634
rect -384 550 -324 634
rect -618 544 -324 550
rect -228 404 -164 412
rect -228 370 -214 404
rect -180 400 -164 404
rect -180 372 6 400
rect -180 370 -164 372
rect -228 360 -164 370
rect -22 316 6 372
rect 764 396 866 402
rect -308 262 -302 314
rect -250 262 -244 314
rect -138 260 -132 312
rect -80 260 -74 312
rect -34 310 18 316
rect -40 258 -34 310
rect 18 258 24 310
rect 682 308 734 314
rect -34 252 18 258
rect 682 250 734 256
rect 764 194 770 396
rect 860 194 866 396
rect 764 188 866 194
rect -618 90 -324 96
rect -618 6 -612 90
rect -384 6 -324 90
rect -618 0 -324 6
rect -228 -66 -164 -58
rect -228 -100 -214 -66
rect -180 -70 -164 -66
rect -180 -98 6 -70
rect -180 -100 -164 -98
rect -228 -110 -164 -100
rect -22 -160 6 -98
rect 764 -98 942 -92
rect 764 -104 872 -98
rect 34 -160 86 -154
rect 682 -160 734 -154
rect -308 -174 -170 -168
rect -308 -210 -296 -174
rect -260 -210 -170 -174
rect -308 -216 -170 -210
rect -138 -216 -132 -164
rect -80 -216 -74 -164
rect -40 -168 34 -160
rect -40 -202 -26 -168
rect 8 -202 34 -168
rect -40 -212 34 -202
rect 86 -212 106 -160
rect -222 -260 -170 -216
rect 34 -218 86 -212
rect 682 -218 734 -212
rect 764 -294 776 -104
rect 854 -294 872 -104
rect 764 -300 872 -294
rect 936 -300 942 -98
rect 764 -306 942 -300
rect -222 -318 -170 -312
rect -618 -454 -324 -448
rect -618 -538 -612 -454
rect -384 -538 -324 -454
rect -618 -544 -324 -538
rect -228 -684 -164 -676
rect -228 -718 -214 -684
rect -180 -688 -164 -684
rect -180 -716 6 -688
rect -180 -718 -164 -716
rect -228 -728 -164 -718
rect -304 -788 -230 -782
rect -304 -826 -292 -788
rect -242 -826 -230 -788
rect -304 -832 -230 -826
rect -138 -828 -132 -776
rect -80 -828 -74 -776
rect -22 -778 6 -716
rect 764 -692 854 -686
rect 102 -778 154 -772
rect -40 -786 102 -778
rect -40 -820 -26 -786
rect 8 -820 102 -786
rect -40 -830 102 -820
rect 154 -830 174 -778
rect 682 -780 734 -774
rect -292 -877 -242 -832
rect 102 -836 154 -830
rect 682 -838 734 -832
rect 456 -876 508 -870
rect -292 -927 456 -877
rect 508 -927 533 -877
rect 764 -894 770 -692
rect 848 -894 854 -692
rect 764 -900 854 -894
rect 456 -934 508 -928
rect -618 -998 -324 -992
rect -618 -1082 -612 -998
rect -384 -1082 -324 -998
rect -618 -1088 -324 -1082
rect -264 -1154 -200 -1146
rect -264 -1188 -250 -1154
rect -216 -1158 -200 -1154
rect -216 -1186 -30 -1158
rect -216 -1188 -200 -1186
rect -264 -1198 -200 -1188
rect -58 -1248 -30 -1186
rect 764 -1186 854 -1180
rect 170 -1248 222 -1242
rect -76 -1250 -12 -1248
rect -184 -1262 -118 -1254
rect -184 -1296 -168 -1262
rect -134 -1296 -118 -1262
rect -184 -1306 -118 -1296
rect -76 -1256 170 -1250
rect -76 -1290 -62 -1256
rect -28 -1290 170 -1256
rect -76 -1300 170 -1290
rect 170 -1306 222 -1300
rect 682 -1248 734 -1242
rect 682 -1306 734 -1300
rect -160 -1348 -118 -1306
rect -160 -1354 -80 -1348
rect -160 -1406 -132 -1354
rect 764 -1388 770 -1186
rect 848 -1388 854 -1186
rect 764 -1394 854 -1388
rect -160 -1412 -80 -1406
rect -618 -1542 -324 -1536
rect -618 -1626 -612 -1542
rect -384 -1626 -324 -1542
rect -618 -1632 -324 -1626
rect -138 -1772 -74 -1764
rect -138 -1806 -124 -1772
rect -90 -1776 -74 -1772
rect -90 -1804 24 -1776
rect -90 -1806 -74 -1804
rect -138 -1816 -74 -1806
rect -308 -1914 -302 -1862
rect -250 -1914 -244 -1862
rect -138 -1914 -132 -1862
rect -80 -1914 -74 -1862
rect -4 -1866 24 -1804
rect 764 -1780 854 -1774
rect 238 -1866 290 -1860
rect -22 -1874 238 -1866
rect -22 -1908 -8 -1874
rect 26 -1908 238 -1874
rect -22 -1918 238 -1908
rect 238 -1924 290 -1918
rect 682 -1868 734 -1862
rect 682 -1926 734 -1920
rect 764 -1982 770 -1780
rect 848 -1982 854 -1780
rect 764 -1988 854 -1982
rect -618 -2086 -324 -2080
rect -618 -2170 -612 -2086
rect -384 -2170 -324 -2086
rect -618 -2176 -324 -2170
rect -308 -2230 -170 -2224
rect -308 -2282 -222 -2230
rect -308 -2288 -170 -2282
rect 764 -2274 854 -2268
rect -308 -2342 -244 -2288
rect 306 -2338 358 -2332
rect -314 -2350 -242 -2342
rect -314 -2386 -296 -2350
rect -260 -2386 -242 -2350
rect -314 -2394 -242 -2386
rect -138 -2394 -132 -2342
rect -80 -2394 -74 -2342
rect -22 -2348 306 -2338
rect -22 -2382 -8 -2348
rect 26 -2382 306 -2348
rect -22 -2390 306 -2382
rect -138 -2510 -74 -2500
rect -138 -2544 -124 -2510
rect -90 -2512 -74 -2510
rect -4 -2512 24 -2390
rect 306 -2396 358 -2390
rect 682 -2338 734 -2332
rect 682 -2396 734 -2390
rect 764 -2476 770 -2274
rect 848 -2476 854 -2274
rect 764 -2482 854 -2476
rect -90 -2540 24 -2512
rect -90 -2544 -74 -2540
rect -138 -2552 -74 -2544
rect -618 -2630 -324 -2624
rect -618 -2714 -612 -2630
rect -384 -2714 -324 -2630
rect -618 -2720 -324 -2714
rect -138 -2800 -74 -2792
rect -138 -2834 -124 -2800
rect -90 -2804 -74 -2800
rect -90 -2832 24 -2804
rect -90 -2834 -74 -2832
rect -138 -2844 -74 -2834
rect -298 -2959 -252 -2947
rect -298 -2993 -292 -2959
rect -258 -2993 -252 -2959
rect -298 -3005 -252 -2993
rect -138 -3002 -132 -2950
rect -80 -3002 -74 -2950
rect -4 -2954 24 -2832
rect 764 -2868 854 -2862
rect 374 -2954 426 -2948
rect -22 -2962 374 -2954
rect -22 -2996 -8 -2962
rect 26 -2996 374 -2962
rect -290 -3082 -261 -3005
rect -22 -3006 374 -2996
rect 374 -3012 426 -3006
rect 682 -2956 734 -2950
rect 682 -3014 734 -3008
rect 764 -3070 770 -2868
rect 848 -3070 854 -2868
rect -143 -3082 -137 -3070
rect -290 -3111 -137 -3082
rect -143 -3122 -137 -3111
rect -85 -3082 -79 -3070
rect 451 -3082 457 -3071
rect -85 -3111 457 -3082
rect -85 -3122 -79 -3111
rect 451 -3123 457 -3111
rect 509 -3123 515 -3071
rect 764 -3076 854 -3070
rect -618 -3174 -324 -3168
rect -618 -3258 -612 -3174
rect -384 -3258 -324 -3174
rect -618 -3264 -324 -3258
rect 414 -3366 964 -3360
rect -312 -3440 -250 -3432
rect -312 -3474 -296 -3440
rect -262 -3474 -250 -3440
rect -312 -3480 -250 -3474
rect -222 -3436 386 -3430
rect -222 -3476 -196 -3436
rect -84 -3476 260 -3436
rect 372 -3476 386 -3436
rect -312 -3562 -252 -3480
rect -222 -3482 386 -3476
rect -312 -3622 -98 -3562
rect -38 -3622 -32 -3562
rect 334 -3620 386 -3482
rect 414 -3546 426 -3366
rect 490 -3546 878 -3366
rect 414 -3566 878 -3546
rect 958 -3566 964 -3366
rect 414 -3572 964 -3566
rect 466 -3620 530 -3614
rect 334 -3672 472 -3620
rect 524 -3672 530 -3620
rect 466 -3678 530 -3672
rect -618 -3718 -324 -3712
rect -618 -3802 -612 -3718
rect -384 -3802 -324 -3718
rect -618 -3808 -324 -3802
rect -308 -3892 -302 -3840
rect -250 -3892 -244 -3840
rect -158 -3848 -106 -3842
rect -158 -3966 -106 -3900
rect 376 -3880 964 -3874
rect -1016 -4006 -70 -3966
rect -314 -4048 -300 -4038
rect -1016 -4088 -300 -4048
rect -314 -4090 -300 -4088
rect -248 -4090 -242 -4038
rect -142 -4048 -70 -4006
rect 376 -3976 878 -3880
rect -142 -4082 -124 -4048
rect -90 -4082 -70 -4048
rect -142 -4090 -70 -4082
rect -34 -4050 18 -4044
rect 376 -4084 388 -3976
rect 472 -3998 878 -3976
rect 958 -3998 964 -3880
rect 472 -4004 964 -3998
rect 472 -4084 486 -4004
rect 376 -4090 486 -4084
rect 792 -4038 844 -4032
rect 792 -4096 844 -4090
rect -34 -4108 18 -4102
rect -618 -4262 -324 -4256
rect -618 -4346 -612 -4262
rect -384 -4346 -324 -4262
rect -618 -4352 -324 -4346
rect 34 -4510 86 -4504
rect -262 -4568 -256 -4516
rect -204 -4568 -198 -4516
rect 792 -4518 844 -4512
rect 34 -4568 86 -4562
rect 376 -4524 486 -4518
rect -188 -4636 -136 -4630
rect -188 -4694 -136 -4688
rect 376 -4632 388 -4524
rect 472 -4604 486 -4524
rect 792 -4576 844 -4570
rect 472 -4610 1016 -4604
rect 472 -4632 930 -4610
rect 376 -4728 930 -4632
rect 1010 -4728 1016 -4610
rect 376 -4734 1016 -4728
rect -618 -4806 -324 -4800
rect -618 -4890 -612 -4806
rect -384 -4890 -324 -4806
rect -618 -4896 -324 -4890
rect 376 -4968 964 -4962
rect 376 -5064 878 -4968
rect -132 -5126 -80 -5120
rect -310 -5180 -304 -5128
rect -252 -5180 -246 -5128
rect -132 -5184 -80 -5178
rect 102 -5126 154 -5120
rect 376 -5172 388 -5064
rect 472 -5086 878 -5064
rect 958 -5086 964 -4968
rect 472 -5092 964 -5086
rect 472 -5172 486 -5092
rect 376 -5178 486 -5172
rect 792 -5126 844 -5120
rect 102 -5184 154 -5178
rect 792 -5184 844 -5178
rect -215 -5219 -163 -5213
rect -215 -5277 -163 -5271
rect -618 -5350 -324 -5344
rect -618 -5434 -612 -5350
rect -384 -5434 -324 -5350
rect -618 -5440 -324 -5434
rect -166 -5492 -106 -5486
rect -266 -5612 -200 -5606
rect -266 -5614 -250 -5612
rect -1016 -5648 -250 -5614
rect -214 -5648 -200 -5612
rect -1016 -5654 -200 -5648
rect 162 -5662 170 -5598
rect 222 -5662 230 -5598
rect 792 -5606 844 -5600
rect 376 -5612 486 -5606
rect -166 -5720 -106 -5714
rect 376 -5720 388 -5612
rect 472 -5692 486 -5612
rect 792 -5664 844 -5658
rect 472 -5698 1016 -5692
rect 472 -5720 930 -5698
rect 376 -5816 930 -5720
rect 1010 -5816 1016 -5698
rect 376 -5822 1016 -5816
rect -618 -5894 -324 -5888
rect -618 -5978 -612 -5894
rect -384 -5978 -324 -5894
rect -618 -5984 -324 -5978
rect 376 -6056 988 -6050
rect -166 -6154 -118 -6142
rect -266 -6222 -200 -6216
rect -266 -6224 -250 -6222
rect -1016 -6258 -250 -6224
rect -214 -6258 -200 -6222
rect -1016 -6264 -200 -6258
rect -166 -6262 -160 -6154
rect -124 -6262 -118 -6154
rect 376 -6152 902 -6056
rect -166 -6332 -118 -6262
rect 238 -6214 290 -6208
rect 376 -6260 388 -6152
rect 472 -6174 902 -6152
rect 982 -6174 988 -6056
rect 472 -6180 988 -6174
rect 472 -6260 486 -6180
rect 376 -6266 486 -6260
rect 792 -6214 844 -6208
rect 238 -6272 290 -6266
rect 792 -6272 844 -6266
rect 464 -6332 470 -6330
rect -166 -6380 470 -6332
rect 464 -6382 470 -6380
rect 522 -6382 528 -6330
rect -618 -6438 -324 -6432
rect -618 -6522 -612 -6438
rect -384 -6522 -324 -6438
rect -618 -6528 -324 -6522
rect 294 -6694 346 -6688
rect 792 -6694 844 -6688
rect 294 -6752 346 -6746
rect 376 -6700 486 -6694
rect 376 -6808 388 -6700
rect 472 -6780 486 -6700
rect 792 -6752 844 -6746
rect 472 -6786 1016 -6780
rect 472 -6808 930 -6786
rect 376 -6904 930 -6808
rect 1010 -6904 1016 -6786
rect 376 -6910 1016 -6904
rect -618 -6982 -44 -6976
rect -618 -7066 -612 -6982
rect -384 -7066 -44 -6982
rect -618 -7072 -44 -7066
rect 376 -7144 1090 -7138
rect 376 -7240 1004 -7144
rect 294 -7310 346 -7304
rect 376 -7348 388 -7240
rect 472 -7262 1004 -7240
rect 1084 -7262 1090 -7144
rect 472 -7268 1090 -7262
rect 472 -7348 486 -7268
rect 376 -7354 486 -7348
rect 792 -7302 844 -7296
rect 792 -7360 844 -7354
rect 294 -7368 346 -7362
rect -618 -7526 -44 -7520
rect -618 -7610 -612 -7526
rect -384 -7610 -44 -7526
rect -618 -7616 -44 -7610
<< via1 >>
rect -612 550 -384 634
rect -302 308 -250 314
rect -302 268 -296 308
rect -296 268 -256 308
rect -256 268 -250 308
rect -302 262 -250 268
rect -132 302 -80 312
rect -132 268 -122 302
rect -122 268 -88 302
rect -88 268 -80 302
rect -132 260 -80 268
rect -34 302 18 310
rect -34 268 -26 302
rect -26 268 8 302
rect 8 268 18 302
rect -34 258 18 268
rect 682 300 734 308
rect 682 264 688 300
rect 688 264 728 300
rect 728 264 734 300
rect 682 256 734 264
rect 770 390 860 396
rect 770 200 776 390
rect 776 200 854 390
rect 854 200 860 390
rect 770 194 860 200
rect -612 6 -384 90
rect -132 -172 -80 -164
rect -132 -206 -122 -172
rect -122 -206 -88 -172
rect -88 -206 -80 -172
rect -132 -216 -80 -206
rect 34 -212 86 -160
rect 682 -168 734 -160
rect 682 -204 688 -168
rect 688 -204 728 -168
rect 728 -204 734 -168
rect 682 -212 734 -204
rect -222 -312 -170 -260
rect 872 -300 936 -98
rect -612 -538 -384 -454
rect -132 -784 -80 -776
rect -132 -818 -122 -784
rect -122 -818 -88 -784
rect -88 -818 -80 -784
rect -132 -828 -80 -818
rect 102 -830 154 -778
rect 682 -788 734 -780
rect 682 -824 688 -788
rect 688 -824 728 -788
rect 728 -824 734 -788
rect 682 -832 734 -824
rect 456 -928 508 -876
rect 770 -698 848 -692
rect 770 -888 776 -698
rect 776 -888 842 -698
rect 842 -888 848 -698
rect 770 -894 848 -888
rect -612 -1082 -384 -998
rect 170 -1300 222 -1248
rect 682 -1256 734 -1248
rect 682 -1292 688 -1256
rect 688 -1292 728 -1256
rect 728 -1292 734 -1256
rect 682 -1300 734 -1292
rect -132 -1406 -80 -1354
rect 770 -1192 848 -1186
rect 770 -1382 776 -1192
rect 776 -1382 842 -1192
rect 842 -1382 848 -1192
rect 770 -1388 848 -1382
rect -612 -1626 -384 -1542
rect -302 -1868 -250 -1862
rect -302 -1908 -296 -1868
rect -296 -1908 -256 -1868
rect -256 -1908 -250 -1868
rect -302 -1914 -250 -1908
rect -132 -1870 -80 -1862
rect -132 -1904 -122 -1870
rect -122 -1904 -88 -1870
rect -88 -1904 -80 -1870
rect -132 -1914 -80 -1904
rect 238 -1918 290 -1866
rect 682 -1876 734 -1868
rect 682 -1912 688 -1876
rect 688 -1912 728 -1876
rect 728 -1912 734 -1876
rect 682 -1920 734 -1912
rect 770 -1786 848 -1780
rect 770 -1976 776 -1786
rect 776 -1976 842 -1786
rect 842 -1976 848 -1786
rect 770 -1982 848 -1976
rect -612 -2170 -384 -2086
rect -222 -2282 -170 -2230
rect -132 -2350 -80 -2342
rect -132 -2384 -122 -2350
rect -122 -2384 -88 -2350
rect -88 -2384 -80 -2350
rect -132 -2394 -80 -2384
rect 306 -2390 358 -2338
rect 682 -2346 734 -2338
rect 682 -2382 688 -2346
rect 688 -2382 728 -2346
rect 728 -2382 734 -2346
rect 682 -2390 734 -2382
rect 770 -2280 848 -2274
rect 770 -2470 776 -2280
rect 776 -2470 842 -2280
rect 842 -2470 848 -2280
rect 770 -2476 848 -2470
rect -612 -2714 -384 -2630
rect -132 -2958 -80 -2950
rect -132 -2992 -122 -2958
rect -122 -2992 -88 -2958
rect -88 -2992 -80 -2958
rect -132 -3002 -80 -2992
rect 374 -3006 426 -2954
rect 682 -2964 734 -2956
rect 682 -3000 688 -2964
rect 688 -3000 728 -2964
rect 728 -3000 734 -2964
rect 682 -3008 734 -3000
rect 770 -2874 848 -2868
rect 770 -3064 776 -2874
rect 776 -3064 842 -2874
rect 842 -3064 848 -2874
rect 770 -3070 848 -3064
rect -137 -3122 -85 -3070
rect 457 -3123 509 -3071
rect -612 -3258 -384 -3174
rect -98 -3622 -38 -3562
rect 878 -3566 958 -3366
rect 472 -3672 524 -3620
rect -612 -3802 -384 -3718
rect -302 -3846 -250 -3840
rect -302 -3886 -296 -3846
rect -296 -3886 -256 -3846
rect -256 -3886 -250 -3846
rect -302 -3892 -250 -3886
rect -158 -3900 -106 -3848
rect -300 -4048 -248 -4038
rect -300 -4082 -294 -4048
rect -294 -4082 -260 -4048
rect -260 -4082 -248 -4048
rect -300 -4090 -248 -4082
rect -34 -4056 18 -4050
rect -34 -4096 -28 -4056
rect -28 -4096 12 -4056
rect 12 -4096 18 -4056
rect 878 -3998 958 -3880
rect 792 -4046 844 -4038
rect 792 -4082 798 -4046
rect 798 -4082 838 -4046
rect 838 -4082 844 -4046
rect 792 -4090 844 -4082
rect -34 -4102 18 -4096
rect -612 -4346 -384 -4262
rect 34 -4516 86 -4510
rect -256 -4522 -204 -4516
rect -256 -4562 -250 -4522
rect -250 -4562 -210 -4522
rect -210 -4562 -204 -4522
rect -256 -4568 -204 -4562
rect 34 -4556 40 -4516
rect 40 -4556 80 -4516
rect 80 -4556 86 -4516
rect 34 -4562 86 -4556
rect -188 -4642 -136 -4636
rect -188 -4682 -182 -4642
rect -182 -4682 -142 -4642
rect -142 -4682 -136 -4642
rect -188 -4688 -136 -4682
rect 792 -4526 844 -4518
rect 792 -4562 798 -4526
rect 798 -4562 838 -4526
rect 838 -4562 844 -4526
rect 792 -4570 844 -4562
rect 930 -4728 1010 -4610
rect -612 -4890 -384 -4806
rect -304 -5136 -252 -5128
rect -304 -5172 -296 -5136
rect -296 -5172 -260 -5136
rect -260 -5172 -252 -5136
rect -304 -5180 -252 -5172
rect -132 -5132 -80 -5126
rect -132 -5172 -126 -5132
rect -126 -5172 -86 -5132
rect -86 -5172 -80 -5132
rect -132 -5178 -80 -5172
rect 102 -5134 154 -5126
rect 102 -5170 110 -5134
rect 110 -5170 146 -5134
rect 146 -5170 154 -5134
rect 102 -5178 154 -5170
rect 878 -5086 958 -4968
rect 792 -5134 844 -5126
rect 792 -5170 798 -5134
rect 798 -5170 838 -5134
rect 838 -5170 844 -5134
rect 792 -5178 844 -5170
rect -215 -5225 -163 -5219
rect -215 -5265 -209 -5225
rect -209 -5265 -169 -5225
rect -169 -5265 -163 -5225
rect -215 -5271 -163 -5265
rect -612 -5434 -384 -5350
rect -166 -5498 -106 -5492
rect -166 -5708 -160 -5498
rect -160 -5708 -112 -5498
rect -112 -5708 -106 -5498
rect 170 -5610 222 -5598
rect 170 -5650 176 -5610
rect 176 -5650 216 -5610
rect 216 -5650 222 -5610
rect 170 -5662 222 -5650
rect -166 -5714 -106 -5708
rect 792 -5614 844 -5606
rect 792 -5650 798 -5614
rect 798 -5650 838 -5614
rect 838 -5650 844 -5614
rect 792 -5658 844 -5650
rect 930 -5816 1010 -5698
rect -612 -5978 -384 -5894
rect 238 -6220 290 -6214
rect 238 -6260 244 -6220
rect 244 -6260 284 -6220
rect 284 -6260 290 -6220
rect 238 -6266 290 -6260
rect 902 -6174 982 -6056
rect 792 -6222 844 -6214
rect 792 -6258 798 -6222
rect 798 -6258 838 -6222
rect 838 -6258 844 -6222
rect 792 -6266 844 -6258
rect 470 -6382 522 -6330
rect -612 -6522 -384 -6438
rect 294 -6700 346 -6694
rect 294 -6740 300 -6700
rect 300 -6740 340 -6700
rect 340 -6740 346 -6700
rect 294 -6746 346 -6740
rect 792 -6702 844 -6694
rect 792 -6738 798 -6702
rect 798 -6738 838 -6702
rect 838 -6738 844 -6702
rect 792 -6746 844 -6738
rect 930 -6904 1010 -6786
rect -612 -7066 -384 -6982
rect 294 -7316 346 -7310
rect 294 -7356 300 -7316
rect 300 -7356 340 -7316
rect 340 -7356 346 -7316
rect 1004 -7262 1084 -7144
rect 792 -7310 844 -7302
rect 792 -7346 798 -7310
rect 798 -7346 838 -7310
rect 838 -7346 844 -7310
rect 792 -7354 844 -7346
rect 294 -7362 346 -7356
rect -612 -7610 -384 -7526
<< metal2 >>
rect -618 634 -378 640
rect -618 550 -612 634
rect -384 550 -378 634
rect -618 544 -378 550
rect 764 396 1010 402
rect -308 262 -302 314
rect -250 262 -244 314
rect -132 312 -80 318
rect -618 90 -378 96
rect -618 6 -612 90
rect -384 6 -378 90
rect -618 0 -378 6
rect -618 -454 -378 -448
rect -618 -538 -612 -454
rect -384 -538 -378 -454
rect -618 -544 -378 -538
rect -618 -998 -378 -992
rect -618 -1082 -612 -998
rect -384 -1082 -378 -998
rect -618 -1088 -378 -1082
rect -618 -1542 -378 -1536
rect -618 -1626 -612 -1542
rect -384 -1626 -378 -1542
rect -618 -1632 -378 -1626
rect -290 -1862 -262 262
rect -132 -164 -80 260
rect -34 310 18 316
rect -34 252 18 258
rect 682 308 734 314
rect -222 -260 -170 -254
rect -222 -318 -170 -312
rect -308 -1914 -302 -1862
rect -250 -1914 -244 -1862
rect -618 -2086 -378 -2080
rect -618 -2170 -612 -2086
rect -384 -2170 -378 -2086
rect -618 -2176 -378 -2170
rect -618 -2630 -378 -2624
rect -618 -2714 -612 -2630
rect -384 -2714 -378 -2630
rect -618 -2720 -378 -2714
rect -618 -3174 -378 -3168
rect -618 -3258 -612 -3174
rect -384 -3258 -378 -3174
rect -618 -3264 -378 -3258
rect -618 -3718 -378 -3712
rect -618 -3802 -612 -3718
rect -384 -3802 -378 -3718
rect -618 -3808 -378 -3802
rect -290 -3840 -262 -1914
rect -210 -2224 -182 -318
rect -132 -776 -80 -216
rect -132 -1354 -80 -828
rect -132 -1862 -80 -1406
rect -222 -2230 -170 -2224
rect -222 -2288 -170 -2282
rect -308 -3892 -302 -3840
rect -250 -3892 -244 -3840
rect -306 -4090 -300 -4038
rect -248 -4090 -242 -4038
rect -618 -4262 -378 -4256
rect -618 -4346 -612 -4262
rect -384 -4346 -378 -4262
rect -618 -4352 -378 -4346
rect -288 -4516 -260 -4090
rect -214 -4416 -186 -2288
rect -132 -2342 -80 -1914
rect -132 -2856 -80 -2394
rect -144 -2866 -68 -2856
rect -144 -2922 -134 -2866
rect -78 -2922 -68 -2866
rect -144 -2932 -68 -2922
rect -132 -2950 -80 -2932
rect -132 -3008 -80 -3002
rect -137 -3070 -85 -3064
rect -137 -3128 -85 -3122
rect -125 -3494 -96 -3128
rect -154 -3522 -96 -3494
rect -22 -3494 6 252
rect 34 -160 86 -154
rect 34 -218 86 -212
rect 682 -160 734 256
rect 764 194 770 396
rect 860 194 1010 396
rect 764 188 1010 194
rect -22 -3522 18 -3494
rect -154 -3676 -126 -3522
rect -98 -3562 -38 -3550
rect -98 -3642 -38 -3630
rect -10 -3676 18 -3522
rect -154 -3704 -50 -3676
rect -158 -3848 -106 -3842
rect -158 -3906 -106 -3900
rect -146 -4214 -118 -3906
rect -78 -3982 -50 -3704
rect -90 -4008 -50 -3982
rect -22 -3704 18 -3676
rect -90 -4137 -62 -4008
rect -22 -4044 6 -3704
rect -34 -4050 18 -4044
rect -34 -4108 18 -4102
rect -90 -4166 -12 -4137
rect -146 -4242 -80 -4214
rect -214 -4444 -142 -4416
rect -288 -4568 -256 -4516
rect -204 -4568 -198 -4516
rect -618 -4806 -378 -4800
rect -618 -4890 -612 -4806
rect -384 -4890 -378 -4806
rect -618 -4896 -378 -4890
rect -288 -5128 -260 -4568
rect -170 -4630 -142 -4444
rect -188 -4636 -136 -4630
rect -188 -4694 -136 -4688
rect -108 -5120 -80 -4242
rect -132 -5126 -80 -5120
rect -310 -5180 -304 -5128
rect -252 -5180 -246 -5128
rect -132 -5184 -80 -5178
rect -221 -5271 -215 -5219
rect -163 -5231 -157 -5219
rect -41 -5231 -12 -4166
rect 46 -4504 74 -218
rect 102 -778 154 -772
rect 102 -836 154 -830
rect 682 -780 734 -212
rect 866 -98 942 -92
rect 866 -300 872 -98
rect 936 -300 942 -98
rect 866 -306 942 -300
rect 894 -408 942 -306
rect 970 -284 1010 188
rect 970 -324 1090 -284
rect 894 -448 1010 -408
rect 34 -4510 86 -4504
rect 34 -4568 86 -4562
rect 114 -5120 142 -836
rect 450 -928 456 -876
rect 508 -928 514 -876
rect 170 -1248 222 -1242
rect 170 -1306 222 -1300
rect 102 -5126 154 -5120
rect 102 -5184 154 -5178
rect -163 -5260 -12 -5231
rect -163 -5271 -157 -5260
rect -618 -5350 -378 -5344
rect -618 -5434 -612 -5350
rect -384 -5434 -378 -5350
rect -618 -5440 -378 -5434
rect -166 -5492 -106 -5486
rect 182 -5592 210 -1306
rect 238 -1866 290 -1860
rect 238 -1924 290 -1918
rect 170 -5598 222 -5592
rect 170 -5668 222 -5662
rect -166 -5720 -106 -5714
rect -618 -5894 -378 -5888
rect -618 -5978 -612 -5894
rect -384 -5978 -378 -5894
rect -618 -5984 -378 -5978
rect 250 -6208 278 -1924
rect 306 -2338 358 -2332
rect 306 -2396 358 -2390
rect 238 -6214 290 -6208
rect 238 -6272 290 -6266
rect -618 -6438 -378 -6432
rect -618 -6522 -612 -6438
rect -384 -6522 -378 -6438
rect -618 -6528 -378 -6522
rect 318 -6688 346 -2396
rect 374 -2954 426 -2948
rect 374 -3012 426 -3006
rect 294 -6694 346 -6688
rect 294 -6752 346 -6746
rect -618 -6982 -378 -6976
rect -618 -7066 -612 -6982
rect -384 -7066 -378 -6982
rect -618 -7072 -378 -7066
rect 294 -7308 346 -7304
rect 386 -7308 414 -3012
rect 468 -3065 497 -928
rect 682 -1248 734 -832
rect 764 -692 854 -686
rect 764 -894 770 -692
rect 848 -860 854 -692
rect 970 -748 1010 -448
rect 970 -788 1090 -748
rect 848 -894 1010 -860
rect 764 -900 1010 -894
rect 682 -1868 734 -1300
rect 764 -1186 854 -1180
rect 764 -1388 770 -1186
rect 848 -1354 854 -1186
rect 970 -1212 1010 -900
rect 970 -1252 1090 -1212
rect 848 -1388 1010 -1354
rect 764 -1394 1010 -1388
rect 970 -1676 1010 -1394
rect 970 -1716 1090 -1676
rect 682 -2338 734 -1920
rect 764 -1780 854 -1774
rect 764 -1982 770 -1780
rect 848 -1948 854 -1780
rect 848 -1982 1010 -1948
rect 764 -1988 1010 -1982
rect 970 -2140 1010 -1988
rect 970 -2180 1090 -2140
rect 682 -2956 734 -2390
rect 764 -2274 854 -2268
rect 764 -2476 770 -2274
rect 848 -2442 854 -2274
rect 848 -2476 1010 -2442
rect 764 -2482 1010 -2476
rect 970 -2604 1010 -2482
rect 970 -2644 1090 -2604
rect 457 -3071 509 -3065
rect 457 -3129 509 -3123
rect 466 -3620 530 -3614
rect 682 -3620 734 -3008
rect 764 -2868 854 -2862
rect 764 -3070 770 -2868
rect 848 -3068 854 -2868
rect 848 -3070 1090 -3068
rect 764 -3108 1090 -3070
rect 872 -3366 964 -3360
rect 872 -3566 878 -3366
rect 958 -3532 964 -3366
rect 958 -3566 1090 -3532
rect 872 -3572 1090 -3566
rect 466 -3672 472 -3620
rect 524 -3672 844 -3620
rect 466 -3678 530 -3672
rect 456 -3906 532 -3896
rect 456 -3962 466 -3906
rect 522 -3962 532 -3906
rect 456 -3972 532 -3962
rect 472 -6324 520 -3972
rect 792 -4038 844 -3672
rect 872 -3880 1004 -3874
rect 872 -3998 878 -3880
rect 958 -3996 1004 -3880
rect 958 -3998 1090 -3996
rect 872 -4004 1090 -3998
rect 964 -4036 1090 -4004
rect 792 -4518 844 -4090
rect 792 -5126 844 -4570
rect 970 -4500 1090 -4460
rect 970 -4604 1016 -4500
rect 924 -4610 1016 -4604
rect 924 -4728 930 -4610
rect 1010 -4728 1016 -4610
rect 924 -4734 1016 -4728
rect 964 -4962 1090 -4924
rect 872 -4964 1090 -4962
rect 872 -4968 1004 -4964
rect 872 -5086 878 -4968
rect 958 -5086 1004 -4968
rect 872 -5092 1004 -5086
rect 792 -5606 844 -5178
rect 792 -6214 844 -5658
rect 970 -5428 1090 -5388
rect 970 -5692 1016 -5428
rect 924 -5698 1016 -5692
rect 924 -5816 930 -5698
rect 1010 -5816 1016 -5698
rect 924 -5822 1016 -5816
rect 942 -5892 1090 -5852
rect 942 -6050 988 -5892
rect 896 -6056 988 -6050
rect 896 -6174 902 -6056
rect 982 -6174 988 -6056
rect 896 -6180 988 -6174
rect 470 -6330 522 -6324
rect 470 -6388 522 -6382
rect 294 -7310 414 -7308
rect 346 -7362 414 -7310
rect 792 -6694 844 -6266
rect 792 -7302 844 -6746
rect 970 -6356 1090 -6316
rect 970 -6780 1016 -6356
rect 924 -6786 1016 -6780
rect 924 -6904 930 -6786
rect 1010 -6904 1016 -6786
rect 924 -6910 1016 -6904
rect 1044 -7138 1090 -6780
rect 998 -7144 1090 -7138
rect 998 -7262 1004 -7144
rect 1084 -7262 1090 -7144
rect 998 -7268 1090 -7262
rect 792 -7360 844 -7354
rect 294 -7364 414 -7362
rect 294 -7368 346 -7364
rect -618 -7526 -378 -7520
rect -618 -7610 -612 -7526
rect -384 -7610 -378 -7526
rect -618 -7616 -378 -7610
<< via2 >>
rect -608 554 -390 630
rect -608 -534 -390 -458
rect -608 -1622 -390 -1546
rect -608 -2166 -390 -2090
rect -608 -2710 -390 -2634
rect -608 -3254 -390 -3178
rect -608 -3798 -390 -3722
rect -608 -4342 -390 -4266
rect -134 -2922 -78 -2866
rect -98 -3622 -38 -3562
rect -98 -3630 -38 -3622
rect -608 -4886 -390 -4810
rect -608 -5430 -390 -5354
rect -164 -5552 -108 -5496
rect -608 -5974 -390 -5898
rect -608 -6518 -390 -6442
rect -608 -7062 -390 -6986
rect 466 -3962 522 -3906
rect -608 -7606 -390 -7530
<< metal3 >>
rect -918 634 -378 640
rect -918 550 -912 634
rect -684 630 -378 634
rect -684 554 -608 630
rect -390 554 -378 630
rect -684 550 -378 554
rect -918 544 -378 550
rect -618 90 -378 96
rect -618 6 -612 90
rect -384 6 -378 90
rect -618 0 -378 6
rect -918 -454 -378 -448
rect -918 -538 -912 -454
rect -684 -458 -378 -454
rect -684 -534 -608 -458
rect -390 -534 -378 -458
rect -684 -538 -378 -534
rect -918 -544 -378 -538
rect -618 -998 -378 -992
rect -618 -1082 -612 -998
rect -384 -1082 -378 -998
rect -618 -1088 -378 -1082
rect -918 -1542 -378 -1536
rect -918 -1626 -912 -1542
rect -684 -1546 -378 -1542
rect -684 -1622 -608 -1546
rect -390 -1622 -378 -1546
rect -684 -1626 -378 -1622
rect -918 -1632 -378 -1626
rect -618 -2086 -378 -2080
rect -618 -2170 -612 -2086
rect -384 -2170 -378 -2086
rect -618 -2176 -378 -2170
rect -918 -2630 -378 -2624
rect -918 -2714 -912 -2630
rect -684 -2634 -378 -2630
rect -684 -2710 -608 -2634
rect -390 -2710 -378 -2634
rect -684 -2714 -378 -2710
rect -918 -2720 -378 -2714
rect -139 -2864 -73 -2861
rect -139 -2866 664 -2864
rect -139 -2922 -134 -2866
rect -78 -2922 664 -2866
rect -139 -2924 664 -2922
rect -139 -2927 -73 -2924
rect -618 -3174 -378 -3168
rect -618 -3258 -612 -3174
rect -384 -3258 -378 -3174
rect -618 -3264 -378 -3258
rect -104 -3562 -32 -3536
rect -104 -3630 -98 -3562
rect -38 -3630 -32 -3562
rect -104 -3658 -32 -3630
rect -918 -3718 -378 -3712
rect -918 -3802 -912 -3718
rect -684 -3722 -378 -3718
rect -684 -3798 -608 -3722
rect -390 -3798 -378 -3722
rect -684 -3802 -378 -3798
rect -918 -3808 -378 -3802
rect -92 -3904 -32 -3658
rect 461 -3904 527 -3901
rect -92 -3906 527 -3904
rect -92 -3962 466 -3906
rect 522 -3962 527 -3906
rect -92 -3964 527 -3962
rect 461 -3967 527 -3964
rect -618 -4262 -378 -4256
rect -618 -4346 -612 -4262
rect -384 -4346 -378 -4262
rect -618 -4352 -378 -4346
rect -918 -4806 -378 -4800
rect -918 -4890 -912 -4806
rect -684 -4810 -378 -4806
rect -684 -4886 -608 -4810
rect -390 -4886 -378 -4810
rect -684 -4890 -378 -4886
rect -918 -4896 -378 -4890
rect -618 -5350 -378 -5344
rect -618 -5434 -612 -5350
rect -384 -5434 -378 -5350
rect -618 -5440 -378 -5434
rect -169 -5494 -103 -5491
rect 604 -5494 664 -2924
rect -169 -5496 664 -5494
rect -169 -5552 -164 -5496
rect -108 -5552 664 -5496
rect -169 -5554 664 -5552
rect -169 -5557 -103 -5554
rect -918 -5894 -378 -5888
rect -918 -5978 -912 -5894
rect -684 -5898 -378 -5894
rect -684 -5974 -608 -5898
rect -390 -5974 -378 -5898
rect -684 -5978 -378 -5974
rect -918 -5984 -378 -5978
rect -618 -6438 -378 -6432
rect -618 -6522 -612 -6438
rect -384 -6522 -378 -6438
rect -618 -6528 -378 -6522
rect -918 -6982 -378 -6976
rect -918 -7066 -912 -6982
rect -684 -6986 -378 -6982
rect -684 -7062 -608 -6986
rect -390 -7062 -378 -6986
rect -684 -7066 -378 -7062
rect -918 -7072 -378 -7066
rect -618 -7526 -378 -7520
rect -618 -7610 -612 -7526
rect -384 -7610 -378 -7526
rect -618 -7616 -378 -7610
<< via3 >>
rect -912 550 -684 634
rect -612 6 -384 90
rect -912 -538 -684 -454
rect -612 -1082 -384 -998
rect -912 -1626 -684 -1542
rect -612 -2090 -384 -2086
rect -612 -2166 -608 -2090
rect -608 -2166 -390 -2090
rect -390 -2166 -384 -2090
rect -612 -2170 -384 -2166
rect -912 -2714 -684 -2630
rect -612 -3178 -384 -3174
rect -612 -3254 -608 -3178
rect -608 -3254 -390 -3178
rect -390 -3254 -384 -3178
rect -612 -3258 -384 -3254
rect -912 -3802 -684 -3718
rect -612 -4266 -384 -4262
rect -612 -4342 -608 -4266
rect -608 -4342 -390 -4266
rect -390 -4342 -384 -4266
rect -612 -4346 -384 -4342
rect -912 -4890 -684 -4806
rect -612 -5354 -384 -5350
rect -612 -5430 -608 -5354
rect -608 -5430 -390 -5354
rect -390 -5430 -384 -5354
rect -612 -5434 -384 -5430
rect -912 -5978 -684 -5894
rect -612 -6442 -384 -6438
rect -612 -6518 -608 -6442
rect -608 -6518 -390 -6442
rect -390 -6518 -384 -6442
rect -612 -6522 -384 -6518
rect -912 -7066 -684 -6982
rect -612 -7530 -384 -7526
rect -612 -7606 -608 -7530
rect -608 -7606 -390 -7530
rect -390 -7606 -384 -7530
rect -612 -7610 -384 -7606
<< metal4 >>
rect -918 634 -678 640
rect -918 550 -912 634
rect -684 550 -678 634
rect -918 -454 -678 550
rect -918 -538 -912 -454
rect -684 -538 -678 -454
rect -918 -1542 -678 -538
rect -918 -1626 -912 -1542
rect -684 -1626 -678 -1542
rect -918 -2630 -678 -1626
rect -918 -2714 -912 -2630
rect -684 -2714 -678 -2630
rect -918 -3718 -678 -2714
rect -918 -3802 -912 -3718
rect -684 -3802 -678 -3718
rect -918 -4806 -678 -3802
rect -918 -4890 -912 -4806
rect -684 -4890 -678 -4806
rect -918 -5894 -678 -4890
rect -918 -5978 -912 -5894
rect -684 -5978 -678 -5894
rect -918 -6982 -678 -5978
rect -918 -7066 -912 -6982
rect -684 -7066 -678 -6982
rect -918 -7616 -678 -7066
rect -618 90 -378 640
rect -618 6 -612 90
rect -384 6 -378 90
rect -618 -998 -378 6
rect -618 -1082 -612 -998
rect -384 -1082 -378 -998
rect -618 -2086 -378 -1082
rect -618 -2170 -612 -2086
rect -384 -2170 -378 -2086
rect -618 -3174 -378 -2170
rect -618 -3258 -612 -3174
rect -384 -3258 -378 -3174
rect -618 -4262 -378 -3258
rect -618 -4346 -612 -4262
rect -384 -4346 -378 -4262
rect -618 -5350 -378 -4346
rect -618 -5434 -612 -5350
rect -384 -5434 -378 -5350
rect -618 -6438 -378 -5434
rect -618 -6522 -612 -6438
rect -384 -6522 -378 -6438
rect -618 -7526 -378 -6522
rect -618 -7610 -612 -7526
rect -384 -7610 -378 -7526
rect -618 -7616 -378 -7610
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 -54 0 -1 -3216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1762784779
transform 1 0 -54 0 1 -4304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1762784779
transform 1 0 -54 0 -1 -4304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1762784779
transform 1 0 -54 0 1 -5392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1762784779
transform 1 0 -54 0 -1 -5392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1762784779
transform 1 0 -54 0 1 -6480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1762784779
transform 1 0 -54 0 -1 -6480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1762784779
transform 1 0 -54 0 1 -7568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn0
timestamp 1762784779
transform 1 0 -54 0 1 48
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn1
timestamp 1762784779
transform 1 0 -54 0 -1 48
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn2
timestamp 1762784779
transform 1 0 -54 0 1 -1040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn3
timestamp 1762784779
transform 1 0 -54 0 -1 -1040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn4
timestamp 1762784779
transform 1 0 -54 0 1 -2128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn5
timestamp 1762784779
transform 1 0 -54 0 -1 -2128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn6
timestamp 1762784779
transform 1 0 -54 0 1 -3216
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  XOTn0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 38 0 1 48
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn1
timestamp 1762784779
transform 1 0 38 0 -1 48
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn2
timestamp 1762784779
transform 1 0 38 0 1 -1040
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn3
timestamp 1762784779
transform 1 0 38 0 -1 -1040
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn4
timestamp 1762784779
transform 1 0 38 0 1 -2128
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn5
timestamp 1762784779
transform 1 0 38 0 -1 -2128
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn6
timestamp 1762784779
transform 1 0 38 0 1 -3216
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  XOTn7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 38 0 -1 -3216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  XOTn8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 866 0 1 -4304
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn9
timestamp 1762784779
transform -1 0 866 0 -1 -4304
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn10
timestamp 1762784779
transform -1 0 866 0 1 -5392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn11
timestamp 1762784779
transform -1 0 866 0 -1 -5392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn12
timestamp 1762784779
transform -1 0 866 0 1 -6480
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn13
timestamp 1762784779
transform -1 0 866 0 -1 -6480
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn14
timestamp 1762784779
transform -1 0 866 0 1 -7568
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  XTA1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 -330 0 1 -4304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  XTA2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 -330 0 -1 -4304
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  XTA3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 -330 0 1 -5392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  XTAN
timestamp 1762784779
transform 1 0 -330 0 -1 -5392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  XTAN2
timestamp 1762784779
transform 1 0 -330 0 1 -6480
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  XTB1
timestamp 1762784779
transform -1 0 -54 0 1 48
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  XTB2
timestamp 1762784779
transform -1 0 -54 0 -1 48
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  XTB3
timestamp 1762784779
transform -1 0 -54 0 1 -1040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  XTB4
timestamp 1762784779
transform -1 0 -54 0 -1 -1040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  XTB5
timestamp 1762784779
transform -1 0 -54 0 1 -2128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  XTB6
timestamp 1762784779
transform -1 0 -54 0 -1 -2128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  XTB7
timestamp 1762784779
transform -1 0 -54 0 1 -3216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  XTBN $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 -330 0 -1 -3216
box -38 -48 314 592
<< labels >>
flabel metal2 1050 -324 1090 -284 0 FreeSans 80 0 0 0 Tn[0]
port 1000 nsew
flabel metal2 1050 -788 1090 -748 0 FreeSans 80 0 0 0 Tn[1]
port 1001 nsew
flabel metal2 1050 -1252 1090 -1212 0 FreeSans 80 0 0 0 Tn[2]
port 1002 nsew
flabel metal2 1050 -1716 1090 -1676 0 FreeSans 80 0 0 0 Tn[3]
port 1003 nsew
flabel metal2 1050 -2180 1090 -2140 0 FreeSans 80 0 0 0 Tn[4]
port 1004 nsew
flabel metal2 1050 -2644 1090 -2604 0 FreeSans 80 0 0 0 Tn[5]
port 1005 nsew
flabel metal2 1050 -3108 1090 -3068 0 FreeSans 80 0 0 0 Tn[6]
port 1006 nsew
flabel metal2 1050 -3572 1090 -3532 0 FreeSans 80 0 0 0 Tn[7]
port 1007 nsew
flabel metal2 1050 -4036 1090 -3996 0 FreeSans 80 0 0 0 Tn[8]
port 1008 nsew
flabel metal2 1050 -4500 1090 -4460 0 FreeSans 80 0 0 0 Tn[9]
port 1009 nsew
flabel metal2 1050 -4964 1090 -4924 0 FreeSans 80 0 0 0 Tn[10]
port 1010 nsew
flabel metal2 1050 -5428 1090 -5388 0 FreeSans 80 0 0 0 Tn[11]
port 1011 nsew
flabel metal2 1050 -5892 1090 -5852 0 FreeSans 80 0 0 0 Tn[12]
port 1012 nsew
flabel metal2 1050 -6356 1090 -6316 0 FreeSans 80 0 0 0 Tn[13]
port 1013 nsew
flabel metal2 1050 -6820 1090 -6780 0 FreeSans 80 0 0 0 Tn[14]
port 1014 nsew
flabel metal1 -1016 -4006 -976 -3966 0 FreeSans 80 0 0 0 d[0]
port 1101 nsew
flabel metal1 -1016 -4088 -976 -4048 0 FreeSans 80 0 0 0 d[1]
port 1102 nsew
flabel metal1 -1016 -5654 -976 -5614 0 FreeSans 80 0 0 0 d[2]
port 1103 nsew
flabel metal1 -1016 -6264 -976 -6224 0 FreeSans 80 0 0 0 d[3]
port 1104 nsew
flabel metal4 -918 -7616 -678 640 0 FreeSans 1600 90 0 0 VPWR
port 90 nsew
flabel metal4 -618 -7616 -378 640 0 FreeSans 1600 90 0 0 VGND
port 91 nsew
<< end >>
