magic
tech sky130A
magscale 1 2
timestamp 1758175872
<< metal1 >>
rect 10676 38319 10756 38324
rect 6845 38311 10756 38319
rect 6845 38259 10691 38311
rect 10743 38259 10756 38311
rect 6845 38249 10756 38259
rect 6860 37812 6900 38249
rect 10676 38244 10756 38249
rect 7450 38167 10756 38180
rect 7450 38115 10691 38167
rect 10743 38115 10756 38167
rect 7450 38100 10756 38115
rect 7470 37808 7510 38100
rect 10676 38029 10756 38038
rect 9026 38025 10756 38029
rect 9026 37973 10691 38025
rect 10743 37973 10756 38025
rect 9026 37968 10756 37973
rect 9036 37812 9076 37968
rect 10676 37958 10756 37968
rect 10676 37889 10756 37898
rect 9108 37885 10756 37889
rect 9108 37833 10691 37885
rect 10743 37833 10756 37885
rect 9108 37828 10756 37833
rect 9118 37812 9158 37828
rect 10676 37818 10756 37828
rect 18744 30729 18824 30734
rect 18734 30721 18824 30729
rect 18734 30669 18759 30721
rect 18811 30669 18824 30721
rect 18734 30659 18824 30669
rect 18744 30654 18824 30659
rect 18734 30577 18824 30590
rect 18734 30525 18759 30577
rect 18811 30525 18824 30577
rect 18734 30510 18824 30525
rect 18744 29039 18824 29048
rect 18734 29035 18824 29039
rect 18734 28983 18759 29035
rect 18811 28983 18824 29035
rect 18734 28978 18824 28983
rect 18744 28968 18824 28978
rect 18744 28487 18824 28496
rect 18734 28483 18824 28487
rect 18734 28431 18759 28483
rect 18811 28431 18824 28483
rect 18734 28426 18824 28431
rect 18744 28416 18824 28426
rect 10676 25605 10756 25610
rect 6845 25597 10756 25605
rect 6845 25545 10691 25597
rect 10743 25545 10756 25597
rect 6845 25535 10756 25545
rect 6860 25098 6900 25535
rect 10676 25530 10756 25535
rect 7450 25453 10756 25466
rect 7450 25401 10691 25453
rect 10743 25401 10756 25453
rect 7450 25386 10756 25401
rect 7470 25094 7510 25386
rect 10676 25315 10756 25324
rect 9026 25311 10756 25315
rect 9026 25259 10691 25311
rect 10743 25259 10756 25311
rect 9026 25254 10756 25259
rect 9036 25098 9076 25254
rect 10676 25244 10756 25254
rect 10676 25175 10756 25184
rect 9108 25171 10756 25175
rect 9108 25119 10691 25171
rect 10743 25119 10756 25171
rect 9108 25114 10756 25119
rect 9118 25098 9158 25114
rect 10676 25104 10756 25114
rect 18744 18015 18824 18020
rect 18734 18007 18824 18015
rect 18734 17955 18759 18007
rect 18811 17955 18824 18007
rect 18734 17945 18824 17955
rect 18744 17940 18824 17945
rect 18734 17863 18824 17876
rect 18734 17811 18759 17863
rect 18811 17811 18824 17863
rect 18734 17796 18824 17811
rect 18744 16325 18824 16334
rect 18734 16321 18824 16325
rect 18734 16269 18759 16321
rect 18811 16269 18824 16321
rect 18734 16264 18824 16269
rect 18744 16254 18824 16264
rect 18744 15773 18824 15782
rect 18734 15769 18824 15773
rect 18734 15717 18759 15769
rect 18811 15717 18824 15769
rect 18734 15712 18824 15717
rect 18744 15702 18824 15712
rect 10676 12891 10756 12896
rect 6845 12883 10756 12891
rect 6845 12831 10691 12883
rect 10743 12831 10756 12883
rect 6845 12821 10756 12831
rect 6860 12384 6900 12821
rect 10676 12816 10756 12821
rect 7450 12739 10756 12752
rect 7450 12687 10691 12739
rect 10743 12687 10756 12739
rect 7450 12672 10756 12687
rect 7470 12380 7510 12672
rect 10676 12601 10756 12610
rect 9026 12597 10756 12601
rect 9026 12545 10691 12597
rect 10743 12545 10756 12597
rect 9026 12540 10756 12545
rect 9036 12384 9076 12540
rect 10676 12530 10756 12540
rect 10676 12461 10756 12470
rect 9108 12457 10756 12461
rect 9108 12405 10691 12457
rect 10743 12405 10756 12457
rect 9108 12400 10756 12405
rect 9118 12384 9158 12400
rect 10676 12390 10756 12400
rect 18744 5301 18824 5306
rect 18734 5293 18824 5301
rect 18734 5241 18759 5293
rect 18811 5241 18824 5293
rect 18734 5231 18824 5241
rect 18744 5226 18824 5231
rect 18734 5149 18824 5162
rect 18734 5097 18759 5149
rect 18811 5097 18824 5149
rect 18734 5082 18824 5097
rect 18744 3611 18824 3620
rect 18734 3607 18824 3611
rect 18734 3555 18759 3607
rect 18811 3555 18824 3607
rect 18734 3550 18824 3555
rect 18744 3540 18824 3550
rect 18744 3059 18824 3068
rect 18734 3055 18824 3059
rect 18734 3003 18759 3055
rect 18811 3003 18824 3055
rect 18734 2998 18824 3003
rect 18744 2988 18824 2998
<< via1 >>
rect 10691 38259 10743 38311
rect 10691 38115 10743 38167
rect 10691 37973 10743 38025
rect 10691 37833 10743 37885
rect 18759 30669 18811 30721
rect 18759 30525 18811 30577
rect 18759 28983 18811 29035
rect 18759 28431 18811 28483
rect 10691 25545 10743 25597
rect 10691 25401 10743 25453
rect 10691 25259 10743 25311
rect 10691 25119 10743 25171
rect 18759 17955 18811 18007
rect 18759 17811 18811 17863
rect 18759 16269 18811 16321
rect 18759 15717 18811 15769
rect 10691 12831 10743 12883
rect 10691 12687 10743 12739
rect 10691 12545 10743 12597
rect 10691 12405 10743 12457
rect 18759 5241 18811 5293
rect 18759 5097 18811 5149
rect 18759 3555 18811 3607
rect 18759 3003 18811 3055
<< metal2 >>
rect 21028 44879 21112 44912
rect 21028 44823 21042 44879
rect 21098 44823 21112 44879
rect 21028 44790 21112 44823
rect 21580 44879 21664 44912
rect 21580 44823 21594 44879
rect 21650 44823 21664 44879
rect 21580 44790 21664 44823
rect 22132 44879 22216 44912
rect 22132 44823 22146 44879
rect 22202 44823 22216 44879
rect 22132 44790 22216 44823
rect 22684 44879 22768 44912
rect 22684 44823 22698 44879
rect 22754 44823 22768 44879
rect 22684 44790 22768 44823
rect 23236 44879 23320 44912
rect 23236 44823 23250 44879
rect 23306 44823 23320 44879
rect 23236 44790 23320 44823
rect 23788 44879 23872 44912
rect 23788 44823 23802 44879
rect 23858 44823 23872 44879
rect 23788 44790 23872 44823
rect 24340 44879 24424 44912
rect 24340 44823 24354 44879
rect 24410 44823 24424 44879
rect 24340 44790 24424 44823
rect 24892 44879 24976 44912
rect 24892 44823 24906 44879
rect 24962 44823 24976 44879
rect 24892 44790 24976 44823
rect 25444 44879 25528 44912
rect 25444 44823 25458 44879
rect 25514 44823 25528 44879
rect 25444 44790 25528 44823
rect 25996 44879 26080 44912
rect 25996 44823 26010 44879
rect 26066 44823 26080 44879
rect 25996 44790 26080 44823
rect 26548 44879 26632 44912
rect 26548 44823 26562 44879
rect 26618 44823 26632 44879
rect 26548 44790 26632 44823
rect 27100 44879 27184 44912
rect 27100 44823 27114 44879
rect 27170 44823 27184 44879
rect 27100 44790 27184 44823
rect 27652 44879 27736 44912
rect 27652 44823 27666 44879
rect 27722 44823 27736 44879
rect 27652 44790 27736 44823
rect 28204 44879 28288 44912
rect 28204 44823 28218 44879
rect 28274 44823 28288 44879
rect 28204 44790 28288 44823
rect 28756 44879 28840 44912
rect 28756 44823 28770 44879
rect 28826 44823 28840 44879
rect 28756 44790 28840 44823
rect 29308 44879 29392 44912
rect 29308 44823 29322 44879
rect 29378 44823 29392 44879
rect 29308 44790 29392 44823
rect 21038 44758 21102 44790
rect 21590 44758 21654 44790
rect 22142 44758 22206 44790
rect 22694 44758 22758 44790
rect 23246 44758 23310 44790
rect 23798 44758 23862 44790
rect 24350 44758 24414 44790
rect 24902 44758 24966 44790
rect 25454 44758 25518 44790
rect 26006 44758 26070 44790
rect 26558 44758 26622 44790
rect 27110 44758 27174 44790
rect 27662 44758 27726 44790
rect 28214 44758 28278 44790
rect 28766 44758 28830 44790
rect 29318 44758 29382 44790
rect 10676 38313 10756 38324
rect 10676 38257 10689 38313
rect 10745 38257 10756 38313
rect 10676 38244 10756 38257
rect 10676 38169 10756 38180
rect 10676 38113 10689 38169
rect 10745 38113 10756 38169
rect 10676 38100 10756 38113
rect 10676 38027 10756 38038
rect 10676 37971 10689 38027
rect 10745 37971 10756 38027
rect 10676 37958 10756 37971
rect 10676 37887 10756 37898
rect 10676 37831 10689 37887
rect 10745 37831 10756 37887
rect 10676 37818 10756 37831
rect 19072 36972 19148 36982
rect 19072 36966 19082 36972
rect 18748 36920 19082 36966
rect 19072 36916 19082 36920
rect 19138 36916 19148 36972
rect 19072 36906 19148 36916
rect 19072 36698 19148 36708
rect 19072 36694 19082 36698
rect 18748 36648 19082 36694
rect 19072 36642 19082 36648
rect 19138 36642 19148 36698
rect 19072 36632 19148 36642
rect 19072 36426 19148 36436
rect 19072 36422 19082 36426
rect 18748 36376 19082 36422
rect 19072 36370 19082 36376
rect 19138 36370 19148 36426
rect 19072 36360 19148 36370
rect 18744 30723 18824 30734
rect 18744 30667 18757 30723
rect 18813 30667 18824 30723
rect 18744 30654 18824 30667
rect 18744 30579 18824 30590
rect 18744 30523 18757 30579
rect 18813 30523 18824 30579
rect 18744 30510 18824 30523
rect 18744 29037 18824 29048
rect 18744 28981 18757 29037
rect 18813 28981 18824 29037
rect 18744 28968 18824 28981
rect 18744 28485 18824 28496
rect 18744 28429 18757 28485
rect 18813 28429 18824 28485
rect 18744 28416 18824 28429
rect 10676 25599 10756 25610
rect 10676 25543 10689 25599
rect 10745 25543 10756 25599
rect 10676 25530 10756 25543
rect 10676 25455 10756 25466
rect 10676 25399 10689 25455
rect 10745 25399 10756 25455
rect 10676 25386 10756 25399
rect 10676 25313 10756 25324
rect 10676 25257 10689 25313
rect 10745 25257 10756 25313
rect 10676 25244 10756 25257
rect 10676 25173 10756 25184
rect 10676 25117 10689 25173
rect 10745 25117 10756 25173
rect 10676 25104 10756 25117
rect 19072 24258 19148 24268
rect 19072 24252 19082 24258
rect 18748 24206 19082 24252
rect 19072 24202 19082 24206
rect 19138 24202 19148 24258
rect 19072 24192 19148 24202
rect 19072 23984 19148 23994
rect 19072 23980 19082 23984
rect 18748 23934 19082 23980
rect 19072 23928 19082 23934
rect 19138 23928 19148 23984
rect 19072 23918 19148 23928
rect 19072 23712 19148 23722
rect 19072 23708 19082 23712
rect 18748 23662 19082 23708
rect 19072 23656 19082 23662
rect 19138 23656 19148 23712
rect 19072 23646 19148 23656
rect 18744 18009 18824 18020
rect 18744 17953 18757 18009
rect 18813 17953 18824 18009
rect 18744 17940 18824 17953
rect 18744 17865 18824 17876
rect 18744 17809 18757 17865
rect 18813 17809 18824 17865
rect 18744 17796 18824 17809
rect 18744 16323 18824 16334
rect 18744 16267 18757 16323
rect 18813 16267 18824 16323
rect 18744 16254 18824 16267
rect 18744 15771 18824 15782
rect 18744 15715 18757 15771
rect 18813 15715 18824 15771
rect 18744 15702 18824 15715
rect 10676 12885 10756 12896
rect 10676 12829 10689 12885
rect 10745 12829 10756 12885
rect 10676 12816 10756 12829
rect 10676 12741 10756 12752
rect 10676 12685 10689 12741
rect 10745 12685 10756 12741
rect 10676 12672 10756 12685
rect 10676 12599 10756 12610
rect 10676 12543 10689 12599
rect 10745 12543 10756 12599
rect 10676 12530 10756 12543
rect 10676 12459 10756 12470
rect 10676 12403 10689 12459
rect 10745 12403 10756 12459
rect 10676 12390 10756 12403
rect 19072 11544 19148 11554
rect 19072 11538 19082 11544
rect 18748 11492 19082 11538
rect 19072 11488 19082 11492
rect 19138 11488 19148 11544
rect 19072 11478 19148 11488
rect 19072 11270 19148 11280
rect 19072 11266 19082 11270
rect 18748 11220 19082 11266
rect 19072 11214 19082 11220
rect 19138 11214 19148 11270
rect 19072 11204 19148 11214
rect 19072 10998 19148 11008
rect 19072 10994 19082 10998
rect 18748 10948 19082 10994
rect 19072 10942 19082 10948
rect 19138 10942 19148 10998
rect 19072 10932 19148 10942
rect 18744 5295 18824 5306
rect 18744 5239 18757 5295
rect 18813 5239 18824 5295
rect 18744 5226 18824 5239
rect 18744 5151 18824 5162
rect 18744 5095 18757 5151
rect 18813 5095 18824 5151
rect 18744 5082 18824 5095
rect 18744 3609 18824 3620
rect 18744 3553 18757 3609
rect 18813 3553 18824 3609
rect 18744 3540 18824 3553
rect 18744 3057 18824 3068
rect 18744 3001 18757 3057
rect 18813 3001 18824 3057
rect 18744 2988 18824 3001
<< via2 >>
rect 21042 44823 21098 44879
rect 21594 44823 21650 44879
rect 22146 44823 22202 44879
rect 22698 44823 22754 44879
rect 23250 44823 23306 44879
rect 23802 44823 23858 44879
rect 24354 44823 24410 44879
rect 24906 44823 24962 44879
rect 25458 44823 25514 44879
rect 26010 44823 26066 44879
rect 26562 44823 26618 44879
rect 27114 44823 27170 44879
rect 27666 44823 27722 44879
rect 28218 44823 28274 44879
rect 28770 44823 28826 44879
rect 29322 44823 29378 44879
rect 10689 38311 10745 38313
rect 10689 38259 10691 38311
rect 10691 38259 10743 38311
rect 10743 38259 10745 38311
rect 10689 38257 10745 38259
rect 10689 38167 10745 38169
rect 10689 38115 10691 38167
rect 10691 38115 10743 38167
rect 10743 38115 10745 38167
rect 10689 38113 10745 38115
rect 10689 38025 10745 38027
rect 10689 37973 10691 38025
rect 10691 37973 10743 38025
rect 10743 37973 10745 38025
rect 10689 37971 10745 37973
rect 10689 37885 10745 37887
rect 10689 37833 10691 37885
rect 10691 37833 10743 37885
rect 10743 37833 10745 37885
rect 10689 37831 10745 37833
rect 19082 36916 19138 36972
rect 19082 36642 19138 36698
rect 19082 36370 19138 36426
rect 18757 30721 18813 30723
rect 18757 30669 18759 30721
rect 18759 30669 18811 30721
rect 18811 30669 18813 30721
rect 18757 30667 18813 30669
rect 18757 30577 18813 30579
rect 18757 30525 18759 30577
rect 18759 30525 18811 30577
rect 18811 30525 18813 30577
rect 18757 30523 18813 30525
rect 18757 29035 18813 29037
rect 18757 28983 18759 29035
rect 18759 28983 18811 29035
rect 18811 28983 18813 29035
rect 18757 28981 18813 28983
rect 18757 28483 18813 28485
rect 18757 28431 18759 28483
rect 18759 28431 18811 28483
rect 18811 28431 18813 28483
rect 18757 28429 18813 28431
rect 10689 25597 10745 25599
rect 10689 25545 10691 25597
rect 10691 25545 10743 25597
rect 10743 25545 10745 25597
rect 10689 25543 10745 25545
rect 10689 25453 10745 25455
rect 10689 25401 10691 25453
rect 10691 25401 10743 25453
rect 10743 25401 10745 25453
rect 10689 25399 10745 25401
rect 10689 25311 10745 25313
rect 10689 25259 10691 25311
rect 10691 25259 10743 25311
rect 10743 25259 10745 25311
rect 10689 25257 10745 25259
rect 10689 25171 10745 25173
rect 10689 25119 10691 25171
rect 10691 25119 10743 25171
rect 10743 25119 10745 25171
rect 10689 25117 10745 25119
rect 19082 24202 19138 24258
rect 19082 23928 19138 23984
rect 19082 23656 19138 23712
rect 18757 18007 18813 18009
rect 18757 17955 18759 18007
rect 18759 17955 18811 18007
rect 18811 17955 18813 18007
rect 18757 17953 18813 17955
rect 18757 17863 18813 17865
rect 18757 17811 18759 17863
rect 18759 17811 18811 17863
rect 18811 17811 18813 17863
rect 18757 17809 18813 17811
rect 18757 16321 18813 16323
rect 18757 16269 18759 16321
rect 18759 16269 18811 16321
rect 18811 16269 18813 16321
rect 18757 16267 18813 16269
rect 18757 15769 18813 15771
rect 18757 15717 18759 15769
rect 18759 15717 18811 15769
rect 18811 15717 18813 15769
rect 18757 15715 18813 15717
rect 10689 12883 10745 12885
rect 10689 12831 10691 12883
rect 10691 12831 10743 12883
rect 10743 12831 10745 12883
rect 10689 12829 10745 12831
rect 10689 12739 10745 12741
rect 10689 12687 10691 12739
rect 10691 12687 10743 12739
rect 10743 12687 10745 12739
rect 10689 12685 10745 12687
rect 10689 12597 10745 12599
rect 10689 12545 10691 12597
rect 10691 12545 10743 12597
rect 10743 12545 10745 12597
rect 10689 12543 10745 12545
rect 10689 12457 10745 12459
rect 10689 12405 10691 12457
rect 10691 12405 10743 12457
rect 10743 12405 10745 12457
rect 10689 12403 10745 12405
rect 19082 11488 19138 11544
rect 19082 11214 19138 11270
rect 19082 10942 19138 10998
rect 18757 5293 18813 5295
rect 18757 5241 18759 5293
rect 18759 5241 18811 5293
rect 18811 5241 18813 5293
rect 18757 5239 18813 5241
rect 18757 5149 18813 5151
rect 18757 5097 18759 5149
rect 18759 5097 18811 5149
rect 18811 5097 18813 5149
rect 18757 5095 18813 5097
rect 18757 3607 18813 3609
rect 18757 3555 18759 3607
rect 18759 3555 18811 3607
rect 18811 3555 18813 3607
rect 18757 3553 18813 3555
rect 18757 3055 18813 3057
rect 18757 3003 18759 3055
rect 18759 3003 18811 3055
rect 18811 3003 18813 3055
rect 18757 3001 18813 3003
<< metal3 >>
rect 9722 44846 9728 44910
rect 9792 44846 9798 44910
rect 21028 44883 21112 44912
rect 9730 44280 9790 44846
rect 21028 44819 21038 44883
rect 21102 44819 21112 44883
rect 21028 44790 21112 44819
rect 21580 44883 21664 44912
rect 21580 44819 21590 44883
rect 21654 44819 21664 44883
rect 21580 44790 21664 44819
rect 22132 44883 22216 44912
rect 22132 44819 22142 44883
rect 22206 44819 22216 44883
rect 22132 44790 22216 44819
rect 22684 44883 22768 44912
rect 22684 44819 22694 44883
rect 22758 44819 22768 44883
rect 22684 44790 22768 44819
rect 23236 44883 23320 44912
rect 23236 44819 23246 44883
rect 23310 44819 23320 44883
rect 23236 44790 23320 44819
rect 23788 44883 23872 44912
rect 23788 44819 23798 44883
rect 23862 44819 23872 44883
rect 23788 44790 23872 44819
rect 24340 44883 24424 44912
rect 24340 44819 24350 44883
rect 24414 44819 24424 44883
rect 24340 44790 24424 44819
rect 24892 44883 24976 44912
rect 24892 44819 24902 44883
rect 24966 44819 24976 44883
rect 24892 44790 24976 44819
rect 25444 44883 25528 44912
rect 25444 44819 25454 44883
rect 25518 44819 25528 44883
rect 25444 44790 25528 44819
rect 25996 44883 26080 44912
rect 25996 44819 26006 44883
rect 26070 44819 26080 44883
rect 25996 44790 26080 44819
rect 26548 44883 26632 44912
rect 26548 44819 26558 44883
rect 26622 44819 26632 44883
rect 26548 44790 26632 44819
rect 27100 44883 27184 44912
rect 27100 44819 27110 44883
rect 27174 44819 27184 44883
rect 27100 44790 27184 44819
rect 27652 44883 27736 44912
rect 27652 44819 27662 44883
rect 27726 44819 27736 44883
rect 27652 44790 27736 44819
rect 28204 44883 28288 44912
rect 28204 44819 28214 44883
rect 28278 44819 28288 44883
rect 28204 44790 28288 44819
rect 28756 44883 28840 44912
rect 28756 44819 28766 44883
rect 28830 44819 28840 44883
rect 28756 44790 28840 44819
rect 29308 44883 29392 44912
rect 29308 44819 29318 44883
rect 29382 44819 29392 44883
rect 29308 44790 29392 44819
rect 24125 44280 24443 44285
rect 30525 44280 30843 44285
rect 380 44279 30844 44280
rect 380 44044 24125 44279
rect 380 43980 746 44044
rect 810 43980 24125 44044
rect 380 43961 24125 43980
rect 24443 44000 30525 44279
rect 24443 43961 24680 44000
rect 380 43960 24680 43961
rect 25180 43961 30525 44000
rect 30843 43961 30844 44279
rect 25180 43960 30844 43961
rect 380 43700 700 43960
rect 24125 43955 24443 43960
rect 30525 43955 30843 43960
rect 380 43400 390 43700
rect 690 43400 700 43700
rect 380 43390 700 43400
rect 13798 42616 20540 42644
rect 13798 42552 18828 42616
rect 18892 42552 20540 42616
rect 13798 42524 20540 42552
rect 13798 42344 20540 42372
rect 13798 42280 18276 42344
rect 18340 42280 20540 42344
rect 13798 42252 20540 42280
rect 13798 42072 20540 42100
rect 13798 42008 17724 42072
rect 17788 42008 20540 42072
rect 13798 41980 20540 42008
rect 13798 41800 20540 41828
rect 13798 41736 17172 41800
rect 17236 41736 20540 41800
rect 13798 41708 20540 41736
rect 13798 41528 20540 41556
rect 13798 41464 16620 41528
rect 16684 41464 20540 41528
rect 13798 41436 20540 41464
rect 13798 41256 20540 41284
rect 13798 41192 16068 41256
rect 16132 41192 20540 41256
rect 13798 41164 20540 41192
rect 13798 40984 20540 41012
rect 13798 40920 15516 40984
rect 15580 40920 20540 40984
rect 13798 40892 20540 40920
rect 13798 40712 20540 40740
rect 13798 40648 14964 40712
rect 15028 40648 20540 40712
rect 13798 40620 20540 40648
rect 13798 40440 20540 40468
rect 13798 40376 14412 40440
rect 14476 40376 20540 40440
rect 13798 40348 20540 40376
rect 13798 40168 20540 40196
rect 13798 40104 13860 40168
rect 13924 40104 20540 40168
rect 13798 40076 20540 40104
rect 10676 38316 10756 38324
rect 10676 38313 20549 38316
rect 10676 38257 10689 38313
rect 10745 38257 20549 38313
rect 10676 38254 20549 38257
rect 10676 38244 10756 38254
rect 10676 38172 10756 38180
rect 10676 38169 20379 38172
rect 10676 38113 10689 38169
rect 10745 38113 20379 38169
rect 10676 38110 20379 38113
rect 10676 38100 10756 38110
rect 10676 38030 10756 38038
rect 10676 38027 20209 38030
rect 10676 37971 10689 38027
rect 10745 37971 20209 38027
rect 10676 37968 20209 37971
rect 10676 37958 10756 37968
rect 10676 37890 10756 37898
rect 10676 37887 19956 37890
rect 10676 37831 10689 37887
rect 10745 37831 19956 37887
rect 10676 37828 19956 37831
rect 10676 37818 10756 37828
rect 200 37734 2380 37754
rect 200 36950 248 37734
rect 872 36950 2380 37734
rect 19894 37179 19956 37828
rect 20147 37453 20209 37968
rect 20317 37737 20379 38110
rect 20487 37933 20549 38254
rect 20317 37675 20547 37737
rect 20147 37391 20531 37453
rect 19894 37117 20551 37179
rect 200 36940 2380 36950
rect 19072 36980 19148 36982
rect 19072 36972 20344 36980
rect 19072 36916 19082 36972
rect 19138 36916 20344 36972
rect 19072 36908 20344 36916
rect 19072 36906 19148 36908
rect 19072 36706 19148 36708
rect 19072 36698 20154 36706
rect 19072 36642 19082 36698
rect 19138 36642 20154 36698
rect 19072 36634 20154 36642
rect 19072 36632 19148 36634
rect 19072 36434 19148 36436
rect 19072 36426 19934 36434
rect 19072 36370 19082 36426
rect 19138 36370 19934 36426
rect 19072 36362 19934 36370
rect 19072 36360 19148 36362
rect 200 35925 2380 35960
rect 200 34981 248 35925
rect 872 34981 2380 35925
rect 19023 35652 19201 35657
rect 17672 35634 19202 35652
rect 17672 35490 17695 35634
rect 17839 35490 19040 35634
rect 19184 35490 19202 35634
rect 17672 35472 19202 35490
rect 19023 35467 19201 35472
rect 19862 35272 19934 36362
rect 20082 35542 20154 36634
rect 20272 35812 20344 36908
rect 20272 35740 20556 35812
rect 20082 35470 20532 35542
rect 19862 35200 20538 35272
rect 200 34936 2380 34981
rect 18744 30726 18824 30734
rect 18744 30723 20541 30726
rect 18744 30667 18757 30723
rect 18813 30667 20541 30723
rect 18744 30664 20541 30667
rect 18744 30654 18824 30664
rect 18744 30582 18824 30590
rect 18744 30579 20389 30582
rect 18744 30523 18757 30579
rect 18813 30523 20389 30579
rect 18744 30520 20389 30523
rect 18744 30510 18824 30520
rect 20327 29551 20389 30520
rect 20479 29765 20541 30664
rect 20327 29489 20513 29551
rect 20123 29213 20521 29275
rect 18744 29040 18824 29048
rect 20123 29040 20185 29213
rect 18744 29037 20185 29040
rect 18744 28981 18757 29037
rect 18813 28981 20185 29037
rect 18744 28978 20185 28981
rect 18744 28968 18824 28978
rect 20327 28951 20537 29013
rect 18744 28488 18824 28496
rect 20327 28488 20389 28951
rect 18744 28485 20389 28488
rect 18744 28429 18757 28485
rect 18813 28429 20389 28485
rect 18744 28426 20389 28429
rect 18744 28416 18824 28426
rect 19829 26722 20007 26727
rect 17594 26704 20008 26722
rect 17594 26560 17617 26704
rect 17761 26560 19846 26704
rect 19990 26560 20008 26704
rect 17594 26542 20008 26560
rect 19829 26537 20007 26542
rect 10676 25602 10756 25610
rect 10676 25599 20545 25602
rect 10676 25543 10689 25599
rect 10745 25543 20545 25599
rect 10676 25540 20545 25543
rect 10676 25530 10756 25540
rect 10676 25458 10756 25466
rect 10676 25455 20377 25458
rect 10676 25399 10689 25455
rect 10745 25399 20377 25455
rect 10676 25396 20377 25399
rect 10676 25386 10756 25396
rect 10676 25316 10756 25324
rect 10676 25313 20219 25316
rect 10676 25257 10689 25313
rect 10745 25257 20219 25313
rect 10676 25254 20219 25257
rect 10676 25244 10756 25254
rect 10676 25176 10756 25184
rect 10676 25173 20049 25176
rect 10676 25117 10689 25173
rect 10745 25117 20049 25173
rect 10676 25114 20049 25117
rect 10676 25104 10756 25114
rect 200 25007 2380 25040
rect 200 24143 248 25007
rect 872 24143 2380 25007
rect 19987 24461 20049 25114
rect 20157 24655 20219 25254
rect 20315 24927 20377 25396
rect 20483 25149 20545 25540
rect 20315 24865 20547 24927
rect 20157 24593 20539 24655
rect 19987 24399 20247 24461
rect 20185 24387 20247 24399
rect 20185 24325 20559 24387
rect 19072 24266 19148 24268
rect 19072 24258 20056 24266
rect 19072 24202 19082 24258
rect 19138 24202 20056 24258
rect 19072 24194 20056 24202
rect 19072 24192 19148 24194
rect 200 24120 2380 24143
rect 19984 24120 20056 24194
rect 19984 24048 20542 24120
rect 19072 23992 19148 23994
rect 19072 23984 19870 23992
rect 19072 23928 19082 23984
rect 19138 23928 19870 23984
rect 19072 23920 19870 23928
rect 19072 23918 19148 23920
rect 19798 23850 19870 23920
rect 19798 23778 20550 23850
rect 19072 23720 19148 23722
rect 19072 23712 19644 23720
rect 19072 23656 19082 23712
rect 19138 23656 19644 23712
rect 19072 23648 19644 23656
rect 19072 23646 19148 23648
rect 19572 23582 19644 23648
rect 19572 23510 20526 23582
rect 200 23118 2380 23140
rect 200 22254 248 23118
rect 872 22254 2380 23118
rect 200 22222 2380 22254
rect 20241 18071 20561 18133
rect 18744 18012 18824 18020
rect 20241 18012 20303 18071
rect 18744 18009 20303 18012
rect 18744 17953 18757 18009
rect 18813 17953 20303 18009
rect 18744 17950 20303 17953
rect 18744 17940 18824 17950
rect 18744 17868 18824 17876
rect 18744 17865 20531 17868
rect 18744 17809 18757 17865
rect 18813 17809 20531 17865
rect 18744 17806 20531 17809
rect 18744 17796 18824 17806
rect 20331 17519 20541 17581
rect 18744 16326 18824 16334
rect 20331 16326 20393 17519
rect 18744 16323 20393 16326
rect 18744 16267 18757 16323
rect 18813 16267 20393 16323
rect 18744 16264 20393 16267
rect 18744 16254 18824 16264
rect 18744 15774 18824 15782
rect 20493 15774 20555 17317
rect 18744 15771 20555 15774
rect 18744 15715 18757 15771
rect 18813 15715 20555 15771
rect 18744 15712 20555 15715
rect 18744 15702 18824 15712
rect 19570 13998 19950 14010
rect 17860 13980 19950 13998
rect 17860 13836 17883 13980
rect 18027 13836 19594 13980
rect 19738 13836 19950 13980
rect 17860 13818 19950 13836
rect 19570 13810 19950 13818
rect 18514 13447 20533 13509
rect 10676 12888 10756 12896
rect 18514 12888 18576 13447
rect 10676 12885 18576 12888
rect 10676 12829 10689 12885
rect 10745 12829 18576 12885
rect 10676 12826 18576 12829
rect 18657 13175 20555 13237
rect 10676 12816 10756 12826
rect 10676 12744 10756 12752
rect 18657 12744 18719 13175
rect 10676 12741 18719 12744
rect 10676 12685 10689 12741
rect 10745 12685 18719 12741
rect 10676 12682 18719 12685
rect 18801 12905 20535 12967
rect 10676 12672 10756 12682
rect 10676 12602 10756 12610
rect 18801 12602 18863 12905
rect 10676 12599 18863 12602
rect 10676 12543 10689 12599
rect 10745 12543 18863 12599
rect 10676 12540 18863 12543
rect 18971 12631 20539 12693
rect 10676 12530 10756 12540
rect 10676 12462 10756 12470
rect 18971 12462 19033 12631
rect 10676 12459 19033 12462
rect 10676 12403 10689 12459
rect 10745 12403 19033 12459
rect 10676 12400 19033 12403
rect 10676 12390 10756 12400
rect 20034 12356 20534 12428
rect 200 12280 2380 12326
rect 200 11416 248 12280
rect 872 11416 2380 12280
rect 19072 11552 19148 11554
rect 20034 11552 20106 12356
rect 19072 11544 20106 11552
rect 19072 11488 19082 11544
rect 19138 11488 20106 11544
rect 19072 11480 20106 11488
rect 20282 12078 20550 12150
rect 19072 11478 19148 11480
rect 200 11380 2380 11416
rect 19072 11278 19148 11280
rect 20282 11278 20354 12078
rect 19072 11270 20354 11278
rect 19072 11214 19082 11270
rect 19138 11214 20354 11270
rect 19072 11206 20354 11214
rect 19072 11204 19148 11206
rect 19072 11006 19148 11008
rect 20502 11006 20574 11878
rect 19072 10998 20574 11006
rect 19072 10942 19082 10998
rect 19138 10942 20574 10998
rect 19072 10934 20574 10942
rect 19072 10932 19148 10934
rect 200 10391 2380 10400
rect 200 9527 248 10391
rect 872 9527 2380 10391
rect 200 9508 2380 9527
rect 19785 6373 20557 6435
rect 18744 5298 18824 5306
rect 19785 5298 19847 6373
rect 18744 5295 19847 5298
rect 18744 5239 18757 5295
rect 18813 5239 19847 5295
rect 18744 5236 19847 5239
rect 19951 6101 20547 6163
rect 18744 5226 18824 5236
rect 18744 5154 18824 5162
rect 19951 5154 20013 6101
rect 18744 5151 20013 5154
rect 18744 5095 18757 5151
rect 18813 5095 20013 5151
rect 18744 5092 20013 5095
rect 20133 5833 20547 5895
rect 18744 5082 18824 5092
rect 18744 3612 18824 3620
rect 20133 3612 20195 5833
rect 18744 3609 20195 3612
rect 18744 3553 18757 3609
rect 18813 3553 20195 3609
rect 18744 3550 20195 3553
rect 20329 5561 20551 5623
rect 18744 3540 18824 3550
rect 18744 3060 18824 3068
rect 20329 3060 20391 5561
rect 18744 3057 20391 3060
rect 18744 3001 18757 3057
rect 18813 3001 20391 3057
rect 18744 2998 20391 3001
rect 18744 2988 18824 2998
rect 19022 2769 19202 2792
rect 19022 2625 19040 2769
rect 19184 2625 19202 2769
rect 19022 830 19202 2625
rect 18770 829 19202 830
rect 18765 812 19202 829
rect 18765 668 18788 812
rect 18932 668 19202 812
rect 18765 651 19202 668
rect 18770 650 19202 651
<< via3 >>
rect 9728 44846 9792 44910
rect 21038 44879 21102 44883
rect 21038 44823 21042 44879
rect 21042 44823 21098 44879
rect 21098 44823 21102 44879
rect 21038 44819 21102 44823
rect 21590 44879 21654 44883
rect 21590 44823 21594 44879
rect 21594 44823 21650 44879
rect 21650 44823 21654 44879
rect 21590 44819 21654 44823
rect 22142 44879 22206 44883
rect 22142 44823 22146 44879
rect 22146 44823 22202 44879
rect 22202 44823 22206 44879
rect 22142 44819 22206 44823
rect 22694 44879 22758 44883
rect 22694 44823 22698 44879
rect 22698 44823 22754 44879
rect 22754 44823 22758 44879
rect 22694 44819 22758 44823
rect 23246 44879 23310 44883
rect 23246 44823 23250 44879
rect 23250 44823 23306 44879
rect 23306 44823 23310 44879
rect 23246 44819 23310 44823
rect 23798 44879 23862 44883
rect 23798 44823 23802 44879
rect 23802 44823 23858 44879
rect 23858 44823 23862 44879
rect 23798 44819 23862 44823
rect 24350 44879 24414 44883
rect 24350 44823 24354 44879
rect 24354 44823 24410 44879
rect 24410 44823 24414 44879
rect 24350 44819 24414 44823
rect 24902 44879 24966 44883
rect 24902 44823 24906 44879
rect 24906 44823 24962 44879
rect 24962 44823 24966 44879
rect 24902 44819 24966 44823
rect 25454 44879 25518 44883
rect 25454 44823 25458 44879
rect 25458 44823 25514 44879
rect 25514 44823 25518 44879
rect 25454 44819 25518 44823
rect 26006 44879 26070 44883
rect 26006 44823 26010 44879
rect 26010 44823 26066 44879
rect 26066 44823 26070 44879
rect 26006 44819 26070 44823
rect 26558 44879 26622 44883
rect 26558 44823 26562 44879
rect 26562 44823 26618 44879
rect 26618 44823 26622 44879
rect 26558 44819 26622 44823
rect 27110 44879 27174 44883
rect 27110 44823 27114 44879
rect 27114 44823 27170 44879
rect 27170 44823 27174 44879
rect 27110 44819 27174 44823
rect 27662 44879 27726 44883
rect 27662 44823 27666 44879
rect 27666 44823 27722 44879
rect 27722 44823 27726 44879
rect 27662 44819 27726 44823
rect 28214 44879 28278 44883
rect 28214 44823 28218 44879
rect 28218 44823 28274 44879
rect 28274 44823 28278 44879
rect 28214 44819 28278 44823
rect 28766 44879 28830 44883
rect 28766 44823 28770 44879
rect 28770 44823 28826 44879
rect 28826 44823 28830 44879
rect 28766 44819 28830 44823
rect 29318 44879 29382 44883
rect 29318 44823 29322 44879
rect 29322 44823 29378 44879
rect 29378 44823 29382 44879
rect 29318 44819 29382 44823
rect 746 43980 810 44044
rect 24125 43961 24443 44279
rect 30525 43961 30843 44279
rect 390 43400 690 43700
rect 18828 42552 18892 42616
rect 18276 42280 18340 42344
rect 17724 42008 17788 42072
rect 17172 41736 17236 41800
rect 16620 41464 16684 41528
rect 16068 41192 16132 41256
rect 15516 40920 15580 40984
rect 14964 40648 15028 40712
rect 14412 40376 14476 40440
rect 13860 40104 13924 40168
rect 248 36950 872 37734
rect 248 34981 872 35925
rect 17695 35490 17839 35634
rect 19040 35490 19184 35634
rect 17617 26560 17761 26704
rect 19846 26560 19990 26704
rect 248 24143 872 25007
rect 248 22254 872 23118
rect 17883 13836 18027 13980
rect 19594 13836 19738 13980
rect 248 11416 872 12280
rect 248 9527 872 10391
rect 19040 2625 19184 2769
rect 18788 668 18932 812
<< metal4 >>
rect 6134 44804 6194 45152
rect 6686 44804 6746 45152
rect 7238 44804 7298 45152
rect 7790 44804 7850 45152
rect 8342 44804 8402 45152
rect 8894 44804 8954 45152
rect 9446 44908 9506 45152
rect 9727 44910 9793 44911
rect 9727 44908 9728 44910
rect 9446 44848 9728 44908
rect 9727 44846 9728 44848
rect 9792 44908 9793 44910
rect 9998 44908 10058 45152
rect 9792 44848 10058 44908
rect 9792 44846 9793 44848
rect 9727 44845 9793 44846
rect 10550 44804 10610 45152
rect 11102 44804 11162 45152
rect 11654 44804 11714 45152
rect 12206 44804 12266 45152
rect 12758 44804 12818 45152
rect 13310 44804 13370 45152
rect 13862 44858 13922 45152
rect 14414 44858 14474 45152
rect 14966 44858 15026 45152
rect 15518 44858 15578 45152
rect 16070 44858 16130 45152
rect 16622 44858 16682 45152
rect 17174 44858 17234 45152
rect 17726 44858 17786 45152
rect 18278 44858 18338 45152
rect 18830 44858 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44912 21098 45152
rect 21590 44912 21650 45152
rect 22142 44912 22202 45152
rect 22694 44912 22754 45152
rect 23246 44912 23306 45152
rect 23798 44912 23858 45152
rect 24350 44912 24410 45152
rect 24902 44912 24962 45152
rect 25454 44912 25514 45152
rect 26006 44912 26066 45152
rect 26558 44912 26618 45152
rect 27110 44912 27170 45152
rect 27662 44912 27722 45152
rect 28214 44912 28274 45152
rect 28766 44912 28826 45152
rect 29318 44912 29378 45152
rect 21028 44883 21112 44912
rect 1120 44704 9360 44804
rect 10144 44704 13440 44804
rect 1120 44556 13440 44704
rect 200 44044 920 44152
rect 200 43980 746 44044
rect 810 43980 920 44044
rect 200 43700 920 43980
rect 200 43400 390 43700
rect 690 43400 920 43700
rect 200 37734 920 43400
rect 200 36950 248 37734
rect 872 36950 920 37734
rect 200 35925 920 36950
rect 200 34981 248 35925
rect 872 34981 920 35925
rect 200 25007 920 34981
rect 200 24143 248 25007
rect 872 24143 920 25007
rect 200 23118 920 24143
rect 200 22254 248 23118
rect 872 22254 920 23118
rect 200 12280 920 22254
rect 200 11416 248 12280
rect 872 11416 920 12280
rect 200 10391 920 11416
rect 200 9527 248 10391
rect 872 9527 920 10391
rect 200 1000 920 9527
rect 1120 43556 1840 44556
rect 1120 43284 1324 43556
rect 1596 43284 1840 43556
rect 1120 1000 1840 43284
rect 13822 40168 13962 44858
rect 13822 40104 13860 40168
rect 13924 40104 13962 40168
rect 13822 40028 13962 40104
rect 14374 40440 14514 44858
rect 14374 40376 14412 40440
rect 14476 40376 14514 40440
rect 14374 40028 14514 40376
rect 14926 40712 15066 44858
rect 14926 40648 14964 40712
rect 15028 40648 15066 40712
rect 14926 40028 15066 40648
rect 15478 40984 15618 44858
rect 15478 40920 15516 40984
rect 15580 40920 15618 40984
rect 15478 40028 15618 40920
rect 16030 41256 16170 44858
rect 16030 41192 16068 41256
rect 16132 41192 16170 41256
rect 16030 40028 16170 41192
rect 16582 41528 16722 44858
rect 16582 41464 16620 41528
rect 16684 41464 16722 41528
rect 16582 40028 16722 41464
rect 17134 41800 17274 44858
rect 17134 41736 17172 41800
rect 17236 41736 17274 41800
rect 17134 40028 17274 41736
rect 17686 42072 17826 44858
rect 17686 42008 17724 42072
rect 17788 42008 17826 42072
rect 17686 40028 17826 42008
rect 18238 42344 18378 44858
rect 18238 42280 18276 42344
rect 18340 42280 18378 42344
rect 18238 40028 18378 42280
rect 18790 42616 18930 44858
rect 21028 44819 21038 44883
rect 21102 44819 21112 44883
rect 21028 44790 21112 44819
rect 21580 44883 21664 44912
rect 21580 44819 21590 44883
rect 21654 44819 21664 44883
rect 21580 44790 21664 44819
rect 22132 44883 22216 44912
rect 22132 44819 22142 44883
rect 22206 44819 22216 44883
rect 22132 44790 22216 44819
rect 22684 44883 22768 44912
rect 22684 44819 22694 44883
rect 22758 44819 22768 44883
rect 22684 44790 22768 44819
rect 23236 44883 23320 44912
rect 23236 44819 23246 44883
rect 23310 44819 23320 44883
rect 23236 44790 23320 44819
rect 23788 44883 23872 44912
rect 23788 44819 23798 44883
rect 23862 44819 23872 44883
rect 23788 44790 23872 44819
rect 24340 44883 24424 44912
rect 24340 44819 24350 44883
rect 24414 44819 24424 44883
rect 24340 44790 24424 44819
rect 24892 44883 24976 44912
rect 24892 44819 24902 44883
rect 24966 44819 24976 44883
rect 24892 44790 24976 44819
rect 25444 44883 25528 44912
rect 25444 44819 25454 44883
rect 25518 44819 25528 44883
rect 25444 44790 25528 44819
rect 25996 44883 26080 44912
rect 25996 44819 26006 44883
rect 26070 44819 26080 44883
rect 25996 44790 26080 44819
rect 26548 44883 26632 44912
rect 26548 44819 26558 44883
rect 26622 44819 26632 44883
rect 26548 44790 26632 44819
rect 27100 44883 27184 44912
rect 27100 44819 27110 44883
rect 27174 44819 27184 44883
rect 27100 44790 27184 44819
rect 27652 44883 27736 44912
rect 27652 44819 27662 44883
rect 27726 44819 27736 44883
rect 27652 44790 27736 44819
rect 28204 44883 28288 44912
rect 28204 44819 28214 44883
rect 28278 44819 28288 44883
rect 28204 44790 28288 44819
rect 28756 44883 28840 44912
rect 28756 44819 28766 44883
rect 28830 44819 28840 44883
rect 28756 44790 28840 44819
rect 29308 44883 29392 44912
rect 29308 44819 29318 44883
rect 29382 44819 29392 44883
rect 29308 44790 29392 44819
rect 18790 42552 18828 42616
rect 18892 42552 18930 42616
rect 18790 40028 18930 42552
rect 24124 44279 24444 44280
rect 24124 43961 24125 44279
rect 24443 43961 24444 44279
rect 17677 35634 17857 35653
rect 15663 35613 17569 35626
rect 17677 35613 17695 35634
rect 15663 35536 17695 35613
rect 17513 35511 17695 35536
rect 17677 35490 17695 35511
rect 17839 35490 17857 35634
rect 17677 35471 17857 35490
rect 19022 35634 19202 35652
rect 19022 35490 19040 35634
rect 19184 35490 19202 35634
rect 17599 26722 17779 26723
rect 15482 26704 17779 26722
rect 15482 26560 17617 26704
rect 17761 26560 17779 26704
rect 15482 26542 17779 26560
rect 17599 26541 17779 26542
rect 17865 13998 18045 13999
rect 15482 13980 18045 13998
rect 15482 13836 17883 13980
rect 18027 13836 18045 13980
rect 15482 13818 18045 13836
rect 17865 13817 18045 13818
rect 19022 2787 19202 35490
rect 19828 26704 20308 26722
rect 19828 26560 19846 26704
rect 19990 26560 20308 26704
rect 19828 26542 20308 26560
rect 19570 13998 19950 14010
rect 19570 13980 19956 13998
rect 19570 13836 19594 13980
rect 19738 13836 19956 13980
rect 19570 13810 19956 13836
rect 19021 2769 19203 2787
rect 19021 2625 19040 2769
rect 19184 2625 19203 2769
rect 19021 2607 19203 2625
rect 15486 1112 19556 1292
rect 18770 812 18950 830
rect 18770 668 18788 812
rect 18932 668 18950 812
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 668
rect 19376 674 19556 1112
rect 19776 996 19956 13810
rect 20128 1308 20308 26542
rect 20128 1128 23796 1308
rect 19776 816 23484 996
rect 19376 494 22814 674
rect 22634 0 22814 494
rect 23304 610 23484 816
rect 23616 894 23796 1128
rect 24124 1000 24444 43961
rect 28258 44140 28318 44280
rect 30524 44279 30844 44280
rect 24784 1000 25104 43960
rect 30524 43961 30525 44279
rect 30843 43961 30844 44279
rect 30524 1000 30844 43961
rect 31184 1000 31504 43960
rect 23616 714 30542 894
rect 23304 430 26678 610
rect 26498 0 26678 430
rect 30362 0 30542 714
<< via4 >>
rect 1324 43284 1596 43556
rect 24784 43960 25104 44280
rect 31184 43960 31504 44280
<< metal5 >>
rect 24760 44280 25128 44304
rect 31160 44280 31528 44304
rect 20280 43960 24784 44280
rect 25104 43960 31184 44280
rect 31504 43960 31528 44280
rect 20280 43580 20600 43960
rect 24760 43936 25128 43960
rect 31160 43936 31528 43960
rect 1300 43556 20600 43580
rect 1300 43284 1324 43556
rect 1596 43284 20600 43556
rect 1300 43260 20600 43284
use controller_wrapper  controller_wrapper_0
timestamp 1758175872
transform 1 0 20468 0 1 900
box 0 496 11394 43900
use csdac255  dac_blue
timestamp 1758175872
transform -1 0 16648 0 1 1000
box -2130 0 14828 11424
use csdac255  dac_green
timestamp 1758175872
transform -1 0 16648 0 1 13714
box -2130 0 14828 11424
use csdac255  dac_red
timestamp 1758175872
transform -1 0 16648 0 1 26428
box -2130 0 14828 11424
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 600 90 0 0 clk
port 1 nsew
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 600 90 0 0 ena
port 2 nsew
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 600 90 0 0 rst_n
port 3 nsew
flabel metal4 s 30362 0 30542 200 0 FreeSans 1200 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 26498 0 26678 200 0 FreeSans 1200 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 22634 0 22814 200 0 FreeSans 1200 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 18770 0 18950 200 0 FreeSans 1200 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 14906 0 15086 200 0 FreeSans 1200 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 11042 0 11222 200 0 FreeSans 1200 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 7178 0 7358 200 0 FreeSans 1200 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 3314 0 3494 200 0 FreeSans 1200 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 600 90 0 0 ui_in[0]
port 12 nsew
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 600 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 600 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 600 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 600 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 600 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 600 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 600 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 600 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 600 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 600 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 600 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 600 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 600 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 600 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 600 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 600 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 600 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 600 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 600 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 600 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 600 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 600 90 0 0 uio_oe[6]
port 34 nsew
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 600 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 600 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 600 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 600 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 600 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 600 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 600 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 600 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 600 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 600 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 600 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 600 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 600 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 600 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 600 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 600 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 600 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 200 1000 920 44152 0 FreeSans 4000 90 0 0 VDPWR
port 52 nsew
flabel metal4 s 1120 1000 1840 44152 0 FreeSans 4000 90 0 0 VGND
port 53 nsew
flabel metal4 s 30524 1000 30844 44200 0 FreeSans 2000 90 0 0 VDPWR
port 52 nsew
flabel metal4 s 24124 1000 24444 44200 0 FreeSans 2000 90 0 0 VDPWR
port 52 nsew
flabel metal4 s 31184 1000 31504 44200 0 FreeSans 2000 90 0 0 VGND
port 53 nsew
flabel metal4 s 24784 1000 25104 44200 0 FreeSans 2000 90 0 0 VGND
port 53 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
string GDS_END 3814346
string GDS_FILE ../gds/tt_um_algofoogle_vga_matrix_dac.gds
string GDS_START 3732774
<< end >>
