* NGSPICE file created from csdac255_parax.ext - technology: sky130A

.subckt csdac255_parax Iout VPWR VGND Vbias data[0] data[1] data[2] data[3] data[4]
+ data[5] data[6] data[7] bias[0] bias[1] bias[2]
X0 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout VGND.t1612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1 VPWR.t1192 XThR.Tn[2].t12 XA.XIR[3].XIC[8].icell.PUM VPWR.t1191 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2 XA.XIR[12].XIC[10].icell.SM XA.XIR[12].XIC[10].icell.Ien Iout.t210 VGND.t1613 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X3 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t946 VPWR.t948 VPWR.t947 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X4 VGND.t1430 XA.Cn[10].t12 XA.XIR[4].XIC[10].icell.PDM VGND.t1429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X5 VGND.t2460 XThR.XTBN.Y a_n997_2667# VGND.t2422 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t953 XThR.Tn[6].t12 XA.XIR[7].XIC[8].icell.PUM VPWR.t952 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X7 XA.XIR[14].XIC[5].icell.Ien XThR.Tn[14].t12 VPWR.t203 VPWR.t202 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X8 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12].t12 XA.XIR[12].XIC[6].icell.Ien VGND.t296 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X9 XA.Cn[6].t7 thermo15c_0.XTBN.Y.t4 VGND.t1341 VGND.t1340 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1926 VGND.t2169 VGND.t2168 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X11 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[9].t12 VGND.t444 VGND.t443 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X12 VGND.t1342 thermo15c_0.XTBN.Y.t5 XA.Cn[5].t11 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 XA.XIR[15].XIC[9].icell.PUM XA.Cn[9].t12 XA.XIR[15].XIC[9].icell.Ien VPWR.t1246 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X14 XA.XIR[9].XIC[0].icell.SM XA.XIR[9].XIC[0].icell.Ien Iout.t216 VGND.t1783 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X15 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[12].t13 VGND.t298 VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X16 VGND.t2462 XA.Cn[11].t12 XA.XIR[12].XIC[11].icell.PDM VGND.t2461 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X17 XA.XIR[12].XIC[1].icell.SM XA.XIR[12].XIC[1].icell.Ien Iout.t167 VGND.t1366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X18 XA.XIR[8].XIC[12].icell.SM XA.XIR[8].XIC[12].icell.Ien Iout.t221 VGND.t1873 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X19 XA.Cn[12].t3 thermo15c_0.XTB5.Y VPWR.t343 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 XA.XIR[8].XIC_15.icell.PDM VPWR.t1927 VGND.t2171 VGND.t2170 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X21 XA.XIR[7].XIC[13].icell.SM XA.XIR[7].XIC[13].icell.Ien Iout.t169 VGND.t1368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X22 XA.XIR[14].XIC[13].icell.PUM XA.Cn[13].t12 XA.XIR[14].XIC[13].icell.Ien VPWR.t1326 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X23 a_2979_9615# thermo15c_0.XTBN.Y.t6 XA.Cn[0].t6 VPWR.t1325 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t944 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t945 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X25 XA.XIR[10].XIC[14].icell.SM XA.XIR[10].XIC[14].icell.Ien Iout.t207 VGND.t1520 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X26 a_4861_9615# thermo15c_0.XTB4.Y.t2 VPWR.t1300 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_5949_9615# thermo15c_0.XTBN.Y.t7 XA.Cn[5].t7 VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6].t13 XA.XIR[6].XIC[10].icell.Ien VGND.t776 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X29 XA.XIR[0].XIC[4].icell.PDM VGND.t1761 VGND.t1763 VGND.t1762 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X30 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[3].t12 VGND.t915 VGND.t914 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X31 XThR.Tn[5].t7 XThR.XTBN.Y a_n1049_5611# VPWR.t1771 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 XA.Cn[4].t3 thermo15c_0.XTB5.Y VGND.t416 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND.t2255 thermo15c_0.XTBN.Y.t8 XA.Cn[2].t5 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 XThR.XTB2.Y XThR.XTB6.A VPWR.t1662 VPWR.t1388 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[6].t14 VGND.t778 VGND.t777 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X36 XA.XIR[6].XIC[11].icell.SM XA.XIR[6].XIC[11].icell.Ien Iout.t168 VGND.t1367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X37 VGND.t830 XA.Cn[2].t12 XA.XIR[12].XIC[2].icell.PDM VGND.t829 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X38 VPWR.t943 VPWR.t941 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t942 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X39 VGND.t2173 VPWR.t1928 XA.XIR[7].XIC_dummy_left.icell.PDM VGND.t2172 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X40 VPWR.t1061 XThR.Tn[3].t13 XA.XIR[4].XIC[11].icell.PUM VPWR.t1060 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X41 VGND.t1272 Vbias.t6 XA.XIR[14].XIC[11].icell.SM VGND.t1271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X42 XA.XIR[2].XIC[1].icell.PUM XA.Cn[1].t12 XA.XIR[2].XIC[1].icell.Ien VPWR.t99 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X43 VGND.t2013 XA.Cn[3].t12 XA.XIR[15].XIC[3].icell.PDM VGND.t2012 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X44 VGND.t2175 VPWR.t1929 XA.XIR[10].XIC_15.icell.PDM VGND.t2174 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X45 VPWR.t1849 XThR.Tn[10].t12 XA.XIR[11].XIC[9].icell.PUM VPWR.t1848 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X46 XA.XIR[0].XIC[14].icell.PUM XA.Cn[14].t12 XA.XIR[0].XIC[14].icell.Ien VPWR.t1626 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X47 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t938 VPWR.t940 VPWR.t939 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X48 a_7651_9569# thermo15c_0.XTB1.Y.t3 XA.Cn[8].t7 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 VGND.t1274 Vbias.t7 XA.XIR[2].XIC[5].icell.SM VGND.t1273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X50 XA.XIR[1].XIC[6].icell.Ien XThR.Tn[1].t12 VPWR.t315 VPWR.t314 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X51 a_10051_9569# thermo15c_0.XTB6.Y XA.Cn[13].t7 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 VGND.t96 XA.Cn[4].t12 XA.XIR[2].XIC[4].icell.PDM VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X53 thermo15c_0.XTB5.Y thermo15c_0.XTB7.B VGND.t1104 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 XA.Cn[7].t3 thermo15c_0.XTBN.Y.t9 VPWR.t1758 VPWR.t1757 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X55 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[9].t13 VGND.t446 VGND.t445 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X56 VGND.t893 XThR.XTB7.Y XThR.Tn[6].t3 VGND.t892 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X57 XA.XIR[4].XIC[7].icell.Ien XThR.Tn[4].t12 VPWR.t1315 VPWR.t1314 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X58 VPWR.t1835 XThR.XTBN.Y XThR.Tn[9].t11 VPWR.t1822 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 XThR.XTB7.Y XThR.XTB7.A VGND.t1455 VGND.t1454 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 XA.XIR[3].XIC[8].icell.Ien XThR.Tn[3].t14 VPWR.t1409 VPWR.t1408 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X61 VPWR.t1411 XThR.Tn[3].t15 XA.XIR[4].XIC[2].icell.PUM VPWR.t1410 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X62 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[12].t14 VGND.t300 VGND.t299 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X63 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[1].t13 XA.XIR[1].XIC[9].icell.Ien VGND.t1809 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X64 VPWR.t1190 XThR.Tn[2].t13 XA.XIR[3].XIC[3].icell.PUM VPWR.t1189 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X65 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout VGND.t1117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X66 VPWR.t221 XThR.Tn[6].t15 XA.XIR[7].XIC[3].icell.PUM VPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X67 VPWR.t937 VPWR.t935 XA.XIR[2].XIC_15.icell.PUM VPWR.t936 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X68 a_6243_9615# thermo15c_0.XTB7.Y VPWR.t1354 VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X69 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11].t12 XA.XIR[11].XIC[14].icell.Ien VGND.t1820 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X70 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11].t13 XA.XIR[11].XIC[8].icell.Ien VGND.t1821 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X71 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[3].t16 VGND.t1509 VGND.t1508 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X72 XThR.Tn[7].t3 XThR.XTBN.Y VPWR.t1834 VPWR.t1833 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[0].t12 VGND.t845 VGND.t844 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X74 a_8963_9569# thermo15c_0.XTBN.Y.t10 VGND.t2256 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X75 VGND.t1276 Vbias.t8 XA.XIR[12].XIC[7].icell.SM VGND.t1275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X76 VGND.t500 XA.Cn[6].t12 XA.XIR[12].XIC[6].icell.PDM VGND.t499 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X77 XA.XIR[6].XIC[9].icell.SM XA.XIR[6].XIC[9].icell.Ien Iout.t70 VGND.t550 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X78 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout VGND.t1282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X79 XA.XIR[3].XIC[11].icell.SM XA.XIR[3].XIC[11].icell.Ien Iout.t139 VGND.t1084 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X80 VGND.t2177 VPWR.t1930 XA.XIR[4].XIC_dummy_left.icell.PDM VGND.t2176 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X81 VGND.t2459 XThR.XTBN.Y XThR.Tn[5].t11 VGND.t2442 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 VGND.t1278 Vbias.t9 XA.XIR[15].XIC[8].icell.SM VGND.t1277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X83 VGND.t1280 Vbias.t10 XA.XIR[14].XIC[9].icell.SM VGND.t1279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X84 VGND.t1019 XA.Cn[7].t8 XA.XIR[15].XIC[7].icell.PDM VGND.t1018 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X85 VGND.t2464 XA.Cn[11].t13 XA.XIR[6].XIC[11].icell.PDM VGND.t2463 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X86 VGND.t204 XA.Cn[1].t13 XA.XIR[3].XIC[1].icell.PDM VGND.t203 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X87 XA.XIR[4].XIC[11].icell.Ien XThR.Tn[4].t13 VPWR.t1317 VPWR.t1316 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X88 VPWR.t552 XThR.XTB6.Y a_n1049_5611# VPWR.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X89 XA.XIR[14].XIC[6].icell.PUM XA.Cn[6].t13 XA.XIR[14].XIC[6].icell.Ien VPWR.t422 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X90 VGND.t239 Vbias.t11 XA.XIR[9].XIC[7].icell.SM VGND.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X91 VGND.t832 XA.Cn[2].t13 XA.XIR[6].XIC[2].icell.PDM VGND.t831 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X92 XA.XIR[11].XIC[9].icell.Ien XThR.Tn[11].t14 VPWR.t1535 VPWR.t1534 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X93 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t1931 XA.XIR[6].XIC_dummy_left.icell.Ien VGND.t2178 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X94 VGND.t1270 Vbias.t3 Vbias.t4 VGND.t1269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X95 a_n1049_7787# XThR.XTB2.Y VPWR.t1670 VPWR.t1092 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X96 VGND.t1172 XA.Cn[9].t13 XA.XIR[14].XIC[9].icell.PDM VGND.t1171 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X97 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8].t12 XA.XIR[8].XIC[11].icell.Ien VGND.t1147 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X98 VGND.t241 Vbias.t12 XA.XIR[2].XIC[0].icell.SM VGND.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X99 XA.XIR[1].XIC[1].icell.Ien XThR.Tn[1].t14 VPWR.t1531 VPWR.t1530 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X100 XA.XIR[13].XIC[4].icell.PUM XA.Cn[4].t13 XA.XIR[13].XIC[4].icell.Ien VPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X101 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t933 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t934 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X102 VGND.t243 Vbias.t13 XA.XIR[0].XIC[13].icell.SM VGND.t242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X103 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[0].t13 VGND.t847 VGND.t846 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X104 XA.XIR[4].XIC[2].icell.Ien XThR.Tn[4].t14 VPWR.t1319 VPWR.t1318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X105 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[8].t13 VGND.t1149 VGND.t1148 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X106 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[8].t14 VGND.t1151 VGND.t1150 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X107 XA.XIR[3].XIC[3].icell.Ien XThR.Tn[3].t17 VPWR.t1413 VPWR.t1412 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X108 VGND.t2640 XA.Cn[12].t12 XA.XIR[0].XIC[12].icell.PDM VGND.t2639 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X109 VPWR.t1013 thermo15c_0.XTB3.Y.t3 a_4067_9615# VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[1].t15 XA.XIR[1].XIC[4].icell.Ien VGND.t1810 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X111 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5].t12 XA.XIR[5].XIC[1].icell.Ien VGND.t1614 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X112 VPWR.t456 data[4].t0 a_n1335_4229# VPWR.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X113 XA.XIR[2].XIC_15.icell.Ien XThR.Tn[2].t14 VPWR.t1188 VPWR.t1187 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X114 XA.XIR[3].XIC[9].icell.SM XA.XIR[3].XIC[9].icell.Ien Iout.t120 VGND.t1006 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X115 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9].t14 XA.XIR[9].XIC[1].icell.Ien VGND.t447 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X116 VGND.t2458 XThR.XTBN.Y XThR.Tn[7].t7 VGND.t2457 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X117 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[4].t15 XA.XIR[4].XIC[5].icell.Ien VGND.t1329 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X118 a_n1319_5317# XThR.XTB7.A VPWR.t1391 VPWR.t1390 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X119 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8].t15 XA.XIR[8].XIC[2].icell.Ien VGND.t902 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X120 VPWR.t104 XThR.Tn[13].t12 XA.XIR[14].XIC[14].icell.PUM VPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X121 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11].t15 XA.XIR[11].XIC[3].icell.Ien VGND.t1816 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X122 XA.XIR[7].XIC[8].icell.PUM XA.Cn[8].t12 XA.XIR[7].XIC[8].icell.Ien VPWR.t465 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X123 XA.Cn[9].t7 thermo15c_0.XTB2.Y VPWR.t1600 VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X124 XA.XIR[15].XIC[4].icell.Ien VPWR.t930 VPWR.t932 VPWR.t931 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X125 VGND.t245 Vbias.t14 XA.XIR[12].XIC[2].icell.SM VGND.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X126 XA.XIR[6].XIC[4].icell.SM XA.XIR[6].XIC[4].icell.Ien Iout.t39 VGND.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X127 VGND.t247 Vbias.t15 XA.XIR[11].XIC_15.icell.SM VGND.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X128 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t927 VPWR.t929 VPWR.t928 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X129 XA.Cn[5].t10 thermo15c_0.XTBN.Y.t11 VGND.t2257 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X130 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout VGND.t665 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X131 VGND.t249 Vbias.t16 XA.XIR[15].XIC[3].icell.SM VGND.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X132 VGND.t251 Vbias.t17 XA.XIR[14].XIC[4].icell.SM VGND.t250 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X133 VGND.t502 XA.Cn[6].t14 XA.XIR[6].XIC[6].icell.PDM VGND.t501 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X134 VPWR.t1039 XThR.Tn[8].t16 XA.XIR[9].XIC[4].icell.PUM VPWR.t1038 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X135 VPWR.t159 XThR.Tn[12].t15 XA.XIR[13].XIC[12].icell.PUM VPWR.t158 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X136 VGND.t1760 VGND.t1758 XA.XIR[13].XIC_dummy_right.icell.SM VGND.t1759 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X137 XThR.Tn[9].t3 XThR.XTB2.Y a_n997_3755# VGND.t1425 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X138 XA.Cn[0].t5 thermo15c_0.XTBN.Y.t12 a_2979_9615# VPWR.t1759 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X139 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1932 VGND.t2180 VGND.t2179 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X140 XA.Cn[5].t6 thermo15c_0.XTBN.Y.t13 a_5949_9615# VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X141 VGND.t415 thermo15c_0.XTB5.Y XA.Cn[4].t2 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X142 XA.XIR[14].XIC[1].icell.PUM XA.Cn[1].t14 XA.XIR[14].XIC[1].icell.Ien VPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X143 VGND.t253 Vbias.t18 XA.XIR[9].XIC[2].icell.SM VGND.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X144 a_9827_9569# thermo15c_0.XTB5.Y XA.Cn[12].t7 VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X145 XA.XIR[13].XIC[0].icell.PUM XA.Cn[0].t12 XA.XIR[13].XIC[0].icell.Ien VPWR.t1710 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X146 XA.Cn[7].t7 thermo15c_0.XTBN.Y.t14 VGND.t2259 VGND.t2258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X147 XA.Cn[2].t4 thermo15c_0.XTBN.Y.t15 VGND.t2260 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X148 VGND.t1432 XA.Cn[10].t13 XA.XIR[0].XIC[10].icell.PDM VGND.t1431 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X149 a_n997_1579# XThR.XTBN.Y VGND.t2456 VGND.t2440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X150 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[5].t13 VGND.t1616 VGND.t1615 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X151 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[5].t14 VGND.t1618 VGND.t1617 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X152 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t925 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t926 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X153 XA.XIR[9].XIC[14].icell.SM XA.XIR[9].XIC[14].icell.Ien Iout.t30 VGND.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X154 VGND.t98 XA.Cn[4].t14 XA.XIR[14].XIC[4].icell.PDM VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X155 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8].t17 XA.XIR[8].XIC[6].icell.Ien VGND.t903 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X156 XA.XIR[1].XIC[7].icell.PUM XA.Cn[7].t9 XA.XIR[1].XIC[7].icell.Ien VPWR.t1090 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X157 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[6].t16 VGND.t351 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X158 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[1].t16 VGND.t1812 VGND.t1811 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X159 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11].t16 XA.XIR[11].XIC[7].icell.Ien VGND.t1817 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X160 XA.XIR[4].XIC[8].icell.PUM XA.Cn[8].t13 XA.XIR[4].XIC[8].icell.Ien VPWR.t466 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X161 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[8].t18 VGND.t905 VGND.t904 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X162 XA.XIR[0].XIC_15.icell.SM XA.XIR[0].XIC_15.icell.Ien Iout.t116 VGND.t880 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X163 XA.XIR[4].XIC[12].icell.SM XA.XIR[4].XIC[12].icell.Ien Iout.t62 VGND.t397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X164 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[13].t13 VGND.t212 VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X165 XA.XIR[11].XIC[12].icell.PUM XA.Cn[12].t13 XA.XIR[11].XIC[12].icell.Ien VPWR.t1916 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X166 XA.XIR[12].XIC[4].icell.Ien XThR.Tn[12].t16 VPWR.t161 VPWR.t160 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X167 XA.XIR[3].XIC[4].icell.SM XA.XIR[3].XIC[4].icell.Ien Iout.t33 VGND.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X168 XA.XIR[15].XIC[0].icell.Ien VPWR.t922 VPWR.t924 VPWR.t923 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X169 VGND.t255 Vbias.t19 XA.XIR[8].XIC_15.icell.SM VGND.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X170 VGND.t1973 XA.Cn[14].t13 XA.XIR[8].XIC[14].icell.PDM VGND.t1972 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X171 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t919 VPWR.t921 VPWR.t920 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X172 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[4].t16 XA.XIR[4].XIC[0].icell.Ien VGND.t1330 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X173 VGND.t552 XA.Cn[8].t14 XA.XIR[8].XIC[8].icell.PDM VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X174 XA.XIR[14].XIC[14].icell.Ien XThR.Tn[14].t13 VPWR.t205 VPWR.t204 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X175 VGND.t2261 thermo15c_0.XTBN.Y.t16 XA.Cn[1].t7 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X176 VGND.t257 Vbias.t20 XA.XIR[1].XIC[5].icell.SM VGND.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X177 VPWR.t163 XThR.Tn[12].t17 XA.XIR[13].XIC[10].icell.PUM VPWR.t162 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X178 XA.XIR[7].XIC[3].icell.PUM XA.Cn[3].t13 XA.XIR[7].XIC[3].icell.Ien VPWR.t1675 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X179 XA.XIR[2].XIC_15.icell.PUM VPWR.t917 XA.XIR[2].XIC_15.icell.Ien VPWR.t918 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X180 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[2].t15 XA.XIR[2].XIC[13].icell.Ien VGND.t2473 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X181 VPWR.t373 XThR.Tn[9].t15 XA.XIR[10].XIC[12].icell.PUM VPWR.t372 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X182 VPWR.t1041 XThR.Tn[8].t19 XA.XIR[9].XIC[0].icell.PUM VPWR.t1040 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X183 VGND.t259 Vbias.t21 XA.XIR[4].XIC[6].icell.SM VGND.t258 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X184 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1933 VGND.t2182 VGND.t2181 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X185 VPWR.t916 VPWR.t914 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t915 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X186 VPWR.t1760 thermo15c_0.XTBN.Y.t17 XA.Cn[10].t11 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X187 VGND.t2455 XThR.XTBN.Y XThR.Tn[3].t11 VGND.t2418 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X188 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[2].t16 VGND.t2472 VGND.t2471 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X189 XA.XIR[6].XIC[8].icell.Ien XThR.Tn[6].t17 VPWR.t223 VPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X190 XThR.Tn[0].t7 XThR.XTBN.Y a_n1049_8581# VPWR.t1832 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X191 XA.XIR[13].XIC[12].icell.Ien XThR.Tn[13].t14 VPWR.t106 VPWR.t105 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X192 XA.XIR[13].XIC[7].icell.SM XA.XIR[13].XIC[7].icell.Ien Iout.t92 VGND.t740 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X193 VPWR.t1479 VGND.t2688 XA.XIR[0].XIC[8].icell.PUM VPWR.t1478 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X194 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10].t13 XA.XIR[10].XIC[14].icell.Ien VGND.t2489 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X195 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10].t14 XA.XIR[10].XIC[8].icell.Ien VGND.t2490 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X196 XA.Cn[12].t2 thermo15c_0.XTB5.Y VPWR.t342 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 XA.XIR[1].XIC[11].icell.PUM XA.Cn[11].t14 XA.XIR[1].XIC[11].icell.Ien VPWR.t997 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X198 XThR.Tn[11].t11 XThR.XTBN.Y VPWR.t1831 VPWR.t1820 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 XA.XIR[0].XIC[7].icell.Ien XThR.Tn[0].t14 VPWR.t996 VPWR.t995 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X200 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[2].t17 VGND.t2470 VGND.t2469 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X201 XA.XIR[8].XIC[9].icell.PUM XA.Cn[9].t14 XA.XIR[8].XIC[9].icell.Ien VPWR.t1247 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X202 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[8].t20 VGND.t907 VGND.t906 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X203 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout VGND.t1116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X204 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[5].t15 VGND.t1620 VGND.t1619 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X205 VGND.t849 XA.Cn[11].t15 XA.XIR[5].XIC[11].icell.PDM VGND.t848 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X206 XA.XIR[11].XIC[10].icell.PUM XA.Cn[10].t14 XA.XIR[11].XIC[10].icell.Ien VPWR.t1377 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X207 XThR.Tn[2].t11 XThR.XTBN.Y VGND.t2454 VGND.t2407 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X208 VGND.t851 XA.Cn[11].t16 XA.XIR[9].XIC[11].icell.PDM VGND.t850 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X209 VGND.t1757 VGND.t1755 XA.XIR[13].XIC_dummy_left.icell.SM VGND.t1756 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X210 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12].t18 VPWR.t165 VPWR.t164 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X211 XA.XIR[1].XIC[2].icell.PUM XA.Cn[2].t14 XA.XIR[1].XIC[2].icell.Ien VPWR.t980 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X212 VPWR.t1830 XThR.XTBN.Y XThR.Tn[12].t11 VPWR.t1781 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X213 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[1].t17 VGND.t1814 VGND.t1813 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X214 thermo15c_0.XTB7.A data[0].t0 VPWR.t949 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X215 VPWR.t375 XThR.Tn[9].t16 XA.XIR[10].XIC[10].icell.PUM VPWR.t374 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X216 XA.XIR[4].XIC[3].icell.PUM XA.Cn[3].t14 XA.XIR[4].XIC[3].icell.Ien VPWR.t1676 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X217 VGND.t261 Vbias.t22 XA.XIR[4].XIC[10].icell.SM VGND.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X218 XA.XIR[0].XIC[13].icell.PDM VGND.t1752 VGND.t1754 VGND.t1753 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X219 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[13].t15 VGND.t1124 VGND.t1123 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X220 VGND.t2184 VPWR.t1934 XA.XIR[0].XIC_dummy_left.icell.PDM VGND.t2183 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X221 VGND.t834 XA.Cn[2].t15 XA.XIR[5].XIC[2].icell.PDM VGND.t833 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X222 VGND.t2563 Vbias.t23 XA.XIR[11].XIC[8].icell.SM VGND.t2562 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X223 XA.Cn[9].t11 thermo15c_0.XTB2.Y a_7875_9569# VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X224 VGND.t1601 XA.Cn[5].t12 XA.XIR[1].XIC[5].icell.PDM VGND.t1600 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X225 XA.XIR[10].XIC[9].icell.Ien XThR.Tn[10].t15 VPWR.t1851 VPWR.t1850 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X226 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1935 VGND.t2186 VGND.t2185 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X227 VGND.t836 XA.Cn[2].t16 XA.XIR[9].XIC[2].icell.PDM VGND.t835 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X228 VGND.t2015 XA.Cn[3].t15 XA.XIR[8].XIC[3].icell.PDM VGND.t2014 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X229 VGND.t2188 VPWR.t1936 XA.XIR[3].XIC_15.icell.PDM VGND.t2187 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X230 a_n1319_5611# XThR.XTB6.A VPWR.t1661 VPWR.t1390 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X231 XA.XIR[13].XIC[10].icell.Ien XThR.Tn[13].t16 VPWR.t1201 VPWR.t1200 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X232 VGND.t2453 XThR.XTBN.Y a_n997_3979# VGND.t2369 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X233 XA.XIR[15].XIC_15.icell.SM XA.XIR[15].XIC_15.icell.Ien Iout.t222 VGND.t1936 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X234 VPWR.t1761 thermo15c_0.XTBN.Y.t18 XA.Cn[14].t3 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X235 VGND.t2565 Vbias.t24 XA.XIR[1].XIC[0].icell.SM VGND.t2564 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X236 VPWR.t167 XThR.Tn[12].t19 XA.XIR[13].XIC[5].icell.PUM VPWR.t166 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X237 XA.XIR[12].XIC[4].icell.PUM XA.Cn[4].t15 XA.XIR[12].XIC[4].icell.Ien VPWR.t31 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X238 VGND.t2567 Vbias.t25 XA.XIR[4].XIC[1].icell.SM VGND.t2566 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X239 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7].t8 XA.XIR[7].XIC[14].icell.Ien VGND.t682 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X240 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7].t9 XA.XIR[7].XIC[8].icell.Ien VGND.t683 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X241 XA.XIR[0].XIC[11].icell.Ien XThR.Tn[0].t15 VPWR.t1616 VPWR.t1615 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X242 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[2].t18 VGND.t2468 VGND.t2467 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X243 XA.XIR[6].XIC[3].icell.Ien XThR.Tn[6].t18 VPWR.t225 VPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X244 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14].t14 XA.XIR[14].XIC[12].icell.Ien VGND.t341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X245 XA.XIR[11].XIC[6].icell.SM XA.XIR[11].XIC[6].icell.Ien Iout.t130 VGND.t1046 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X246 XA.XIR[1].XIC_15.icell.Ien XThR.Tn[1].t18 VPWR.t1533 VPWR.t1532 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X247 VGND.t2569 Vbias.t26 XA.XIR[2].XIC[14].icell.SM VGND.t2568 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X248 VGND.t1344 XA.Cn[13].t13 XA.XIR[2].XIC[13].icell.PDM VGND.t1343 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X249 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[5].t16 VGND.t1622 VGND.t1621 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X250 VPWR.t1488 XThR.XTB4.Y.t2 a_n1049_6699# VPWR.t1240 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X251 VGND.t2190 VPWR.t1937 XA.XIR[15].XIC_dummy_right.icell.PDM VGND.t2189 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X252 XA.XIR[13].XIC[2].icell.SM XA.XIR[13].XIC[2].icell.Ien Iout.t142 VGND.t1106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X253 VPWR.t1477 VGND.t2689 XA.XIR[0].XIC[3].icell.PUM VPWR.t1476 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X254 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10].t16 XA.XIR[10].XIC[3].icell.Ien VGND.t2491 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X255 VPWR.t1037 thermo15c_0.XTB6.Y a_5949_9615# VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X256 VPWR.t1376 XThR.XTB1.Y a_n1049_8581# VPWR.t1375 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X257 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5].t17 XA.XIR[5].XIC_15.icell.Ien VGND.t1770 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X258 VPWR.t1537 XThR.Tn[11].t17 XA.XIR[12].XIC[7].icell.PUM VPWR.t1536 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X259 XA.XIR[0].XIC[2].icell.Ien XThR.Tn[0].t16 VPWR.t1618 VPWR.t1617 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X260 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9].t17 XA.XIR[9].XIC_15.icell.Ien VGND.t448 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X261 XA.XIR[0].XIC[8].icell.SM XA.XIR[0].XIC[8].icell.Ien Iout.t90 VGND.t738 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X262 VGND.t2571 Vbias.t27 XA.XIR[5].XIC[7].icell.SM VGND.t2570 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X263 XA.XIR[11].XIC[5].icell.PUM XA.Cn[5].t13 XA.XIR[11].XIC[5].icell.Ien VPWR.t1436 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X264 VGND.t504 XA.Cn[6].t15 XA.XIR[5].XIC[6].icell.PDM VGND.t503 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X265 VGND.t1139 XThR.XTB7.B a_n1335_8107# VGND.t1133 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X266 VPWR.t500 XThR.Tn[7].t10 XA.XIR[8].XIC[4].icell.PUM VPWR.t499 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X267 XA.XIR[0].XIC[5].icell.PDM XThR.Tn[0].t17 XA.XIR[0].XIC[5].icell.Ien VGND.t1959 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X268 VPWR.t913 VPWR.t911 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t912 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X269 VGND.t506 XA.Cn[6].t16 XA.XIR[9].XIC[6].icell.PDM VGND.t505 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X270 VGND.t2573 Vbias.t28 XA.XIR[8].XIC[8].icell.SM VGND.t2572 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X271 XA.XIR[7].XIC[9].icell.Ien XThR.Tn[7].t11 VPWR.t502 VPWR.t501 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X272 thermo15c_0.XTB4.Y.t0 thermo15c_0.XTB7.B VPWR.t1130 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X273 VGND.t1751 VGND.t1749 XA.XIR[12].XIC_dummy_right.icell.SM VGND.t1750 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X274 VGND.t1021 XA.Cn[7].t10 XA.XIR[8].XIC[7].icell.PDM VGND.t1020 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X275 VPWR.t910 VPWR.t908 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t909 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X276 XThR.Tn[2].t2 XThR.XTB3.Y.t3 VGND.t1030 VGND.t1029 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X277 VGND.t2450 XThR.XTBN.Y a_n997_2891# VGND.t2403 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X278 VPWR.t436 XThR.Tn[9].t18 XA.XIR[10].XIC[5].icell.PUM VPWR.t435 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X279 XA.XIR[5].XIC[5].icell.SM XA.XIR[5].XIC[5].icell.Ien Iout.t214 VGND.t1781 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X280 VPWR.t1243 XThR.XTB5.Y XThR.Tn[12].t7 VPWR.t1242 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X281 XA.XIR[12].XIC[0].icell.PUM XA.Cn[0].t13 XA.XIR[12].XIC[0].icell.Ien VPWR.t1711 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X282 VGND.t1925 XA.Cn[0].t14 XA.XIR[1].XIC[0].icell.PDM VGND.t1924 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X283 VGND.t2575 Vbias.t29 XA.XIR[11].XIC[3].icell.SM VGND.t2574 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X284 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14].t15 XA.XIR[14].XIC[10].icell.Ien VGND.t342 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X285 XA.XIR[11].XIC[10].icell.SM XA.XIR[11].XIC[10].icell.Ien Iout.t242 VGND.t2162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X286 VGND.t2452 XThR.XTBN.Y XThR.Tn[6].t11 VGND.t2451 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X287 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[11].t18 VGND.t1819 VGND.t1818 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X288 VPWR.t1829 XThR.XTBN.Y XThR.Tn[9].t10 VPWR.t1815 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X289 XA.XIR[8].XIC[6].icell.SM XA.XIR[8].XIC[6].icell.Ien Iout.t172 VGND.t1371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X290 XA.XIR[13].XIC[5].icell.Ien XThR.Tn[13].t17 VPWR.t1203 VPWR.t1202 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X291 VGND.t1748 VGND.t1746 XA.XIR[9].XIC_dummy_right.icell.SM VGND.t1747 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X292 XA.XIR[14].XIC_15.icell.PUM VPWR.t906 XA.XIR[14].XIC_15.icell.Ien VPWR.t907 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X293 a_n997_715# XThR.XTBN.Y VGND.t2449 VGND.t2448 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X294 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10].t17 XA.XIR[10].XIC[7].icell.Ien VGND.t2492 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X295 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7].t12 XA.XIR[7].XIC[3].icell.Ien VGND.t684 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X296 XA.Cn[1].t6 thermo15c_0.XTBN.Y.t19 VGND.t392 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X297 VPWR.t1539 XThR.Tn[11].t19 XA.XIR[12].XIC[11].icell.PUM VPWR.t1538 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X298 XA.XIR[6].XIC[4].icell.PUM XA.Cn[4].t16 XA.XIR[6].XIC[4].icell.Ien VPWR.t32 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X299 XThR.Tn[14].t3 XThR.XTB7.Y VPWR.t1022 VPWR.t537 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X300 XA.XIR[10].XIC[12].icell.PUM XA.Cn[12].t14 XA.XIR[10].XIC[12].icell.Ien VPWR.t1917 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X301 XA.XIR[2].XIC[5].icell.SM XA.XIR[2].XIC[5].icell.Ien Iout.t95 VGND.t743 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X302 XA.XIR[11].XIC[1].icell.SM XA.XIR[11].XIC[1].icell.Ien Iout.t148 VGND.t1120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X303 XA.XIR[7].XIC_15.icell.PDM VPWR.t1938 VGND.t2192 VGND.t2191 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X304 XA.XIR[6].XIC[13].icell.SM XA.XIR[6].XIC[13].icell.Ien Iout.t51 VGND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X305 XA.XIR[13].XIC[13].icell.PUM XA.Cn[13].t14 XA.XIR[13].XIC[13].icell.Ien VPWR.t1327 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X306 VGND.t2577 Vbias.t30 XA.XIR[15].XIC[12].icell.SM VGND.t2576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X307 VGND.t2579 Vbias.t31 XA.XIR[14].XIC[13].icell.SM VGND.t2578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X308 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[2].t19 XA.XIR[2].XIC[1].icell.Ien VGND.t2466 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X309 VPWR.t273 XThR.Tn[7].t13 XA.XIR[8].XIC[0].icell.PUM VPWR.t272 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X310 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[1].t19 XA.XIR[1].XIC[13].icell.Ien VGND.t1815 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X311 VPWR.t1241 XThR.XTB5.Y a_n1049_6405# VPWR.t1240 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X312 VPWR.t1541 XThR.Tn[11].t20 XA.XIR[12].XIC[2].icell.PUM VPWR.t1540 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X313 XThR.XTB7.B data[6].t0 VPWR.t1012 VPWR.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X314 XA.XIR[0].XIC[8].icell.PUM XA.Cn[8].t15 XA.XIR[0].XIC[8].icell.Ien VPWR.t467 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X315 VPWR.t1301 thermo15c_0.XTB4.Y.t3 a_4861_9615# VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X316 XA.XIR[0].XIC[3].icell.SM XA.XIR[0].XIC[3].icell.Ien Iout.t201 VGND.t1504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X317 VGND.t2581 Vbias.t32 XA.XIR[5].XIC[2].icell.SM VGND.t2580 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X318 XA.XIR[8].XIC[4].icell.Ien XThR.Tn[8].t21 VPWR.t1043 VPWR.t1042 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X319 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t903 VPWR.t905 VPWR.t904 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X320 VGND.t2002 XThR.XTB2.Y XThR.Tn[1].t3 VGND.t1418 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X321 XA.XIR[0].XIC[0].icell.PDM XThR.Tn[0].t18 XA.XIR[0].XIC[0].icell.Ien VGND.t1960 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X322 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[11].t21 VGND.t2478 VGND.t2477 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X323 XA.XIR[12].XIC[7].icell.SM XA.XIR[12].XIC[7].icell.Ien Iout.t82 VGND.t669 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X324 XThR.XTB7.A data[4].t1 a_n1331_2891# VGND.t540 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X325 XA.XIR[8].XIC[10].icell.SM XA.XIR[8].XIC[10].icell.Ien Iout.t218 VGND.t1785 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X326 VGND.t2583 Vbias.t33 XA.XIR[8].XIC[3].icell.SM VGND.t2582 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X327 XA.XIR[15].XIC[13].icell.Ien VPWR.t900 VPWR.t902 VPWR.t901 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X328 XA.XIR[15].XIC[8].icell.SM XA.XIR[15].XIC[8].icell.Ien Iout.t106 VGND.t824 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X329 VPWR.t1493 XThR.Tn[5].t18 XA.XIR[6].XIC[12].icell.PUM VPWR.t1492 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X330 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1939 XA.XIR[11].XIC_dummy_right.icell.Ien VGND.t2193 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X331 VPWR.t317 XThR.Tn[8].t22 XA.XIR[9].XIC[13].icell.PUM VPWR.t316 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X332 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7].t14 XA.XIR[7].XIC[7].icell.Ien VGND.t378 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X333 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t7 VPWR.t1814 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X334 XA.XIR[5].XIC[0].icell.SM XA.XIR[5].XIC[0].icell.Ien Iout.t252 VGND.t2628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X335 XA.XIR[10].XIC[10].icell.PUM XA.Cn[10].t15 XA.XIR[10].XIC[10].icell.Ien VPWR.t1378 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X336 VGND.t393 thermo15c_0.XTBN.Y.t20 XA.Cn[4].t11 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X337 XA.XIR[6].XIC[0].icell.PUM XA.Cn[0].t15 XA.XIR[6].XIC[0].icell.Ien VPWR.t1587 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X338 XA.XIR[8].XIC[1].icell.SM XA.XIR[8].XIC[1].icell.Ien Iout.t243 VGND.t2364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X339 XA.XIR[3].XIC[13].icell.SM XA.XIR[3].XIC[13].icell.Ien Iout.t3 VGND.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X340 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t898 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t899 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X341 VGND.t1745 VGND.t1743 XA.XIR[12].XIC_dummy_left.icell.SM VGND.t1744 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X342 thermo15c_0.XTB5.A data[1].t0 a_7331_10587# VPWR.t524 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X343 VGND.t714 data[1].t1 a_8739_10571# VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X344 XA.XIR[0].XIC[1].icell.PDM VGND.t1740 VGND.t1742 VGND.t1741 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X345 VPWR.t1669 XThR.XTB2.Y XThR.Tn[9].t7 VPWR.t1244 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X346 VGND.t2447 XThR.XTBN.Y XThR.Tn[7].t6 VGND.t2446 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X347 VGND.t1346 XA.Cn[13].t15 XA.XIR[14].XIC[13].icell.PDM VGND.t1345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X348 XA.XIR[2].XIC[0].icell.SM XA.XIR[2].XIC[0].icell.Ien Iout.t197 VGND.t1499 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X349 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1940 XA.XIR[14].XIC_dummy_left.icell.Ien VGND.t2194 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X350 XThR.Tn[13].t11 XThR.XTBN.Y VPWR.t1828 VPWR.t1791 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X351 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[10].t18 VGND.t1089 VGND.t1088 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X352 XA.XIR[14].XIC_15.icell.SM XA.XIR[14].XIC_15.icell.Ien Iout.t138 VGND.t1083 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X353 VGND.t2585 Vbias.t34 XA.XIR[10].XIC[11].icell.SM VGND.t2584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X354 VGND.t1739 VGND.t1737 XA.XIR[9].XIC_dummy_left.icell.SM VGND.t1738 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X355 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8].t23 VPWR.t319 VPWR.t318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X356 VPWR.t1186 XThR.Tn[2].t20 XA.XIR[3].XIC[9].icell.PUM VPWR.t1185 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X357 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t895 VPWR.t897 VPWR.t896 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X358 XA.XIR[12].XIC[13].icell.Ien XThR.Tn[12].t20 VPWR.t171 VPWR.t170 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X359 VPWR.t227 XThR.Tn[6].t19 XA.XIR[7].XIC[9].icell.PUM VPWR.t226 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X360 XA.XIR[0].XIC[3].icell.PUM XA.Cn[3].t16 XA.XIR[0].XIC[3].icell.Ien VPWR.t1677 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X361 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t892 VPWR.t894 VPWR.t893 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X362 VPWR.t1495 XThR.Tn[5].t19 XA.XIR[6].XIC[10].icell.PUM VPWR.t1494 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X363 VGND.t206 XA.Cn[1].t15 XA.XIR[2].XIC[1].icell.PDM VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X364 VGND.t756 XThR.XTB6.Y XThR.Tn[5].t3 VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X365 XA.XIR[13].XIC[6].icell.PUM XA.Cn[6].t17 XA.XIR[13].XIC[6].icell.Ien VPWR.t423 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X366 XThR.Tn[9].t2 XThR.XTB2.Y a_n997_3755# VGND.t1422 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X367 VGND.t983 Vbias.t35 XA.XIR[1].XIC[14].icell.SM VGND.t982 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X368 XThR.XTB6.Y XThR.XTB6.A VGND.t1998 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X369 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t1941 VGND.t2196 VGND.t2195 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X370 XA.XIR[12].XIC[2].icell.SM XA.XIR[12].XIC[2].icell.Ien Iout.t245 VGND.t2475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X371 a_n997_1579# XThR.XTBN.Y VGND.t2445 VGND.t2435 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X372 VGND.t1174 XA.Cn[9].t15 XA.XIR[13].XIC[9].icell.PDM VGND.t1173 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X373 XA.XIR[15].XIC[3].icell.SM XA.XIR[15].XIC[3].icell.Ien Iout.t56 VGND.t199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X374 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[3].t18 XA.XIR[3].XIC[14].icell.Ien VGND.t1510 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X375 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[3].t19 XA.XIR[3].XIC[8].icell.Ien VGND.t1511 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X376 VPWR.t207 XThR.Tn[14].t16 XA.XIR[15].XIC[7].icell.PUM VPWR.t206 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X377 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t890 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t891 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X378 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout VGND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X379 VPWR.t1205 XThR.Tn[13].t18 XA.XIR[14].XIC[8].icell.PUM VPWR.t1204 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X380 XA.XIR[10].XIC[5].icell.PUM XA.Cn[5].t14 XA.XIR[10].XIC[5].icell.Ien VPWR.t1437 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X381 XA.XIR[15].XIC[6].icell.Ien VPWR.t887 VPWR.t889 VPWR.t888 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X382 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t1942 VGND.t2198 VGND.t2197 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X383 VGND.t985 Vbias.t36 XA.XIR[10].XIC[9].icell.SM VGND.t984 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X384 VPWR.t173 XThR.Tn[12].t21 XA.XIR[13].XIC[14].icell.PUM VPWR.t172 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X385 VPWR.t321 XThR.Tn[8].t24 XA.XIR[9].XIC[6].icell.PUM VPWR.t320 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X386 XA.XIR[15].XIC[9].icell.PDM VPWR.t1943 XA.XIR[15].XIC[9].icell.Ien VGND.t2199 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X387 XA.XIR[3].XIC[9].icell.Ien XThR.Tn[3].t20 VPWR.t1415 VPWR.t1414 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X388 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[10].t19 VGND.t1091 VGND.t1090 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X389 XA.XIR[15].XIC[12].icell.PDM XThR.Tn[14].t17 VGND.t344 VGND.t343 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X390 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1944 VGND.t2201 VGND.t2200 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X391 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[13].t19 VGND.t1126 VGND.t1125 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X392 VPWR.t1894 XThR.XTBN.A XThR.XTBN.Y VPWR.t1893 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X393 VPWR.t1497 XThR.Tn[5].t20 XA.XIR[6].XIC[5].icell.PUM VPWR.t1496 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X394 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[4].t17 XA.XIR[4].XIC[11].icell.Ien VGND.t1331 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X395 XA.XIR[5].XIC[4].icell.PUM XA.Cn[4].t17 XA.XIR[5].XIC[4].icell.Ien VPWR.t33 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X396 VPWR.t209 XThR.Tn[14].t18 XA.XIR[15].XIC[11].icell.PUM VPWR.t208 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X397 XA.XIR[1].XIC[5].icell.SM XA.XIR[1].XIC[5].icell.Ien Iout.t87 VGND.t716 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X398 XA.XIR[13].XIC[1].icell.PUM XA.Cn[1].t16 XA.XIR[13].XIC[1].icell.Ien VPWR.t101 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X399 XA.XIR[9].XIC[4].icell.PUM XA.Cn[4].t18 XA.XIR[9].XIC[4].icell.Ien VPWR.t34 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X400 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t885 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t886 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X401 a_3523_10575# thermo15c_0.XTB7.B VGND.t1103 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X402 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[4].t18 VGND.t1802 VGND.t1801 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X403 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[4].t19 VGND.t1804 VGND.t1803 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X404 XA.XIR[12].XIC[13].icell.PUM XA.Cn[13].t16 XA.XIR[12].XIC[13].icell.Ien VPWR.t1328 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X405 XA.XIR[4].XIC[6].icell.SM XA.XIR[4].XIC[6].icell.Ien Iout.t255 VGND.t2687 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X406 XA.XIR[11].XIC[14].icell.PUM XA.Cn[14].t14 XA.XIR[11].XIC[14].icell.Ien VPWR.t81 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X407 VPWR.t301 thermo15c_0.XTBN.Y.t21 XA.Cn[13].t11 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[1].t20 XA.XIR[1].XIC[1].icell.Ien VGND.t699 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X409 VGND.t987 Vbias.t37 XA.XIR[13].XIC[5].icell.SM VGND.t986 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X410 VGND.t100 XA.Cn[4].t19 XA.XIR[13].XIC[4].icell.PDM VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X411 XA.XIR[12].XIC[6].icell.Ien XThR.Tn[12].t22 VPWR.t175 VPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X412 XA.Cn[5].t3 thermo15c_0.XTB6.Y VGND.t900 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 XA.Cn[4].t1 thermo15c_0.XTB5.Y VGND.t414 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X414 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[4].t20 XA.XIR[4].XIC[2].icell.Ien VGND.t1805 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X415 VGND.t2203 VPWR.t1945 XA.XIR[8].XIC_dummy_right.icell.PDM VGND.t2202 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X416 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[3].t21 XA.XIR[3].XIC[3].icell.Ien VGND.t1512 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X417 XA.XIR[14].XIC[8].icell.Ien XThR.Tn[14].t19 VPWR.t185 VPWR.t184 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X418 VPWR.t187 XThR.Tn[14].t20 XA.XIR[15].XIC[2].icell.PUM VPWR.t186 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X419 XA.XIR[2].XIC_15.icell.PDM XThR.Tn[2].t21 XA.XIR[2].XIC_15.icell.Ien VGND.t2602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X420 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t7 VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X421 VPWR.t1207 XThR.Tn[13].t20 XA.XIR[14].XIC[3].icell.PUM VPWR.t1206 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X422 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12].t23 XA.XIR[12].XIC[9].icell.Ien VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X423 VPWR.t438 XThR.Tn[9].t19 XA.XIR[10].XIC[14].icell.PUM VPWR.t437 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X424 XA.XIR[15].XIC[1].icell.Ien VPWR.t879 VPWR.t881 VPWR.t880 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X425 VGND.t989 Vbias.t38 XA.XIR[11].XIC[12].icell.SM VGND.t988 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X426 VGND.t991 Vbias.t39 XA.XIR[7].XIC_15.icell.SM VGND.t990 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X427 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t882 VPWR.t884 VPWR.t883 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X428 VGND.t166 XA.Cn[14].t15 XA.XIR[7].XIC[14].icell.PDM VGND.t165 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X429 VGND.t554 XA.Cn[8].t16 XA.XIR[7].XIC[8].icell.PDM VGND.t553 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X430 a_7875_9569# thermo15c_0.XTB2.Y XA.Cn[9].t10 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X431 XA.Cn[4].t10 thermo15c_0.XTBN.Y.t22 VGND.t394 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X432 VPWR.t1620 XThR.Tn[0].t19 XA.XIR[1].XIC[4].icell.PUM VPWR.t1619 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X433 a_n1049_5317# XThR.XTB7.Y VPWR.t1021 VPWR.t549 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X434 XA.XIR[13].XIC[14].icell.Ien XThR.Tn[13].t21 VPWR.t1582 VPWR.t1581 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X435 XA.XIR[14].XIC[8].icell.SM XA.XIR[14].XIC[8].icell.Ien Iout.t0 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X436 XA.XIR[15].XIC[10].icell.PDM XThR.Tn[14].t21 VGND.t318 VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X437 VGND.t993 Vbias.t40 XA.XIR[10].XIC[4].icell.SM VGND.t992 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X438 VGND.t1736 VGND.t1734 XA.XIR[5].XIC_dummy_right.icell.SM VGND.t1735 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X439 VPWR.t323 XThR.Tn[8].t25 XA.XIR[9].XIC[1].icell.PUM VPWR.t322 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X440 VPWR.t1527 XThR.Tn[4].t21 XA.XIR[5].XIC[4].icell.PUM VPWR.t1526 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X441 thermo15c_0.XTB6.Y thermo15c_0.XTB7.B VGND.t1102 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X442 VPWR.t878 VPWR.t876 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t877 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X443 XA.XIR[15].XIC[4].icell.PDM VPWR.t1946 XA.XIR[15].XIC[4].icell.Ien VGND.t2204 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X444 VPWR.t275 XThR.Tn[7].t15 XA.XIR[8].XIC[13].icell.PUM VPWR.t274 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X445 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t1947 XA.XIR[10].XIC_dummy_right.icell.Ien VGND.t2205 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X446 a_6243_9615# thermo15c_0.XTBN.Y.t23 XA.Cn[6].t3 VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X447 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout VGND.t668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X448 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[1].t21 VGND.t701 VGND.t700 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X449 XA.XIR[5].XIC[0].icell.PUM XA.Cn[0].t16 XA.XIR[5].XIC[0].icell.Ien VPWR.t1588 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X450 XA.XIR[4].XIC[10].icell.SM XA.XIR[4].XIC[10].icell.Ien Iout.t8 VGND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X451 XA.XIR[9].XIC[0].icell.PUM XA.Cn[0].t17 XA.XIR[9].XIC[0].icell.Ien VPWR.t1589 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X452 XA.Cn[13].t3 thermo15c_0.XTB6.Y VPWR.t1036 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X453 XA.XIR[5].XIC[14].icell.SM XA.XIR[5].XIC[14].icell.Ien Iout.t20 VGND.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X454 VGND.t395 thermo15c_0.XTBN.Y.t24 XA.Cn[0].t10 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X455 XThR.Tn[3].t7 XThR.XTBN.Y a_n1049_6699# VPWR.t1827 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X456 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[4].t22 XA.XIR[4].XIC[6].icell.Ien VGND.t1806 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X457 VGND.t208 XA.Cn[1].t17 XA.XIR[14].XIC[1].icell.PDM VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X458 VGND.t1769 XThR.XTB4.Y.t3 XThR.Tn[3].t3 VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X459 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[3].t22 XA.XIR[3].XIC[7].icell.Ien VGND.t1513 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X460 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[1].t22 VGND.t703 VGND.t702 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X461 XA.XIR[7].XIC[9].icell.PUM XA.Cn[9].t16 XA.XIR[7].XIC[9].icell.Ien VPWR.t1248 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X462 XA.XIR[1].XIC[0].icell.SM XA.XIR[1].XIC[0].icell.Ien Iout.t128 VGND.t1035 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X463 XA.XIR[3].XIC[12].icell.PUM XA.Cn[12].t15 XA.XIR[3].XIC[12].icell.Ien VPWR.t1918 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X464 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[4].t23 VGND.t1808 VGND.t1807 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X465 XA.XIR[0].XIC[12].icell.SM XA.XIR[0].XIC[12].icell.Ien Iout.t55 VGND.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X466 XA.XIR[0].XIC_15.icell.PDM VPWR.t1948 VGND.t2207 VGND.t2206 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X467 XA.XIR[4].XIC[1].icell.SM XA.XIR[4].XIC[1].icell.Ien Iout.t31 VGND.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X468 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[9].t20 VGND.t526 VGND.t525 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X469 VGND.t995 Vbias.t41 XA.XIR[13].XIC[0].icell.SM VGND.t994 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X470 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12].t24 VPWR.t177 VPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X471 XA.XIR[6].XIC[13].icell.PUM XA.Cn[13].t17 XA.XIR[6].XIC[13].icell.Ien VPWR.t1329 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X472 VGND.t997 Vbias.t42 XA.XIR[8].XIC[12].icell.SM VGND.t996 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X473 XA.XIR[2].XIC[14].icell.SM XA.XIR[2].XIC[14].icell.Ien Iout.t89 VGND.t737 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X474 XThR.Tn[11].t6 XThR.XTB4.Y.t4 VPWR.t1489 VPWR.t1234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X475 VGND.t1050 XA.Cn[8].t17 XA.XIR[4].XIC[8].icell.PDM VGND.t1049 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X476 VGND.t168 XA.Cn[14].t16 XA.XIR[4].XIC[14].icell.PDM VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X477 XA.Cn[14].t11 thermo15c_0.XTB7.Y a_10915_9569# VGND.t1400 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X478 VPWR.t1622 XThR.Tn[0].t20 XA.XIR[1].XIC[0].icell.PUM VPWR.t1621 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X479 XA.XIR[14].XIC[3].icell.Ien XThR.Tn[14].t22 VPWR.t189 VPWR.t188 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X480 VGND.t2642 XA.Cn[12].t16 XA.XIR[11].XIC[12].icell.PDM VGND.t2641 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X481 VPWR.t1529 XThR.Tn[4].t24 XA.XIR[5].XIC[0].icell.PUM VPWR.t1528 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X482 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12].t25 XA.XIR[12].XIC[4].icell.Ien VGND.t304 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X483 XA.XIR[12].XIC[6].icell.PUM XA.Cn[6].t18 XA.XIR[12].XIC[6].icell.Ien VPWR.t424 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X484 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t1949 XA.XIR[7].XIC_dummy_right.icell.Ien VGND.t2208 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X485 VPWR.t875 VPWR.t873 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t874 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X486 XA.XIR[15].XIC[7].icell.PUM XA.Cn[7].t11 XA.XIR[15].XIC[7].icell.Ien VPWR.t1091 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X487 VGND.t1294 thermo15c_0.XTB4.Y.t4 XA.Cn[3].t3 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X488 VPWR.t1599 thermo15c_0.XTB2.Y XA.Cn[9].t6 VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X489 XA.XIR[5].XIC[12].icell.Ien XThR.Tn[5].t21 VPWR.t1499 VPWR.t1498 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X490 VGND.t2017 XA.Cn[3].t17 XA.XIR[7].XIC[3].icell.PDM VGND.t2016 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X491 VGND.t999 Vbias.t43 XA.XIR[6].XIC[11].icell.SM VGND.t998 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X492 VGND.t2210 VPWR.t1950 XA.XIR[2].XIC_15.icell.PDM VGND.t2209 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X493 VPWR.t1239 XThR.XTB5.Y XThR.Tn[12].t6 VPWR.t1238 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 VGND.t1176 XA.Cn[9].t17 XA.XIR[12].XIC[9].icell.PDM VGND.t1175 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X495 XA.XIR[14].XIC[3].icell.SM XA.XIR[14].XIC[3].icell.Ien Iout.t54 VGND.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X496 XA.XIR[9].XIC[12].icell.Ien XThR.Tn[9].t21 VPWR.t440 VPWR.t439 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X497 XA.XIR[8].XIC[13].icell.Ien XThR.Tn[8].t26 VPWR.t325 VPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X498 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout VGND.t2519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X499 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6].t20 XA.XIR[6].XIC[14].icell.Ien VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X500 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6].t21 XA.XIR[6].XIC[8].icell.Ien VGND.t353 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X501 VPWR.t1020 XThR.XTB7.Y XThR.Tn[14].t2 VPWR.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X502 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[1].t23 VGND.t705 VGND.t704 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X503 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13].t22 XA.XIR[13].XIC[12].icell.Ien VGND.t1920 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X504 XA.XIR[4].XIC[9].icell.PUM XA.Cn[9].t18 XA.XIR[4].XIC[9].icell.Ien VPWR.t1249 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X505 XThR.Tn[8].t7 XThR.XTB1.Y a_n997_3979# VGND.t1425 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X506 XA.XIR[3].XIC[10].icell.PUM XA.Cn[10].t16 XA.XIR[3].XIC[10].icell.Ien VPWR.t1379 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X507 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[4].t25 VGND.t215 VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X508 VGND.t853 XA.Cn[11].t17 XA.XIR[1].XIC[11].icell.PDM VGND.t852 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X509 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1951 VGND.t2212 VGND.t2211 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X510 VPWR.t277 XThR.Tn[7].t16 XA.XIR[8].XIC[6].icell.PUM VPWR.t276 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X511 VPWR.t1 data[2].t0 thermo15c_0.XTB7.B VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X512 VGND.t1733 VGND.t1731 XA.XIR[5].XIC_dummy_left.icell.SM VGND.t1732 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X513 VPWR.t1119 XThR.Tn[10].t20 XA.XIR[11].XIC[7].icell.PUM VPWR.t1118 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X514 VGND.t1434 XA.Cn[10].t17 XA.XIR[11].XIC[10].icell.PDM VGND.t1433 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X515 XA.Cn[13].t6 thermo15c_0.XTB6.Y a_10051_9569# VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X516 XThR.Tn[4].t11 XThR.XTBN.Y a_n1049_6405# VPWR.t1827 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X517 XThR.XTB5.Y XThR.XTB7.B a_n1319_6405# VPWR.t1218 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X518 VGND.t1001 Vbias.t44 XA.XIR[4].XIC[7].icell.SM VGND.t1000 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X519 XA.Cn[8].t11 thermo15c_0.XTBN.Y.t25 VPWR.t304 VPWR.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X520 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[13].t23 VGND.t1922 VGND.t1921 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X521 XA.XIR[15].XIC[11].icell.PUM XA.Cn[11].t18 XA.XIR[15].XIC[11].icell.Ien VPWR.t998 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X522 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[9].t22 VGND.t528 VGND.t527 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X523 a_n1335_4229# data[5].t0 XThR.XTB5.A VPWR.t1407 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X524 VGND.t838 XA.Cn[2].t17 XA.XIR[1].XIC[2].icell.PDM VGND.t837 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X525 VGND.t1003 Vbias.t45 XA.XIR[7].XIC[8].icell.SM VGND.t1002 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X526 XA.XIR[6].XIC[9].icell.Ien XThR.Tn[6].t22 VPWR.t229 VPWR.t228 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X527 XA.XIR[5].XIC[10].icell.Ien XThR.Tn[5].t22 VPWR.t1501 VPWR.t1500 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X528 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[12].t26 VGND.t306 VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X529 VGND.t1023 XA.Cn[7].t12 XA.XIR[7].XIC[7].icell.PDM VGND.t1022 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X530 VGND.t1005 Vbias.t46 XA.XIR[6].XIC[9].icell.SM VGND.t1004 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X531 VGND.t786 Vbias.t47 XA.XIR[3].XIC[11].icell.SM VGND.t785 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X532 XA.Cn[8].t6 thermo15c_0.XTB1.Y.t4 a_7651_9569# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X533 XA.Cn[13].t10 thermo15c_0.XTBN.Y.t26 VPWR.t305 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X534 VGND.t2019 XA.Cn[3].t18 XA.XIR[4].XIC[3].icell.PDM VGND.t2018 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X535 XA.XIR[9].XIC[10].icell.Ien XThR.Tn[9].t23 VPWR.t442 VPWR.t441 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X536 XA.XIR[7].XIC_15.icell.SM XA.XIR[7].XIC_15.icell.Ien Iout.t143 VGND.t1107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X537 XA.XIR[15].XIC[12].icell.SM XA.XIR[15].XIC[12].icell.Ien Iout.t144 VGND.t1108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X538 VPWR.t1475 VGND.t2690 XA.XIR[0].XIC[9].icell.PUM VPWR.t1474 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X539 VGND.t899 thermo15c_0.XTB6.Y XA.Cn[5].t2 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X540 XA.XIR[12].XIC[1].icell.PUM XA.Cn[1].t18 XA.XIR[12].XIC[1].icell.Ien VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X541 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t870 VPWR.t872 VPWR.t871 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X542 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[3].t23 VGND.t1515 VGND.t1514 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X543 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[3].t24 VGND.t1517 VGND.t1516 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X544 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13].t24 XA.XIR[13].XIC[10].icell.Ien VGND.t1923 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X545 XA.XIR[15].XIC[2].icell.PUM XA.Cn[2].t18 XA.XIR[15].XIC[2].icell.Ien VPWR.t119 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X546 XA.XIR[6].XIC[6].icell.PUM XA.Cn[6].t19 XA.XIR[6].XIC[6].icell.Ien VPWR.t425 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X547 XA.XIR[10].XIC[14].icell.PUM XA.Cn[14].t17 XA.XIR[10].XIC[14].icell.Ien VPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X548 VGND.t788 Vbias.t48 XA.XIR[12].XIC[5].icell.SM VGND.t787 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X549 VGND.t51 XA.Cn[4].t20 XA.XIR[12].XIC[4].icell.PDM VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X550 a_n1049_5611# XThR.XTB6.Y VPWR.t550 VPWR.t549 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X551 XA.XIR[13].XIC_15.icell.PUM VPWR.t868 XA.XIR[13].XIC_15.icell.Ien VPWR.t869 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X552 XThR.Tn[10].t7 XThR.XTB3.Y.t4 a_n997_2891# VGND.t1226 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X553 VGND.t790 Vbias.t49 XA.XIR[15].XIC[6].icell.SM VGND.t789 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X554 XA.XIR[0].XIC[11].icell.PDM XThR.Tn[0].t21 XA.XIR[0].XIC[11].icell.Ien VGND.t1961 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X555 VGND.t1603 XA.Cn[5].t15 XA.XIR[15].XIC[5].icell.PDM VGND.t1602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X556 VGND.t1178 XA.Cn[9].t19 XA.XIR[6].XIC[9].icell.PDM VGND.t1177 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X557 VPWR.t307 thermo15c_0.XTBN.Y.t27 XA.Cn[7].t2 VPWR.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X558 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6].t23 XA.XIR[6].XIC[3].icell.Ien VGND.t354 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X559 XA.XIR[1].XIC_15.icell.PDM XThR.Tn[1].t24 XA.XIR[1].XIC_15.icell.Ien VGND.t706 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X560 VPWR.t1121 XThR.Tn[10].t21 XA.XIR[11].XIC[11].icell.PUM VPWR.t1120 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X561 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t866 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t867 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X562 VPWR.t1668 XThR.XTB2.Y XThR.Tn[9].t6 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X563 VPWR.t1473 VGND.t2691 Vbias.t5 VPWR.t93 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X564 XA.Cn[6].t2 thermo15c_0.XTBN.Y.t28 a_6243_9615# VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X565 XA.XIR[3].XIC[5].icell.PUM XA.Cn[5].t16 XA.XIR[3].XIC[5].icell.Ien VPWR.t1438 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X566 VGND.t792 Vbias.t50 XA.XIR[9].XIC[5].icell.SM VGND.t791 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X567 XA.XIR[8].XIC[6].icell.Ien XThR.Tn[8].t27 VPWR.t327 VPWR.t326 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X568 VGND.t508 XA.Cn[6].t20 XA.XIR[1].XIC[6].icell.PDM VGND.t507 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X569 VPWR.t1045 XThR.Tn[3].t25 XA.XIR[4].XIC[4].icell.PUM VPWR.t1044 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X570 VPWR.t279 XThR.Tn[7].t17 XA.XIR[8].XIC[1].icell.PUM VPWR.t278 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X571 XA.XIR[0].XIC[2].icell.PDM XThR.Tn[0].t22 XA.XIR[0].XIC[2].icell.Ien VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X572 XA.XIR[11].XIC[7].icell.Ien XThR.Tn[11].t22 VPWR.t1840 VPWR.t1839 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X573 VGND.t794 Vbias.t51 XA.XIR[3].XIC[9].icell.SM VGND.t793 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X574 VGND.t1025 XA.Cn[7].t13 XA.XIR[4].XIC[7].icell.PDM VGND.t1024 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X575 XA.XIR[15].XIC_15.icell.Ien VPWR.t863 VPWR.t865 VPWR.t864 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X576 VPWR.t1123 XThR.Tn[10].t22 XA.XIR[11].XIC[2].icell.PUM VPWR.t1122 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X577 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout VGND.t1047 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X578 VPWR.t1503 XThR.Tn[5].t23 XA.XIR[6].XIC[14].icell.PUM VPWR.t1502 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X579 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t7 VPWR.t1774 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X580 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8].t28 XA.XIR[8].XIC[9].icell.Ien VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X581 XA.Cn[0].t9 thermo15c_0.XTBN.Y.t29 VGND.t396 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X582 VGND.t796 Vbias.t52 XA.XIR[4].XIC[2].icell.SM VGND.t795 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X583 VPWR.t862 VPWR.t860 XA.XIR[9].XIC_15.icell.PUM VPWR.t861 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X584 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[0].t23 VGND.t42 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X585 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[0].t24 VGND.t44 VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X586 VGND.t798 Vbias.t53 XA.XIR[7].XIC[3].icell.SM VGND.t797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X587 a_4067_9615# thermo15c_0.XTBN.Y.t30 XA.Cn[2].t9 VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X588 XThR.Tn[0].t3 XThR.XTB1.Y VGND.t1424 VGND.t1423 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X589 VGND.t2444 XThR.XTBN.Y XThR.Tn[5].t10 VGND.t2430 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X590 XA.XIR[11].XIC[7].icell.SM XA.XIR[11].XIC[7].icell.Ien Iout.t181 VGND.t1388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X591 XA.XIR[5].XIC[5].icell.Ien XThR.Tn[5].t24 VPWR.t1505 VPWR.t1504 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X592 VGND.t800 Vbias.t54 XA.XIR[6].XIC[4].icell.SM VGND.t799 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X593 XThR.Tn[14].t7 XThR.XTB7.Y a_n997_715# VGND.t891 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X594 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[12].t27 VGND.t308 VGND.t307 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X595 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[7].t18 VGND.t380 VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X596 VGND.t802 Vbias.t55 XA.XIR[15].XIC[10].icell.SM VGND.t801 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X597 XA.XIR[9].XIC[5].icell.Ien XThR.Tn[9].t24 VPWR.t444 VPWR.t443 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X598 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[10].t23 VGND.t1093 VGND.t1092 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X599 XA.XIR[10].XIC[11].icell.SM XA.XIR[10].XIC[11].icell.Ien Iout.t232 VGND.t2003 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X600 VGND.t2214 VPWR.t1952 XA.XIR[11].XIC_dummy_left.icell.PDM VGND.t2213 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X601 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6].t24 XA.XIR[6].XIC[7].icell.Ien VGND.t355 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X602 VGND.t2443 XThR.XTBN.Y XThR.Tn[4].t7 VGND.t2442 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X603 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[3].t26 VGND.t909 VGND.t908 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X604 XA.XIR[6].XIC[1].icell.PUM XA.Cn[1].t19 XA.XIR[6].XIC[1].icell.Ien VPWR.t1878 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X605 VGND.t2216 VPWR.t1953 XA.XIR[14].XIC_15.icell.PDM VGND.t2215 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X606 a_8963_9569# thermo15c_0.XTB4.Y.t5 XA.Cn[11].t6 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X607 XA.XIR[5].XIC[13].icell.PUM XA.Cn[13].t18 XA.XIR[5].XIC[13].icell.Ien VPWR.t1330 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X608 VGND.t804 Vbias.t56 XA.XIR[12].XIC[0].icell.SM VGND.t803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X609 XA.XIR[1].XIC[14].icell.SM XA.XIR[1].XIC[14].icell.Ien Iout.t196 VGND.t1498 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X610 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t858 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t859 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X611 XA.XIR[9].XIC[13].icell.PUM XA.Cn[13].t19 XA.XIR[9].XIC[13].icell.Ien VPWR.t1331 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X612 VGND.t806 Vbias.t57 XA.XIR[15].XIC[1].icell.SM VGND.t805 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X613 XA.XIR[0].XIC[6].icell.PDM XThR.Tn[0].t25 XA.XIR[0].XIC[6].icell.Ien VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X614 VGND.t53 XA.Cn[4].t21 XA.XIR[6].XIC[4].icell.PDM VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X615 VGND.t1927 XA.Cn[0].t18 XA.XIR[15].XIC[0].icell.PDM VGND.t1926 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X616 VGND.t808 Vbias.t58 XA.XIR[10].XIC[13].icell.SM VGND.t807 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X617 XA.XIR[11].XIC[11].icell.Ien XThR.Tn[11].t23 VPWR.t1842 VPWR.t1841 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X618 VGND.t2644 XA.Cn[12].t17 XA.XIR[10].XIC[12].icell.PDM VGND.t2643 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X619 VPWR.t1047 XThR.Tn[3].t27 XA.XIR[4].XIC[0].icell.PUM VPWR.t1046 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X620 VGND.t1296 Vbias.t59 XA.XIR[13].XIC[14].icell.SM VGND.t1295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X621 XA.XIR[12].XIC_15.icell.Ien XThR.Tn[12].t28 VPWR.t179 VPWR.t178 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X622 VGND.t496 thermo15c_0.XTBN.Y.t31 a_8739_9569# VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X623 VGND.t1348 XA.Cn[13].t20 XA.XIR[13].XIC[13].icell.PDM VGND.t1347 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X624 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t1954 XA.XIR[13].XIC_dummy_left.icell.Ien VGND.t2217 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X625 VPWR.t94 bias[0].t0 Vbias.t0 VPWR.t93 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X626 VGND.t1298 Vbias.t60 XA.XIR[9].XIC[0].icell.SM VGND.t1297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X627 XA.XIR[4].XIC[4].icell.Ien XThR.Tn[4].t26 VPWR.t108 VPWR.t107 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X628 XA.XIR[8].XIC[1].icell.Ien XThR.Tn[8].t29 VPWR.t1112 VPWR.t1111 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X629 VGND.t1300 Vbias.t61 XA.XIR[0].XIC_15.icell.SM VGND.t1299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X630 VGND.t1052 XA.Cn[8].t18 XA.XIR[0].XIC[8].icell.PDM VGND.t1051 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X631 VGND.t170 XA.Cn[14].t18 XA.XIR[0].XIC[14].icell.PDM VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X632 XA.XIR[11].XIC[2].icell.Ien XThR.Tn[11].t24 VPWR.t1844 VPWR.t1843 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X633 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[7].t19 VGND.t382 VGND.t381 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X634 XA.XIR[8].XIC[7].icell.SM XA.XIR[8].XIC[7].icell.Ien Iout.t104 VGND.t818 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X635 a_9827_9569# thermo15c_0.XTBN.Y.t32 VGND.t497 VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X636 VGND.t1302 Vbias.t62 XA.XIR[3].XIC[4].icell.SM VGND.t1301 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X637 XA.XIR[7].XIC[8].icell.SM XA.XIR[7].XIC[8].icell.Ien Iout.t123 VGND.t1028 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X638 VPWR.t515 XThR.Tn[1].t25 XA.XIR[2].XIC[12].icell.PUM VPWR.t514 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X639 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8].t30 XA.XIR[8].XIC[4].icell.Ien VGND.t1065 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X640 VPWR.t17 XThR.Tn[0].t26 XA.XIR[1].XIC[13].icell.PUM VPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X641 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t1955 XA.XIR[3].XIC_dummy_right.icell.Ien VGND.t2218 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X642 XA.XIR[10].XIC[9].icell.SM XA.XIR[10].XIC[9].icell.Ien Iout.t189 VGND.t1428 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X643 VPWR.t110 XThR.Tn[4].t27 XA.XIR[5].XIC[13].icell.PUM VPWR.t109 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X644 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11].t25 XA.XIR[11].XIC[5].icell.Ien VGND.t2479 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X645 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[3].t28 VGND.t911 VGND.t910 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X646 VPWR.t857 VPWR.t855 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t856 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X647 XA.XIR[15].XIC[13].icell.PDM VPWR.t1956 XA.XIR[15].XIC[13].icell.Ien VGND.t2219 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X648 VGND.t369 thermo15c_0.XTB1.Y.t5 XA.Cn[0].t2 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[0].t27 VGND.t47 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X650 XA.XIR[11].XIC[2].icell.SM XA.XIR[11].XIC[2].icell.Ien Iout.t146 VGND.t1118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X651 XThR.XTB7.A data[5].t1 VPWR.t1908 VPWR.t1907 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X652 VGND.t1436 XA.Cn[10].t18 XA.XIR[10].XIC[10].icell.PDM VGND.t1435 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X653 VPWR.t181 XThR.Tn[12].t29 XA.XIR[13].XIC[8].icell.PUM VPWR.t180 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X654 VGND.t822 thermo15c_0.XTBN.A thermo15c_0.XTBN.Y.t3 VGND.t821 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X655 XA.XIR[0].XIC[9].icell.PUM XA.Cn[9].t20 XA.XIR[0].XIC[9].icell.Ien VPWR.t1250 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X656 VPWR.t1217 XThR.XTB7.B XThR.XTB1.Y VPWR.t1216 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X657 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t6 VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X658 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[2].t22 VGND.t2601 VGND.t2600 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X659 XA.XIR[4].XIC[0].icell.Ien XThR.Tn[4].t28 VPWR.t112 VPWR.t111 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X660 XA.XIR[14].XIC[12].icell.SM XA.XIR[14].XIC[12].icell.Ien Iout.t186 VGND.t1413 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X661 XA.XIR[14].XIC_15.icell.PDM VPWR.t1957 VGND.t2221 VGND.t2220 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X662 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t852 VPWR.t854 VPWR.t853 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X663 XA.XIR[13].XIC[5].icell.SM XA.XIR[13].XIC[5].icell.Ien Iout.t163 VGND.t1281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X664 VPWR.t517 XThR.Tn[1].t26 XA.XIR[2].XIC[10].icell.PUM VPWR.t516 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X665 XA.XIR[5].XIC[6].icell.PUM XA.Cn[6].t21 XA.XIR[5].XIC[6].icell.Ien VPWR.t426 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X666 XA.Cn[7].t1 thermo15c_0.XTBN.Y.t33 VPWR.t419 VPWR.t418 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X667 VGND.t1138 XThR.XTB7.B a_n1335_7243# VGND.t1137 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X668 XA.XIR[9].XIC[6].icell.PUM XA.Cn[6].t22 XA.XIR[9].XIC[6].icell.Ien VPWR.t427 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X669 XA.XIR[8].XIC[7].icell.PUM XA.Cn[7].t14 XA.XIR[8].XIC[7].icell.Ien VPWR.t1086 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X670 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[0].t28 VGND.t49 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X671 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1958 VGND.t2223 VGND.t2222 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X672 XA.XIR[12].XIC_15.icell.PUM VPWR.t850 XA.XIR[12].XIC_15.icell.Ien VPWR.t851 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X673 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[8].t31 VGND.t1067 VGND.t1066 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X674 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12].t30 XA.XIR[12].XIC[13].icell.Ien VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X675 VGND.t2523 XA.Cn[3].t19 XA.XIR[0].XIC[3].icell.PDM VGND.t2522 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X676 XA.XIR[11].XIC[8].icell.PUM XA.Cn[8].t19 XA.XIR[11].XIC[8].icell.Ien VPWR.t1098 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X677 VGND.t1180 XA.Cn[9].t21 XA.XIR[5].XIC[9].icell.PDM VGND.t1179 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X678 XA.XIR[8].XIC[2].icell.SM XA.XIR[8].XIC[2].icell.Ien Iout.t100 VGND.t773 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X679 XA.XIR[2].XIC[12].icell.Ien XThR.Tn[2].t23 VPWR.t1184 VPWR.t1183 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X680 XA.XIR[7].XIC[3].icell.SM XA.XIR[7].XIC[3].icell.Ien Iout.t101 VGND.t774 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X681 XA.Cn[11].t7 thermo15c_0.XTB4.Y.t6 VPWR.t1888 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X682 VGND.t1182 XA.Cn[9].t22 XA.XIR[9].XIC[9].icell.PDM VGND.t1181 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X683 XA.XIR[10].XIC[4].icell.SM XA.XIR[10].XIC[4].icell.Ien Iout.t250 VGND.t2618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X684 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t847 VPWR.t849 VPWR.t848 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X685 a_n997_1803# XThR.XTBN.Y VGND.t2441 VGND.t2440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X686 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11].t26 XA.XIR[11].XIC[0].icell.Ien VGND.t2480 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X687 XThR.Tn[3].t6 XThR.XTBN.Y a_n1049_6699# VPWR.t1826 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X688 VPWR.t446 XThR.Tn[9].t25 XA.XIR[10].XIC[8].icell.PUM VPWR.t445 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X689 VGND.t2439 XThR.XTBN.Y XThR.Tn[3].t10 VGND.t2405 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X690 VGND.t1304 Vbias.t63 XA.XIR[11].XIC[6].icell.SM VGND.t1303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X691 XA.XIR[10].XIC[7].icell.Ien XThR.Tn[10].t24 VPWR.t1125 VPWR.t1124 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X692 VGND.t2225 VPWR.t1959 XA.XIR[7].XIC_dummy_right.icell.PDM VGND.t2224 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X693 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1960 VGND.t2227 VGND.t2226 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X694 XA.Cn[2].t8 thermo15c_0.XTBN.Y.t34 a_4067_9615# VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X695 VPWR.t984 XThR.Tn[0].t29 XA.XIR[1].XIC[6].icell.PUM VPWR.t983 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X696 XA.XIR[13].XIC[8].icell.Ien XThR.Tn[13].t25 VPWR.t1584 VPWR.t1583 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X697 VPWR.t114 XThR.Tn[4].t29 XA.XIR[5].XIC[6].icell.PUM VPWR.t113 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X698 VPWR.t183 XThR.Tn[12].t31 XA.XIR[13].XIC[3].icell.PUM VPWR.t182 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X699 XThR.Tn[11].t7 XThR.XTB4.Y.t5 VPWR.t1490 VPWR.t1230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X700 VPWR.t846 VPWR.t844 XA.XIR[8].XIC_15.icell.PUM VPWR.t845 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X701 VPWR.t1598 thermo15c_0.XTB2.Y a_3773_9615# VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X702 a_n1049_8581# XThR.XTB1.Y VPWR.t1374 VPWR.t1373 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X703 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t842 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t843 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X704 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[2].t24 VGND.t2599 VGND.t2598 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X705 XA.XIR[8].XIC[11].icell.PUM XA.Cn[11].t19 XA.XIR[8].XIC[11].icell.Ien VPWR.t999 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X706 VGND.t1306 Vbias.t64 XA.XIR[0].XIC[8].icell.SM VGND.t1305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X707 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[10].t25 VGND.t1095 VGND.t1094 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X708 VGND.t1013 XA.Cn[7].t15 XA.XIR[0].XIC[7].icell.PDM VGND.t1012 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X709 VGND.t1730 VGND.t1728 XA.XIR[4].XIC_dummy_right.icell.SM VGND.t1729 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X710 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[5].t25 VGND.t1772 VGND.t1771 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X711 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[9].t26 VGND.t530 VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X712 XA.XIR[9].XIC[11].icell.SM XA.XIR[9].XIC[11].icell.Ien Iout.t126 VGND.t1033 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X713 XA.XIR[2].XIC[10].icell.Ien XThR.Tn[2].t25 VPWR.t1176 VPWR.t1175 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X714 XA.XIR[13].XIC[0].icell.SM XA.XIR[13].XIC[0].icell.Ien Iout.t80 VGND.t666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X715 VGND.t2229 VPWR.t1961 XA.XIR[10].XIC_dummy_left.icell.PDM VGND.t2228 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X716 VPWR.t1209 thermo15c_0.XTB6.A a_5949_10571# VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X717 VPWR.t1648 XThR.Tn[1].t27 XA.XIR[2].XIC[5].icell.PUM VPWR.t1647 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X718 XA.XIR[1].XIC[4].icell.PUM XA.Cn[4].t22 XA.XIR[1].XIC[4].icell.Ien VPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X719 XA.XIR[5].XIC[1].icell.PUM XA.Cn[1].t20 XA.XIR[5].XIC[1].icell.Ien VPWR.t1879 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X720 VGND.t302 XThR.XTB3.Y.t5 XThR.Tn[2].t1 VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X721 VPWR.t1586 XThR.Tn[13].t26 XA.XIR[14].XIC[9].icell.PUM VPWR.t1585 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X722 XA.XIR[9].XIC[1].icell.PUM XA.Cn[1].t21 XA.XIR[9].XIC[1].icell.Ien VPWR.t1880 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X723 XA.XIR[8].XIC[2].icell.PUM XA.Cn[2].t19 XA.XIR[8].XIC[2].icell.Ien VPWR.t120 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X724 XA.XIR[3].XIC[14].icell.PUM XA.Cn[14].t19 XA.XIR[3].XIC[14].icell.Ien VPWR.t83 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X725 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[8].t32 VGND.t1069 VGND.t1068 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X726 XA.XIR[0].XIC[6].icell.SM XA.XIR[0].XIC[6].icell.Ien Iout.t34 VGND.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X727 thermo15c_0.XTBN.Y.t1 thermo15c_0.XTBN.A VPWR.t979 VPWR.t978 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X728 VGND.t1308 Vbias.t65 XA.XIR[5].XIC[5].icell.SM VGND.t1307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X729 XA.XIR[11].XIC[3].icell.PUM XA.Cn[3].t20 XA.XIR[11].XIC[3].icell.Ien VPWR.t1852 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X730 VGND.t55 XA.Cn[4].t23 XA.XIR[5].XIC[4].icell.PDM VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X731 VGND.t1310 Vbias.t66 XA.XIR[11].XIC[10].icell.SM VGND.t1309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X732 XA.XIR[10].XIC[11].icell.Ien XThR.Tn[10].t26 VPWR.t1509 VPWR.t1508 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X733 XThR.Tn[8].t6 XThR.XTB1.Y a_n997_3979# VGND.t1422 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X734 XA.XIR[6].XIC_15.icell.PUM VPWR.t840 XA.XIR[6].XIC_15.icell.Ien VPWR.t841 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X735 VGND.t2553 XA.Cn[1].t22 XA.XIR[13].XIC[1].icell.PDM VGND.t2552 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X736 VGND.t1312 Vbias.t67 XA.XIR[12].XIC[14].icell.SM VGND.t1311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X737 VGND.t57 XA.Cn[4].t24 XA.XIR[9].XIC[4].icell.PDM VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X738 VGND.t1314 Vbias.t68 XA.XIR[8].XIC[6].icell.SM VGND.t1313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X739 XA.XIR[7].XIC[7].icell.Ien XThR.Tn[7].t20 VPWR.t532 VPWR.t531 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X740 VGND.t2231 VPWR.t1962 XA.XIR[4].XIC_dummy_right.icell.PDM VGND.t2230 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X741 VGND.t1605 XA.Cn[5].t17 XA.XIR[8].XIC[5].icell.PDM VGND.t1604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X742 VGND.t81 XA.Cn[13].t21 XA.XIR[12].XIC[13].icell.PDM VGND.t80 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X743 VGND.t498 thermo15c_0.XTBN.Y.t35 a_9827_9569# VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X744 XA.XIR[2].XIC[12].icell.PUM XA.Cn[12].t18 XA.XIR[2].XIC[12].icell.Ien VPWR.t1919 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X745 VPWR.t448 XThR.Tn[9].t27 XA.XIR[10].XIC[3].icell.PUM VPWR.t447 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X746 VPWR.t1353 thermo15c_0.XTB7.Y XA.Cn[14].t7 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X747 XThR.Tn[4].t10 XThR.XTBN.Y a_n1049_6405# VPWR.t1826 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X748 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14].t23 XA.XIR[14].XIC[8].icell.Ien VGND.t319 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X749 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14].t24 XA.XIR[14].XIC[14].icell.Ien VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X750 VGND.t1316 Vbias.t69 XA.XIR[11].XIC[1].icell.SM VGND.t1315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X751 XA.XIR[10].XIC[2].icell.Ien XThR.Tn[10].t27 VPWR.t1511 VPWR.t1510 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X752 VGND.t1318 Vbias.t70 XA.XIR[7].XIC[12].icell.SM VGND.t1317 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X753 VPWR.t1491 XThR.XTB4.Y.t6 a_n1049_6699# VPWR.t1236 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X754 XA.XIR[5].XIC[14].icell.Ien XThR.Tn[5].t26 VPWR.t1286 VPWR.t1285 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X755 VGND.t2662 Vbias.t71 XA.XIR[6].XIC[13].icell.SM VGND.t2661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X756 VPWR.t986 XThR.Tn[0].t30 XA.XIR[1].XIC[1].icell.PUM VPWR.t985 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X757 XA.XIR[13].XIC[3].icell.Ien XThR.Tn[13].t27 VPWR.t1083 VPWR.t1082 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X758 XA.XIR[9].XIC[14].icell.Ien XThR.Tn[9].t28 VPWR.t450 VPWR.t449 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X759 VGND.t2664 Vbias.t72 XA.XIR[9].XIC[14].icell.SM VGND.t2663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X760 VPWR.t116 XThR.Tn[4].t30 XA.XIR[5].XIC[1].icell.PUM VPWR.t115 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X761 XA.XIR[9].XIC[9].icell.SM XA.XIR[9].XIC[9].icell.Ien Iout.t233 VGND.t2125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X762 XA.XIR[8].XIC_15.icell.Ien XThR.Tn[8].t33 VPWR.t1114 VPWR.t1113 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X763 XA.XIR[15].XIC[1].icell.PDM VPWR.t1963 XA.XIR[15].XIC[1].icell.Ien VGND.t2232 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X764 VPWR.t1049 XThR.Tn[3].t29 XA.XIR[4].XIC[13].icell.PUM VPWR.t1048 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X765 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10].t28 XA.XIR[10].XIC[5].icell.Ien VGND.t1774 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X766 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1964 XA.XIR[6].XIC_dummy_right.icell.Ien VGND.t2233 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X767 XA.XIR[0].XIC[4].icell.Ien XThR.Tn[0].t31 VPWR.t988 VPWR.t987 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X768 XA.XIR[1].XIC[0].icell.PUM XA.Cn[0].t19 XA.XIR[1].XIC[0].icell.Ien VPWR.t1590 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X769 VGND.t2666 Vbias.t73 XA.XIR[0].XIC[3].icell.SM VGND.t2665 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X770 XA.XIR[4].XIC[7].icell.SM XA.XIR[4].XIC[7].icell.Ien Iout.t134 VGND.t1059 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X771 XA.XIR[0].XIC[10].icell.SM XA.XIR[0].XIC[10].icell.Ien Iout.t43 VGND.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X772 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[5].t27 VGND.t1262 VGND.t1261 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X773 XA.XIR[2].XIC[5].icell.Ien XThR.Tn[2].t26 VPWR.t1182 VPWR.t1181 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X774 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout VGND.t2167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X775 VGND.t2668 Vbias.t74 XA.XIR[8].XIC[10].icell.SM VGND.t2667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X776 VPWR.t1825 XThR.XTBN.Y XThR.Tn[8].t11 VPWR.t1824 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X777 XA.XIR[7].XIC[11].icell.Ien XThR.Tn[7].t21 VPWR.t534 VPWR.t533 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X778 XThR.Tn[10].t6 XThR.XTB3.Y.t6 a_n997_2891# VGND.t1228 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X779 XA.XIR[14].XIC[9].icell.Ien XThR.Tn[14].t25 VPWR.t191 VPWR.t190 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X780 XA.XIR[2].XIC[10].icell.PUM XA.Cn[10].t19 XA.XIR[2].XIC[10].icell.Ien VPWR.t1380 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X781 thermo15c_0.XTB3.Y.t0 thermo15c_0.XTB7.B VPWR.t1129 VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X782 XA.XIR[0].XIC[1].icell.SM XA.XIR[0].XIC[1].icell.Ien Iout.t205 VGND.t1518 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X783 VGND.t2670 Vbias.t75 XA.XIR[5].XIC[0].icell.SM VGND.t2669 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X784 VGND.t1727 VGND.t1725 XA.XIR[4].XIC_dummy_left.icell.SM VGND.t1726 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X785 VGND.t2672 Vbias.t76 XA.XIR[8].XIC[1].icell.SM VGND.t2671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X786 VPWR.t1208 thermo15c_0.XTB6.A thermo15c_0.XTB2.Y VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X787 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[11].t27 VGND.t2482 VGND.t2481 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X788 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[11].t28 VGND.t105 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X789 XA.XIR[12].XIC[5].icell.SM XA.XIR[12].XIC[5].icell.Ien Iout.t25 VGND.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X790 XA.XIR[7].XIC[2].icell.Ien XThR.Tn[7].t22 VPWR.t536 VPWR.t535 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X791 VGND.t2674 Vbias.t77 XA.XIR[3].XIC[13].icell.SM VGND.t2673 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X792 VGND.t1929 XA.Cn[0].t20 XA.XIR[8].XIC[0].icell.PDM VGND.t1928 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X793 VGND.t2646 XA.Cn[12].t19 XA.XIR[3].XIC[12].icell.PDM VGND.t2645 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X794 XThR.XTB3.Y.t2 XThR.XTB7.A VPWR.t1389 VPWR.t1388 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X795 XA.XIR[15].XIC[6].icell.SM XA.XIR[15].XIC[6].icell.Ien Iout.t11 VGND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X796 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12].t32 XA.XIR[12].XIC[1].icell.Ien VGND.t310 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X797 VGND.t83 XA.Cn[13].t22 XA.XIR[6].XIC[13].icell.PDM VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X798 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7].t23 XA.XIR[7].XIC[5].icell.Ien VGND.t731 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X799 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1965 VGND.t2235 VGND.t2234 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X800 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t6 VGND.t890 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X801 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14].t26 XA.XIR[14].XIC[3].icell.Ien VGND.t321 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X802 XA.XIR[10].XIC[8].icell.PUM XA.Cn[8].t20 XA.XIR[10].XIC[8].icell.Ien VPWR.t1099 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X803 XA.XIR[1].XIC[12].icell.Ien XThR.Tn[1].t28 VPWR.t1650 VPWR.t1649 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X804 VGND.t2676 Vbias.t78 XA.XIR[2].XIC[11].icell.SM VGND.t2675 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X805 XA.XIR[6].XIC_15.icell.SM XA.XIR[6].XIC_15.icell.Ien Iout.t75 VGND.t565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X806 XA.XIR[0].XIC[0].icell.Ien XThR.Tn[0].t32 VPWR.t990 VPWR.t989 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X807 XThR.Tn[0].t11 XThR.XTBN.Y VGND.t2438 VGND.t2381 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X808 VPWR.t1237 XThR.XTB5.Y a_n1049_6405# VPWR.t1236 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X809 XA.XIR[4].XIC[13].icell.Ien XThR.Tn[4].t31 VPWR.t118 VPWR.t117 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X810 VGND.t2678 Vbias.t79 XA.XIR[14].XIC_15.icell.SM VGND.t2677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X811 XA.XIR[9].XIC[4].icell.SM XA.XIR[9].XIC[4].icell.Ien Iout.t13 VGND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X812 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10].t29 XA.XIR[10].XIC[0].icell.Ien VGND.t1775 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X813 XA.Cn[10].t1 thermo15c_0.XTB3.Y.t4 VPWR.t1014 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X814 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5].t28 XA.XIR[5].XIC[12].icell.Ien VGND.t1263 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X815 VPWR.t1823 XThR.XTBN.Y XThR.Tn[10].t11 VPWR.t1822 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X816 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout VGND.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X817 VPWR.t36 XThR.Tn[11].t29 XA.XIR[12].XIC[4].icell.PUM VPWR.t35 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X818 VPWR.t420 thermo15c_0.XTBN.Y.t36 XA.Cn[13].t9 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X819 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9].t29 XA.XIR[9].XIC[12].icell.Ien VGND.t531 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X820 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8].t34 XA.XIR[8].XIC[13].icell.Ien VGND.t1070 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X821 a_3773_9615# thermo15c_0.XTB2.Y VPWR.t1597 VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X822 XA.Cn[5].t1 thermo15c_0.XTB6.Y VGND.t898 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X823 XA.XIR[4].XIC[2].icell.SM XA.XIR[4].XIC[2].icell.Ien Iout.t162 VGND.t1170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X824 XA.Cn[2].t0 thermo15c_0.XTB3.Y.t5 VGND.t873 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X825 VPWR.t1051 XThR.Tn[3].t30 XA.XIR[4].XIC[6].icell.PUM VPWR.t1050 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X826 VPWR.t1180 XThR.Tn[2].t27 XA.XIR[3].XIC[7].icell.PUM VPWR.t1179 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X827 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[12].t33 VGND.t312 VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X828 VGND.t1438 XA.Cn[10].t20 XA.XIR[3].XIC[10].icell.PDM VGND.t1437 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X829 VPWR.t231 XThR.Tn[6].t25 XA.XIR[7].XIC[7].icell.PUM VPWR.t230 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X830 XA.XIR[15].XIC[10].icell.SM XA.XIR[15].XIC[10].icell.Ien Iout.t125 VGND.t1032 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X831 VPWR.t1288 XThR.Tn[5].t29 XA.XIR[6].XIC[8].icell.PUM VPWR.t1287 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X832 VGND.t2437 XThR.XTBN.Y a_n997_3755# VGND.t2426 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X833 XA.XIR[2].XIC[5].icell.PUM XA.Cn[5].t18 XA.XIR[2].XIC[5].icell.Ien VPWR.t1439 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X834 VPWR.t259 thermo15c_0.XTB1.Y.t6 a_2979_9615# VPWR.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X835 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[9].t30 VGND.t533 VGND.t532 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X836 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1966 VGND.t2237 VGND.t2236 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X837 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14].t27 XA.XIR[14].XIC[7].icell.Ien VGND.t322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X838 XA.XIR[1].XIC[10].icell.Ien XThR.Tn[1].t29 VPWR.t1652 VPWR.t1651 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X839 VGND.t2680 Vbias.t80 XA.XIR[2].XIC[9].icell.SM VGND.t2679 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X840 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[12].t34 VGND.t314 VGND.t313 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X841 XA.XIR[12].XIC[0].icell.SM XA.XIR[12].XIC[0].icell.Ien Iout.t68 VGND.t548 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X842 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[11].t30 VGND.t107 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X843 XA.XIR[3].XIC_15.icell.SM XA.XIR[3].XIC_15.icell.Ien Iout.t6 VGND.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X844 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout VGND.t1521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X845 XA.XIR[7].XIC[12].icell.SM XA.XIR[7].XIC[12].icell.Ien Iout.t18 VGND.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X846 XA.XIR[14].XIC[12].icell.PUM XA.Cn[12].t20 XA.XIR[14].XIC[12].icell.Ien VPWR.t1920 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X847 XA.XIR[15].XIC[1].icell.SM XA.XIR[15].XIC[1].icell.Ien Iout.t17 VGND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X848 VGND.t855 XA.Cn[11].t20 XA.XIR[15].XIC[11].icell.PDM VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X849 XA.XIR[11].XIC_15.icell.PDM VPWR.t1967 VGND.t2239 VGND.t2238 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X850 XA.XIR[10].XIC[13].icell.SM XA.XIR[10].XIC[13].icell.Ien Iout.t156 VGND.t1157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X851 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5].t30 XA.XIR[5].XIC[10].icell.Ien VGND.t1264 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X852 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7].t24 XA.XIR[7].XIC[0].icell.Ien VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X853 XA.XIR[13].XIC[14].icell.SM XA.XIR[13].XIC[14].icell.Ien Iout.t102 VGND.t809 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X854 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9].t31 XA.XIR[9].XIC[10].icell.Ien VGND.t534 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X855 XA.XIR[10].XIC[3].icell.PUM XA.Cn[3].t21 XA.XIR[10].XIC[3].icell.Ien VPWR.t1853 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X856 a_5155_9615# thermo15c_0.XTB5.Y VPWR.t341 VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X857 XA.XIR[5].XIC_15.icell.PUM VPWR.t838 XA.XIR[5].XIC_15.icell.Ien VPWR.t839 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X858 VPWR.t38 XThR.Tn[11].t31 XA.XIR[12].XIC[0].icell.PUM VPWR.t37 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X859 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[6].t26 VGND.t357 VGND.t356 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X860 a_n1049_7493# XThR.XTB3.Y.t7 VPWR.t1093 VPWR.t1092 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X861 VGND.t2555 XA.Cn[1].t23 XA.XIR[12].XIC[1].icell.PDM VGND.t2554 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X862 XA.XIR[9].XIC_15.icell.PUM VPWR.t836 XA.XIR[9].XIC_15.icell.Ien VPWR.t837 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X863 VGND.t217 XA.Cn[2].t20 XA.XIR[15].XIC[2].icell.PDM VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X864 VPWR.t1178 XThR.Tn[2].t28 XA.XIR[3].XIC[11].icell.PUM VPWR.t1177 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X865 VPWR.t233 XThR.Tn[6].t27 XA.XIR[7].XIC[11].icell.PUM VPWR.t232 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X866 VGND.t2241 VPWR.t1968 XA.XIR[13].XIC_15.icell.PDM VGND.t2240 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X867 XA.Cn[8].t3 thermo15c_0.XTB1.Y.t7 VPWR.t261 VPWR.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X868 Vbias.t1 bias[2].t0 VPWR.t267 VPWR.t266 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X869 XA.XIR[4].XIC[6].icell.Ien XThR.Tn[4].t32 VPWR.t1602 VPWR.t1601 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X870 XA.XIR[3].XIC[7].icell.Ien XThR.Tn[3].t31 VPWR.t1053 VPWR.t1052 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X871 VGND.t1168 XThR.XTB5.Y XThR.Tn[4].t3 VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X872 a_5155_9615# thermo15c_0.XTBN.Y.t37 XA.Cn[4].t7 VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X873 VGND.t2243 VPWR.t1969 XA.XIR[0].XIC_dummy_right.icell.PDM VGND.t2242 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X874 VPWR.t1055 XThR.Tn[3].t32 XA.XIR[4].XIC[1].icell.PUM VPWR.t1054 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X875 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[12].t35 VGND.t316 VGND.t315 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X876 VPWR.t1174 XThR.Tn[2].t29 XA.XIR[3].XIC[2].icell.PUM VPWR.t1173 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X877 XThR.XTB5.Y XThR.XTB5.A VGND.t20 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X878 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[11].t32 VGND.t109 VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X879 VPWR.t235 XThR.Tn[6].t28 XA.XIR[7].XIC[2].icell.PUM VPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X880 VPWR.t1654 XThR.Tn[1].t30 XA.XIR[2].XIC[14].icell.PUM VPWR.t1653 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X881 VPWR.t1290 XThR.Tn[5].t31 XA.XIR[6].XIC[3].icell.PUM VPWR.t1289 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X882 XA.XIR[14].XIC[10].icell.PUM XA.Cn[10].t21 XA.XIR[14].XIC[10].icell.Ien VPWR.t1381 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X883 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout VGND.t1045 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X884 VPWR.t835 VPWR.t833 XA.XIR[1].XIC_15.icell.PUM VPWR.t834 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X885 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[4].t33 XA.XIR[4].XIC[9].icell.Ien VGND.t1945 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X886 VPWR.t832 VPWR.t830 XA.XIR[5].XIC_15.icell.PUM VPWR.t831 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X887 XA.XIR[15].XIC_15.icell.PDM VPWR.t1970 XA.XIR[15].XIC_15.icell.Ien VGND.t2244 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X888 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[6].t29 VGND.t359 VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X889 XA.XIR[1].XIC[5].icell.Ien XThR.Tn[1].t31 VPWR.t1656 VPWR.t1655 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X890 VGND.t2682 Vbias.t81 XA.XIR[2].XIC[4].icell.SM VGND.t2681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X891 XA.XIR[6].XIC[8].icell.SM XA.XIR[6].XIC[8].icell.Ien Iout.t191 VGND.t1452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X892 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[2].t30 VGND.t1572 VGND.t1571 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X893 VGND.t2684 Vbias.t82 XA.XIR[15].XIC[7].icell.SM VGND.t2683 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X894 VGND.t2246 VPWR.t1971 XA.XIR[3].XIC_dummy_left.icell.PDM VGND.t2245 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X895 VGND.t263 Vbias.t83 XA.XIR[14].XIC[8].icell.SM VGND.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X896 VGND.t510 XA.Cn[6].t23 XA.XIR[15].XIC[6].icell.PDM VGND.t509 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X897 VPWR.t829 VPWR.t827 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t828 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X898 XA.Cn[14].t10 thermo15c_0.XTB7.Y a_10915_9569# VGND.t1399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X899 thermo15c_0.XTB3.Y.t1 thermo15c_0.XTB7.A a_4387_10575# VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X900 a_n997_1803# XThR.XTBN.Y VGND.t2436 VGND.t2435 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X901 XA.XIR[1].XIC[13].icell.PUM XA.Cn[13].t23 XA.XIR[1].XIC[13].icell.Ien VPWR.t25 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X902 XA.XIR[3].XIC[11].icell.Ien XThR.Tn[3].t33 VPWR.t1057 VPWR.t1056 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X903 XA.XIR[15].XIC[14].icell.PDM XThR.Tn[14].t28 VGND.t324 VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X904 a_3773_9615# thermo15c_0.XTBN.Y.t38 XA.Cn[1].t3 VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X905 VGND.t2557 XA.Cn[1].t24 XA.XIR[6].XIC[1].icell.PDM VGND.t2556 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X906 XA.XIR[14].XIC[6].icell.SM XA.XIR[14].XIC[6].icell.Ien Iout.t97 VGND.t757 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X907 XA.XIR[15].XIC[8].icell.PDM XThR.Tn[14].t29 VGND.t326 VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X908 VGND.t265 Vbias.t84 XA.XIR[5].XIC[14].icell.SM VGND.t264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X909 VGND.t85 XA.Cn[13].t24 XA.XIR[5].XIC[13].icell.PDM VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X910 VPWR.t1838 thermo15c_0.XTB5.A thermo15c_0.XTB1.Y.t2 VPWR.t1837 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X911 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1972 XA.XIR[5].XIC_dummy_left.icell.Ien VGND.t2247 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X912 VGND.t87 XA.Cn[13].t25 XA.XIR[9].XIC[13].icell.PDM VGND.t86 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X913 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t1973 XA.XIR[9].XIC_dummy_left.icell.Ien VGND.t2248 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X914 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[1].t32 VGND.t1987 VGND.t1986 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X915 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11].t33 XA.XIR[11].XIC[11].icell.Ien VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X916 VGND.t267 Vbias.t85 XA.XIR[1].XIC[11].icell.SM VGND.t266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X917 XA.XIR[4].XIC[1].icell.Ien XThR.Tn[4].t34 VPWR.t1604 VPWR.t1603 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X918 VGND.t269 Vbias.t86 XA.XIR[0].XIC[12].icell.SM VGND.t268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X919 XA.XIR[3].XIC[2].icell.Ien XThR.Tn[3].t34 VPWR.t1059 VPWR.t1058 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X920 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12].t36 XA.XIR[12].XIC_15.icell.Ien VGND.t112 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X921 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t825 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t826 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X922 XA.XIR[2].XIC[14].icell.Ien XThR.Tn[2].t31 VPWR.t1172 VPWR.t1171 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X923 XA.XIR[3].XIC[8].icell.SM XA.XIR[3].XIC[8].icell.Ien Iout.t192 VGND.t1456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X924 VGND.t874 thermo15c_0.XTB3.Y.t6 XA.Cn[2].t1 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X925 XA.XIR[14].XIC[5].icell.PUM XA.Cn[5].t19 XA.XIR[14].XIC[5].icell.Ien VPWR.t1440 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X926 a_8739_9569# thermo15c_0.XTB3.Y.t7 XA.Cn[10].t6 VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X927 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8].t35 XA.XIR[8].XIC[1].icell.Ien VGND.t1071 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X928 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[4].t35 XA.XIR[4].XIC[4].icell.Ien VGND.t1946 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X929 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[3].t35 XA.XIR[3].XIC[5].icell.Ien VGND.t912 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X930 a_n1319_6405# XThR.XTB5.A VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X931 VPWR.t193 XThR.Tn[14].t30 XA.XIR[15].XIC[4].icell.PUM VPWR.t192 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X932 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11].t34 XA.XIR[11].XIC[2].icell.Ien VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X933 XA.XIR[7].XIC[7].icell.PUM XA.Cn[7].t16 XA.XIR[7].XIC[7].icell.Ien VPWR.t1087 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X934 VPWR.t824 VPWR.t822 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t823 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X935 XA.XIR[6].XIC[3].icell.SM XA.XIR[6].XIC[3].icell.Ien Iout.t114 VGND.t878 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X936 a_2979_9615# thermo15c_0.XTB1.Y.t8 VPWR.t263 VPWR.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X937 XA.XIR[0].XIC[13].icell.Ien XThR.Tn[0].t33 VPWR.t992 VPWR.t991 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X938 VGND.t271 Vbias.t87 XA.XIR[15].XIC[2].icell.SM VGND.t270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X939 VGND.t273 Vbias.t88 XA.XIR[14].XIC[3].icell.SM VGND.t272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X940 XThR.Tn[12].t10 XThR.XTBN.Y VPWR.t1821 VPWR.t1820 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X941 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout VGND.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X942 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t819 VPWR.t821 VPWR.t820 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X943 XA.XIR[14].XIC[10].icell.SM XA.XIR[14].XIC[10].icell.Ien Iout.t85 VGND.t695 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X944 XA.Cn[11].t5 thermo15c_0.XTBN.Y.t39 VPWR.t421 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X945 VGND.t542 data[4].t2 XThR.XTB5.A VGND.t541 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X946 XThR.XTBN.Y XThR.XTBN.A VGND.t2609 VGND.t2608 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X947 VGND.t686 data[3].t0 thermo15c_0.XTBN.A VGND.t685 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X948 VGND.t275 Vbias.t89 XA.XIR[1].XIC[9].icell.SM VGND.t274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X949 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1974 VGND.t2250 VGND.t2249 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X950 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[8].t36 VGND.t708 VGND.t707 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X951 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t3 VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X952 XA.XIR[15].XIC[3].icell.PDM XThR.Tn[14].t31 VGND.t328 VGND.t327 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X953 XA.XIR[14].XIC[1].icell.SM XA.XIR[14].XIC[1].icell.Ien Iout.t1 VGND.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X954 XA.XIR[10].XIC_15.icell.PDM VPWR.t1975 VGND.t2252 VGND.t2251 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X955 XA.XIR[9].XIC[13].icell.SM XA.XIR[9].XIC[13].icell.Ien Iout.t57 VGND.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X956 a_n997_2667# XThR.XTBN.Y VGND.t2434 VGND.t2393 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X957 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t817 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t818 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X958 XA.XIR[12].XIC[14].icell.SM XA.XIR[12].XIC[14].icell.Ien Iout.t27 VGND.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X959 XA.XIR[1].XIC[6].icell.PUM XA.Cn[6].t24 XA.XIR[1].XIC[6].icell.Ien VPWR.t428 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X960 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[1].t33 VGND.t1989 VGND.t1988 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X961 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11].t35 XA.XIR[11].XIC[6].icell.Ien VGND.t811 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X962 XA.XIR[7].XIC[11].icell.PUM XA.Cn[11].t21 XA.XIR[7].XIC[11].icell.Ien VPWR.t1000 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X963 XA.XIR[4].XIC[7].icell.PUM XA.Cn[7].t17 XA.XIR[4].XIC[7].icell.Ien VPWR.t1088 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X964 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[4].t36 VGND.t1948 VGND.t1947 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X965 VPWR.t195 XThR.Tn[14].t32 XA.XIR[15].XIC[0].icell.PUM VPWR.t194 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X966 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[8].t37 VGND.t710 VGND.t709 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X967 XA.XIR[3].XIC[8].icell.PUM XA.Cn[8].t21 XA.XIR[3].XIC[8].icell.Ien VPWR.t1100 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X968 VGND.t1184 XA.Cn[9].t23 XA.XIR[1].XIC[9].icell.PDM VGND.t1183 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X969 XA.XIR[3].XIC[3].icell.SM XA.XIR[3].XIC[3].icell.Ien Iout.t185 VGND.t1404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X970 XA.Cn[4].t6 thermo15c_0.XTBN.Y.t40 a_5155_9615# VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X971 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[3].t36 XA.XIR[3].XIC[0].icell.Ien VGND.t920 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X972 VGND.t2254 VPWR.t1976 XA.XIR[12].XIC_15.icell.PDM VGND.t2253 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X973 VPWR.t40 XThR.Tn[12].t37 XA.XIR[13].XIC[9].icell.PUM VPWR.t39 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X974 VPWR.t1819 XThR.XTBN.Y XThR.Tn[8].t10 VPWR.t1818 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X975 VGND.t172 XA.Cn[14].t20 XA.XIR[11].XIC[14].icell.PDM VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X976 VGND.t1054 XA.Cn[8].t22 XA.XIR[11].XIC[8].icell.PDM VGND.t1053 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X977 XA.XIR[7].XIC[2].icell.PUM XA.Cn[2].t21 XA.XIR[7].XIC[2].icell.Ien VPWR.t121 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X978 XA.XIR[2].XIC[14].icell.PUM XA.Cn[14].t21 XA.XIR[2].XIC[14].icell.Ien VPWR.t84 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X979 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t814 VPWR.t816 VPWR.t815 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X980 a_7651_9569# thermo15c_0.XTB1.Y.t9 XA.Cn[8].t5 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X981 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[2].t32 XA.XIR[2].XIC[12].icell.Ien VGND.t1570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X982 VGND.t277 Vbias.t90 XA.XIR[4].XIC[5].icell.SM VGND.t276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X983 VPWR.t340 thermo15c_0.XTB5.Y XA.Cn[12].t1 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X984 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t1977 XA.XIR[14].XIC_dummy_right.icell.Ien VGND.t2265 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X985 VPWR.t961 XThR.Tn[11].t36 XA.XIR[12].XIC[13].icell.PUM VPWR.t960 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X986 VPWR.t813 VPWR.t811 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t812 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X987 VGND.t279 Vbias.t91 XA.XIR[7].XIC[6].icell.SM VGND.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X988 XA.XIR[6].XIC[7].icell.Ien XThR.Tn[6].t30 VPWR.t237 VPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X989 XA.XIR[5].XIC[8].icell.Ien XThR.Tn[5].t32 VPWR.t1292 VPWR.t1291 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X990 VGND.t2021 XA.Cn[5].t20 XA.XIR[7].XIC[5].icell.PDM VGND.t2020 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X991 VGND.t2433 XThR.XTBN.Y XThR.Tn[1].t11 VGND.t2391 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X992 XA.XIR[15].XIC[7].icell.PDM XThR.Tn[14].t33 VGND.t330 VGND.t329 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X993 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[5].t33 VGND.t1266 VGND.t1265 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X994 XA.XIR[9].XIC[8].icell.Ien XThR.Tn[9].t32 VPWR.t349 VPWR.t348 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X995 VPWR.t1472 VGND.t2692 XA.XIR[0].XIC[7].icell.PUM VPWR.t1471 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X996 VPWR.t810 VPWR.t808 XA.XIR[4].XIC_15.icell.PUM VPWR.t809 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X997 XA.XIR[0].XIC[6].icell.Ien XThR.Tn[0].t34 VPWR.t994 VPWR.t993 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X998 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13].t28 XA.XIR[13].XIC[14].icell.Ien VGND.t1008 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X999 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13].t29 XA.XIR[13].XIC[8].icell.Ien VGND.t1009 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1000 VGND.t281 Vbias.t92 XA.XIR[1].XIC[4].icell.SM VGND.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1001 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[2].t33 VGND.t1569 VGND.t1568 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1002 XThR.Tn[6].t2 XThR.XTB7.Y VGND.t889 VGND.t888 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1003 a_9827_9569# thermo15c_0.XTBN.Y.t41 VGND.t438 VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1004 XA.XIR[4].XIC[11].icell.PUM XA.Cn[11].t22 XA.XIR[4].XIC[11].icell.Ien VPWR.t1001 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1005 XThR.Tn[9].t9 XThR.XTBN.Y VPWR.t1817 VPWR.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1006 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[8].t38 VGND.t712 VGND.t711 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1007 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[5].t34 VGND.t1268 VGND.t1267 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1008 XA.XIR[11].XIC[9].icell.PUM XA.Cn[9].t24 XA.XIR[11].XIC[9].icell.Ien VPWR.t1003 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1009 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout VGND.t1161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1010 XA.XIR[5].XIC[11].icell.SM XA.XIR[5].XIC[11].icell.Ien Iout.t239 VGND.t2149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1011 XA.XIR[0].XIC[9].icell.PDM XThR.Tn[0].t35 XA.XIR[0].XIC[9].icell.Ien VGND.t842 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1012 XA.Cn[1].t2 thermo15c_0.XTBN.Y.t42 a_3773_9615# VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1013 VGND.t857 XA.Cn[11].t23 XA.XIR[8].XIC[11].icell.PDM VGND.t856 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1014 XThR.Tn[0].t10 XThR.XTBN.Y VGND.t2432 VGND.t2373 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1015 XA.Cn[13].t5 thermo15c_0.XTB6.Y a_10051_9569# VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1016 XA.XIR[1].XIC[1].icell.PUM XA.Cn[1].t25 XA.XIR[1].XIC[1].icell.Ien VPWR.t1881 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1017 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[2].t34 XA.XIR[2].XIC[10].icell.Ien VGND.t2603 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1018 XA.XIR[4].XIC[2].icell.PUM XA.Cn[2].t22 XA.XIR[4].XIC[2].icell.Ien VPWR.t122 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1019 VPWR.t1816 XThR.XTBN.Y XThR.Tn[10].t10 VPWR.t1815 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1020 VPWR.t351 XThR.Tn[9].t33 XA.XIR[10].XIC[9].icell.PUM VPWR.t350 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1021 XA.XIR[3].XIC[3].icell.PUM XA.Cn[3].t22 XA.XIR[3].XIC[3].icell.Ien VPWR.t1854 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1022 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[4].t37 VGND.t1950 VGND.t1949 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1023 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t805 VPWR.t807 VPWR.t806 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1024 XA.XIR[0].XIC[12].icell.PDM VGND.t1722 VGND.t1724 VGND.t1723 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1025 VGND.t59 XA.Cn[4].t25 XA.XIR[1].XIC[4].icell.PDM VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1026 VGND.t2559 XA.Cn[1].t26 XA.XIR[5].XIC[1].icell.PDM VGND.t2558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1027 VGND.t283 Vbias.t93 XA.XIR[11].XIC[7].icell.SM VGND.t282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1028 VGND.t285 Vbias.t94 XA.XIR[7].XIC[10].icell.SM VGND.t284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1029 XA.XIR[6].XIC[11].icell.Ien XThR.Tn[6].t31 VPWR.t239 VPWR.t238 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1030 VPWR.t1352 thermo15c_0.XTB7.Y a_6243_9615# VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1031 XA.XIR[2].XIC[11].icell.SM XA.XIR[2].XIC[11].icell.Ien Iout.t200 VGND.t1503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1032 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1978 VGND.t2267 VGND.t2266 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1033 VGND.t2561 XA.Cn[1].t27 XA.XIR[9].XIC[1].icell.PDM VGND.t2560 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1034 VGND.t2023 XA.Cn[5].t21 XA.XIR[4].XIC[5].icell.PDM VGND.t2022 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1035 XA.XIR[13].XIC[9].icell.Ien XThR.Tn[13].t30 VPWR.t1085 VPWR.t1084 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1036 VGND.t219 XA.Cn[2].t23 XA.XIR[8].XIC[2].icell.PDM VGND.t218 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1037 VPWR.t1470 VGND.t2693 XA.XIR[0].XIC[11].icell.PUM VPWR.t1469 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1038 VGND.t2525 XA.Cn[3].t23 XA.XIR[11].XIC[3].icell.PDM VGND.t2524 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1039 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10].t30 XA.XIR[10].XIC[11].icell.Ien VGND.t1776 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1040 VGND.t2269 VPWR.t1979 XA.XIR[6].XIC_15.icell.PDM VGND.t2268 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1041 VGND.t439 thermo15c_0.XTBN.Y.t43 a_8963_9569# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1042 VGND.t1236 Vbias.t95 XA.XIR[4].XIC[0].icell.SM VGND.t1235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1043 XA.XIR[15].XIC[4].icell.PUM XA.Cn[4].t26 XA.XIR[15].XIC[4].icell.Ien VPWR.t19 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1044 VPWR.t1372 XThR.XTB1.Y XThR.Tn[8].t3 VPWR.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1045 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t803 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t804 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1046 VGND.t1238 Vbias.t96 XA.XIR[7].XIC[1].icell.SM VGND.t1237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1047 VGND.t1240 Vbias.t97 XA.XIR[2].XIC[13].icell.SM VGND.t1239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1048 XA.XIR[6].XIC[2].icell.Ien XThR.Tn[6].t32 VPWR.t1858 VPWR.t1857 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1049 XA.XIR[11].XIC[5].icell.SM XA.XIR[11].XIC[5].icell.Ien Iout.t36 VGND.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1050 VGND.t1931 XA.Cn[0].t21 XA.XIR[7].XIC[0].icell.PDM VGND.t1930 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1051 XA.XIR[1].XIC[14].icell.Ien XThR.Tn[1].t34 VPWR.t125 VPWR.t124 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1052 XA.XIR[5].XIC[3].icell.Ien XThR.Tn[5].t35 VPWR.t1342 VPWR.t1341 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1053 VGND.t2648 XA.Cn[12].t21 XA.XIR[2].XIC[12].icell.PDM VGND.t2647 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1054 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[5].t36 VGND.t1380 VGND.t1379 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1055 XThR.XTBN.A data[7].t0 VPWR.t526 VPWR.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1056 XA.XIR[9].XIC[3].icell.Ien XThR.Tn[9].t34 VPWR.t353 VPWR.t352 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1057 XA.XIR[4].XIC_15.icell.Ien XThR.Tn[4].t38 VPWR.t1606 VPWR.t1605 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1058 XA.XIR[5].XIC[9].icell.SM XA.XIR[5].XIC[9].icell.Ien Iout.t45 VGND.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1059 a_6243_10571# thermo15c_0.XTB7.B thermo15c_0.XTB7.Y VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1060 VPWR.t1468 VGND.t2694 XA.XIR[0].XIC[2].icell.PUM VPWR.t1467 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1061 VPWR.t1667 XThR.XTB2.Y a_n1049_7787# VPWR.t1355 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1062 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10].t31 XA.XIR[10].XIC[2].icell.Ien VGND.t1777 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1063 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6].t33 XA.XIR[6].XIC[5].icell.Ien VGND.t2531 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1064 XA.XIR[0].XIC[1].icell.Ien XThR.Tn[0].t36 VPWR.t64 VPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1065 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13].t31 XA.XIR[13].XIC[3].icell.Ien VGND.t1010 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1066 VPWR.t963 XThR.Tn[11].t37 XA.XIR[12].XIC[6].icell.PUM VPWR.t962 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1067 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8].t39 XA.XIR[8].XIC_15.icell.Ien VGND.t713 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1068 XA.XIR[0].XIC[7].icell.SM XA.XIR[0].XIC[7].icell.Ien Iout.t81 VGND.t667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1069 XA.XIR[0].XIC[10].icell.PDM VGND.t1719 VGND.t1721 VGND.t1720 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1070 XA.XIR[0].XIC[4].icell.PDM XThR.Tn[0].t37 XA.XIR[0].XIC[4].icell.Ien VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1071 VGND.t1242 Vbias.t98 XA.XIR[8].XIC[7].icell.SM VGND.t1241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1072 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t6 VPWR.t1814 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1073 XA.XIR[2].XIC[9].icell.SM XA.XIR[2].XIC[9].icell.Ien Iout.t38 VGND.t173 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1074 VGND.t512 XA.Cn[6].t25 XA.XIR[8].XIC[6].icell.PDM VGND.t511 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1075 XA.Cn[8].t2 thermo15c_0.XTB1.Y.t10 VPWR.t265 VPWR.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1076 VPWR.t1513 XThR.Tn[10].t32 XA.XIR[11].XIC[4].icell.PUM VPWR.t1512 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1077 VPWR.t802 VPWR.t800 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t801 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1078 VGND.t1718 VGND.t1716 XA.XIR[15].XIC_dummy_right.icell.SM VGND.t1717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1079 VGND.t1015 XA.Cn[7].t18 XA.XIR[11].XIC[7].icell.PDM VGND.t1014 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1080 XThR.Tn[0].t2 XThR.XTB1.Y VGND.t1421 VGND.t1420 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1081 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7].t25 XA.XIR[7].XIC[11].icell.Ien VGND.t733 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1082 VGND.t1244 Vbias.t99 XA.XIR[11].XIC[2].icell.SM VGND.t1243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1083 XA.XIR[15].XIC[0].icell.PUM XA.Cn[0].t22 XA.XIR[15].XIC[0].icell.Ien VPWR.t1591 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1084 VPWR.t1245 XThR.XTB3.Y.t8 XThR.Tn[10].t4 VPWR.t1244 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1085 VGND.t1440 XA.Cn[10].t22 XA.XIR[2].XIC[10].icell.PDM VGND.t1439 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1086 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[7].t26 VGND.t735 VGND.t734 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1087 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[7].t27 VGND.t371 VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1088 XA.XIR[8].XIC[5].icell.SM XA.XIR[8].XIC[5].icell.Ien Iout.t213 VGND.t1780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1089 VPWR.t1596 thermo15c_0.XTB2.Y a_3773_9615# VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1090 VGND.t1933 XA.Cn[0].t23 XA.XIR[4].XIC[0].icell.PDM VGND.t1932 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1091 VGND.t2431 XThR.XTBN.Y XThR.Tn[4].t6 VGND.t2430 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1092 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t798 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t799 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1093 XA.XIR[7].XIC[6].icell.SM XA.XIR[7].XIC[6].icell.Ien Iout.t149 VGND.t1121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1094 XA.XIR[14].XIC[14].icell.PUM XA.Cn[14].t22 XA.XIR[14].XIC[14].icell.Ien VPWR.t1657 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1095 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10].t33 XA.XIR[10].XIC[6].icell.Ien VGND.t1778 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1096 VPWR.t365 thermo15c_0.XTBN.Y.t44 XA.Cn[9].t3 VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1097 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t1980 XA.XIR[2].XIC_dummy_left.icell.Ien VGND.t2270 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1098 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7].t28 XA.XIR[7].XIC[2].icell.Ien VGND.t372 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1099 VGND.t441 thermo15c_0.XTBN.Y.t45 XA.Cn[5].t9 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1100 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[3].t37 VGND.t922 VGND.t921 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1101 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13].t32 XA.XIR[13].XIC[7].icell.Ien VGND.t1011 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1102 XA.XIR[11].XIC[0].icell.SM XA.XIR[11].XIC[0].icell.Ien Iout.t244 VGND.t2474 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1103 XA.XIR[6].XIC[12].icell.SM XA.XIR[6].XIC[12].icell.Ien Iout.t41 VGND.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1104 VGND.t2429 XThR.XTBN.Y a_n997_1579# VGND.t2412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1105 XA.XIR[13].XIC[12].icell.PUM XA.Cn[12].t22 XA.XIR[13].XIC[12].icell.Ien VPWR.t57 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1106 XA.XIR[5].XIC[4].icell.SM XA.XIR[5].XIC[4].icell.Ien Iout.t66 VGND.t463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1107 VGND.t1246 Vbias.t100 XA.XIR[14].XIC[12].icell.SM VGND.t1245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1108 VGND.t1248 Vbias.t101 XA.XIR[10].XIC_15.icell.SM VGND.t1247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1109 a_2979_9615# thermo15c_0.XTBN.Y.t46 XA.Cn[0].t4 VPWR.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1110 VGND.t1991 XA.Cn[14].t23 XA.XIR[10].XIC[14].icell.PDM VGND.t1990 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1111 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6].t34 XA.XIR[6].XIC[0].icell.Ien VGND.t2532 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1112 VGND.t1056 XA.Cn[8].t23 XA.XIR[10].XIC[8].icell.PDM VGND.t1055 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1113 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[1].t35 XA.XIR[1].XIC[12].icell.Ien VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1114 VPWR.t965 XThR.Tn[11].t38 XA.XIR[12].XIC[1].icell.PUM VPWR.t964 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1115 XA.XIR[0].XIC[7].icell.PUM XA.Cn[7].t19 XA.XIR[0].XIC[7].icell.Ien VPWR.t1089 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1116 XA.Cn[12].t6 thermo15c_0.XTB5.Y a_9827_9569# VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1117 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[4].t39 XA.XIR[4].XIC[13].icell.Ien VGND.t2073 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1118 VPWR.t1515 XThR.Tn[10].t34 XA.XIR[11].XIC[0].icell.PUM VPWR.t1514 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1119 XThR.XTB6.A data[5].t2 VPWR.t1742 VPWR.t1741 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1120 XA.XIR[0].XIC[2].icell.SM XA.XIR[0].XIC[2].icell.Ien Iout.t174 VGND.t1373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1121 VPWR.t797 VPWR.t795 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t796 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1122 XThR.Tn[14].t5 XThR.XTB7.Y a_n997_715# VGND.t887 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1123 VPWR.t197 XThR.Tn[14].t34 XA.XIR[15].XIC[13].icell.PUM VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1124 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t7 VPWR.t1812 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1125 XA.XIR[11].XIC[4].icell.Ien XThR.Tn[11].t39 VPWR.t967 VPWR.t966 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1126 VGND.t1250 Vbias.t102 XA.XIR[8].XIC[2].icell.SM VGND.t1249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1127 XA.XIR[2].XIC[4].icell.SM XA.XIR[2].XIC[4].icell.Ien Iout.t241 VGND.t2161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1128 XA.XIR[15].XIC[12].icell.Ien VPWR.t792 VPWR.t794 VPWR.t793 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1129 XA.XIR[7].XIC[10].icell.SM XA.XIR[7].XIC[10].icell.Ien Iout.t203 VGND.t1506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1130 XA.XIR[15].XIC[7].icell.SM XA.XIR[15].XIC[7].icell.Ien Iout.t145 VGND.t1115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1131 VPWR.t127 XThR.Tn[1].t36 XA.XIR[2].XIC[8].icell.PUM VPWR.t126 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1132 VPWR.t519 XThR.Tn[8].t40 XA.XIR[9].XIC[12].icell.PUM VPWR.t518 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1133 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7].t29 XA.XIR[7].XIC[6].icell.Ien VGND.t373 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1134 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1981 VGND.t2272 VGND.t2271 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1135 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[0].t38 VGND.t140 VGND.t139 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1136 XA.XIR[10].XIC[9].icell.PUM XA.Cn[9].t25 XA.XIR[10].XIC[9].icell.Ien VPWR.t1004 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1137 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[7].t30 VGND.t375 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1138 XA.XIR[8].XIC[0].icell.SM XA.XIR[8].XIC[0].icell.Ien Iout.t2 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1139 XA.XIR[3].XIC[12].icell.SM XA.XIR[3].XIC[12].icell.Ien Iout.t129 VGND.t1036 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1140 XA.XIR[3].XIC_15.icell.PDM VPWR.t1982 VGND.t2274 VGND.t2273 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1141 XA.XIR[13].XIC[10].icell.PUM XA.Cn[10].t23 XA.XIR[13].XIC[10].icell.Ien VPWR.t1382 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1142 XA.XIR[7].XIC[1].icell.SM XA.XIR[7].XIC[1].icell.Ien Iout.t108 VGND.t826 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1143 a_6243_9615# thermo15c_0.XTB7.Y VPWR.t1351 VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1144 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t790 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t791 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1145 VGND.t1715 VGND.t1713 XA.XIR[15].XIC_dummy_left.icell.SM VGND.t1714 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1146 XA.Cn[10].t0 thermo15c_0.XTBN.Y.t47 VPWR.t368 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1147 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[1].t37 XA.XIR[1].XIC[10].icell.Ien VGND.t225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1148 XA.XIR[0].XIC[11].icell.PUM XA.Cn[11].t24 XA.XIR[0].XIC[11].icell.Ien VPWR.t1002 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1149 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[3].t38 VGND.t924 VGND.t923 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1150 VGND.t124 XA.Cn[12].t23 XA.XIR[14].XIC[12].icell.PDM VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1151 XA.XIR[1].XIC_15.icell.PUM VPWR.t788 XA.XIR[1].XIC_15.icell.Ien VPWR.t789 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1152 XA.Cn[10].t7 thermo15c_0.XTB3.Y.t8 a_8739_9569# VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1153 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[1].t38 VGND.t227 VGND.t226 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1154 VGND.t1398 thermo15c_0.XTB7.Y XA.Cn[6].t11 VGND.t1397 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1155 XA.XIR[1].XIC[11].icell.SM XA.XIR[1].XIC[11].icell.Ien Iout.t133 VGND.t1058 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1156 VGND.t2276 VPWR.t1983 XA.XIR[2].XIC_dummy_left.icell.PDM VGND.t2275 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1157 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1984 VGND.t2278 VGND.t2277 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1158 XThR.Tn[11].t10 XThR.XTBN.Y VPWR.t1813 VPWR.t1794 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1159 VGND.t2527 XA.Cn[3].t24 XA.XIR[10].XIC[3].icell.PDM VGND.t2526 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1160 VPWR.t369 thermo15c_0.XTBN.Y.t48 XA.Cn[12].t11 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1161 VGND.t2280 VPWR.t1985 XA.XIR[5].XIC_15.icell.PDM VGND.t2279 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1162 XA.XIR[15].XIC[10].icell.Ien VPWR.t785 VPWR.t787 VPWR.t786 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1163 VGND.t1252 Vbias.t103 XA.XIR[13].XIC[11].icell.SM VGND.t1251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1164 XA.XIR[12].XIC[12].icell.Ien XThR.Tn[12].t38 VPWR.t42 VPWR.t41 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1165 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11].t40 VPWR.t969 VPWR.t968 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1166 VGND.t2282 VPWR.t1986 XA.XIR[9].XIC_15.icell.PDM VGND.t2281 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1167 VPWR.t1344 XThR.Tn[5].t37 XA.XIR[6].XIC[9].icell.PUM VPWR.t1343 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1168 XA.XIR[0].XIC[2].icell.PUM XA.Cn[2].t24 XA.XIR[0].XIC[2].icell.Ien VPWR.t123 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1169 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t782 VPWR.t784 VPWR.t783 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1170 VPWR.t521 XThR.Tn[8].t41 XA.XIR[9].XIC[10].icell.PUM VPWR.t520 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1171 VGND.t1254 Vbias.t104 XA.XIR[1].XIC[13].icell.SM VGND.t1253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1172 VGND.t1256 Vbias.t105 XA.XIR[0].XIC[6].icell.SM VGND.t1255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1173 VGND.t2025 XA.Cn[5].t22 XA.XIR[0].XIC[5].icell.PDM VGND.t2024 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1174 VGND.t1258 Vbias.t106 XA.XIR[4].XIC[14].icell.SM VGND.t1257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1175 VGND.t2160 thermo15c_0.XTB7.A thermo15c_0.XTB7.Y VGND.t2159 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1176 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[7].t31 VGND.t377 VGND.t376 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1177 XA.XIR[2].XIC[8].icell.Ien XThR.Tn[2].t35 VPWR.t1170 VPWR.t1169 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1178 VPWR.t129 XThR.Tn[1].t39 XA.XIR[2].XIC[3].icell.PUM VPWR.t128 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1179 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t2 VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1180 XA.XIR[15].XIC[2].icell.SM XA.XIR[15].XIC[2].icell.Ien Iout.t79 VGND.t640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1181 a_n997_2667# XThR.XTBN.Y VGND.t2428 VGND.t2383 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1182 VPWR.t390 XThR.Tn[14].t35 XA.XIR[15].XIC[6].icell.PUM VPWR.t389 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1183 VPWR.t486 XThR.Tn[13].t33 XA.XIR[14].XIC[7].icell.PUM VPWR.t485 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1184 a_7875_9569# thermo15c_0.XTBN.Y.t49 VGND.t442 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1185 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[0].t39 VGND.t142 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1186 VGND.t1442 XA.Cn[10].t24 XA.XIR[14].XIC[10].icell.PDM VGND.t1441 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1187 VGND.t2427 XThR.XTBN.Y a_n997_3979# VGND.t2426 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1188 XA.XIR[0].XIC_15.icell.Ien XThR.Tn[0].t40 VPWR.t66 VPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1189 XA.XIR[1].XIC[9].icell.SM XA.XIR[1].XIC[9].icell.Ien Iout.t178 VGND.t1377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1190 XA.XIR[13].XIC[5].icell.PUM XA.Cn[5].t23 XA.XIR[13].XIC[5].icell.Ien VPWR.t1678 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1191 XA.Cn[14].t2 thermo15c_0.XTBN.Y.t50 VPWR.t371 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1192 a_n1049_6699# XThR.XTB4.Y.t7 VPWR.t1283 VPWR.t1232 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1193 a_4861_9615# thermo15c_0.XTBN.Y.t51 XA.Cn[3].t7 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1194 VGND.t642 Vbias.t107 XA.XIR[10].XIC[8].icell.SM VGND.t641 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1195 VGND.t1017 XA.Cn[7].t20 XA.XIR[10].XIC[7].icell.PDM VGND.t1016 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1196 VGND.t644 Vbias.t108 XA.XIR[13].XIC[9].icell.SM VGND.t643 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1197 XA.XIR[12].XIC[10].icell.Ien XThR.Tn[12].t39 VPWR.t44 VPWR.t43 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1198 XA.Cn[2].t10 thermo15c_0.XTB3.Y.t9 VGND.t1575 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1199 XA.Cn[9].t2 thermo15c_0.XTBN.Y.t52 VPWR.t386 VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1200 XA.Cn[5].t8 thermo15c_0.XTBN.Y.t53 VGND.t464 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1201 a_n1335_8107# XThR.XTB6.A XThR.XTB2.Y VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1202 VGND.t646 Vbias.t109 XA.XIR[0].XIC[10].icell.SM VGND.t645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1203 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[13].t34 VGND.t672 VGND.t671 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1204 VGND.t89 XA.Cn[13].t26 XA.XIR[1].XIC[13].icell.PDM VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1205 XA.XIR[15].XIC[5].icell.Ien VPWR.t779 VPWR.t781 VPWR.t780 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1206 VGND.t1712 VGND.t1710 XA.XIR[11].XIC_dummy_right.icell.SM VGND.t1711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1207 VPWR.t141 thermo15c_0.XTB1.Y.t11 a_2979_9615# VPWR.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1208 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1987 XA.XIR[1].XIC_dummy_left.icell.Ien VGND.t2283 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1209 XA.Cn[0].t3 thermo15c_0.XTBN.Y.t54 a_2979_9615# VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1210 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[3].t39 XA.XIR[3].XIC[11].icell.Ien VGND.t925 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1211 VPWR.t523 XThR.Tn[8].t42 XA.XIR[9].XIC[5].icell.PUM VPWR.t522 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1212 VPWR.t488 XThR.Tn[13].t35 XA.XIR[14].XIC[11].icell.PUM VPWR.t487 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1213 XThR.Tn[12].t5 XThR.XTB5.Y VPWR.t1235 VPWR.t1234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1214 XA.XIR[8].XIC[4].icell.PUM XA.Cn[4].t27 XA.XIR[8].XIC[4].icell.Ien VPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1215 XA.XIR[12].XIC[12].icell.PUM XA.Cn[12].t24 XA.XIR[12].XIC[12].icell.Ien VPWR.t58 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1216 VGND.t648 Vbias.t110 XA.XIR[0].XIC[1].icell.SM VGND.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1217 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t777 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t778 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1218 XA.XIR[4].XIC[5].icell.SM XA.XIR[4].XIC[5].icell.Ien Iout.t83 VGND.t670 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1219 VGND.t1935 XA.Cn[0].t24 XA.XIR[0].XIC[0].icell.PDM VGND.t1934 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1220 XThR.Tn[6].t10 XThR.XTBN.Y VGND.t2425 VGND.t2424 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1221 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t6 VPWR.t1812 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1222 XA.XIR[15].XIC[13].icell.PUM XA.Cn[13].t27 XA.XIR[15].XIC[13].icell.Ien VPWR.t26 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1223 VGND.t2423 XThR.XTBN.Y a_n997_2891# VGND.t2422 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1224 VGND.t1136 XThR.XTB7.B XThR.XTB7.Y VGND.t1135 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1225 XA.XIR[2].XIC[3].icell.Ien XThR.Tn[2].t36 VPWR.t1168 VPWR.t1167 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1226 XA.XIR[11].XIC[14].icell.SM XA.XIR[11].XIC[14].icell.Ien Iout.t91 VGND.t739 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1227 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[4].t40 XA.XIR[4].XIC[1].icell.Ien VGND.t2074 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1228 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[3].t40 XA.XIR[3].XIC[2].icell.Ien VGND.t926 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1229 XA.XIR[14].XIC[7].icell.Ien XThR.Tn[14].t36 VPWR.t392 VPWR.t391 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1230 VPWR.t394 XThR.Tn[14].t37 XA.XIR[15].XIC[1].icell.PUM VPWR.t393 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1231 VGND.t2285 VPWR.t1988 XA.XIR[11].XIC_dummy_right.icell.PDM VGND.t2284 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1232 XA.XIR[2].XIC[8].icell.PUM XA.Cn[8].t24 XA.XIR[2].XIC[8].icell.Ien VPWR.t1196 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1233 VPWR.t490 XThR.Tn[13].t36 XA.XIR[14].XIC[2].icell.PUM VPWR.t489 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1234 a_n997_2667# XThR.XTB4.Y.t8 XThR.Tn[11].t4 VGND.t913 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1235 VPWR.t776 VPWR.t774 XA.XIR[12].XIC_15.icell.PUM VPWR.t775 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1236 XA.XIR[1].XIC[4].icell.SM XA.XIR[1].XIC[4].icell.Ien Iout.t219 VGND.t1786 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1237 XA.XIR[10].XIC[4].icell.Ien XThR.Tn[10].t35 VPWR.t1744 VPWR.t1743 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1238 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t771 VPWR.t773 VPWR.t772 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1239 VGND.t650 Vbias.t111 XA.XIR[6].XIC_15.icell.SM VGND.t649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1240 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout VGND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1241 XA.XIR[14].XIC[7].icell.SM XA.XIR[14].XIC[7].icell.Ien Iout.t236 VGND.t2128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1242 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[13].t37 VGND.t674 VGND.t673 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1243 VGND.t652 Vbias.t112 XA.XIR[10].XIC[3].icell.SM VGND.t651 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1244 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t768 VPWR.t770 VPWR.t769 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1245 VGND.t465 thermo15c_0.XTBN.Y.t55 XA.Cn[1].t5 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1246 a_n1049_6405# XThR.XTB5.Y VPWR.t1233 VPWR.t1232 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1247 VGND.t654 Vbias.t113 XA.XIR[13].XIC[4].icell.SM VGND.t653 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1248 XA.XIR[12].XIC[5].icell.Ien XThR.Tn[12].t40 VPWR.t46 VPWR.t45 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1249 VPWR.t269 XThR.Tn[7].t32 XA.XIR[8].XIC[12].icell.PUM VPWR.t268 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1250 XA.XIR[0].XIC[13].icell.PDM XThR.Tn[0].t41 XA.XIR[0].XIC[13].icell.Ien VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1251 VGND.t1709 VGND.t1707 XA.XIR[8].XIC_dummy_right.icell.SM VGND.t1708 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1252 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1989 XA.XIR[13].XIC_dummy_right.icell.Ien VGND.t2286 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1253 VGND.t2288 VPWR.t1990 XA.XIR[14].XIC_dummy_left.icell.PDM VGND.t2287 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1254 VPWR.t1746 XThR.Tn[10].t36 XA.XIR[11].XIC[13].icell.PUM VPWR.t1745 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1255 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[4].t41 VGND.t2076 VGND.t2075 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1256 XA.XIR[12].XIC[10].icell.PUM XA.Cn[10].t25 XA.XIR[12].XIC[10].icell.Ien VPWR.t1383 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1257 VPWR.t1370 XThR.XTB1.Y XThR.Tn[8].t2 VPWR.t1369 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1258 XA.XIR[8].XIC[0].icell.PUM XA.Cn[0].t25 XA.XIR[8].XIC[0].icell.Ien VPWR.t1592 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1259 XA.XIR[5].XIC[13].icell.SM XA.XIR[5].XIC[13].icell.Ien Iout.t93 VGND.t741 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1260 VPWR.t1811 XThR.XTBN.Y XThR.Tn[7].t2 VPWR.t1810 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1261 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t766 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t767 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1262 VGND.t1941 thermo15c_0.XTB2.Y XA.Cn[1].t11 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1263 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t764 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t765 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1264 XA.XIR[8].XIC[14].icell.SM XA.XIR[8].XIC[14].icell.Ien Iout.t72 VGND.t562 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1265 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[3].t41 XA.XIR[3].XIC[6].icell.Ien VGND.t927 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1266 XA.Cn[12].t10 thermo15c_0.XTBN.Y.t56 VPWR.t388 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1267 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[1].t40 VGND.t229 VGND.t228 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1268 XA.XIR[14].XIC[11].icell.Ien XThR.Tn[14].t38 VPWR.t396 VPWR.t395 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1269 VGND.t2001 XThR.XTB2.Y XThR.Tn[1].t2 VGND.t1415 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1270 XThR.Tn[1].t6 XThR.XTBN.Y a_n1049_7787# VPWR.t1790 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1271 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[4].t42 VGND.t2078 VGND.t2077 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1272 XA.XIR[4].XIC[0].icell.SM XA.XIR[4].XIC[0].icell.Ien Iout.t158 VGND.t1160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1273 XA.XIR[6].XIC[12].icell.PUM XA.Cn[12].t25 XA.XIR[6].XIC[12].icell.Ien VPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1274 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[12].t41 VGND.t114 VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1275 VGND.t859 XA.Cn[11].t25 XA.XIR[7].XIC[11].icell.PDM VGND.t858 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1276 XA.XIR[2].XIC[13].icell.SM XA.XIR[2].XIC[13].icell.Ien Iout.t188 VGND.t1427 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1277 XA.XIR[7].XIC[4].icell.Ien XThR.Tn[7].t33 VPWR.t271 VPWR.t270 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1278 VGND.t656 Vbias.t114 XA.XIR[3].XIC_15.icell.SM VGND.t655 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1279 VGND.t658 Vbias.t115 XA.XIR[12].XIC[11].icell.SM VGND.t657 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1280 VGND.t1706 VGND.t1704 XA.XIR[11].XIC_dummy_left.icell.SM VGND.t1705 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1281 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10].t37 VPWR.t1748 VPWR.t1747 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1282 VGND.t1110 XA.Cn[8].t25 XA.XIR[3].XIC[8].icell.PDM VGND.t1109 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1283 VGND.t1993 XA.Cn[14].t24 XA.XIR[3].XIC[14].icell.PDM VGND.t1992 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1284 XA.XIR[14].XIC[2].icell.Ien XThR.Tn[14].t39 VPWR.t398 VPWR.t397 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1285 XThR.Tn[9].t5 XThR.XTB2.Y VPWR.t1666 VPWR.t1226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1286 XThR.Tn[7].t5 XThR.XTBN.Y VGND.t2421 VGND.t2420 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1287 VPWR.t1906 data[1].t2 thermo15c_0.XTB6.A VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1288 XA.XIR[2].XIC[3].icell.PUM XA.Cn[3].t25 XA.XIR[2].XIC[3].icell.Ien VPWR.t1855 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1289 VPWR.t247 XThR.Tn[7].t34 XA.XIR[8].XIC[10].icell.PUM VPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1290 XA.XIR[15].XIC[6].icell.PUM XA.Cn[6].t26 XA.XIR[15].XIC[6].icell.Ien VPWR.t429 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1291 VPWR.t763 VPWR.t761 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t762 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1292 VGND.t466 thermo15c_0.XTBN.Y.t57 a_7875_9569# VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1293 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14].t40 XA.XIR[14].XIC[5].icell.Ien VGND.t471 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1294 VPWR.t1809 XThR.XTBN.Y XThR.Tn[13].t10 VPWR.t1797 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1295 XA.XIR[1].XIC[8].icell.Ien XThR.Tn[1].t41 VPWR.t507 VPWR.t506 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1296 VPWR.t760 VPWR.t758 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t759 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1297 VGND.t221 XA.Cn[2].t25 XA.XIR[7].XIC[2].icell.PDM VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1298 a_8739_10571# data[0].t1 thermo15c_0.XTB7.A VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1299 XA.XIR[14].XIC[2].icell.SM XA.XIR[14].XIC[2].icell.Ien Iout.t228 VGND.t1957 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1300 VGND.t660 Vbias.t116 XA.XIR[9].XIC[11].icell.SM VGND.t659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1301 VPWR.t3 XThR.XTB3.Y.t9 XThR.Tn[10].t0 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1302 XA.XIR[8].XIC[12].icell.Ien XThR.Tn[8].t43 VPWR.t68 VPWR.t67 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1303 VGND.t863 XA.Cn[9].t26 XA.XIR[15].XIC[9].icell.PDM VGND.t862 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1304 XA.Cn[3].t6 thermo15c_0.XTBN.Y.t58 a_4861_9615# VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1305 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5].t38 XA.XIR[5].XIC[8].icell.Ien VGND.t1381 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1306 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5].t39 XA.XIR[5].XIC[14].icell.Ien VGND.t1382 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1307 XA.XIR[11].XIC[13].icell.Ien XThR.Tn[11].t41 VPWR.t971 VPWR.t970 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1308 XThR.Tn[5].t2 XThR.XTB6.Y VGND.t752 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1309 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9].t35 XA.XIR[9].XIC[14].icell.Ien VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1310 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9].t36 XA.XIR[9].XIC[8].icell.Ien VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1311 VPWR.t1215 XThR.XTB7.B XThR.XTB4.Y.t0 VPWR.t1214 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1312 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout VGND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1313 XA.XIR[3].XIC[9].icell.PUM XA.Cn[9].t27 XA.XIR[3].XIC[9].icell.Ien VPWR.t1005 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1314 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[4].t43 VGND.t2080 VGND.t2079 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1315 XA.XIR[12].XIC[5].icell.PUM XA.Cn[5].t24 XA.XIR[12].XIC[5].icell.Ien VPWR.t1679 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1316 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1991 VGND.t2290 VGND.t2289 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1317 XA.XIR[6].XIC[10].icell.PUM XA.Cn[10].t26 XA.XIR[6].XIC[10].icell.Ien VPWR.t1332 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1318 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout VGND.t1146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1319 VGND.t662 Vbias.t117 XA.XIR[12].XIC[9].icell.SM VGND.t661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1320 VGND.t861 XA.Cn[11].t26 XA.XIR[4].XIC[11].icell.PDM VGND.t860 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1321 VPWR.t1750 XThR.Tn[10].t38 XA.XIR[11].XIC[6].icell.PUM VPWR.t1749 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1322 VGND.t1703 VGND.t1701 XA.XIR[8].XIC_dummy_left.icell.SM VGND.t1702 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1323 XA.XIR[7].XIC[0].icell.Ien XThR.Tn[7].t35 VPWR.t249 VPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1324 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t4 VGND.t886 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1325 VGND.t2545 XA.Cn[1].t28 XA.XIR[1].XIC[1].icell.PDM VGND.t2544 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1326 VGND.t664 Vbias.t118 XA.XIR[7].XIC[7].icell.SM VGND.t663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1327 XA.XIR[5].XIC[9].icell.Ien XThR.Tn[5].t40 VPWR.t1346 VPWR.t1345 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1328 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[12].t42 VGND.t116 VGND.t115 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1329 VGND.t514 XA.Cn[6].t27 XA.XIR[7].XIC[6].icell.PDM VGND.t513 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1330 VGND.t1538 Vbias.t119 XA.XIR[6].XIC[8].icell.SM VGND.t1537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1331 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[11].t42 VGND.t676 VGND.t675 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1332 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t1992 VGND.t2292 VGND.t2291 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1333 VGND.t223 XA.Cn[2].t26 XA.XIR[4].XIC[2].icell.PDM VGND.t222 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1334 XA.XIR[9].XIC[9].icell.Ien XThR.Tn[9].t37 VPWR.t355 VPWR.t354 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1335 VGND.t2529 XA.Cn[3].t26 XA.XIR[3].XIC[3].icell.PDM VGND.t2528 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1336 XA.XIR[14].XIC[8].icell.PUM XA.Cn[8].t26 XA.XIR[14].XIC[8].icell.Ien VPWR.t1197 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1337 VGND.t1540 Vbias.t120 XA.XIR[9].XIC[9].icell.SM VGND.t1539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1338 XA.XIR[8].XIC[10].icell.Ien XThR.Tn[8].t44 VPWR.t70 VPWR.t69 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1339 XA.XIR[10].XIC_15.icell.SM XA.XIR[10].XIC_15.icell.Ien Iout.t98 VGND.t771 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1340 VPWR.t251 XThR.Tn[7].t36 XA.XIR[8].XIC[5].icell.PUM VPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1341 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6].t35 XA.XIR[6].XIC[11].icell.Ien VGND.t2533 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1342 XA.XIR[15].XIC[1].icell.PUM XA.Cn[1].t29 XA.XIR[15].XIC[1].icell.Ien VPWR.t1873 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1343 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14].t41 XA.XIR[14].XIC[0].icell.Ien VGND.t472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1344 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[6].t36 VGND.t2535 VGND.t2534 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1345 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[6].t37 VGND.t2537 VGND.t2536 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1346 XA.XIR[1].XIC[3].icell.Ien XThR.Tn[1].t42 VPWR.t509 VPWR.t508 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1347 XA.XIR[6].XIC[6].icell.SM XA.XIR[6].XIC[6].icell.Ien Iout.t173 VGND.t1372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1348 XA.XIR[13].XIC[14].icell.PUM XA.Cn[14].t25 XA.XIR[13].XIC[14].icell.Ien VPWR.t1658 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1349 VGND.t1542 Vbias.t121 XA.XIR[15].XIC[5].icell.SM VGND.t1541 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1350 VGND.t1544 Vbias.t122 XA.XIR[14].XIC[6].icell.SM VGND.t1543 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1351 VGND.t61 XA.Cn[4].t28 XA.XIR[15].XIC[4].icell.PDM VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1352 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6].t38 XA.XIR[6].XIC[2].icell.Ien VGND.t2538 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1353 VGND.t2294 VPWR.t1993 XA.XIR[10].XIC_dummy_right.icell.PDM VGND.t2293 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1354 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5].t41 XA.XIR[5].XIC[3].icell.Ien VGND.t1383 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1355 XA.Cn[1].t4 thermo15c_0.XTBN.Y.t59 VGND.t467 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1356 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9].t38 XA.XIR[9].XIC[3].icell.Ien VGND.t431 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1357 XA.XIR[4].XIC_15.icell.PDM XThR.Tn[4].t44 XA.XIR[4].XIC_15.icell.Ien VGND.t2081 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1358 VPWR.t757 VPWR.t755 XA.XIR[15].XIC_15.icell.PUM VPWR.t756 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1359 XA.XIR[6].XIC[5].icell.PUM XA.Cn[5].t25 XA.XIR[6].XIC[5].icell.Ien VPWR.t1680 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1360 XA.XIR[0].XIC[1].icell.PDM XThR.Tn[0].t42 XA.XIR[0].XIC[1].icell.Ien VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1361 XA.XIR[11].XIC[6].icell.Ien XThR.Tn[11].t43 VPWR.t494 VPWR.t493 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1362 a_7875_9569# thermo15c_0.XTB2.Y XA.Cn[9].t9 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1363 VPWR.t1166 XThR.Tn[2].t37 XA.XIR[3].XIC[4].icell.PUM VPWR.t1165 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1364 VGND.t1546 Vbias.t123 XA.XIR[3].XIC[8].icell.SM VGND.t1545 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1365 VGND.t516 XA.Cn[6].t28 XA.XIR[4].XIC[6].icell.PDM VGND.t515 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1366 XA.XIR[15].XIC[14].icell.Ien VPWR.t752 VPWR.t754 VPWR.t753 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1367 VGND.t1548 Vbias.t124 XA.XIR[12].XIC[4].icell.SM VGND.t1547 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1368 VPWR.t1752 XThR.Tn[10].t39 XA.XIR[11].XIC[1].icell.PUM VPWR.t1751 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1369 VGND.t688 XA.Cn[7].t21 XA.XIR[3].XIC[7].icell.PDM VGND.t687 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1370 VPWR.t1860 XThR.Tn[6].t39 XA.XIR[7].XIC[4].icell.PUM VPWR.t1859 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1371 VPWR.t748 VPWR.t746 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t747 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1372 XThR.Tn[13].t5 XThR.XTB6.Y a_n997_1579# VGND.t750 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1373 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t6 VPWR.t1808 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1374 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout VGND.t1026 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1375 VPWR.t72 XThR.Tn[8].t45 XA.XIR[9].XIC[14].icell.PUM VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1376 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11].t44 XA.XIR[11].XIC[9].icell.Ien VGND.t677 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1377 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[3].t42 VGND.t929 VGND.t928 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1378 VGND.t1550 Vbias.t125 XA.XIR[7].XIC[2].icell.SM VGND.t1549 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1379 VGND.t1552 Vbias.t126 XA.XIR[6].XIC[3].icell.SM VGND.t1551 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1380 XA.XIR[6].XIC[10].icell.SM XA.XIR[6].XIC[10].icell.Ien Iout.t206 VGND.t1519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1381 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[11].t45 VGND.t679 VGND.t678 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1382 XA.XIR[3].XIC[6].icell.SM XA.XIR[3].XIC[6].icell.Ien Iout.t215 VGND.t1782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1383 XA.XIR[14].XIC[3].icell.PUM XA.Cn[3].t27 XA.XIR[14].XIC[3].icell.Ien VPWR.t1856 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1384 VGND.t1554 Vbias.t127 XA.XIR[9].XIC[4].icell.SM VGND.t1553 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1385 XA.XIR[8].XIC[5].icell.Ien XThR.Tn[8].t46 VPWR.t74 VPWR.t73 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1386 VGND.t1556 Vbias.t128 XA.XIR[14].XIC[10].icell.SM VGND.t1555 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1387 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[10].t40 VGND.t2164 VGND.t2163 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1388 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6].t40 XA.XIR[6].XIC[6].icell.Ien VGND.t2539 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1389 VGND.t7 data[2].t1 thermo15c_0.XTB7.B VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1390 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5].t42 XA.XIR[5].XIC[7].icell.Ien VGND.t1384 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1391 VGND.t2419 XThR.XTBN.Y XThR.Tn[2].t10 VGND.t2418 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1392 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[3].t43 VGND.t931 VGND.t930 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1393 XA.XIR[13].XIC[11].icell.SM XA.XIR[13].XIC[11].icell.Ien Iout.t230 VGND.t1974 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1394 a_n1049_5317# XThR.XTB7.Y VPWR.t1019 VPWR.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1395 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9].t39 XA.XIR[9].XIC[7].icell.Ien VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1396 VGND.t468 thermo15c_0.XTBN.Y.t60 XA.Cn[4].t9 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1397 XA.XIR[5].XIC[12].icell.PUM XA.Cn[12].t26 XA.XIR[5].XIC[12].icell.Ien VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1398 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[6].t41 VGND.t2541 VGND.t2540 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1399 XA.XIR[2].XIC_15.icell.PDM VPWR.t1994 VGND.t2296 VGND.t2295 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1400 XA.XIR[6].XIC[1].icell.SM XA.XIR[6].XIC[1].icell.Ien Iout.t249 VGND.t2615 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1401 XA.XIR[1].XIC[13].icell.SM XA.XIR[1].XIC[13].icell.Ien Iout.t58 VGND.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1402 XA.XIR[9].XIC[12].icell.PUM XA.Cn[12].t27 XA.XIR[9].XIC[12].icell.Ien VPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1403 VGND.t1558 Vbias.t129 XA.XIR[15].XIC[0].icell.SM VGND.t1557 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1404 XA.XIR[8].XIC[13].icell.PUM XA.Cn[13].t28 XA.XIR[8].XIC[13].icell.Ien VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1405 VGND.t1560 Vbias.t130 XA.XIR[14].XIC[1].icell.SM VGND.t1559 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1406 VGND.t1577 Vbias.t131 XA.XIR[10].XIC[12].icell.SM VGND.t1576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1407 XA.XIR[4].XIC[14].icell.SM XA.XIR[4].XIC[14].icell.Ien Iout.t254 VGND.t2686 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1408 XThR.Tn[3].t1 XThR.XTB4.Y.t9 VGND.t1259 VGND.t1140 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1409 VGND.t1579 Vbias.t132 XA.XIR[13].XIC[13].icell.SM VGND.t1578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1410 VPWR.t1164 XThR.Tn[2].t38 XA.XIR[3].XIC[0].icell.PUM VPWR.t1163 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1411 VGND.t126 XA.Cn[12].t28 XA.XIR[13].XIC[12].icell.PDM VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1412 XA.XIR[12].XIC[14].icell.Ien XThR.Tn[12].t43 VPWR.t48 VPWR.t47 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1413 VPWR.t1862 XThR.Tn[6].t42 XA.XIR[7].XIC[0].icell.PUM VPWR.t1861 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1414 VPWR.t1350 thermo15c_0.XTB7.Y a_6243_9615# VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1415 VPWR.t1035 thermo15c_0.XTB6.Y XA.Cn[13].t2 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1416 VPWR.t751 VPWR.t749 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t750 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1417 VGND.t1500 data[1].t3 thermo15c_0.XTB5.A VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1418 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[0].t43 VGND.t759 VGND.t758 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1419 XA.XIR[3].XIC[4].icell.Ien XThR.Tn[3].t44 VPWR.t1079 VPWR.t1078 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1420 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[8].t47 VGND.t146 VGND.t145 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1421 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11].t46 VPWR.t496 VPWR.t495 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1422 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t743 VPWR.t745 VPWR.t744 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1423 VGND.t1581 Vbias.t133 XA.XIR[3].XIC[3].icell.SM VGND.t1580 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1424 XA.XIR[7].XIC[7].icell.SM XA.XIR[7].XIC[7].icell.Ien Iout.t147 VGND.t1119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1425 XA.XIR[3].XIC[10].icell.SM XA.XIR[3].XIC[10].icell.Ien Iout.t154 VGND.t1155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1426 XA.XIR[10].XIC[13].icell.Ien XThR.Tn[10].t41 VPWR.t1754 VPWR.t1753 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1427 VPWR.t554 XThR.Tn[0].t44 XA.XIR[1].XIC[12].icell.PUM VPWR.t553 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1428 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[10].t42 VGND.t2166 VGND.t2165 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1429 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout VGND.t543 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1430 XA.XIR[10].XIC[8].icell.SM XA.XIR[10].XIC[8].icell.Ien Iout.t117 VGND.t881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1431 VGND.t470 thermo15c_0.XTBN.Y.t61 XA.Cn[7].t6 VGND.t469 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1432 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[3].t45 VGND.t933 VGND.t932 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1433 VPWR.t1700 XThR.Tn[4].t45 XA.XIR[5].XIC[12].icell.PUM VPWR.t1699 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1434 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11].t47 XA.XIR[11].XIC[4].icell.Ien VGND.t680 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1435 XA.XIR[13].XIC[9].icell.SM XA.XIR[13].XIC[9].icell.Ien Iout.t220 VGND.t1822 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1436 XA.XIR[15].XIC[12].icell.PDM VPWR.t1995 XA.XIR[15].XIC[12].icell.Ien VGND.t2297 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1437 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[0].t45 VGND.t761 VGND.t760 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1438 XA.XIR[5].XIC[10].icell.PUM XA.Cn[10].t27 XA.XIR[5].XIC[10].icell.Ien VPWR.t1333 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1439 XThR.Tn[12].t4 XThR.XTB5.Y VPWR.t1231 VPWR.t1230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1440 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[6].t43 VGND.t2543 VGND.t2542 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1441 a_10915_9569# thermo15c_0.XTBN.Y.t62 VGND.t63 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1442 XA.XIR[3].XIC[1].icell.SM XA.XIR[3].XIC[1].icell.Ien Iout.t166 VGND.t1365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1443 XA.XIR[9].XIC[10].icell.PUM XA.Cn[10].t28 XA.XIR[9].XIC[10].icell.Ien VPWR.t1334 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1444 XThR.Tn[6].t9 XThR.XTBN.Y VGND.t2417 VGND.t2416 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1445 VPWR.t50 XThR.Tn[12].t44 XA.XIR[13].XIC[7].icell.PUM VPWR.t49 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1446 XA.Cn[3].t2 thermo15c_0.XTB4.Y.t7 VGND.t2604 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1447 XA.Cn[9].t5 thermo15c_0.XTB2.Y VPWR.t1595 VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1448 VGND.t1350 XA.Cn[10].t29 XA.XIR[13].XIC[10].icell.PDM VGND.t1349 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1449 a_n997_2667# XThR.XTB4.Y.t10 XThR.Tn[11].t5 VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1450 VGND.t401 XA.Cn[11].t27 XA.XIR[0].XIC[11].icell.PDM VGND.t400 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1451 XA.XIR[15].XIC[5].icell.PDM XThR.Tn[14].t42 VGND.t474 VGND.t473 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1452 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[5].t43 VGND.t1386 VGND.t1385 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1453 VGND.t1583 Vbias.t134 XA.XIR[5].XIC[11].icell.SM VGND.t1582 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1454 XA.XIR[3].XIC[0].icell.Ien XThR.Tn[3].t46 VPWR.t1081 VPWR.t1080 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1455 XA.XIR[9].XIC_15.icell.SM XA.XIR[9].XIC_15.icell.Ien Iout.t175 VGND.t1374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1456 VGND.t2299 VPWR.t1996 XA.XIR[1].XIC_15.icell.PDM VGND.t2298 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1457 VPWR.t511 XThR.Tn[1].t43 XA.XIR[2].XIC[9].icell.PUM VPWR.t510 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1458 VPWR.t556 XThR.Tn[0].t46 XA.XIR[1].XIC[10].icell.PUM VPWR.t555 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1459 XA.XIR[7].XIC[13].icell.Ien XThR.Tn[7].t37 VPWR.t253 VPWR.t252 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1460 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t740 VPWR.t742 VPWR.t741 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1461 VPWR.t1553 XThR.Tn[4].t46 XA.XIR[5].XIC[10].icell.PUM VPWR.t1552 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1462 XA.XIR[15].XIC[10].icell.PDM VPWR.t1997 XA.XIR[15].XIC[10].icell.Ien VGND.t2300 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1463 XA.XIR[12].XIC[14].icell.PUM XA.Cn[14].t26 XA.XIR[12].XIC[14].icell.Ien VPWR.t1659 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1464 XA.XIR[8].XIC[6].icell.PUM XA.Cn[6].t29 XA.XIR[8].XIC[6].icell.Ien VPWR.t430 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1465 VGND.t1134 XThR.XTB7.B a_n1335_8331# VGND.t1133 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1466 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[0].t47 VGND.t763 VGND.t762 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1467 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12].t45 XA.XIR[12].XIC[12].icell.Ien VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1468 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[8].t48 VGND.t148 VGND.t147 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1469 VGND.t1333 XA.Cn[2].t27 XA.XIR[0].XIC[2].icell.PDM VGND.t1332 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1470 XA.XIR[11].XIC[7].icell.PUM XA.Cn[7].t22 XA.XIR[11].XIC[7].icell.Ien VPWR.t503 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1471 VPWR.t22 thermo15c_0.XTBN.Y.t63 XA.Cn[9].t1 VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1472 XA.XIR[15].XIC_15.icell.PUM VPWR.t738 XA.XIR[15].XIC_15.icell.Ien VPWR.t739 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1473 XA.XIR[7].XIC[2].icell.SM XA.XIR[7].XIC[2].icell.Ien Iout.t26 VGND.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1474 a_10051_9569# thermo15c_0.XTBN.Y.t64 VGND.t65 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1475 VGND.t865 XA.Cn[9].t28 XA.XIR[8].XIC[9].icell.PDM VGND.t864 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1476 XA.XIR[10].XIC[3].icell.SM XA.XIR[10].XIC[3].icell.Ien Iout.t132 VGND.t1057 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1477 VPWR.t1807 XThR.XTBN.Y XThR.Tn[7].t1 VPWR.t1806 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1478 VPWR.t52 XThR.Tn[12].t46 XA.XIR[13].XIC[11].icell.PUM VPWR.t51 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1479 XA.XIR[7].XIC[4].icell.PUM XA.Cn[4].t29 XA.XIR[7].XIC[4].icell.Ien VPWR.t1909 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1480 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t736 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t737 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1481 XA.XIR[13].XIC[4].icell.SM XA.XIR[13].XIC[4].icell.Ien Iout.t226 VGND.t1944 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1482 VPWR.t357 XThR.Tn[9].t40 XA.XIR[10].XIC[7].icell.PUM VPWR.t356 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1483 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[2].t39 XA.XIR[2].XIC[8].icell.Ien VGND.t566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1484 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[2].t40 XA.XIR[2].XIC[14].icell.Ien VGND.t1574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1485 XA.Cn[11].t8 thermo15c_0.XTB4.Y.t8 VPWR.t1889 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1486 VGND.t2415 XThR.XTBN.Y XThR.Tn[1].t10 VGND.t2371 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1487 XThR.Tn[1].t5 XThR.XTBN.Y a_n1049_7787# VPWR.t1787 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1488 a_7651_9569# thermo15c_0.XTBN.Y.t65 VGND.t67 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1489 XA.XIR[5].XIC[5].icell.PUM XA.Cn[5].t26 XA.XIR[5].XIC[5].icell.Ien VPWR.t1681 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1490 VGND.t1585 Vbias.t135 XA.XIR[11].XIC[5].icell.SM VGND.t1584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1491 XA.XIR[10].XIC[6].icell.Ien XThR.Tn[10].t43 VPWR.t1756 VPWR.t1755 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1492 XA.XIR[9].XIC[5].icell.PUM XA.Cn[5].t27 XA.XIR[9].XIC[5].icell.Ien VPWR.t1682 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1493 XA.XIR[13].XIC[7].icell.Ien XThR.Tn[13].t38 VPWR.t492 VPWR.t491 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1494 VGND.t1587 Vbias.t136 XA.XIR[5].XIC[9].icell.SM VGND.t1586 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1495 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t1998 VGND.t2302 VGND.t2301 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1496 VPWR.t54 XThR.Tn[12].t47 XA.XIR[13].XIC[2].icell.PUM VPWR.t53 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1497 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout VGND.t2476 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1498 VPWR.t255 XThR.Tn[7].t38 XA.XIR[8].XIC[14].icell.PUM VPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1499 XA.XIR[0].XIC_15.icell.PDM XThR.Tn[0].t48 XA.XIR[0].XIC_15.icell.Ien VGND.t764 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1500 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10].t44 XA.XIR[10].XIC[9].icell.Ien VGND.t331 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1501 XThR.Tn[6].t1 XThR.XTB7.Y VGND.t885 VGND.t884 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1502 a_n1049_5611# XThR.XTB6.Y VPWR.t548 VPWR.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1503 XThR.Tn[9].t4 XThR.XTB2.Y VPWR.t1665 VPWR.t1506 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1504 VPWR.t735 VPWR.t733 XA.XIR[11].XIC_15.icell.PUM VPWR.t734 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1505 VGND.t1589 Vbias.t137 XA.XIR[0].XIC[7].icell.SM VGND.t1588 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1506 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12].t48 XA.XIR[12].XIC[10].icell.Ien VGND.t118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1507 XA.Cn[4].t8 thermo15c_0.XTBN.Y.t66 VGND.t69 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1508 VGND.t518 XA.Cn[6].t30 XA.XIR[0].XIC[6].icell.PDM VGND.t517 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1509 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[5].t44 VGND.t1230 VGND.t1229 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1510 XA.XIR[15].XIC[0].icell.PDM XThR.Tn[14].t43 VGND.t476 VGND.t475 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1511 XA.XIR[11].XIC[11].icell.PUM XA.Cn[11].t28 XA.XIR[11].XIC[11].icell.Ien VPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1512 VPWR.t1805 XThR.XTBN.Y XThR.Tn[13].t9 VPWR.t1783 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1513 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[9].t41 VGND.t434 VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1514 XA.XIR[2].XIC[9].icell.Ien XThR.Tn[2].t41 VPWR.t1162 VPWR.t1161 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1515 VGND.t1700 VGND.t1698 XA.XIR[7].XIC_dummy_right.icell.SM VGND.t1699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1516 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[12].t49 VGND.t120 VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1517 XA.XIR[12].XIC[11].icell.SM XA.XIR[12].XIC[11].icell.Ien Iout.t209 VGND.t1611 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1518 VPWR.t558 XThR.Tn[0].t49 XA.XIR[1].XIC[5].icell.PUM VPWR.t557 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1519 VGND.t2304 VPWR.t1999 XA.XIR[13].XIC_dummy_left.icell.PDM VGND.t2303 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1520 VPWR.t1555 XThR.Tn[4].t47 XA.XIR[5].XIC[5].icell.PUM VPWR.t1554 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1521 VPWR.t359 XThR.Tn[9].t42 XA.XIR[10].XIC[11].icell.PUM VPWR.t358 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1522 XA.XIR[8].XIC[1].icell.PUM XA.Cn[1].t30 XA.XIR[8].XIC[1].icell.Ien VPWR.t1874 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1523 XA.XIR[4].XIC[4].icell.PUM XA.Cn[4].t30 XA.XIR[4].XIC[4].icell.Ien VPWR.t1910 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1524 VGND.t1419 XThR.XTB1.Y XThR.Tn[0].t1 VGND.t1418 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1525 XA.XIR[0].XIC[5].icell.SM XA.XIR[0].XIC[5].icell.Ien Iout.t211 VGND.t1773 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1526 XThR.Tn[5].t9 XThR.XTBN.Y VGND.t2414 VGND.t2400 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1527 XA.XIR[7].XIC[0].icell.PUM XA.Cn[0].t26 XA.XIR[7].XIC[0].icell.Ien VPWR.t1251 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1528 XA.XIR[0].XIC[8].icell.PDM VGND.t1695 VGND.t1697 VGND.t1696 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1529 XA.XIR[0].XIC[14].icell.PDM VGND.t1692 VGND.t1694 VGND.t1693 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1530 VGND.t1132 XThR.XTB7.B XThR.XTB6.Y VGND.t1130 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 XA.XIR[11].XIC[2].icell.PUM XA.Cn[2].t28 XA.XIR[11].XIC[2].icell.Ien VPWR.t1320 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1532 XA.XIR[6].XIC[14].icell.PUM XA.Cn[14].t27 XA.XIR[6].XIC[14].icell.Ien VPWR.t1660 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1533 VGND.t71 thermo15c_0.XTBN.Y.t67 XA.Cn[0].t8 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1534 VGND.t1591 Vbias.t138 XA.XIR[8].XIC[5].icell.SM VGND.t1590 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1535 XA.XIR[7].XIC[6].icell.Ien XThR.Tn[7].t39 VPWR.t257 VPWR.t256 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1536 XA.XIR[13].XIC[11].icell.Ien XThR.Tn[13].t39 VPWR.t973 VPWR.t972 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1537 VGND.t1593 Vbias.t139 XA.XIR[12].XIC[13].icell.SM VGND.t1592 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1538 VGND.t2621 XA.Cn[4].t31 XA.XIR[8].XIC[4].icell.PDM VGND.t2620 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1539 VGND.t2306 VPWR.t2000 XA.XIR[3].XIC_dummy_right.icell.PDM VGND.t2305 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1540 VGND.t128 XA.Cn[12].t29 XA.XIR[12].XIC[12].icell.PDM VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1541 VGND.t73 thermo15c_0.XTBN.Y.t68 XA.Cn[3].t11 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1542 VGND.t1595 Vbias.t140 XA.XIR[15].XIC[14].icell.SM VGND.t1594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1543 VGND.t2027 XA.Cn[5].t28 XA.XIR[11].XIC[5].icell.PDM VGND.t2026 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1544 VGND.t91 XA.Cn[13].t29 XA.XIR[15].XIC[13].icell.PDM VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1545 VPWR.t361 XThR.Tn[9].t43 XA.XIR[10].XIC[2].icell.PUM VPWR.t360 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1546 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[2].t42 XA.XIR[2].XIC[3].icell.Ien VGND.t1573 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1547 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t2001 XA.XIR[15].XIC_dummy_left.icell.Ien VGND.t2307 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1548 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7].t40 XA.XIR[7].XIC[9].icell.Ien VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1549 XA.Cn[7].t5 thermo15c_0.XTBN.Y.t69 VGND.t75 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1550 VPWR.t24 thermo15c_0.XTBN.Y.t70 XA.Cn[12].t9 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1551 VGND.t1597 Vbias.t141 XA.XIR[11].XIC[0].icell.SM VGND.t1596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1552 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10].t45 VPWR.t199 VPWR.t198 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1553 XA.XIR[6].XIC[4].icell.Ien XThR.Tn[6].t44 VPWR.t1864 VPWR.t1863 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1554 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t730 VPWR.t732 VPWR.t731 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1555 VGND.t1599 Vbias.t142 XA.XIR[2].XIC_15.icell.SM VGND.t1598 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1556 VGND.t2050 Vbias.t143 XA.XIR[6].XIC[12].icell.SM VGND.t2049 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1557 VGND.t1112 XA.Cn[8].t27 XA.XIR[2].XIC[8].icell.PDM VGND.t1111 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1558 VGND.t1995 XA.Cn[14].t28 XA.XIR[2].XIC[14].icell.PDM VGND.t1994 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1559 VPWR.t1664 XThR.XTB2.Y a_n1049_7787# VPWR.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1560 XA.XIR[13].XIC[2].icell.Ien XThR.Tn[13].t40 VPWR.t975 VPWR.t974 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1561 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[9].t44 VGND.t436 VGND.t435 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1562 VGND.t2052 Vbias.t144 XA.XIR[5].XIC[4].icell.SM VGND.t2051 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1563 VGND.t2054 Vbias.t145 XA.XIR[9].XIC[13].icell.SM VGND.t2053 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1564 XA.XIR[9].XIC[8].icell.SM XA.XIR[9].XIC[8].icell.Ien Iout.t157 VGND.t1158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1565 XA.XIR[8].XIC[14].icell.Ien XThR.Tn[8].t49 VPWR.t76 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1566 VGND.t77 thermo15c_0.XTBN.Y.t71 a_10915_9569# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1567 VPWR.t1466 VGND.t2695 XA.XIR[0].XIC[4].icell.PUM VPWR.t1465 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1568 VPWR.t1063 XThR.Tn[3].t47 XA.XIR[4].XIC[12].icell.PUM VPWR.t1062 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1569 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10].t46 XA.XIR[10].XIC[4].icell.Ien VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1570 VPWR.t1160 XThR.Tn[2].t43 XA.XIR[3].XIC[13].icell.PUM VPWR.t1159 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1571 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t2002 XA.XIR[5].XIC_dummy_right.icell.Ien VGND.t2308 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1572 XA.XIR[12].XIC[9].icell.SM XA.XIR[12].XIC[9].icell.Ien Iout.t119 VGND.t901 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1573 XA.XIR[11].XIC_15.icell.Ien XThR.Tn[11].t48 VPWR.t498 VPWR.t497 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1574 XA.Cn[11].t9 thermo15c_0.XTB4.Y.t9 a_8963_9569# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1575 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13].t41 XA.XIR[13].XIC[5].icell.Ien VGND.t812 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1576 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t2003 XA.XIR[9].XIC_dummy_right.icell.Ien VGND.t2309 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1577 VPWR.t1866 XThR.Tn[6].t45 XA.XIR[7].XIC[13].icell.PUM VPWR.t1865 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1578 VGND.t2605 thermo15c_0.XTB4.Y.t10 XA.Cn[3].t1 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1579 VGND.t2056 Vbias.t146 XA.XIR[0].XIC[2].icell.SM VGND.t2055 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1580 XThR.Tn[14].t11 XThR.XTBN.Y VPWR.t1804 VPWR.t1785 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1581 XA.XIR[4].XIC[0].icell.PUM XA.Cn[0].t27 XA.XIR[4].XIC[0].icell.Ien VPWR.t1252 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1582 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t728 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t729 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1583 a_7875_9569# thermo15c_0.XTBN.Y.t72 VGND.t79 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1584 VPWR.t546 XThR.XTB6.Y XThR.Tn[13].t3 VPWR.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1585 VGND.t1352 XA.Cn[10].t30 XA.XIR[12].XIC[10].icell.PDM VGND.t1351 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1586 XA.XIR[2].XIC[9].icell.PUM XA.Cn[9].t29 XA.XIR[2].XIC[9].icell.Ien VPWR.t1006 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1587 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[2].t44 XA.XIR[2].XIC[7].icell.Ien VGND.t567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1588 XA.XIR[0].XIC[0].icell.SM XA.XIR[0].XIC[0].icell.Ien Iout.t182 VGND.t1401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1589 XA.XIR[0].XIC[3].icell.PDM VGND.t1689 VGND.t1691 VGND.t1690 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1590 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t2004 XA.XIR[12].XIC_dummy_left.icell.Ien VGND.t2310 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1591 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14].t44 XA.XIR[14].XIC[11].icell.Ien VGND.t477 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1592 XA.Cn[11].t10 thermo15c_0.XTB4.Y.t11 a_8963_9569# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1593 VGND.t2058 Vbias.t147 XA.XIR[8].XIC[0].icell.SM VGND.t2057 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1594 XA.XIR[7].XIC[1].icell.Ien XThR.Tn[7].t41 VPWR.t955 VPWR.t954 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1595 VGND.t2060 Vbias.t148 XA.XIR[3].XIC[12].icell.SM VGND.t2059 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1596 XA.XIR[6].XIC[0].icell.Ien XThR.Tn[6].t46 VPWR.t1868 VPWR.t1867 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1597 VGND.t1688 VGND.t1686 XA.XIR[7].XIC_dummy_left.icell.SM VGND.t1687 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1598 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t726 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t727 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1599 XA.Cn[0].t0 thermo15c_0.XTB1.Y.t12 VGND.t235 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1600 XA.XIR[15].XIC[5].icell.SM XA.XIR[15].XIC[5].icell.Ien Iout.t42 VGND.t177 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1601 VGND.t1074 thermo15c_0.XTBN.Y.t73 a_10051_9569# VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1602 VGND.t1210 XA.Cn[0].t28 XA.XIR[11].XIC[0].icell.PDM VGND.t1209 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1603 VPWR.t1065 XThR.Tn[3].t48 XA.XIR[4].XIC[10].icell.PUM VPWR.t1064 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1604 VGND.t130 XA.Cn[12].t30 XA.XIR[6].XIC[12].icell.PDM VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1605 XThR.XTB1.Y XThR.XTB5.A VPWR.t13 VPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1606 VPWR.t1464 VGND.t2696 XA.XIR[0].XIC[0].icell.PUM VPWR.t1463 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1607 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7].t42 XA.XIR[7].XIC[4].icell.Ien VGND.t779 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1608 XThR.Tn[13].t4 XThR.XTB6.Y a_n997_1579# VGND.t749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1609 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14].t45 XA.XIR[14].XIC[2].icell.Ien VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1610 XA.XIR[10].XIC[7].icell.PUM XA.Cn[7].t23 XA.XIR[10].XIC[7].icell.Ien VPWR.t504 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1611 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2005 VGND.t2312 VGND.t2311 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1612 VGND.t2140 XA.Cn[3].t28 XA.XIR[2].XIC[3].icell.PDM VGND.t2139 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1613 XA.XIR[13].XIC[8].icell.PUM XA.Cn[8].t28 XA.XIR[13].XIC[8].icell.Ien VPWR.t1198 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1614 VGND.t1075 thermo15c_0.XTBN.Y.t74 a_7651_9569# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1615 XA.XIR[4].XIC[12].icell.Ien XThR.Tn[4].t48 VPWR.t1557 VPWR.t1556 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1616 XA.XIR[9].XIC[3].icell.SM XA.XIR[9].XIC[3].icell.Ien Iout.t202 VGND.t1505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1617 thermo15c_0.XTBN.Y.t2 thermo15c_0.XTBN.A VGND.t820 VGND.t819 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1618 XA.XIR[3].XIC[13].icell.Ien XThR.Tn[3].t49 VPWR.t1067 VPWR.t1066 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1619 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t723 VPWR.t725 VPWR.t724 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1620 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[1].t44 XA.XIR[1].XIC[14].icell.Ien VGND.t696 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1621 XA.XIR[12].XIC[4].icell.SM XA.XIR[12].XIC[4].icell.Ien Iout.t32 VGND.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1622 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[1].t45 XA.XIR[1].XIC[8].icell.Ien VGND.t697 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1623 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout VGND.t1159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1624 a_n1335_7243# XThR.XTB7.A XThR.XTB3.Y.t1 VGND.t1453 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1625 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13].t42 XA.XIR[13].XIC[0].icell.Ien VGND.t813 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1626 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8].t50 XA.XIR[8].XIC[12].icell.Ien VGND.t765 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1627 XA.XIR[0].XIC[7].icell.PDM VGND.t1683 VGND.t1685 VGND.t1684 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1628 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t6 VPWR.t1801 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1629 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11].t49 XA.XIR[11].XIC[13].icell.Ien VGND.t1405 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1630 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2006 VGND.t2314 VGND.t2313 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1631 a_4067_9615# thermo15c_0.XTB3.Y.t10 VPWR.t1434 VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1632 VPWR.t1116 thermo15c_0.XTBN.Y.t75 XA.Cn[7].t0 VPWR.t1115 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1633 VPWR.t1158 XThR.Tn[2].t45 XA.XIR[3].XIC[6].icell.PUM VPWR.t1157 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1634 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[11].t50 VGND.t1407 VGND.t1406 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1635 XA.XIR[15].XIC[8].icell.Ien VPWR.t720 VPWR.t722 VPWR.t721 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1636 VPWR.t1870 XThR.Tn[6].t47 XA.XIR[7].XIC[6].icell.PUM VPWR.t1869 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1637 VGND.t2413 XThR.XTBN.Y a_n997_1803# VGND.t2412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1638 VPWR.t1272 XThR.Tn[5].t45 XA.XIR[6].XIC[7].icell.PUM VPWR.t1271 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1639 XThR.Tn[3].t9 XThR.XTBN.Y VGND.t2411 VGND.t2365 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1640 VGND.t1354 XA.Cn[10].t31 XA.XIR[6].XIC[10].icell.PDM VGND.t1353 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1641 VPWR.t560 XThR.Tn[8].t51 XA.XIR[9].XIC[8].icell.PUM VPWR.t559 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1642 VPWR.t1890 thermo15c_0.XTB4.Y.t12 XA.Cn[11].t11 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14].t46 XA.XIR[14].XIC[6].icell.Ien VGND.t479 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1644 XA.XIR[10].XIC[11].icell.PUM XA.Cn[11].t29 XA.XIR[10].XIC[11].icell.Ien VPWR.t329 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1645 VGND.t2062 Vbias.t149 XA.XIR[2].XIC[8].icell.SM VGND.t2061 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1646 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[12].t50 VGND.t122 VGND.t121 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1647 XA.XIR[1].XIC[9].icell.Ien XThR.Tn[1].t46 VPWR.t513 VPWR.t512 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1648 VGND.t690 XA.Cn[7].t24 XA.XIR[2].XIC[7].icell.PDM VGND.t689 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1649 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[11].t51 VGND.t1409 VGND.t1408 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1650 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[7].t43 VGND.t781 VGND.t780 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1651 XA.XIR[4].XIC[10].icell.Ien XThR.Tn[4].t49 VPWR.t1559 VPWR.t1558 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1652 XA.XIR[15].XIC[0].icell.SM XA.XIR[15].XIC[0].icell.Ien Iout.t223 VGND.t1937 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1653 VGND.t2316 VPWR.t2007 XA.XIR[12].XIC_dummy_left.icell.PDM VGND.t2315 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1654 XA.Cn[0].t7 thermo15c_0.XTBN.Y.t76 VGND.t1076 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1655 XA.XIR[10].XIC[12].icell.SM XA.XIR[10].XIC[12].icell.Ien Iout.t94 VGND.t742 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1656 VPWR.t1069 XThR.Tn[3].t50 XA.XIR[4].XIC[5].icell.PUM VPWR.t1068 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1657 XA.XIR[13].XIC[13].icell.SM XA.XIR[13].XIC[13].icell.Ien Iout.t253 VGND.t2629 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1658 XA.Cn[3].t10 thermo15c_0.XTBN.Y.t77 VGND.t1077 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1659 VGND.t1114 XA.Cn[8].t29 XA.XIR[14].XIC[8].icell.PDM VGND.t1113 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1660 VGND.t1997 XA.Cn[14].t29 XA.XIR[14].XIC[14].icell.PDM VGND.t1996 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1661 XA.XIR[10].XIC[2].icell.PUM XA.Cn[2].t29 XA.XIR[10].XIC[2].icell.Ien VPWR.t1321 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1662 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8].t52 XA.XIR[8].XIC[10].icell.Ien VGND.t766 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1663 XA.XIR[5].XIC[14].icell.PUM XA.Cn[14].t30 XA.XIR[5].XIC[14].icell.Ien VPWR.t1623 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1664 XA.XIR[13].XIC[3].icell.PUM XA.Cn[3].t29 XA.XIR[13].XIC[3].icell.Ien VPWR.t1722 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1665 XA.XIR[9].XIC[14].icell.PUM XA.Cn[14].t31 XA.XIR[9].XIC[14].icell.Ien VPWR.t1624 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1666 XA.XIR[8].XIC_15.icell.PUM VPWR.t718 XA.XIR[8].XIC_15.icell.Ien VPWR.t719 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1667 a_n1049_8581# XThR.XTB1.Y VPWR.t1368 VPWR.t1367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1668 VGND.t2547 XA.Cn[1].t31 XA.XIR[15].XIC[1].icell.PDM VGND.t2546 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1669 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[8].t53 VGND.t768 VGND.t767 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1670 VPWR.t717 VPWR.t715 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t716 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1671 VGND.t2064 Vbias.t150 XA.XIR[10].XIC[6].icell.SM VGND.t2063 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1672 VGND.t2029 XA.Cn[5].t29 XA.XIR[10].XIC[5].icell.PDM VGND.t2028 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1673 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[1].t47 XA.XIR[1].XIC[3].icell.Ien VGND.t698 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1674 XA.XIR[12].XIC[8].icell.Ien XThR.Tn[12].t51 VPWR.t56 VPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1675 VPWR.t1274 XThR.Tn[5].t46 XA.XIR[6].XIC[11].icell.PUM VPWR.t1273 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1676 XA.XIR[0].XIC[4].icell.PUM XA.Cn[4].t32 XA.XIR[0].XIC[4].icell.Ien VPWR.t1911 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1677 VGND.t2066 Vbias.t151 XA.XIR[1].XIC_15.icell.SM VGND.t2065 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1678 XA.XIR[7].XIC[13].icell.PUM XA.Cn[13].t30 XA.XIR[7].XIC[13].icell.Ien VPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1679 thermo15c_0.XTB1.Y.t1 thermo15c_0.XTB5.A a_3299_10575# VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1680 XA.XIR[3].XIC[6].icell.Ien XThR.Tn[3].t51 VPWR.t1071 VPWR.t1070 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1681 VPWR.t1156 XThR.Tn[2].t46 XA.XIR[3].XIC[1].icell.PUM VPWR.t1155 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1682 VGND.t39 XThR.XTB3.Y.t10 XThR.Tn[2].t0 VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1683 XA.XIR[15].XIC[3].icell.Ien VPWR.t712 VPWR.t714 VPWR.t713 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1684 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[11].t52 VGND.t1411 VGND.t1410 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1685 VGND.t2068 Vbias.t152 XA.XIR[11].XIC[14].icell.SM VGND.t2067 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1686 XA.XIR[10].XIC_15.icell.Ien XThR.Tn[10].t47 VPWR.t201 VPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1687 XA.XIR[14].XIC[9].icell.PUM XA.Cn[9].t30 XA.XIR[14].XIC[9].icell.Ien VPWR.t1007 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1688 VPWR.t1872 XThR.Tn[6].t48 XA.XIR[7].XIC[1].icell.PUM VPWR.t1871 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1689 VPWR.t1276 XThR.Tn[5].t47 XA.XIR[6].XIC[2].icell.PUM VPWR.t1275 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1690 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout VGND.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1691 VPWR.t1102 XThR.Tn[0].t50 XA.XIR[1].XIC[14].icell.PUM VPWR.t1101 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1692 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[3].t52 XA.XIR[3].XIC[9].icell.Ien VGND.t916 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1693 VPWR.t1561 XThR.Tn[4].t50 XA.XIR[5].XIC[14].icell.PUM VPWR.t1560 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1694 VPWR.t562 XThR.Tn[8].t54 XA.XIR[9].XIC[3].icell.PUM VPWR.t561 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1695 VGND.t1079 thermo15c_0.XTBN.Y.t78 XA.Cn[6].t6 VGND.t1078 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1696 VGND.t2070 Vbias.t153 XA.XIR[2].XIC[3].icell.SM VGND.t2069 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1697 XA.XIR[6].XIC[7].icell.SM XA.XIR[6].XIC[7].icell.Ien Iout.t141 VGND.t1105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1698 XA.Cn[10].t8 thermo15c_0.XTB3.Y.t11 VPWR.t1435 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1699 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[7].t44 VGND.t783 VGND.t782 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1700 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[2].t47 VGND.t571 VGND.t570 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1701 XA.XIR[4].XIC[5].icell.Ien XThR.Tn[4].t51 VPWR.t1563 VPWR.t1562 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1702 VGND.t1682 VGND.t1680 XA.XIR[0].XIC_dummy_right.icell.SM VGND.t1681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1703 VGND.t2072 Vbias.t154 XA.XIR[14].XIC[7].icell.SM VGND.t2071 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1704 VGND.t1473 Vbias.t155 XA.XIR[10].XIC[10].icell.SM VGND.t1472 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1705 XA.Cn[14].t6 thermo15c_0.XTB7.Y VPWR.t1349 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1706 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[5].t48 VGND.t1232 VGND.t1231 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1707 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[1].t48 XA.XIR[1].XIC[7].icell.Ien VGND.t1952 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1708 VGND.t2318 VPWR.t2008 XA.XIR[6].XIC_dummy_left.icell.PDM VGND.t2317 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1709 VGND.t236 thermo15c_0.XTB1.Y.t13 XA.Cn[0].t1 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1710 VGND.t2142 XA.Cn[3].t30 XA.XIR[14].XIC[3].icell.PDM VGND.t2141 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1711 XA.XIR[0].XIC[0].icell.PUM XA.Cn[0].t29 XA.XIR[0].XIC[0].icell.Ien VPWR.t1253 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1712 XA.XIR[1].XIC[12].icell.PUM XA.Cn[12].t31 XA.XIR[1].XIC[12].icell.Ien VPWR.t62 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1713 XA.XIR[4].XIC[13].icell.PUM XA.Cn[13].t31 XA.XIR[4].XIC[13].icell.Ien VPWR.t29 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1714 VGND.t1475 Vbias.t156 XA.XIR[10].XIC[1].icell.SM VGND.t1474 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1715 XThR.Tn[8].t9 XThR.XTBN.Y VPWR.t1803 VPWR.t1802 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1716 XA.XIR[0].XIC[14].icell.SM XA.XIR[0].XIC[14].icell.Ien Iout.t199 VGND.t1502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1717 VGND.t1477 Vbias.t157 XA.XIR[5].XIC[13].icell.SM VGND.t1476 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1718 XA.XIR[14].XIC[5].icell.SM XA.XIR[14].XIC[5].icell.Ien Iout.t179 VGND.t1378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1719 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[13].t43 VGND.t815 VGND.t814 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1720 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[13].t44 VGND.t817 VGND.t816 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1721 VGND.t1212 XA.Cn[0].t30 XA.XIR[10].XIC[0].icell.PDM VGND.t1211 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1722 VGND.t132 XA.Cn[12].t32 XA.XIR[5].XIC[12].icell.PDM VGND.t131 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1723 XA.XIR[12].XIC[3].icell.Ien XThR.Tn[12].t52 VPWR.t281 VPWR.t280 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1724 VGND.t134 XA.Cn[12].t33 XA.XIR[9].XIC[12].icell.PDM VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1725 VGND.t1479 Vbias.t158 XA.XIR[8].XIC[14].icell.SM VGND.t1478 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1726 XA.XIR[7].XIC_15.icell.Ien XThR.Tn[7].t45 VPWR.t957 VPWR.t956 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1727 VGND.t93 XA.Cn[13].t32 XA.XIR[8].XIC[13].icell.PDM VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1728 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t2009 XA.XIR[8].XIC_dummy_left.icell.Ien VGND.t2319 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1729 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t5 VPWR.t1801 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1730 XA.XIR[3].XIC[1].icell.Ien XThR.Tn[3].t53 VPWR.t1073 VPWR.t1072 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1731 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[4].t52 VGND.t1824 VGND.t1823 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1732 XA.XIR[12].XIC[8].icell.PUM XA.Cn[8].t30 XA.XIR[12].XIC[8].icell.Ien VPWR.t1199 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1733 VGND.t1481 Vbias.t159 XA.XIR[4].XIC[11].icell.SM VGND.t1480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1734 XA.XIR[3].XIC[7].icell.SM XA.XIR[3].XIC[7].icell.Ien Iout.t248 VGND.t2530 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1735 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[2].t48 VGND.t569 VGND.t568 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1736 XThR.XTBN.A data[7].t1 VGND.t2005 VGND.t2004 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1737 XA.XIR[6].XIC[13].icell.Ien XThR.Tn[6].t49 VPWR.t1686 VPWR.t1685 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1738 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[3].t54 XA.XIR[3].XIC[4].icell.Ien VGND.t917 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1739 XA.Cn[14].t5 thermo15c_0.XTB7.Y VPWR.t1348 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1740 VPWR.t528 XThR.Tn[13].t45 XA.XIR[14].XIC[4].icell.PUM VPWR.t527 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1741 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11].t53 XA.XIR[11].XIC[1].icell.Ien VGND.t1412 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1742 XA.XIR[7].XIC[6].icell.PUM XA.Cn[6].t31 XA.XIR[7].XIC[6].icell.Ien VPWR.t431 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1743 VPWR.t1462 VGND.t2697 XA.XIR[0].XIC[13].icell.PUM VPWR.t1461 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1744 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2010 XA.XIR[2].XIC_dummy_right.icell.Ien VGND.t2320 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1745 VGND.t692 XA.Cn[7].t25 XA.XIR[14].XIC[7].icell.PDM VGND.t691 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1746 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10].t48 XA.XIR[10].XIC[13].icell.Ien VGND.t333 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1747 thermo15c_0.XTB2.Y thermo15c_0.XTB7.B VPWR.t1128 VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1748 XA.XIR[1].XIC[10].icell.PUM XA.Cn[10].t32 XA.XIR[1].XIC[10].icell.Ien VPWR.t1335 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1749 XA.XIR[6].XIC[2].icell.SM XA.XIR[6].XIC[2].icell.Ien Iout.t183 VGND.t1402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1750 XA.XIR[0].XIC[12].icell.Ien XThR.Tn[0].t51 VPWR.t1104 VPWR.t1103 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1751 XThR.Tn[5].t8 XThR.XTBN.Y VGND.t2410 VGND.t2389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1752 VGND.t867 XA.Cn[9].t31 XA.XIR[7].XIC[9].icell.PDM VGND.t866 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1753 XA.XIR[15].XIC[11].icell.PDM XThR.Tn[14].t47 VGND.t481 VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1754 VGND.t1483 Vbias.t160 XA.XIR[14].XIC[2].icell.SM VGND.t1482 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1755 VGND.t1356 XA.Cn[10].t33 XA.XIR[5].XIC[10].icell.PDM VGND.t1355 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1756 XThR.Tn[10].t9 XThR.XTBN.Y VPWR.t1800 VPWR.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1757 VPWR.t959 XThR.Tn[7].t46 XA.XIR[8].XIC[8].icell.PUM VPWR.t958 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1758 VGND.t1358 XA.Cn[10].t34 XA.XIR[9].XIC[10].icell.PDM VGND.t1357 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1759 a_5949_9615# thermo15c_0.XTB6.Y VPWR.t1034 VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1760 VGND.t1485 Vbias.t161 XA.XIR[1].XIC[8].icell.SM VGND.t1484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1761 VGND.t1487 Vbias.t162 XA.XIR[4].XIC[9].icell.SM VGND.t1486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1762 XA.XIR[14].XIC[0].icell.SM XA.XIR[14].XIC[0].icell.Ien Iout.t124 VGND.t1031 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1763 XA.XIR[15].XIC[2].icell.PDM XThR.Tn[14].t48 VGND.t483 VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1764 VPWR.t1193 thermo15c_0.XTB3.Y.t12 XA.Cn[10].t2 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1765 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[13].t46 VGND.t726 VGND.t725 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1766 VGND.t1679 VGND.t1677 XA.XIR[0].XIC_dummy_left.icell.SM VGND.t1678 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1767 XA.XIR[5].XIC_15.icell.SM XA.XIR[5].XIC_15.icell.Ien Iout.t187 VGND.t1426 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1768 XA.XIR[9].XIC[12].icell.SM XA.XIR[9].XIC[12].icell.Ien Iout.t153 VGND.t1154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1769 XA.Cn[13].t8 thermo15c_0.XTBN.Y.t79 VPWR.t1117 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1770 XA.XIR[13].XIC_15.icell.PDM VPWR.t2011 VGND.t2322 VGND.t2321 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1771 a_n997_3755# XThR.XTBN.Y VGND.t2409 VGND.t2395 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1772 XA.XIR[12].XIC[13].icell.SM XA.XIR[12].XIC[13].icell.Ien Iout.t9 VGND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1773 VPWR.t1798 XThR.XTBN.Y XThR.Tn[14].t10 VPWR.t1797 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 XA.XIR[15].XIC[14].icell.SM XA.XIR[15].XIC[14].icell.Ien Iout.t37 VGND.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1775 XA.XIR[4].XIC[6].icell.PUM XA.Cn[6].t32 XA.XIR[4].XIC[6].icell.Ien VPWR.t432 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1776 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[8].t55 VGND.t770 VGND.t769 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1777 XA.XIR[3].XIC[7].icell.PUM XA.Cn[7].t26 XA.XIR[3].XIC[7].icell.Ien VPWR.t505 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1778 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[4].t53 VGND.t1915 VGND.t1914 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1779 XA.XIR[12].XIC[3].icell.PUM XA.Cn[3].t31 XA.XIR[12].XIC[3].icell.Ien VPWR.t1723 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1780 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2012 VGND.t2324 VGND.t2323 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1781 VPWR.t530 XThR.Tn[13].t47 XA.XIR[14].XIC[0].icell.PUM VPWR.t529 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1782 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7].t47 XA.XIR[7].XIC[13].icell.Ien VGND.t784 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1783 XA.XIR[0].XIC[10].icell.Ien XThR.Tn[0].t52 VPWR.t1106 VPWR.t1105 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1784 XA.XIR[3].XIC[2].icell.SM XA.XIR[3].XIC[2].icell.Ien Iout.t73 VGND.t563 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1785 XA.XIR[6].XIC[8].icell.PUM XA.Cn[8].t31 XA.XIR[6].XIC[8].icell.Ien VPWR.t1671 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1786 XA.XIR[11].XIC[11].icell.SM XA.XIR[11].XIC[11].icell.Ien Iout.t177 VGND.t1376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1787 XThR.Tn[7].t4 XThR.XTBN.Y VGND.t2398 VGND.t2397 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1788 XA.XIR[2].XIC_15.icell.SM XA.XIR[2].XIC_15.icell.Ien Iout.t52 VGND.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1789 VPWR.t711 VPWR.t709 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t710 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1790 VGND.t869 XA.Cn[9].t32 XA.XIR[4].XIC[9].icell.PDM VGND.t868 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1791 XA.XIR[14].XIC[4].icell.Ien XThR.Tn[14].t49 VPWR.t400 VPWR.t399 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1792 XA.XIR[7].XIC[1].icell.PUM XA.Cn[1].t32 XA.XIR[7].XIC[1].icell.Ien VPWR.t1875 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1793 VGND.t2326 VPWR.t2013 XA.XIR[15].XIC_15.icell.PDM VGND.t2325 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1794 thermo15c_0.XTB4.Y.t1 thermo15c_0.XTB7.B VGND.t1101 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1795 VPWR.t544 XThR.XTB6.Y XThR.Tn[13].t2 VPWR.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VPWR.t1356 XThR.XTB3.Y.t11 a_n1049_7493# VPWR.t1355 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1797 XA.XIR[1].XIC[5].icell.PUM XA.Cn[5].t30 XA.XIR[1].XIC[5].icell.Ien VPWR.t1683 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1798 VPWR.t1358 XThR.Tn[11].t54 XA.XIR[12].XIC[12].icell.PUM VPWR.t1357 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1799 VGND.t1489 Vbias.t163 XA.XIR[7].XIC[5].icell.SM VGND.t1488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1800 XA.XIR[6].XIC[6].icell.Ien XThR.Tn[6].t50 VPWR.t1688 VPWR.t1687 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1801 XA.XIR[5].XIC[7].icell.Ien XThR.Tn[5].t49 VPWR.t1278 VPWR.t1277 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1802 VPWR.t458 data[4].t3 XThR.XTB7.A VPWR.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1803 VGND.t2623 XA.Cn[4].t33 XA.XIR[7].XIC[4].icell.PDM VGND.t2622 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1804 VGND.t1491 Vbias.t164 XA.XIR[6].XIC[6].icell.SM VGND.t1490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1805 VGND.t2328 VPWR.t2014 XA.XIR[2].XIC_dummy_right.icell.PDM VGND.t2327 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1806 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2015 VGND.t2330 VGND.t2329 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1807 XA.XIR[15].XIC[6].icell.PDM XThR.Tn[14].t50 VGND.t485 VGND.t484 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1808 XA.Cn[6].t5 thermo15c_0.XTBN.Y.t80 VGND.t1081 VGND.t1080 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1809 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[13].t48 VGND.t728 VGND.t727 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1810 XA.XIR[9].XIC[7].icell.Ien XThR.Tn[9].t45 VPWR.t363 VPWR.t362 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1811 XA.XIR[8].XIC[8].icell.Ien XThR.Tn[8].t56 VPWR.t564 VPWR.t563 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1812 VPWR.t1460 VGND.t2698 XA.XIR[0].XIC[6].icell.PUM VPWR.t1459 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1813 VPWR.t1075 XThR.Tn[3].t55 XA.XIR[4].XIC[14].icell.PUM VPWR.t1074 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1814 XThR.Tn[5].t1 XThR.XTB6.Y VGND.t748 VGND.t747 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1815 VPWR.t1385 XThR.Tn[7].t48 XA.XIR[8].XIC[3].icell.PUM VPWR.t1384 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1816 VPWR.t339 thermo15c_0.XTB5.Y a_5155_9615# VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1817 VPWR.t708 VPWR.t706 XA.XIR[3].XIC_15.icell.PUM VPWR.t707 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1818 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6].t51 XA.XIR[6].XIC[9].icell.Ien VGND.t2034 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1819 VPWR.t705 VPWR.t703 XA.XIR[7].XIC_15.icell.PUM VPWR.t704 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1820 VGND.t1493 Vbias.t165 XA.XIR[1].XIC[3].icell.SM VGND.t1492 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1821 XA.XIR[3].XIC[11].icell.PUM XA.Cn[11].t30 XA.XIR[3].XIC[11].icell.Ien VPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1822 XThR.Tn[4].t2 XThR.XTB5.Y VGND.t1167 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1823 a_4861_9615# thermo15c_0.XTB4.Y.t13 VPWR.t155 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1824 a_5949_9615# thermo15c_0.XTBN.Y.t81 XA.Cn[5].t5 VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1825 VGND.t1495 Vbias.t166 XA.XIR[4].XIC[4].icell.SM VGND.t1494 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1826 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[5].t50 VGND.t1234 VGND.t1233 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1827 VGND.t2332 VPWR.t2016 XA.XIR[5].XIC_dummy_left.icell.PDM VGND.t2331 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1828 XA.XIR[11].XIC[9].icell.SM XA.XIR[11].XIC[9].icell.Ien Iout.t53 VGND.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1829 VGND.t1082 thermo15c_0.XTBN.Y.t82 XA.Cn[2].t3 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1830 VGND.t2334 VPWR.t2017 XA.XIR[9].XIC_dummy_left.icell.PDM VGND.t2333 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1831 XA.XIR[8].XIC[11].icell.SM XA.XIR[8].XIC[11].icell.Ien Iout.t121 VGND.t1007 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1832 VPWR.t143 thermo15c_0.XTB1.Y.t14 XA.Cn[8].t1 VPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1833 VGND.t403 XA.Cn[11].t31 XA.XIR[11].XIC[11].icell.PDM VGND.t402 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1834 a_5155_10571# thermo15c_0.XTB7.B thermo15c_0.XTB5.Y VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1835 a_10915_9569# thermo15c_0.XTBN.Y.t83 VGND.t2358 VGND.t2357 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1836 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14].t51 VPWR.t1628 VPWR.t1627 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1837 XA.XIR[4].XIC[1].icell.PUM XA.Cn[1].t33 XA.XIR[4].XIC[1].icell.Ien VPWR.t1876 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1838 XA.XIR[3].XIC[2].icell.PUM XA.Cn[2].t30 XA.XIR[3].XIC[2].icell.Ien VPWR.t1322 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1839 VPWR.t1360 XThR.Tn[11].t55 XA.XIR[12].XIC[10].icell.PUM VPWR.t1359 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1840 XA.XIR[0].XIC[5].icell.Ien XThR.Tn[0].t53 VPWR.t1108 VPWR.t1107 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1841 XA.XIR[6].XIC[3].icell.PUM XA.Cn[3].t32 XA.XIR[6].XIC[3].icell.Ien VPWR.t1724 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1842 VGND.t959 Vbias.t167 XA.XIR[6].XIC[10].icell.SM VGND.t958 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1843 XA.XIR[5].XIC[11].icell.Ien XThR.Tn[5].t51 VPWR.t1280 VPWR.t1279 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1844 XA.Cn[3].t0 thermo15c_0.XTB4.Y.t14 VGND.t295 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1845 VGND.t961 Vbias.t168 XA.XIR[3].XIC[6].icell.SM VGND.t960 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1846 VGND.t2625 XA.Cn[4].t34 XA.XIR[4].XIC[4].icell.PDM VGND.t2624 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1847 VGND.t2549 XA.Cn[1].t34 XA.XIR[8].XIC[1].icell.PDM VGND.t2548 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1848 VGND.t2031 XA.Cn[5].t31 XA.XIR[3].XIC[5].icell.PDM VGND.t2030 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1849 XA.XIR[9].XIC[11].icell.Ien XThR.Tn[9].t46 VPWR.t377 VPWR.t376 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1850 VGND.t1335 XA.Cn[2].t31 XA.XIR[11].XIC[2].icell.PDM VGND.t1334 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1851 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[3].t56 VGND.t919 VGND.t918 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1852 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13].t49 XA.XIR[13].XIC[11].icell.Ien VGND.t729 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1853 XThR.Tn[3].t8 XThR.XTBN.Y VGND.t2408 VGND.t2407 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1854 XA.XIR[0].XIC[13].icell.PUM XA.Cn[13].t33 XA.XIR[0].XIC[13].icell.Ien VPWR.t1921 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1855 XA.XIR[6].XIC[1].icell.Ien XThR.Tn[6].t52 VPWR.t1690 VPWR.t1689 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1856 VGND.t963 Vbias.t169 XA.XIR[7].XIC[0].icell.SM VGND.t962 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1857 VGND.t965 Vbias.t170 XA.XIR[2].XIC[12].icell.SM VGND.t964 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1858 XA.XIR[5].XIC[2].icell.Ien XThR.Tn[5].t52 VPWR.t1282 VPWR.t1281 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1859 VGND.t967 Vbias.t171 XA.XIR[6].XIC[1].icell.SM VGND.t966 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1860 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t701 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t702 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1861 a_10915_9569# thermo15c_0.XTB7.Y XA.Cn[14].t9 VGND.t1396 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1862 XA.XIR[9].XIC[2].icell.Ien XThR.Tn[9].t47 VPWR.t379 VPWR.t378 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1863 a_4387_10575# thermo15c_0.XTB7.B VGND.t1100 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1864 XA.XIR[4].XIC[14].icell.Ien XThR.Tn[4].t54 VPWR.t1576 VPWR.t1575 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1865 XA.XIR[5].XIC[8].icell.SM XA.XIR[5].XIC[8].icell.Ien Iout.t78 VGND.t636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1866 XA.XIR[8].XIC[3].icell.Ien XThR.Tn[8].t57 VPWR.t1220 VPWR.t1219 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1867 VPWR.t1458 VGND.t2699 XA.XIR[0].XIC[1].icell.PUM VPWR.t1457 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1868 XA.XIR[3].XIC_15.icell.Ien XThR.Tn[3].t57 VPWR.t1077 VPWR.t1076 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1869 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10].t49 XA.XIR[10].XIC[1].icell.Ien VGND.t334 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1870 XA.XIR[8].XIC[9].icell.SM XA.XIR[8].XIC[9].icell.Ien Iout.t176 VGND.t1375 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1871 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6].t53 XA.XIR[6].XIC[4].icell.Ien VGND.t2035 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1872 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t2018 XA.XIR[1].XIC_dummy_right.icell.Ien VGND.t2335 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1873 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5].t53 XA.XIR[5].XIC[5].icell.Ien VGND.t1764 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1874 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13].t50 XA.XIR[13].XIC[2].icell.Ien VGND.t730 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1875 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9].t48 XA.XIR[9].XIC[5].icell.Ien VGND.t449 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1876 a_10051_9569# thermo15c_0.XTBN.Y.t84 VGND.t2359 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1877 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11].t56 XA.XIR[11].XIC_15.icell.Ien VGND.t1606 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1878 thermo15c_0.XTB1.Y.t0 thermo15c_0.XTB7.B VPWR.t1127 VPWR.t1126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1879 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t5 VPWR.t1793 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1880 XA.XIR[2].XIC[8].icell.SM XA.XIR[2].XIC[8].icell.Ien Iout.t110 VGND.t828 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1881 XA.XIR[11].XIC[4].icell.SM XA.XIR[11].XIC[4].icell.Ien Iout.t161 VGND.t1169 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1882 VGND.t969 Vbias.t172 XA.XIR[3].XIC[10].icell.SM VGND.t968 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1883 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t698 VPWR.t700 VPWR.t699 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1884 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout VGND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1885 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t5 VPWR.t1796 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1886 a_7651_9569# thermo15c_0.XTBN.Y.t85 VGND.t2360 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1887 VGND.t1676 VGND.t1674 XA.XIR[14].XIC_dummy_right.icell.SM VGND.t1675 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1888 VGND.t520 XA.Cn[6].t33 XA.XIR[11].XIC[6].icell.PDM VGND.t519 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1889 VPWR.t1740 thermo15c_0.XTB7.A a_6243_10571# VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1890 VPWR.t697 VPWR.t695 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t696 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1891 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[0].t54 VGND.t1062 VGND.t1061 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1892 VPWR.t1442 XThR.Tn[11].t57 XA.XIR[12].XIC[5].icell.PUM VPWR.t1441 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1893 XA.Cn[10].t3 thermo15c_0.XTB3.Y.t13 a_8739_9569# VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1894 VGND.t971 Vbias.t173 XA.XIR[3].XIC[1].icell.SM VGND.t970 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1895 XA.XIR[7].XIC[5].icell.SM XA.XIR[7].XIC[5].icell.Ien Iout.t151 VGND.t1152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1896 VGND.t1214 XA.Cn[0].t31 XA.XIR[3].XIC[0].icell.PDM VGND.t1213 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1897 VGND.t2406 XThR.XTBN.Y XThR.Tn[2].t9 VGND.t2405 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1898 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[10].t50 VGND.t336 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1899 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[10].t51 VGND.t338 VGND.t337 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1900 XA.XIR[10].XIC[6].icell.SM XA.XIR[10].XIC[6].icell.Ien Iout.t40 VGND.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1901 XThR.XTB5.A data[5].t3 VGND.t1087 VGND.t1086 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1902 XA.XIR[14].XIC[14].icell.SM XA.XIR[14].XIC[14].icell.Ien Iout.t217 VGND.t1784 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1903 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t693 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t694 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1904 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[3].t58 VGND.t287 VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1905 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7].t49 XA.XIR[7].XIC[1].icell.Ien VGND.t1444 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1906 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13].t51 XA.XIR[13].XIC[6].icell.Ien VGND.t1530 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1907 XThR.Tn[12].t9 XThR.XTBN.Y VPWR.t1795 VPWR.t1794 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1908 VGND.t2337 VPWR.t2019 XA.XIR[14].XIC_dummy_right.icell.PDM VGND.t2336 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1909 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[6].t54 VGND.t2037 VGND.t2036 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1910 XA.XIR[5].XIC[8].icell.PUM XA.Cn[8].t32 XA.XIR[5].XIC[8].icell.Ien VPWR.t1672 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1911 XThR.Tn[12].t1 XThR.XTB5.Y a_n997_1803# VGND.t750 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1912 XA.XIR[1].XIC_15.icell.SM XA.XIR[1].XIC_15.icell.Ien Iout.t115 VGND.t879 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1913 XA.XIR[9].XIC[8].icell.PUM XA.Cn[8].t33 XA.XIR[9].XIC[8].icell.Ien VPWR.t1673 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1914 XThR.Tn[3].t2 XThR.XTB4.Y.t11 VGND.t1260 VGND.t1029 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1915 XA.XIR[5].XIC[3].icell.SM XA.XIR[5].XIC[3].icell.Ien Iout.t159 VGND.t1163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1916 VGND.t2404 XThR.XTBN.Y a_n997_2667# VGND.t2403 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1917 XA.XIR[9].XIC_15.icell.PDM VPWR.t2020 VGND.t2339 VGND.t2338 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1918 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5].t54 XA.XIR[5].XIC[0].icell.Ien VGND.t1765 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1919 XA.XIR[8].XIC[4].icell.SM XA.XIR[8].XIC[4].icell.Ien Iout.t240 VGND.t2158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1920 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout VGND.t1162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1921 VGND.t973 Vbias.t174 XA.XIR[13].XIC_15.icell.SM VGND.t972 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1922 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t690 VPWR.t692 VPWR.t691 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1923 XA.XIR[0].XIC[6].icell.PUM XA.Cn[6].t34 XA.XIR[0].XIC[6].icell.Ien VPWR.t433 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1924 VGND.t1963 XA.Cn[14].t32 XA.XIR[13].XIC[14].icell.PDM VGND.t1962 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1925 VGND.t2007 XA.Cn[8].t34 XA.XIR[13].XIC[8].icell.PDM VGND.t2006 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1926 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9].t49 XA.XIR[9].XIC[0].icell.Ien VGND.t450 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1927 a_5155_9615# thermo15c_0.XTB5.Y VPWR.t338 VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1928 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[4].t55 XA.XIR[4].XIC[12].icell.Ien VGND.t1916 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1929 VPWR.t337 thermo15c_0.XTB5.Y XA.Cn[12].t0 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1930 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[3].t59 XA.XIR[3].XIC[13].icell.Ien VGND.t288 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1931 VPWR.t1630 XThR.Tn[14].t52 XA.XIR[15].XIC[12].icell.PUM VPWR.t1629 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1932 XA.XIR[7].XIC_15.icell.PUM VPWR.t688 XA.XIR[7].XIC_15.icell.Ien VPWR.t689 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1933 VPWR.t1419 XThR.Tn[13].t52 XA.XIR[14].XIC[13].icell.PUM VPWR.t1418 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1934 VPWR.t687 VPWR.t685 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t686 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1935 VGND.t871 XA.Cn[9].t33 XA.XIR[0].XIC[9].icell.PDM VGND.t870 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1936 XA.Cn[5].t4 thermo15c_0.XTBN.Y.t86 a_5949_9615# VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1937 XA.XIR[2].XIC[3].icell.SM XA.XIR[2].XIC[3].icell.Ien Iout.t71 VGND.t561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1938 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[7].t50 VGND.t1446 VGND.t1445 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1939 VGND.t413 thermo15c_0.XTB5.Y XA.Cn[4].t0 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1940 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t9 VPWR.t1793 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1941 VPWR.t1608 XThR.Tn[1].t49 XA.XIR[2].XIC[7].icell.PUM VPWR.t1607 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1942 VPWR.t1110 XThR.Tn[0].t55 XA.XIR[1].XIC[8].icell.PUM VPWR.t1109 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1943 XA.XIR[10].XIC[10].icell.SM XA.XIR[10].XIC[10].icell.Ien Iout.t63 VGND.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1944 XA.Cn[2].t2 thermo15c_0.XTBN.Y.t87 VGND.t2361 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1945 VPWR.t1578 XThR.Tn[4].t56 XA.XIR[5].XIC[8].icell.PUM VPWR.t1577 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1946 XA.XIR[15].XIC[14].icell.PDM VPWR.t2021 XA.XIR[15].XIC[14].icell.Ien VGND.t2340 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1947 XA.XIR[15].XIC[8].icell.PDM VPWR.t2022 XA.XIR[15].XIC[8].icell.Ien VGND.t2341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1948 a_5155_9615# thermo15c_0.XTBN.Y.t88 XA.Cn[4].t5 VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1949 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[0].t56 VGND.t1064 VGND.t1063 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1950 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[7].t51 VGND.t1448 VGND.t1447 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1951 XA.XIR[13].XIC[9].icell.PUM XA.Cn[9].t34 XA.XIR[13].XIC[9].icell.Ien VPWR.t1008 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1952 XA.XIR[7].XIC[0].icell.SM XA.XIR[7].XIC[0].icell.Ien Iout.t238 VGND.t2148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1953 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout VGND.t2630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1954 VPWR.t1213 XThR.XTB7.B XThR.XTB2.Y VPWR.t1210 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1955 XA.Cn[8].t4 thermo15c_0.XTB1.Y.t15 a_7651_9569# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1956 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[10].t52 VGND.t340 VGND.t339 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1957 VGND.t405 XA.Cn[11].t32 XA.XIR[10].XIC[11].icell.PDM VGND.t404 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1958 XA.XIR[10].XIC[1].icell.SM XA.XIR[10].XIC[1].icell.Ien Iout.t86 VGND.t715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1959 XA.XIR[6].XIC_15.icell.PDM VPWR.t2023 VGND.t2343 VGND.t2342 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1960 VGND.t2465 thermo15c_0.XTB5.A thermo15c_0.XTB5.Y VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1961 VGND.t1673 VGND.t1671 XA.XIR[14].XIC_dummy_left.icell.SM VGND.t1672 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1962 VGND.t883 XThR.XTB7.Y XThR.Tn[6].t0 VGND.t882 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1963 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[4].t57 XA.XIR[4].XIC[10].icell.Ien VGND.t1917 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1964 XA.XIR[1].XIC[14].icell.PUM XA.Cn[14].t33 XA.XIR[1].XIC[14].icell.Ien VPWR.t1625 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1965 XA.XIR[5].XIC[3].icell.PUM XA.Cn[3].t33 XA.XIR[5].XIC[3].icell.Ien VPWR.t1725 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1966 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[6].t55 VGND.t2039 VGND.t2038 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1967 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[1].t50 VGND.t1954 VGND.t1953 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1968 VPWR.t1632 XThR.Tn[14].t53 XA.XIR[15].XIC[10].icell.PUM VPWR.t1631 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1969 XA.XIR[9].XIC[3].icell.PUM XA.Cn[3].t34 XA.XIR[9].XIC[3].icell.Ien VPWR.t1726 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1970 XA.XIR[4].XIC_15.icell.PUM VPWR.t683 XA.XIR[4].XIC_15.icell.Ien VPWR.t684 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1971 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[4].t58 VGND.t1919 VGND.t1918 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1972 XA.XIR[4].XIC[11].icell.SM XA.XIR[4].XIC[11].icell.Ien Iout.t109 VGND.t827 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1973 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2024 VGND.t2345 VGND.t2344 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1974 XA.XIR[15].XIC[9].icell.Ien VPWR.t680 VPWR.t682 VPWR.t681 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1975 VGND.t1337 XA.Cn[2].t32 XA.XIR[10].XIC[2].icell.PDM VGND.t1336 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1976 XThR.Tn[9].t8 XThR.XTBN.Y VPWR.t1789 VPWR.t1772 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1977 VGND.t2362 thermo15c_0.XTBN.Y.t89 a_9827_9569# VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1978 XA.XIR[0].XIC[1].icell.PUM XA.Cn[1].t35 XA.XIR[0].XIC[1].icell.Ien VPWR.t1877 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1979 VPWR.t1610 XThR.Tn[1].t51 XA.XIR[2].XIC[11].icell.PUM VPWR.t1609 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1980 VGND.t2144 XA.Cn[3].t35 XA.XIR[13].XIC[3].icell.PDM VGND.t2143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1981 VGND.t2347 VPWR.t2025 XA.XIR[8].XIC_15.icell.PDM VGND.t2346 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1982 VPWR.t1222 XThR.Tn[8].t58 XA.XIR[9].XIC[9].icell.PUM VPWR.t1221 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1983 VGND.t975 Vbias.t175 XA.XIR[1].XIC[12].icell.SM VGND.t974 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1984 XA.XIR[14].XIC[13].icell.Ien XThR.Tn[14].t54 VPWR.t1634 VPWR.t1633 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1985 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t677 VPWR.t679 VPWR.t678 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1986 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12].t53 XA.XIR[12].XIC[14].icell.Ien VGND.t383 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1987 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t675 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t676 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1988 XA.Cn[0].t11 thermo15c_0.XTB1.Y.t16 VGND.t2147 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1989 VGND.t977 Vbias.t176 XA.XIR[0].XIC[5].icell.SM VGND.t976 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1990 VGND.t979 Vbias.t177 XA.XIR[4].XIC[13].icell.SM VGND.t978 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1991 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12].t54 XA.XIR[12].XIC[8].icell.Ien VGND.t384 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1992 VGND.t2627 XA.Cn[4].t35 XA.XIR[0].XIC[4].icell.PDM VGND.t2626 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1993 a_10051_9569# thermo15c_0.XTB6.Y XA.Cn[13].t4 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1994 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[7].t52 VGND.t1450 VGND.t1449 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1995 XA.XIR[2].XIC[7].icell.Ien XThR.Tn[2].t49 VPWR.t1154 VPWR.t1153 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1996 VGND.t981 Vbias.t178 XA.XIR[7].XIC[14].icell.SM VGND.t980 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1997 XA.XIR[6].XIC_15.icell.Ien XThR.Tn[6].t56 VPWR.t1692 VPWR.t1691 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1998 VPWR.t1612 XThR.Tn[1].t52 XA.XIR[2].XIC[2].icell.PUM VPWR.t1611 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1999 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[10].t53 VGND.t638 VGND.t637 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2000 VGND.t2650 XA.Cn[13].t34 XA.XIR[7].XIC[13].icell.PDM VGND.t2649 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2001 VPWR.t86 XThR.Tn[0].t57 XA.XIR[1].XIC[3].icell.PUM VPWR.t85 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2002 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout VGND.t1085 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2003 XThR.Tn[14].t9 XThR.XTBN.Y VPWR.t1792 VPWR.t1791 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2004 VPWR.t1580 XThR.Tn[4].t59 XA.XIR[5].XIC[3].icell.PUM VPWR.t1579 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2005 VPWR.t674 VPWR.t672 XA.XIR[0].XIC_15.icell.PUM VPWR.t673 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2006 VPWR.t1421 XThR.Tn[13].t53 XA.XIR[14].XIC[6].icell.PUM VPWR.t1420 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2007 XA.XIR[15].XIC[3].icell.PDM VPWR.t2026 XA.XIR[15].XIC[3].icell.Ien VGND.t2348 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2008 a_n997_3755# XThR.XTBN.Y VGND.t2402 VGND.t2387 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2009 XThR.Tn[8].t1 XThR.XTB1.Y VPWR.t1366 VPWR.t1365 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2010 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10].t54 XA.XIR[10].XIC_15.icell.Ien VGND.t639 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2011 XA.XIR[0].XIC[14].icell.Ien XThR.Tn[0].t58 VPWR.t88 VPWR.t87 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2012 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[1].t53 VGND.t1956 VGND.t1955 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2013 XA.XIR[1].XIC[8].icell.SM XA.XIR[1].XIC[8].icell.Ien Iout.t229 VGND.t1958 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2014 VGND.t2102 Vbias.t179 XA.XIR[10].XIC[7].icell.SM VGND.t2101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2015 a_n1049_7787# XThR.XTB2.Y VPWR.t1663 VPWR.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2016 XA.XIR[4].XIC[9].icell.SM XA.XIR[4].XIC[9].icell.Ien Iout.t7 VGND.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2017 VGND.t522 XA.Cn[6].t35 XA.XIR[10].XIC[6].icell.PDM VGND.t521 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2018 VPWR.t283 XThR.Tn[12].t55 XA.XIR[13].XIC[4].icell.PUM VPWR.t282 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2019 a_n1331_2891# data[5].t4 VGND.t1977 VGND.t1976 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2020 VGND.t2104 Vbias.t180 XA.XIR[13].XIC[8].icell.SM VGND.t2103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2021 XA.XIR[12].XIC[9].icell.Ien XThR.Tn[12].t56 VPWR.t285 VPWR.t284 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2022 VPWR.t671 VPWR.t669 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t670 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2023 VGND.t694 XA.Cn[7].t27 XA.XIR[13].XIC[7].icell.PDM VGND.t693 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2024 VPWR.t1636 XThR.Tn[14].t55 XA.XIR[15].XIC[5].icell.PUM VPWR.t1635 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2025 XThR.XTB7.B data[6].t1 VGND.t876 VGND.t875 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2026 XThR.Tn[2].t5 XThR.XTBN.Y a_n1049_7493# VPWR.t1790 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2027 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[9].t50 VGND.t452 VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2028 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[9].t51 VGND.t454 VGND.t453 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2029 XA.XIR[2].XIC[11].icell.Ien XThR.Tn[2].t50 VPWR.t1152 VPWR.t1151 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2030 XA.XIR[9].XIC[6].icell.SM XA.XIR[9].XIC[6].icell.Ien Iout.t29 VGND.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2031 VGND.t1458 XA.Cn[12].t34 XA.XIR[1].XIC[12].icell.PDM VGND.t1457 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2032 VGND.t2652 XA.Cn[13].t35 XA.XIR[4].XIC[13].icell.PDM VGND.t2651 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2033 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t2027 XA.XIR[4].XIC_dummy_left.icell.Ien VGND.t2349 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2034 XA.XIR[15].XIC[7].icell.PDM VPWR.t2028 XA.XIR[15].XIC[7].icell.Ien VGND.t2350 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2035 VGND.t2106 Vbias.t181 XA.XIR[0].XIC[0].icell.SM VGND.t2105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2036 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12].t57 XA.XIR[12].XIC[3].icell.Ien VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2037 VPWR.t1765 thermo15c_0.XTBN.Y.t90 XA.Cn[8].t10 VPWR.t1764 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2038 XThR.Tn[10].t3 XThR.XTB3.Y.t12 VPWR.t1227 VPWR.t1226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2039 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7].t53 XA.XIR[7].XIC_15.icell.Ien VGND.t1451 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2040 XA.XIR[11].XIC[4].icell.PUM XA.Cn[4].t36 XA.XIR[11].XIC[4].icell.Ien VPWR.t1912 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2041 XThR.Tn[4].t5 XThR.XTBN.Y VGND.t2401 VGND.t2400 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2042 XA.XIR[15].XIC[12].icell.PUM XA.Cn[12].t35 XA.XIR[15].XIC[12].icell.Ien VPWR.t1392 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2043 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t667 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t668 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2044 XA.XIR[2].XIC[2].icell.Ien XThR.Tn[2].t51 VPWR.t1150 VPWR.t1149 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2045 XA.XIR[11].XIC[13].icell.SM XA.XIR[11].XIC[13].icell.Ien Iout.t112 VGND.t843 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2046 VGND.t1131 XThR.XTB7.B XThR.XTB5.Y VGND.t1130 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2047 VGND.t2108 Vbias.t182 XA.XIR[12].XIC_15.icell.SM VGND.t2107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2048 VGND.t1965 XA.Cn[14].t34 XA.XIR[12].XIC[14].icell.PDM VGND.t1964 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2049 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[3].t60 XA.XIR[3].XIC[1].icell.Ien VGND.t289 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2050 XA.XIR[14].XIC[6].icell.Ien XThR.Tn[14].t56 VPWR.t1638 VPWR.t1637 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2051 VGND.t2009 XA.Cn[8].t35 XA.XIR[12].XIC[8].icell.PDM VGND.t2008 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2052 VPWR.t1423 XThR.Tn[13].t54 XA.XIR[14].XIC[1].icell.PUM VPWR.t1422 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2053 XA.XIR[2].XIC[7].icell.PUM XA.Cn[7].t28 XA.XIR[2].XIC[7].icell.Ien VPWR.t1517 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2054 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[2].t52 XA.XIR[2].XIC[5].icell.Ien VGND.t572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2055 VPWR.t287 XThR.Tn[12].t58 XA.XIR[13].XIC[0].icell.PUM VPWR.t286 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2056 VPWR.t381 XThR.Tn[9].t52 XA.XIR[10].XIC[4].icell.PUM VPWR.t380 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2057 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6].t57 XA.XIR[6].XIC[13].icell.Ien VGND.t2040 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2058 XA.XIR[1].XIC[3].icell.SM XA.XIR[1].XIC[3].icell.Ien Iout.t61 VGND.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2059 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14].t57 XA.XIR[14].XIC[9].icell.Ien VGND.t1978 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2060 VPWR.t1444 XThR.Tn[11].t58 XA.XIR[12].XIC[14].icell.PUM VPWR.t1443 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2061 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t1 VGND.t1417 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2062 XA.Cn[4].t4 thermo15c_0.XTBN.Y.t91 a_5155_9615# VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2063 XA.XIR[13].XIC[4].icell.Ien XThR.Tn[13].t55 VPWR.t1425 VPWR.t1424 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2064 VGND.t2110 Vbias.t183 XA.XIR[10].XIC[2].icell.SM VGND.t2109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2065 XA.XIR[4].XIC[4].icell.SM XA.XIR[4].XIC[4].icell.Ien Iout.t77 VGND.t635 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2066 VGND.t2112 Vbias.t184 XA.XIR[9].XIC_15.icell.SM VGND.t2111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2067 XA.XIR[9].XIC[10].icell.SM XA.XIR[9].XIC[10].icell.Ien Iout.t65 VGND.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2068 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t664 VPWR.t666 VPWR.t665 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2069 VGND.t1360 XA.Cn[10].t35 XA.XIR[1].XIC[10].icell.PDM VGND.t1359 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2070 VGND.t2114 Vbias.t185 XA.XIR[13].XIC[3].icell.SM VGND.t2113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2071 XA.XIR[0].XIC[12].icell.PDM XThR.Tn[0].t59 XA.XIR[0].XIC[12].icell.Ien VGND.t182 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2072 VPWR.t145 XThR.Tn[3].t61 XA.XIR[4].XIC[8].icell.PUM VPWR.t144 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2073 VGND.t2399 XThR.XTBN.Y a_n997_1579# VGND.t2379 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2074 VPWR.t472 XThR.Tn[10].t55 XA.XIR[11].XIC[12].icell.PUM VPWR.t471 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2075 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2029 VGND.t2352 VGND.t2351 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2076 XA.XIR[12].XIC[9].icell.PUM XA.Cn[9].t35 XA.XIR[12].XIC[9].icell.Ien VPWR.t1009 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2077 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12].t59 XA.XIR[12].XIC[7].icell.Ien VGND.t386 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2078 XA.XIR[15].XIC[10].icell.PUM XA.Cn[10].t36 XA.XIR[15].XIC[10].icell.Ien VPWR.t1336 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2079 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[9].t53 VGND.t456 VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2080 XA.XIR[5].XIC[12].icell.SM XA.XIR[5].XIC[12].icell.Ien Iout.t14 VGND.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2081 XA.XIR[9].XIC[1].icell.SM XA.XIR[9].XIC[1].icell.Ien Iout.t225 VGND.t1943 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2082 a_9827_9569# thermo15c_0.XTB5.Y XA.Cn[12].t5 VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2083 XA.XIR[11].XIC[0].icell.PUM XA.Cn[0].t32 XA.XIR[11].XIC[0].icell.Ien VPWR.t1254 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2084 XA.XIR[8].XIC[13].icell.SM XA.XIR[8].XIC[13].icell.Ien Iout.t247 VGND.t2518 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2085 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t662 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t663 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2086 XA.XIR[7].XIC[14].icell.SM XA.XIR[7].XIC[14].icell.Ien Iout.t5 VGND.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2087 XA.XIR[2].XIC[11].icell.PUM XA.Cn[11].t33 XA.XIR[2].XIC[11].icell.Ien VPWR.t331 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2088 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[4].t60 VGND.t1320 VGND.t1319 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2089 XA.XIR[0].XIC[5].icell.PDM VGND.t1668 VGND.t1670 VGND.t1669 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2090 VPWR.t383 XThR.Tn[9].t54 XA.XIR[10].XIC[0].icell.PUM VPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2091 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[3].t62 VGND.t291 VGND.t290 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2092 XA.XIR[2].XIC[12].icell.SM XA.XIR[2].XIC[12].icell.Ien Iout.t165 VGND.t1293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2093 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[11].t59 VGND.t1608 VGND.t1607 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2094 VGND.t2146 XA.Cn[3].t36 XA.XIR[12].XIC[3].icell.PDM VGND.t2145 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2095 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14].t58 VPWR.t1640 VPWR.t1639 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2096 XThR.XTBN.Y XThR.XTBN.A VPWR.t1892 VPWR.t1891 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2097 VGND.t2116 Vbias.t186 XA.XIR[15].XIC[11].icell.SM VGND.t2115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2098 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13].t56 VPWR.t1427 VPWR.t1426 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2099 VPWR.t1387 XThR.Tn[7].t54 XA.XIR[8].XIC[9].icell.PUM VPWR.t1386 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2100 VGND.t1967 XA.Cn[14].t35 XA.XIR[6].XIC[14].icell.PDM VGND.t1966 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2101 XA.XIR[0].XIC[10].icell.PDM XThR.Tn[0].t60 XA.XIR[0].XIC[10].icell.Ien VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2102 XA.XIR[2].XIC[2].icell.PUM XA.Cn[2].t33 XA.XIR[2].XIC[2].icell.Ien VPWR.t1323 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2103 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[2].t53 XA.XIR[2].XIC[0].icell.Ien VGND.t2597 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2104 VGND.t2011 XA.Cn[8].t36 XA.XIR[6].XIC[8].icell.PDM VGND.t2010 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2105 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t659 VPWR.t661 VPWR.t660 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2106 VPWR.t474 XThR.Tn[10].t56 XA.XIR[11].XIC[10].icell.PUM VPWR.t473 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2107 XA.XIR[0].XIC_15.icell.PUM VPWR.t657 XA.XIR[0].XIC_15.icell.Ien VPWR.t658 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2108 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14].t59 XA.XIR[14].XIC[4].icell.Ien VGND.t1979 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2109 XA.XIR[1].XIC[7].icell.Ien XThR.Tn[1].t54 VPWR.t1614 VPWR.t1613 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2110 VGND.t2118 Vbias.t187 XA.XIR[2].XIC[6].icell.SM VGND.t2117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2111 VGND.t2551 XA.Cn[1].t36 XA.XIR[7].XIC[1].icell.PDM VGND.t2550 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2112 VGND.t2033 XA.Cn[5].t32 XA.XIR[2].XIC[5].icell.PDM VGND.t2032 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2113 VPWR.t1788 XThR.XTBN.Y XThR.Tn[11].t9 VPWR.t1768 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2114 XA.XIR[4].XIC[8].icell.Ien XThR.Tn[4].t61 VPWR.t1303 VPWR.t1302 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2115 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[9].t55 VGND.t458 VGND.t457 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2116 VPWR.t1516 data[1].t4 thermo15c_0.XTB7.A VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2117 VPWR.t147 XThR.Tn[3].t63 XA.XIR[4].XIC[3].icell.PUM VPWR.t146 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2118 XA.XIR[11].XIC[12].icell.Ien XThR.Tn[11].t60 VPWR.t1446 VPWR.t1445 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2119 a_8739_9569# thermo15c_0.XTBN.Y.t92 VGND.t2363 VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2120 VGND.t2607 XThR.XTBN.A XThR.XTBN.Y VGND.t2606 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 XA.Cn[6].t10 thermo15c_0.XTB7.Y VGND.t1395 VGND.t1394 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2122 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8].t59 XA.XIR[8].XIC[14].icell.Ien VGND.t1142 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2123 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8].t60 XA.XIR[8].XIC[8].icell.Ien VGND.t1143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2124 XA.XIR[15].XIC[5].icell.PUM XA.Cn[5].t33 XA.XIR[15].XIC[5].icell.Ien VPWR.t1684 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2125 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[0].t61 VGND.t185 VGND.t184 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2126 XA.XIR[6].XIC[9].icell.PUM XA.Cn[9].t36 XA.XIR[6].XIC[9].icell.Ien VPWR.t1010 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2127 XThR.Tn[12].t0 XThR.XTB5.Y a_n997_1803# VGND.t749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2128 VGND.t2354 VPWR.t2030 XA.XIR[1].XIC_dummy_left.icell.PDM VGND.t2353 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2129 VGND.t2120 Vbias.t188 XA.XIR[12].XIC[8].icell.SM VGND.t2119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2130 VGND.t407 XA.Cn[11].t34 XA.XIR[3].XIC[11].icell.PDM VGND.t406 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2131 VGND.t1788 XA.Cn[7].t29 XA.XIR[12].XIC[7].icell.PDM VGND.t1787 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2132 VGND.t2122 Vbias.t189 XA.XIR[15].XIC[9].icell.SM VGND.t2121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2133 a_n997_3979# XThR.XTBN.Y VGND.t2396 VGND.t2395 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2134 thermo15c_0.XTB7.Y thermo15c_0.XTB7.B VGND.t1099 VGND.t1098 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2135 XA.XIR[0].XIC[0].icell.PDM VGND.t1665 VGND.t1667 VGND.t1666 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2136 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t654 VPWR.t656 VPWR.t655 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2137 VGND.t2124 Vbias.t190 XA.XIR[6].XIC[7].icell.SM VGND.t2123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2138 XA.XIR[1].XIC[11].icell.Ien XThR.Tn[1].t55 VPWR.t1707 VPWR.t1706 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2139 VGND.t935 Vbias.t191 XA.XIR[2].XIC[10].icell.SM VGND.t934 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2140 XA.Cn[8].t9 thermo15c_0.XTBN.Y.t93 VPWR.t1767 VPWR.t1766 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2141 VGND.t2132 XA.Cn[1].t37 XA.XIR[4].XIC[1].icell.PDM VGND.t2131 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2142 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[11].t61 VGND.t1610 VGND.t1609 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2143 VGND.t1339 XA.Cn[2].t34 XA.XIR[3].XIC[2].icell.PDM VGND.t1338 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2144 VGND.t937 Vbias.t192 XA.XIR[9].XIC[8].icell.SM VGND.t936 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2145 XA.XIR[14].XIC[7].icell.PUM XA.Cn[7].t30 XA.XIR[14].XIC[7].icell.Ien VPWR.t1518 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2146 XA.XIR[8].XIC[9].icell.Ien XThR.Tn[8].t61 VPWR.t1224 VPWR.t1223 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2147 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t2031 VGND.t2356 VGND.t2355 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2148 VGND.t1883 XA.Cn[3].t37 XA.XIR[6].XIC[3].icell.PDM VGND.t1882 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2149 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5].t55 XA.XIR[5].XIC[11].icell.Ien VGND.t1766 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2150 XA.XIR[11].XIC[10].icell.Ien XThR.Tn[11].t62 VPWR.t1448 VPWR.t1447 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2151 a_n1049_6699# XThR.XTB4.Y.t12 VPWR.t1284 VPWR.t1228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2152 XA.XIR[13].XIC_15.icell.SM XA.XIR[13].XIC_15.icell.Ien Iout.t4 VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2153 VPWR.t476 XThR.Tn[10].t57 XA.XIR[11].XIC[5].icell.PUM VPWR.t475 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2154 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9].t56 XA.XIR[9].XIC[11].icell.Ien VGND.t459 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2155 XA.XIR[10].XIC[4].icell.PUM XA.Cn[4].t37 XA.XIR[10].XIC[4].icell.Ien VPWR.t1913 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2156 XA.XIR[1].XIC[2].icell.Ien XThR.Tn[1].t56 VPWR.t1709 VPWR.t1708 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2157 VGND.t939 Vbias.t193 XA.XIR[2].XIC[1].icell.SM VGND.t938 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2158 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t652 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t653 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2159 XA.XIR[6].XIC[5].icell.SM XA.XIR[6].XIC[5].icell.Ien Iout.t160 VGND.t1164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2160 VGND.t1216 XA.Cn[0].t33 XA.XIR[2].XIC[0].icell.PDM VGND.t1215 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2161 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t650 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t651 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2162 XA.XIR[4].XIC[3].icell.Ien XThR.Tn[4].t62 VPWR.t1305 VPWR.t1304 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2163 VGND.t941 Vbias.t194 XA.XIR[0].XIC[14].icell.SM VGND.t940 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2164 VGND.t943 Vbias.t195 XA.XIR[14].XIC[5].icell.SM VGND.t942 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2165 VGND.t2654 XA.Cn[13].t36 XA.XIR[0].XIC[13].icell.PDM VGND.t2653 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2166 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6].t58 XA.XIR[6].XIC[1].icell.Ien VGND.t2041 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2167 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t2032 XA.XIR[0].XIC_dummy_left.icell.Ien VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2168 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[1].t57 XA.XIR[1].XIC[5].icell.Ien VGND.t2088 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2169 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5].t56 XA.XIR[5].XIC[2].icell.Ien VGND.t1767 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2170 VGND.t576 VPWR.t2033 XA.XIR[13].XIC_dummy_right.icell.PDM VGND.t575 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2171 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9].t57 XA.XIR[9].XIC[2].icell.Ien VGND.t460 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2172 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8].t62 XA.XIR[8].XIC[3].icell.Ien VGND.t1144 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2173 XA.XIR[3].XIC_15.icell.PDM XThR.Tn[3].t64 XA.XIR[3].XIC_15.icell.Ien VGND.t292 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2174 VGND.t2264 data[1].t5 thermo15c_0.XTB6.A VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2175 VPWR.t1642 XThR.Tn[14].t60 XA.XIR[15].XIC[14].icell.PUM VPWR.t1641 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2176 VPWR.t649 VPWR.t647 XA.XIR[14].XIC_15.icell.PUM VPWR.t648 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2177 a_n997_2891# XThR.XTBN.Y VGND.t2394 VGND.t2393 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2178 VGND.t945 Vbias.t196 XA.XIR[12].XIC[3].icell.SM VGND.t944 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2179 VGND.t947 Vbias.t197 XA.XIR[3].XIC[7].icell.SM VGND.t946 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2180 VGND.t524 XA.Cn[6].t36 XA.XIR[3].XIC[6].icell.PDM VGND.t523 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2181 XA.XIR[14].XIC[11].icell.PUM XA.Cn[11].t35 XA.XIR[14].XIC[11].icell.Ien VPWR.t332 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2182 VPWR.t1481 XThR.Tn[5].t57 XA.XIR[6].XIC[4].icell.PUM VPWR.t1480 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2183 VPWR.t646 VPWR.t644 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t645 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2184 VGND.t949 Vbias.t198 XA.XIR[15].XIC[4].icell.SM VGND.t948 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2185 VGND.t1664 VGND.t1662 XA.XIR[10].XIC_dummy_right.icell.SM VGND.t1663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2186 VGND.t1790 XA.Cn[7].t31 XA.XIR[6].XIC[7].icell.PDM VGND.t1789 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2187 VPWR.t643 VPWR.t641 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t642 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2188 VPWR.t289 XThR.Tn[12].t60 XA.XIR[13].XIC[13].icell.PUM VPWR.t288 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2189 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t2034 XA.XIR[15].XIC_dummy_right.icell.Ien VGND.t577 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2190 XThR.Tn[11].t0 XThR.XTB4.Y.t13 a_n997_2667# VGND.t1226 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2191 VGND.t951 Vbias.t199 XA.XIR[6].XIC[2].icell.SM VGND.t950 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2192 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[6].t59 VGND.t2043 VGND.t2042 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2193 VPWR.t336 thermo15c_0.XTB5.Y a_5155_9615# VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2194 XA.XIR[10].XIC[0].icell.PUM XA.Cn[0].t34 XA.XIR[10].XIC[0].icell.Ien VPWR.t1255 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2195 XA.XIR[3].XIC[5].icell.SM XA.XIR[3].XIC[5].icell.Ien Iout.t23 VGND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2196 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[2].t54 VGND.t2596 VGND.t2595 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2197 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[2].t55 VGND.t2594 VGND.t2593 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2198 VGND.t953 Vbias.t200 XA.XIR[9].XIC[3].icell.SM VGND.t952 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2199 XA.XIR[14].XIC[2].icell.PUM XA.Cn[2].t35 XA.XIR[14].XIC[2].icell.Ien VPWR.t1324 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2200 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5].t58 XA.XIR[5].XIC[6].icell.Ien VGND.t1768 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2201 XA.XIR[11].XIC[5].icell.Ien XThR.Tn[11].t63 VPWR.t1896 VPWR.t1895 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2202 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[3].t65 VGND.t294 VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2203 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9].t58 XA.XIR[9].XIC[6].icell.Ien VGND.t461 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2204 VGND.t418 XA.Cn[5].t34 XA.XIR[14].XIC[5].icell.PDM VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2205 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8].t63 XA.XIR[8].XIC[7].icell.Ien VGND.t1145 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2206 VGND.t2392 XThR.XTBN.Y XThR.Tn[0].t9 VGND.t2391 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2207 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[6].t60 VGND.t2045 VGND.t2044 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2208 XA.XIR[1].XIC[8].icell.PUM XA.Cn[8].t37 XA.XIR[1].XIC[8].icell.Ien VPWR.t1674 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2209 a_n1049_6405# XThR.XTB5.Y VPWR.t1229 VPWR.t1228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2210 XA.XIR[6].XIC[0].icell.SM XA.XIR[6].XIC[0].icell.Ien Iout.t35 VGND.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2211 XThR.Tn[8].t0 XThR.XTB1.Y VPWR.t1364 VPWR.t1363 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2212 XA.XIR[1].XIC[12].icell.SM XA.XIR[1].XIC[12].icell.Ien Iout.t251 VGND.t2619 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2213 XA.XIR[8].XIC[12].icell.PUM XA.Cn[12].t36 XA.XIR[8].XIC[12].icell.Ien VPWR.t1393 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2214 VGND.t955 Vbias.t201 XA.XIR[14].XIC[0].icell.SM VGND.t954 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2215 XA.XIR[15].XIC[9].icell.PDM XThR.Tn[14].t61 VGND.t1981 VGND.t1980 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2216 XA.XIR[4].XIC[13].icell.SM XA.XIR[4].XIC[13].icell.Ien Iout.t84 VGND.t681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2217 XA.XIR[5].XIC_15.icell.PDM VPWR.t2035 VGND.t579 VGND.t578 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2218 VGND.t957 Vbias.t202 XA.XIR[5].XIC_15.icell.SM VGND.t956 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2219 XA.XIR[11].XIC[13].icell.PUM XA.Cn[13].t37 XA.XIR[11].XIC[13].icell.Ien VPWR.t1922 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2220 VGND.t1038 XA.Cn[8].t38 XA.XIR[5].XIC[8].icell.PDM VGND.t1037 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2221 VGND.t1969 XA.Cn[14].t36 XA.XIR[5].XIC[14].icell.PDM VGND.t1968 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2222 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[1].t58 XA.XIR[1].XIC[0].icell.Ien VGND.t2089 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2223 VGND.t2495 Vbias.t203 XA.XIR[13].XIC[12].icell.SM VGND.t2494 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2224 XThR.Tn[1].t1 XThR.XTB2.Y VGND.t2000 VGND.t1423 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2225 VGND.t1971 XA.Cn[14].t37 XA.XIR[9].XIC[14].icell.PDM VGND.t1970 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2226 VGND.t1040 XA.Cn[8].t39 XA.XIR[9].XIC[8].icell.PDM VGND.t1039 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2227 VPWR.t1483 XThR.Tn[5].t59 XA.XIR[6].XIC[0].icell.PUM VPWR.t1482 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2228 VGND.t1284 thermo15c_0.XTBN.Y.t94 a_8739_9569# VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2229 XA.XIR[14].XIC_15.icell.Ien XThR.Tn[14].t62 VPWR.t1644 VPWR.t1643 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2230 VGND.t2497 Vbias.t204 XA.XIR[1].XIC[6].icell.SM VGND.t2496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2231 VPWR.t640 VPWR.t638 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t639 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2232 XA.Cn[1].t10 thermo15c_0.XTB2.Y VGND.t1940 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2233 VGND.t1393 thermo15c_0.XTB7.Y XA.Cn[6].t9 VGND.t1392 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2234 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t2036 XA.XIR[12].XIC_dummy_right.icell.Ien VGND.t580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2235 VPWR.t385 XThR.Tn[9].t59 XA.XIR[10].XIC[13].icell.PUM VPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2236 VPWR.t637 VPWR.t635 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t636 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2237 a_6243_9615# thermo15c_0.XTBN.Y.t95 XA.Cn[6].t1 VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2238 VGND.t2499 Vbias.t205 XA.XIR[3].XIC[2].icell.SM VGND.t2498 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2239 VGND.t2501 Vbias.t206 XA.XIR[11].XIC[11].icell.SM VGND.t2500 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2240 XA.XIR[10].XIC[12].icell.Ien XThR.Tn[10].t58 VPWR.t478 VPWR.t477 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2241 XThR.Tn[2].t4 XThR.XTBN.Y a_n1049_7493# VPWR.t1787 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2242 VGND.t582 VPWR.t2037 XA.XIR[7].XIC_15.icell.PDM VGND.t581 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2243 XA.XIR[10].XIC[7].icell.SM XA.XIR[10].XIC[7].icell.Ien Iout.t122 VGND.t1027 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2244 XA.XIR[13].XIC[13].icell.Ien XThR.Tn[13].t57 VPWR.t1429 VPWR.t1428 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2245 XA.XIR[13].XIC[8].icell.SM XA.XIR[13].XIC[8].icell.Ien Iout.t150 VGND.t1122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2246 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[0].t62 VGND.t187 VGND.t186 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2247 XThR.Tn[13].t8 XThR.XTBN.Y VPWR.t1786 VPWR.t1785 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2248 XA.XIR[5].XIC[9].icell.PUM XA.Cn[9].t37 XA.XIR[5].XIC[9].icell.Ien VPWR.t1011 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2249 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[6].t61 VGND.t2047 VGND.t2046 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2250 XA.XIR[0].XIC[8].icell.Ien XThR.Tn[0].t63 VPWR.t90 VPWR.t89 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2251 XA.XIR[3].XIC[0].icell.SM XA.XIR[3].XIC[0].icell.Ien Iout.t135 VGND.t1060 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2252 XA.XIR[9].XIC[9].icell.PUM XA.Cn[9].t38 XA.XIR[9].XIC[9].icell.Ien VPWR.t1570 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2253 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[2].t56 VGND.t2592 VGND.t2591 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2254 XThR.Tn[10].t5 XThR.XTB3.Y.t13 VPWR.t1507 VPWR.t1506 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2255 XA.XIR[8].XIC[10].icell.PUM XA.Cn[10].t37 XA.XIR[8].XIC[10].icell.Ien VPWR.t1337 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2256 XThR.Tn[4].t4 XThR.XTBN.Y VGND.t2390 VGND.t2389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2257 VPWR.t291 XThR.Tn[12].t61 XA.XIR[13].XIC[6].icell.PUM VPWR.t290 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2258 VGND.t1661 VGND.t1659 XA.XIR[10].XIC_dummy_left.icell.SM VGND.t1660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2259 VGND.t746 XThR.XTB6.Y XThR.Tn[5].t0 VGND.t745 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2260 VGND.t1218 XA.Cn[0].t35 XA.XIR[14].XIC[0].icell.PDM VGND.t1217 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2261 XA.XIR[1].XIC[3].icell.PUM XA.Cn[3].t38 XA.XIR[1].XIC[3].icell.Ien VPWR.t1572 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2262 VGND.t2503 Vbias.t207 XA.XIR[1].XIC[10].icell.SM VGND.t2502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2263 a_4861_9615# thermo15c_0.XTBN.Y.t96 XA.Cn[3].t5 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2264 XA.XIR[15].XIC[4].icell.PDM XThR.Tn[14].t63 VGND.t1983 VGND.t1982 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2265 XA.XIR[0].XIC[11].icell.SM XA.XIR[0].XIC[11].icell.Ien Iout.t22 VGND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2266 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[13].t58 VGND.t1532 VGND.t1531 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2267 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2038 VGND.t584 VGND.t583 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2268 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t0 VGND.t1414 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2269 VGND.t1885 XA.Cn[3].t39 XA.XIR[5].XIC[3].icell.PDM VGND.t1884 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2270 VGND.t2505 Vbias.t208 XA.XIR[11].XIC[9].icell.SM VGND.t2504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2271 XA.XIR[10].XIC[10].icell.Ien XThR.Tn[10].t59 VPWR.t480 VPWR.t479 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2272 XA.XIR[12].XIC_15.icell.SM XA.XIR[12].XIC_15.icell.Ien Iout.t76 VGND.t573 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2273 VGND.t1887 XA.Cn[3].t40 XA.XIR[9].XIC[3].icell.PDM VGND.t1886 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2274 VGND.t2507 Vbias.t209 XA.XIR[8].XIC[11].icell.SM VGND.t2506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2275 XA.XIR[7].XIC[12].icell.Ien XThR.Tn[7].t55 VPWR.t1398 VPWR.t1397 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2276 VPWR.t460 XThR.Tn[0].t64 XA.XIR[1].XIC[9].icell.PUM VPWR.t459 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2277 VGND.t586 VPWR.t2039 XA.XIR[4].XIC_15.icell.PDM VGND.t585 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2278 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t632 VPWR.t634 VPWR.t633 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2279 VGND.t2509 Vbias.t210 XA.XIR[1].XIC[1].icell.SM VGND.t2508 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2280 VPWR.t1307 XThR.Tn[4].t63 XA.XIR[5].XIC[9].icell.PUM VPWR.t1306 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2281 VGND.t2134 XA.Cn[1].t38 XA.XIR[0].XIC[1].icell.PDM VGND.t2133 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2282 XA.XIR[11].XIC[6].icell.PUM XA.Cn[6].t37 XA.XIR[11].XIC[6].icell.Ien VPWR.t434 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2283 XA.XIR[15].XIC[14].icell.PUM XA.Cn[14].t38 XA.XIR[15].XIC[14].icell.Ien VPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2284 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[2].t57 VGND.t2590 VGND.t2589 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2285 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14].t64 XA.XIR[14].XIC[13].icell.Ien VGND.t1984 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2286 VGND.t588 VPWR.t2040 XA.XIR[12].XIC_dummy_right.icell.PDM VGND.t587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2287 XA.XIR[10].XIC[2].icell.SM XA.XIR[10].XIC[2].icell.Ien Iout.t231 VGND.t1975 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2288 VGND.t1875 XA.Cn[9].t39 XA.XIR[11].XIC[9].icell.PDM VGND.t1874 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2289 VPWR.t454 XThR.XTB3.Y.t14 a_n1049_7493# VPWR.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2290 XA.XIR[13].XIC[3].icell.SM XA.XIR[13].XIC[3].icell.Ien Iout.t171 VGND.t1370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2291 VPWR.t402 XThR.Tn[9].t60 XA.XIR[10].XIC[6].icell.PUM VPWR.t401 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2292 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6].t62 XA.XIR[6].XIC_15.icell.Ien VGND.t2048 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2293 VPWR.t1898 XThR.Tn[11].t64 XA.XIR[12].XIC[8].icell.PUM VPWR.t1897 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2294 XA.XIR[0].XIC[3].icell.Ien XThR.Tn[0].t65 VPWR.t462 VPWR.t461 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2295 XA.XIR[8].XIC[5].icell.PUM XA.Cn[5].t35 XA.XIR[8].XIC[5].icell.Ien VPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2296 XA.XIR[13].XIC[6].icell.Ien XThR.Tn[13].t59 VPWR.t1431 VPWR.t1430 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2297 XA.XIR[0].XIC[9].icell.SM XA.XIR[0].XIC[9].icell.Ien Iout.t28 VGND.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2298 VGND.t2511 Vbias.t211 XA.XIR[5].XIC[8].icell.SM VGND.t2510 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2299 VGND.t1792 XA.Cn[7].t32 XA.XIR[5].XIC[7].icell.PDM VGND.t1791 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2300 VPWR.t293 XThR.Tn[12].t62 XA.XIR[13].XIC[1].icell.PUM VPWR.t292 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2301 thermo15c_0.XTB2.Y thermo15c_0.XTB6.A a_3523_10575# VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2302 VPWR.t631 VPWR.t629 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t630 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2303 VGND.t1794 XA.Cn[7].t33 XA.XIR[9].XIC[7].icell.PDM VGND.t1793 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2304 VGND.t2513 Vbias.t212 XA.XIR[8].XIC[9].icell.SM VGND.t2512 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2305 XA.XIR[7].XIC[10].icell.Ien XThR.Tn[7].t56 VPWR.t1400 VPWR.t1399 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2306 XThR.Tn[4].t1 XThR.XTB5.Y VGND.t1166 VGND.t747 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2307 VPWR.t1784 XThR.XTBN.Y XThR.Tn[14].t8 VPWR.t1783 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2308 VPWR.t482 XThR.Tn[10].t60 XA.XIR[11].XIC[14].icell.PUM VPWR.t481 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2309 XA.Cn[13].t1 thermo15c_0.XTB6.Y VPWR.t1033 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2310 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13].t60 XA.XIR[13].XIC[9].icell.Ien VGND.t1533 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2311 VGND.t897 thermo15c_0.XTB6.Y XA.Cn[5].t0 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2312 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[13].t61 VGND.t1535 VGND.t1534 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2313 XA.XIR[5].XIC[6].icell.SM XA.XIR[5].XIC[6].icell.Ien Iout.t74 VGND.t564 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2314 VPWR.t1782 XThR.XTBN.Y XThR.Tn[11].t8 VPWR.t1781 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2315 VGND.t2515 Vbias.t213 XA.XIR[11].XIC[4].icell.SM VGND.t2514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2316 XA.XIR[10].XIC[5].icell.Ien XThR.Tn[10].t61 VPWR.t484 VPWR.t483 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2317 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[12].t63 VGND.t388 VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2318 VGND.t1658 VGND.t1656 XA.XIR[6].XIC_dummy_right.icell.SM VGND.t1657 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2319 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[11].t65 VGND.t2611 VGND.t2610 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2320 XA.XIR[15].XIC[11].icell.SM XA.XIR[15].XIC[11].icell.Ien Iout.t21 VGND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2321 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[2].t58 XA.XIR[2].XIC[11].icell.Ien VGND.t2588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2322 XA.XIR[3].XIC[4].icell.PUM XA.Cn[4].t38 XA.XIR[3].XIC[4].icell.Ien VPWR.t1845 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2323 XA.Cn[9].t8 thermo15c_0.XTB2.Y a_7875_9569# VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2324 XA.XIR[4].XIC_15.icell.PDM VPWR.t2041 VGND.t590 VGND.t589 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2325 XA.XIR[11].XIC[1].icell.PUM XA.Cn[1].t39 XA.XIR[11].XIC[1].icell.Ien VPWR.t1719 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2326 VGND.t1127 thermo15c_0.XTB6.A thermo15c_0.XTB6.Y VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2327 VGND.t1939 thermo15c_0.XTB2.Y XA.Cn[1].t9 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 XA.XIR[10].XIC[13].icell.PUM XA.Cn[13].t38 XA.XIR[10].XIC[13].icell.Ien VPWR.t1923 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2329 XA.XIR[2].XIC[6].icell.SM XA.XIR[2].XIC[6].icell.Ien Iout.t64 VGND.t437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2330 VGND.t2517 Vbias.t214 XA.XIR[12].XIC[12].icell.SM VGND.t2516 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2331 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t627 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t628 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2332 XA.Cn[6].t0 thermo15c_0.XTBN.Y.t97 a_6243_9615# VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2333 XA.XIR[6].XIC[14].icell.SM XA.XIR[6].XIC[14].icell.Ien Iout.t19 VGND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2334 VGND.t1186 Vbias.t215 XA.XIR[15].XIC[13].icell.SM VGND.t1185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2335 VGND.t1188 Vbias.t216 XA.XIR[14].XIC[14].icell.SM VGND.t1187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2336 VGND.t1460 XA.Cn[12].t37 XA.XIR[15].XIC[12].icell.PDM VGND.t1459 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2337 VGND.t2484 XA.Cn[4].t39 XA.XIR[11].XIC[4].icell.PDM VGND.t2483 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2338 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[2].t59 XA.XIR[2].XIC[2].icell.Ien VGND.t2587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2339 VPWR.t1018 XThR.XTB7.Y a_n1049_5317# VPWR.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2340 VPWR.t404 XThR.Tn[9].t61 XA.XIR[10].XIC[1].icell.PUM VPWR.t403 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2341 VGND.t592 VPWR.t2042 XA.XIR[6].XIC_dummy_right.icell.PDM VGND.t591 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2342 VPWR.t1032 thermo15c_0.XTB6.Y XA.Cn[13].t0 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2343 VPWR.t1900 XThR.Tn[11].t66 XA.XIR[12].XIC[3].icell.PUM VPWR.t1899 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2344 a_n997_3979# XThR.XTBN.Y VGND.t2388 VGND.t2387 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2345 XA.XIR[5].XIC[4].icell.Ien XThR.Tn[5].t60 VPWR.t1485 VPWR.t1484 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2346 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13].t62 VPWR.t1433 VPWR.t1432 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2347 XA.XIR[9].XIC[4].icell.Ien XThR.Tn[9].t62 VPWR.t406 VPWR.t405 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2348 XA.XIR[0].XIC[4].icell.SM XA.XIR[0].XIC[4].icell.Ien Iout.t103 VGND.t810 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2349 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t624 VPWR.t626 VPWR.t625 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2350 VGND.t1190 Vbias.t217 XA.XIR[5].XIC[3].icell.SM VGND.t1189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2351 VGND.t1192 Vbias.t218 XA.XIR[9].XIC[12].icell.SM VGND.t1191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2352 XA.XIR[9].XIC[7].icell.SM XA.XIR[9].XIC[7].icell.Ien Iout.t127 VGND.t1034 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2353 VGND.t1227 XThR.XTB4.Y.t14 XThR.Tn[3].t0 VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2354 XA.XIR[5].XIC[10].icell.SM XA.XIR[5].XIC[10].icell.Ien Iout.t180 VGND.t1387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2355 a_7331_10587# data[0].t2 VPWR.t951 VPWR.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2356 a_4067_9615# thermo15c_0.XTBN.Y.t98 XA.Cn[2].t7 VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2357 VPWR.t1148 XThR.Tn[2].t60 XA.XIR[3].XIC[12].icell.PUM VPWR.t1147 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2358 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[12].t64 VGND.t390 VGND.t389 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2359 XA.XIR[12].XIC[8].icell.SM XA.XIR[12].XIC[8].icell.Ien Iout.t24 VGND.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2360 XA.XIR[11].XIC[14].icell.Ien XThR.Tn[11].t67 VPWR.t1902 VPWR.t1901 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2361 VGND.t1194 Vbias.t219 XA.XIR[8].XIC[4].icell.SM VGND.t1193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2362 VGND.t1655 VGND.t1653 XA.XIR[3].XIC_dummy_right.icell.SM VGND.t1654 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2363 XA.XIR[7].XIC[5].icell.Ien XThR.Tn[7].t57 VPWR.t1402 VPWR.t1401 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2364 VPWR.t1694 XThR.Tn[6].t63 XA.XIR[7].XIC[12].icell.PUM VPWR.t1693 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2365 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13].t63 XA.XIR[13].XIC[4].icell.Ien VGND.t1522 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2366 XA.XIR[15].XIC[9].icell.SM XA.XIR[15].XIC[9].icell.Ien Iout.t170 VGND.t1369 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2367 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t2043 XA.XIR[8].XIC_dummy_right.icell.Ien VGND.t593 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2368 VPWR.t1487 XThR.Tn[5].t61 XA.XIR[6].XIC[13].icell.PUM VPWR.t1486 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2369 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t4 VPWR.t1780 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2370 XA.XIR[0].XIC[11].icell.PDM VGND.t1650 VGND.t1652 VGND.t1651 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2371 XA.XIR[3].XIC[0].icell.PUM XA.Cn[0].t36 XA.XIR[3].XIC[0].icell.Ien VPWR.t1256 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2372 XA.XIR[1].XIC_15.icell.PDM VPWR.t2044 VGND.t595 VGND.t594 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2373 XA.XIR[5].XIC[1].icell.SM XA.XIR[5].XIC[1].icell.Ien Iout.t107 VGND.t825 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2374 XA.XIR[2].XIC[10].icell.SM XA.XIR[2].XIC[10].icell.Ien Iout.t111 VGND.t839 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2375 XA.Cn[3].t4 thermo15c_0.XTBN.Y.t99 a_4861_9615# VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2376 XA.XIR[3].XIC[14].icell.SM XA.XIR[3].XIC[14].icell.Ien Iout.t88 VGND.t736 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2377 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t622 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t623 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2378 thermo15c_0.XTB5.A data[0].t3 VGND.t775 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2379 VGND.t1362 XA.Cn[10].t38 XA.XIR[15].XIC[10].icell.PDM VGND.t1361 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2380 VPWR.t1269 XThR.XTB4.Y.t15 XThR.Tn[11].t1 VPWR.t1242 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2381 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[2].t61 XA.XIR[2].XIC[6].icell.Ien VGND.t1561 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2382 XA.XIR[0].XIC[2].icell.PDM VGND.t1647 VGND.t1649 VGND.t1648 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2383 XA.XIR[2].XIC[1].icell.SM XA.XIR[2].XIC[1].icell.Ien Iout.t96 VGND.t744 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2384 VGND.t409 XA.Cn[11].t36 XA.XIR[2].XIC[11].icell.PDM VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2385 VGND.t2386 XThR.XTBN.Y a_n997_715# VGND.t2385 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2386 a_n997_2891# XThR.XTBN.Y VGND.t2384 VGND.t2383 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2387 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[7].t58 VGND.t1468 VGND.t1467 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2388 VGND.t1646 VGND.t1644 XA.XIR[6].XIC_dummy_left.icell.SM VGND.t1645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2389 XA.XIR[5].XIC[0].icell.Ien XThR.Tn[5].t62 VPWR.t1258 VPWR.t1257 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2390 VPWR.t149 XThR.Tn[3].t66 XA.XIR[4].XIC[9].icell.PUM VPWR.t148 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2391 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9].t63 VPWR.t408 VPWR.t407 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2392 VPWR.t1146 XThR.Tn[2].t62 XA.XIR[3].XIC[10].icell.PUM VPWR.t1145 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2393 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t619 VPWR.t621 VPWR.t620 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2394 VPWR.t1696 XThR.Tn[6].t64 XA.XIR[7].XIC[10].icell.PUM VPWR.t1695 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2395 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14].t65 XA.XIR[14].XIC[1].icell.Ien VGND.t1985 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2396 XA.XIR[10].XIC[6].icell.PUM XA.Cn[6].t38 XA.XIR[10].XIC[6].icell.Ien VPWR.t468 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2397 XThR.Tn[11].t2 XThR.XTB4.Y.t16 a_n997_2667# VGND.t1228 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2398 VPWR.t618 VPWR.t616 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t617 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2399 VGND.t2083 XA.Cn[2].t36 XA.XIR[2].XIC[2].icell.PDM VGND.t2082 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2400 XA.XIR[13].XIC[7].icell.PUM XA.Cn[7].t34 XA.XIR[13].XIC[7].icell.Ien VPWR.t1519 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2401 XA.XIR[9].XIC[2].icell.SM XA.XIR[9].XIC[2].icell.Ien Iout.t155 VGND.t1156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2402 VPWR.t1594 thermo15c_0.XTB2.Y XA.Cn[9].t4 VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2403 XA.XIR[3].XIC[12].icell.Ien XThR.Tn[3].t67 VPWR.t151 VPWR.t150 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2404 a_n997_3979# XThR.XTB1.Y XThR.Tn[8].t5 VGND.t1417 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2405 VGND.t597 VPWR.t2045 XA.XIR[0].XIC_15.icell.PDM VGND.t596 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2406 VGND.t1877 XA.Cn[9].t40 XA.XIR[10].XIC[9].icell.PDM VGND.t1876 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2407 XA.XIR[12].XIC[3].icell.SM XA.XIR[12].XIC[3].icell.Ien Iout.t190 VGND.t1443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2408 VPWR.t1294 thermo15c_0.XTBN.Y.t100 XA.Cn[8].t8 VPWR.t1293 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2409 XA.XIR[15].XIC[4].icell.SM XA.XIR[15].XIC[4].icell.Ien Iout.t224 VGND.t1942 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2410 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[4].t64 XA.XIR[4].XIC[8].icell.Ien VGND.t1321 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2411 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[4].t65 XA.XIR[4].XIC[14].icell.Ien VGND.t1322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2412 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout VGND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2413 a_n1335_8331# XThR.XTB5.A XThR.XTB1.Y VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2414 VPWR.t1646 XThR.Tn[14].t66 XA.XIR[15].XIC[8].icell.PUM VPWR.t1645 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2415 XA.XIR[0].XIC[6].icell.PDM VGND.t1641 VGND.t1643 VGND.t1642 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2416 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11].t68 XA.XIR[11].XIC[12].icell.Ien VGND.t2612 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2417 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t8 VPWR.t1780 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2418 XA.XIR[15].XIC[7].icell.Ien VPWR.t613 VPWR.t615 VPWR.t614 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2419 XThR.Tn[7].t0 XThR.XTBN.Y VPWR.t1779 VPWR.t1778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2420 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2046 VGND.t599 VGND.t598 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2421 VPWR.t1260 XThR.Tn[5].t63 XA.XIR[6].XIC[6].icell.PUM VPWR.t1259 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2422 VGND.t1640 VGND.t1638 XA.XIR[3].XIC_dummy_left.icell.SM VGND.t1639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2423 VPWR.t131 XThR.Tn[8].t64 XA.XIR[9].XIC[7].icell.PUM VPWR.t130 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2424 XA.Cn[9].t0 thermo15c_0.XTBN.Y.t101 VPWR.t1295 VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2425 XThR.Tn[1].t9 XThR.XTBN.Y VGND.t2382 VGND.t2381 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2426 VPWR.t599 VPWR.t597 XA.XIR[13].XIC_15.icell.PUM VPWR.t598 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2427 VGND.t1196 Vbias.t220 XA.XIR[2].XIC[7].icell.SM VGND.t1195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2428 VGND.t556 XA.Cn[6].t39 XA.XIR[2].XIC[6].icell.PDM VGND.t555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2429 XA.XIR[13].XIC[11].icell.PUM XA.Cn[11].t37 XA.XIR[13].XIC[11].icell.Ien VPWR.t333 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2430 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[11].t69 VGND.t2614 VGND.t2613 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2431 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[7].t59 VGND.t1470 VGND.t1469 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2432 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2047 VGND.t601 VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2433 XA.XIR[4].XIC[9].icell.Ien XThR.Tn[4].t66 VPWR.t1309 VPWR.t1308 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2434 XA.XIR[3].XIC[10].icell.Ien XThR.Tn[3].t68 VPWR.t153 VPWR.t152 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2435 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[10].t62 VGND.t2151 VGND.t2150 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2436 XA.XIR[14].XIC[11].icell.SM XA.XIR[14].XIC[11].icell.Ien Iout.t47 VGND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2437 XA.XIR[15].XIC[13].icell.PDM XThR.Tn[14].t67 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2438 VPWR.t1296 thermo15c_0.XTBN.Y.t102 XA.Cn[11].t4 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2439 VPWR.t1144 XThR.Tn[2].t63 XA.XIR[3].XIC[5].icell.PUM VPWR.t1143 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2440 VPWR.t542 XThR.XTB6.Y a_n1049_5611# VPWR.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2441 VGND.t603 VPWR.t2048 XA.XIR[15].XIC_dummy_left.icell.PDM VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2442 a_n997_2891# XThR.XTB3.Y.t15 XThR.Tn[10].t2 VGND.t913 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2443 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[1].t59 XA.XIR[1].XIC[11].icell.Ien VGND.t2090 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2444 XA.XIR[13].XIC[12].icell.SM XA.XIR[13].XIC[12].icell.Ien Iout.t140 VGND.t1096 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2445 VPWR.t1698 XThR.Tn[6].t65 XA.XIR[7].XIC[5].icell.PUM VPWR.t1697 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2446 XA.XIR[10].XIC[1].icell.PUM XA.Cn[1].t40 XA.XIR[10].XIC[1].icell.Ien VPWR.t1720 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2447 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t611 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t612 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2448 XA.XIR[1].XIC[6].icell.SM XA.XIR[1].XIC[6].icell.Ien Iout.t118 VGND.t896 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2449 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[1].t60 VGND.t2092 VGND.t2091 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2450 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[1].t61 VGND.t2094 VGND.t2093 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2451 XA.XIR[13].XIC[2].icell.PUM XA.Cn[2].t37 XA.XIR[13].XIC[2].icell.Ien VPWR.t1701 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2452 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11].t70 XA.XIR[11].XIC[10].icell.Ien VGND.t2586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2453 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[8].t65 VGND.t232 VGND.t231 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2454 XA.XIR[8].XIC[14].icell.PUM XA.Cn[14].t39 XA.XIR[8].XIC[14].icell.Ien VPWR.t78 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2455 VGND.t1198 Vbias.t221 XA.XIR[10].XIC[5].icell.SM VGND.t1197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2456 XA.XIR[15].XIC[11].icell.Ien VPWR.t608 VPWR.t610 VPWR.t609 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2457 VGND.t2486 XA.Cn[4].t40 XA.XIR[10].XIC[4].icell.PDM VGND.t2485 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2458 VGND.t605 VPWR.t2049 XA.XIR[5].XIC_dummy_right.icell.PDM VGND.t604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2459 XA.XIR[11].XIC_15.icell.PUM VPWR.t606 XA.XIR[11].XIC_15.icell.Ien VPWR.t607 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2460 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[1].t62 XA.XIR[1].XIC[2].icell.Ien VGND.t2095 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2461 VGND.t1200 Vbias.t222 XA.XIR[13].XIC[6].icell.SM VGND.t1199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2462 XA.XIR[12].XIC[7].icell.Ien XThR.Tn[12].t65 VPWR.t295 VPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2463 VGND.t420 XA.Cn[5].t36 XA.XIR[13].XIC[5].icell.PDM VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2464 VGND.t607 VPWR.t2050 XA.XIR[9].XIC_dummy_right.icell.PDM VGND.t606 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2465 XA.Cn[2].t6 thermo15c_0.XTBN.Y.t103 a_4067_9615# VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2466 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[4].t67 XA.XIR[4].XIC[3].icell.Ien VGND.t1795 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2467 VPWR.t133 XThR.Tn[8].t66 XA.XIR[9].XIC[11].icell.PUM VPWR.t132 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2468 VPWR.t5 XThR.Tn[14].t68 XA.XIR[15].XIC[3].icell.PUM VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2469 XA.XIR[7].XIC[12].icell.PUM XA.Cn[12].t38 XA.XIR[7].XIC[12].icell.Ien VPWR.t1394 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2470 VGND.t1129 XThR.XTB7.B XThR.XTB4.Y.t1 VGND.t1128 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2471 VPWR.t605 VPWR.t603 XA.XIR[10].XIC_15.icell.PUM VPWR.t604 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2472 VGND.t1202 Vbias.t223 XA.XIR[4].XIC_15.icell.SM VGND.t1201 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2473 XA.XIR[15].XIC[2].icell.Ien VPWR.t600 VPWR.t602 VPWR.t601 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2474 VGND.t1204 Vbias.t224 XA.XIR[11].XIC[13].icell.SM VGND.t1203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2475 XA.XIR[10].XIC[14].icell.Ien XThR.Tn[10].t63 VPWR.t1732 VPWR.t1731 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2476 VGND.t1416 XThR.XTB1.Y XThR.Tn[0].t0 VGND.t1415 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2477 VPWR.t1713 XThR.Tn[1].t63 XA.XIR[2].XIC[4].icell.PUM VPWR.t1712 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2478 VPWR.t1262 XThR.Tn[5].t64 XA.XIR[6].XIC[1].icell.PUM VPWR.t1261 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2479 XA.XIR[13].XIC_15.icell.Ien XThR.Tn[13].t64 VPWR.t1417 VPWR.t1416 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2480 XA.XIR[14].XIC[9].icell.SM XA.XIR[14].XIC[9].icell.Ien Iout.t137 VGND.t1073 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2481 VPWR.t135 XThR.Tn[8].t67 XA.XIR[9].XIC[2].icell.PUM VPWR.t134 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2482 XA.XIR[15].XIC[5].icell.PDM VPWR.t2051 XA.XIR[15].XIC[5].icell.Ien VGND.t608 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2483 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout VGND.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2484 VGND.t411 XA.Cn[11].t38 XA.XIR[14].XIC[11].icell.PDM VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2485 VGND.t1206 Vbias.t225 XA.XIR[2].XIC[2].icell.SM VGND.t1205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2486 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t594 VPWR.t596 VPWR.t595 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2487 XA.XIR[1].XIC[10].icell.SM XA.XIR[1].XIC[10].icell.Ien Iout.t235 VGND.t2127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2488 a_8739_9569# thermo15c_0.XTBN.Y.t104 VGND.t1285 VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2489 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[8].t68 VGND.t234 VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2490 XA.Cn[6].t8 thermo15c_0.XTB7.Y VGND.t1391 VGND.t1390 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2491 XA.XIR[3].XIC[5].icell.Ien XThR.Tn[3].t69 VPWR.t1024 VPWR.t1023 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2492 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[10].t64 VGND.t2153 VGND.t2152 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2493 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[5].t65 VGND.t1222 VGND.t1221 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2494 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[1].t64 XA.XIR[1].XIC[6].icell.Ien VGND.t2096 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2495 VGND.t1208 Vbias.t226 XA.XIR[13].XIC[10].icell.SM VGND.t1207 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2496 VGND.t1324 thermo15c_0.XTBN.Y.t105 XA.Cn[7].t4 VGND.t1323 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2497 XA.Cn[12].t8 thermo15c_0.XTBN.Y.t106 VPWR.t1310 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2498 XA.XIR[12].XIC[11].icell.Ien XThR.Tn[12].t66 VPWR.t297 VPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2499 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[4].t68 XA.XIR[4].XIC[7].icell.Ien VGND.t1796 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2500 VGND.t2085 XA.Cn[2].t38 XA.XIR[14].XIC[2].icell.PDM VGND.t2084 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2501 XA.Cn[12].t4 thermo15c_0.XTB5.Y a_9827_9569# VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2502 XA.XIR[1].XIC[1].icell.SM XA.XIR[1].XIC[1].icell.Ien Iout.t60 VGND.t213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2503 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[1].t65 VGND.t2098 VGND.t2097 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2504 XA.XIR[7].XIC[10].icell.PUM XA.Cn[10].t39 XA.XIR[7].XIC[10].icell.Ien VPWR.t1338 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2505 XA.XIR[4].XIC[12].icell.PUM XA.Cn[12].t39 XA.XIR[4].XIC[12].icell.Ien VPWR.t1395 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2506 a_8963_9569# thermo15c_0.XTB4.Y.t15 XA.Cn[11].t0 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2507 XA.XIR[0].XIC[13].icell.SM XA.XIR[0].XIC[13].icell.Ien Iout.t212 VGND.t1779 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2508 XA.XIR[3].XIC[13].icell.PUM XA.Cn[13].t39 XA.XIR[3].XIC[13].icell.Ien VPWR.t1924 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2509 VGND.t1891 Vbias.t227 XA.XIR[10].XIC[0].icell.SM VGND.t1890 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2510 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t592 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t593 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2511 VGND.t1893 Vbias.t228 XA.XIR[5].XIC[12].icell.SM VGND.t1892 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2512 VGND.t1042 XA.Cn[8].t40 XA.XIR[1].XIC[8].icell.PDM VGND.t1041 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2513 VGND.t161 XA.Cn[14].t40 XA.XIR[1].XIC[14].icell.PDM VGND.t160 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2514 XThR.Tn[13].t1 XThR.XTB6.Y VPWR.t540 VPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2515 VGND.t1895 Vbias.t229 XA.XIR[13].XIC[1].icell.SM VGND.t1894 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2516 XA.XIR[12].XIC[2].icell.Ien XThR.Tn[12].t67 VPWR.t299 VPWR.t298 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2517 VGND.t1220 XA.Cn[0].t37 XA.XIR[13].XIC[0].icell.PDM VGND.t1219 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2518 VGND.t1897 Vbias.t230 XA.XIR[8].XIC[13].icell.SM VGND.t1896 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2519 XA.XIR[7].XIC[14].icell.Ien XThR.Tn[7].t60 VPWR.t1404 VPWR.t1403 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2520 VGND.t1462 XA.Cn[12].t40 XA.XIR[8].XIC[12].icell.PDM VGND.t1461 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2521 VPWR.t1715 XThR.Tn[1].t66 XA.XIR[2].XIC[0].icell.PUM VPWR.t1714 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2522 VGND.t2656 XA.Cn[13].t40 XA.XIR[11].XIC[13].icell.PDM VGND.t2655 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2523 XA.XIR[12].XIC[7].icell.PUM XA.Cn[7].t35 XA.XIR[12].XIC[7].icell.Ien VPWR.t95 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2524 VGND.t1325 thermo15c_0.XTBN.Y.t107 a_7875_9569# VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2525 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12].t68 XA.XIR[12].XIC[5].icell.Ien VGND.t717 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2526 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2052 XA.XIR[11].XIC_dummy_left.icell.Ien VGND.t609 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2527 XA.XIR[15].XIC[8].icell.PUM XA.Cn[8].t41 XA.XIR[15].XIC[8].icell.Ien VPWR.t1096 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2528 XA.XIR[2].XIC[4].icell.Ien XThR.Tn[2].t64 VPWR.t1142 VPWR.t1141 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2529 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14].t69 XA.XIR[14].XIC_15.icell.Ien VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2530 XA.XIR[11].XIC_15.icell.SM XA.XIR[11].XIC_15.icell.Ien Iout.t246 VGND.t2493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2531 VGND.t1899 Vbias.t231 XA.XIR[7].XIC[11].icell.SM VGND.t1898 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2532 XA.XIR[6].XIC[12].icell.Ien XThR.Tn[6].t66 VPWR.t211 VPWR.t210 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2533 XA.XIR[5].XIC[13].icell.Ien XThR.Tn[5].t66 VPWR.t1264 VPWR.t1263 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2534 XA.XIR[14].XIC[4].icell.SM XA.XIR[14].XIC[4].icell.Ien Iout.t198 VGND.t1501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2535 XA.XIR[9].XIC[13].icell.Ien XThR.Tn[9].t64 VPWR.t410 VPWR.t409 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2536 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[5].t67 VGND.t1224 VGND.t1223 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2537 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout VGND.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2538 VPWR.t1456 VGND.t2700 XA.XIR[0].XIC[12].icell.PUM VPWR.t1455 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2539 XA.XIR[15].XIC[0].icell.PDM VPWR.t2053 XA.XIR[15].XIC[0].icell.Ien VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2540 a_8963_9569# thermo15c_0.XTBN.Y.t108 VGND.t1326 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2541 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10].t65 XA.XIR[10].XIC[12].icell.Ien VGND.t2154 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2542 VGND.t558 XA.Cn[6].t40 XA.XIR[14].XIC[6].icell.PDM VGND.t557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2543 XA.XIR[1].XIC[9].icell.PUM XA.Cn[9].t41 XA.XIR[1].XIC[9].icell.Ien VPWR.t1571 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2544 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[1].t67 VGND.t2100 VGND.t2099 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2545 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13].t65 XA.XIR[13].XIC[13].icell.Ien VGND.t1523 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2546 VPWR.t591 VPWR.t589 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t590 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2547 XA.XIR[4].XIC[10].icell.PUM XA.Cn[10].t40 XA.XIR[4].XIC[10].icell.Ien VPWR.t1339 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2548 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[13].t66 VGND.t1525 VGND.t1524 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2549 XA.XIR[0].XIC[8].icell.PDM XThR.Tn[0].t66 XA.XIR[0].XIC[8].icell.Ien VGND.t544 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2550 XA.XIR[0].XIC[14].icell.PDM XThR.Tn[0].t67 XA.XIR[0].XIC[14].icell.Ien VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2551 VPWR.t1406 XThR.Tn[7].t61 XA.XIR[8].XIC[7].icell.PUM VPWR.t1405 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2552 VGND.t1364 XA.Cn[10].t41 XA.XIR[8].XIC[10].icell.PDM VGND.t1363 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2553 XA.Cn[11].t3 thermo15c_0.XTBN.Y.t109 VPWR.t1311 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2554 VPWR.t1734 XThR.Tn[10].t66 XA.XIR[11].XIC[8].icell.PUM VPWR.t1733 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2555 VGND.t1901 Vbias.t232 XA.XIR[1].XIC[7].icell.SM VGND.t1900 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2556 XThR.Tn[6].t5 XThR.XTBN.Y a_n1049_5317# VPWR.t1775 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2557 XA.XIR[7].XIC[5].icell.PUM XA.Cn[5].t37 XA.XIR[7].XIC[5].icell.Ien VPWR.t345 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2558 VPWR.t156 thermo15c_0.XTB4.Y.t16 XA.Cn[11].t1 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2559 XThR.XTB7.Y XThR.XTB7.B a_n1319_5317# VPWR.t1212 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2560 XA.XIR[12].XIC[11].icell.PUM XA.Cn[11].t39 XA.XIR[12].XIC[11].icell.Ien VPWR.t334 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2561 VGND.t1903 Vbias.t233 XA.XIR[4].XIC[8].icell.SM VGND.t1902 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2562 XA.XIR[15].XIC[1].icell.PDM XThR.Tn[14].t70 VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2563 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[13].t67 VGND.t1527 VGND.t1526 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2564 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[9].t65 VGND.t487 VGND.t486 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2565 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2054 VGND.t612 VGND.t611 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2566 VGND.t1889 XA.Cn[3].t41 XA.XIR[1].XIC[3].icell.PDM VGND.t1888 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2567 VGND.t1905 Vbias.t234 XA.XIR[7].XIC[9].icell.SM VGND.t1904 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2568 XA.XIR[6].XIC[10].icell.Ien XThR.Tn[6].t67 VPWR.t213 VPWR.t212 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2569 XA.XIR[2].XIC[0].icell.Ien XThR.Tn[2].t65 VPWR.t1140 VPWR.t1139 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2570 XA.XIR[12].XIC_15.icell.PDM VPWR.t2055 VGND.t614 VGND.t613 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2571 XA.XIR[12].XIC[12].icell.SM XA.XIR[12].XIC[12].icell.Ien Iout.t46 VGND.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2572 XA.XIR[8].XIC_15.icell.SM XA.XIR[8].XIC_15.icell.Ien Iout.t234 VGND.t2126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2573 XA.XIR[15].XIC[13].icell.SM XA.XIR[15].XIC[13].icell.Ien Iout.t105 VGND.t823 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2574 VPWR.t1454 VGND.t2701 XA.XIR[0].XIC[10].icell.PUM VPWR.t1453 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2575 VPWR.t1194 thermo15c_0.XTB3.Y.t14 a_4067_9615# VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2576 XA.XIR[3].XIC[6].icell.PUM XA.Cn[6].t41 XA.XIR[3].XIC[6].icell.Ien VPWR.t469 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2577 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12].t69 XA.XIR[12].XIC[0].icell.Ien VGND.t718 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2578 XA.XIR[12].XIC[2].icell.PUM XA.Cn[2].t39 XA.XIR[12].XIC[2].icell.Ien VPWR.t1702 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2579 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10].t67 XA.XIR[10].XIC[10].icell.Ien VGND.t2155 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2580 VGND.t2380 XThR.XTBN.Y a_n997_1803# VGND.t2379 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2581 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7].t62 XA.XIR[7].XIC[12].icell.Ien VGND.t360 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2582 XA.XIR[0].XIC[9].icell.Ien XThR.Tn[0].t68 VPWR.t464 VPWR.t463 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2583 XA.XIR[15].XIC[3].icell.PUM XA.Cn[3].t42 XA.XIR[15].XIC[3].icell.Ien VPWR.t1573 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2584 XA.XIR[6].XIC[7].icell.PUM XA.Cn[7].t36 XA.XIR[6].XIC[7].icell.Ien VPWR.t96 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2585 XA.XIR[10].XIC_15.icell.PUM VPWR.t587 XA.XIR[10].XIC_15.icell.Ien VPWR.t588 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2586 a_3773_9615# thermo15c_0.XTB2.Y VPWR.t1593 VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2587 VPWR.t586 VPWR.t584 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t585 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2588 VGND.t1907 Vbias.t235 XA.XIR[12].XIC[6].icell.SM VGND.t1906 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2589 VGND.t1879 XA.Cn[9].t42 XA.XIR[3].XIC[9].icell.PDM VGND.t1878 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2590 VGND.t422 XA.Cn[5].t38 XA.XIR[12].XIC[5].icell.PDM VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2591 VPWR.t241 XThR.Tn[7].t63 XA.XIR[8].XIC[11].icell.PUM VPWR.t240 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2592 XA.XIR[2].XIC[4].icell.PUM XA.Cn[4].t41 XA.XIR[2].XIC[4].icell.Ien VPWR.t1846 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2593 VPWR.t1270 XThR.XTB4.Y.t17 XThR.Tn[11].t3 VPWR.t1238 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2594 a_n997_715# XThR.XTBN.Y VGND.t2378 VGND.t2377 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2595 VGND.t1909 Vbias.t236 XA.XIR[6].XIC[5].icell.SM VGND.t1908 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2596 VPWR.t1362 XThR.XTB1.Y a_n1049_8581# VPWR.t1361 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2597 XA.XIR[4].XIC[5].icell.PUM XA.Cn[5].t39 XA.XIR[4].XIC[5].icell.Ien VPWR.t346 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2598 XA.XIR[5].XIC[6].icell.Ien XThR.Tn[5].t68 VPWR.t1266 VPWR.t1265 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2599 XThR.Tn[14].t1 XThR.XTB7.Y VPWR.t1017 VPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2600 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[13].t68 VGND.t1529 VGND.t1528 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2601 XA.XIR[9].XIC[6].icell.Ien XThR.Tn[9].t66 VPWR.t412 VPWR.t411 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2602 VGND.t1911 Vbias.t237 XA.XIR[9].XIC[6].icell.SM VGND.t1910 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2603 VGND.t1327 thermo15c_0.XTBN.Y.t110 XA.Cn[3].t9 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2604 XA.XIR[8].XIC[7].icell.Ien XThR.Tn[8].t69 VPWR.t137 VPWR.t136 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2605 VGND.t202 XA.Cn[7].t37 XA.XIR[1].XIC[7].icell.PDM VGND.t201 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2606 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2056 VGND.t616 VGND.t615 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2607 XA.XIR[0].XIC[3].icell.PDM XThR.Tn[0].t69 XA.XIR[0].XIC[3].icell.Ien VGND.t546 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2608 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout VGND.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2609 VPWR.t243 XThR.Tn[7].t64 XA.XIR[8].XIC[2].icell.PUM VPWR.t242 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2610 XA.Cn[1].t8 thermo15c_0.XTB2.Y VGND.t1938 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2611 VPWR.t1138 XThR.Tn[2].t66 XA.XIR[3].XIC[14].icell.PUM VPWR.t1137 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2612 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5].t69 XA.XIR[5].XIC[9].icell.Ien VGND.t1225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2613 XA.XIR[11].XIC[8].icell.Ien XThR.Tn[11].t71 VPWR.t1883 VPWR.t1882 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2614 VPWR.t977 thermo15c_0.XTBN.A thermo15c_0.XTBN.Y.t0 VPWR.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2615 VPWR.t1736 XThR.Tn[10].t68 XA.XIR[11].XIC[3].icell.PUM VPWR.t1735 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2616 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9].t67 XA.XIR[9].XIC[9].icell.Ien VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2617 VPWR.t215 XThR.Tn[6].t68 XA.XIR[7].XIC[14].icell.PUM VPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2618 VGND.t1913 Vbias.t238 XA.XIR[1].XIC[2].icell.SM VGND.t1912 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2619 VPWR.t583 VPWR.t581 XA.XIR[6].XIC_15.icell.PUM VPWR.t582 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2620 VGND.t1848 Vbias.t239 XA.XIR[4].XIC[3].icell.SM VGND.t1847 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2621 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7].t65 XA.XIR[7].XIC[10].icell.Ien VGND.t361 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2622 XThR.Tn[2].t3 XThR.XTB3.Y.t16 VGND.t1141 VGND.t1140 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2623 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[9].t68 VGND.t490 VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2624 XA.XIR[6].XIC[11].icell.PUM XA.Cn[11].t40 XA.XIR[6].XIC[11].icell.Ien VPWR.t1903 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2625 XA.XIR[11].XIC[8].icell.SM XA.XIR[11].XIC[8].icell.Ien Iout.t227 VGND.t1951 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2626 VGND.t1850 Vbias.t240 XA.XIR[7].XIC[4].icell.SM VGND.t1849 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2627 XA.XIR[6].XIC[5].icell.Ien XThR.Tn[6].t69 VPWR.t217 VPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2628 VGND.t1637 VGND.t1635 XA.XIR[2].XIC_dummy_right.icell.SM VGND.t1636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2629 VGND.t1852 Vbias.t241 XA.XIR[12].XIC[10].icell.SM VGND.t1851 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2630 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[7].t66 VGND.t363 VGND.t362 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2631 a_n997_3979# XThR.XTB1.Y XThR.Tn[8].t4 VGND.t1414 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2632 XA.XIR[7].XIC[11].icell.SM XA.XIR[7].XIC[11].icell.Ien Iout.t136 VGND.t1072 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2633 a_3299_10575# thermo15c_0.XTB7.B VGND.t1097 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2634 VGND.t618 VPWR.t2057 XA.XIR[8].XIC_dummy_left.icell.PDM VGND.t617 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2635 VGND.t2376 XThR.XTBN.Y XThR.Tn[6].t8 VGND.t2375 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2636 VPWR.t1452 VGND.t2702 XA.XIR[0].XIC[5].icell.PUM VPWR.t1451 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2637 XA.XIR[3].XIC[1].icell.PUM XA.Cn[1].t41 XA.XIR[3].XIC[1].icell.Ien VPWR.t1721 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2638 XA.XIR[2].XIC[0].icell.PUM XA.Cn[0].t38 XA.XIR[2].XIC[0].icell.Ien VPWR.t1914 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2639 VPWR.t1885 XThR.Tn[11].t72 XA.XIR[12].XIC[9].icell.PUM VPWR.t1884 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2640 XA.XIR[6].XIC[2].icell.PUM XA.Cn[2].t40 XA.XIR[6].XIC[2].icell.Ien VPWR.t1703 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2641 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t578 VPWR.t580 VPWR.t579 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2642 VGND.t1854 Vbias.t242 XA.XIR[12].XIC[1].icell.SM VGND.t1853 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2643 VGND.t1856 Vbias.t243 XA.XIR[3].XIC[5].icell.SM VGND.t1855 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2644 VGND.t2632 XA.Cn[0].t39 XA.XIR[12].XIC[0].icell.PDM VGND.t2631 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2645 VGND.t2488 XA.Cn[4].t42 XA.XIR[3].XIC[4].icell.PDM VGND.t2487 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2646 VGND.t1858 Vbias.t244 XA.XIR[9].XIC[10].icell.SM VGND.t1857 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2647 XA.XIR[8].XIC[11].icell.Ien XThR.Tn[8].t70 VPWR.t139 VPWR.t138 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2648 VGND.t2136 XA.Cn[1].t42 XA.XIR[11].XIC[1].icell.PDM VGND.t2135 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2649 VGND.t1860 Vbias.t245 XA.XIR[10].XIC[14].icell.SM VGND.t1859 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2650 XA.XIR[0].XIC[7].icell.PDM XThR.Tn[0].t70 XA.XIR[0].XIC[7].icell.Ien VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2651 VGND.t424 XA.Cn[5].t40 XA.XIR[6].XIC[5].icell.PDM VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2652 VPWR.t1312 thermo15c_0.XTBN.Y.t111 XA.Cn[10].t5 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2653 VGND.t2658 XA.Cn[13].t41 XA.XIR[10].XIC[13].icell.PDM VGND.t2657 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2654 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2058 XA.XIR[10].XIC_dummy_left.icell.Ien VGND.t619 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2655 XA.XIR[0].XIC[12].icell.PUM XA.Cn[12].t41 XA.XIR[0].XIC[12].icell.Ien VPWR.t1396 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2656 VGND.t1328 thermo15c_0.XTBN.Y.t112 a_8963_9569# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2657 XA.XIR[5].XIC[1].icell.Ien XThR.Tn[5].t70 VPWR.t1268 VPWR.t1267 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2658 VGND.t1862 Vbias.t246 XA.XIR[6].XIC[0].icell.SM VGND.t1861 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2659 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[6].t70 VGND.t346 VGND.t345 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2660 VPWR.t1836 thermo15c_0.XTB5.A a_5155_10571# VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2661 VPWR.t1347 thermo15c_0.XTB7.Y XA.Cn[14].t4 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2662 XThR.Tn[1].t8 XThR.XTBN.Y VGND.t2374 VGND.t2373 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2663 XA.XIR[1].XIC[4].icell.Ien XThR.Tn[1].t68 VPWR.t1717 VPWR.t1716 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2664 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9].t69 VPWR.t414 VPWR.t413 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2665 VGND.t1864 Vbias.t247 XA.XIR[9].XIC[1].icell.SM VGND.t1863 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2666 XA.XIR[8].XIC[2].icell.Ien XThR.Tn[8].t71 VPWR.t982 VPWR.t981 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2667 XA.XIR[3].XIC[14].icell.Ien XThR.Tn[3].t70 VPWR.t1026 VPWR.t1025 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2668 XA.XIR[5].XIC[7].icell.SM XA.XIR[5].XIC[7].icell.Ien Iout.t99 VGND.t772 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2669 VPWR.t1739 thermo15c_0.XTB7.A thermo15c_0.XTB3.Y.t2 VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2670 XA.XIR[11].XIC[3].icell.Ien XThR.Tn[11].t73 VPWR.t1887 VPWR.t1886 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2671 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5].t71 XA.XIR[5].XIC[4].icell.Ien VGND.t2262 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2672 XA.XIR[8].XIC[8].icell.SM XA.XIR[8].XIC[8].icell.Ien Iout.t194 VGND.t1496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2673 XA.XIR[7].XIC[9].icell.SM XA.XIR[7].XIC[9].icell.Ien Iout.t164 VGND.t1283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2674 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13].t69 XA.XIR[13].XIC[1].icell.Ien VGND.t1871 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2675 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9].t70 XA.XIR[9].XIC[4].icell.Ien VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2676 XThR.Tn[8].t8 XThR.XTBN.Y VPWR.t1777 VPWR.t1776 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2677 VPWR.t1543 XThR.Tn[1].t69 XA.XIR[2].XIC[13].icell.PUM VPWR.t1542 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2678 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t2059 XA.XIR[4].XIC_dummy_right.icell.Ien VGND.t620 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2679 XThR.Tn[5].t4 XThR.XTBN.Y a_n1049_5611# VPWR.t1775 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2680 a_n997_2891# XThR.XTB3.Y.t17 XThR.Tn[10].t1 VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2681 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8].t72 XA.XIR[8].XIC[5].icell.Ien VGND.t840 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2682 XThR.XTB6.Y XThR.XTB7.B a_n1319_5611# VPWR.t1212 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2683 VPWR.t577 VPWR.t575 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t576 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2684 XA.XIR[2].XIC[7].icell.SM XA.XIR[2].XIC[7].icell.Ien Iout.t208 VGND.t1536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2685 XA.XIR[11].XIC[3].icell.SM XA.XIR[11].XIC[3].icell.Ien Iout.t59 VGND.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2686 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t4 VPWR.t1774 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2687 a_3773_9615# thermo15c_0.XTBN.Y.t113 XA.Cn[1].t1 VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2688 VPWR.t1211 XThR.XTB7.B XThR.XTB3.Y.t0 VPWR.t1210 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2689 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t2060 XA.XIR[7].XIC_dummy_left.icell.Ien VGND.t621 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2690 XA.XIR[0].XIC[10].icell.PUM XA.Cn[10].t42 XA.XIR[0].XIC[10].icell.Ien VPWR.t1340 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2691 a_4067_9615# thermo15c_0.XTB3.Y.t15 VPWR.t1195 VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2692 VGND.t1866 Vbias.t248 XA.XIR[3].XIC[0].icell.SM VGND.t1865 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2693 VPWR.t1718 thermo15c_0.XTB3.Y.t16 XA.Cn[10].t9 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2694 VPWR.t1313 thermo15c_0.XTBN.Y.t114 XA.Cn[14].t1 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2695 XA.XIR[1].XIC[0].icell.Ien XThR.Tn[1].t70 VPWR.t1545 VPWR.t1544 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2696 VGND.t1634 VGND.t1632 XA.XIR[2].XIC_dummy_left.icell.SM VGND.t1633 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2697 XA.XIR[14].XIC[4].icell.PUM XA.Cn[4].t43 XA.XIR[14].XIC[4].icell.Ien VPWR.t1847 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2698 XA.XIR[15].XIC_15.icell.PDM VPWR.t2061 VGND.t623 VGND.t622 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2699 XA.XIR[10].XIC[5].icell.SM XA.XIR[10].XIC[5].icell.Ien Iout.t10 VGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2700 VGND.t2634 XA.Cn[0].t40 XA.XIR[6].XIC[0].icell.PDM VGND.t2633 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2701 XA.XIR[14].XIC[13].icell.SM XA.XIR[14].XIC[13].icell.Ien Iout.t67 VGND.t539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2702 VGND.t2372 XThR.XTBN.Y XThR.Tn[0].t8 VGND.t2371 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2703 XA.XIR[13].XIC[6].icell.SM XA.XIR[13].XIC[6].icell.Ien Iout.t16 VGND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2704 VGND.t2130 thermo15c_0.XTB3.Y.t17 XA.Cn[2].t11 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2705 XA.XIR[5].XIC[7].icell.PUM XA.Cn[7].t38 XA.XIR[5].XIC[7].icell.Ien VPWR.t97 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2706 XThR.Tn[10].t8 XThR.XTBN.Y VPWR.t1773 VPWR.t1772 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2707 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[6].t71 VGND.t348 VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2708 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2062 VGND.t625 VGND.t624 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2709 XA.XIR[9].XIC[7].icell.PUM XA.Cn[7].t39 XA.XIR[9].XIC[7].icell.Ien VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2710 XA.XIR[5].XIC[2].icell.SM XA.XIR[5].XIC[2].icell.Ien Iout.t195 VGND.t1497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2711 XA.XIR[8].XIC[8].icell.PUM XA.Cn[8].t42 XA.XIR[8].XIC[8].icell.Ien VPWR.t1097 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2712 VGND.t1868 Vbias.t249 XA.XIR[0].XIC[11].icell.SM VGND.t1867 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2713 VPWR.t1031 thermo15c_0.XTB6.Y a_5949_9615# VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2714 XThR.Tn[1].t0 XThR.XTB2.Y VGND.t1999 VGND.t1420 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2715 XA.XIR[4].XIC_15.icell.SM XA.XIR[4].XIC_15.icell.Ien Iout.t44 VGND.t179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2716 VGND.t2370 XThR.XTBN.Y a_n997_3755# VGND.t2369 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2717 VPWR.t1225 data[3].t1 thermo15c_0.XTBN.A VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2718 XA.XIR[8].XIC[3].icell.SM XA.XIR[8].XIC[3].icell.Ien Iout.t204 VGND.t1507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2719 a_2979_9615# thermo15c_0.XTB1.Y.t17 VPWR.t1728 VPWR.t1727 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2720 XA.Cn[3].t8 thermo15c_0.XTBN.Y.t115 VGND.t1286 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2721 XA.XIR[2].XIC[13].icell.Ien XThR.Tn[2].t67 VPWR.t1136 VPWR.t1135 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2722 XA.XIR[7].XIC[4].icell.SM XA.XIR[7].XIC[4].icell.Ien Iout.t48 VGND.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2723 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8].t73 XA.XIR[8].XIC[0].icell.Ien VGND.t841 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2724 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[3].t71 XA.XIR[3].XIC[12].icell.Ien VGND.t894 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2725 XA.XIR[7].XIC[14].icell.PUM XA.Cn[14].t41 XA.XIR[7].XIC[14].icell.Ien VPWR.t79 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2726 VPWR.t1565 XThR.Tn[13].t70 XA.XIR[14].XIC[12].icell.PUM VPWR.t1564 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2727 XA.XIR[2].XIC[2].icell.SM XA.XIR[2].XIC[2].icell.Ien Iout.t49 VGND.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2728 XA.XIR[10].XIC[8].icell.Ien XThR.Tn[10].t69 VPWR.t1738 VPWR.t1737 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2729 a_5949_10571# thermo15c_0.XTB7.B thermo15c_0.XTB6.Y VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2730 VPWR.t1547 XThR.Tn[1].t71 XA.XIR[2].XIC[6].icell.PUM VPWR.t1546 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2731 VPWR.t309 XThR.Tn[0].t71 XA.XIR[1].XIC[7].icell.PUM VPWR.t308 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2732 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[10].t70 VGND.t2157 VGND.t2156 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2733 XA.XIR[14].XIC[0].icell.PUM XA.Cn[0].t41 XA.XIR[14].XIC[0].icell.Ien VPWR.t1915 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2734 XThR.Tn[13].t0 XThR.XTB6.Y VPWR.t538 VPWR.t537 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2735 VPWR.t1521 XThR.Tn[4].t69 XA.XIR[5].XIC[7].icell.PUM VPWR.t1520 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2736 XA.XIR[13].XIC[10].icell.SM XA.XIR[13].XIC[10].icell.Ien Iout.t152 VGND.t1153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2737 a_n1049_7493# XThR.XTB3.Y.t18 VPWR.t92 VPWR.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2738 XA.XIR[0].XIC[5].icell.PUM XA.Cn[5].t41 XA.XIR[0].XIC[5].icell.Ien VPWR.t347 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2739 XA.XIR[5].XIC[11].icell.PUM XA.Cn[11].t41 XA.XIR[5].XIC[11].icell.Ien VPWR.t1904 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2740 XA.XIR[9].XIC[11].icell.PUM XA.Cn[11].t42 XA.XIR[9].XIC[11].icell.Ien VPWR.t1905 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2741 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[7].t67 VGND.t365 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2742 VGND.t1631 VGND.t1629 XA.XIR[1].XIC_dummy_right.icell.SM VGND.t1630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2743 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[2].t68 VGND.t1563 VGND.t1562 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2744 VGND.t1870 Vbias.t250 XA.XIR[0].XIC[9].icell.SM VGND.t1869 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2745 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[10].t71 VGND.t536 VGND.t535 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2746 XA.XIR[10].XIC[0].icell.SM XA.XIR[10].XIC[0].icell.Ien Iout.t113 VGND.t877 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2747 VPWR.t1730 thermo15c_0.XTB1.Y.t18 XA.Cn[8].t0 VPWR.t1729 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2748 VGND.t2617 XA.Cn[11].t43 XA.XIR[13].XIC[11].icell.PDM VGND.t2616 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2749 XA.XIR[13].XIC[1].icell.SM XA.XIR[13].XIC[1].icell.Ien Iout.t12 VGND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2750 VGND.t1165 XThR.XTB5.Y XThR.Tn[4].t0 VGND.t745 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2751 XA.Cn[10].t4 thermo15c_0.XTBN.Y.t116 VPWR.t1297 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2752 VGND.t1288 thermo15c_0.XTBN.Y.t117 XA.Cn[6].t4 VGND.t1287 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2753 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[3].t72 XA.XIR[3].XIC[10].icell.Ien VGND.t895 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2754 XA.XIR[5].XIC[2].icell.PUM XA.Cn[2].t41 XA.XIR[5].XIC[2].icell.Ien VPWR.t1704 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2755 VPWR.t7 XThR.Tn[14].t71 XA.XIR[15].XIC[9].icell.PUM VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2756 VPWR.t1567 XThR.Tn[13].t71 XA.XIR[14].XIC[10].icell.PUM VPWR.t1566 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2757 XA.XIR[9].XIC[2].icell.PUM XA.Cn[2].t42 XA.XIR[9].XIC[2].icell.Ien VPWR.t1705 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2758 XA.XIR[4].XIC[14].icell.PUM XA.Cn[14].t42 XA.XIR[4].XIC[14].icell.Ien VPWR.t80 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2759 XA.XIR[8].XIC[3].icell.PUM XA.Cn[3].t43 XA.XIR[8].XIC[3].icell.Ien VPWR.t1574 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2760 XA.XIR[3].XIC_15.icell.PUM VPWR.t573 XA.XIR[3].XIC_15.icell.Ien VPWR.t574 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2761 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[4].t70 VGND.t1798 VGND.t1797 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2762 VGND.t1826 Vbias.t251 XA.XIR[5].XIC[6].icell.SM VGND.t1825 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2763 VGND.t2138 XA.Cn[1].t43 XA.XIR[10].XIC[1].icell.PDM VGND.t2137 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2764 VGND.t627 VPWR.t2063 XA.XIR[1].XIC_dummy_right.icell.PDM VGND.t626 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2765 VGND.t426 XA.Cn[5].t42 XA.XIR[5].XIC[5].icell.PDM VGND.t425 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2766 VGND.t2087 XA.Cn[2].t43 XA.XIR[13].XIC[2].icell.PDM VGND.t2086 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2767 VGND.t428 XA.Cn[5].t43 XA.XIR[9].XIC[5].icell.PDM VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2768 VPWR.t311 XThR.Tn[0].t72 XA.XIR[1].XIC[11].icell.PUM VPWR.t310 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2769 XA.XIR[7].XIC[8].icell.Ien XThR.Tn[7].t68 VPWR.t245 VPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2770 VPWR.t157 thermo15c_0.XTB4.Y.t17 a_4861_9615# VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2771 VPWR.t1523 XThR.Tn[4].t71 XA.XIR[5].XIC[11].icell.PUM VPWR.t1522 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2772 XA.XIR[14].XIC[12].icell.Ien XThR.Tn[14].t72 VPWR.t9 VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2773 XA.XIR[15].XIC[11].icell.PDM VPWR.t2064 XA.XIR[15].XIC[11].icell.Ien VGND.t628 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2774 VGND.t630 VPWR.t2065 XA.XIR[11].XIC_15.icell.PDM VGND.t629 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2775 XA.XIR[2].XIC[13].icell.PUM XA.Cn[13].t42 XA.XIR[2].XIC[13].icell.Ien VPWR.t1925 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2776 VGND.t1828 Vbias.t252 XA.XIR[4].XIC[12].icell.SM VGND.t1827 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2777 XThR.Tn[6].t4 XThR.XTBN.Y a_n1049_5317# VPWR.t1771 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2778 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t571 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t572 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2779 a_10915_9569# thermo15c_0.XTB7.Y XA.Cn[14].t8 VGND.t1389 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2780 XA.XIR[2].XIC[6].icell.Ien XThR.Tn[2].t69 VPWR.t1134 VPWR.t1133 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2781 XA.XIR[10].XIC[3].icell.Ien XThR.Tn[10].t72 VPWR.t452 VPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2782 VGND.t1830 Vbias.t253 XA.XIR[7].XIC[13].icell.SM VGND.t1829 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2783 XA.XIR[6].XIC[14].icell.Ien XThR.Tn[6].t72 VPWR.t219 VPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2784 VGND.t1290 thermo15c_0.XTBN.Y.t118 a_10915_9569# VGND.t1289 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2785 VPWR.t1549 XThR.Tn[1].t72 XA.XIR[2].XIC[1].icell.PUM VPWR.t1548 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2786 XA.XIR[5].XIC_15.icell.Ien XThR.Tn[5].t72 VPWR.t1763 VPWR.t1762 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2787 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[10].t73 VGND.t538 VGND.t537 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2788 VGND.t1464 XA.Cn[12].t42 XA.XIR[7].XIC[12].icell.PDM VGND.t1463 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2789 VGND.t1832 Vbias.t254 XA.XIR[6].XIC[14].icell.SM VGND.t1831 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2790 VPWR.t313 XThR.Tn[0].t73 XA.XIR[1].XIC[2].icell.PUM VPWR.t312 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2791 XA.XIR[9].XIC_15.icell.Ien XThR.Tn[9].t71 VPWR.t416 VPWR.t415 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2792 VPWR.t1525 XThR.Tn[4].t72 XA.XIR[5].XIC[2].icell.PUM VPWR.t1524 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2793 VPWR.t1450 VGND.t2703 XA.XIR[0].XIC[14].icell.PUM VPWR.t1449 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2794 XA.XIR[15].XIC[2].icell.PDM VPWR.t2066 XA.XIR[15].XIC[2].icell.Ien VGND.t631 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2795 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[2].t70 XA.XIR[2].XIC[9].icell.Ien VGND.t1567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2796 XA.Cn[1].t0 thermo15c_0.XTBN.Y.t119 a_3773_9615# VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2797 XA.XIR[1].XIC[7].icell.SM XA.XIR[1].XIC[7].icell.Ien Iout.t237 VGND.t2129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2798 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13].t72 XA.XIR[13].XIC_15.icell.Ien VGND.t1872 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2799 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[2].t71 VGND.t1566 VGND.t1565 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2800 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[4].t73 VGND.t1800 VGND.t1799 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2801 VGND.t1834 Vbias.t255 XA.XIR[0].XIC[4].icell.SM VGND.t1833 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2802 XA.XIR[4].XIC[8].icell.SM XA.XIR[4].XIC[8].icell.Ien Iout.t131 VGND.t1048 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2803 XA.Cn[14].t0 thermo15c_0.XTBN.Y.t120 VPWR.t1298 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2804 VGND.t1836 Vbias.t256 XA.XIR[5].XIC[10].icell.SM VGND.t1835 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2805 VGND.t1838 Vbias.t257 XA.XIR[13].XIC[7].icell.SM VGND.t1837 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2806 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2067 XA.XIR[0].XIC_dummy_right.icell.Ien VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2807 VGND.t560 XA.Cn[6].t42 XA.XIR[13].XIC[6].icell.PDM VGND.t559 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2808 VGND.t2368 XThR.XTBN.Y a_n997_715# VGND.t2367 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2809 VPWR.t570 VPWR.t568 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t569 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2810 XA.XIR[14].XIC[10].icell.Ien XThR.Tn[14].t73 VPWR.t11 VPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2811 VPWR.t1569 XThR.Tn[13].t73 XA.XIR[14].XIC[5].icell.PUM VPWR.t1568 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2812 VPWR.t1016 XThR.XTB7.Y XThR.Tn[14].t0 VPWR.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2813 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12].t70 XA.XIR[12].XIC[11].icell.Ien VGND.t719 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2814 VGND.t1628 VGND.t1626 XA.XIR[1].XIC_dummy_left.icell.SM VGND.t1627 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2815 VGND.t1840 Vbias.t258 XA.XIR[5].XIC[1].icell.SM VGND.t1839 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2816 XA.XIR[9].XIC[5].icell.SM XA.XIR[9].XIC[5].icell.Ien Iout.t15 VGND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2817 XThR.XTB6.A data[5].t5 VGND.t368 VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2818 XThR.Tn[0].t4 XThR.XTBN.Y a_n1049_8581# VPWR.t1770 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2819 VGND.t2636 XA.Cn[0].t42 XA.XIR[5].XIC[0].icell.PDM VGND.t2635 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2820 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[12].t71 VGND.t721 VGND.t720 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2821 a_5949_9615# thermo15c_0.XTB6.Y VPWR.t1030 VPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2822 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[12].t72 VGND.t723 VGND.t722 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2823 XA.XIR[12].XIC[6].icell.SM XA.XIR[12].XIC[6].icell.Ien Iout.t193 VGND.t1471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2824 VGND.t2638 XA.Cn[0].t43 XA.XIR[9].XIC[0].icell.PDM VGND.t2637 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2825 VGND.t2521 XA.Cn[10].t43 XA.XIR[7].XIC[10].icell.PDM VGND.t2520 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2826 XA.XIR[7].XIC[3].icell.Ien XThR.Tn[7].t69 VPWR.t169 VPWR.t168 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2827 VGND.t1291 thermo15c_0.XTBN.Y.t121 a_10051_9569# VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2828 VGND.t1842 Vbias.t259 XA.XIR[3].XIC[14].icell.SM VGND.t1841 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2829 VGND.t1466 XA.Cn[12].t43 XA.XIR[4].XIC[12].icell.PDM VGND.t1465 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2830 VGND.t2660 XA.Cn[13].t43 XA.XIR[3].XIC[13].icell.PDM VGND.t2659 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2831 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2068 XA.XIR[3].XIC_dummy_left.icell.Ien VGND.t633 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2832 XA.XIR[15].XIC[6].icell.PDM VPWR.t2069 XA.XIR[15].XIC[6].icell.Ien VGND.t634 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2833 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12].t73 XA.XIR[12].XIC[2].icell.Ien VGND.t724 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2834 XA.XIR[0].XIC[9].icell.PDM VGND.t1623 VGND.t1625 VGND.t1624 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2835 VPWR.t1299 thermo15c_0.XTBN.Y.t122 XA.Cn[11].t2 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2836 VGND.t1292 thermo15c_0.XTBN.Y.t123 a_7651_9569# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2837 XA.XIR[2].XIC[1].icell.Ien XThR.Tn[2].t72 VPWR.t1132 VPWR.t1131 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2838 Vbias.t2 bias[1].t0 VPWR.t1095 VPWR.t1094 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
X2839 XA.XIR[11].XIC[12].icell.SM XA.XIR[11].XIC[12].icell.Ien Iout.t50 VGND.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2840 XA.XIR[1].XIC[13].icell.Ien XThR.Tn[1].t73 VPWR.t1551 VPWR.t1550 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2841 XThR.Tn[2].t8 XThR.XTBN.Y VGND.t2366 VGND.t2365 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2842 VPWR.t1015 XThR.XTB7.Y a_n1049_5317# VPWR.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2843 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout VGND.t2685 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2844 VGND.t1844 Vbias.t260 XA.XIR[15].XIC_15.icell.SM VGND.t1843 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2845 a_8739_9569# thermo15c_0.XTB3.Y.t18 XA.Cn[10].t10 VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2846 XA.XIR[2].XIC[6].icell.PUM XA.Cn[6].t43 XA.XIR[2].XIC[6].icell.Ien VPWR.t470 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2847 VGND.t163 XA.Cn[14].t43 XA.XIR[15].XIC[14].icell.PDM VGND.t162 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2848 VGND.t1044 XA.Cn[8].t43 XA.XIR[15].XIC[8].icell.PDM VGND.t1043 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2849 VPWR.t1769 XThR.XTBN.Y XThR.Tn[12].t8 VPWR.t1768 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2850 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[2].t73 XA.XIR[2].XIC[4].icell.Ien VGND.t1564 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2851 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6].t73 XA.XIR[6].XIC[12].icell.Ien VGND.t349 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2852 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5].t73 XA.XIR[5].XIC[13].icell.Ien VGND.t2263 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2853 XA.XIR[1].XIC[2].icell.SM XA.XIR[1].XIC[2].icell.Ien Iout.t69 VGND.t549 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2854 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9].t72 XA.XIR[9].XIC[13].icell.Ien VGND.t492 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2855 VPWR.t567 VPWR.t565 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t566 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2856 VGND.t1881 XA.Cn[9].t43 XA.XIR[2].XIC[9].icell.PDM VGND.t1880 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2857 XA.XIR[4].XIC[3].icell.SM XA.XIR[4].XIC[3].icell.Ien Iout.t184 VGND.t1403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2858 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[9].t73 VGND.t494 VGND.t493 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2859 VGND.t1846 Vbias.t261 XA.XIR[13].XIC[2].icell.SM VGND.t1845 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2860 VPWR.t1028 XThR.Tn[3].t73 XA.XIR[4].XIC[7].icell.PUM VPWR.t1027 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
R0 VGND.n3019 VGND.n3018 15660.6
R1 VGND.n196 VGND.n195 13477
R2 VGND.n3018 VGND.n7 11578
R3 VGND.n195 VGND.n7 10429.6
R4 VGND.n3012 VGND.n8 9309.26
R5 VGND.n200 VGND.n199 9223.7
R6 VGND.n198 VGND.n197 9223.7
R7 VGND.n197 VGND.n196 9223.7
R8 VGND.n2969 VGND.n200 9223.7
R9 VGND.n2969 VGND.n2968 7447.41
R10 VGND.n2249 VGND.n2248 7387.65
R11 VGND.n2250 VGND.n2249 7387.65
R12 VGND.n2285 VGND.n2284 7387.65
R13 VGND.n3017 VGND.n3016 7387.65
R14 VGND.n3016 VGND.n3015 7387.65
R15 VGND.n3015 VGND.n3014 7387.65
R16 VGND.n3014 VGND.n3013 7387.65
R17 VGND.n3013 VGND.n3012 7387.65
R18 VGND.n2351 VGND.n2285 6674.35
R19 VGND.n1386 VGND.t685 6324.96
R20 VGND.n199 VGND.n198 5231.11
R21 VGND.n1336 VGND.t2323 5168.13
R22 VGND.n2967 VGND.n8 5074.71
R23 VGND.n3018 VGND.n3017 5063.19
R24 VGND.n1154 VGND.n806 4539.15
R25 VGND VGND.n8 4240.58
R26 VGND.t1627 VGND.t1146 4212.19
R27 VGND.t1633 VGND.t1116 4212.19
R28 VGND.t1639 VGND.t1282 4212.19
R29 VGND.t1726 VGND.t1085 4212.19
R30 VGND.t1732 VGND.t1161 4212.19
R31 VGND.t1645 VGND.t1117 4212.19
R32 VGND.t1687 VGND.t2630 4212.19
R33 VGND.t1045 VGND.t1738 4212.19
R34 VGND.t151 VGND.t1660 4212.19
R35 VGND.t152 VGND.t1705 4212.19
R36 VGND.t1521 VGND.t1744 4212.19
R37 VGND.t1047 VGND.t1756 4212.19
R38 VGND.t668 VGND.t1672 4212.19
R39 VGND.t2476 VGND.t1714 4212.19
R40 VGND.n2919 VGND.n222 4077.12
R41 VGND.n1340 VGND.n1338 3417.39
R42 VGND.n1340 VGND.n1339 3417.39
R43 VGND.n1388 VGND.n1387 3417.39
R44 VGND.n2180 VGND.n504 3417.39
R45 VGND.n503 VGND.n473 3417.39
R46 VGND.n2353 VGND.n2352 3417.39
R47 VGND.n2920 VGND.n2919 3331.79
R48 VGND.n2921 VGND.n2920 3331.79
R49 VGND.n2922 VGND.n2921 3331.79
R50 VGND.n2923 VGND.n2922 3331.79
R51 VGND.n2924 VGND.n2923 3331.79
R52 VGND.n2925 VGND.n2924 3331.79
R53 VGND.n2926 VGND.n2925 3331.79
R54 VGND.n2927 VGND.n2926 3331.79
R55 VGND.n2928 VGND.n2927 3331.79
R56 VGND.n2929 VGND.n2928 3331.79
R57 VGND.n2930 VGND.n2929 3331.79
R58 VGND.n2931 VGND.n2930 3331.79
R59 VGND.n2932 VGND.n2931 3331.79
R60 VGND.n2933 VGND.n2932 3331.79
R61 VGND.n2934 VGND.n2933 3331.79
R62 VGND.n1339 VGND.n806 3273.91
R63 VGND.n2181 VGND.n539 3265.22
R64 VGND.n2934 VGND.n201 2725.63
R65 VGND.n197 VGND.t2442 2655.17
R66 VGND.n196 VGND.t2418 2655.17
R67 VGND.n2353 VGND.n2285 2517.39
R68 VGND.t1026 VGND.n201 2334.15
R69 VGND.t574 VGND.n2701 2307.69
R70 VGND.n359 VGND.t2283 2307.69
R71 VGND.n360 VGND.t2270 2307.69
R72 VGND.n370 VGND.t633 2307.69
R73 VGND.n371 VGND.t2349 2307.69
R74 VGND.n381 VGND.t2247 2307.69
R75 VGND.n382 VGND.t2178 2307.69
R76 VGND.t621 VGND.n327 2307.69
R77 VGND.n2705 VGND.t2319 2307.69
R78 VGND.n2728 VGND.t2248 2307.69
R79 VGND.n2738 VGND.t619 2307.69
R80 VGND.t609 VGND.n2737 2307.69
R81 VGND.n2731 VGND.t2310 2307.69
R82 VGND.n2776 VGND.t2217 2307.69
R83 VGND.t2194 VGND.n2775 2307.69
R84 VGND.n2943 VGND.t2307 2307.69
R85 VGND.t1678 VGND.n2703 2280.49
R86 VGND.n3020 VGND.n5 2229.43
R87 VGND.n3020 VGND.n6 2229.43
R88 VGND.n2348 VGND.n6 2229.43
R89 VGND.n2348 VGND.n5 2229.43
R90 VGND.n1338 VGND.n1337 2173.91
R91 VGND.n2704 VGND.t101 2132.93
R92 VGND.n2701 VGND.t2181 2123.08
R93 VGND.t2351 VGND.n359 2123.08
R94 VGND.n360 VGND.t2329 2123.08
R95 VGND.t2179 VGND.n370 2123.08
R96 VGND.n371 VGND.t2168 2123.08
R97 VGND.t615 VGND.n381 2123.08
R98 VGND.n382 VGND.t2249 2123.08
R99 VGND.n2705 VGND.t611 2123.08
R100 VGND.t2313 VGND.n2728 2123.08
R101 VGND.n2738 VGND.t2301 2123.08
R102 VGND.n2737 VGND.t2197 2123.08
R103 VGND.n2731 VGND.t598 2123.08
R104 VGND.n2776 VGND.t2289 2123.08
R105 VGND.n2775 VGND.t2211 2123.08
R106 VGND.n2704 VGND.t1702 2079.27
R107 VGND.t1146 VGND.t1678 2012.2
R108 VGND.t1116 VGND.t1627 2012.2
R109 VGND.t1282 VGND.t1633 2012.2
R110 VGND.t1085 VGND.t1639 2012.2
R111 VGND.t1161 VGND.t1726 2012.2
R112 VGND.t1117 VGND.t1732 2012.2
R113 VGND.t2630 VGND.t1645 2012.2
R114 VGND.t101 VGND.t1687 2012.2
R115 VGND.t1702 VGND.t1045 2012.2
R116 VGND.t1738 VGND.t151 2012.2
R117 VGND.t1660 VGND.t152 2012.2
R118 VGND.t1705 VGND.t1521 2012.2
R119 VGND.t1744 VGND.t1047 2012.2
R120 VGND.t1756 VGND.t668 2012.2
R121 VGND.t1672 VGND.t2476 2012.2
R122 VGND.t1714 VGND.t1026 2012.2
R123 VGND.n199 VGND 1997.7
R124 VGND.n200 VGND 1997.7
R125 VGND VGND.n2969 1997.7
R126 VGND.n2968 VGND.n2944 1907.51
R127 VGND.n2284 VGND.n2251 1831.57
R128 VGND.n198 VGND.t2375 1807.04
R129 VGND.n2970 VGND.t2004 1785.51
R130 VGND.n2352 VGND.n2351 1760.87
R131 VGND.n2702 VGND.t2271 1738.46
R132 VGND.n2250 VGND.n504 1691.3
R133 VGND.n2351 VGND.n2350 1656.52
R134 VGND.t1425 VGND.n66 1618.39
R135 VGND.n3011 VGND.t1226 1618.39
R136 VGND.n2971 VGND.t750 1618.39
R137 VGND.n2702 VGND.n7 1604.17
R138 VGND.n2350 VGND.n328 1517.39
R139 VGND.n195 VGND.t2391 1517.24
R140 VGND.n2248 VGND.n540 1513.49
R141 VGND.t2226 VGND.n2704 1507.69
R142 VGND.n2703 VGND.n2702 1441.28
R143 VGND.n1386 VGND.n540 1370.36
R144 VGND.t2271 VGND.t2183 1353.85
R145 VGND.t2183 VGND.t574 1353.85
R146 VGND.t2353 VGND.t2181 1353.85
R147 VGND.t2283 VGND.t2353 1353.85
R148 VGND.t2275 VGND.t2351 1353.85
R149 VGND.t2270 VGND.t2275 1353.85
R150 VGND.t2329 VGND.t2245 1353.85
R151 VGND.t2245 VGND.t633 1353.85
R152 VGND.t2176 VGND.t2179 1353.85
R153 VGND.t2349 VGND.t2176 1353.85
R154 VGND.t2168 VGND.t2331 1353.85
R155 VGND.t2331 VGND.t2247 1353.85
R156 VGND.t2317 VGND.t615 1353.85
R157 VGND.t2178 VGND.t2317 1353.85
R158 VGND.t2249 VGND.t2172 1353.85
R159 VGND.t2172 VGND.t621 1353.85
R160 VGND.t617 VGND.t2226 1353.85
R161 VGND.t2319 VGND.t617 1353.85
R162 VGND.t611 VGND.t2333 1353.85
R163 VGND.t2333 VGND.t2248 1353.85
R164 VGND.t2228 VGND.t2313 1353.85
R165 VGND.t619 VGND.t2228 1353.85
R166 VGND.t2301 VGND.t2213 1353.85
R167 VGND.t2213 VGND.t609 1353.85
R168 VGND.t2315 VGND.t2197 1353.85
R169 VGND.t2310 VGND.t2315 1353.85
R170 VGND.t598 VGND.t2303 1353.85
R171 VGND.t2303 VGND.t2217 1353.85
R172 VGND.t2289 VGND.t2287 1353.85
R173 VGND.t2287 VGND.t2194 1353.85
R174 VGND.t2211 VGND.t602 1353.85
R175 VGND.t602 VGND.t2307 1353.85
R176 VGND.n2944 VGND.n201 1301.35
R177 VGND.n2703 VGND.n328 1278.26
R178 VGND.t1624 VGND.n540 1270.28
R179 VGND.n1127 VGND.t64 1268.93
R180 VGND.n1127 VGND.t412 1268.93
R181 VGND.n502 VGND.t391 1253.59
R182 VGND.t70 VGND.n502 1253.59
R183 VGND.n2283 VGND.t72 1253.59
R184 VGND.t872 VGND.n2283 1253.59
R185 VGND.n538 VGND.t440 1253.59
R186 VGND.t68 VGND.n538 1253.59
R187 VGND.n2247 VGND.t78 1253.59
R188 VGND.t66 VGND.n2247 1253.59
R189 VGND.n1385 VGND.t6 1253.59
R190 VGND.t495 VGND.n1385 1253.59
R191 VGND.n1337 VGND.n1336 1243.48
R192 VGND.n2251 VGND.t1669 1237.71
R193 VGND.n66 VGND.t541 1213.79
R194 VGND.n2967 VGND.n2966 1198.25
R195 VGND.n1155 VGND.n1154 1198.25
R196 VGND.n2943 VGND.n2942 1180.79
R197 VGND.n2936 VGND.n2935 1180.79
R198 VGND.n2534 VGND.n208 1180.79
R199 VGND.n2529 VGND.n209 1180.79
R200 VGND.n2817 VGND.n210 1180.79
R201 VGND.n1989 VGND.n211 1180.79
R202 VGND.n1996 VGND.n212 1180.79
R203 VGND.n2842 VGND.n213 1180.79
R204 VGND.n1829 VGND.n214 1180.79
R205 VGND.n1836 VGND.n215 1180.79
R206 VGND.n2867 VGND.n216 1180.79
R207 VGND.n1655 VGND.n217 1180.79
R208 VGND.n1650 VGND.n218 1180.79
R209 VGND.n2892 VGND.n219 1180.79
R210 VGND.n1607 VGND.n220 1180.79
R211 VGND.n2912 VGND.n221 1180.79
R212 VGND.n1282 VGND.n222 1180.79
R213 VGND.n2918 VGND.n2917 1180.79
R214 VGND.n1335 VGND.n1334 1180.46
R215 VGND.n929 VGND.n890 1180.46
R216 VGND.n934 VGND.n933 1180.46
R217 VGND.n939 VGND.n938 1180.46
R218 VGND.n944 VGND.n943 1180.46
R219 VGND.n949 VGND.n948 1180.46
R220 VGND.n954 VGND.n953 1180.46
R221 VGND.n959 VGND.n958 1180.46
R222 VGND.n964 VGND.n963 1180.46
R223 VGND.n969 VGND.n968 1180.46
R224 VGND.n974 VGND.n973 1180.46
R225 VGND.n979 VGND.n978 1180.46
R226 VGND.n984 VGND.n983 1180.46
R227 VGND.n989 VGND.n988 1180.46
R228 VGND.n991 VGND.n990 1180.46
R229 VGND.n1279 VGND.n1278 1180.46
R230 VGND.n1277 VGND.n1276 1180.46
R231 VGND.n1234 VGND.n1233 1180.46
R232 VGND.n1239 VGND.n1238 1180.46
R233 VGND.n1241 VGND.n1240 1180.46
R234 VGND.n1246 VGND.n1245 1180.46
R235 VGND.n1248 VGND.n1247 1180.46
R236 VGND.n1220 VGND.n1219 1180.46
R237 VGND.n1209 VGND.n1208 1180.46
R238 VGND.n1207 VGND.n1206 1180.46
R239 VGND.n1190 VGND.n1189 1180.46
R240 VGND.n1188 VGND.n1187 1180.46
R241 VGND.n1177 VGND.n1176 1180.46
R242 VGND.n1175 VGND.n1174 1180.46
R243 VGND.n1167 VGND.n1166 1180.46
R244 VGND.n2775 VGND.n2774 1180.46
R245 VGND.n2777 VGND.n2776 1180.46
R246 VGND.n2732 VGND.n2731 1180.46
R247 VGND.n2737 VGND.n2736 1180.46
R248 VGND.n2739 VGND.n2738 1180.46
R249 VGND.n2728 VGND.n2727 1180.46
R250 VGND.n2706 VGND.n2705 1180.46
R251 VGND.n388 VGND.n327 1180.46
R252 VGND.n383 VGND.n382 1180.46
R253 VGND.n381 VGND.n380 1180.46
R254 VGND.n372 VGND.n371 1180.46
R255 VGND.n370 VGND.n369 1180.46
R256 VGND.n361 VGND.n360 1180.46
R257 VGND.n359 VGND.n333 1180.46
R258 VGND.n2701 VGND.n2700 1180.46
R259 VGND.n2641 VGND.n2640 1180.46
R260 VGND.n2646 VGND.n2645 1180.46
R261 VGND.n2651 VGND.n2650 1180.46
R262 VGND.n2656 VGND.n2655 1180.46
R263 VGND.n2661 VGND.n2660 1180.46
R264 VGND.n2666 VGND.n2665 1180.46
R265 VGND.n2671 VGND.n2670 1180.46
R266 VGND.n2673 VGND.n2672 1180.46
R267 VGND.n2717 VGND.n2716 1180.46
R268 VGND.n2719 VGND.n2718 1180.46
R269 VGND.n2750 VGND.n2749 1180.46
R270 VGND.n2757 VGND.n2756 1180.46
R271 VGND.n2755 VGND.n2754 1180.46
R272 VGND.n2790 VGND.n2789 1180.46
R273 VGND.n2792 VGND.n2791 1180.46
R274 VGND.n2345 VGND.n2344 1180.46
R275 VGND.n2340 VGND.n2339 1180.46
R276 VGND.n2335 VGND.n2334 1180.46
R277 VGND.n2330 VGND.n2329 1180.46
R278 VGND.n2325 VGND.n2324 1180.46
R279 VGND.n2320 VGND.n2319 1180.46
R280 VGND.n2315 VGND.n2314 1180.46
R281 VGND.n2310 VGND.n2309 1180.46
R282 VGND.n2305 VGND.n2304 1180.46
R283 VGND.n2300 VGND.n2299 1180.46
R284 VGND.n2295 VGND.n2294 1180.46
R285 VGND.n2290 VGND.n2289 1180.46
R286 VGND.n2545 VGND.n2544 1180.46
R287 VGND.n2543 VGND.n2542 1180.46
R288 VGND.n2538 VGND.n2537 1180.46
R289 VGND.n2355 VGND.n2354 1180.46
R290 VGND.n2379 VGND.n2378 1180.46
R291 VGND.n2381 VGND.n2380 1180.46
R292 VGND.n2405 VGND.n2404 1180.46
R293 VGND.n2407 VGND.n2406 1180.46
R294 VGND.n2431 VGND.n2430 1180.46
R295 VGND.n2433 VGND.n2432 1180.46
R296 VGND.n2457 VGND.n2456 1180.46
R297 VGND.n2459 VGND.n2458 1180.46
R298 VGND.n2483 VGND.n2482 1180.46
R299 VGND.n2485 VGND.n2484 1180.46
R300 VGND.n2514 VGND.n2513 1180.46
R301 VGND.n2519 VGND.n2518 1180.46
R302 VGND.n2524 VGND.n2523 1180.46
R303 VGND.n2526 VGND.n2525 1180.46
R304 VGND.n2366 VGND.n2365 1180.46
R305 VGND.n2368 VGND.n2367 1180.46
R306 VGND.n2392 VGND.n2391 1180.46
R307 VGND.n2394 VGND.n2393 1180.46
R308 VGND.n2418 VGND.n2417 1180.46
R309 VGND.n2420 VGND.n2419 1180.46
R310 VGND.n2444 VGND.n2443 1180.46
R311 VGND.n2446 VGND.n2445 1180.46
R312 VGND.n2470 VGND.n2469 1180.46
R313 VGND.n2472 VGND.n2471 1180.46
R314 VGND.n2496 VGND.n2495 1180.46
R315 VGND.n2503 VGND.n2502 1180.46
R316 VGND.n2501 VGND.n2500 1180.46
R317 VGND.n2812 VGND.n2811 1180.46
R318 VGND.n2814 VGND.n2813 1180.46
R319 VGND.n1913 VGND.n1912 1180.46
R320 VGND.n1915 VGND.n1914 1180.46
R321 VGND.n1924 VGND.n1923 1180.46
R322 VGND.n1926 VGND.n1925 1180.46
R323 VGND.n1935 VGND.n1934 1180.46
R324 VGND.n1937 VGND.n1936 1180.46
R325 VGND.n1946 VGND.n1945 1180.46
R326 VGND.n1948 VGND.n1947 1180.46
R327 VGND.n1957 VGND.n1956 1180.46
R328 VGND.n1959 VGND.n1958 1180.46
R329 VGND.n1968 VGND.n1967 1180.46
R330 VGND.n1970 VGND.n1969 1180.46
R331 VGND.n1979 VGND.n1978 1180.46
R332 VGND.n1984 VGND.n1983 1180.46
R333 VGND.n1986 VGND.n1985 1180.46
R334 VGND.n599 VGND.n598 1180.46
R335 VGND.n2060 VGND.n2059 1180.46
R336 VGND.n2058 VGND.n2057 1180.46
R337 VGND.n2053 VGND.n2052 1180.46
R338 VGND.n2048 VGND.n2047 1180.46
R339 VGND.n2043 VGND.n2042 1180.46
R340 VGND.n2038 VGND.n2037 1180.46
R341 VGND.n2033 VGND.n2032 1180.46
R342 VGND.n2028 VGND.n2027 1180.46
R343 VGND.n2023 VGND.n2022 1180.46
R344 VGND.n2018 VGND.n2017 1180.46
R345 VGND.n2013 VGND.n2012 1180.46
R346 VGND.n2008 VGND.n2007 1180.46
R347 VGND.n2003 VGND.n2002 1180.46
R348 VGND.n602 VGND.n601 1180.46
R349 VGND.n2072 VGND.n2071 1180.46
R350 VGND.n2077 VGND.n2076 1180.46
R351 VGND.n2082 VGND.n2081 1180.46
R352 VGND.n2087 VGND.n2086 1180.46
R353 VGND.n2092 VGND.n2091 1180.46
R354 VGND.n2097 VGND.n2096 1180.46
R355 VGND.n2102 VGND.n2101 1180.46
R356 VGND.n2107 VGND.n2106 1180.46
R357 VGND.n2112 VGND.n2111 1180.46
R358 VGND.n2117 VGND.n2116 1180.46
R359 VGND.n2122 VGND.n2121 1180.46
R360 VGND.n2129 VGND.n2128 1180.46
R361 VGND.n2127 VGND.n2126 1180.46
R362 VGND.n2837 VGND.n2836 1180.46
R363 VGND.n2839 VGND.n2838 1180.46
R364 VGND.n2179 VGND.n2178 1180.46
R365 VGND.n1754 VGND.n550 1180.46
R366 VGND.n1764 VGND.n1763 1180.46
R367 VGND.n1766 VGND.n1765 1180.46
R368 VGND.n1775 VGND.n1774 1180.46
R369 VGND.n1777 VGND.n1776 1180.46
R370 VGND.n1786 VGND.n1785 1180.46
R371 VGND.n1788 VGND.n1787 1180.46
R372 VGND.n1797 VGND.n1796 1180.46
R373 VGND.n1799 VGND.n1798 1180.46
R374 VGND.n1808 VGND.n1807 1180.46
R375 VGND.n1810 VGND.n1809 1180.46
R376 VGND.n1819 VGND.n1818 1180.46
R377 VGND.n1824 VGND.n1823 1180.46
R378 VGND.n1826 VGND.n1825 1180.46
R379 VGND.n1681 VGND.n1680 1180.46
R380 VGND.n1683 VGND.n1682 1180.46
R381 VGND.n1692 VGND.n1691 1180.46
R382 VGND.n1697 VGND.n1696 1180.46
R383 VGND.n1702 VGND.n1701 1180.46
R384 VGND.n1707 VGND.n1706 1180.46
R385 VGND.n1712 VGND.n1711 1180.46
R386 VGND.n1717 VGND.n1716 1180.46
R387 VGND.n1722 VGND.n1721 1180.46
R388 VGND.n1727 VGND.n1726 1180.46
R389 VGND.n1732 VGND.n1731 1180.46
R390 VGND.n1850 VGND.n1849 1180.46
R391 VGND.n1848 VGND.n1847 1180.46
R392 VGND.n1843 VGND.n1842 1180.46
R393 VGND.n1735 VGND.n1734 1180.46
R394 VGND.n672 VGND.n671 1180.46
R395 VGND.n677 VGND.n676 1180.46
R396 VGND.n682 VGND.n681 1180.46
R397 VGND.n687 VGND.n686 1180.46
R398 VGND.n692 VGND.n691 1180.46
R399 VGND.n697 VGND.n696 1180.46
R400 VGND.n702 VGND.n701 1180.46
R401 VGND.n707 VGND.n706 1180.46
R402 VGND.n712 VGND.n711 1180.46
R403 VGND.n717 VGND.n716 1180.46
R404 VGND.n722 VGND.n721 1180.46
R405 VGND.n729 VGND.n728 1180.46
R406 VGND.n727 VGND.n726 1180.46
R407 VGND.n2862 VGND.n2861 1180.46
R408 VGND.n2864 VGND.n2863 1180.46
R409 VGND.n1355 VGND.n1354 1180.46
R410 VGND.n877 VGND.n876 1180.46
R411 VGND.n872 VGND.n871 1180.46
R412 VGND.n821 VGND.n808 1180.46
R413 VGND.n826 VGND.n825 1180.46
R414 VGND.n831 VGND.n830 1180.46
R415 VGND.n836 VGND.n835 1180.46
R416 VGND.n841 VGND.n840 1180.46
R417 VGND.n846 VGND.n845 1180.46
R418 VGND.n851 VGND.n850 1180.46
R419 VGND.n858 VGND.n857 1180.46
R420 VGND.n856 VGND.n855 1180.46
R421 VGND.n1666 VGND.n1665 1180.46
R422 VGND.n1664 VGND.n1663 1180.46
R423 VGND.n1659 VGND.n1658 1180.46
R424 VGND.n1393 VGND.n1392 1180.46
R425 VGND.n1398 VGND.n1397 1180.46
R426 VGND.n1400 VGND.n1399 1180.46
R427 VGND.n1493 VGND.n1492 1180.46
R428 VGND.n1495 VGND.n1494 1180.46
R429 VGND.n1519 VGND.n1518 1180.46
R430 VGND.n1521 VGND.n1520 1180.46
R431 VGND.n1545 VGND.n1544 1180.46
R432 VGND.n1550 VGND.n1549 1180.46
R433 VGND.n1557 VGND.n1556 1180.46
R434 VGND.n1555 VGND.n1554 1180.46
R435 VGND.n1635 VGND.n1634 1180.46
R436 VGND.n1640 VGND.n1639 1180.46
R437 VGND.n1645 VGND.n1644 1180.46
R438 VGND.n1647 VGND.n1646 1180.46
R439 VGND.n1413 VGND.n1412 1180.46
R440 VGND.n1415 VGND.n1414 1180.46
R441 VGND.n1480 VGND.n1479 1180.46
R442 VGND.n1482 VGND.n1481 1180.46
R443 VGND.n1506 VGND.n1505 1180.46
R444 VGND.n1508 VGND.n1507 1180.46
R445 VGND.n1532 VGND.n1531 1180.46
R446 VGND.n1534 VGND.n1533 1180.46
R447 VGND.n1569 VGND.n1568 1180.46
R448 VGND.n1586 VGND.n1585 1180.46
R449 VGND.n1584 VGND.n1583 1180.46
R450 VGND.n1579 VGND.n1578 1180.46
R451 VGND.n1574 VGND.n1573 1180.46
R452 VGND.n2887 VGND.n2886 1180.46
R453 VGND.n2889 VGND.n2888 1180.46
R454 VGND.n1342 VGND.n1341 1180.46
R455 VGND.n1426 VGND.n1425 1180.46
R456 VGND.n1431 VGND.n1430 1180.46
R457 VGND.n1436 VGND.n1435 1180.46
R458 VGND.n1441 VGND.n1440 1180.46
R459 VGND.n1446 VGND.n1445 1180.46
R460 VGND.n1451 VGND.n1450 1180.46
R461 VGND.n1456 VGND.n1455 1180.46
R462 VGND.n1463 VGND.n1462 1180.46
R463 VGND.n1461 VGND.n1460 1180.46
R464 VGND.n1598 VGND.n1597 1180.46
R465 VGND.n1603 VGND.n1602 1180.46
R466 VGND.n1618 VGND.n1617 1180.46
R467 VGND.n1616 VGND.n1615 1180.46
R468 VGND.n1611 VGND.n1610 1180.46
R469 VGND.n1034 VGND.n1033 1180.46
R470 VGND.n1039 VGND.n1038 1180.46
R471 VGND.n1099 VGND.n1098 1180.46
R472 VGND.n1097 VGND.n1096 1180.46
R473 VGND.n1092 VGND.n1091 1180.46
R474 VGND.n1087 VGND.n1086 1180.46
R475 VGND.n1082 VGND.n1081 1180.46
R476 VGND.n1077 VGND.n1076 1180.46
R477 VGND.n1072 VGND.n1071 1180.46
R478 VGND.n1050 VGND.n1041 1180.46
R479 VGND.n1055 VGND.n1054 1180.46
R480 VGND.n1060 VGND.n1059 1180.46
R481 VGND.n1062 VGND.n1061 1180.46
R482 VGND.n2907 VGND.n2906 1180.46
R483 VGND.n2909 VGND.n2908 1180.46
R484 VGND.t540 VGND.n3011 1180.08
R485 VGND.n1387 VGND.n1386 1169.57
R486 VGND.n3015 VGND.t19 1146.36
R487 VGND.n3017 VGND.t18 1112.64
R488 VGND.n3016 VGND.t1453 1112.64
R489 VGND.n2351 VGND.n2349 1070.21
R490 VGND.n2968 VGND 1055.35
R491 VGND.n2251 VGND.n2250 1052.29
R492 VGND.t1340 VGND.n2181 1032.59
R493 VGND.t141 VGND.n2641 988.926
R494 VGND.t1813 VGND.n2646 988.926
R495 VGND.t1565 VGND.n2651 988.926
R496 VGND.t923 VGND.n2656 988.926
R497 VGND.t1949 VGND.n2661 988.926
R498 VGND.t1261 VGND.n2666 988.926
R499 VGND.t2038 VGND.n2671 988.926
R500 VGND.n2672 VGND.t782 988.926
R501 VGND.t1068 VGND.n2717 988.926
R502 VGND.n2718 VGND.t489 988.926
R503 VGND.t2152 VGND.n2750 988.926
R504 VGND.n2756 VGND.t678 988.926
R505 VGND.n2755 VGND.t307 988.926
R506 VGND.t1534 VGND.n2790 988.926
R507 VGND.n2791 VGND.t475 988.926
R508 VGND.n2345 VGND.t186 988.926
R509 VGND.n2340 VGND.t228 988.926
R510 VGND.n2335 VGND.t1568 988.926
R511 VGND.n2330 VGND.t293 988.926
R512 VGND.n2325 VGND.t1319 988.926
R513 VGND.n2320 VGND.t1233 988.926
R514 VGND.n2315 VGND.t350 988.926
R515 VGND.n2310 VGND.t364 988.926
R516 VGND.n2305 VGND.t769 988.926
R517 VGND.n2300 VGND.t532 988.926
R518 VGND.n2295 VGND.t1094 988.926
R519 VGND.n2290 VGND.t2613 988.926
R520 VGND.n2544 VGND.t121 988.926
R521 VGND.n2543 VGND.t1921 988.926
R522 VGND.n2538 VGND.t12 988.926
R523 VGND.n2354 VGND.t760 988.926
R524 VGND.t702 VGND.n2379 988.926
R525 VGND.n2380 VGND.t2469 988.926
R526 VGND.t930 VGND.n2405 988.926
R527 VGND.n2406 VGND.t2077 988.926
R528 VGND.t1267 VGND.n2431 988.926
R529 VGND.n2432 VGND.t2044 988.926
R530 VGND.t1447 VGND.n2457 988.926
R531 VGND.n2458 VGND.t709 988.926
R532 VGND.t443 VGND.n2483 988.926
R533 VGND.n2484 VGND.t535 988.926
R534 VGND.t1408 VGND.n2514 988.926
R535 VGND.t313 VGND.n2519 988.926
R536 VGND.t1526 VGND.n2524 988.926
R537 VGND.n2525 VGND.t482 988.926
R538 VGND.t46 VGND.n2366 988.926
R539 VGND.n2367 VGND.t2097 988.926
R540 VGND.t2591 VGND.n2392 988.926
R541 VGND.n2393 VGND.t908 988.926
R542 VGND.t1807 VGND.n2418 988.926
R543 VGND.n2419 VGND.t1619 988.926
R544 VGND.t2540 VGND.n2444 988.926
R545 VGND.n2445 VGND.t374 988.926
R546 VGND.t904 VGND.n2470 988.926
R547 VGND.n2471 VGND.t455 988.926
R548 VGND.t339 VGND.n2496 988.926
R549 VGND.n2502 VGND.t106 988.926
R550 VGND.n2501 VGND.t297 988.926
R551 VGND.t725 VGND.n2812 988.926
R552 VGND.n2813 VGND.t327 988.926
R553 VGND.t1063 VGND.n1913 988.926
R554 VGND.n1914 VGND.t1988 988.926
R555 VGND.t2598 VGND.n1924 988.926
R556 VGND.n1925 VGND.t286 988.926
R557 VGND.t1914 VGND.n1935 988.926
R558 VGND.n1936 VGND.t1229 988.926
R559 VGND.t347 VGND.n1946 988.926
R560 VGND.n1947 VGND.t1469 988.926
R561 VGND.t147 VGND.n1957 988.926
R562 VGND.n1958 VGND.t527 988.926
R563 VGND.t1090 VGND.n1968 988.926
R564 VGND.n1969 VGND.t1609 988.926
R565 VGND.t115 VGND.n1979 988.926
R566 VGND.t1123 VGND.n1984 988.926
R567 VGND.n1985 VGND.t1982 988.926
R568 VGND.t139 VGND.n599 988.926
R569 VGND.n2059 VGND.t1811 988.926
R570 VGND.n2058 VGND.t1562 988.926
R571 VGND.n2053 VGND.t921 988.926
R572 VGND.n2048 VGND.t1947 988.926
R573 VGND.n2043 VGND.t1771 988.926
R574 VGND.n2038 VGND.t2036 988.926
R575 VGND.n2033 VGND.t780 988.926
R576 VGND.n2028 VGND.t1066 988.926
R577 VGND.n2023 VGND.t486 988.926
R578 VGND.n2018 VGND.t2150 988.926
R579 VGND.n2013 VGND.t675 988.926
R580 VGND.n2008 VGND.t305 988.926
R581 VGND.n2003 VGND.t1531 988.926
R582 VGND.n601 VGND.t473 988.926
R583 VGND.t762 VGND.n2072 988.926
R584 VGND.t704 VGND.n2077 988.926
R585 VGND.t2467 VGND.n2082 988.926
R586 VGND.t932 VGND.n2087 988.926
R587 VGND.t2079 VGND.n2092 988.926
R588 VGND.t1379 VGND.n2097 988.926
R589 VGND.t2046 VGND.n2102 988.926
R590 VGND.t1449 VGND.n2107 988.926
R591 VGND.t711 VGND.n2112 988.926
R592 VGND.t445 VGND.n2117 988.926
R593 VGND.t537 VGND.n2122 988.926
R594 VGND.n2128 VGND.t1410 988.926
R595 VGND.n2127 VGND.t315 988.926
R596 VGND.t1528 VGND.n2837 988.926
R597 VGND.n2838 VGND.t484 988.926
R598 VGND.n2179 VGND.t48 988.926
R599 VGND.t2099 VGND.n1754 988.926
R600 VGND.t2589 VGND.n1764 988.926
R601 VGND.n1765 VGND.t910 988.926
R602 VGND.t214 VGND.n1775 988.926
R603 VGND.n1776 VGND.t1621 988.926
R604 VGND.t2542 VGND.n1786 988.926
R605 VGND.n1787 VGND.t376 988.926
R606 VGND.t906 VGND.n1797 988.926
R607 VGND.n1798 VGND.t457 988.926
R608 VGND.t637 VGND.n1808 988.926
R609 VGND.n1809 VGND.t108 988.926
R610 VGND.t299 VGND.n1819 988.926
R611 VGND.t727 VGND.n1824 988.926
R612 VGND.n1825 VGND.t329 988.926
R613 VGND.t41 VGND.n1681 988.926
R614 VGND.n1682 VGND.t2091 988.926
R615 VGND.t2595 VGND.n1692 988.926
R616 VGND.t1514 VGND.n1697 988.926
R617 VGND.t1801 VGND.n1702 988.926
R618 VGND.t1617 VGND.n1707 988.926
R619 VGND.t2536 VGND.n1712 988.926
R620 VGND.t370 VGND.n1717 988.926
R621 VGND.t1150 VGND.n1722 988.926
R622 VGND.t453 VGND.n1727 988.926
R623 VGND.t337 VGND.n1732 988.926
R624 VGND.n1849 VGND.t104 988.926
R625 VGND.n1848 VGND.t722 988.926
R626 VGND.n1843 VGND.t814 988.926
R627 VGND.n1734 VGND.t325 988.926
R628 VGND.t1061 VGND.n672 988.926
R629 VGND.t1986 VGND.n677 988.926
R630 VGND.t2600 VGND.n682 988.926
R631 VGND.t918 VGND.n687 988.926
R632 VGND.t1823 VGND.n692 988.926
R633 VGND.t1385 VGND.n697 988.926
R634 VGND.t345 VGND.n702 988.926
R635 VGND.t1467 VGND.n707 988.926
R636 VGND.t145 VGND.n712 988.926
R637 VGND.t525 VGND.n717 988.926
R638 VGND.t1088 VGND.n722 988.926
R639 VGND.n728 VGND.t1607 988.926
R640 VGND.n727 VGND.t113 988.926
R641 VGND.t211 VGND.n2862 988.926
R642 VGND.n2863 VGND.t1980 988.926
R643 VGND.n1355 VGND.t846 988.926
R644 VGND.n877 VGND.t1955 988.926
R645 VGND.n872 VGND.t568 988.926
R646 VGND.t1508 VGND.n821 988.926
R647 VGND.t1799 VGND.n826 988.926
R648 VGND.t1223 VGND.n831 988.926
R649 VGND.t358 VGND.n836 988.926
R650 VGND.t381 VGND.n841 988.926
R651 VGND.t233 VGND.n846 988.926
R652 VGND.t435 VGND.n851 988.926
R653 VGND.n857 VGND.t2165 988.926
R654 VGND.n856 VGND.t2477 988.926
R655 VGND.n1665 VGND.t389 988.926
R656 VGND.n1664 VGND.t673 988.926
R657 VGND.n1659 VGND.t317 988.926
R658 VGND.t758 VGND.n1393 988.926
R659 VGND.t700 VGND.n1398 988.926
R660 VGND.n1399 VGND.t2471 988.926
R661 VGND.t928 VGND.n1493 988.926
R662 VGND.n1494 VGND.t2075 988.926
R663 VGND.t1265 VGND.n1519 988.926
R664 VGND.n1520 VGND.t2042 988.926
R665 VGND.t1445 VGND.n1545 988.926
R666 VGND.t707 VGND.n1550 988.926
R667 VGND.n1556 VGND.t493 988.926
R668 VGND.n1555 VGND.t2156 988.926
R669 VGND.t1406 VGND.n1635 988.926
R670 VGND.t311 VGND.n1640 988.926
R671 VGND.t1524 VGND.n1645 988.926
R672 VGND.n1646 VGND.t480 988.926
R673 VGND.t844 VGND.n1413 988.926
R674 VGND.n1414 VGND.t1953 988.926
R675 VGND.t570 VGND.n1480 988.926
R676 VGND.n1481 VGND.t914 988.926
R677 VGND.t1797 VGND.n1506 988.926
R678 VGND.n1507 VGND.t1221 988.926
R679 VGND.t356 VGND.n1532 988.926
R680 VGND.n1533 VGND.t379 988.926
R681 VGND.t231 VGND.n1569 988.926
R682 VGND.n1585 VGND.t433 988.926
R683 VGND.n1584 VGND.t2163 988.926
R684 VGND.n1579 VGND.t1818 988.926
R685 VGND.n1574 VGND.t387 988.926
R686 VGND.t671 VGND.n2887 988.926
R687 VGND.n2888 VGND.t343 988.926
R688 VGND.n1341 VGND.t184 988.926
R689 VGND.t226 VGND.n1426 988.926
R690 VGND.t1571 VGND.n1431 988.926
R691 VGND.t290 VGND.n1436 988.926
R692 VGND.t1918 VGND.n1441 988.926
R693 VGND.t1231 VGND.n1446 988.926
R694 VGND.t777 VGND.n1451 988.926
R695 VGND.t362 VGND.n1456 988.926
R696 VGND.n1462 VGND.t767 988.926
R697 VGND.n1461 VGND.t529 988.926
R698 VGND.t1092 VGND.n1598 988.926
R699 VGND.t2610 VGND.n1603 988.926
R700 VGND.n1617 VGND.t119 988.926
R701 VGND.n1616 VGND.t1125 988.926
R702 VGND.n1611 VGND.t9 988.926
R703 VGND.t43 VGND.n1034 988.926
R704 VGND.t2093 VGND.n1039 988.926
R705 VGND.n1098 VGND.t2593 988.926
R706 VGND.n1097 VGND.t1516 988.926
R707 VGND.n1092 VGND.t1803 988.926
R708 VGND.n1087 VGND.t1615 988.926
R709 VGND.n1082 VGND.t2534 988.926
R710 VGND.n1077 VGND.t734 988.926
R711 VGND.n1072 VGND.t1148 988.926
R712 VGND.t451 VGND.n1050 988.926
R713 VGND.t335 VGND.n1055 988.926
R714 VGND.t2481 VGND.n1060 988.926
R715 VGND.n1061 VGND.t720 988.926
R716 VGND.t816 VGND.n2907 988.926
R717 VGND.n2908 VGND.t323 988.926
R718 VGND.n1335 VGND.t594 988.926
R719 VGND.t2295 VGND.n929 988.926
R720 VGND.t2273 VGND.n934 988.926
R721 VGND.t589 VGND.n939 988.926
R722 VGND.t578 VGND.n944 988.926
R723 VGND.t2342 VGND.n949 988.926
R724 VGND.t2191 VGND.n954 988.926
R725 VGND.t2170 VGND.n959 988.926
R726 VGND.t2338 VGND.n964 988.926
R727 VGND.t2251 VGND.n969 988.926
R728 VGND.t2238 VGND.n974 988.926
R729 VGND.t613 VGND.n979 988.926
R730 VGND.t2321 VGND.n984 988.926
R731 VGND.t2220 VGND.n989 988.926
R732 VGND.n990 VGND.t622 988.926
R733 VGND.n2248 VGND.n539 934.784
R734 VGND.n116 VGND 927.203
R735 VGND.n134 VGND 927.203
R736 VGND.n2182 VGND 918.774
R737 VGND.n194 VGND 910.346
R738 VGND.n165 VGND 910.346
R739 VGND.t891 VGND.n2967 909.365
R740 VGND.n2285 VGND.n473 900
R741 VGND.n2641 VGND.t1401 852.769
R742 VGND.n2646 VGND.t1035 852.769
R743 VGND.n2651 VGND.t1499 852.769
R744 VGND.n2656 VGND.t1060 852.769
R745 VGND.n2661 VGND.t1160 852.769
R746 VGND.n2666 VGND.t2628 852.769
R747 VGND.n2671 VGND.t158 852.769
R748 VGND.n2672 VGND.t2148 852.769
R749 VGND.n2717 VGND.t2 852.769
R750 VGND.n2718 VGND.t1783 852.769
R751 VGND.n2750 VGND.t877 852.769
R752 VGND.n2756 VGND.t2474 852.769
R753 VGND.t548 VGND.n2755 852.769
R754 VGND.n2790 VGND.t666 852.769
R755 VGND.n2791 VGND.t1031 852.769
R756 VGND.n2935 VGND.t1937 852.769
R757 VGND.t1518 VGND.n2345 852.769
R758 VGND.t213 VGND.n2340 852.769
R759 VGND.t744 VGND.n2335 852.769
R760 VGND.t1365 VGND.n2330 852.769
R761 VGND.t154 VGND.n2325 852.769
R762 VGND.t825 VGND.n2320 852.769
R763 VGND.t2615 VGND.n2315 852.769
R764 VGND.t826 VGND.n2310 852.769
R765 VGND.t2364 VGND.n2305 852.769
R766 VGND.t1943 VGND.n2300 852.769
R767 VGND.t715 VGND.n2295 852.769
R768 VGND.t1120 VGND.n2290 852.769
R769 VGND.n2544 VGND.t1366 852.769
R770 VGND.t24 VGND.n2543 852.769
R771 VGND.t1 VGND.n2538 852.769
R772 VGND.t29 VGND.n208 852.769
R773 VGND.n2354 VGND.t1373 852.769
R774 VGND.n2379 VGND.t549 852.769
R775 VGND.n2380 VGND.t192 852.769
R776 VGND.n2405 VGND.t563 852.769
R777 VGND.n2406 VGND.t1170 852.769
R778 VGND.n2431 VGND.t1497 852.769
R779 VGND.n2432 VGND.t1402 852.769
R780 VGND.n2457 VGND.t103 852.769
R781 VGND.n2458 VGND.t773 852.769
R782 VGND.n2483 VGND.t1156 852.769
R783 VGND.n2484 VGND.t1975 852.769
R784 VGND.n2514 VGND.t1118 852.769
R785 VGND.n2519 VGND.t2475 852.769
R786 VGND.n2524 VGND.t1106 852.769
R787 VGND.n2525 VGND.t1957 852.769
R788 VGND.t640 VGND.n209 852.769
R789 VGND.n2366 VGND.t1504 852.769
R790 VGND.n2367 VGND.t237 852.769
R791 VGND.n2392 VGND.t561 852.769
R792 VGND.n2393 VGND.t1404 852.769
R793 VGND.n2418 VGND.t1403 852.769
R794 VGND.n2419 VGND.t1163 852.769
R795 VGND.n2444 VGND.t878 852.769
R796 VGND.n2445 VGND.t774 852.769
R797 VGND.n2470 VGND.t1507 852.769
R798 VGND.n2471 VGND.t1505 852.769
R799 VGND.n2496 VGND.t1057 852.769
R800 VGND.n2502 VGND.t210 852.769
R801 VGND.t1443 VGND.n2501 852.769
R802 VGND.n2812 VGND.t1370 852.769
R803 VGND.n2813 VGND.t197 852.769
R804 VGND.t199 VGND.n210 852.769
R805 VGND.n1913 VGND.t810 852.769
R806 VGND.n1914 VGND.t1786 852.769
R807 VGND.n1924 VGND.t2161 852.769
R808 VGND.n1925 VGND.t156 852.769
R809 VGND.n1935 VGND.t635 852.769
R810 VGND.n1936 VGND.t463 852.769
R811 VGND.n1946 VGND.t174 852.769
R812 VGND.n1947 VGND.t191 852.769
R813 VGND.n1957 VGND.t2158 852.769
R814 VGND.n1958 VGND.t25 852.769
R815 VGND.n1968 VGND.t2618 852.769
R816 VGND.n1969 VGND.t1169 852.769
R817 VGND.n1979 VGND.t155 852.769
R818 VGND.n1984 VGND.t1944 852.769
R819 VGND.n1985 VGND.t1501 852.769
R820 VGND.t1942 VGND.n211 852.769
R821 VGND.n599 VGND.t1773 852.769
R822 VGND.n2059 VGND.t716 852.769
R823 VGND.t743 VGND.n2058 852.769
R824 VGND.t37 VGND.n2053 852.769
R825 VGND.t670 VGND.n2048 852.769
R826 VGND.t1781 VGND.n2043 852.769
R827 VGND.t1164 VGND.n2038 852.769
R828 VGND.t1152 VGND.n2033 852.769
R829 VGND.t1780 VGND.n2028 852.769
R830 VGND.t27 VGND.n2023 852.769
R831 VGND.t22 VGND.n2018 852.769
R832 VGND.t159 VGND.n2013 852.769
R833 VGND.t102 VGND.n2008 852.769
R834 VGND.t1281 VGND.n2003 852.769
R835 VGND.n601 VGND.t1378 852.769
R836 VGND.t177 VGND.n212 852.769
R837 VGND.n2072 VGND.t157 852.769
R838 VGND.n2077 VGND.t896 852.769
R839 VGND.n2082 VGND.t437 852.769
R840 VGND.n2087 VGND.t1782 852.769
R841 VGND.n2092 VGND.t2687 852.769
R842 VGND.n2097 VGND.t564 852.769
R843 VGND.n2102 VGND.t1372 852.769
R844 VGND.n2107 VGND.t1121 852.769
R845 VGND.n2112 VGND.t1371 852.769
R846 VGND.n2117 VGND.t137 852.769
R847 VGND.n2122 VGND.t175 852.769
R848 VGND.n2128 VGND.t1046 852.769
R849 VGND.t1471 VGND.n2127 852.769
R850 VGND.n2837 VGND.t28 852.769
R851 VGND.n2838 VGND.t757 852.769
R852 VGND.t23 VGND.n213 852.769
R853 VGND.t667 VGND.n2179 852.769
R854 VGND.n1754 VGND.t2129 852.769
R855 VGND.n1764 VGND.t1536 852.769
R856 VGND.n1765 VGND.t2530 852.769
R857 VGND.n1775 VGND.t1059 852.769
R858 VGND.n1776 VGND.t772 852.769
R859 VGND.n1786 VGND.t1105 852.769
R860 VGND.n1787 VGND.t1119 852.769
R861 VGND.n1797 VGND.t818 852.769
R862 VGND.n1798 VGND.t1034 852.769
R863 VGND.n1808 VGND.t1027 852.769
R864 VGND.n1809 VGND.t1388 852.769
R865 VGND.n1819 VGND.t669 852.769
R866 VGND.n1824 VGND.t740 852.769
R867 VGND.n1825 VGND.t2128 852.769
R868 VGND.t1115 VGND.n214 852.769
R869 VGND.n1681 VGND.t738 852.769
R870 VGND.n1682 VGND.t1958 852.769
R871 VGND.n1692 VGND.t828 852.769
R872 VGND.n1697 VGND.t1456 852.769
R873 VGND.n1702 VGND.t1048 852.769
R874 VGND.n1707 VGND.t636 852.769
R875 VGND.n1712 VGND.t1452 852.769
R876 VGND.n1717 VGND.t1028 852.769
R877 VGND.n1722 VGND.t1496 852.769
R878 VGND.n1727 VGND.t1158 852.769
R879 VGND.n1732 VGND.t881 852.769
R880 VGND.n1849 VGND.t1951 852.769
R881 VGND.t94 VGND.n1848 852.769
R882 VGND.t1122 VGND.n1843 852.769
R883 VGND.n1734 VGND.t0 852.769
R884 VGND.t824 VGND.n215 852.769
R885 VGND.n672 VGND.t136 852.769
R886 VGND.n677 VGND.t1377 852.769
R887 VGND.n682 VGND.t173 852.769
R888 VGND.n687 VGND.t1006 852.769
R889 VGND.n692 VGND.t16 852.769
R890 VGND.n697 VGND.t180 852.769
R891 VGND.n702 VGND.t550 852.769
R892 VGND.n707 VGND.t1283 852.769
R893 VGND.n712 VGND.t1375 852.769
R894 VGND.n717 VGND.t2125 852.769
R895 VGND.n722 VGND.t1428 852.769
R896 VGND.n728 VGND.t196 852.769
R897 VGND.t901 VGND.n727 852.769
R898 VGND.n2862 VGND.t1822 852.769
R899 VGND.n2863 VGND.t1073 852.769
R900 VGND.t1369 VGND.n216 852.769
R901 VGND.t178 VGND.n1355 852.769
R902 VGND.t2127 VGND.n877 852.769
R903 VGND.t839 VGND.n872 852.769
R904 VGND.n821 VGND.t1155 852.769
R905 VGND.n826 VGND.t17 852.769
R906 VGND.n831 VGND.t1387 852.769
R907 VGND.n836 VGND.t1519 852.769
R908 VGND.n841 VGND.t1506 852.769
R909 VGND.n846 VGND.t1785 852.769
R910 VGND.n851 VGND.t462 852.769
R911 VGND.n857 VGND.t398 852.769
R912 VGND.t2162 VGND.n856 852.769
R913 VGND.n1665 VGND.t1613 852.769
R914 VGND.t1153 VGND.n1664 852.769
R915 VGND.t695 VGND.n1659 852.769
R916 VGND.t1032 VGND.n217 852.769
R917 VGND.n1393 VGND.t36 852.769
R918 VGND.n1398 VGND.t1058 852.769
R919 VGND.n1399 VGND.t1503 852.769
R920 VGND.n1493 VGND.t1084 852.769
R921 VGND.n1494 VGND.t827 852.769
R922 VGND.n1519 VGND.t2149 852.769
R923 VGND.n1520 VGND.t1367 852.769
R924 VGND.n1545 VGND.t1072 852.769
R925 VGND.n1550 VGND.t1007 852.769
R926 VGND.n1556 VGND.t1033 852.769
R927 VGND.t2003 VGND.n1555 852.769
R928 VGND.n1635 VGND.t1376 852.769
R929 VGND.n1640 VGND.t1611 852.769
R930 VGND.n1645 VGND.t1974 852.769
R931 VGND.n1646 VGND.t190 852.769
R932 VGND.t34 VGND.n218 852.769
R933 VGND.n1413 VGND.t198 852.769
R934 VGND.n1414 VGND.t2619 852.769
R935 VGND.n1480 VGND.t1293 852.769
R936 VGND.n1481 VGND.t1036 852.769
R937 VGND.n1506 VGND.t397 852.769
R938 VGND.n1507 VGND.t26 852.769
R939 VGND.n1532 VGND.t176 852.769
R940 VGND.n1533 VGND.t31 852.769
R941 VGND.n1569 VGND.t1873 852.769
R942 VGND.n1585 VGND.t1154 852.769
R943 VGND.t742 VGND.n1584 852.769
R944 VGND.t193 VGND.n1579 852.769
R945 VGND.t189 VGND.n1574 852.769
R946 VGND.n2887 VGND.t1096 852.769
R947 VGND.n2888 VGND.t1413 852.769
R948 VGND.t1108 VGND.n219 852.769
R949 VGND.n1341 VGND.t1779 852.769
R950 VGND.n1426 VGND.t209 852.769
R951 VGND.n1431 VGND.t1427 852.769
R952 VGND.n1436 VGND.t3 852.769
R953 VGND.n1441 VGND.t681 852.769
R954 VGND.n1446 VGND.t741 852.769
R955 VGND.n1451 VGND.t194 852.769
R956 VGND.n1456 VGND.t1368 852.769
R957 VGND.n1462 VGND.t2518 852.769
R958 VGND.t200 VGND.n1461 852.769
R959 VGND.n1598 VGND.t1157 852.769
R960 VGND.n1603 VGND.t843 852.769
R961 VGND.n1617 VGND.t21 852.769
R962 VGND.t2629 VGND.n1616 852.769
R963 VGND.t539 VGND.n1611 852.769
R964 VGND.t823 VGND.n220 852.769
R965 VGND.n1034 VGND.t1502 852.769
R966 VGND.n1039 VGND.t1498 852.769
R967 VGND.n1098 VGND.t737 852.769
R968 VGND.t736 VGND.n1097 852.769
R969 VGND.t2686 VGND.n1092 852.769
R970 VGND.t33 VGND.n1087 852.769
R971 VGND.t32 VGND.n1082 852.769
R972 VGND.t5 VGND.n1077 852.769
R973 VGND.t562 VGND.n1072 852.769
R974 VGND.n1050 VGND.t153 852.769
R975 VGND.n1055 VGND.t1520 852.769
R976 VGND.n1060 VGND.t739 852.769
R977 VGND.n1061 VGND.t135 852.769
R978 VGND.n2907 VGND.t809 852.769
R979 VGND.n2908 VGND.t1784 852.769
R980 VGND.t164 VGND.n221 852.769
R981 VGND.t880 VGND.n1335 852.769
R982 VGND.n929 VGND.t879 852.769
R983 VGND.n934 VGND.t195 852.769
R984 VGND.n939 VGND.t15 852.769
R985 VGND.n944 VGND.t179 852.769
R986 VGND.n949 VGND.t1426 852.769
R987 VGND.n954 VGND.t565 852.769
R988 VGND.n959 VGND.t1107 852.769
R989 VGND.n964 VGND.t2126 852.769
R990 VGND.n969 VGND.t1374 852.769
R991 VGND.n974 VGND.t771 852.769
R992 VGND.n979 VGND.t2493 852.769
R993 VGND.n984 VGND.t573 852.769
R994 VGND.n989 VGND.t4 852.769
R995 VGND.n990 VGND.t1083 852.769
R996 VGND.n2918 VGND.t1936 852.769
R997 VGND.n2249 VGND 851.341
R998 VGND.n2944 VGND.n2943 846.154
R999 VGND.n2350 VGND.t1666 809.773
R1000 VGND.n2352 VGND.t1741 809.773
R1001 VGND.t1648 VGND.n2353 809.773
R1002 VGND.n473 VGND.t1690 809.773
R1003 VGND.t1762 VGND.n503 809.773
R1004 VGND.t1642 VGND.n504 809.773
R1005 VGND.n2180 VGND.t1684 809.773
R1006 VGND.t1696 VGND.n539 809.773
R1007 VGND.n1387 VGND.t1720 809.773
R1008 VGND.t1651 VGND.n1388 809.773
R1009 VGND.n1339 VGND.t1723 809.773
R1010 VGND.t1753 VGND.n1340 809.773
R1011 VGND.n1338 VGND.t1693 809.773
R1012 VGND.n1336 VGND.t2206 809.773
R1013 VGND.t2391 VGND.t2373 708.047
R1014 VGND.t2373 VGND.t2371 708.047
R1015 VGND.t2371 VGND.t2381 708.047
R1016 VGND.t2381 VGND.t1415 708.047
R1017 VGND.t1415 VGND.t1423 708.047
R1018 VGND.t1423 VGND.t1418 708.047
R1019 VGND.t1418 VGND.t1420 708.047
R1020 VGND.t1133 VGND.t18 708.047
R1021 VGND.t2387 VGND.t2426 708.047
R1022 VGND.t2426 VGND.t2395 708.047
R1023 VGND.t2395 VGND.t2369 708.047
R1024 VGND.t2369 VGND.t1414 708.047
R1025 VGND.t1414 VGND.t1422 708.047
R1026 VGND.t1422 VGND.t1417 708.047
R1027 VGND.t1417 VGND.t1425 708.047
R1028 VGND.t2442 VGND.t2389 708.047
R1029 VGND.t2389 VGND.t2430 708.047
R1030 VGND.t2430 VGND.t2400 708.047
R1031 VGND.t2400 VGND.t755 708.047
R1032 VGND.t755 VGND.t751 708.047
R1033 VGND.t751 VGND.t745 708.047
R1034 VGND.t745 VGND.t747 708.047
R1035 VGND.t1130 VGND.t19 708.047
R1036 VGND.t2418 VGND.t2407 708.047
R1037 VGND.t2407 VGND.t2405 708.047
R1038 VGND.t2405 VGND.t2365 708.047
R1039 VGND.t2365 VGND.t38 708.047
R1040 VGND.t38 VGND.t1140 708.047
R1041 VGND.t1140 VGND.t301 708.047
R1042 VGND.t301 VGND.t1029 708.047
R1043 VGND.t2383 VGND.t2422 708.047
R1044 VGND.t2422 VGND.t2393 708.047
R1045 VGND.t2393 VGND.t2403 708.047
R1046 VGND.t2403 VGND.t181 708.047
R1047 VGND.t181 VGND.t1228 708.047
R1048 VGND.t1228 VGND.t913 708.047
R1049 VGND.t913 VGND.t1226 708.047
R1050 VGND.t2379 VGND.t2435 708.047
R1051 VGND.t2440 VGND.t2379 708.047
R1052 VGND.t2412 VGND.t2440 708.047
R1053 VGND.t753 VGND.t2412 708.047
R1054 VGND.t749 VGND.t753 708.047
R1055 VGND.t754 VGND.t749 708.047
R1056 VGND.t750 VGND.t754 708.047
R1057 VGND.n2971 VGND.n2970 708.047
R1058 VGND.t2606 VGND.t1454 691.188
R1059 VGND.t819 VGND.t2159 691.188
R1060 VGND.t2446 VGND.t2424 657.471
R1061 VGND.t2420 VGND.t892 657.471
R1062 VGND.t2457 VGND.t888 657.471
R1063 VGND.t2397 VGND.t882 657.471
R1064 VGND.t469 VGND.t1394 657.471
R1065 VGND.t74 VGND.t1392 657.471
R1066 VGND.t1323 VGND.t1390 657.471
R1067 VGND.t2258 VGND.t1078 657.471
R1068 VGND.t2424 VGND.t2451 654.197
R1069 VGND.t1078 VGND.t1080 654.197
R1070 VGND VGND.n194 640.614
R1071 VGND VGND.n134 640.614
R1072 VGND VGND.n165 640.614
R1073 VGND.n2182 VGND 640.614
R1074 VGND.n116 VGND 632.184
R1075 VGND.t1934 VGND.t1960 630.62
R1076 VGND.t2089 VGND.t1924 630.62
R1077 VGND.t2597 VGND.t1215 630.62
R1078 VGND.t920 VGND.t1213 630.62
R1079 VGND.t1330 VGND.t1932 630.62
R1080 VGND.t1765 VGND.t2635 630.62
R1081 VGND.t2532 VGND.t2633 630.62
R1082 VGND.t732 VGND.t1930 630.62
R1083 VGND.t1928 VGND.t841 630.62
R1084 VGND.t450 VGND.t2637 630.62
R1085 VGND.t1211 VGND.t1775 630.62
R1086 VGND.t2480 VGND.t1209 630.62
R1087 VGND.t2631 VGND.t718 630.62
R1088 VGND.t1219 VGND.t813 630.62
R1089 VGND.t472 VGND.t1217 630.62
R1090 VGND.t1926 VGND.t610 630.62
R1091 VGND.t2133 VGND.t144 630.62
R1092 VGND.t2544 VGND.t699 630.62
R1093 VGND.t205 VGND.t2466 630.62
R1094 VGND.t203 VGND.t289 630.62
R1095 VGND.t2131 VGND.t2074 630.62
R1096 VGND.t2558 VGND.t1614 630.62
R1097 VGND.t2556 VGND.t2041 630.62
R1098 VGND.t2550 VGND.t1444 630.62
R1099 VGND.t2548 VGND.t1071 630.62
R1100 VGND.t2560 VGND.t447 630.62
R1101 VGND.t2137 VGND.t334 630.62
R1102 VGND.t2135 VGND.t1412 630.62
R1103 VGND.t2554 VGND.t310 630.62
R1104 VGND.t2552 VGND.t1871 630.62
R1105 VGND.t207 VGND.t1985 630.62
R1106 VGND.t2546 VGND.t2232 630.62
R1107 VGND.t40 VGND.t1332 630.62
R1108 VGND.t837 VGND.t2095 630.62
R1109 VGND.t2587 VGND.t2082 630.62
R1110 VGND.t1338 VGND.t926 630.62
R1111 VGND.t1805 VGND.t222 630.62
R1112 VGND.t833 VGND.t1767 630.62
R1113 VGND.t2538 VGND.t831 630.62
R1114 VGND.t220 VGND.t372 630.62
R1115 VGND.t902 VGND.t218 630.62
R1116 VGND.t835 VGND.t460 630.62
R1117 VGND.t1777 VGND.t1336 630.62
R1118 VGND.t1334 VGND.t111 630.62
R1119 VGND.t724 VGND.t829 630.62
R1120 VGND.t730 VGND.t2086 630.62
R1121 VGND.t478 VGND.t2084 630.62
R1122 VGND.t216 VGND.t631 630.62
R1123 VGND.t2522 VGND.t546 630.62
R1124 VGND.t698 VGND.t1888 630.62
R1125 VGND.t2139 VGND.t1573 630.62
R1126 VGND.t1512 VGND.t2528 630.62
R1127 VGND.t2018 VGND.t1795 630.62
R1128 VGND.t1383 VGND.t1884 630.62
R1129 VGND.t1882 VGND.t354 630.62
R1130 VGND.t684 VGND.t2016 630.62
R1131 VGND.t2014 VGND.t1144 630.62
R1132 VGND.t431 VGND.t1886 630.62
R1133 VGND.t2526 VGND.t2491 630.62
R1134 VGND.t1816 VGND.t2524 630.62
R1135 VGND.t2145 VGND.t385 630.62
R1136 VGND.t2143 VGND.t1010 630.62
R1137 VGND.t321 VGND.t2141 630.62
R1138 VGND.t2012 VGND.t2348 630.62
R1139 VGND.t138 VGND.t2626 630.62
R1140 VGND.t1810 VGND.t58 630.62
R1141 VGND.t95 VGND.t1564 630.62
R1142 VGND.t917 VGND.t2487 630.62
R1143 VGND.t2624 VGND.t1946 630.62
R1144 VGND.t2262 VGND.t54 630.62
R1145 VGND.t52 VGND.t2035 630.62
R1146 VGND.t779 VGND.t2622 630.62
R1147 VGND.t2620 VGND.t1065 630.62
R1148 VGND.t491 VGND.t56 630.62
R1149 VGND.t2485 VGND.t332 630.62
R1150 VGND.t680 VGND.t2483 630.62
R1151 VGND.t50 VGND.t304 630.62
R1152 VGND.t1522 VGND.t99 630.62
R1153 VGND.t1979 VGND.t97 630.62
R1154 VGND.t60 VGND.t2204 630.62
R1155 VGND.t1959 VGND.t2024 630.62
R1156 VGND.t2088 VGND.t1600 630.62
R1157 VGND.t2032 VGND.t572 630.62
R1158 VGND.t2030 VGND.t912 630.62
R1159 VGND.t2022 VGND.t1329 630.62
R1160 VGND.t425 VGND.t1764 630.62
R1161 VGND.t423 VGND.t2531 630.62
R1162 VGND.t2020 VGND.t731 630.62
R1163 VGND.t1604 VGND.t840 630.62
R1164 VGND.t427 VGND.t449 630.62
R1165 VGND.t2028 VGND.t1774 630.62
R1166 VGND.t2026 VGND.t2479 630.62
R1167 VGND.t421 VGND.t717 630.62
R1168 VGND.t419 VGND.t812 630.62
R1169 VGND.t471 VGND.t417 630.62
R1170 VGND.t1602 VGND.t608 630.62
R1171 VGND.t45 VGND.t517 630.62
R1172 VGND.t2096 VGND.t507 630.62
R1173 VGND.t1561 VGND.t555 630.62
R1174 VGND.t927 VGND.t523 630.62
R1175 VGND.t1806 VGND.t515 630.62
R1176 VGND.t1768 VGND.t503 630.62
R1177 VGND.t2539 VGND.t501 630.62
R1178 VGND.t373 VGND.t513 630.62
R1179 VGND.t903 VGND.t511 630.62
R1180 VGND.t461 VGND.t505 630.62
R1181 VGND.t1778 VGND.t521 630.62
R1182 VGND.t811 VGND.t519 630.62
R1183 VGND.t499 VGND.t296 630.62
R1184 VGND.t559 VGND.t1530 630.62
R1185 VGND.t479 VGND.t557 630.62
R1186 VGND.t509 VGND.t634 630.62
R1187 VGND.t1012 VGND.t547 630.62
R1188 VGND.t1952 VGND.t201 630.62
R1189 VGND.t567 VGND.t689 630.62
R1190 VGND.t1513 VGND.t687 630.62
R1191 VGND.t1024 VGND.t1796 630.62
R1192 VGND.t1384 VGND.t1791 630.62
R1193 VGND.t1789 VGND.t355 630.62
R1194 VGND.t378 VGND.t1022 630.62
R1195 VGND.t1020 VGND.t1145 630.62
R1196 VGND.t432 VGND.t1793 630.62
R1197 VGND.t1016 VGND.t2492 630.62
R1198 VGND.t1817 VGND.t1014 630.62
R1199 VGND.t1787 VGND.t386 630.62
R1200 VGND.t1011 VGND.t693 630.62
R1201 VGND.t322 VGND.t691 630.62
R1202 VGND.t1018 VGND.t2350 630.62
R1203 VGND.t544 VGND.t1051 630.62
R1204 VGND.t697 VGND.t1041 630.62
R1205 VGND.t1111 VGND.t566 630.62
R1206 VGND.t1511 VGND.t1109 630.62
R1207 VGND.t1321 VGND.t1049 630.62
R1208 VGND.t1381 VGND.t1037 630.62
R1209 VGND.t353 VGND.t2010 630.62
R1210 VGND.t683 VGND.t553 630.62
R1211 VGND.t1143 VGND.t551 630.62
R1212 VGND.t430 VGND.t1039 630.62
R1213 VGND.t2490 VGND.t1055 630.62
R1214 VGND.t1821 VGND.t1053 630.62
R1215 VGND.t2008 VGND.t384 630.62
R1216 VGND.t2006 VGND.t1009 630.62
R1217 VGND.t319 VGND.t1113 630.62
R1218 VGND.t1043 VGND.t2341 630.62
R1219 VGND.t842 VGND.t870 630.62
R1220 VGND.t1809 VGND.t1183 630.62
R1221 VGND.t1567 VGND.t1880 630.62
R1222 VGND.t916 VGND.t1878 630.62
R1223 VGND.t1945 VGND.t868 630.62
R1224 VGND.t1225 VGND.t1179 630.62
R1225 VGND.t2034 VGND.t1177 630.62
R1226 VGND.t366 VGND.t866 630.62
R1227 VGND.t399 VGND.t864 630.62
R1228 VGND.t488 VGND.t1181 630.62
R1229 VGND.t331 VGND.t1876 630.62
R1230 VGND.t677 VGND.t1874 630.62
R1231 VGND.t1175 VGND.t303 630.62
R1232 VGND.t1173 VGND.t1533 630.62
R1233 VGND.t1978 VGND.t1171 630.62
R1234 VGND.t862 VGND.t2199 630.62
R1235 VGND.t1431 VGND.t183 630.62
R1236 VGND.t1359 VGND.t225 630.62
R1237 VGND.t1439 VGND.t2603 630.62
R1238 VGND.t895 VGND.t1437 630.62
R1239 VGND.t1917 VGND.t1429 630.62
R1240 VGND.t1264 VGND.t1355 630.62
R1241 VGND.t776 VGND.t1353 630.62
R1242 VGND.t361 VGND.t2520 630.62
R1243 VGND.t766 VGND.t1363 630.62
R1244 VGND.t534 VGND.t1357 630.62
R1245 VGND.t2155 VGND.t1435 630.62
R1246 VGND.t1433 VGND.t2586 630.62
R1247 VGND.t1351 VGND.t118 630.62
R1248 VGND.t1349 VGND.t1923 630.62
R1249 VGND.t1441 VGND.t342 630.62
R1250 VGND.t1361 VGND.t2300 630.62
R1251 VGND.t1961 VGND.t400 630.62
R1252 VGND.t2090 VGND.t852 630.62
R1253 VGND.t2588 VGND.t408 630.62
R1254 VGND.t406 VGND.t925 630.62
R1255 VGND.t1331 VGND.t860 630.62
R1256 VGND.t848 VGND.t1766 630.62
R1257 VGND.t2533 VGND.t2463 630.62
R1258 VGND.t858 VGND.t733 630.62
R1259 VGND.t1147 VGND.t856 630.62
R1260 VGND.t459 VGND.t850 630.62
R1261 VGND.t404 VGND.t1776 630.62
R1262 VGND.t402 VGND.t110 630.62
R1263 VGND.t719 VGND.t2461 630.62
R1264 VGND.t729 VGND.t2616 630.62
R1265 VGND.t477 VGND.t410 630.62
R1266 VGND.t854 VGND.t628 630.62
R1267 VGND.t2639 VGND.t182 630.62
R1268 VGND.t224 VGND.t1457 630.62
R1269 VGND.t2647 VGND.t1570 630.62
R1270 VGND.t894 VGND.t2645 630.62
R1271 VGND.t1465 VGND.t1916 630.62
R1272 VGND.t1263 VGND.t131 630.62
R1273 VGND.t129 VGND.t349 630.62
R1274 VGND.t360 VGND.t1463 630.62
R1275 VGND.t1461 VGND.t765 630.62
R1276 VGND.t531 VGND.t133 630.62
R1277 VGND.t2643 VGND.t2154 630.62
R1278 VGND.t2641 VGND.t2612 630.62
R1279 VGND.t127 VGND.t117 630.62
R1280 VGND.t125 VGND.t1920 630.62
R1281 VGND.t341 VGND.t123 630.62
R1282 VGND.t1459 VGND.t2297 630.62
R1283 VGND.t143 VGND.t2653 630.62
R1284 VGND.t88 VGND.t1815 630.62
R1285 VGND.t2473 VGND.t1343 630.62
R1286 VGND.t288 VGND.t2659 630.62
R1287 VGND.t2073 VGND.t2651 630.62
R1288 VGND.t2263 VGND.t84 630.62
R1289 VGND.t2040 VGND.t82 630.62
R1290 VGND.t784 VGND.t2649 630.62
R1291 VGND.t1070 VGND.t92 630.62
R1292 VGND.t86 VGND.t492 630.62
R1293 VGND.t2657 VGND.t333 630.62
R1294 VGND.t1405 VGND.t2655 630.62
R1295 VGND.t309 VGND.t80 630.62
R1296 VGND.t1347 VGND.t1523 630.62
R1297 VGND.t1345 VGND.t1984 630.62
R1298 VGND.t90 VGND.t2219 630.62
R1299 VGND.t545 VGND.t169 630.62
R1300 VGND.t696 VGND.t160 630.62
R1301 VGND.t1574 VGND.t1994 630.62
R1302 VGND.t1992 VGND.t1510 630.62
R1303 VGND.t167 VGND.t1322 630.62
R1304 VGND.t1968 VGND.t1382 630.62
R1305 VGND.t1966 VGND.t352 630.62
R1306 VGND.t165 VGND.t682 630.62
R1307 VGND.t1972 VGND.t1142 630.62
R1308 VGND.t429 VGND.t1970 630.62
R1309 VGND.t2489 VGND.t1990 630.62
R1310 VGND.t1820 VGND.t171 630.62
R1311 VGND.t383 VGND.t1964 630.62
R1312 VGND.t1962 VGND.t1008 630.62
R1313 VGND.t320 VGND.t1996 630.62
R1314 VGND.t162 VGND.t2340 630.62
R1315 VGND.t596 VGND.t764 630.62
R1316 VGND.t706 VGND.t2298 630.62
R1317 VGND.t2602 VGND.t2209 630.62
R1318 VGND.t292 VGND.t2187 630.62
R1319 VGND.t2081 VGND.t585 630.62
R1320 VGND.t1770 VGND.t2279 630.62
R1321 VGND.t2048 VGND.t2268 630.62
R1322 VGND.t1451 VGND.t581 630.62
R1323 VGND.t713 VGND.t2346 630.62
R1324 VGND.t448 VGND.t2281 630.62
R1325 VGND.t639 VGND.t2174 630.62
R1326 VGND.t1606 VGND.t629 630.62
R1327 VGND.t112 VGND.t2253 630.62
R1328 VGND.t1872 VGND.t2240 630.62
R1329 VGND.t11 VGND.t2215 630.62
R1330 VGND.t2325 VGND.t2244 630.62
R1331 VGND.n2704 VGND.n327 615.385
R1332 VGND.n2349 VGND.t1269 602.708
R1333 VGND.n3019 VGND.t1269 602.708
R1334 VGND.n3011 VGND.n3010 599.125
R1335 VGND.n194 VGND.n193 599.125
R1336 VGND.n66 VGND.n65 599.125
R1337 VGND.n117 VGND.n116 599.125
R1338 VGND.n134 VGND.n133 599.125
R1339 VGND.n165 VGND.n164 599.125
R1340 VGND.n2210 VGND.n2182 599.125
R1341 VGND.n2972 VGND.n2971 599.125
R1342 VGND VGND.t1976 581.61
R1343 VGND.t1420 VGND 573.181
R1344 VGND VGND.t884 573.181
R1345 VGND.t747 VGND 573.181
R1346 VGND.t1029 VGND 573.181
R1347 VGND.n3013 VGND 564.751
R1348 VGND.t2608 VGND 564.751
R1349 VGND.n3014 VGND 564.751
R1350 VGND.n3012 VGND 556.322
R1351 VGND.t1086 VGND 539.465
R1352 VGND VGND.t1098 539.465
R1353 VGND.t64 VGND.n806 494.779
R1354 VGND.n1166 VGND.t2236 492.058
R1355 VGND.t624 VGND.n1175 492.058
R1356 VGND.n1176 VGND.t600 492.058
R1357 VGND.t2234 VGND.n1188 492.058
R1358 VGND.n1189 VGND.t2222 492.058
R1359 VGND.t2200 VGND.n1207 492.058
R1360 VGND.n1208 VGND.t2311 492.058
R1361 VGND.t2291 VGND.n1220 492.058
R1362 VGND.n1247 VGND.t2195 492.058
R1363 VGND.n1246 VGND.t583 492.058
R1364 VGND.n1240 VGND.t2355 492.058
R1365 VGND.n1239 VGND.t2266 492.058
R1366 VGND.n1233 VGND.t2185 492.058
R1367 VGND.t2344 VGND.n1277 492.058
R1368 VGND.n1278 VGND.t2277 492.058
R1369 VGND.t2416 VGND.t2375 481.877
R1370 VGND.t2451 VGND.t2416 481.877
R1371 VGND.t1080 VGND.t1287 481.877
R1372 VGND.t1287 VGND.t1340 481.877
R1373 VGND.t685 VGND 452.382
R1374 VGND.n1166 VGND.t30 424.312
R1375 VGND.n1175 VGND.t665 424.312
R1376 VGND.n1176 VGND.t1612 424.312
R1377 VGND.n1188 VGND.t1162 424.312
R1378 VGND.n1189 VGND.t150 424.312
R1379 VGND.n1207 VGND.t2685 424.312
R1380 VGND.n1208 VGND.t14 424.312
R1381 VGND.n1220 VGND.t1159 424.312
R1382 VGND.n1247 VGND.t188 424.312
R1383 VGND.t230 VGND.n1246 424.312
R1384 VGND.n1240 VGND.t35 424.312
R1385 VGND.t2167 VGND.n1239 424.312
R1386 VGND.n1233 VGND.t2519 424.312
R1387 VGND.n1277 VGND.t8 424.312
R1388 VGND.n1278 VGND.t543 424.312
R1389 VGND.t149 VGND.n222 424.312
R1390 VGND.t412 VGND 419.68
R1391 VGND.n2284 VGND.n503 413.043
R1392 VGND.t1666 VGND.t2105 408.469
R1393 VGND.t2564 VGND.t141 408.469
R1394 VGND.t240 VGND.t1813 408.469
R1395 VGND.t1865 VGND.t1565 408.469
R1396 VGND.t1235 VGND.t923 408.469
R1397 VGND.t2669 VGND.t1949 408.469
R1398 VGND.t1861 VGND.t1261 408.469
R1399 VGND.t962 VGND.t2038 408.469
R1400 VGND.t782 VGND.t2057 408.469
R1401 VGND.t1297 VGND.t1068 408.469
R1402 VGND.t489 VGND.t1890 408.469
R1403 VGND.t1596 VGND.t2152 408.469
R1404 VGND.t678 VGND.t803 408.469
R1405 VGND.t307 VGND.t994 408.469
R1406 VGND.t954 VGND.t1534 408.469
R1407 VGND.t475 VGND.t1557 408.469
R1408 VGND.t1741 VGND.t647 408.469
R1409 VGND.t186 VGND.t2508 408.469
R1410 VGND.t228 VGND.t938 408.469
R1411 VGND.t1568 VGND.t970 408.469
R1412 VGND.t293 VGND.t2566 408.469
R1413 VGND.t1319 VGND.t1839 408.469
R1414 VGND.t1233 VGND.t966 408.469
R1415 VGND.t350 VGND.t1237 408.469
R1416 VGND.t364 VGND.t2671 408.469
R1417 VGND.t769 VGND.t1863 408.469
R1418 VGND.t532 VGND.t1474 408.469
R1419 VGND.t1094 VGND.t1315 408.469
R1420 VGND.t2613 VGND.t1853 408.469
R1421 VGND.t121 VGND.t1894 408.469
R1422 VGND.t1921 VGND.t1559 408.469
R1423 VGND.t12 VGND.t805 408.469
R1424 VGND.t2055 VGND.t1648 408.469
R1425 VGND.t760 VGND.t1912 408.469
R1426 VGND.t1205 VGND.t702 408.469
R1427 VGND.t2469 VGND.t2498 408.469
R1428 VGND.t795 VGND.t930 408.469
R1429 VGND.t2077 VGND.t2580 408.469
R1430 VGND.t950 VGND.t1267 408.469
R1431 VGND.t2044 VGND.t1549 408.469
R1432 VGND.t1249 VGND.t1447 408.469
R1433 VGND.t709 VGND.t252 408.469
R1434 VGND.t2109 VGND.t443 408.469
R1435 VGND.t535 VGND.t1243 408.469
R1436 VGND.t244 VGND.t1408 408.469
R1437 VGND.t1845 VGND.t313 408.469
R1438 VGND.t1482 VGND.t1526 408.469
R1439 VGND.t482 VGND.t270 408.469
R1440 VGND.t1690 VGND.t2665 408.469
R1441 VGND.t1492 VGND.t46 408.469
R1442 VGND.t2097 VGND.t2069 408.469
R1443 VGND.t1580 VGND.t2591 408.469
R1444 VGND.t908 VGND.t1847 408.469
R1445 VGND.t1189 VGND.t1807 408.469
R1446 VGND.t1619 VGND.t1551 408.469
R1447 VGND.t797 VGND.t2540 408.469
R1448 VGND.t374 VGND.t2582 408.469
R1449 VGND.t952 VGND.t904 408.469
R1450 VGND.t455 VGND.t651 408.469
R1451 VGND.t2574 VGND.t339 408.469
R1452 VGND.t106 VGND.t944 408.469
R1453 VGND.t297 VGND.t2113 408.469
R1454 VGND.t272 VGND.t725 408.469
R1455 VGND.t327 VGND.t248 408.469
R1456 VGND.t1833 VGND.t1762 408.469
R1457 VGND.t280 VGND.t1063 408.469
R1458 VGND.t1988 VGND.t2681 408.469
R1459 VGND.t1301 VGND.t2598 408.469
R1460 VGND.t286 VGND.t1494 408.469
R1461 VGND.t2051 VGND.t1914 408.469
R1462 VGND.t1229 VGND.t799 408.469
R1463 VGND.t1849 VGND.t347 408.469
R1464 VGND.t1469 VGND.t1193 408.469
R1465 VGND.t1553 VGND.t147 408.469
R1466 VGND.t527 VGND.t992 408.469
R1467 VGND.t2514 VGND.t1090 408.469
R1468 VGND.t1609 VGND.t1547 408.469
R1469 VGND.t653 VGND.t115 408.469
R1470 VGND.t250 VGND.t1123 408.469
R1471 VGND.t1982 VGND.t948 408.469
R1472 VGND.t976 VGND.t1669 408.469
R1473 VGND.t256 VGND.t139 408.469
R1474 VGND.t1811 VGND.t1273 408.469
R1475 VGND.t1562 VGND.t1855 408.469
R1476 VGND.t921 VGND.t276 408.469
R1477 VGND.t1947 VGND.t1307 408.469
R1478 VGND.t1771 VGND.t1908 408.469
R1479 VGND.t2036 VGND.t1488 408.469
R1480 VGND.t780 VGND.t1590 408.469
R1481 VGND.t1066 VGND.t791 408.469
R1482 VGND.t486 VGND.t1197 408.469
R1483 VGND.t2150 VGND.t1584 408.469
R1484 VGND.t675 VGND.t787 408.469
R1485 VGND.t305 VGND.t986 408.469
R1486 VGND.t942 VGND.t1531 408.469
R1487 VGND.t473 VGND.t1541 408.469
R1488 VGND.t1255 VGND.t1642 408.469
R1489 VGND.t2496 VGND.t762 408.469
R1490 VGND.t2117 VGND.t704 408.469
R1491 VGND.t960 VGND.t2467 408.469
R1492 VGND.t258 VGND.t932 408.469
R1493 VGND.t1825 VGND.t2079 408.469
R1494 VGND.t1490 VGND.t1379 408.469
R1495 VGND.t278 VGND.t2046 408.469
R1496 VGND.t1313 VGND.t1449 408.469
R1497 VGND.t1910 VGND.t711 408.469
R1498 VGND.t2063 VGND.t445 408.469
R1499 VGND.t1303 VGND.t537 408.469
R1500 VGND.t1410 VGND.t1906 408.469
R1501 VGND.t315 VGND.t1199 408.469
R1502 VGND.t1543 VGND.t1528 408.469
R1503 VGND.t484 VGND.t789 408.469
R1504 VGND.t1684 VGND.t1588 408.469
R1505 VGND.t1900 VGND.t48 408.469
R1506 VGND.t1195 VGND.t2099 408.469
R1507 VGND.t946 VGND.t2589 408.469
R1508 VGND.t910 VGND.t1000 408.469
R1509 VGND.t2570 VGND.t214 408.469
R1510 VGND.t1621 VGND.t2123 408.469
R1511 VGND.t663 VGND.t2542 408.469
R1512 VGND.t376 VGND.t1241 408.469
R1513 VGND.t238 VGND.t906 408.469
R1514 VGND.t457 VGND.t2101 408.469
R1515 VGND.t282 VGND.t637 408.469
R1516 VGND.t108 VGND.t1275 408.469
R1517 VGND.t1837 VGND.t299 408.469
R1518 VGND.t2071 VGND.t727 408.469
R1519 VGND.t329 VGND.t2683 408.469
R1520 VGND.t1305 VGND.t1696 408.469
R1521 VGND.t1484 VGND.t41 408.469
R1522 VGND.t2091 VGND.t2061 408.469
R1523 VGND.t1545 VGND.t2595 408.469
R1524 VGND.t1902 VGND.t1514 408.469
R1525 VGND.t2510 VGND.t1801 408.469
R1526 VGND.t1537 VGND.t1617 408.469
R1527 VGND.t1002 VGND.t2536 408.469
R1528 VGND.t2572 VGND.t370 408.469
R1529 VGND.t936 VGND.t1150 408.469
R1530 VGND.t641 VGND.t453 408.469
R1531 VGND.t2562 VGND.t337 408.469
R1532 VGND.t104 VGND.t2119 408.469
R1533 VGND.t722 VGND.t2103 408.469
R1534 VGND.t262 VGND.t814 408.469
R1535 VGND.t325 VGND.t1277 408.469
R1536 VGND.t1869 VGND.t1624 408.469
R1537 VGND.t274 VGND.t1061 408.469
R1538 VGND.t2679 VGND.t1986 408.469
R1539 VGND.t793 VGND.t2600 408.469
R1540 VGND.t1486 VGND.t918 408.469
R1541 VGND.t1586 VGND.t1823 408.469
R1542 VGND.t1004 VGND.t1385 408.469
R1543 VGND.t1904 VGND.t345 408.469
R1544 VGND.t2512 VGND.t1467 408.469
R1545 VGND.t1539 VGND.t145 408.469
R1546 VGND.t984 VGND.t525 408.469
R1547 VGND.t2504 VGND.t1088 408.469
R1548 VGND.t1607 VGND.t661 408.469
R1549 VGND.t113 VGND.t643 408.469
R1550 VGND.t1279 VGND.t211 408.469
R1551 VGND.t1980 VGND.t2121 408.469
R1552 VGND.t1720 VGND.t645 408.469
R1553 VGND.t846 VGND.t2502 408.469
R1554 VGND.t1955 VGND.t934 408.469
R1555 VGND.t968 VGND.t568 408.469
R1556 VGND.t260 VGND.t1508 408.469
R1557 VGND.t1835 VGND.t1799 408.469
R1558 VGND.t958 VGND.t1223 408.469
R1559 VGND.t284 VGND.t358 408.469
R1560 VGND.t2667 VGND.t381 408.469
R1561 VGND.t1857 VGND.t233 408.469
R1562 VGND.t1472 VGND.t435 408.469
R1563 VGND.t2165 VGND.t1309 408.469
R1564 VGND.t2477 VGND.t1851 408.469
R1565 VGND.t389 VGND.t1207 408.469
R1566 VGND.t673 VGND.t1555 408.469
R1567 VGND.t317 VGND.t801 408.469
R1568 VGND.t1867 VGND.t1651 408.469
R1569 VGND.t266 VGND.t758 408.469
R1570 VGND.t2675 VGND.t700 408.469
R1571 VGND.t2471 VGND.t785 408.469
R1572 VGND.t1480 VGND.t928 408.469
R1573 VGND.t2075 VGND.t1582 408.469
R1574 VGND.t998 VGND.t1265 408.469
R1575 VGND.t2042 VGND.t1898 408.469
R1576 VGND.t2506 VGND.t1445 408.469
R1577 VGND.t659 VGND.t707 408.469
R1578 VGND.t493 VGND.t2584 408.469
R1579 VGND.t2156 VGND.t2500 408.469
R1580 VGND.t657 VGND.t1406 408.469
R1581 VGND.t1251 VGND.t311 408.469
R1582 VGND.t1271 VGND.t1524 408.469
R1583 VGND.t480 VGND.t2115 408.469
R1584 VGND.t1723 VGND.t268 408.469
R1585 VGND.t974 VGND.t844 408.469
R1586 VGND.t1953 VGND.t964 408.469
R1587 VGND.t2059 VGND.t570 408.469
R1588 VGND.t914 VGND.t1827 408.469
R1589 VGND.t1892 VGND.t1797 408.469
R1590 VGND.t1221 VGND.t2049 408.469
R1591 VGND.t1317 VGND.t356 408.469
R1592 VGND.t379 VGND.t996 408.469
R1593 VGND.t1191 VGND.t231 408.469
R1594 VGND.t433 VGND.t1576 408.469
R1595 VGND.t2163 VGND.t988 408.469
R1596 VGND.t1818 VGND.t2516 408.469
R1597 VGND.t387 VGND.t2494 408.469
R1598 VGND.t1245 VGND.t671 408.469
R1599 VGND.t343 VGND.t2576 408.469
R1600 VGND.t242 VGND.t1753 408.469
R1601 VGND.t184 VGND.t1253 408.469
R1602 VGND.t1239 VGND.t226 408.469
R1603 VGND.t2673 VGND.t1571 408.469
R1604 VGND.t978 VGND.t290 408.469
R1605 VGND.t1476 VGND.t1918 408.469
R1606 VGND.t2661 VGND.t1231 408.469
R1607 VGND.t1829 VGND.t777 408.469
R1608 VGND.t1896 VGND.t362 408.469
R1609 VGND.t767 VGND.t2053 408.469
R1610 VGND.t529 VGND.t807 408.469
R1611 VGND.t1203 VGND.t1092 408.469
R1612 VGND.t1592 VGND.t2610 408.469
R1613 VGND.t119 VGND.t1578 408.469
R1614 VGND.t1125 VGND.t2578 408.469
R1615 VGND.t9 VGND.t1185 408.469
R1616 VGND.t940 VGND.t1693 408.469
R1617 VGND.t982 VGND.t43 408.469
R1618 VGND.t2568 VGND.t2093 408.469
R1619 VGND.t2593 VGND.t1841 408.469
R1620 VGND.t1516 VGND.t1257 408.469
R1621 VGND.t1803 VGND.t264 408.469
R1622 VGND.t1615 VGND.t1831 408.469
R1623 VGND.t2534 VGND.t980 408.469
R1624 VGND.t734 VGND.t1478 408.469
R1625 VGND.t2663 VGND.t1148 408.469
R1626 VGND.t1859 VGND.t451 408.469
R1627 VGND.t2067 VGND.t335 408.469
R1628 VGND.t1311 VGND.t2481 408.469
R1629 VGND.t720 VGND.t1295 408.469
R1630 VGND.t1187 VGND.t816 408.469
R1631 VGND.t323 VGND.t1594 408.469
R1632 VGND.t2206 VGND.t1299 408.469
R1633 VGND.t2065 VGND.t594 408.469
R1634 VGND.t1598 VGND.t2295 408.469
R1635 VGND.t655 VGND.t2273 408.469
R1636 VGND.t1201 VGND.t589 408.469
R1637 VGND.t956 VGND.t578 408.469
R1638 VGND.t649 VGND.t2342 408.469
R1639 VGND.t990 VGND.t2191 408.469
R1640 VGND.t254 VGND.t2170 408.469
R1641 VGND.t2111 VGND.t2338 408.469
R1642 VGND.t1247 VGND.t2251 408.469
R1643 VGND.t246 VGND.t2238 408.469
R1644 VGND.t2107 VGND.t613 408.469
R1645 VGND.t972 VGND.t2321 408.469
R1646 VGND.t2677 VGND.t2220 408.469
R1647 VGND.t622 VGND.t1843 408.469
R1648 VGND.t2448 VGND.t2367 397.848
R1649 VGND.t2367 VGND.t2377 397.848
R1650 VGND.t2377 VGND.t2385 397.848
R1651 VGND.t2385 VGND.t886 397.848
R1652 VGND.t886 VGND.t887 397.848
R1653 VGND.t887 VGND.t890 397.848
R1654 VGND.t890 VGND.t891 397.848
R1655 VGND.t1128 VGND.t1453 396.17
R1656 VGND.t875 VGND.t540 396.17
R1657 VGND.n2935 VGND.n2934 394.137
R1658 VGND.n2933 VGND.n208 394.137
R1659 VGND.n2932 VGND.n209 394.137
R1660 VGND.n2931 VGND.n210 394.137
R1661 VGND.n2930 VGND.n211 394.137
R1662 VGND.n2929 VGND.n212 394.137
R1663 VGND.n2928 VGND.n213 394.137
R1664 VGND.n2927 VGND.n214 394.137
R1665 VGND.n2926 VGND.n215 394.137
R1666 VGND.n2925 VGND.n216 394.137
R1667 VGND.n2924 VGND.n217 394.137
R1668 VGND.n2923 VGND.n218 394.137
R1669 VGND.n2922 VGND.n219 394.137
R1670 VGND.n2921 VGND.n220 394.137
R1671 VGND.n2920 VGND.n221 394.137
R1672 VGND.n2919 VGND.n2918 394.137
R1673 VGND.n2285 VGND.t391 387.421
R1674 VGND.n2284 VGND.t72 387.421
R1675 VGND.n2250 VGND.t440 387.421
R1676 VGND.n2248 VGND.t78 387.421
R1677 VGND.n1386 VGND.t6 387.421
R1678 VGND.t541 VGND.t367 362.452
R1679 VGND.t367 VGND.t1086 345.594
R1680 VGND VGND.t70 328.616
R1681 VGND VGND.t872 328.616
R1682 VGND VGND.t68 328.616
R1683 VGND VGND.t66 328.616
R1684 VGND VGND.t495 328.616
R1685 VGND.t632 VGND.t2242 313.776
R1686 VGND.t626 VGND.t2335 313.776
R1687 VGND.t2320 VGND.t2327 313.776
R1688 VGND.t2305 VGND.t2218 313.776
R1689 VGND.t620 VGND.t2230 313.776
R1690 VGND.t604 VGND.t2308 313.776
R1691 VGND.t2233 VGND.t591 313.776
R1692 VGND.t2224 VGND.t2208 313.776
R1693 VGND.t593 VGND.t2202 313.776
R1694 VGND.t606 VGND.t2309 313.776
R1695 VGND.t2205 VGND.t2293 313.776
R1696 VGND.t2284 VGND.t2193 313.776
R1697 VGND.t580 VGND.t587 313.776
R1698 VGND.t575 VGND.t2286 313.776
R1699 VGND.t2265 VGND.t2336 313.776
R1700 VGND.t2189 VGND.t577 313.776
R1701 VGND.t1137 VGND.t1128 311.877
R1702 VGND.t1976 VGND.t875 311.877
R1703 VGND VGND.t1133 303.449
R1704 VGND VGND.t1137 295.019
R1705 VGND.n101 VGND.t2376 287.832
R1706 VGND VGND.t1397 286.591
R1707 VGND.n93 VGND.t2398 282.327
R1708 VGND.n2184 VGND.t470 282.327
R1709 VGND.n104 VGND.t2447 281.13
R1710 VGND.n2189 VGND.t2259 281.13
R1711 VGND.n177 VGND.t2392 280.978
R1712 VGND.n177 VGND.t2433 280.978
R1713 VGND.n78 VGND.t2443 280.978
R1714 VGND.n78 VGND.t2459 280.978
R1715 VGND.n146 VGND.t2419 280.978
R1716 VGND.n146 VGND.t2455 280.978
R1717 VGND.n482 VGND.t1076 280.978
R1718 VGND.n482 VGND.t467 280.978
R1719 VGND.n2263 VGND.t2260 280.978
R1720 VGND.n2263 VGND.t1286 280.978
R1721 VGND.n518 VGND.t69 280.978
R1722 VGND.n518 VGND.t464 280.978
R1723 VGND.n2194 VGND.t1341 280.978
R1724 VGND.t821 VGND 278.161
R1725 VGND.n2970 VGND 271.014
R1726 VGND.n3021 VGND.n4 259.389
R1727 VGND.n2347 VGND.n4 259.389
R1728 VGND.n3022 VGND.n3 252.988
R1729 VGND VGND.t2387 252.875
R1730 VGND VGND.t1135 252.875
R1731 VGND VGND.t1130 252.875
R1732 VGND VGND.t2383 252.875
R1733 VGND.t2435 VGND 252.875
R1734 VGND.n887 VGND.t1300 241.393
R1735 VGND.n330 VGND.t1679 241.393
R1736 VGND.n396 VGND.t2106 241.393
R1737 VGND.n400 VGND.t648 241.393
R1738 VGND.n469 VGND.t2056 241.393
R1739 VGND.n466 VGND.t2666 241.393
R1740 VGND.n625 VGND.t1834 241.393
R1741 VGND.n590 VGND.t977 241.393
R1742 VGND.n587 VGND.t1256 241.393
R1743 VGND.n547 VGND.t1589 241.393
R1744 VGND.n628 VGND.t1306 241.393
R1745 VGND.n632 VGND.t1870 241.393
R1746 VGND.n879 VGND.t646 241.393
R1747 VGND.n800 VGND.t1868 241.393
R1748 VGND.n797 VGND.t269 241.393
R1749 VGND.n882 VGND.t243 241.393
R1750 VGND.n1024 VGND.t941 241.393
R1751 VGND.n1014 VGND.t1682 241.393
R1752 VGND.n1333 VGND.t2066 241.284
R1753 VGND.n894 VGND.t1599 241.284
R1754 VGND.n932 VGND.t656 241.284
R1755 VGND.n937 VGND.t1202 241.284
R1756 VGND.n942 VGND.t957 241.284
R1757 VGND.n947 VGND.t650 241.284
R1758 VGND.n952 VGND.t991 241.284
R1759 VGND.n957 VGND.t255 241.284
R1760 VGND.n962 VGND.t2112 241.284
R1761 VGND.n967 VGND.t1248 241.284
R1762 VGND.n972 VGND.t247 241.284
R1763 VGND.n977 VGND.t2108 241.284
R1764 VGND.n982 VGND.t973 241.284
R1765 VGND.n987 VGND.t2678 241.284
R1766 VGND.n1280 VGND.t1718 241.284
R1767 VGND.n1275 VGND.t1676 241.284
R1768 VGND.n1232 VGND.t1760 241.284
R1769 VGND.n1237 VGND.t1751 241.284
R1770 VGND.n1225 VGND.t1712 241.284
R1771 VGND.n1244 VGND.t1664 241.284
R1772 VGND.n1001 VGND.t1748 241.284
R1773 VGND.n1218 VGND.t1709 241.284
R1774 VGND.n1210 VGND.t1700 241.284
R1775 VGND.n1205 VGND.t1658 241.284
R1776 VGND.n1009 VGND.t1736 241.284
R1777 VGND.n1186 VGND.t1730 241.284
R1778 VGND.n1178 VGND.t1655 241.284
R1779 VGND.n1173 VGND.t1637 241.284
R1780 VGND.n1168 VGND.t1631 241.284
R1781 VGND.n2773 VGND.t1715 241.284
R1782 VGND.n294 VGND.t1673 241.284
R1783 VGND.n2730 VGND.t1757 241.284
R1784 VGND.n2735 VGND.t1745 241.284
R1785 VGND.n312 VGND.t1706 241.284
R1786 VGND.n2726 VGND.t1661 241.284
R1787 VGND.n326 VGND.t1739 241.284
R1788 VGND.n387 VGND.t1703 241.284
R1789 VGND.n384 VGND.t1688 241.284
R1790 VGND.n379 VGND.t1646 241.284
R1791 VGND.n373 VGND.t1733 241.284
R1792 VGND.n368 VGND.t1727 241.284
R1793 VGND.n362 VGND.t1640 241.284
R1794 VGND.n355 VGND.t1634 241.284
R1795 VGND.n2699 VGND.t1628 241.284
R1796 VGND.n2639 VGND.t2565 241.284
R1797 VGND.n2644 VGND.t241 241.284
R1798 VGND.n2649 VGND.t1866 241.284
R1799 VGND.n2654 VGND.t1236 241.284
R1800 VGND.n2659 VGND.t2670 241.284
R1801 VGND.n2664 VGND.t1862 241.284
R1802 VGND.n2669 VGND.t963 241.284
R1803 VGND.n394 VGND.t2058 241.284
R1804 VGND.n2715 VGND.t1298 241.284
R1805 VGND.n320 VGND.t1891 241.284
R1806 VGND.n2748 VGND.t1597 241.284
R1807 VGND.n304 VGND.t804 241.284
R1808 VGND.n2753 VGND.t995 241.284
R1809 VGND.n2788 VGND.t955 241.284
R1810 VGND.n287 VGND.t1558 241.284
R1811 VGND.n2343 VGND.t2509 241.284
R1812 VGND.n2338 VGND.t939 241.284
R1813 VGND.n2333 VGND.t971 241.284
R1814 VGND.n2328 VGND.t2567 241.284
R1815 VGND.n2323 VGND.t1840 241.284
R1816 VGND.n2318 VGND.t967 241.284
R1817 VGND.n2313 VGND.t1238 241.284
R1818 VGND.n2308 VGND.t2672 241.284
R1819 VGND.n2303 VGND.t1864 241.284
R1820 VGND.n2298 VGND.t1475 241.284
R1821 VGND.n2293 VGND.t1316 241.284
R1822 VGND.n2288 VGND.t1854 241.284
R1823 VGND.n415 VGND.t1895 241.284
R1824 VGND.n2541 VGND.t1560 241.284
R1825 VGND.n2536 VGND.t806 241.284
R1826 VGND.n472 VGND.t1913 241.284
R1827 VGND.n2377 VGND.t1206 241.284
R1828 VGND.n460 VGND.t2499 241.284
R1829 VGND.n2403 VGND.t796 241.284
R1830 VGND.n452 VGND.t2581 241.284
R1831 VGND.n2429 VGND.t951 241.284
R1832 VGND.n444 VGND.t1550 241.284
R1833 VGND.n2455 VGND.t1250 241.284
R1834 VGND.n436 VGND.t253 241.284
R1835 VGND.n2481 VGND.t2110 241.284
R1836 VGND.n428 VGND.t1244 241.284
R1837 VGND.n2512 VGND.t245 241.284
R1838 VGND.n2517 VGND.t1846 241.284
R1839 VGND.n2522 VGND.t1483 241.284
R1840 VGND.n2527 VGND.t271 241.284
R1841 VGND.n2364 VGND.t1493 241.284
R1842 VGND.n464 VGND.t2070 241.284
R1843 VGND.n2390 VGND.t1581 241.284
R1844 VGND.n456 VGND.t1848 241.284
R1845 VGND.n2416 VGND.t1190 241.284
R1846 VGND.n448 VGND.t1552 241.284
R1847 VGND.n2442 VGND.t798 241.284
R1848 VGND.n440 VGND.t2583 241.284
R1849 VGND.n2468 VGND.t953 241.284
R1850 VGND.n432 VGND.t652 241.284
R1851 VGND.n2494 VGND.t2575 241.284
R1852 VGND.n424 VGND.t945 241.284
R1853 VGND.n2499 VGND.t2114 241.284
R1854 VGND.n2810 VGND.t273 241.284
R1855 VGND.n2815 VGND.t249 241.284
R1856 VGND.n1911 VGND.t281 241.284
R1857 VGND.n623 VGND.t2682 241.284
R1858 VGND.n1922 VGND.t1302 241.284
R1859 VGND.n620 VGND.t1495 241.284
R1860 VGND.n1933 VGND.t2052 241.284
R1861 VGND.n617 VGND.t800 241.284
R1862 VGND.n1944 VGND.t1850 241.284
R1863 VGND.n614 VGND.t1194 241.284
R1864 VGND.n1955 VGND.t1554 241.284
R1865 VGND.n611 VGND.t993 241.284
R1866 VGND.n1966 VGND.t2515 241.284
R1867 VGND.n608 VGND.t1548 241.284
R1868 VGND.n1977 VGND.t654 241.284
R1869 VGND.n1982 VGND.t251 241.284
R1870 VGND.n1987 VGND.t949 241.284
R1871 VGND.n597 VGND.t257 241.284
R1872 VGND.n594 VGND.t1274 241.284
R1873 VGND.n2056 VGND.t1856 241.284
R1874 VGND.n2051 VGND.t277 241.284
R1875 VGND.n2046 VGND.t1308 241.284
R1876 VGND.n2041 VGND.t1909 241.284
R1877 VGND.n2036 VGND.t1489 241.284
R1878 VGND.n2031 VGND.t1591 241.284
R1879 VGND.n2026 VGND.t792 241.284
R1880 VGND.n2021 VGND.t1198 241.284
R1881 VGND.n2016 VGND.t1585 241.284
R1882 VGND.n2011 VGND.t788 241.284
R1883 VGND.n2006 VGND.t987 241.284
R1884 VGND.n2001 VGND.t943 241.284
R1885 VGND.n1994 VGND.t1542 241.284
R1886 VGND.n2070 VGND.t2497 241.284
R1887 VGND.n2075 VGND.t2118 241.284
R1888 VGND.n2080 VGND.t961 241.284
R1889 VGND.n2085 VGND.t259 241.284
R1890 VGND.n2090 VGND.t1826 241.284
R1891 VGND.n2095 VGND.t1491 241.284
R1892 VGND.n2100 VGND.t279 241.284
R1893 VGND.n2105 VGND.t1314 241.284
R1894 VGND.n2110 VGND.t1911 241.284
R1895 VGND.n2115 VGND.t2064 241.284
R1896 VGND.n2120 VGND.t1304 241.284
R1897 VGND.n585 VGND.t1907 241.284
R1898 VGND.n2125 VGND.t1200 241.284
R1899 VGND.n2835 VGND.t1544 241.284
R1900 VGND.n2840 VGND.t790 241.284
R1901 VGND.n2177 VGND.t1901 241.284
R1902 VGND.n1756 VGND.t1196 241.284
R1903 VGND.n1762 VGND.t947 241.284
R1904 VGND.n1753 VGND.t1001 241.284
R1905 VGND.n1773 VGND.t2571 241.284
R1906 VGND.n1750 VGND.t2124 241.284
R1907 VGND.n1784 VGND.t664 241.284
R1908 VGND.n1747 VGND.t1242 241.284
R1909 VGND.n1795 VGND.t239 241.284
R1910 VGND.n1744 VGND.t2102 241.284
R1911 VGND.n1806 VGND.t283 241.284
R1912 VGND.n1741 VGND.t1276 241.284
R1913 VGND.n1817 VGND.t1838 241.284
R1914 VGND.n1822 VGND.t2072 241.284
R1915 VGND.n1827 VGND.t2684 241.284
R1916 VGND.n1679 VGND.t1485 241.284
R1917 VGND.n1676 VGND.t2062 241.284
R1918 VGND.n1690 VGND.t1546 241.284
R1919 VGND.n1695 VGND.t1903 241.284
R1920 VGND.n1700 VGND.t2511 241.284
R1921 VGND.n1705 VGND.t1538 241.284
R1922 VGND.n1710 VGND.t1003 241.284
R1923 VGND.n1715 VGND.t2573 241.284
R1924 VGND.n1720 VGND.t937 241.284
R1925 VGND.n1725 VGND.t642 241.284
R1926 VGND.n1730 VGND.t2563 241.284
R1927 VGND.n1673 VGND.t2120 241.284
R1928 VGND.n1846 VGND.t2104 241.284
R1929 VGND.n1841 VGND.t263 241.284
R1930 VGND.n1834 VGND.t1278 241.284
R1931 VGND.n670 VGND.t275 241.284
R1932 VGND.n675 VGND.t2680 241.284
R1933 VGND.n680 VGND.t794 241.284
R1934 VGND.n685 VGND.t1487 241.284
R1935 VGND.n690 VGND.t1587 241.284
R1936 VGND.n695 VGND.t1005 241.284
R1937 VGND.n700 VGND.t1905 241.284
R1938 VGND.n705 VGND.t2513 241.284
R1939 VGND.n710 VGND.t1540 241.284
R1940 VGND.n715 VGND.t985 241.284
R1941 VGND.n720 VGND.t2505 241.284
R1942 VGND.n667 VGND.t662 241.284
R1943 VGND.n725 VGND.t644 241.284
R1944 VGND.n2860 VGND.t1280 241.284
R1945 VGND.n2865 VGND.t2122 241.284
R1946 VGND.n1353 VGND.t2503 241.284
R1947 VGND.n875 VGND.t935 241.284
R1948 VGND.n870 VGND.t969 241.284
R1949 VGND.n810 VGND.t261 241.284
R1950 VGND.n824 VGND.t1836 241.284
R1951 VGND.n829 VGND.t959 241.284
R1952 VGND.n834 VGND.t285 241.284
R1953 VGND.n839 VGND.t2668 241.284
R1954 VGND.n844 VGND.t1858 241.284
R1955 VGND.n849 VGND.t1473 241.284
R1956 VGND.n820 VGND.t1310 241.284
R1957 VGND.n854 VGND.t1852 241.284
R1958 VGND.n735 VGND.t1208 241.284
R1959 VGND.n1662 VGND.t1556 241.284
R1960 VGND.n1657 VGND.t802 241.284
R1961 VGND.n1391 VGND.t267 241.284
R1962 VGND.n1396 VGND.t2676 241.284
R1963 VGND.n805 VGND.t786 241.284
R1964 VGND.n1491 VGND.t1481 241.284
R1965 VGND.n777 VGND.t1583 241.284
R1966 VGND.n1517 VGND.t999 241.284
R1967 VGND.n769 VGND.t1899 241.284
R1968 VGND.n1543 VGND.t2507 241.284
R1969 VGND.n1548 VGND.t660 241.284
R1970 VGND.n761 VGND.t2585 241.284
R1971 VGND.n1553 VGND.t2501 241.284
R1972 VGND.n1633 VGND.t658 241.284
R1973 VGND.n1638 VGND.t1252 241.284
R1974 VGND.n1643 VGND.t1272 241.284
R1975 VGND.n1648 VGND.t2116 241.284
R1976 VGND.n1411 VGND.t975 241.284
R1977 VGND.n795 VGND.t965 241.284
R1978 VGND.n1478 VGND.t2060 241.284
R1979 VGND.n781 VGND.t1828 241.284
R1980 VGND.n1504 VGND.t1893 241.284
R1981 VGND.n773 VGND.t2050 241.284
R1982 VGND.n1530 VGND.t1318 241.284
R1983 VGND.n765 VGND.t997 241.284
R1984 VGND.n1567 VGND.t1192 241.284
R1985 VGND.n756 VGND.t1577 241.284
R1986 VGND.n1582 VGND.t989 241.284
R1987 VGND.n1577 VGND.t2517 241.284
R1988 VGND.n1572 VGND.t2495 241.284
R1989 VGND.n2885 VGND.t1246 241.284
R1990 VGND.n2890 VGND.t2577 241.284
R1991 VGND.n885 VGND.t1254 241.284
R1992 VGND.n1424 VGND.t1240 241.284
R1993 VGND.n1429 VGND.t2674 241.284
R1994 VGND.n1434 VGND.t979 241.284
R1995 VGND.n1439 VGND.t1477 241.284
R1996 VGND.n1444 VGND.t2662 241.284
R1997 VGND.n1449 VGND.t1830 241.284
R1998 VGND.n1454 VGND.t1897 241.284
R1999 VGND.n791 VGND.t2054 241.284
R2000 VGND.n1459 VGND.t808 241.284
R2001 VGND.n1596 VGND.t1204 241.284
R2002 VGND.n1601 VGND.t1593 241.284
R2003 VGND.n750 VGND.t1579 241.284
R2004 VGND.n1614 VGND.t2579 241.284
R2005 VGND.n1609 VGND.t1186 241.284
R2006 VGND.n1032 VGND.t983 241.284
R2007 VGND.n1037 VGND.t2569 241.284
R2008 VGND.n1029 VGND.t1842 241.284
R2009 VGND.n1095 VGND.t1258 241.284
R2010 VGND.n1090 VGND.t265 241.284
R2011 VGND.n1085 VGND.t1832 241.284
R2012 VGND.n1080 VGND.t981 241.284
R2013 VGND.n1075 VGND.t1479 241.284
R2014 VGND.n1070 VGND.t2664 241.284
R2015 VGND.n1043 VGND.t1860 241.284
R2016 VGND.n1053 VGND.t2068 241.284
R2017 VGND.n1058 VGND.t1312 241.284
R2018 VGND.n1049 VGND.t1296 241.284
R2019 VGND.n2905 VGND.t1188 241.284
R2020 VGND.n2910 VGND.t1595 241.284
R2021 VGND.n928 VGND.t1844 241.284
R2022 VGND.t2105 VGND.t1934 222.15
R2023 VGND.t1960 VGND.t1401 222.15
R2024 VGND.t1924 VGND.t2564 222.15
R2025 VGND.t1035 VGND.t2089 222.15
R2026 VGND.t1215 VGND.t240 222.15
R2027 VGND.t1499 VGND.t2597 222.15
R2028 VGND.t1213 VGND.t1865 222.15
R2029 VGND.t1060 VGND.t920 222.15
R2030 VGND.t1932 VGND.t1235 222.15
R2031 VGND.t1160 VGND.t1330 222.15
R2032 VGND.t2635 VGND.t2669 222.15
R2033 VGND.t2628 VGND.t1765 222.15
R2034 VGND.t2633 VGND.t1861 222.15
R2035 VGND.t158 VGND.t2532 222.15
R2036 VGND.t1930 VGND.t962 222.15
R2037 VGND.t2148 VGND.t732 222.15
R2038 VGND.t2057 VGND.t1928 222.15
R2039 VGND.t841 VGND.t2 222.15
R2040 VGND.t2637 VGND.t1297 222.15
R2041 VGND.t1783 VGND.t450 222.15
R2042 VGND.t1890 VGND.t1211 222.15
R2043 VGND.t1775 VGND.t877 222.15
R2044 VGND.t1209 VGND.t1596 222.15
R2045 VGND.t2474 VGND.t2480 222.15
R2046 VGND.t803 VGND.t2631 222.15
R2047 VGND.t718 VGND.t548 222.15
R2048 VGND.t994 VGND.t1219 222.15
R2049 VGND.t813 VGND.t666 222.15
R2050 VGND.t1217 VGND.t954 222.15
R2051 VGND.t1031 VGND.t472 222.15
R2052 VGND.t1557 VGND.t1926 222.15
R2053 VGND.t610 VGND.t1937 222.15
R2054 VGND.t647 VGND.t2133 222.15
R2055 VGND.t144 VGND.t1518 222.15
R2056 VGND.t2508 VGND.t2544 222.15
R2057 VGND.t699 VGND.t213 222.15
R2058 VGND.t938 VGND.t205 222.15
R2059 VGND.t2466 VGND.t744 222.15
R2060 VGND.t970 VGND.t203 222.15
R2061 VGND.t289 VGND.t1365 222.15
R2062 VGND.t2566 VGND.t2131 222.15
R2063 VGND.t2074 VGND.t154 222.15
R2064 VGND.t1839 VGND.t2558 222.15
R2065 VGND.t1614 VGND.t825 222.15
R2066 VGND.t966 VGND.t2556 222.15
R2067 VGND.t2041 VGND.t2615 222.15
R2068 VGND.t1237 VGND.t2550 222.15
R2069 VGND.t1444 VGND.t826 222.15
R2070 VGND.t2671 VGND.t2548 222.15
R2071 VGND.t1071 VGND.t2364 222.15
R2072 VGND.t1863 VGND.t2560 222.15
R2073 VGND.t447 VGND.t1943 222.15
R2074 VGND.t1474 VGND.t2137 222.15
R2075 VGND.t334 VGND.t715 222.15
R2076 VGND.t1315 VGND.t2135 222.15
R2077 VGND.t1412 VGND.t1120 222.15
R2078 VGND.t1853 VGND.t2554 222.15
R2079 VGND.t310 VGND.t1366 222.15
R2080 VGND.t1894 VGND.t2552 222.15
R2081 VGND.t1871 VGND.t24 222.15
R2082 VGND.t1559 VGND.t207 222.15
R2083 VGND.t1985 VGND.t1 222.15
R2084 VGND.t805 VGND.t2546 222.15
R2085 VGND.t2232 VGND.t29 222.15
R2086 VGND.t1332 VGND.t2055 222.15
R2087 VGND.t1373 VGND.t40 222.15
R2088 VGND.t1912 VGND.t837 222.15
R2089 VGND.t2095 VGND.t549 222.15
R2090 VGND.t2082 VGND.t1205 222.15
R2091 VGND.t192 VGND.t2587 222.15
R2092 VGND.t2498 VGND.t1338 222.15
R2093 VGND.t926 VGND.t563 222.15
R2094 VGND.t222 VGND.t795 222.15
R2095 VGND.t1170 VGND.t1805 222.15
R2096 VGND.t2580 VGND.t833 222.15
R2097 VGND.t1767 VGND.t1497 222.15
R2098 VGND.t831 VGND.t950 222.15
R2099 VGND.t1402 VGND.t2538 222.15
R2100 VGND.t1549 VGND.t220 222.15
R2101 VGND.t372 VGND.t103 222.15
R2102 VGND.t218 VGND.t1249 222.15
R2103 VGND.t773 VGND.t902 222.15
R2104 VGND.t252 VGND.t835 222.15
R2105 VGND.t460 VGND.t1156 222.15
R2106 VGND.t1336 VGND.t2109 222.15
R2107 VGND.t1975 VGND.t1777 222.15
R2108 VGND.t1243 VGND.t1334 222.15
R2109 VGND.t111 VGND.t1118 222.15
R2110 VGND.t829 VGND.t244 222.15
R2111 VGND.t2475 VGND.t724 222.15
R2112 VGND.t2086 VGND.t1845 222.15
R2113 VGND.t1106 VGND.t730 222.15
R2114 VGND.t2084 VGND.t1482 222.15
R2115 VGND.t1957 VGND.t478 222.15
R2116 VGND.t270 VGND.t216 222.15
R2117 VGND.t631 VGND.t640 222.15
R2118 VGND.t2665 VGND.t2522 222.15
R2119 VGND.t546 VGND.t1504 222.15
R2120 VGND.t1888 VGND.t1492 222.15
R2121 VGND.t237 VGND.t698 222.15
R2122 VGND.t2069 VGND.t2139 222.15
R2123 VGND.t1573 VGND.t561 222.15
R2124 VGND.t2528 VGND.t1580 222.15
R2125 VGND.t1404 VGND.t1512 222.15
R2126 VGND.t1847 VGND.t2018 222.15
R2127 VGND.t1795 VGND.t1403 222.15
R2128 VGND.t1884 VGND.t1189 222.15
R2129 VGND.t1163 VGND.t1383 222.15
R2130 VGND.t1551 VGND.t1882 222.15
R2131 VGND.t354 VGND.t878 222.15
R2132 VGND.t2016 VGND.t797 222.15
R2133 VGND.t774 VGND.t684 222.15
R2134 VGND.t2582 VGND.t2014 222.15
R2135 VGND.t1144 VGND.t1507 222.15
R2136 VGND.t1886 VGND.t952 222.15
R2137 VGND.t1505 VGND.t431 222.15
R2138 VGND.t651 VGND.t2526 222.15
R2139 VGND.t2491 VGND.t1057 222.15
R2140 VGND.t2524 VGND.t2574 222.15
R2141 VGND.t210 VGND.t1816 222.15
R2142 VGND.t944 VGND.t2145 222.15
R2143 VGND.t385 VGND.t1443 222.15
R2144 VGND.t2113 VGND.t2143 222.15
R2145 VGND.t1010 VGND.t1370 222.15
R2146 VGND.t2141 VGND.t272 222.15
R2147 VGND.t197 VGND.t321 222.15
R2148 VGND.t248 VGND.t2012 222.15
R2149 VGND.t2348 VGND.t199 222.15
R2150 VGND.t2626 VGND.t1833 222.15
R2151 VGND.t810 VGND.t138 222.15
R2152 VGND.t58 VGND.t280 222.15
R2153 VGND.t1786 VGND.t1810 222.15
R2154 VGND.t2681 VGND.t95 222.15
R2155 VGND.t1564 VGND.t2161 222.15
R2156 VGND.t2487 VGND.t1301 222.15
R2157 VGND.t156 VGND.t917 222.15
R2158 VGND.t1494 VGND.t2624 222.15
R2159 VGND.t1946 VGND.t635 222.15
R2160 VGND.t54 VGND.t2051 222.15
R2161 VGND.t463 VGND.t2262 222.15
R2162 VGND.t799 VGND.t52 222.15
R2163 VGND.t2035 VGND.t174 222.15
R2164 VGND.t2622 VGND.t1849 222.15
R2165 VGND.t191 VGND.t779 222.15
R2166 VGND.t1193 VGND.t2620 222.15
R2167 VGND.t1065 VGND.t2158 222.15
R2168 VGND.t56 VGND.t1553 222.15
R2169 VGND.t25 VGND.t491 222.15
R2170 VGND.t992 VGND.t2485 222.15
R2171 VGND.t332 VGND.t2618 222.15
R2172 VGND.t2483 VGND.t2514 222.15
R2173 VGND.t1169 VGND.t680 222.15
R2174 VGND.t1547 VGND.t50 222.15
R2175 VGND.t304 VGND.t155 222.15
R2176 VGND.t99 VGND.t653 222.15
R2177 VGND.t1944 VGND.t1522 222.15
R2178 VGND.t97 VGND.t250 222.15
R2179 VGND.t1501 VGND.t1979 222.15
R2180 VGND.t948 VGND.t60 222.15
R2181 VGND.t2204 VGND.t1942 222.15
R2182 VGND.t2024 VGND.t976 222.15
R2183 VGND.t1773 VGND.t1959 222.15
R2184 VGND.t1600 VGND.t256 222.15
R2185 VGND.t716 VGND.t2088 222.15
R2186 VGND.t1273 VGND.t2032 222.15
R2187 VGND.t572 VGND.t743 222.15
R2188 VGND.t1855 VGND.t2030 222.15
R2189 VGND.t912 VGND.t37 222.15
R2190 VGND.t276 VGND.t2022 222.15
R2191 VGND.t1329 VGND.t670 222.15
R2192 VGND.t1307 VGND.t425 222.15
R2193 VGND.t1764 VGND.t1781 222.15
R2194 VGND.t1908 VGND.t423 222.15
R2195 VGND.t2531 VGND.t1164 222.15
R2196 VGND.t1488 VGND.t2020 222.15
R2197 VGND.t731 VGND.t1152 222.15
R2198 VGND.t1590 VGND.t1604 222.15
R2199 VGND.t840 VGND.t1780 222.15
R2200 VGND.t791 VGND.t427 222.15
R2201 VGND.t449 VGND.t27 222.15
R2202 VGND.t1197 VGND.t2028 222.15
R2203 VGND.t1774 VGND.t22 222.15
R2204 VGND.t1584 VGND.t2026 222.15
R2205 VGND.t2479 VGND.t159 222.15
R2206 VGND.t787 VGND.t421 222.15
R2207 VGND.t717 VGND.t102 222.15
R2208 VGND.t986 VGND.t419 222.15
R2209 VGND.t812 VGND.t1281 222.15
R2210 VGND.t417 VGND.t942 222.15
R2211 VGND.t1378 VGND.t471 222.15
R2212 VGND.t1541 VGND.t1602 222.15
R2213 VGND.t608 VGND.t177 222.15
R2214 VGND.t517 VGND.t1255 222.15
R2215 VGND.t157 VGND.t45 222.15
R2216 VGND.t507 VGND.t2496 222.15
R2217 VGND.t896 VGND.t2096 222.15
R2218 VGND.t555 VGND.t2117 222.15
R2219 VGND.t437 VGND.t1561 222.15
R2220 VGND.t523 VGND.t960 222.15
R2221 VGND.t1782 VGND.t927 222.15
R2222 VGND.t515 VGND.t258 222.15
R2223 VGND.t2687 VGND.t1806 222.15
R2224 VGND.t503 VGND.t1825 222.15
R2225 VGND.t564 VGND.t1768 222.15
R2226 VGND.t501 VGND.t1490 222.15
R2227 VGND.t1372 VGND.t2539 222.15
R2228 VGND.t513 VGND.t278 222.15
R2229 VGND.t1121 VGND.t373 222.15
R2230 VGND.t511 VGND.t1313 222.15
R2231 VGND.t1371 VGND.t903 222.15
R2232 VGND.t505 VGND.t1910 222.15
R2233 VGND.t137 VGND.t461 222.15
R2234 VGND.t521 VGND.t2063 222.15
R2235 VGND.t175 VGND.t1778 222.15
R2236 VGND.t519 VGND.t1303 222.15
R2237 VGND.t1046 VGND.t811 222.15
R2238 VGND.t1906 VGND.t499 222.15
R2239 VGND.t296 VGND.t1471 222.15
R2240 VGND.t1199 VGND.t559 222.15
R2241 VGND.t1530 VGND.t28 222.15
R2242 VGND.t557 VGND.t1543 222.15
R2243 VGND.t757 VGND.t479 222.15
R2244 VGND.t789 VGND.t509 222.15
R2245 VGND.t634 VGND.t23 222.15
R2246 VGND.t1588 VGND.t1012 222.15
R2247 VGND.t547 VGND.t667 222.15
R2248 VGND.t201 VGND.t1900 222.15
R2249 VGND.t2129 VGND.t1952 222.15
R2250 VGND.t689 VGND.t1195 222.15
R2251 VGND.t1536 VGND.t567 222.15
R2252 VGND.t687 VGND.t946 222.15
R2253 VGND.t2530 VGND.t1513 222.15
R2254 VGND.t1000 VGND.t1024 222.15
R2255 VGND.t1796 VGND.t1059 222.15
R2256 VGND.t1791 VGND.t2570 222.15
R2257 VGND.t772 VGND.t1384 222.15
R2258 VGND.t2123 VGND.t1789 222.15
R2259 VGND.t355 VGND.t1105 222.15
R2260 VGND.t1022 VGND.t663 222.15
R2261 VGND.t1119 VGND.t378 222.15
R2262 VGND.t1241 VGND.t1020 222.15
R2263 VGND.t1145 VGND.t818 222.15
R2264 VGND.t1793 VGND.t238 222.15
R2265 VGND.t1034 VGND.t432 222.15
R2266 VGND.t2101 VGND.t1016 222.15
R2267 VGND.t2492 VGND.t1027 222.15
R2268 VGND.t1014 VGND.t282 222.15
R2269 VGND.t1388 VGND.t1817 222.15
R2270 VGND.t1275 VGND.t1787 222.15
R2271 VGND.t386 VGND.t669 222.15
R2272 VGND.t693 VGND.t1837 222.15
R2273 VGND.t740 VGND.t1011 222.15
R2274 VGND.t691 VGND.t2071 222.15
R2275 VGND.t2128 VGND.t322 222.15
R2276 VGND.t2683 VGND.t1018 222.15
R2277 VGND.t2350 VGND.t1115 222.15
R2278 VGND.t1051 VGND.t1305 222.15
R2279 VGND.t738 VGND.t544 222.15
R2280 VGND.t1041 VGND.t1484 222.15
R2281 VGND.t1958 VGND.t697 222.15
R2282 VGND.t2061 VGND.t1111 222.15
R2283 VGND.t566 VGND.t828 222.15
R2284 VGND.t1109 VGND.t1545 222.15
R2285 VGND.t1456 VGND.t1511 222.15
R2286 VGND.t1049 VGND.t1902 222.15
R2287 VGND.t1048 VGND.t1321 222.15
R2288 VGND.t1037 VGND.t2510 222.15
R2289 VGND.t636 VGND.t1381 222.15
R2290 VGND.t2010 VGND.t1537 222.15
R2291 VGND.t1452 VGND.t353 222.15
R2292 VGND.t553 VGND.t1002 222.15
R2293 VGND.t1028 VGND.t683 222.15
R2294 VGND.t551 VGND.t2572 222.15
R2295 VGND.t1496 VGND.t1143 222.15
R2296 VGND.t1039 VGND.t936 222.15
R2297 VGND.t1158 VGND.t430 222.15
R2298 VGND.t1055 VGND.t641 222.15
R2299 VGND.t881 VGND.t2490 222.15
R2300 VGND.t1053 VGND.t2562 222.15
R2301 VGND.t1951 VGND.t1821 222.15
R2302 VGND.t2119 VGND.t2008 222.15
R2303 VGND.t384 VGND.t94 222.15
R2304 VGND.t2103 VGND.t2006 222.15
R2305 VGND.t1009 VGND.t1122 222.15
R2306 VGND.t1113 VGND.t262 222.15
R2307 VGND.t0 VGND.t319 222.15
R2308 VGND.t1277 VGND.t1043 222.15
R2309 VGND.t2341 VGND.t824 222.15
R2310 VGND.t870 VGND.t1869 222.15
R2311 VGND.t136 VGND.t842 222.15
R2312 VGND.t1183 VGND.t274 222.15
R2313 VGND.t1377 VGND.t1809 222.15
R2314 VGND.t1880 VGND.t2679 222.15
R2315 VGND.t173 VGND.t1567 222.15
R2316 VGND.t1878 VGND.t793 222.15
R2317 VGND.t1006 VGND.t916 222.15
R2318 VGND.t868 VGND.t1486 222.15
R2319 VGND.t16 VGND.t1945 222.15
R2320 VGND.t1179 VGND.t1586 222.15
R2321 VGND.t180 VGND.t1225 222.15
R2322 VGND.t1177 VGND.t1004 222.15
R2323 VGND.t550 VGND.t2034 222.15
R2324 VGND.t866 VGND.t1904 222.15
R2325 VGND.t1283 VGND.t366 222.15
R2326 VGND.t864 VGND.t2512 222.15
R2327 VGND.t1375 VGND.t399 222.15
R2328 VGND.t1181 VGND.t1539 222.15
R2329 VGND.t2125 VGND.t488 222.15
R2330 VGND.t1876 VGND.t984 222.15
R2331 VGND.t1428 VGND.t331 222.15
R2332 VGND.t1874 VGND.t2504 222.15
R2333 VGND.t196 VGND.t677 222.15
R2334 VGND.t661 VGND.t1175 222.15
R2335 VGND.t303 VGND.t901 222.15
R2336 VGND.t643 VGND.t1173 222.15
R2337 VGND.t1533 VGND.t1822 222.15
R2338 VGND.t1171 VGND.t1279 222.15
R2339 VGND.t1073 VGND.t1978 222.15
R2340 VGND.t2121 VGND.t862 222.15
R2341 VGND.t2199 VGND.t1369 222.15
R2342 VGND.t645 VGND.t1431 222.15
R2343 VGND.t183 VGND.t178 222.15
R2344 VGND.t2502 VGND.t1359 222.15
R2345 VGND.t225 VGND.t2127 222.15
R2346 VGND.t934 VGND.t1439 222.15
R2347 VGND.t2603 VGND.t839 222.15
R2348 VGND.t1437 VGND.t968 222.15
R2349 VGND.t1155 VGND.t895 222.15
R2350 VGND.t1429 VGND.t260 222.15
R2351 VGND.t17 VGND.t1917 222.15
R2352 VGND.t1355 VGND.t1835 222.15
R2353 VGND.t1387 VGND.t1264 222.15
R2354 VGND.t1353 VGND.t958 222.15
R2355 VGND.t1519 VGND.t776 222.15
R2356 VGND.t2520 VGND.t284 222.15
R2357 VGND.t1506 VGND.t361 222.15
R2358 VGND.t1363 VGND.t2667 222.15
R2359 VGND.t1785 VGND.t766 222.15
R2360 VGND.t1357 VGND.t1857 222.15
R2361 VGND.t462 VGND.t534 222.15
R2362 VGND.t1435 VGND.t1472 222.15
R2363 VGND.t398 VGND.t2155 222.15
R2364 VGND.t1309 VGND.t1433 222.15
R2365 VGND.t2586 VGND.t2162 222.15
R2366 VGND.t1851 VGND.t1351 222.15
R2367 VGND.t118 VGND.t1613 222.15
R2368 VGND.t1207 VGND.t1349 222.15
R2369 VGND.t1923 VGND.t1153 222.15
R2370 VGND.t1555 VGND.t1441 222.15
R2371 VGND.t342 VGND.t695 222.15
R2372 VGND.t801 VGND.t1361 222.15
R2373 VGND.t2300 VGND.t1032 222.15
R2374 VGND.t400 VGND.t1867 222.15
R2375 VGND.t36 VGND.t1961 222.15
R2376 VGND.t852 VGND.t266 222.15
R2377 VGND.t1058 VGND.t2090 222.15
R2378 VGND.t408 VGND.t2675 222.15
R2379 VGND.t1503 VGND.t2588 222.15
R2380 VGND.t785 VGND.t406 222.15
R2381 VGND.t925 VGND.t1084 222.15
R2382 VGND.t860 VGND.t1480 222.15
R2383 VGND.t827 VGND.t1331 222.15
R2384 VGND.t1582 VGND.t848 222.15
R2385 VGND.t1766 VGND.t2149 222.15
R2386 VGND.t2463 VGND.t998 222.15
R2387 VGND.t1367 VGND.t2533 222.15
R2388 VGND.t1898 VGND.t858 222.15
R2389 VGND.t733 VGND.t1072 222.15
R2390 VGND.t856 VGND.t2506 222.15
R2391 VGND.t1007 VGND.t1147 222.15
R2392 VGND.t850 VGND.t659 222.15
R2393 VGND.t1033 VGND.t459 222.15
R2394 VGND.t2584 VGND.t404 222.15
R2395 VGND.t1776 VGND.t2003 222.15
R2396 VGND.t2500 VGND.t402 222.15
R2397 VGND.t110 VGND.t1376 222.15
R2398 VGND.t2461 VGND.t657 222.15
R2399 VGND.t1611 VGND.t719 222.15
R2400 VGND.t2616 VGND.t1251 222.15
R2401 VGND.t1974 VGND.t729 222.15
R2402 VGND.t410 VGND.t1271 222.15
R2403 VGND.t190 VGND.t477 222.15
R2404 VGND.t2115 VGND.t854 222.15
R2405 VGND.t628 VGND.t34 222.15
R2406 VGND.t268 VGND.t2639 222.15
R2407 VGND.t182 VGND.t198 222.15
R2408 VGND.t1457 VGND.t974 222.15
R2409 VGND.t2619 VGND.t224 222.15
R2410 VGND.t964 VGND.t2647 222.15
R2411 VGND.t1570 VGND.t1293 222.15
R2412 VGND.t2645 VGND.t2059 222.15
R2413 VGND.t1036 VGND.t894 222.15
R2414 VGND.t1827 VGND.t1465 222.15
R2415 VGND.t1916 VGND.t397 222.15
R2416 VGND.t131 VGND.t1892 222.15
R2417 VGND.t26 VGND.t1263 222.15
R2418 VGND.t2049 VGND.t129 222.15
R2419 VGND.t349 VGND.t176 222.15
R2420 VGND.t1463 VGND.t1317 222.15
R2421 VGND.t31 VGND.t360 222.15
R2422 VGND.t996 VGND.t1461 222.15
R2423 VGND.t765 VGND.t1873 222.15
R2424 VGND.t133 VGND.t1191 222.15
R2425 VGND.t1154 VGND.t531 222.15
R2426 VGND.t1576 VGND.t2643 222.15
R2427 VGND.t2154 VGND.t742 222.15
R2428 VGND.t988 VGND.t2641 222.15
R2429 VGND.t2612 VGND.t193 222.15
R2430 VGND.t2516 VGND.t127 222.15
R2431 VGND.t117 VGND.t189 222.15
R2432 VGND.t2494 VGND.t125 222.15
R2433 VGND.t1920 VGND.t1096 222.15
R2434 VGND.t123 VGND.t1245 222.15
R2435 VGND.t1413 VGND.t341 222.15
R2436 VGND.t2576 VGND.t1459 222.15
R2437 VGND.t2297 VGND.t1108 222.15
R2438 VGND.t2653 VGND.t242 222.15
R2439 VGND.t1779 VGND.t143 222.15
R2440 VGND.t1253 VGND.t88 222.15
R2441 VGND.t1815 VGND.t209 222.15
R2442 VGND.t1343 VGND.t1239 222.15
R2443 VGND.t1427 VGND.t2473 222.15
R2444 VGND.t2659 VGND.t2673 222.15
R2445 VGND.t3 VGND.t288 222.15
R2446 VGND.t2651 VGND.t978 222.15
R2447 VGND.t681 VGND.t2073 222.15
R2448 VGND.t84 VGND.t1476 222.15
R2449 VGND.t741 VGND.t2263 222.15
R2450 VGND.t82 VGND.t2661 222.15
R2451 VGND.t194 VGND.t2040 222.15
R2452 VGND.t2649 VGND.t1829 222.15
R2453 VGND.t1368 VGND.t784 222.15
R2454 VGND.t92 VGND.t1896 222.15
R2455 VGND.t2518 VGND.t1070 222.15
R2456 VGND.t2053 VGND.t86 222.15
R2457 VGND.t492 VGND.t200 222.15
R2458 VGND.t807 VGND.t2657 222.15
R2459 VGND.t333 VGND.t1157 222.15
R2460 VGND.t2655 VGND.t1203 222.15
R2461 VGND.t843 VGND.t1405 222.15
R2462 VGND.t80 VGND.t1592 222.15
R2463 VGND.t21 VGND.t309 222.15
R2464 VGND.t1578 VGND.t1347 222.15
R2465 VGND.t1523 VGND.t2629 222.15
R2466 VGND.t2578 VGND.t1345 222.15
R2467 VGND.t1984 VGND.t539 222.15
R2468 VGND.t1185 VGND.t90 222.15
R2469 VGND.t2219 VGND.t823 222.15
R2470 VGND.t169 VGND.t940 222.15
R2471 VGND.t1502 VGND.t545 222.15
R2472 VGND.t160 VGND.t982 222.15
R2473 VGND.t1498 VGND.t696 222.15
R2474 VGND.t1994 VGND.t2568 222.15
R2475 VGND.t737 VGND.t1574 222.15
R2476 VGND.t1841 VGND.t1992 222.15
R2477 VGND.t1510 VGND.t736 222.15
R2478 VGND.t1257 VGND.t167 222.15
R2479 VGND.t1322 VGND.t2686 222.15
R2480 VGND.t264 VGND.t1968 222.15
R2481 VGND.t1382 VGND.t33 222.15
R2482 VGND.t1831 VGND.t1966 222.15
R2483 VGND.t352 VGND.t32 222.15
R2484 VGND.t980 VGND.t165 222.15
R2485 VGND.t682 VGND.t5 222.15
R2486 VGND.t1478 VGND.t1972 222.15
R2487 VGND.t1142 VGND.t562 222.15
R2488 VGND.t1970 VGND.t2663 222.15
R2489 VGND.t153 VGND.t429 222.15
R2490 VGND.t1990 VGND.t1859 222.15
R2491 VGND.t1520 VGND.t2489 222.15
R2492 VGND.t171 VGND.t2067 222.15
R2493 VGND.t739 VGND.t1820 222.15
R2494 VGND.t1964 VGND.t1311 222.15
R2495 VGND.t135 VGND.t383 222.15
R2496 VGND.t1295 VGND.t1962 222.15
R2497 VGND.t1008 VGND.t809 222.15
R2498 VGND.t1996 VGND.t1187 222.15
R2499 VGND.t1784 VGND.t320 222.15
R2500 VGND.t1594 VGND.t162 222.15
R2501 VGND.t2340 VGND.t164 222.15
R2502 VGND.t1299 VGND.t596 222.15
R2503 VGND.t764 VGND.t880 222.15
R2504 VGND.t2298 VGND.t2065 222.15
R2505 VGND.t879 VGND.t706 222.15
R2506 VGND.t2209 VGND.t1598 222.15
R2507 VGND.t195 VGND.t2602 222.15
R2508 VGND.t2187 VGND.t655 222.15
R2509 VGND.t15 VGND.t292 222.15
R2510 VGND.t585 VGND.t1201 222.15
R2511 VGND.t179 VGND.t2081 222.15
R2512 VGND.t2279 VGND.t956 222.15
R2513 VGND.t1426 VGND.t1770 222.15
R2514 VGND.t2268 VGND.t649 222.15
R2515 VGND.t565 VGND.t2048 222.15
R2516 VGND.t581 VGND.t990 222.15
R2517 VGND.t1107 VGND.t1451 222.15
R2518 VGND.t2346 VGND.t254 222.15
R2519 VGND.t2126 VGND.t713 222.15
R2520 VGND.t2281 VGND.t2111 222.15
R2521 VGND.t1374 VGND.t448 222.15
R2522 VGND.t2174 VGND.t1247 222.15
R2523 VGND.t771 VGND.t639 222.15
R2524 VGND.t629 VGND.t246 222.15
R2525 VGND.t2493 VGND.t1606 222.15
R2526 VGND.t2253 VGND.t2107 222.15
R2527 VGND.t573 VGND.t112 222.15
R2528 VGND.t2240 VGND.t972 222.15
R2529 VGND.t4 VGND.t1872 222.15
R2530 VGND.t2215 VGND.t2677 222.15
R2531 VGND.t1083 VGND.t11 222.15
R2532 VGND.t1843 VGND.t2325 222.15
R2533 VGND.t2244 VGND.t1936 222.15
R2534 VGND.n2346 VGND.n3 218.73
R2535 VGND.n489 VGND.n487 214.365
R2536 VGND.n489 VGND.n488 214.365
R2537 VGND.n479 VGND.n477 214.365
R2538 VGND.n479 VGND.n478 214.365
R2539 VGND.n497 VGND.n495 214.365
R2540 VGND.n497 VGND.n496 214.365
R2541 VGND.n2270 VGND.n2268 214.365
R2542 VGND.n2270 VGND.n2269 214.365
R2543 VGND.n2260 VGND.n2258 214.365
R2544 VGND.n2260 VGND.n2259 214.365
R2545 VGND.n2278 VGND.n2276 214.365
R2546 VGND.n2278 VGND.n2277 214.365
R2547 VGND.n525 VGND.n523 214.365
R2548 VGND.n525 VGND.n524 214.365
R2549 VGND.n515 VGND.n513 214.365
R2550 VGND.n515 VGND.n514 214.365
R2551 VGND.n533 VGND.n531 214.365
R2552 VGND.n533 VGND.n532 214.365
R2553 VGND.n2191 VGND.n2190 214.365
R2554 VGND.n1140 VGND.n1139 213.613
R2555 VGND.n1142 VGND.n1141 213.613
R2556 VGND.n1112 VGND.n1110 213.613
R2557 VGND.n1112 VGND.n1111 213.613
R2558 VGND.n1115 VGND.n1113 213.613
R2559 VGND.n1115 VGND.n1114 213.613
R2560 VGND.n2236 VGND.n2229 213.613
R2561 VGND.n2236 VGND.n2230 213.613
R2562 VGND.n2234 VGND.n2231 213.613
R2563 VGND.n2234 VGND.n2233 213.613
R2564 VGND.n1374 VGND.n1367 213.613
R2565 VGND.n1374 VGND.n1368 213.613
R2566 VGND.n1372 VGND.n1369 213.613
R2567 VGND.n1372 VGND.n1371 213.613
R2568 VGND.n1154 VGND.t1389 211.359
R2569 VGND.n179 VGND.n175 207.965
R2570 VGND.n179 VGND.n176 207.965
R2571 VGND.n173 VGND.n171 207.965
R2572 VGND.n173 VGND.n172 207.965
R2573 VGND.n186 VGND.n169 207.965
R2574 VGND.n186 VGND.n170 207.965
R2575 VGND.n98 VGND.n97 207.965
R2576 VGND.n110 VGND.n95 207.965
R2577 VGND.n102 VGND.n100 207.965
R2578 VGND.n80 VGND.n76 207.965
R2579 VGND.n80 VGND.n77 207.965
R2580 VGND.n74 VGND.n72 207.965
R2581 VGND.n74 VGND.n73 207.965
R2582 VGND.n87 VGND.n70 207.965
R2583 VGND.n87 VGND.n71 207.965
R2584 VGND.n148 VGND.n144 207.965
R2585 VGND.n148 VGND.n145 207.965
R2586 VGND.n142 VGND.n140 207.965
R2587 VGND.n142 VGND.n141 207.965
R2588 VGND.n155 VGND.n138 207.965
R2589 VGND.n155 VGND.n139 207.965
R2590 VGND.n2188 VGND.n2187 207.965
R2591 VGND.n2205 VGND.n2185 207.965
R2592 VGND.n2981 VGND.n2979 207.213
R2593 VGND.n2981 VGND.n2980 207.213
R2594 VGND.n2985 VGND.n2976 207.213
R2595 VGND.n2985 VGND.n2977 207.213
R2596 VGND.n18 VGND.n16 207.213
R2597 VGND.n18 VGND.n17 207.213
R2598 VGND.n22 VGND.n14 207.213
R2599 VGND.n22 VGND.n15 207.213
R2600 VGND.n2951 VGND.n2950 207.213
R2601 VGND.n2955 VGND.n2949 207.213
R2602 VGND.n44 VGND.n42 207.213
R2603 VGND.n44 VGND.n43 207.213
R2604 VGND.n48 VGND.n40 207.213
R2605 VGND.n48 VGND.n41 207.213
R2606 VGND.n109 VGND.n96 207.213
R2607 VGND.n2204 VGND.n2186 207.213
R2608 VGND.t1681 VGND.t2323 203.242
R2609 VGND.t2236 VGND.t1630 203.242
R2610 VGND.t1636 VGND.t624 203.242
R2611 VGND.t600 VGND.t1654 203.242
R2612 VGND.t1729 VGND.t2234 203.242
R2613 VGND.t2222 VGND.t1735 203.242
R2614 VGND.t1657 VGND.t2200 203.242
R2615 VGND.t2311 VGND.t1699 203.242
R2616 VGND.t1708 VGND.t2291 203.242
R2617 VGND.t2195 VGND.t1747 203.242
R2618 VGND.t1663 VGND.t583 203.242
R2619 VGND.t2355 VGND.t1711 203.242
R2620 VGND.t1750 VGND.t2266 203.242
R2621 VGND.t2185 VGND.t1759 203.242
R2622 VGND.t1675 VGND.t2344 203.242
R2623 VGND.t2277 VGND.t1717 203.242
R2624 VGND VGND.n332 194.419
R2625 VGND VGND.n356 194.419
R2626 VGND VGND.n363 194.419
R2627 VGND VGND.n366 194.419
R2628 VGND VGND.n374 194.419
R2629 VGND VGND.n377 194.419
R2630 VGND VGND.n385 194.419
R2631 VGND VGND.n324 194.419
R2632 VGND VGND.n313 194.419
R2633 VGND VGND.n308 194.419
R2634 VGND VGND.n310 194.419
R2635 VGND VGND.n2729 194.419
R2636 VGND VGND.n292 194.419
R2637 VGND VGND.n295 194.419
R2638 VGND VGND.n202 194.419
R2639 VGND.n887 VGND.n886 194.391
R2640 VGND.n1332 VGND.n889 194.391
R2641 VGND.n895 VGND.n893 194.391
R2642 VGND.n931 VGND.n930 194.391
R2643 VGND.n936 VGND.n935 194.391
R2644 VGND.n941 VGND.n940 194.391
R2645 VGND.n946 VGND.n945 194.391
R2646 VGND.n951 VGND.n950 194.391
R2647 VGND.n956 VGND.n955 194.391
R2648 VGND.n961 VGND.n960 194.391
R2649 VGND.n966 VGND.n965 194.391
R2650 VGND.n971 VGND.n970 194.391
R2651 VGND.n976 VGND.n975 194.391
R2652 VGND.n981 VGND.n980 194.391
R2653 VGND.n986 VGND.n985 194.391
R2654 VGND.n1281 VGND.n996 194.391
R2655 VGND.n1274 VGND.n1273 194.391
R2656 VGND.n1231 VGND.n1230 194.391
R2657 VGND.n1236 VGND.n1229 194.391
R2658 VGND.n1227 VGND.n1226 194.391
R2659 VGND.n1243 VGND.n1224 194.391
R2660 VGND.n1222 VGND.n1221 194.391
R2661 VGND.n1217 VGND.n1216 194.391
R2662 VGND.n1211 VGND.n1002 194.391
R2663 VGND.n1204 VGND.n1203 194.391
R2664 VGND.n1008 VGND.n1007 194.391
R2665 VGND.n1185 VGND.n1184 194.391
R2666 VGND.n1179 VGND.n1010 194.391
R2667 VGND.n1172 VGND.n1171 194.391
R2668 VGND.n1169 VGND.n1012 194.391
R2669 VGND.n330 VGND.n329 194.391
R2670 VGND.n396 VGND.n395 194.391
R2671 VGND.n2638 VGND.n2637 194.391
R2672 VGND.n2643 VGND.n2642 194.391
R2673 VGND.n2648 VGND.n2647 194.391
R2674 VGND.n2653 VGND.n2652 194.391
R2675 VGND.n2658 VGND.n2657 194.391
R2676 VGND.n2663 VGND.n2662 194.391
R2677 VGND.n2668 VGND.n2667 194.391
R2678 VGND.n393 VGND.n392 194.391
R2679 VGND.n2714 VGND.n2713 194.391
R2680 VGND.n319 VGND.n318 194.391
R2681 VGND.n2747 VGND.n2746 194.391
R2682 VGND.n303 VGND.n302 194.391
R2683 VGND.n2752 VGND.n2751 194.391
R2684 VGND.n2787 VGND.n2786 194.391
R2685 VGND.n286 VGND.n285 194.391
R2686 VGND.n400 VGND.n399 194.391
R2687 VGND.n2342 VGND.n2341 194.391
R2688 VGND.n2337 VGND.n2336 194.391
R2689 VGND.n2332 VGND.n2331 194.391
R2690 VGND.n2327 VGND.n2326 194.391
R2691 VGND.n2322 VGND.n2321 194.391
R2692 VGND.n2317 VGND.n2316 194.391
R2693 VGND.n2312 VGND.n2311 194.391
R2694 VGND.n2307 VGND.n2306 194.391
R2695 VGND.n2302 VGND.n2301 194.391
R2696 VGND.n2297 VGND.n2296 194.391
R2697 VGND.n2292 VGND.n2291 194.391
R2698 VGND.n2287 VGND.n2286 194.391
R2699 VGND.n414 VGND.n413 194.391
R2700 VGND.n2540 VGND.n2539 194.391
R2701 VGND.n2535 VGND.n416 194.391
R2702 VGND.n469 VGND.n468 194.391
R2703 VGND.n471 VGND.n470 194.391
R2704 VGND.n2376 VGND.n2375 194.391
R2705 VGND.n459 VGND.n458 194.391
R2706 VGND.n2402 VGND.n2401 194.391
R2707 VGND.n451 VGND.n450 194.391
R2708 VGND.n2428 VGND.n2427 194.391
R2709 VGND.n443 VGND.n442 194.391
R2710 VGND.n2454 VGND.n2453 194.391
R2711 VGND.n435 VGND.n434 194.391
R2712 VGND.n2480 VGND.n2479 194.391
R2713 VGND.n427 VGND.n426 194.391
R2714 VGND.n2511 VGND.n2510 194.391
R2715 VGND.n2516 VGND.n2515 194.391
R2716 VGND.n2521 VGND.n2520 194.391
R2717 VGND.n2528 VGND.n418 194.391
R2718 VGND.n466 VGND.n465 194.391
R2719 VGND.n2363 VGND.n2362 194.391
R2720 VGND.n463 VGND.n462 194.391
R2721 VGND.n2389 VGND.n2388 194.391
R2722 VGND.n455 VGND.n454 194.391
R2723 VGND.n2415 VGND.n2414 194.391
R2724 VGND.n447 VGND.n446 194.391
R2725 VGND.n2441 VGND.n2440 194.391
R2726 VGND.n439 VGND.n438 194.391
R2727 VGND.n2467 VGND.n2466 194.391
R2728 VGND.n431 VGND.n430 194.391
R2729 VGND.n2493 VGND.n2492 194.391
R2730 VGND.n423 VGND.n422 194.391
R2731 VGND.n2498 VGND.n2497 194.391
R2732 VGND.n2809 VGND.n2808 194.391
R2733 VGND.n2816 VGND.n276 194.391
R2734 VGND.n625 VGND.n624 194.391
R2735 VGND.n1910 VGND.n1909 194.391
R2736 VGND.n622 VGND.n621 194.391
R2737 VGND.n1921 VGND.n1920 194.391
R2738 VGND.n619 VGND.n618 194.391
R2739 VGND.n1932 VGND.n1931 194.391
R2740 VGND.n616 VGND.n615 194.391
R2741 VGND.n1943 VGND.n1942 194.391
R2742 VGND.n613 VGND.n612 194.391
R2743 VGND.n1954 VGND.n1953 194.391
R2744 VGND.n610 VGND.n609 194.391
R2745 VGND.n1965 VGND.n1964 194.391
R2746 VGND.n607 VGND.n606 194.391
R2747 VGND.n1976 VGND.n1975 194.391
R2748 VGND.n1981 VGND.n1980 194.391
R2749 VGND.n1988 VGND.n605 194.391
R2750 VGND.n590 VGND.n589 194.391
R2751 VGND.n596 VGND.n595 194.391
R2752 VGND.n593 VGND.n592 194.391
R2753 VGND.n2055 VGND.n2054 194.391
R2754 VGND.n2050 VGND.n2049 194.391
R2755 VGND.n2045 VGND.n2044 194.391
R2756 VGND.n2040 VGND.n2039 194.391
R2757 VGND.n2035 VGND.n2034 194.391
R2758 VGND.n2030 VGND.n2029 194.391
R2759 VGND.n2025 VGND.n2024 194.391
R2760 VGND.n2020 VGND.n2019 194.391
R2761 VGND.n2015 VGND.n2014 194.391
R2762 VGND.n2010 VGND.n2009 194.391
R2763 VGND.n2005 VGND.n2004 194.391
R2764 VGND.n2000 VGND.n600 194.391
R2765 VGND.n1995 VGND.n1993 194.391
R2766 VGND.n587 VGND.n586 194.391
R2767 VGND.n2069 VGND.n2068 194.391
R2768 VGND.n2074 VGND.n2073 194.391
R2769 VGND.n2079 VGND.n2078 194.391
R2770 VGND.n2084 VGND.n2083 194.391
R2771 VGND.n2089 VGND.n2088 194.391
R2772 VGND.n2094 VGND.n2093 194.391
R2773 VGND.n2099 VGND.n2098 194.391
R2774 VGND.n2104 VGND.n2103 194.391
R2775 VGND.n2109 VGND.n2108 194.391
R2776 VGND.n2114 VGND.n2113 194.391
R2777 VGND.n2119 VGND.n2118 194.391
R2778 VGND.n584 VGND.n583 194.391
R2779 VGND.n2124 VGND.n2123 194.391
R2780 VGND.n2834 VGND.n2833 194.391
R2781 VGND.n2841 VGND.n264 194.391
R2782 VGND.n547 VGND.n546 194.391
R2783 VGND.n2176 VGND.n549 194.391
R2784 VGND.n1757 VGND.n1755 194.391
R2785 VGND.n1761 VGND.n1760 194.391
R2786 VGND.n1752 VGND.n1751 194.391
R2787 VGND.n1772 VGND.n1771 194.391
R2788 VGND.n1749 VGND.n1748 194.391
R2789 VGND.n1783 VGND.n1782 194.391
R2790 VGND.n1746 VGND.n1745 194.391
R2791 VGND.n1794 VGND.n1793 194.391
R2792 VGND.n1743 VGND.n1742 194.391
R2793 VGND.n1805 VGND.n1804 194.391
R2794 VGND.n1740 VGND.n1739 194.391
R2795 VGND.n1816 VGND.n1815 194.391
R2796 VGND.n1821 VGND.n1820 194.391
R2797 VGND.n1828 VGND.n1738 194.391
R2798 VGND.n628 VGND.n627 194.391
R2799 VGND.n1678 VGND.n1677 194.391
R2800 VGND.n1675 VGND.n1674 194.391
R2801 VGND.n1689 VGND.n1688 194.391
R2802 VGND.n1694 VGND.n1693 194.391
R2803 VGND.n1699 VGND.n1698 194.391
R2804 VGND.n1704 VGND.n1703 194.391
R2805 VGND.n1709 VGND.n1708 194.391
R2806 VGND.n1714 VGND.n1713 194.391
R2807 VGND.n1719 VGND.n1718 194.391
R2808 VGND.n1724 VGND.n1723 194.391
R2809 VGND.n1729 VGND.n1728 194.391
R2810 VGND.n1672 VGND.n1671 194.391
R2811 VGND.n1845 VGND.n1844 194.391
R2812 VGND.n1840 VGND.n1733 194.391
R2813 VGND.n1835 VGND.n1833 194.391
R2814 VGND.n632 VGND.n631 194.391
R2815 VGND.n669 VGND.n668 194.391
R2816 VGND.n674 VGND.n673 194.391
R2817 VGND.n679 VGND.n678 194.391
R2818 VGND.n684 VGND.n683 194.391
R2819 VGND.n689 VGND.n688 194.391
R2820 VGND.n694 VGND.n693 194.391
R2821 VGND.n699 VGND.n698 194.391
R2822 VGND.n704 VGND.n703 194.391
R2823 VGND.n709 VGND.n708 194.391
R2824 VGND.n714 VGND.n713 194.391
R2825 VGND.n719 VGND.n718 194.391
R2826 VGND.n666 VGND.n665 194.391
R2827 VGND.n724 VGND.n723 194.391
R2828 VGND.n2859 VGND.n2858 194.391
R2829 VGND.n2866 VGND.n252 194.391
R2830 VGND.n879 VGND.n878 194.391
R2831 VGND.n1352 VGND.n1351 194.391
R2832 VGND.n874 VGND.n873 194.391
R2833 VGND.n869 VGND.n807 194.391
R2834 VGND.n811 VGND.n809 194.391
R2835 VGND.n823 VGND.n822 194.391
R2836 VGND.n828 VGND.n827 194.391
R2837 VGND.n833 VGND.n832 194.391
R2838 VGND.n838 VGND.n837 194.391
R2839 VGND.n843 VGND.n842 194.391
R2840 VGND.n848 VGND.n847 194.391
R2841 VGND.n819 VGND.n818 194.391
R2842 VGND.n853 VGND.n852 194.391
R2843 VGND.n734 VGND.n733 194.391
R2844 VGND.n1661 VGND.n1660 194.391
R2845 VGND.n1656 VGND.n736 194.391
R2846 VGND.n800 VGND.n799 194.391
R2847 VGND.n1390 VGND.n1389 194.391
R2848 VGND.n1395 VGND.n1394 194.391
R2849 VGND.n804 VGND.n803 194.391
R2850 VGND.n1490 VGND.n1489 194.391
R2851 VGND.n776 VGND.n775 194.391
R2852 VGND.n1516 VGND.n1515 194.391
R2853 VGND.n768 VGND.n767 194.391
R2854 VGND.n1542 VGND.n1541 194.391
R2855 VGND.n1547 VGND.n1546 194.391
R2856 VGND.n760 VGND.n759 194.391
R2857 VGND.n1552 VGND.n1551 194.391
R2858 VGND.n1632 VGND.n1631 194.391
R2859 VGND.n1637 VGND.n1636 194.391
R2860 VGND.n1642 VGND.n1641 194.391
R2861 VGND.n1649 VGND.n739 194.391
R2862 VGND.n797 VGND.n796 194.391
R2863 VGND.n1410 VGND.n1409 194.391
R2864 VGND.n794 VGND.n793 194.391
R2865 VGND.n1477 VGND.n1476 194.391
R2866 VGND.n780 VGND.n779 194.391
R2867 VGND.n1503 VGND.n1502 194.391
R2868 VGND.n772 VGND.n771 194.391
R2869 VGND.n1529 VGND.n1528 194.391
R2870 VGND.n764 VGND.n763 194.391
R2871 VGND.n1566 VGND.n1565 194.391
R2872 VGND.n755 VGND.n754 194.391
R2873 VGND.n1581 VGND.n1580 194.391
R2874 VGND.n1576 VGND.n1575 194.391
R2875 VGND.n1571 VGND.n1570 194.391
R2876 VGND.n2884 VGND.n2883 194.391
R2877 VGND.n2891 VGND.n239 194.391
R2878 VGND.n882 VGND.n881 194.391
R2879 VGND.n884 VGND.n883 194.391
R2880 VGND.n1423 VGND.n1422 194.391
R2881 VGND.n1428 VGND.n1427 194.391
R2882 VGND.n1433 VGND.n1432 194.391
R2883 VGND.n1438 VGND.n1437 194.391
R2884 VGND.n1443 VGND.n1442 194.391
R2885 VGND.n1448 VGND.n1447 194.391
R2886 VGND.n1453 VGND.n1452 194.391
R2887 VGND.n790 VGND.n789 194.391
R2888 VGND.n1458 VGND.n1457 194.391
R2889 VGND.n1595 VGND.n1594 194.391
R2890 VGND.n1600 VGND.n1599 194.391
R2891 VGND.n749 VGND.n748 194.391
R2892 VGND.n1613 VGND.n1612 194.391
R2893 VGND.n1608 VGND.n1604 194.391
R2894 VGND.n1024 VGND.n1023 194.391
R2895 VGND.n1031 VGND.n1030 194.391
R2896 VGND.n1036 VGND.n1035 194.391
R2897 VGND.n1028 VGND.n1027 194.391
R2898 VGND.n1094 VGND.n1093 194.391
R2899 VGND.n1089 VGND.n1088 194.391
R2900 VGND.n1084 VGND.n1083 194.391
R2901 VGND.n1079 VGND.n1078 194.391
R2902 VGND.n1074 VGND.n1073 194.391
R2903 VGND.n1069 VGND.n1040 194.391
R2904 VGND.n1044 VGND.n1042 194.391
R2905 VGND.n1052 VGND.n1051 194.391
R2906 VGND.n1057 VGND.n1056 194.391
R2907 VGND.n1048 VGND.n1047 194.391
R2908 VGND.n2904 VGND.n2903 194.391
R2909 VGND.n2911 VGND.n227 194.391
R2910 VGND.n1014 VGND.n1013 194.391
R2911 VGND.n927 VGND.n926 194.391
R2912 VGND.n2606 VGND.n2605 161.308
R2913 VGND.n2603 VGND.n2602 161.308
R2914 VGND.n2600 VGND.n2599 161.308
R2915 VGND.n2597 VGND.n2596 161.308
R2916 VGND.n2594 VGND.n2593 161.308
R2917 VGND.n2591 VGND.n2590 161.308
R2918 VGND.n2588 VGND.n2587 161.308
R2919 VGND.n2585 VGND.n2584 161.308
R2920 VGND.n2582 VGND.n2581 161.308
R2921 VGND.n2579 VGND.n2578 161.308
R2922 VGND.n2576 VGND.n2575 161.308
R2923 VGND.n2573 VGND.n2572 161.308
R2924 VGND.n2570 VGND.n2569 161.308
R2925 VGND.n2567 VGND.n2566 161.308
R2926 VGND.n2564 VGND.n2563 161.308
R2927 VGND.n2605 VGND.t2696 159.978
R2928 VGND.n2602 VGND.t2699 159.978
R2929 VGND.n2599 VGND.t2694 159.978
R2930 VGND.n2596 VGND.t2689 159.978
R2931 VGND.n2593 VGND.t2695 159.978
R2932 VGND.n2590 VGND.t2702 159.978
R2933 VGND.n2587 VGND.t2698 159.978
R2934 VGND.n2584 VGND.t2692 159.978
R2935 VGND.n2581 VGND.t2688 159.978
R2936 VGND.n2578 VGND.t2690 159.978
R2937 VGND.n2575 VGND.t2701 159.978
R2938 VGND.n2572 VGND.t2693 159.978
R2939 VGND.n2569 VGND.t2700 159.978
R2940 VGND.n2566 VGND.t2697 159.978
R2941 VGND.n2563 VGND.t2703 159.978
R2942 VGND.n123 VGND.t2609 159.315
R2943 VGND.n2216 VGND.t822 159.315
R2944 VGND.n1132 VGND.t686 158.361
R2945 VGND.n2999 VGND.t2005 158.361
R2946 VGND.n121 VGND.t2607 157.291
R2947 VGND.n544 VGND.t820 157.291
R2948 VGND.n68 VGND.t1131 156.915
R2949 VGND.n506 VGND.t1104 156.915
R2950 VGND.n68 VGND.t1132 156.915
R2951 VGND.n506 VGND.t1102 156.915
R2952 VGND.n36 VGND.t542 154.131
R2953 VGND.n123 VGND.t1455 154.131
R2954 VGND.n128 VGND.t1998 154.131
R2955 VGND.n128 VGND.t20 154.131
R2956 VGND.n508 VGND.t2465 154.131
R2957 VGND.n508 VGND.t1127 154.131
R2958 VGND.n2216 VGND.t2160 154.131
R2959 VGND.n541 VGND.t775 154.131
R2960 VGND.n3005 VGND.t876 153.631
R2961 VGND.n60 VGND.t368 153.631
R2962 VGND.n160 VGND.t1129 153.631
R2963 VGND.n2255 VGND.t1101 153.631
R2964 VGND.n2222 VGND.t2264 153.631
R2965 VGND.n1360 VGND.t7 153.631
R2966 VGND.n59 VGND.t1087 152.757
R2967 VGND.n2221 VGND.t1500 152.757
R2968 VGND.n92 VGND.t1136 152.381
R2969 VGND.n2211 VGND.t1099 152.381
R2970 VGND.n2181 VGND.n2180 152.174
R2971 VGND.n167 VGND.t1139 150.922
R2972 VGND.n167 VGND.t1134 150.922
R2973 VGND.n475 VGND.t1103 150.922
R2974 VGND.n475 VGND.t1097 150.922
R2975 VGND.n166 VGND.t1999 150.922
R2976 VGND.n67 VGND.t748 150.922
R2977 VGND.n135 VGND.t1260 150.922
R2978 VGND.n474 VGND.t1941 150.922
R2979 VGND.n2253 VGND.t1294 150.922
R2980 VGND.n505 VGND.t897 150.922
R2981 VGND.n166 VGND.t1421 150.922
R2982 VGND.n67 VGND.t1166 150.922
R2983 VGND.n135 VGND.t1030 150.922
R2984 VGND.n474 VGND.t369 150.922
R2985 VGND.n2253 VGND.t2130 150.922
R2986 VGND.n505 VGND.t413 150.922
R2987 VGND.n3004 VGND.t1977 147.411
R2988 VGND.n159 VGND.t1138 147.411
R2989 VGND.n2254 VGND.t1100 147.411
R2990 VGND.n1359 VGND.t714 147.411
R2991 VGND.n115 VGND.t885 146.964
R2992 VGND.n545 VGND.t1398 146.964
R2993 VGND.n2605 VGND.t1665 143.911
R2994 VGND.n2602 VGND.t1740 143.911
R2995 VGND.n2599 VGND.t1647 143.911
R2996 VGND.n2596 VGND.t1689 143.911
R2997 VGND.n2593 VGND.t1761 143.911
R2998 VGND.n2590 VGND.t1668 143.911
R2999 VGND.n2587 VGND.t1641 143.911
R3000 VGND.n2584 VGND.t1683 143.911
R3001 VGND.n2581 VGND.t1695 143.911
R3002 VGND.n2578 VGND.t1623 143.911
R3003 VGND.n2575 VGND.t1719 143.911
R3004 VGND.n2572 VGND.t1650 143.911
R3005 VGND.n2569 VGND.t1722 143.911
R3006 VGND.n2566 VGND.t1752 143.911
R3007 VGND.n2563 VGND.t1692 143.911
R3008 VGND.n1388 VGND.n806 143.478
R3009 VGND VGND.t2448 142.089
R3010 VGND.n1021 VGND.t1680 119.309
R3011 VGND.n994 VGND.t1716 119.309
R3012 VGND.n2630 VGND.t1677 119.309
R3013 VGND.n204 VGND.t1713 119.309
R3014 VGND.n334 VGND.t1626 119.309
R3015 VGND.n2626 VGND.t1632 119.309
R3016 VGND.n2623 VGND.t1638 119.309
R3017 VGND.n2620 VGND.t1725 119.309
R3018 VGND.n2617 VGND.t1731 119.309
R3019 VGND.n2614 VGND.t1644 119.309
R3020 VGND.n2611 VGND.t1686 119.309
R3021 VGND.n322 VGND.t1701 119.309
R3022 VGND.n315 VGND.t1737 119.309
R3023 VGND.n306 VGND.t1659 119.309
R3024 VGND.n299 VGND.t1704 119.309
R3025 VGND.n2765 VGND.t1743 119.309
R3026 VGND.n290 VGND.t1755 119.309
R3027 VGND.n297 VGND.t1671 119.309
R3028 VGND.n1018 VGND.t1629 119.309
R3029 VGND.n1015 VGND.t1635 119.309
R3030 VGND.n1180 VGND.t1653 119.309
R3031 VGND.n1006 VGND.t1728 119.309
R3032 VGND.n1004 VGND.t1734 119.309
R3033 VGND.n1195 VGND.t1656 119.309
R3034 VGND.n1212 VGND.t1698 119.309
R3035 VGND.n1000 VGND.t1707 119.309
R3036 VGND.n1253 VGND.t1746 119.309
R3037 VGND.n1256 VGND.t1662 119.309
R3038 VGND.n1259 VGND.t1710 119.309
R3039 VGND.n1262 VGND.t1749 119.309
R3040 VGND.n998 VGND.t1758 119.309
R3041 VGND.n1265 VGND.t1674 119.309
R3042 VGND.n5 VGND.n3 117.001
R3043 VGND.t1269 VGND.n5 117.001
R3044 VGND.n6 VGND.n4 117.001
R3045 VGND.n328 VGND.n6 117.001
R3046 VGND.t2242 VGND.t1681 110.535
R3047 VGND.t30 VGND.t632 110.535
R3048 VGND.t1630 VGND.t626 110.535
R3049 VGND.t2335 VGND.t665 110.535
R3050 VGND.t2327 VGND.t1636 110.535
R3051 VGND.t1612 VGND.t2320 110.535
R3052 VGND.t1654 VGND.t2305 110.535
R3053 VGND.t2218 VGND.t1162 110.535
R3054 VGND.t2230 VGND.t1729 110.535
R3055 VGND.t150 VGND.t620 110.535
R3056 VGND.t1735 VGND.t604 110.535
R3057 VGND.t2308 VGND.t2685 110.535
R3058 VGND.t591 VGND.t1657 110.535
R3059 VGND.t14 VGND.t2233 110.535
R3060 VGND.t1699 VGND.t2224 110.535
R3061 VGND.t2208 VGND.t1159 110.535
R3062 VGND.t2202 VGND.t1708 110.535
R3063 VGND.t188 VGND.t593 110.535
R3064 VGND.t1747 VGND.t606 110.535
R3065 VGND.t2309 VGND.t230 110.535
R3066 VGND.t2293 VGND.t1663 110.535
R3067 VGND.t35 VGND.t2205 110.535
R3068 VGND.t1711 VGND.t2284 110.535
R3069 VGND.t2193 VGND.t2167 110.535
R3070 VGND.t587 VGND.t1750 110.535
R3071 VGND.t2519 VGND.t580 110.535
R3072 VGND.t1759 VGND.t575 110.535
R3073 VGND.t2286 VGND.t8 110.535
R3074 VGND.t2336 VGND.t1675 110.535
R3075 VGND.t543 VGND.t2265 110.535
R3076 VGND.t1717 VGND.t2189 110.535
R3077 VGND.t577 VGND.t149 110.535
R3078 VGND.t1389 VGND.t1399 92.4699
R3079 VGND.t1399 VGND.t1396 92.4699
R3080 VGND.t1396 VGND.t1400 92.4699
R3081 VGND.t1400 VGND.t62 92.4699
R3082 VGND.t62 VGND.t76 92.4699
R3083 VGND.t76 VGND.t2357 92.4699
R3084 VGND.t2357 VGND.t1289 92.4699
R3085 VGND VGND.n806 80.9529
R3086 VGND VGND.n806 75.1009
R3087 VGND.n1337 VGND 74.8566
R3088 VGND.t1289 VGND 70.4533
R3089 VGND.n2285 VGND 58.8055
R3090 VGND.n2284 VGND 58.8055
R3091 VGND.n2250 VGND 58.8055
R3092 VGND.n2248 VGND 58.8055
R3093 VGND.n1386 VGND 58.8055
R3094 VGND.n2348 VGND.n2347 53.1823
R3095 VGND.n2349 VGND.n2348 53.1823
R3096 VGND.n3021 VGND.n3020 53.1823
R3097 VGND.n3020 VGND.n3019 53.1823
R3098 VGND.t892 VGND.t2446 50.5752
R3099 VGND.t888 VGND.t2420 50.5752
R3100 VGND.t882 VGND.t2457 50.5752
R3101 VGND.t884 VGND.t2397 50.5752
R3102 VGND.t1397 VGND.t469 50.5752
R3103 VGND.t1394 VGND.t74 50.5752
R3104 VGND.t1392 VGND.t1323 50.5752
R3105 VGND.t1390 VGND.t2258 50.5752
R3106 VGND VGND.n2981 43.2063
R3107 VGND VGND.n18 43.2063
R3108 VGND VGND.n2951 43.2063
R3109 VGND VGND.n44 43.2063
R3110 VGND.n2347 VGND.n2346 40.6593
R3111 VGND.n886 VGND.t2207 34.8005
R3112 VGND.n886 VGND.t597 34.8005
R3113 VGND.n889 VGND.t595 34.8005
R3114 VGND.n889 VGND.t2299 34.8005
R3115 VGND.n893 VGND.t2296 34.8005
R3116 VGND.n893 VGND.t2210 34.8005
R3117 VGND.n930 VGND.t2274 34.8005
R3118 VGND.n930 VGND.t2188 34.8005
R3119 VGND.n935 VGND.t590 34.8005
R3120 VGND.n935 VGND.t586 34.8005
R3121 VGND.n940 VGND.t579 34.8005
R3122 VGND.n940 VGND.t2280 34.8005
R3123 VGND.n945 VGND.t2343 34.8005
R3124 VGND.n945 VGND.t2269 34.8005
R3125 VGND.n950 VGND.t2192 34.8005
R3126 VGND.n950 VGND.t582 34.8005
R3127 VGND.n955 VGND.t2171 34.8005
R3128 VGND.n955 VGND.t2347 34.8005
R3129 VGND.n960 VGND.t2339 34.8005
R3130 VGND.n960 VGND.t2282 34.8005
R3131 VGND.n965 VGND.t2252 34.8005
R3132 VGND.n965 VGND.t2175 34.8005
R3133 VGND.n970 VGND.t2239 34.8005
R3134 VGND.n970 VGND.t630 34.8005
R3135 VGND.n975 VGND.t614 34.8005
R3136 VGND.n975 VGND.t2254 34.8005
R3137 VGND.n980 VGND.t2322 34.8005
R3138 VGND.n980 VGND.t2241 34.8005
R3139 VGND.n985 VGND.t2221 34.8005
R3140 VGND.n985 VGND.t2216 34.8005
R3141 VGND.n996 VGND.t2278 34.8005
R3142 VGND.n996 VGND.t2190 34.8005
R3143 VGND.n1273 VGND.t2345 34.8005
R3144 VGND.n1273 VGND.t2337 34.8005
R3145 VGND.n1230 VGND.t2186 34.8005
R3146 VGND.n1230 VGND.t576 34.8005
R3147 VGND.n1229 VGND.t2267 34.8005
R3148 VGND.n1229 VGND.t588 34.8005
R3149 VGND.n1226 VGND.t2356 34.8005
R3150 VGND.n1226 VGND.t2285 34.8005
R3151 VGND.n1224 VGND.t584 34.8005
R3152 VGND.n1224 VGND.t2294 34.8005
R3153 VGND.n1221 VGND.t2196 34.8005
R3154 VGND.n1221 VGND.t607 34.8005
R3155 VGND.n1216 VGND.t2292 34.8005
R3156 VGND.n1216 VGND.t2203 34.8005
R3157 VGND.n1002 VGND.t2312 34.8005
R3158 VGND.n1002 VGND.t2225 34.8005
R3159 VGND.n1203 VGND.t2201 34.8005
R3160 VGND.n1203 VGND.t592 34.8005
R3161 VGND.n1007 VGND.t2223 34.8005
R3162 VGND.n1007 VGND.t605 34.8005
R3163 VGND.n1184 VGND.t2235 34.8005
R3164 VGND.n1184 VGND.t2231 34.8005
R3165 VGND.n1010 VGND.t601 34.8005
R3166 VGND.n1010 VGND.t2306 34.8005
R3167 VGND.n1171 VGND.t625 34.8005
R3168 VGND.n1171 VGND.t2328 34.8005
R3169 VGND.n1012 VGND.t2237 34.8005
R3170 VGND.n1012 VGND.t627 34.8005
R3171 VGND.n329 VGND.t2272 34.8005
R3172 VGND.n329 VGND.t2184 34.8005
R3173 VGND.n332 VGND.t2182 34.8005
R3174 VGND.n332 VGND.t2354 34.8005
R3175 VGND.n356 VGND.t2352 34.8005
R3176 VGND.n356 VGND.t2276 34.8005
R3177 VGND.n363 VGND.t2330 34.8005
R3178 VGND.n363 VGND.t2246 34.8005
R3179 VGND.n366 VGND.t2180 34.8005
R3180 VGND.n366 VGND.t2177 34.8005
R3181 VGND.n374 VGND.t2169 34.8005
R3182 VGND.n374 VGND.t2332 34.8005
R3183 VGND.n377 VGND.t616 34.8005
R3184 VGND.n377 VGND.t2318 34.8005
R3185 VGND.n385 VGND.t2250 34.8005
R3186 VGND.n385 VGND.t2173 34.8005
R3187 VGND.n324 VGND.t2227 34.8005
R3188 VGND.n324 VGND.t618 34.8005
R3189 VGND.n313 VGND.t612 34.8005
R3190 VGND.n313 VGND.t2334 34.8005
R3191 VGND.n308 VGND.t2314 34.8005
R3192 VGND.n308 VGND.t2229 34.8005
R3193 VGND.n310 VGND.t2302 34.8005
R3194 VGND.n310 VGND.t2214 34.8005
R3195 VGND.n2729 VGND.t2198 34.8005
R3196 VGND.n2729 VGND.t2316 34.8005
R3197 VGND.n292 VGND.t599 34.8005
R3198 VGND.n292 VGND.t2304 34.8005
R3199 VGND.n295 VGND.t2290 34.8005
R3200 VGND.n295 VGND.t2288 34.8005
R3201 VGND.n202 VGND.t2212 34.8005
R3202 VGND.n202 VGND.t603 34.8005
R3203 VGND.n395 VGND.t1667 34.8005
R3204 VGND.n395 VGND.t1935 34.8005
R3205 VGND.n2637 VGND.t142 34.8005
R3206 VGND.n2637 VGND.t1925 34.8005
R3207 VGND.n2642 VGND.t1814 34.8005
R3208 VGND.n2642 VGND.t1216 34.8005
R3209 VGND.n2647 VGND.t1566 34.8005
R3210 VGND.n2647 VGND.t1214 34.8005
R3211 VGND.n2652 VGND.t924 34.8005
R3212 VGND.n2652 VGND.t1933 34.8005
R3213 VGND.n2657 VGND.t1950 34.8005
R3214 VGND.n2657 VGND.t2636 34.8005
R3215 VGND.n2662 VGND.t1262 34.8005
R3216 VGND.n2662 VGND.t2634 34.8005
R3217 VGND.n2667 VGND.t2039 34.8005
R3218 VGND.n2667 VGND.t1931 34.8005
R3219 VGND.n392 VGND.t783 34.8005
R3220 VGND.n392 VGND.t1929 34.8005
R3221 VGND.n2713 VGND.t1069 34.8005
R3222 VGND.n2713 VGND.t2638 34.8005
R3223 VGND.n318 VGND.t490 34.8005
R3224 VGND.n318 VGND.t1212 34.8005
R3225 VGND.n2746 VGND.t2153 34.8005
R3226 VGND.n2746 VGND.t1210 34.8005
R3227 VGND.n302 VGND.t679 34.8005
R3228 VGND.n302 VGND.t2632 34.8005
R3229 VGND.n2751 VGND.t308 34.8005
R3230 VGND.n2751 VGND.t1220 34.8005
R3231 VGND.n2786 VGND.t1535 34.8005
R3232 VGND.n2786 VGND.t1218 34.8005
R3233 VGND.n285 VGND.t476 34.8005
R3234 VGND.n285 VGND.t1927 34.8005
R3235 VGND.n399 VGND.t1742 34.8005
R3236 VGND.n399 VGND.t2134 34.8005
R3237 VGND.n2341 VGND.t187 34.8005
R3238 VGND.n2341 VGND.t2545 34.8005
R3239 VGND.n2336 VGND.t229 34.8005
R3240 VGND.n2336 VGND.t206 34.8005
R3241 VGND.n2331 VGND.t1569 34.8005
R3242 VGND.n2331 VGND.t204 34.8005
R3243 VGND.n2326 VGND.t294 34.8005
R3244 VGND.n2326 VGND.t2132 34.8005
R3245 VGND.n2321 VGND.t1320 34.8005
R3246 VGND.n2321 VGND.t2559 34.8005
R3247 VGND.n2316 VGND.t1234 34.8005
R3248 VGND.n2316 VGND.t2557 34.8005
R3249 VGND.n2311 VGND.t351 34.8005
R3250 VGND.n2311 VGND.t2551 34.8005
R3251 VGND.n2306 VGND.t365 34.8005
R3252 VGND.n2306 VGND.t2549 34.8005
R3253 VGND.n2301 VGND.t770 34.8005
R3254 VGND.n2301 VGND.t2561 34.8005
R3255 VGND.n2296 VGND.t533 34.8005
R3256 VGND.n2296 VGND.t2138 34.8005
R3257 VGND.n2291 VGND.t1095 34.8005
R3258 VGND.n2291 VGND.t2136 34.8005
R3259 VGND.n2286 VGND.t2614 34.8005
R3260 VGND.n2286 VGND.t2555 34.8005
R3261 VGND.n413 VGND.t122 34.8005
R3262 VGND.n413 VGND.t2553 34.8005
R3263 VGND.n2539 VGND.t1922 34.8005
R3264 VGND.n2539 VGND.t208 34.8005
R3265 VGND.n416 VGND.t13 34.8005
R3266 VGND.n416 VGND.t2547 34.8005
R3267 VGND.n468 VGND.t1649 34.8005
R3268 VGND.n468 VGND.t1333 34.8005
R3269 VGND.n470 VGND.t761 34.8005
R3270 VGND.n470 VGND.t838 34.8005
R3271 VGND.n2375 VGND.t703 34.8005
R3272 VGND.n2375 VGND.t2083 34.8005
R3273 VGND.n458 VGND.t2470 34.8005
R3274 VGND.n458 VGND.t1339 34.8005
R3275 VGND.n2401 VGND.t931 34.8005
R3276 VGND.n2401 VGND.t223 34.8005
R3277 VGND.n450 VGND.t2078 34.8005
R3278 VGND.n450 VGND.t834 34.8005
R3279 VGND.n2427 VGND.t1268 34.8005
R3280 VGND.n2427 VGND.t832 34.8005
R3281 VGND.n442 VGND.t2045 34.8005
R3282 VGND.n442 VGND.t221 34.8005
R3283 VGND.n2453 VGND.t1448 34.8005
R3284 VGND.n2453 VGND.t219 34.8005
R3285 VGND.n434 VGND.t710 34.8005
R3286 VGND.n434 VGND.t836 34.8005
R3287 VGND.n2479 VGND.t444 34.8005
R3288 VGND.n2479 VGND.t1337 34.8005
R3289 VGND.n426 VGND.t536 34.8005
R3290 VGND.n426 VGND.t1335 34.8005
R3291 VGND.n2510 VGND.t1409 34.8005
R3292 VGND.n2510 VGND.t830 34.8005
R3293 VGND.n2515 VGND.t314 34.8005
R3294 VGND.n2515 VGND.t2087 34.8005
R3295 VGND.n2520 VGND.t1527 34.8005
R3296 VGND.n2520 VGND.t2085 34.8005
R3297 VGND.n418 VGND.t483 34.8005
R3298 VGND.n418 VGND.t217 34.8005
R3299 VGND.n465 VGND.t1691 34.8005
R3300 VGND.n465 VGND.t2523 34.8005
R3301 VGND.n2362 VGND.t47 34.8005
R3302 VGND.n2362 VGND.t1889 34.8005
R3303 VGND.n462 VGND.t2098 34.8005
R3304 VGND.n462 VGND.t2140 34.8005
R3305 VGND.n2388 VGND.t2592 34.8005
R3306 VGND.n2388 VGND.t2529 34.8005
R3307 VGND.n454 VGND.t909 34.8005
R3308 VGND.n454 VGND.t2019 34.8005
R3309 VGND.n2414 VGND.t1808 34.8005
R3310 VGND.n2414 VGND.t1885 34.8005
R3311 VGND.n446 VGND.t1620 34.8005
R3312 VGND.n446 VGND.t1883 34.8005
R3313 VGND.n2440 VGND.t2541 34.8005
R3314 VGND.n2440 VGND.t2017 34.8005
R3315 VGND.n438 VGND.t375 34.8005
R3316 VGND.n438 VGND.t2015 34.8005
R3317 VGND.n2466 VGND.t905 34.8005
R3318 VGND.n2466 VGND.t1887 34.8005
R3319 VGND.n430 VGND.t456 34.8005
R3320 VGND.n430 VGND.t2527 34.8005
R3321 VGND.n2492 VGND.t340 34.8005
R3322 VGND.n2492 VGND.t2525 34.8005
R3323 VGND.n422 VGND.t107 34.8005
R3324 VGND.n422 VGND.t2146 34.8005
R3325 VGND.n2497 VGND.t298 34.8005
R3326 VGND.n2497 VGND.t2144 34.8005
R3327 VGND.n2808 VGND.t726 34.8005
R3328 VGND.n2808 VGND.t2142 34.8005
R3329 VGND.n276 VGND.t328 34.8005
R3330 VGND.n276 VGND.t2013 34.8005
R3331 VGND.n624 VGND.t1763 34.8005
R3332 VGND.n624 VGND.t2627 34.8005
R3333 VGND.n1909 VGND.t1064 34.8005
R3334 VGND.n1909 VGND.t59 34.8005
R3335 VGND.n621 VGND.t1989 34.8005
R3336 VGND.n621 VGND.t96 34.8005
R3337 VGND.n1920 VGND.t2599 34.8005
R3338 VGND.n1920 VGND.t2488 34.8005
R3339 VGND.n618 VGND.t287 34.8005
R3340 VGND.n618 VGND.t2625 34.8005
R3341 VGND.n1931 VGND.t1915 34.8005
R3342 VGND.n1931 VGND.t55 34.8005
R3343 VGND.n615 VGND.t1230 34.8005
R3344 VGND.n615 VGND.t53 34.8005
R3345 VGND.n1942 VGND.t348 34.8005
R3346 VGND.n1942 VGND.t2623 34.8005
R3347 VGND.n612 VGND.t1470 34.8005
R3348 VGND.n612 VGND.t2621 34.8005
R3349 VGND.n1953 VGND.t148 34.8005
R3350 VGND.n1953 VGND.t57 34.8005
R3351 VGND.n609 VGND.t528 34.8005
R3352 VGND.n609 VGND.t2486 34.8005
R3353 VGND.n1964 VGND.t1091 34.8005
R3354 VGND.n1964 VGND.t2484 34.8005
R3355 VGND.n606 VGND.t1610 34.8005
R3356 VGND.n606 VGND.t51 34.8005
R3357 VGND.n1975 VGND.t116 34.8005
R3358 VGND.n1975 VGND.t100 34.8005
R3359 VGND.n1980 VGND.t1124 34.8005
R3360 VGND.n1980 VGND.t98 34.8005
R3361 VGND.n605 VGND.t1983 34.8005
R3362 VGND.n605 VGND.t61 34.8005
R3363 VGND.n589 VGND.t1670 34.8005
R3364 VGND.n589 VGND.t2025 34.8005
R3365 VGND.n595 VGND.t140 34.8005
R3366 VGND.n595 VGND.t1601 34.8005
R3367 VGND.n592 VGND.t1812 34.8005
R3368 VGND.n592 VGND.t2033 34.8005
R3369 VGND.n2054 VGND.t1563 34.8005
R3370 VGND.n2054 VGND.t2031 34.8005
R3371 VGND.n2049 VGND.t922 34.8005
R3372 VGND.n2049 VGND.t2023 34.8005
R3373 VGND.n2044 VGND.t1948 34.8005
R3374 VGND.n2044 VGND.t426 34.8005
R3375 VGND.n2039 VGND.t1772 34.8005
R3376 VGND.n2039 VGND.t424 34.8005
R3377 VGND.n2034 VGND.t2037 34.8005
R3378 VGND.n2034 VGND.t2021 34.8005
R3379 VGND.n2029 VGND.t781 34.8005
R3380 VGND.n2029 VGND.t1605 34.8005
R3381 VGND.n2024 VGND.t1067 34.8005
R3382 VGND.n2024 VGND.t428 34.8005
R3383 VGND.n2019 VGND.t487 34.8005
R3384 VGND.n2019 VGND.t2029 34.8005
R3385 VGND.n2014 VGND.t2151 34.8005
R3386 VGND.n2014 VGND.t2027 34.8005
R3387 VGND.n2009 VGND.t676 34.8005
R3388 VGND.n2009 VGND.t422 34.8005
R3389 VGND.n2004 VGND.t306 34.8005
R3390 VGND.n2004 VGND.t420 34.8005
R3391 VGND.n600 VGND.t1532 34.8005
R3392 VGND.n600 VGND.t418 34.8005
R3393 VGND.n1993 VGND.t474 34.8005
R3394 VGND.n1993 VGND.t1603 34.8005
R3395 VGND.n586 VGND.t1643 34.8005
R3396 VGND.n586 VGND.t518 34.8005
R3397 VGND.n2068 VGND.t763 34.8005
R3398 VGND.n2068 VGND.t508 34.8005
R3399 VGND.n2073 VGND.t705 34.8005
R3400 VGND.n2073 VGND.t556 34.8005
R3401 VGND.n2078 VGND.t2468 34.8005
R3402 VGND.n2078 VGND.t524 34.8005
R3403 VGND.n2083 VGND.t933 34.8005
R3404 VGND.n2083 VGND.t516 34.8005
R3405 VGND.n2088 VGND.t2080 34.8005
R3406 VGND.n2088 VGND.t504 34.8005
R3407 VGND.n2093 VGND.t1380 34.8005
R3408 VGND.n2093 VGND.t502 34.8005
R3409 VGND.n2098 VGND.t2047 34.8005
R3410 VGND.n2098 VGND.t514 34.8005
R3411 VGND.n2103 VGND.t1450 34.8005
R3412 VGND.n2103 VGND.t512 34.8005
R3413 VGND.n2108 VGND.t712 34.8005
R3414 VGND.n2108 VGND.t506 34.8005
R3415 VGND.n2113 VGND.t446 34.8005
R3416 VGND.n2113 VGND.t522 34.8005
R3417 VGND.n2118 VGND.t538 34.8005
R3418 VGND.n2118 VGND.t520 34.8005
R3419 VGND.n583 VGND.t1411 34.8005
R3420 VGND.n583 VGND.t500 34.8005
R3421 VGND.n2123 VGND.t316 34.8005
R3422 VGND.n2123 VGND.t560 34.8005
R3423 VGND.n2833 VGND.t1529 34.8005
R3424 VGND.n2833 VGND.t558 34.8005
R3425 VGND.n264 VGND.t485 34.8005
R3426 VGND.n264 VGND.t510 34.8005
R3427 VGND.n546 VGND.t1685 34.8005
R3428 VGND.n546 VGND.t1013 34.8005
R3429 VGND.n549 VGND.t49 34.8005
R3430 VGND.n549 VGND.t202 34.8005
R3431 VGND.n1755 VGND.t2100 34.8005
R3432 VGND.n1755 VGND.t690 34.8005
R3433 VGND.n1760 VGND.t2590 34.8005
R3434 VGND.n1760 VGND.t688 34.8005
R3435 VGND.n1751 VGND.t911 34.8005
R3436 VGND.n1751 VGND.t1025 34.8005
R3437 VGND.n1771 VGND.t215 34.8005
R3438 VGND.n1771 VGND.t1792 34.8005
R3439 VGND.n1748 VGND.t1622 34.8005
R3440 VGND.n1748 VGND.t1790 34.8005
R3441 VGND.n1782 VGND.t2543 34.8005
R3442 VGND.n1782 VGND.t1023 34.8005
R3443 VGND.n1745 VGND.t377 34.8005
R3444 VGND.n1745 VGND.t1021 34.8005
R3445 VGND.n1793 VGND.t907 34.8005
R3446 VGND.n1793 VGND.t1794 34.8005
R3447 VGND.n1742 VGND.t458 34.8005
R3448 VGND.n1742 VGND.t1017 34.8005
R3449 VGND.n1804 VGND.t638 34.8005
R3450 VGND.n1804 VGND.t1015 34.8005
R3451 VGND.n1739 VGND.t109 34.8005
R3452 VGND.n1739 VGND.t1788 34.8005
R3453 VGND.n1815 VGND.t300 34.8005
R3454 VGND.n1815 VGND.t694 34.8005
R3455 VGND.n1820 VGND.t728 34.8005
R3456 VGND.n1820 VGND.t692 34.8005
R3457 VGND.n1738 VGND.t330 34.8005
R3458 VGND.n1738 VGND.t1019 34.8005
R3459 VGND.n627 VGND.t1697 34.8005
R3460 VGND.n627 VGND.t1052 34.8005
R3461 VGND.n1677 VGND.t42 34.8005
R3462 VGND.n1677 VGND.t1042 34.8005
R3463 VGND.n1674 VGND.t2092 34.8005
R3464 VGND.n1674 VGND.t1112 34.8005
R3465 VGND.n1688 VGND.t2596 34.8005
R3466 VGND.n1688 VGND.t1110 34.8005
R3467 VGND.n1693 VGND.t1515 34.8005
R3468 VGND.n1693 VGND.t1050 34.8005
R3469 VGND.n1698 VGND.t1802 34.8005
R3470 VGND.n1698 VGND.t1038 34.8005
R3471 VGND.n1703 VGND.t1618 34.8005
R3472 VGND.n1703 VGND.t2011 34.8005
R3473 VGND.n1708 VGND.t2537 34.8005
R3474 VGND.n1708 VGND.t554 34.8005
R3475 VGND.n1713 VGND.t371 34.8005
R3476 VGND.n1713 VGND.t552 34.8005
R3477 VGND.n1718 VGND.t1151 34.8005
R3478 VGND.n1718 VGND.t1040 34.8005
R3479 VGND.n1723 VGND.t454 34.8005
R3480 VGND.n1723 VGND.t1056 34.8005
R3481 VGND.n1728 VGND.t338 34.8005
R3482 VGND.n1728 VGND.t1054 34.8005
R3483 VGND.n1671 VGND.t105 34.8005
R3484 VGND.n1671 VGND.t2009 34.8005
R3485 VGND.n1844 VGND.t723 34.8005
R3486 VGND.n1844 VGND.t2007 34.8005
R3487 VGND.n1733 VGND.t815 34.8005
R3488 VGND.n1733 VGND.t1114 34.8005
R3489 VGND.n1833 VGND.t326 34.8005
R3490 VGND.n1833 VGND.t1044 34.8005
R3491 VGND.n631 VGND.t1625 34.8005
R3492 VGND.n631 VGND.t871 34.8005
R3493 VGND.n668 VGND.t1062 34.8005
R3494 VGND.n668 VGND.t1184 34.8005
R3495 VGND.n673 VGND.t1987 34.8005
R3496 VGND.n673 VGND.t1881 34.8005
R3497 VGND.n678 VGND.t2601 34.8005
R3498 VGND.n678 VGND.t1879 34.8005
R3499 VGND.n683 VGND.t919 34.8005
R3500 VGND.n683 VGND.t869 34.8005
R3501 VGND.n688 VGND.t1824 34.8005
R3502 VGND.n688 VGND.t1180 34.8005
R3503 VGND.n693 VGND.t1386 34.8005
R3504 VGND.n693 VGND.t1178 34.8005
R3505 VGND.n698 VGND.t346 34.8005
R3506 VGND.n698 VGND.t867 34.8005
R3507 VGND.n703 VGND.t1468 34.8005
R3508 VGND.n703 VGND.t865 34.8005
R3509 VGND.n708 VGND.t146 34.8005
R3510 VGND.n708 VGND.t1182 34.8005
R3511 VGND.n713 VGND.t526 34.8005
R3512 VGND.n713 VGND.t1877 34.8005
R3513 VGND.n718 VGND.t1089 34.8005
R3514 VGND.n718 VGND.t1875 34.8005
R3515 VGND.n665 VGND.t1608 34.8005
R3516 VGND.n665 VGND.t1176 34.8005
R3517 VGND.n723 VGND.t114 34.8005
R3518 VGND.n723 VGND.t1174 34.8005
R3519 VGND.n2858 VGND.t212 34.8005
R3520 VGND.n2858 VGND.t1172 34.8005
R3521 VGND.n252 VGND.t1981 34.8005
R3522 VGND.n252 VGND.t863 34.8005
R3523 VGND.n878 VGND.t1721 34.8005
R3524 VGND.n878 VGND.t1432 34.8005
R3525 VGND.n1351 VGND.t847 34.8005
R3526 VGND.n1351 VGND.t1360 34.8005
R3527 VGND.n873 VGND.t1956 34.8005
R3528 VGND.n873 VGND.t1440 34.8005
R3529 VGND.n807 VGND.t569 34.8005
R3530 VGND.n807 VGND.t1438 34.8005
R3531 VGND.n809 VGND.t1509 34.8005
R3532 VGND.n809 VGND.t1430 34.8005
R3533 VGND.n822 VGND.t1800 34.8005
R3534 VGND.n822 VGND.t1356 34.8005
R3535 VGND.n827 VGND.t1224 34.8005
R3536 VGND.n827 VGND.t1354 34.8005
R3537 VGND.n832 VGND.t359 34.8005
R3538 VGND.n832 VGND.t2521 34.8005
R3539 VGND.n837 VGND.t382 34.8005
R3540 VGND.n837 VGND.t1364 34.8005
R3541 VGND.n842 VGND.t234 34.8005
R3542 VGND.n842 VGND.t1358 34.8005
R3543 VGND.n847 VGND.t436 34.8005
R3544 VGND.n847 VGND.t1436 34.8005
R3545 VGND.n818 VGND.t2166 34.8005
R3546 VGND.n818 VGND.t1434 34.8005
R3547 VGND.n852 VGND.t2478 34.8005
R3548 VGND.n852 VGND.t1352 34.8005
R3549 VGND.n733 VGND.t390 34.8005
R3550 VGND.n733 VGND.t1350 34.8005
R3551 VGND.n1660 VGND.t674 34.8005
R3552 VGND.n1660 VGND.t1442 34.8005
R3553 VGND.n736 VGND.t318 34.8005
R3554 VGND.n736 VGND.t1362 34.8005
R3555 VGND.n799 VGND.t1652 34.8005
R3556 VGND.n799 VGND.t401 34.8005
R3557 VGND.n1389 VGND.t759 34.8005
R3558 VGND.n1389 VGND.t853 34.8005
R3559 VGND.n1394 VGND.t701 34.8005
R3560 VGND.n1394 VGND.t409 34.8005
R3561 VGND.n803 VGND.t2472 34.8005
R3562 VGND.n803 VGND.t407 34.8005
R3563 VGND.n1489 VGND.t929 34.8005
R3564 VGND.n1489 VGND.t861 34.8005
R3565 VGND.n775 VGND.t2076 34.8005
R3566 VGND.n775 VGND.t849 34.8005
R3567 VGND.n1515 VGND.t1266 34.8005
R3568 VGND.n1515 VGND.t2464 34.8005
R3569 VGND.n767 VGND.t2043 34.8005
R3570 VGND.n767 VGND.t859 34.8005
R3571 VGND.n1541 VGND.t1446 34.8005
R3572 VGND.n1541 VGND.t857 34.8005
R3573 VGND.n1546 VGND.t708 34.8005
R3574 VGND.n1546 VGND.t851 34.8005
R3575 VGND.n759 VGND.t494 34.8005
R3576 VGND.n759 VGND.t405 34.8005
R3577 VGND.n1551 VGND.t2157 34.8005
R3578 VGND.n1551 VGND.t403 34.8005
R3579 VGND.n1631 VGND.t1407 34.8005
R3580 VGND.n1631 VGND.t2462 34.8005
R3581 VGND.n1636 VGND.t312 34.8005
R3582 VGND.n1636 VGND.t2617 34.8005
R3583 VGND.n1641 VGND.t1525 34.8005
R3584 VGND.n1641 VGND.t411 34.8005
R3585 VGND.n739 VGND.t481 34.8005
R3586 VGND.n739 VGND.t855 34.8005
R3587 VGND.n796 VGND.t1724 34.8005
R3588 VGND.n796 VGND.t2640 34.8005
R3589 VGND.n1409 VGND.t845 34.8005
R3590 VGND.n1409 VGND.t1458 34.8005
R3591 VGND.n793 VGND.t1954 34.8005
R3592 VGND.n793 VGND.t2648 34.8005
R3593 VGND.n1476 VGND.t571 34.8005
R3594 VGND.n1476 VGND.t2646 34.8005
R3595 VGND.n779 VGND.t915 34.8005
R3596 VGND.n779 VGND.t1466 34.8005
R3597 VGND.n1502 VGND.t1798 34.8005
R3598 VGND.n1502 VGND.t132 34.8005
R3599 VGND.n771 VGND.t1222 34.8005
R3600 VGND.n771 VGND.t130 34.8005
R3601 VGND.n1528 VGND.t357 34.8005
R3602 VGND.n1528 VGND.t1464 34.8005
R3603 VGND.n763 VGND.t380 34.8005
R3604 VGND.n763 VGND.t1462 34.8005
R3605 VGND.n1565 VGND.t232 34.8005
R3606 VGND.n1565 VGND.t134 34.8005
R3607 VGND.n754 VGND.t434 34.8005
R3608 VGND.n754 VGND.t2644 34.8005
R3609 VGND.n1580 VGND.t2164 34.8005
R3610 VGND.n1580 VGND.t2642 34.8005
R3611 VGND.n1575 VGND.t1819 34.8005
R3612 VGND.n1575 VGND.t128 34.8005
R3613 VGND.n1570 VGND.t388 34.8005
R3614 VGND.n1570 VGND.t126 34.8005
R3615 VGND.n2883 VGND.t672 34.8005
R3616 VGND.n2883 VGND.t124 34.8005
R3617 VGND.n239 VGND.t344 34.8005
R3618 VGND.n239 VGND.t1460 34.8005
R3619 VGND.n881 VGND.t1754 34.8005
R3620 VGND.n881 VGND.t2654 34.8005
R3621 VGND.n883 VGND.t185 34.8005
R3622 VGND.n883 VGND.t89 34.8005
R3623 VGND.n1422 VGND.t227 34.8005
R3624 VGND.n1422 VGND.t1344 34.8005
R3625 VGND.n1427 VGND.t1572 34.8005
R3626 VGND.n1427 VGND.t2660 34.8005
R3627 VGND.n1432 VGND.t291 34.8005
R3628 VGND.n1432 VGND.t2652 34.8005
R3629 VGND.n1437 VGND.t1919 34.8005
R3630 VGND.n1437 VGND.t85 34.8005
R3631 VGND.n1442 VGND.t1232 34.8005
R3632 VGND.n1442 VGND.t83 34.8005
R3633 VGND.n1447 VGND.t778 34.8005
R3634 VGND.n1447 VGND.t2650 34.8005
R3635 VGND.n1452 VGND.t363 34.8005
R3636 VGND.n1452 VGND.t93 34.8005
R3637 VGND.n789 VGND.t768 34.8005
R3638 VGND.n789 VGND.t87 34.8005
R3639 VGND.n1457 VGND.t530 34.8005
R3640 VGND.n1457 VGND.t2658 34.8005
R3641 VGND.n1594 VGND.t1093 34.8005
R3642 VGND.n1594 VGND.t2656 34.8005
R3643 VGND.n1599 VGND.t2611 34.8005
R3644 VGND.n1599 VGND.t81 34.8005
R3645 VGND.n748 VGND.t120 34.8005
R3646 VGND.n748 VGND.t1348 34.8005
R3647 VGND.n1612 VGND.t1126 34.8005
R3648 VGND.n1612 VGND.t1346 34.8005
R3649 VGND.n1604 VGND.t10 34.8005
R3650 VGND.n1604 VGND.t91 34.8005
R3651 VGND.n1023 VGND.t1694 34.8005
R3652 VGND.n1023 VGND.t170 34.8005
R3653 VGND.n1030 VGND.t44 34.8005
R3654 VGND.n1030 VGND.t161 34.8005
R3655 VGND.n1035 VGND.t2094 34.8005
R3656 VGND.n1035 VGND.t1995 34.8005
R3657 VGND.n1027 VGND.t2594 34.8005
R3658 VGND.n1027 VGND.t1993 34.8005
R3659 VGND.n1093 VGND.t1517 34.8005
R3660 VGND.n1093 VGND.t168 34.8005
R3661 VGND.n1088 VGND.t1804 34.8005
R3662 VGND.n1088 VGND.t1969 34.8005
R3663 VGND.n1083 VGND.t1616 34.8005
R3664 VGND.n1083 VGND.t1967 34.8005
R3665 VGND.n1078 VGND.t2535 34.8005
R3666 VGND.n1078 VGND.t166 34.8005
R3667 VGND.n1073 VGND.t735 34.8005
R3668 VGND.n1073 VGND.t1973 34.8005
R3669 VGND.n1040 VGND.t1149 34.8005
R3670 VGND.n1040 VGND.t1971 34.8005
R3671 VGND.n1042 VGND.t452 34.8005
R3672 VGND.n1042 VGND.t1991 34.8005
R3673 VGND.n1051 VGND.t336 34.8005
R3674 VGND.n1051 VGND.t172 34.8005
R3675 VGND.n1056 VGND.t2482 34.8005
R3676 VGND.n1056 VGND.t1965 34.8005
R3677 VGND.n1047 VGND.t721 34.8005
R3678 VGND.n1047 VGND.t1963 34.8005
R3679 VGND.n2903 VGND.t817 34.8005
R3680 VGND.n2903 VGND.t1997 34.8005
R3681 VGND.n227 VGND.t324 34.8005
R3682 VGND.n227 VGND.t163 34.8005
R3683 VGND.n1013 VGND.t2324 34.8005
R3684 VGND.n1013 VGND.t2243 34.8005
R3685 VGND.n926 VGND.t623 34.8005
R3686 VGND.n926 VGND.t2326 34.8005
R3687 VGND.n105 VGND.n103 34.6358
R3688 VGND.n2984 VGND.n2978 34.6358
R3689 VGND.n2987 VGND.n2986 34.6358
R3690 VGND.n2987 VGND.n2974 34.6358
R3691 VGND.n2991 VGND.n2974 34.6358
R3692 VGND.n2992 VGND.n2991 34.6358
R3693 VGND.n2993 VGND.n2992 34.6358
R3694 VGND.n21 VGND.n20 34.6358
R3695 VGND.n23 VGND.n12 34.6358
R3696 VGND.n27 VGND.n12 34.6358
R3697 VGND.n28 VGND.n27 34.6358
R3698 VGND.n29 VGND.n28 34.6358
R3699 VGND.n29 VGND.n9 34.6358
R3700 VGND.n3006 VGND.n10 34.6358
R3701 VGND.n181 VGND.n180 34.6358
R3702 VGND.n185 VGND.n184 34.6358
R3703 VGND.n2954 VGND.n2953 34.6358
R3704 VGND.n2956 VGND.n2947 34.6358
R3705 VGND.n2960 VGND.n2947 34.6358
R3706 VGND.n2961 VGND.n2960 34.6358
R3707 VGND.n2962 VGND.n2961 34.6358
R3708 VGND.n2962 VGND.n2945 34.6358
R3709 VGND.n47 VGND.n46 34.6358
R3710 VGND.n49 VGND.n38 34.6358
R3711 VGND.n53 VGND.n38 34.6358
R3712 VGND.n54 VGND.n53 34.6358
R3713 VGND.n55 VGND.n54 34.6358
R3714 VGND.n55 VGND.n35 34.6358
R3715 VGND.n109 VGND.n108 34.6358
R3716 VGND.n82 VGND.n81 34.6358
R3717 VGND.n86 VGND.n85 34.6358
R3718 VGND.n150 VGND.n149 34.6358
R3719 VGND.n154 VGND.n153 34.6358
R3720 VGND.n1153 VGND.n1135 34.6358
R3721 VGND.n1149 VGND.n1135 34.6358
R3722 VGND.n1149 VGND.n1148 34.6358
R3723 VGND.n1148 VGND.n1147 34.6358
R3724 VGND.n1147 VGND.n1137 34.6358
R3725 VGND.n1131 VGND.n1105 34.6358
R3726 VGND.n1126 VGND.n1106 34.6358
R3727 VGND.n1122 VGND.n1106 34.6358
R3728 VGND.n1122 VGND.n1121 34.6358
R3729 VGND.n1121 VGND.n1120 34.6358
R3730 VGND.n1120 VGND.n1108 34.6358
R3731 VGND.n486 VGND.n481 34.6358
R3732 VGND.n491 VGND.n490 34.6358
R3733 VGND.n2267 VGND.n2262 34.6358
R3734 VGND.n2272 VGND.n2271 34.6358
R3735 VGND.n522 VGND.n517 34.6358
R3736 VGND.n527 VGND.n526 34.6358
R3737 VGND.n2196 VGND.n2195 34.6358
R3738 VGND.n2204 VGND.n2203 34.6358
R3739 VGND.n2200 VGND.n2199 34.6358
R3740 VGND.n2243 VGND.n542 34.6358
R3741 VGND.n2243 VGND.n2242 34.6358
R3742 VGND.n2242 VGND.n2241 34.6358
R3743 VGND.n2241 VGND.n2227 34.6358
R3744 VGND.n2237 VGND.n2227 34.6358
R3745 VGND.n1361 VGND.n1356 34.6358
R3746 VGND.n1381 VGND.n1357 34.6358
R3747 VGND.n1381 VGND.n1380 34.6358
R3748 VGND.n1380 VGND.n1379 34.6358
R3749 VGND.n1379 VGND.n1365 34.6358
R3750 VGND.n1375 VGND.n1365 34.6358
R3751 VGND.n2998 VGND.n2997 34.6358
R3752 VGND.n2 VGND.t1270 34.4422
R3753 VGND.n122 VGND.n121 33.1299
R3754 VGND.n2215 VGND.n544 33.1299
R3755 VGND.n111 VGND.n93 32.377
R3756 VGND.n187 VGND.n186 32.377
R3757 VGND.n111 VGND.n110 32.377
R3758 VGND.n88 VGND.n87 32.377
R3759 VGND.n156 VGND.n155 32.377
R3760 VGND.n2206 VGND.n2205 32.377
R3761 VGND.n2206 VGND.n2184 32.0005
R3762 VGND.n497 VGND.n494 30.4946
R3763 VGND.n2278 VGND.n2275 30.4946
R3764 VGND.n533 VGND.n530 30.4946
R3765 VGND.n190 VGND.n167 29.8709
R3766 VGND.n1143 VGND.n1142 28.9887
R3767 VGND.n1116 VGND.n1115 28.9887
R3768 VGND.n2235 VGND.n2234 28.9887
R3769 VGND.n1373 VGND.n1372 28.9887
R3770 VGND.n2985 VGND.n2984 27.8593
R3771 VGND.n22 VGND.n21 27.8593
R3772 VGND.n2955 VGND.n2954 27.8593
R3773 VGND.n48 VGND.n47 27.8593
R3774 VGND.n2256 VGND.n2255 27.0003
R3775 VGND.n161 VGND.n160 26.8591
R3776 VGND.n184 VGND.n173 26.3534
R3777 VGND.n108 VGND.n98 26.3534
R3778 VGND.n85 VGND.n74 26.3534
R3779 VGND.n153 VGND.n142 26.3534
R3780 VGND.n2203 VGND.n2188 26.3534
R3781 VGND.n129 VGND.n68 25.977
R3782 VGND.n498 VGND.n497 25.977
R3783 VGND.n2279 VGND.n2278 25.977
R3784 VGND.n534 VGND.n533 25.977
R3785 VGND.n509 VGND.n506 25.977
R3786 VGND.n2980 VGND.t2445 24.9236
R3787 VGND.n2980 VGND.t2399 24.9236
R3788 VGND.n2979 VGND.t2436 24.9236
R3789 VGND.n2979 VGND.t2380 24.9236
R3790 VGND.n2977 VGND.t2456 24.9236
R3791 VGND.n2977 VGND.t2429 24.9236
R3792 VGND.n2976 VGND.t2441 24.9236
R3793 VGND.n2976 VGND.t2413 24.9236
R3794 VGND.n17 VGND.t2428 24.9236
R3795 VGND.n17 VGND.t2460 24.9236
R3796 VGND.n16 VGND.t2384 24.9236
R3797 VGND.n16 VGND.t2423 24.9236
R3798 VGND.n15 VGND.t2434 24.9236
R3799 VGND.n15 VGND.t2404 24.9236
R3800 VGND.n14 VGND.t2394 24.9236
R3801 VGND.n14 VGND.t2450 24.9236
R3802 VGND.n176 VGND.t2374 24.9236
R3803 VGND.n176 VGND.t2415 24.9236
R3804 VGND.n175 VGND.t2432 24.9236
R3805 VGND.n175 VGND.t2372 24.9236
R3806 VGND.n172 VGND.t2382 24.9236
R3807 VGND.n172 VGND.t2001 24.9236
R3808 VGND.n171 VGND.t2438 24.9236
R3809 VGND.n171 VGND.t1416 24.9236
R3810 VGND.n170 VGND.t2000 24.9236
R3811 VGND.n170 VGND.t2002 24.9236
R3812 VGND.n169 VGND.t1424 24.9236
R3813 VGND.n169 VGND.t1419 24.9236
R3814 VGND.n2950 VGND.t2449 24.9236
R3815 VGND.n2950 VGND.t2368 24.9236
R3816 VGND.n2949 VGND.t2378 24.9236
R3817 VGND.n2949 VGND.t2386 24.9236
R3818 VGND.n43 VGND.t2402 24.9236
R3819 VGND.n43 VGND.t2437 24.9236
R3820 VGND.n42 VGND.t2388 24.9236
R3821 VGND.n42 VGND.t2427 24.9236
R3822 VGND.n41 VGND.t2409 24.9236
R3823 VGND.n41 VGND.t2370 24.9236
R3824 VGND.n40 VGND.t2396 24.9236
R3825 VGND.n40 VGND.t2453 24.9236
R3826 VGND.n96 VGND.t2421 24.9236
R3827 VGND.n96 VGND.t2458 24.9236
R3828 VGND.n97 VGND.t2425 24.9236
R3829 VGND.n97 VGND.t893 24.9236
R3830 VGND.n95 VGND.t889 24.9236
R3831 VGND.n95 VGND.t883 24.9236
R3832 VGND.n100 VGND.t2417 24.9236
R3833 VGND.n100 VGND.t2452 24.9236
R3834 VGND.n77 VGND.t2410 24.9236
R3835 VGND.n77 VGND.t2444 24.9236
R3836 VGND.n76 VGND.t2390 24.9236
R3837 VGND.n76 VGND.t2431 24.9236
R3838 VGND.n73 VGND.t2414 24.9236
R3839 VGND.n73 VGND.t756 24.9236
R3840 VGND.n72 VGND.t2401 24.9236
R3841 VGND.n72 VGND.t1168 24.9236
R3842 VGND.n71 VGND.t752 24.9236
R3843 VGND.n71 VGND.t746 24.9236
R3844 VGND.n70 VGND.t1167 24.9236
R3845 VGND.n70 VGND.t1165 24.9236
R3846 VGND.n145 VGND.t2408 24.9236
R3847 VGND.n145 VGND.t2439 24.9236
R3848 VGND.n144 VGND.t2454 24.9236
R3849 VGND.n144 VGND.t2406 24.9236
R3850 VGND.n141 VGND.t2411 24.9236
R3851 VGND.n141 VGND.t1769 24.9236
R3852 VGND.n140 VGND.t2366 24.9236
R3853 VGND.n140 VGND.t39 24.9236
R3854 VGND.n139 VGND.t1259 24.9236
R3855 VGND.n139 VGND.t1227 24.9236
R3856 VGND.n138 VGND.t1141 24.9236
R3857 VGND.n138 VGND.t302 24.9236
R3858 VGND.n1139 VGND.t63 24.9236
R3859 VGND.n1139 VGND.t77 24.9236
R3860 VGND.n1141 VGND.t2358 24.9236
R3861 VGND.n1141 VGND.t1290 24.9236
R3862 VGND.n1111 VGND.t497 24.9236
R3863 VGND.n1111 VGND.t498 24.9236
R3864 VGND.n1110 VGND.t65 24.9236
R3865 VGND.n1110 VGND.t1074 24.9236
R3866 VGND.n1114 VGND.t438 24.9236
R3867 VGND.n1114 VGND.t2362 24.9236
R3868 VGND.n1113 VGND.t2359 24.9236
R3869 VGND.n1113 VGND.t1291 24.9236
R3870 VGND.n488 VGND.t396 24.9236
R3871 VGND.n488 VGND.t71 24.9236
R3872 VGND.n487 VGND.t392 24.9236
R3873 VGND.n487 VGND.t465 24.9236
R3874 VGND.n478 VGND.t2147 24.9236
R3875 VGND.n478 VGND.t395 24.9236
R3876 VGND.n477 VGND.t1938 24.9236
R3877 VGND.n477 VGND.t2261 24.9236
R3878 VGND.n496 VGND.t235 24.9236
R3879 VGND.n496 VGND.t236 24.9236
R3880 VGND.n495 VGND.t1940 24.9236
R3881 VGND.n495 VGND.t1939 24.9236
R3882 VGND.n2269 VGND.t2361 24.9236
R3883 VGND.n2269 VGND.t2255 24.9236
R3884 VGND.n2268 VGND.t1077 24.9236
R3885 VGND.n2268 VGND.t1327 24.9236
R3886 VGND.n2259 VGND.t1575 24.9236
R3887 VGND.n2259 VGND.t1082 24.9236
R3888 VGND.n2258 VGND.t295 24.9236
R3889 VGND.n2258 VGND.t73 24.9236
R3890 VGND.n2277 VGND.t873 24.9236
R3891 VGND.n2277 VGND.t874 24.9236
R3892 VGND.n2276 VGND.t2604 24.9236
R3893 VGND.n2276 VGND.t2605 24.9236
R3894 VGND.n524 VGND.t394 24.9236
R3895 VGND.n524 VGND.t468 24.9236
R3896 VGND.n523 VGND.t2257 24.9236
R3897 VGND.n523 VGND.t441 24.9236
R3898 VGND.n514 VGND.t414 24.9236
R3899 VGND.n514 VGND.t393 24.9236
R3900 VGND.n513 VGND.t898 24.9236
R3901 VGND.n513 VGND.t1342 24.9236
R3902 VGND.n532 VGND.t416 24.9236
R3903 VGND.n532 VGND.t415 24.9236
R3904 VGND.n531 VGND.t900 24.9236
R3905 VGND.n531 VGND.t899 24.9236
R3906 VGND.n2186 VGND.t75 24.9236
R3907 VGND.n2186 VGND.t1324 24.9236
R3908 VGND.n2187 VGND.t1391 24.9236
R3909 VGND.n2187 VGND.t1079 24.9236
R3910 VGND.n2185 VGND.t1395 24.9236
R3911 VGND.n2185 VGND.t1393 24.9236
R3912 VGND.n2190 VGND.t1081 24.9236
R3913 VGND.n2190 VGND.t1288 24.9236
R3914 VGND.n2230 VGND.t67 24.9236
R3915 VGND.n2230 VGND.t1075 24.9236
R3916 VGND.n2229 VGND.t442 24.9236
R3917 VGND.n2229 VGND.t466 24.9236
R3918 VGND.n2233 VGND.t2360 24.9236
R3919 VGND.n2233 VGND.t1292 24.9236
R3920 VGND.n2231 VGND.t79 24.9236
R3921 VGND.n2231 VGND.t1325 24.9236
R3922 VGND.n1368 VGND.t2363 24.9236
R3923 VGND.n1368 VGND.t1284 24.9236
R3924 VGND.n1367 VGND.t1326 24.9236
R3925 VGND.n1367 VGND.t1328 24.9236
R3926 VGND.n1371 VGND.t1285 24.9236
R3927 VGND.n1371 VGND.t496 24.9236
R3928 VGND.n1369 VGND.t2256 24.9236
R3929 VGND.n1369 VGND.t439 24.9236
R3930 VGND.n187 VGND.n166 24.4711
R3931 VGND.n61 VGND.n36 24.4711
R3932 VGND.n123 VGND.n122 24.4711
R3933 VGND.n88 VGND.n67 24.4711
R3934 VGND.n129 VGND.n128 24.4711
R3935 VGND.n156 VGND.n135 24.4711
R3936 VGND.n498 VGND.n474 24.4711
R3937 VGND.n2279 VGND.n2253 24.4711
R3938 VGND.n534 VGND.n505 24.4711
R3939 VGND.n509 VGND.n508 24.4711
R3940 VGND.n2216 VGND.n2215 24.4711
R3941 VGND.n2223 VGND.n541 24.4711
R3942 VGND.n164 VGND.n136 23.7181
R3943 VGND.n2993 VGND.n2972 23.7181
R3944 VGND.n3010 VGND.n9 23.7181
R3945 VGND.n3010 VGND.n10 23.7181
R3946 VGND.n2966 VGND.n2945 23.7181
R3947 VGND.n65 VGND.n35 23.7181
R3948 VGND.n1155 VGND.n1153 23.7181
R3949 VGND.n1127 VGND.n1105 23.7181
R3950 VGND.n1127 VGND.n1126 23.7181
R3951 VGND.n2283 VGND.n2252 23.7181
R3952 VGND.n2210 VGND.n545 23.7181
R3953 VGND.n2247 VGND.n542 23.7181
R3954 VGND.n1385 VGND.n1356 23.7181
R3955 VGND.n1385 VGND.n1357 23.7181
R3956 VGND.n2997 VGND.n2972 23.7181
R3957 VGND.n117 VGND.n115 23.3417
R3958 VGND.n117 VGND.n92 23.3417
R3959 VGND.n2211 VGND.n2210 23.3417
R3960 VGND.n1143 VGND.n1140 21.4593
R3961 VGND.n1116 VGND.n1112 21.4593
R3962 VGND.n2236 VGND.n2235 21.4593
R3963 VGND.n1374 VGND.n1373 21.4593
R3964 VGND.n179 VGND.n178 21.0905
R3965 VGND.n102 VGND.n101 21.0905
R3966 VGND.n80 VGND.n79 21.0905
R3967 VGND.n148 VGND.n147 21.0905
R3968 VGND.n180 VGND.n179 20.3299
R3969 VGND.n103 VGND.n102 20.3299
R3970 VGND.n81 VGND.n80 20.3299
R3971 VGND.n149 VGND.n148 20.3299
R3972 VGND.n494 VGND.n479 19.9534
R3973 VGND.n2275 VGND.n2260 19.9534
R3974 VGND.n530 VGND.n515 19.9534
R3975 VGND.n3006 VGND.n3005 19.2005
R3976 VGND.n61 VGND.n60 19.2005
R3977 VGND.n2223 VGND.n2222 19.2005
R3978 VGND.n1361 VGND.n1360 19.2005
R3979 VGND.t1135 VGND.t2606 16.8587
R3980 VGND.t1454 VGND.t2608 16.8587
R3981 VGND.t2159 VGND.t821 16.8587
R3982 VGND.t1098 VGND.t819 16.8587
R3983 VGND.n1133 VGND.n1132 16.077
R3984 VGND.n3000 VGND.n2999 16.077
R3985 VGND.n60 VGND.n59 15.4358
R3986 VGND.n2222 VGND.n2221 15.4358
R3987 VGND.n3005 VGND.n3004 14.6829
R3988 VGND.n160 VGND.n159 14.6829
R3989 VGND.n2255 VGND.n2254 14.6829
R3990 VGND.n1360 VGND.n1359 14.6829
R3991 VGND.n483 VGND.n482 14.5711
R3992 VGND.n2264 VGND.n2263 14.5711
R3993 VGND.n519 VGND.n518 14.5711
R3994 VGND.n2194 VGND.n2193 14.5711
R3995 VGND.n133 VGND.n68 14.3064
R3996 VGND.n538 VGND.n506 14.3064
R3997 VGND.n490 VGND.n489 13.9299
R3998 VGND.n2271 VGND.n2270 13.9299
R3999 VGND.n526 VGND.n525 13.9299
R4000 VGND.n2199 VGND.n2191 13.9299
R4001 VGND.n65 VGND.n36 13.5534
R4002 VGND.n2247 VGND.n541 13.5534
R4003 VGND.n193 VGND.n166 13.177
R4004 VGND.n133 VGND.n67 13.177
R4005 VGND.n164 VGND.n135 13.177
R4006 VGND.n502 VGND.n474 13.177
R4007 VGND.n2283 VGND.n2253 13.177
R4008 VGND.n538 VGND.n505 13.177
R4009 VGND.n193 VGND.n167 12.8005
R4010 VGND.n502 VGND.n475 12.8005
R4011 VGND.n3023 VGND.t2691 12.5645
R4012 VGND.n1132 VGND.n1131 10.5417
R4013 VGND.n2999 VGND.n2998 10.5417
R4014 VGND.n3004 VGND.n3003 10.0534
R4015 VGND.n1359 VGND.n1358 10.0534
R4016 VGND.n20 VGND.n19 9.3005
R4017 VGND.n21 VGND.n13 9.3005
R4018 VGND.n24 VGND.n23 9.3005
R4019 VGND.n25 VGND.n12 9.3005
R4020 VGND.n27 VGND.n26 9.3005
R4021 VGND.n28 VGND.n11 9.3005
R4022 VGND.n30 VGND.n29 9.3005
R4023 VGND.n31 VGND.n9 9.3005
R4024 VGND.n3008 VGND.n10 9.3005
R4025 VGND.n3007 VGND.n3006 9.3005
R4026 VGND.n3010 VGND.n3009 9.3005
R4027 VGND.n191 VGND.n167 9.3005
R4028 VGND.n180 VGND.n174 9.3005
R4029 VGND.n182 VGND.n181 9.3005
R4030 VGND.n184 VGND.n183 9.3005
R4031 VGND.n185 VGND.n168 9.3005
R4032 VGND.n188 VGND.n187 9.3005
R4033 VGND.n189 VGND.n166 9.3005
R4034 VGND.n193 VGND.n192 9.3005
R4035 VGND.n2953 VGND.n2952 9.3005
R4036 VGND.n2954 VGND.n2948 9.3005
R4037 VGND.n2957 VGND.n2956 9.3005
R4038 VGND.n2958 VGND.n2947 9.3005
R4039 VGND.n2960 VGND.n2959 9.3005
R4040 VGND.n2961 VGND.n2946 9.3005
R4041 VGND.n2963 VGND.n2962 9.3005
R4042 VGND.n2964 VGND.n2945 9.3005
R4043 VGND.n2966 VGND.n2965 9.3005
R4044 VGND.n59 VGND.n58 9.3005
R4045 VGND.n46 VGND.n45 9.3005
R4046 VGND.n47 VGND.n39 9.3005
R4047 VGND.n50 VGND.n49 9.3005
R4048 VGND.n51 VGND.n38 9.3005
R4049 VGND.n53 VGND.n52 9.3005
R4050 VGND.n54 VGND.n37 9.3005
R4051 VGND.n56 VGND.n55 9.3005
R4052 VGND.n57 VGND.n35 9.3005
R4053 VGND.n63 VGND.n36 9.3005
R4054 VGND.n62 VGND.n61 9.3005
R4055 VGND.n65 VGND.n64 9.3005
R4056 VGND.n124 VGND.n123 9.3005
R4057 VGND.n103 VGND.n99 9.3005
R4058 VGND.n106 VGND.n105 9.3005
R4059 VGND.n108 VGND.n107 9.3005
R4060 VGND.n109 VGND.n94 9.3005
R4061 VGND.n112 VGND.n111 9.3005
R4062 VGND.n114 VGND.n113 9.3005
R4063 VGND.n120 VGND.n119 9.3005
R4064 VGND.n122 VGND.n91 9.3005
R4065 VGND.n118 VGND.n117 9.3005
R4066 VGND.n128 VGND.n127 9.3005
R4067 VGND.n81 VGND.n75 9.3005
R4068 VGND.n83 VGND.n82 9.3005
R4069 VGND.n85 VGND.n84 9.3005
R4070 VGND.n86 VGND.n69 9.3005
R4071 VGND.n89 VGND.n88 9.3005
R4072 VGND.n90 VGND.n67 9.3005
R4073 VGND.n131 VGND.n68 9.3005
R4074 VGND.n130 VGND.n129 9.3005
R4075 VGND.n133 VGND.n132 9.3005
R4076 VGND.n162 VGND.n136 9.3005
R4077 VGND.n149 VGND.n143 9.3005
R4078 VGND.n151 VGND.n150 9.3005
R4079 VGND.n153 VGND.n152 9.3005
R4080 VGND.n154 VGND.n137 9.3005
R4081 VGND.n157 VGND.n156 9.3005
R4082 VGND.n158 VGND.n135 9.3005
R4083 VGND.n164 VGND.n163 9.3005
R4084 VGND.n1144 VGND.n1143 9.3005
R4085 VGND.n1145 VGND.n1137 9.3005
R4086 VGND.n1147 VGND.n1146 9.3005
R4087 VGND.n1148 VGND.n1136 9.3005
R4088 VGND.n1150 VGND.n1149 9.3005
R4089 VGND.n1151 VGND.n1135 9.3005
R4090 VGND.n1153 VGND.n1152 9.3005
R4091 VGND.n1156 VGND.n1155 9.3005
R4092 VGND.n1117 VGND.n1116 9.3005
R4093 VGND.n1118 VGND.n1108 9.3005
R4094 VGND.n1120 VGND.n1119 9.3005
R4095 VGND.n1121 VGND.n1107 9.3005
R4096 VGND.n1123 VGND.n1122 9.3005
R4097 VGND.n1124 VGND.n1106 9.3005
R4098 VGND.n1126 VGND.n1125 9.3005
R4099 VGND.n1129 VGND.n1105 9.3005
R4100 VGND.n1131 VGND.n1130 9.3005
R4101 VGND.n1128 VGND.n1127 9.3005
R4102 VGND.n500 VGND.n474 9.3005
R4103 VGND.n484 VGND.n481 9.3005
R4104 VGND.n486 VGND.n485 9.3005
R4105 VGND.n490 VGND.n480 9.3005
R4106 VGND.n492 VGND.n491 9.3005
R4107 VGND.n494 VGND.n493 9.3005
R4108 VGND.n497 VGND.n476 9.3005
R4109 VGND.n499 VGND.n498 9.3005
R4110 VGND.n502 VGND.n501 9.3005
R4111 VGND.n2281 VGND.n2253 9.3005
R4112 VGND.n2265 VGND.n2262 9.3005
R4113 VGND.n2267 VGND.n2266 9.3005
R4114 VGND.n2271 VGND.n2261 9.3005
R4115 VGND.n2273 VGND.n2272 9.3005
R4116 VGND.n2275 VGND.n2274 9.3005
R4117 VGND.n2278 VGND.n2257 9.3005
R4118 VGND.n2280 VGND.n2279 9.3005
R4119 VGND.n2256 VGND.n2252 9.3005
R4120 VGND.n2283 VGND.n2282 9.3005
R4121 VGND.n508 VGND.n507 9.3005
R4122 VGND.n511 VGND.n506 9.3005
R4123 VGND.n536 VGND.n505 9.3005
R4124 VGND.n520 VGND.n517 9.3005
R4125 VGND.n522 VGND.n521 9.3005
R4126 VGND.n526 VGND.n516 9.3005
R4127 VGND.n528 VGND.n527 9.3005
R4128 VGND.n530 VGND.n529 9.3005
R4129 VGND.n533 VGND.n512 9.3005
R4130 VGND.n535 VGND.n534 9.3005
R4131 VGND.n510 VGND.n509 9.3005
R4132 VGND.n538 VGND.n537 9.3005
R4133 VGND.n2217 VGND.n2216 9.3005
R4134 VGND.n2208 VGND.n545 9.3005
R4135 VGND.n2195 VGND.n2192 9.3005
R4136 VGND.n2197 VGND.n2196 9.3005
R4137 VGND.n2199 VGND.n2198 9.3005
R4138 VGND.n2201 VGND.n2200 9.3005
R4139 VGND.n2203 VGND.n2202 9.3005
R4140 VGND.n2204 VGND.n2183 9.3005
R4141 VGND.n2207 VGND.n2206 9.3005
R4142 VGND.n2213 VGND.n2212 9.3005
R4143 VGND.n2215 VGND.n2214 9.3005
R4144 VGND.n2210 VGND.n2209 9.3005
R4145 VGND.n2235 VGND.n2228 9.3005
R4146 VGND.n2238 VGND.n2237 9.3005
R4147 VGND.n2239 VGND.n2227 9.3005
R4148 VGND.n2241 VGND.n2240 9.3005
R4149 VGND.n2242 VGND.n2226 9.3005
R4150 VGND.n2244 VGND.n2243 9.3005
R4151 VGND.n2245 VGND.n542 9.3005
R4152 VGND.n2225 VGND.n541 9.3005
R4153 VGND.n2224 VGND.n2223 9.3005
R4154 VGND.n2221 VGND.n2220 9.3005
R4155 VGND.n2247 VGND.n2246 9.3005
R4156 VGND.n1373 VGND.n1366 9.3005
R4157 VGND.n1376 VGND.n1375 9.3005
R4158 VGND.n1377 VGND.n1365 9.3005
R4159 VGND.n1379 VGND.n1378 9.3005
R4160 VGND.n1380 VGND.n1364 9.3005
R4161 VGND.n1382 VGND.n1381 9.3005
R4162 VGND.n1383 VGND.n1357 9.3005
R4163 VGND.n1363 VGND.n1356 9.3005
R4164 VGND.n1362 VGND.n1361 9.3005
R4165 VGND.n1385 VGND.n1384 9.3005
R4166 VGND.n2982 VGND.n2978 9.3005
R4167 VGND.n2984 VGND.n2983 9.3005
R4168 VGND.n2986 VGND.n2975 9.3005
R4169 VGND.n2988 VGND.n2987 9.3005
R4170 VGND.n2989 VGND.n2974 9.3005
R4171 VGND.n2991 VGND.n2990 9.3005
R4172 VGND.n2992 VGND.n2973 9.3005
R4173 VGND.n2994 VGND.n2993 9.3005
R4174 VGND.n2995 VGND.n2972 9.3005
R4175 VGND.n2997 VGND.n2996 9.3005
R4176 VGND.n2998 VGND.n34 9.3005
R4177 VGND.n181 VGND.n173 8.28285
R4178 VGND.n82 VGND.n74 8.28285
R4179 VGND.n150 VGND.n142 8.28285
R4180 VGND.n2636 VGND.n2635 7.9105
R4181 VGND.n2693 VGND.n337 7.9105
R4182 VGND.n2692 VGND.n338 7.9105
R4183 VGND.n2687 VGND.n343 7.9105
R4184 VGND.n2686 VGND.n344 7.9105
R4185 VGND.n2681 VGND.n349 7.9105
R4186 VGND.n2680 VGND.n350 7.9105
R4187 VGND.n2675 VGND.n2674 7.9105
R4188 VGND.n2712 VGND.n2711 7.9105
R4189 VGND.n2721 VGND.n2720 7.9105
R4190 VGND.n2745 VGND.n2744 7.9105
R4191 VGND.n2759 VGND.n2758 7.9105
R4192 VGND.n2783 VGND.n288 7.9105
R4193 VGND.n2785 VGND.n2784 7.9105
R4194 VGND.n2794 VGND.n2793 7.9105
R4195 VGND.n2937 VGND.n2936 7.9105
R4196 VGND.n2559 VGND.n401 7.9105
R4197 VGND.n2558 VGND.n402 7.9105
R4198 VGND.n2557 VGND.n403 7.9105
R4199 VGND.n2556 VGND.n404 7.9105
R4200 VGND.n2555 VGND.n405 7.9105
R4201 VGND.n2554 VGND.n406 7.9105
R4202 VGND.n2553 VGND.n407 7.9105
R4203 VGND.n2552 VGND.n408 7.9105
R4204 VGND.n2551 VGND.n409 7.9105
R4205 VGND.n2550 VGND.n410 7.9105
R4206 VGND.n2549 VGND.n411 7.9105
R4207 VGND.n2548 VGND.n412 7.9105
R4208 VGND.n2547 VGND.n2546 7.9105
R4209 VGND.n2798 VGND.n282 7.9105
R4210 VGND.n2797 VGND.n283 7.9105
R4211 VGND.n2534 VGND.n2533 7.9105
R4212 VGND.n2357 VGND.n2356 7.9105
R4213 VGND.n2374 VGND.n2373 7.9105
R4214 VGND.n2383 VGND.n2382 7.9105
R4215 VGND.n2400 VGND.n2399 7.9105
R4216 VGND.n2409 VGND.n2408 7.9105
R4217 VGND.n2426 VGND.n2425 7.9105
R4218 VGND.n2435 VGND.n2434 7.9105
R4219 VGND.n2452 VGND.n2451 7.9105
R4220 VGND.n2461 VGND.n2460 7.9105
R4221 VGND.n2478 VGND.n2477 7.9105
R4222 VGND.n2487 VGND.n2486 7.9105
R4223 VGND.n2509 VGND.n2508 7.9105
R4224 VGND.n2802 VGND.n279 7.9105
R4225 VGND.n2801 VGND.n280 7.9105
R4226 VGND.n420 VGND.n419 7.9105
R4227 VGND.n2530 VGND.n2529 7.9105
R4228 VGND.n2361 VGND.n2360 7.9105
R4229 VGND.n2370 VGND.n2369 7.9105
R4230 VGND.n2387 VGND.n2386 7.9105
R4231 VGND.n2396 VGND.n2395 7.9105
R4232 VGND.n2413 VGND.n2412 7.9105
R4233 VGND.n2422 VGND.n2421 7.9105
R4234 VGND.n2439 VGND.n2438 7.9105
R4235 VGND.n2448 VGND.n2447 7.9105
R4236 VGND.n2465 VGND.n2464 7.9105
R4237 VGND.n2474 VGND.n2473 7.9105
R4238 VGND.n2491 VGND.n2490 7.9105
R4239 VGND.n2505 VGND.n2504 7.9105
R4240 VGND.n2805 VGND.n277 7.9105
R4241 VGND.n2807 VGND.n2806 7.9105
R4242 VGND.n2819 VGND.n273 7.9105
R4243 VGND.n2818 VGND.n2817 7.9105
R4244 VGND.n1908 VGND.n1907 7.9105
R4245 VGND.n1917 VGND.n1916 7.9105
R4246 VGND.n1919 VGND.n1918 7.9105
R4247 VGND.n1928 VGND.n1927 7.9105
R4248 VGND.n1930 VGND.n1929 7.9105
R4249 VGND.n1939 VGND.n1938 7.9105
R4250 VGND.n1941 VGND.n1940 7.9105
R4251 VGND.n1950 VGND.n1949 7.9105
R4252 VGND.n1952 VGND.n1951 7.9105
R4253 VGND.n1961 VGND.n1960 7.9105
R4254 VGND.n1963 VGND.n1962 7.9105
R4255 VGND.n1972 VGND.n1971 7.9105
R4256 VGND.n1974 VGND.n1973 7.9105
R4257 VGND.n2823 VGND.n270 7.9105
R4258 VGND.n2822 VGND.n271 7.9105
R4259 VGND.n1990 VGND.n1989 7.9105
R4260 VGND.n2063 VGND.n591 7.9105
R4261 VGND.n2062 VGND.n2061 7.9105
R4262 VGND.n2167 VGND.n556 7.9105
R4263 VGND.n2166 VGND.n557 7.9105
R4264 VGND.n2159 VGND.n562 7.9105
R4265 VGND.n2158 VGND.n563 7.9105
R4266 VGND.n2151 VGND.n568 7.9105
R4267 VGND.n2150 VGND.n569 7.9105
R4268 VGND.n2143 VGND.n574 7.9105
R4269 VGND.n2142 VGND.n575 7.9105
R4270 VGND.n2135 VGND.n580 7.9105
R4271 VGND.n2134 VGND.n581 7.9105
R4272 VGND.n2827 VGND.n267 7.9105
R4273 VGND.n2826 VGND.n268 7.9105
R4274 VGND.n1999 VGND.n1998 7.9105
R4275 VGND.n1997 VGND.n1996 7.9105
R4276 VGND.n2067 VGND.n2066 7.9105
R4277 VGND.n2171 VGND.n553 7.9105
R4278 VGND.n2170 VGND.n554 7.9105
R4279 VGND.n2163 VGND.n559 7.9105
R4280 VGND.n2162 VGND.n560 7.9105
R4281 VGND.n2155 VGND.n565 7.9105
R4282 VGND.n2154 VGND.n566 7.9105
R4283 VGND.n2147 VGND.n571 7.9105
R4284 VGND.n2146 VGND.n572 7.9105
R4285 VGND.n2139 VGND.n577 7.9105
R4286 VGND.n2138 VGND.n578 7.9105
R4287 VGND.n2131 VGND.n2130 7.9105
R4288 VGND.n2830 VGND.n265 7.9105
R4289 VGND.n2832 VGND.n2831 7.9105
R4290 VGND.n2844 VGND.n261 7.9105
R4291 VGND.n2843 VGND.n2842 7.9105
R4292 VGND.n1901 VGND.n548 7.9105
R4293 VGND.n2175 VGND.n2174 7.9105
R4294 VGND.n1759 VGND.n1758 7.9105
R4295 VGND.n1768 VGND.n1767 7.9105
R4296 VGND.n1770 VGND.n1769 7.9105
R4297 VGND.n1779 VGND.n1778 7.9105
R4298 VGND.n1781 VGND.n1780 7.9105
R4299 VGND.n1790 VGND.n1789 7.9105
R4300 VGND.n1792 VGND.n1791 7.9105
R4301 VGND.n1801 VGND.n1800 7.9105
R4302 VGND.n1803 VGND.n1802 7.9105
R4303 VGND.n1812 VGND.n1811 7.9105
R4304 VGND.n1814 VGND.n1813 7.9105
R4305 VGND.n2848 VGND.n258 7.9105
R4306 VGND.n2847 VGND.n259 7.9105
R4307 VGND.n1830 VGND.n1829 7.9105
R4308 VGND.n1899 VGND.n629 7.9105
R4309 VGND.n1685 VGND.n1684 7.9105
R4310 VGND.n1687 VGND.n1686 7.9105
R4311 VGND.n1884 VGND.n643 7.9105
R4312 VGND.n1883 VGND.n644 7.9105
R4313 VGND.n1876 VGND.n649 7.9105
R4314 VGND.n1875 VGND.n650 7.9105
R4315 VGND.n1868 VGND.n655 7.9105
R4316 VGND.n1867 VGND.n656 7.9105
R4317 VGND.n1860 VGND.n661 7.9105
R4318 VGND.n1859 VGND.n662 7.9105
R4319 VGND.n1852 VGND.n1851 7.9105
R4320 VGND.n2852 VGND.n255 7.9105
R4321 VGND.n2851 VGND.n256 7.9105
R4322 VGND.n1839 VGND.n1838 7.9105
R4323 VGND.n1837 VGND.n1836 7.9105
R4324 VGND.n1896 VGND.n633 7.9105
R4325 VGND.n1895 VGND.n634 7.9105
R4326 VGND.n1888 VGND.n640 7.9105
R4327 VGND.n1887 VGND.n641 7.9105
R4328 VGND.n1880 VGND.n646 7.9105
R4329 VGND.n1879 VGND.n647 7.9105
R4330 VGND.n1872 VGND.n652 7.9105
R4331 VGND.n1871 VGND.n653 7.9105
R4332 VGND.n1864 VGND.n658 7.9105
R4333 VGND.n1863 VGND.n659 7.9105
R4334 VGND.n1856 VGND.n664 7.9105
R4335 VGND.n1855 VGND.n730 7.9105
R4336 VGND.n2855 VGND.n253 7.9105
R4337 VGND.n2857 VGND.n2856 7.9105
R4338 VGND.n2869 VGND.n249 7.9105
R4339 VGND.n2868 VGND.n2867 7.9105
R4340 VGND.n1350 VGND.n1349 7.9105
R4341 VGND.n1892 VGND.n636 7.9105
R4342 VGND.n1891 VGND.n637 7.9105
R4343 VGND.n868 VGND.n867 7.9105
R4344 VGND.n866 VGND.n812 7.9105
R4345 VGND.n865 VGND.n813 7.9105
R4346 VGND.n864 VGND.n814 7.9105
R4347 VGND.n863 VGND.n815 7.9105
R4348 VGND.n862 VGND.n816 7.9105
R4349 VGND.n861 VGND.n817 7.9105
R4350 VGND.n860 VGND.n859 7.9105
R4351 VGND.n1669 VGND.n732 7.9105
R4352 VGND.n1668 VGND.n1667 7.9105
R4353 VGND.n2873 VGND.n246 7.9105
R4354 VGND.n2872 VGND.n247 7.9105
R4355 VGND.n1655 VGND.n1654 7.9105
R4356 VGND.n1404 VGND.n801 7.9105
R4357 VGND.n1403 VGND.n802 7.9105
R4358 VGND.n1402 VGND.n1401 7.9105
R4359 VGND.n1488 VGND.n1487 7.9105
R4360 VGND.n1497 VGND.n1496 7.9105
R4361 VGND.n1514 VGND.n1513 7.9105
R4362 VGND.n1523 VGND.n1522 7.9105
R4363 VGND.n1540 VGND.n1539 7.9105
R4364 VGND.n1560 VGND.n758 7.9105
R4365 VGND.n1559 VGND.n1558 7.9105
R4366 VGND.n1628 VGND.n742 7.9105
R4367 VGND.n1630 VGND.n1629 7.9105
R4368 VGND.n2877 VGND.n243 7.9105
R4369 VGND.n2876 VGND.n244 7.9105
R4370 VGND.n741 VGND.n740 7.9105
R4371 VGND.n1651 VGND.n1650 7.9105
R4372 VGND.n1408 VGND.n1407 7.9105
R4373 VGND.n1417 VGND.n1416 7.9105
R4374 VGND.n1475 VGND.n1474 7.9105
R4375 VGND.n1484 VGND.n1483 7.9105
R4376 VGND.n1501 VGND.n1500 7.9105
R4377 VGND.n1510 VGND.n1509 7.9105
R4378 VGND.n1527 VGND.n1526 7.9105
R4379 VGND.n1536 VGND.n1535 7.9105
R4380 VGND.n1564 VGND.n1563 7.9105
R4381 VGND.n1588 VGND.n1587 7.9105
R4382 VGND.n1625 VGND.n744 7.9105
R4383 VGND.n1624 VGND.n745 7.9105
R4384 VGND.n2880 VGND.n240 7.9105
R4385 VGND.n2882 VGND.n2881 7.9105
R4386 VGND.n2894 VGND.n236 7.9105
R4387 VGND.n2893 VGND.n2892 7.9105
R4388 VGND.n1344 VGND.n1343 7.9105
R4389 VGND.n1421 VGND.n1420 7.9105
R4390 VGND.n1471 VGND.n783 7.9105
R4391 VGND.n1470 VGND.n784 7.9105
R4392 VGND.n1469 VGND.n785 7.9105
R4393 VGND.n1468 VGND.n786 7.9105
R4394 VGND.n1467 VGND.n787 7.9105
R4395 VGND.n1466 VGND.n788 7.9105
R4396 VGND.n1465 VGND.n1464 7.9105
R4397 VGND.n1591 VGND.n751 7.9105
R4398 VGND.n1593 VGND.n1592 7.9105
R4399 VGND.n1621 VGND.n747 7.9105
R4400 VGND.n1620 VGND.n1619 7.9105
R4401 VGND.n2898 VGND.n231 7.9105
R4402 VGND.n2897 VGND.n232 7.9105
R4403 VGND.n1607 VGND.n1606 7.9105
R4404 VGND.n1103 VGND.n1025 7.9105
R4405 VGND.n1102 VGND.n1026 7.9105
R4406 VGND.n1101 VGND.n1100 7.9105
R4407 VGND.n1321 VGND.n899 7.9105
R4408 VGND.n1320 VGND.n900 7.9105
R4409 VGND.n1313 VGND.n905 7.9105
R4410 VGND.n1312 VGND.n906 7.9105
R4411 VGND.n1305 VGND.n911 7.9105
R4412 VGND.n1304 VGND.n912 7.9105
R4413 VGND.n1068 VGND.n1067 7.9105
R4414 VGND.n1066 VGND.n1045 7.9105
R4415 VGND.n1065 VGND.n1046 7.9105
R4416 VGND.n1064 VGND.n1063 7.9105
R4417 VGND.n2902 VGND.n2901 7.9105
R4418 VGND.n233 VGND.n228 7.9105
R4419 VGND.n2913 VGND.n2912 7.9105
R4420 VGND.n1161 VGND.n888 7.9105
R4421 VGND.n1331 VGND.n1330 7.9105
R4422 VGND.n1325 VGND.n896 7.9105
R4423 VGND.n1324 VGND.n897 7.9105
R4424 VGND.n1317 VGND.n902 7.9105
R4425 VGND.n1316 VGND.n903 7.9105
R4426 VGND.n1309 VGND.n908 7.9105
R4427 VGND.n1308 VGND.n909 7.9105
R4428 VGND.n1301 VGND.n914 7.9105
R4429 VGND.n1300 VGND.n915 7.9105
R4430 VGND.n1295 VGND.n919 7.9105
R4431 VGND.n1294 VGND.n920 7.9105
R4432 VGND.n1289 VGND.n924 7.9105
R4433 VGND.n1288 VGND.n925 7.9105
R4434 VGND.n1287 VGND.n992 7.9105
R4435 VGND.n2917 VGND.n2916 7.9105
R4436 VGND.n489 VGND.n486 7.90638
R4437 VGND.n482 VGND.n481 7.90638
R4438 VGND.n2270 VGND.n2267 7.90638
R4439 VGND.n2263 VGND.n2262 7.90638
R4440 VGND.n525 VGND.n522 7.90638
R4441 VGND.n518 VGND.n517 7.90638
R4442 VGND.n2196 VGND.n2191 7.90638
R4443 VGND.n2195 VGND.n2194 7.90638
R4444 VGND.n1142 VGND.n1138 7.4049
R4445 VGND.n1115 VGND.n1109 7.4049
R4446 VGND.n2234 VGND.n2232 7.4049
R4447 VGND.n1372 VGND.n1370 7.4049
R4448 VGND VGND.n475 7.12482
R4449 VGND.n178 VGND.n177 6.85473
R4450 VGND.n79 VGND.n78 6.85473
R4451 VGND.n147 VGND.n146 6.85473
R4452 VGND.n2986 VGND.n2985 6.77697
R4453 VGND.n23 VGND.n22 6.77697
R4454 VGND.n2956 VGND.n2955 6.77697
R4455 VGND.n49 VGND.n48 6.77697
R4456 VGND.n3022 VGND.n3021 6.4005
R4457 VGND.n104 VGND.n98 5.27109
R4458 VGND.n2189 VGND.n2188 5.27109
R4459 VGND.n2565 VGND.n2564 4.5005
R4460 VGND.n2568 VGND.n2567 4.5005
R4461 VGND.n2571 VGND.n2570 4.5005
R4462 VGND.n2574 VGND.n2573 4.5005
R4463 VGND.n2577 VGND.n2576 4.5005
R4464 VGND.n2580 VGND.n2579 4.5005
R4465 VGND.n2583 VGND.n2582 4.5005
R4466 VGND.n2586 VGND.n2585 4.5005
R4467 VGND.n2589 VGND.n2588 4.5005
R4468 VGND.n2592 VGND.n2591 4.5005
R4469 VGND.n2595 VGND.n2594 4.5005
R4470 VGND.n2598 VGND.n2597 4.5005
R4471 VGND.n2601 VGND.n2600 4.5005
R4472 VGND.n2604 VGND.n2603 4.5005
R4473 VGND.n2607 VGND.n2606 4.5005
R4474 VGND.n335 VGND.n334 4.5005
R4475 VGND.n2627 VGND.n2626 4.5005
R4476 VGND.n2624 VGND.n2623 4.5005
R4477 VGND.n2621 VGND.n2620 4.5005
R4478 VGND.n2618 VGND.n2617 4.5005
R4479 VGND.n2615 VGND.n2614 4.5005
R4480 VGND.n2612 VGND.n2611 4.5005
R4481 VGND.n323 VGND.n322 4.5005
R4482 VGND.n316 VGND.n315 4.5005
R4483 VGND.n307 VGND.n306 4.5005
R4484 VGND.n2763 VGND.n299 4.5005
R4485 VGND.n2766 VGND.n2765 4.5005
R4486 VGND.n291 VGND.n290 4.5005
R4487 VGND.n2770 VGND.n297 4.5005
R4488 VGND.n205 VGND.n204 4.5005
R4489 VGND.n2631 VGND.n2630 4.5005
R4490 VGND.n2632 VGND.n331 4.5005
R4491 VGND.n2697 VGND.n2696 4.5005
R4492 VGND.n358 VGND.n340 4.5005
R4493 VGND.n365 VGND.n341 4.5005
R4494 VGND.n354 VGND.n346 4.5005
R4495 VGND.n376 VGND.n347 4.5005
R4496 VGND.n353 VGND.n352 4.5005
R4497 VGND.n390 VGND.n389 4.5005
R4498 VGND.n2708 VGND.n2707 4.5005
R4499 VGND.n2725 VGND.n2724 4.5005
R4500 VGND.n2741 VGND.n2740 4.5005
R4501 VGND.n2762 VGND.n300 4.5005
R4502 VGND.n2733 VGND.n289 4.5005
R4503 VGND.n2779 VGND.n2778 4.5005
R4504 VGND.n2772 VGND.n2771 4.5005
R4505 VGND.n2942 VGND.n2941 4.5005
R4506 VGND.n1019 VGND.n1018 4.5005
R4507 VGND.n1016 VGND.n1015 4.5005
R4508 VGND.n1181 VGND.n1180 4.5005
R4509 VGND.n1193 VGND.n1006 4.5005
R4510 VGND.n1200 VGND.n1004 4.5005
R4511 VGND.n1197 VGND.n1195 4.5005
R4512 VGND.n1213 VGND.n1212 4.5005
R4513 VGND.n1251 VGND.n1000 4.5005
R4514 VGND.n1254 VGND.n1253 4.5005
R4515 VGND.n1257 VGND.n1256 4.5005
R4516 VGND.n1260 VGND.n1259 4.5005
R4517 VGND.n1263 VGND.n1262 4.5005
R4518 VGND.n1269 VGND.n998 4.5005
R4519 VGND.n1266 VGND.n1265 4.5005
R4520 VGND.n995 VGND.n994 4.5005
R4521 VGND.n1022 VGND.n1021 4.5005
R4522 VGND.n1165 VGND.n1164 4.5005
R4523 VGND.n1170 VGND.n891 4.5005
R4524 VGND.n1011 VGND.n892 4.5005
R4525 VGND.n1183 VGND.n1182 4.5005
R4526 VGND.n1192 VGND.n1191 4.5005
R4527 VGND.n1202 VGND.n1201 4.5005
R4528 VGND.n1196 VGND.n1003 4.5005
R4529 VGND.n1215 VGND.n1214 4.5005
R4530 VGND.n1250 VGND.n1249 4.5005
R4531 VGND.n1223 VGND.n916 4.5005
R4532 VGND.n1242 VGND.n917 4.5005
R4533 VGND.n1228 VGND.n921 4.5005
R4534 VGND.n1235 VGND.n922 4.5005
R4535 VGND.n1272 VGND.n1271 4.5005
R4536 VGND.n997 VGND.n993 4.5005
R4537 VGND.n1283 VGND.n1282 4.5005
R4538 VGND.n1157 VGND.n1156 4.41365
R4539 VGND VGND.n33 4.35375
R4540 VGND.n1134 VGND.n1133 4.05427
R4541 VGND.n507 VGND.n0 4.05427
R4542 VGND.n2218 VGND.n2217 4.05427
R4543 VGND.n2220 VGND.n2219 4.05427
R4544 VGND.n1358 VGND.n543 4.05427
R4545 VGND VGND.n3002 3.99438
R4546 VGND VGND.n32 3.99438
R4547 VGND.n125 VGND 3.99438
R4548 VGND VGND.n126 3.99438
R4549 VGND.n3001 VGND 3.99437
R4550 VGND.n1284 VGND.n223 3.77268
R4551 VGND.n2940 VGND.n206 3.77268
R4552 VGND.n1163 VGND.n1162 3.77268
R4553 VGND.n2634 VGND.n2633 3.77268
R4554 VGND.n1327 VGND.n1326 3.77268
R4555 VGND.n2691 VGND.n2690 3.77268
R4556 VGND.n1323 VGND.n898 3.77268
R4557 VGND.n2689 VGND.n2688 3.77268
R4558 VGND.n1318 VGND.n901 3.77268
R4559 VGND.n2685 VGND.n2684 3.77268
R4560 VGND.n1315 VGND.n904 3.77268
R4561 VGND.n2683 VGND.n2682 3.77268
R4562 VGND.n1310 VGND.n907 3.77268
R4563 VGND.n2679 VGND.n2678 3.77268
R4564 VGND.n1307 VGND.n910 3.77268
R4565 VGND.n2677 VGND.n2676 3.77268
R4566 VGND.n1302 VGND.n913 3.77268
R4567 VGND.n2710 VGND.n2709 3.77268
R4568 VGND.n1299 VGND.n1298 3.77268
R4569 VGND.n2723 VGND.n2722 3.77268
R4570 VGND.n1297 VGND.n1296 3.77268
R4571 VGND.n2743 VGND.n2742 3.77268
R4572 VGND.n1293 VGND.n1292 3.77268
R4573 VGND.n2761 VGND.n2760 3.77268
R4574 VGND.n1291 VGND.n1290 3.77268
R4575 VGND.n2782 VGND.n2781 3.77268
R4576 VGND.n1270 VGND.n229 3.77268
R4577 VGND.n2780 VGND.n281 3.77268
R4578 VGND.n1286 VGND.n1285 3.77268
R4579 VGND.n2795 VGND.n284 3.77268
R4580 VGND.n1329 VGND.n1328 3.77268
R4581 VGND.n2695 VGND.n2694 3.77268
R4582 VGND.n2769 VGND.n205 3.75914
R4583 VGND.n2631 VGND.n2629 3.75914
R4584 VGND.n1267 VGND.n995 3.75914
R4585 VGND.n1022 VGND.n1020 3.75914
R4586 VGND.n2771 VGND.n284 3.4105
R4587 VGND.n2780 VGND.n2779 3.4105
R4588 VGND.n2781 VGND.n289 3.4105
R4589 VGND.n2762 VGND.n2761 3.4105
R4590 VGND.n2742 VGND.n2741 3.4105
R4591 VGND.n2724 VGND.n2723 3.4105
R4592 VGND.n2709 VGND.n2708 3.4105
R4593 VGND.n2677 VGND.n390 3.4105
R4594 VGND.n2678 VGND.n352 3.4105
R4595 VGND.n2683 VGND.n347 3.4105
R4596 VGND.n2684 VGND.n346 3.4105
R4597 VGND.n2689 VGND.n341 3.4105
R4598 VGND.n2690 VGND.n340 3.4105
R4599 VGND.n2696 VGND.n2695 3.4105
R4600 VGND.n2941 VGND.n2940 3.4105
R4601 VGND.n2770 VGND.n2769 3.4105
R4602 VGND.n2768 VGND.n291 3.4105
R4603 VGND.n2767 VGND.n2766 3.4105
R4604 VGND.n2764 VGND.n2763 3.4105
R4605 VGND.n307 VGND.n298 3.4105
R4606 VGND.n2609 VGND.n316 3.4105
R4607 VGND.n2610 VGND.n323 3.4105
R4608 VGND.n2613 VGND.n2612 3.4105
R4609 VGND.n2616 VGND.n2615 3.4105
R4610 VGND.n2619 VGND.n2618 3.4105
R4611 VGND.n2622 VGND.n2621 3.4105
R4612 VGND.n2625 VGND.n2624 3.4105
R4613 VGND.n2628 VGND.n2627 3.4105
R4614 VGND.n2629 VGND.n335 3.4105
R4615 VGND.n2633 VGND.n2632 3.4105
R4616 VGND.n2937 VGND.n206 3.4105
R4617 VGND.n2635 VGND.n2634 3.4105
R4618 VGND.n2559 VGND.n397 3.4105
R4619 VGND.n2533 VGND.n2532 3.4105
R4620 VGND.n2557 VGND.n339 3.4105
R4621 VGND.n2692 VGND.n2691 3.4105
R4622 VGND.n2384 VGND.n2383 3.4105
R4623 VGND.n2358 VGND.n2357 3.4105
R4624 VGND.n2531 VGND.n2530 3.4105
R4625 VGND.n2399 VGND.n2398 3.4105
R4626 VGND.n2556 VGND.n342 3.4105
R4627 VGND.n2688 VGND.n2687 3.4105
R4628 VGND.n2397 VGND.n2396 3.4105
R4629 VGND.n2386 VGND.n2385 3.4105
R4630 VGND.n2360 VGND.n2359 3.4105
R4631 VGND.n2818 VGND.n274 3.4105
R4632 VGND.n2412 VGND.n2411 3.4105
R4633 VGND.n2410 VGND.n2409 3.4105
R4634 VGND.n2555 VGND.n345 3.4105
R4635 VGND.n2686 VGND.n2685 3.4105
R4636 VGND.n1929 VGND.n449 3.4105
R4637 VGND.n1928 VGND.n453 3.4105
R4638 VGND.n1918 VGND.n457 3.4105
R4639 VGND.n1907 VGND.n467 3.4105
R4640 VGND.n1990 VGND.n604 3.4105
R4641 VGND.n1939 VGND.n445 3.4105
R4642 VGND.n2423 VGND.n2422 3.4105
R4643 VGND.n2425 VGND.n2424 3.4105
R4644 VGND.n2554 VGND.n348 3.4105
R4645 VGND.n2682 VGND.n2681 3.4105
R4646 VGND.n2158 VGND.n2157 3.4105
R4647 VGND.n2160 VGND.n2159 3.4105
R4648 VGND.n2166 VGND.n2165 3.4105
R4649 VGND.n2168 VGND.n2167 3.4105
R4650 VGND.n2064 VGND.n2063 3.4105
R4651 VGND.n1997 VGND.n603 3.4105
R4652 VGND.n2152 VGND.n2151 3.4105
R4653 VGND.n1940 VGND.n441 3.4105
R4654 VGND.n2438 VGND.n2437 3.4105
R4655 VGND.n2436 VGND.n2435 3.4105
R4656 VGND.n2553 VGND.n351 3.4105
R4657 VGND.n2680 VGND.n2679 3.4105
R4658 VGND.n2154 VGND.n2153 3.4105
R4659 VGND.n2156 VGND.n2155 3.4105
R4660 VGND.n2162 VGND.n2161 3.4105
R4661 VGND.n2164 VGND.n2163 3.4105
R4662 VGND.n2170 VGND.n2169 3.4105
R4663 VGND.n2066 VGND.n2065 3.4105
R4664 VGND.n2843 VGND.n262 3.4105
R4665 VGND.n2148 VGND.n2147 3.4105
R4666 VGND.n2150 VGND.n2149 3.4105
R4667 VGND.n1950 VGND.n437 3.4105
R4668 VGND.n2449 VGND.n2448 3.4105
R4669 VGND.n2451 VGND.n2450 3.4105
R4670 VGND.n2552 VGND.n391 3.4105
R4671 VGND.n2676 VGND.n2675 3.4105
R4672 VGND.n1790 VGND.n570 3.4105
R4673 VGND.n1780 VGND.n567 3.4105
R4674 VGND.n1779 VGND.n564 3.4105
R4675 VGND.n1769 VGND.n561 3.4105
R4676 VGND.n1768 VGND.n558 3.4105
R4677 VGND.n1758 VGND.n555 3.4105
R4678 VGND.n1901 VGND.n588 3.4105
R4679 VGND.n1830 VGND.n1737 3.4105
R4680 VGND.n1791 VGND.n573 3.4105
R4681 VGND.n2146 VGND.n2145 3.4105
R4682 VGND.n2144 VGND.n2143 3.4105
R4683 VGND.n1951 VGND.n433 3.4105
R4684 VGND.n2464 VGND.n2463 3.4105
R4685 VGND.n2462 VGND.n2461 3.4105
R4686 VGND.n2551 VGND.n321 3.4105
R4687 VGND.n2711 VGND.n2710 3.4105
R4688 VGND.n1867 VGND.n1866 3.4105
R4689 VGND.n1869 VGND.n1868 3.4105
R4690 VGND.n1875 VGND.n1874 3.4105
R4691 VGND.n1877 VGND.n1876 3.4105
R4692 VGND.n1883 VGND.n1882 3.4105
R4693 VGND.n1885 VGND.n1884 3.4105
R4694 VGND.n1686 VGND.n639 3.4105
R4695 VGND.n1899 VGND.n1898 3.4105
R4696 VGND.n1837 VGND.n1736 3.4105
R4697 VGND.n1861 VGND.n1860 3.4105
R4698 VGND.n1801 VGND.n576 3.4105
R4699 VGND.n2140 VGND.n2139 3.4105
R4700 VGND.n2142 VGND.n2141 3.4105
R4701 VGND.n1961 VGND.n429 3.4105
R4702 VGND.n2475 VGND.n2474 3.4105
R4703 VGND.n2477 VGND.n2476 3.4105
R4704 VGND.n2550 VGND.n317 3.4105
R4705 VGND.n2722 VGND.n2721 3.4105
R4706 VGND.n1863 VGND.n1862 3.4105
R4707 VGND.n1865 VGND.n1864 3.4105
R4708 VGND.n1871 VGND.n1870 3.4105
R4709 VGND.n1873 VGND.n1872 3.4105
R4710 VGND.n1879 VGND.n1878 3.4105
R4711 VGND.n1881 VGND.n1880 3.4105
R4712 VGND.n1887 VGND.n1886 3.4105
R4713 VGND.n1889 VGND.n1888 3.4105
R4714 VGND.n1897 VGND.n1896 3.4105
R4715 VGND.n2868 VGND.n250 3.4105
R4716 VGND.n1857 VGND.n1856 3.4105
R4717 VGND.n1859 VGND.n1858 3.4105
R4718 VGND.n1802 VGND.n579 3.4105
R4719 VGND.n2138 VGND.n2137 3.4105
R4720 VGND.n2136 VGND.n2135 3.4105
R4721 VGND.n1962 VGND.n425 3.4105
R4722 VGND.n2490 VGND.n2489 3.4105
R4723 VGND.n2488 VGND.n2487 3.4105
R4724 VGND.n2549 VGND.n305 3.4105
R4725 VGND.n2744 VGND.n2743 3.4105
R4726 VGND.n860 VGND.n663 3.4105
R4727 VGND.n861 VGND.n660 3.4105
R4728 VGND.n862 VGND.n657 3.4105
R4729 VGND.n863 VGND.n654 3.4105
R4730 VGND.n864 VGND.n651 3.4105
R4731 VGND.n865 VGND.n648 3.4105
R4732 VGND.n866 VGND.n645 3.4105
R4733 VGND.n867 VGND.n642 3.4105
R4734 VGND.n1891 VGND.n1890 3.4105
R4735 VGND.n1349 VGND.n630 3.4105
R4736 VGND.n1654 VGND.n737 3.4105
R4737 VGND.n1670 VGND.n1669 3.4105
R4738 VGND.n1855 VGND.n1854 3.4105
R4739 VGND.n1853 VGND.n1852 3.4105
R4740 VGND.n1812 VGND.n582 3.4105
R4741 VGND.n2132 VGND.n2131 3.4105
R4742 VGND.n2134 VGND.n2133 3.4105
R4743 VGND.n1972 VGND.n421 3.4105
R4744 VGND.n2506 VGND.n2505 3.4105
R4745 VGND.n2508 VGND.n2507 3.4105
R4746 VGND.n2548 VGND.n301 3.4105
R4747 VGND.n2760 VGND.n2759 3.4105
R4748 VGND.n1629 VGND.n731 3.4105
R4749 VGND.n1628 VGND.n1627 3.4105
R4750 VGND.n1559 VGND.n753 3.4105
R4751 VGND.n1561 VGND.n1560 3.4105
R4752 VGND.n1539 VGND.n1538 3.4105
R4753 VGND.n1524 VGND.n1523 3.4105
R4754 VGND.n1513 VGND.n1512 3.4105
R4755 VGND.n1498 VGND.n1497 3.4105
R4756 VGND.n1487 VGND.n1486 3.4105
R4757 VGND.n1402 VGND.n638 3.4105
R4758 VGND.n1405 VGND.n1404 3.4105
R4759 VGND.n1651 VGND.n738 3.4105
R4760 VGND.n2878 VGND.n2877 3.4105
R4761 VGND.n1668 VGND.n242 3.4105
R4762 VGND.n2855 VGND.n2854 3.4105
R4763 VGND.n2853 VGND.n2852 3.4105
R4764 VGND.n1813 VGND.n254 3.4105
R4765 VGND.n2830 VGND.n2829 3.4105
R4766 VGND.n2828 VGND.n2827 3.4105
R4767 VGND.n1973 VGND.n266 3.4105
R4768 VGND.n2805 VGND.n2804 3.4105
R4769 VGND.n2803 VGND.n2802 3.4105
R4770 VGND.n2547 VGND.n278 3.4105
R4771 VGND.n2783 VGND.n2782 3.4105
R4772 VGND.n2880 VGND.n2879 3.4105
R4773 VGND.n1624 VGND.n1623 3.4105
R4774 VGND.n1626 VGND.n1625 3.4105
R4775 VGND.n1589 VGND.n1588 3.4105
R4776 VGND.n1563 VGND.n1562 3.4105
R4777 VGND.n1537 VGND.n1536 3.4105
R4778 VGND.n1526 VGND.n1525 3.4105
R4779 VGND.n1511 VGND.n1510 3.4105
R4780 VGND.n1500 VGND.n1499 3.4105
R4781 VGND.n1485 VGND.n1484 3.4105
R4782 VGND.n1474 VGND.n1473 3.4105
R4783 VGND.n1407 VGND.n1406 3.4105
R4784 VGND.n2893 VGND.n237 3.4105
R4785 VGND.n2881 VGND.n230 3.4105
R4786 VGND.n2876 VGND.n2875 3.4105
R4787 VGND.n2874 VGND.n2873 3.4105
R4788 VGND.n2856 VGND.n245 3.4105
R4789 VGND.n2851 VGND.n2850 3.4105
R4790 VGND.n2849 VGND.n2848 3.4105
R4791 VGND.n2831 VGND.n257 3.4105
R4792 VGND.n2826 VGND.n2825 3.4105
R4793 VGND.n2824 VGND.n2823 3.4105
R4794 VGND.n2806 VGND.n269 3.4105
R4795 VGND.n2801 VGND.n2800 3.4105
R4796 VGND.n2799 VGND.n2798 3.4105
R4797 VGND.n2784 VGND.n281 3.4105
R4798 VGND.n2899 VGND.n2898 3.4105
R4799 VGND.n1620 VGND.n241 3.4105
R4800 VGND.n1622 VGND.n1621 3.4105
R4801 VGND.n1592 VGND.n743 3.4105
R4802 VGND.n1591 VGND.n1590 3.4105
R4803 VGND.n1465 VGND.n757 3.4105
R4804 VGND.n1466 VGND.n762 3.4105
R4805 VGND.n1467 VGND.n766 3.4105
R4806 VGND.n1468 VGND.n770 3.4105
R4807 VGND.n1469 VGND.n774 3.4105
R4808 VGND.n1470 VGND.n778 3.4105
R4809 VGND.n1472 VGND.n1471 3.4105
R4810 VGND.n1344 VGND.n798 3.4105
R4811 VGND.n1606 VGND.n1605 3.4105
R4812 VGND.n2897 VGND.n2896 3.4105
R4813 VGND.n2895 VGND.n2894 3.4105
R4814 VGND.n740 VGND.n235 3.4105
R4815 VGND.n2872 VGND.n2871 3.4105
R4816 VGND.n2870 VGND.n2869 3.4105
R4817 VGND.n1838 VGND.n248 3.4105
R4818 VGND.n2847 VGND.n2846 3.4105
R4819 VGND.n2845 VGND.n2844 3.4105
R4820 VGND.n1998 VGND.n260 3.4105
R4821 VGND.n2822 VGND.n2821 3.4105
R4822 VGND.n2820 VGND.n2819 3.4105
R4823 VGND.n419 VGND.n272 3.4105
R4824 VGND.n2797 VGND.n2796 3.4105
R4825 VGND.n2795 VGND.n2794 3.4105
R4826 VGND.n234 VGND.n233 3.4105
R4827 VGND.n2901 VGND.n2900 3.4105
R4828 VGND.n1064 VGND.n923 3.4105
R4829 VGND.n1065 VGND.n746 3.4105
R4830 VGND.n1066 VGND.n918 3.4105
R4831 VGND.n1067 VGND.n752 3.4105
R4832 VGND.n1304 VGND.n1303 3.4105
R4833 VGND.n1306 VGND.n1305 3.4105
R4834 VGND.n1312 VGND.n1311 3.4105
R4835 VGND.n1314 VGND.n1313 3.4105
R4836 VGND.n1320 VGND.n1319 3.4105
R4837 VGND.n1322 VGND.n1321 3.4105
R4838 VGND.n1101 VGND.n782 3.4105
R4839 VGND.n1104 VGND.n1103 3.4105
R4840 VGND.n2913 VGND.n226 3.4105
R4841 VGND.n1102 VGND.n792 3.4105
R4842 VGND.n1420 VGND.n1419 3.4105
R4843 VGND.n1418 VGND.n1417 3.4105
R4844 VGND.n1403 VGND.n635 3.4105
R4845 VGND.n1893 VGND.n1892 3.4105
R4846 VGND.n1895 VGND.n1894 3.4105
R4847 VGND.n1685 VGND.n551 3.4105
R4848 VGND.n2174 VGND.n2173 3.4105
R4849 VGND.n2172 VGND.n2171 3.4105
R4850 VGND.n2062 VGND.n552 3.4105
R4851 VGND.n1917 VGND.n461 3.4105
R4852 VGND.n2371 VGND.n2370 3.4105
R4853 VGND.n2373 VGND.n2372 3.4105
R4854 VGND.n2558 VGND.n336 3.4105
R4855 VGND.n2694 VGND.n2693 3.4105
R4856 VGND.n1285 VGND.n993 3.4105
R4857 VGND.n1271 VGND.n1270 3.4105
R4858 VGND.n1291 VGND.n922 3.4105
R4859 VGND.n1292 VGND.n921 3.4105
R4860 VGND.n1297 VGND.n917 3.4105
R4861 VGND.n1298 VGND.n916 3.4105
R4862 VGND.n1250 VGND.n913 3.4105
R4863 VGND.n1214 VGND.n910 3.4105
R4864 VGND.n1196 VGND.n907 3.4105
R4865 VGND.n1201 VGND.n904 3.4105
R4866 VGND.n1192 VGND.n901 3.4105
R4867 VGND.n1182 VGND.n898 3.4105
R4868 VGND.n1327 VGND.n892 3.4105
R4869 VGND.n1328 VGND.n891 3.4105
R4870 VGND.n1284 VGND.n1283 3.4105
R4871 VGND.n1267 VGND.n1266 3.4105
R4872 VGND.n1269 VGND.n1268 3.4105
R4873 VGND.n1264 VGND.n1263 3.4105
R4874 VGND.n1261 VGND.n1260 3.4105
R4875 VGND.n1258 VGND.n1257 3.4105
R4876 VGND.n1255 VGND.n1254 3.4105
R4877 VGND.n1252 VGND.n1251 3.4105
R4878 VGND.n1213 VGND.n999 3.4105
R4879 VGND.n1198 VGND.n1197 3.4105
R4880 VGND.n1200 VGND.n1199 3.4105
R4881 VGND.n1194 VGND.n1193 3.4105
R4882 VGND.n1181 VGND.n1005 3.4105
R4883 VGND.n1017 VGND.n1016 3.4105
R4884 VGND.n1020 VGND.n1019 3.4105
R4885 VGND.n1164 VGND.n1163 3.4105
R4886 VGND.n1287 VGND.n1286 3.4105
R4887 VGND.n1288 VGND.n229 3.4105
R4888 VGND.n1290 VGND.n1289 3.4105
R4889 VGND.n1294 VGND.n1293 3.4105
R4890 VGND.n1296 VGND.n1295 3.4105
R4891 VGND.n1300 VGND.n1299 3.4105
R4892 VGND.n1302 VGND.n1301 3.4105
R4893 VGND.n1308 VGND.n1307 3.4105
R4894 VGND.n1310 VGND.n1309 3.4105
R4895 VGND.n1316 VGND.n1315 3.4105
R4896 VGND.n1318 VGND.n1317 3.4105
R4897 VGND.n1324 VGND.n1323 3.4105
R4898 VGND.n1326 VGND.n1325 3.4105
R4899 VGND.n1330 VGND.n1329 3.4105
R4900 VGND.n1162 VGND.n1161 3.4105
R4901 VGND.n2916 VGND.n223 3.4105
R4902 VGND.n105 VGND.n104 3.01226
R4903 VGND.n2200 VGND.n2189 3.01226
R4904 VGND.n2184 VGND.n545 2.63579
R4905 VGND.n2565 VGND 2.52282
R4906 VGND.n2568 VGND 2.52282
R4907 VGND.n2571 VGND 2.52282
R4908 VGND.n2574 VGND 2.52282
R4909 VGND.n2577 VGND 2.52282
R4910 VGND.n2580 VGND 2.52282
R4911 VGND.n2583 VGND 2.52282
R4912 VGND.n2586 VGND 2.52282
R4913 VGND.n2589 VGND 2.52282
R4914 VGND.n2592 VGND 2.52282
R4915 VGND.n2595 VGND 2.52282
R4916 VGND.n2598 VGND 2.52282
R4917 VGND.n2601 VGND 2.52282
R4918 VGND.n2604 VGND 2.52282
R4919 VGND.n2607 VGND 2.52282
R4920 VGND.n186 VGND.n185 2.25932
R4921 VGND.n114 VGND.n93 2.25932
R4922 VGND.n110 VGND.n109 2.25932
R4923 VGND.n87 VGND.n86 2.25932
R4924 VGND.n155 VGND.n154 2.25932
R4925 VGND.n2205 VGND.n2204 2.25932
R4926 VGND.n491 VGND.n479 1.88285
R4927 VGND.n2272 VGND.n2260 1.88285
R4928 VGND.n527 VGND.n515 1.88285
R4929 VGND.n2608 VGND 1.79514
R4930 VGND.n1158 VGND.n224 1.76378
R4931 VGND.n2608 VGND 1.57193
R4932 VGND.n2940 VGND.n2939 1.54254
R4933 VGND.n2938 VGND.n2937 1.54254
R4934 VGND.n2533 VGND.n207 1.54254
R4935 VGND.n2530 VGND.n417 1.54254
R4936 VGND.n2818 VGND.n275 1.54254
R4937 VGND.n1991 VGND.n1990 1.54254
R4938 VGND.n1997 VGND.n1992 1.54254
R4939 VGND.n2843 VGND.n263 1.54254
R4940 VGND.n1831 VGND.n1830 1.54254
R4941 VGND.n1837 VGND.n1832 1.54254
R4942 VGND.n2868 VGND.n251 1.54254
R4943 VGND.n1654 VGND.n1653 1.54254
R4944 VGND.n1652 VGND.n1651 1.54254
R4945 VGND.n2893 VGND.n238 1.54254
R4946 VGND.n1606 VGND.n225 1.54254
R4947 VGND.n2914 VGND.n2913 1.54254
R4948 VGND.n1284 VGND.n224 1.54254
R4949 VGND.n2916 VGND.n2915 1.54254
R4950 VGND.n121 VGND.n120 1.50638
R4951 VGND.n2212 VGND.n544 1.50638
R4952 VGND VGND.n2562 1.3946
R4953 VGND.n2561 VGND 1.3946
R4954 VGND.n2560 VGND 1.3946
R4955 VGND VGND.n398 1.3946
R4956 VGND.n1905 VGND 1.3946
R4957 VGND VGND.n1906 1.3946
R4958 VGND.n1904 VGND 1.3946
R4959 VGND.n1903 VGND 1.3946
R4960 VGND.n1902 VGND 1.3946
R4961 VGND.n1900 VGND 1.3946
R4962 VGND VGND.n626 1.3946
R4963 VGND VGND.n1348 1.3946
R4964 VGND.n1347 VGND 1.3946
R4965 VGND.n1346 VGND 1.3946
R4966 VGND.n1345 VGND 1.3946
R4967 VGND VGND.n880 1.3946
R4968 VGND.n1159 VGND 1.3946
R4969 VGND VGND.n1160 1.3946
R4970 VGND.n1158 VGND.n1157 1.04899
R4971 VGND.n2696 VGND.n335 1.00149
R4972 VGND.n2627 VGND.n340 1.00149
R4973 VGND.n2624 VGND.n341 1.00149
R4974 VGND.n2621 VGND.n346 1.00149
R4975 VGND.n2618 VGND.n347 1.00149
R4976 VGND.n2615 VGND.n352 1.00149
R4977 VGND.n2612 VGND.n390 1.00149
R4978 VGND.n2708 VGND.n323 1.00149
R4979 VGND.n2724 VGND.n316 1.00149
R4980 VGND.n2741 VGND.n307 1.00149
R4981 VGND.n2763 VGND.n2762 1.00149
R4982 VGND.n2766 VGND.n289 1.00149
R4983 VGND.n2779 VGND.n291 1.00149
R4984 VGND.n2771 VGND.n2770 1.00149
R4985 VGND.n2941 VGND.n205 1.00149
R4986 VGND.n1019 VGND.n891 1.00149
R4987 VGND.n1016 VGND.n892 1.00149
R4988 VGND.n1182 VGND.n1181 1.00149
R4989 VGND.n1193 VGND.n1192 1.00149
R4990 VGND.n1201 VGND.n1200 1.00149
R4991 VGND.n1197 VGND.n1196 1.00149
R4992 VGND.n1214 VGND.n1213 1.00149
R4993 VGND.n1251 VGND.n1250 1.00149
R4994 VGND.n1254 VGND.n916 1.00149
R4995 VGND.n1257 VGND.n917 1.00149
R4996 VGND.n1260 VGND.n921 1.00149
R4997 VGND.n1263 VGND.n922 1.00149
R4998 VGND.n1271 VGND.n1269 1.00149
R4999 VGND.n1266 VGND.n993 1.00149
R5000 VGND.n1283 VGND.n995 1.00149
R5001 VGND.n1164 VGND.n1022 1.00149
R5002 VGND.n2632 VGND.n2631 0.973133
R5003 VGND.n2346 VGND.n2 0.9305
R5004 VGND.n178 VGND.n174 0.929432
R5005 VGND.n101 VGND.n99 0.929432
R5006 VGND.n79 VGND.n75 0.929432
R5007 VGND.n147 VGND.n143 0.929432
R5008 VGND.n126 VGND.n1 0.916608
R5009 VGND VGND.n2565 0.839786
R5010 VGND VGND.n2568 0.839786
R5011 VGND VGND.n2571 0.839786
R5012 VGND VGND.n2574 0.839786
R5013 VGND VGND.n2577 0.839786
R5014 VGND VGND.n2580 0.839786
R5015 VGND VGND.n2583 0.839786
R5016 VGND VGND.n2586 0.839786
R5017 VGND VGND.n2589 0.839786
R5018 VGND VGND.n2592 0.839786
R5019 VGND VGND.n2595 0.839786
R5020 VGND VGND.n2598 0.839786
R5021 VGND VGND.n2601 0.839786
R5022 VGND VGND.n2604 0.839786
R5023 VGND VGND.n2607 0.839786
R5024 VGND.n3023 VGND.n3022 0.7755
R5025 VGND.n3024 VGND.n3023 0.774207
R5026 VGND.n2981 VGND.n2978 0.753441
R5027 VGND.n20 VGND.n18 0.753441
R5028 VGND.n2953 VGND.n2951 0.753441
R5029 VGND.n46 VGND.n44 0.753441
R5030 VGND.n159 VGND.n136 0.753441
R5031 VGND.n2254 VGND.n2252 0.753441
R5032 VGND.n3025 VGND 0.706681
R5033 VGND VGND.n0 0.542567
R5034 VGND.n3025 VGND.n1 0.507317
R5035 VGND.n2939 VGND.n33 0.404308
R5036 VGND.n115 VGND.n114 0.376971
R5037 VGND.n120 VGND.n92 0.376971
R5038 VGND.n1140 VGND.n1137 0.376971
R5039 VGND.n1112 VGND.n1108 0.376971
R5040 VGND.n2212 VGND.n2211 0.376971
R5041 VGND.n2237 VGND.n2236 0.376971
R5042 VGND.n1375 VGND.n1374 0.376971
R5043 VGND VGND.n3025 0.37415
R5044 VGND.n226 VGND.n223 0.362676
R5045 VGND.n1605 VGND.n226 0.362676
R5046 VGND.n1605 VGND.n237 0.362676
R5047 VGND.n738 VGND.n237 0.362676
R5048 VGND.n738 VGND.n737 0.362676
R5049 VGND.n737 VGND.n250 0.362676
R5050 VGND.n1736 VGND.n250 0.362676
R5051 VGND.n1737 VGND.n1736 0.362676
R5052 VGND.n1737 VGND.n262 0.362676
R5053 VGND.n603 VGND.n262 0.362676
R5054 VGND.n604 VGND.n603 0.362676
R5055 VGND.n604 VGND.n274 0.362676
R5056 VGND.n2531 VGND.n274 0.362676
R5057 VGND.n2532 VGND.n2531 0.362676
R5058 VGND.n2532 VGND.n206 0.362676
R5059 VGND.n1162 VGND.n1104 0.362676
R5060 VGND.n1104 VGND.n798 0.362676
R5061 VGND.n1406 VGND.n798 0.362676
R5062 VGND.n1406 VGND.n1405 0.362676
R5063 VGND.n1405 VGND.n630 0.362676
R5064 VGND.n1897 VGND.n630 0.362676
R5065 VGND.n1898 VGND.n1897 0.362676
R5066 VGND.n1898 VGND.n588 0.362676
R5067 VGND.n2065 VGND.n588 0.362676
R5068 VGND.n2065 VGND.n2064 0.362676
R5069 VGND.n2064 VGND.n467 0.362676
R5070 VGND.n2359 VGND.n467 0.362676
R5071 VGND.n2359 VGND.n2358 0.362676
R5072 VGND.n2358 VGND.n397 0.362676
R5073 VGND.n2634 VGND.n397 0.362676
R5074 VGND.n1326 VGND.n782 0.362676
R5075 VGND.n1472 VGND.n782 0.362676
R5076 VGND.n1473 VGND.n1472 0.362676
R5077 VGND.n1473 VGND.n638 0.362676
R5078 VGND.n1890 VGND.n638 0.362676
R5079 VGND.n1890 VGND.n1889 0.362676
R5080 VGND.n1889 VGND.n639 0.362676
R5081 VGND.n639 VGND.n555 0.362676
R5082 VGND.n2169 VGND.n555 0.362676
R5083 VGND.n2169 VGND.n2168 0.362676
R5084 VGND.n2168 VGND.n457 0.362676
R5085 VGND.n2385 VGND.n457 0.362676
R5086 VGND.n2385 VGND.n2384 0.362676
R5087 VGND.n2384 VGND.n339 0.362676
R5088 VGND.n2691 VGND.n339 0.362676
R5089 VGND.n1323 VGND.n1322 0.362676
R5090 VGND.n1322 VGND.n778 0.362676
R5091 VGND.n1485 VGND.n778 0.362676
R5092 VGND.n1486 VGND.n1485 0.362676
R5093 VGND.n1486 VGND.n642 0.362676
R5094 VGND.n1886 VGND.n642 0.362676
R5095 VGND.n1886 VGND.n1885 0.362676
R5096 VGND.n1885 VGND.n558 0.362676
R5097 VGND.n2164 VGND.n558 0.362676
R5098 VGND.n2165 VGND.n2164 0.362676
R5099 VGND.n2165 VGND.n453 0.362676
R5100 VGND.n2397 VGND.n453 0.362676
R5101 VGND.n2398 VGND.n2397 0.362676
R5102 VGND.n2398 VGND.n342 0.362676
R5103 VGND.n2688 VGND.n342 0.362676
R5104 VGND.n1319 VGND.n1318 0.362676
R5105 VGND.n1319 VGND.n774 0.362676
R5106 VGND.n1499 VGND.n774 0.362676
R5107 VGND.n1499 VGND.n1498 0.362676
R5108 VGND.n1498 VGND.n645 0.362676
R5109 VGND.n1881 VGND.n645 0.362676
R5110 VGND.n1882 VGND.n1881 0.362676
R5111 VGND.n1882 VGND.n561 0.362676
R5112 VGND.n2161 VGND.n561 0.362676
R5113 VGND.n2161 VGND.n2160 0.362676
R5114 VGND.n2160 VGND.n449 0.362676
R5115 VGND.n2411 VGND.n449 0.362676
R5116 VGND.n2411 VGND.n2410 0.362676
R5117 VGND.n2410 VGND.n345 0.362676
R5118 VGND.n2685 VGND.n345 0.362676
R5119 VGND.n1315 VGND.n1314 0.362676
R5120 VGND.n1314 VGND.n770 0.362676
R5121 VGND.n1511 VGND.n770 0.362676
R5122 VGND.n1512 VGND.n1511 0.362676
R5123 VGND.n1512 VGND.n648 0.362676
R5124 VGND.n1878 VGND.n648 0.362676
R5125 VGND.n1878 VGND.n1877 0.362676
R5126 VGND.n1877 VGND.n564 0.362676
R5127 VGND.n2156 VGND.n564 0.362676
R5128 VGND.n2157 VGND.n2156 0.362676
R5129 VGND.n2157 VGND.n445 0.362676
R5130 VGND.n2423 VGND.n445 0.362676
R5131 VGND.n2424 VGND.n2423 0.362676
R5132 VGND.n2424 VGND.n348 0.362676
R5133 VGND.n2682 VGND.n348 0.362676
R5134 VGND.n1311 VGND.n1310 0.362676
R5135 VGND.n1311 VGND.n766 0.362676
R5136 VGND.n1525 VGND.n766 0.362676
R5137 VGND.n1525 VGND.n1524 0.362676
R5138 VGND.n1524 VGND.n651 0.362676
R5139 VGND.n1873 VGND.n651 0.362676
R5140 VGND.n1874 VGND.n1873 0.362676
R5141 VGND.n1874 VGND.n567 0.362676
R5142 VGND.n2153 VGND.n567 0.362676
R5143 VGND.n2153 VGND.n2152 0.362676
R5144 VGND.n2152 VGND.n441 0.362676
R5145 VGND.n2437 VGND.n441 0.362676
R5146 VGND.n2437 VGND.n2436 0.362676
R5147 VGND.n2436 VGND.n351 0.362676
R5148 VGND.n2679 VGND.n351 0.362676
R5149 VGND.n1307 VGND.n1306 0.362676
R5150 VGND.n1306 VGND.n762 0.362676
R5151 VGND.n1537 VGND.n762 0.362676
R5152 VGND.n1538 VGND.n1537 0.362676
R5153 VGND.n1538 VGND.n654 0.362676
R5154 VGND.n1870 VGND.n654 0.362676
R5155 VGND.n1870 VGND.n1869 0.362676
R5156 VGND.n1869 VGND.n570 0.362676
R5157 VGND.n2148 VGND.n570 0.362676
R5158 VGND.n2149 VGND.n2148 0.362676
R5159 VGND.n2149 VGND.n437 0.362676
R5160 VGND.n2449 VGND.n437 0.362676
R5161 VGND.n2450 VGND.n2449 0.362676
R5162 VGND.n2450 VGND.n391 0.362676
R5163 VGND.n2676 VGND.n391 0.362676
R5164 VGND.n1303 VGND.n1302 0.362676
R5165 VGND.n1303 VGND.n757 0.362676
R5166 VGND.n1562 VGND.n757 0.362676
R5167 VGND.n1562 VGND.n1561 0.362676
R5168 VGND.n1561 VGND.n657 0.362676
R5169 VGND.n1865 VGND.n657 0.362676
R5170 VGND.n1866 VGND.n1865 0.362676
R5171 VGND.n1866 VGND.n573 0.362676
R5172 VGND.n2145 VGND.n573 0.362676
R5173 VGND.n2145 VGND.n2144 0.362676
R5174 VGND.n2144 VGND.n433 0.362676
R5175 VGND.n2463 VGND.n433 0.362676
R5176 VGND.n2463 VGND.n2462 0.362676
R5177 VGND.n2462 VGND.n321 0.362676
R5178 VGND.n2710 VGND.n321 0.362676
R5179 VGND.n1299 VGND.n752 0.362676
R5180 VGND.n1590 VGND.n752 0.362676
R5181 VGND.n1590 VGND.n1589 0.362676
R5182 VGND.n1589 VGND.n753 0.362676
R5183 VGND.n753 VGND.n660 0.362676
R5184 VGND.n1862 VGND.n660 0.362676
R5185 VGND.n1862 VGND.n1861 0.362676
R5186 VGND.n1861 VGND.n576 0.362676
R5187 VGND.n2140 VGND.n576 0.362676
R5188 VGND.n2141 VGND.n2140 0.362676
R5189 VGND.n2141 VGND.n429 0.362676
R5190 VGND.n2475 VGND.n429 0.362676
R5191 VGND.n2476 VGND.n2475 0.362676
R5192 VGND.n2476 VGND.n317 0.362676
R5193 VGND.n2722 VGND.n317 0.362676
R5194 VGND.n1296 VGND.n918 0.362676
R5195 VGND.n918 VGND.n743 0.362676
R5196 VGND.n1626 VGND.n743 0.362676
R5197 VGND.n1627 VGND.n1626 0.362676
R5198 VGND.n1627 VGND.n663 0.362676
R5199 VGND.n1857 VGND.n663 0.362676
R5200 VGND.n1858 VGND.n1857 0.362676
R5201 VGND.n1858 VGND.n579 0.362676
R5202 VGND.n2137 VGND.n579 0.362676
R5203 VGND.n2137 VGND.n2136 0.362676
R5204 VGND.n2136 VGND.n425 0.362676
R5205 VGND.n2489 VGND.n425 0.362676
R5206 VGND.n2489 VGND.n2488 0.362676
R5207 VGND.n2488 VGND.n305 0.362676
R5208 VGND.n2743 VGND.n305 0.362676
R5209 VGND.n1293 VGND.n746 0.362676
R5210 VGND.n1622 VGND.n746 0.362676
R5211 VGND.n1623 VGND.n1622 0.362676
R5212 VGND.n1623 VGND.n731 0.362676
R5213 VGND.n1670 VGND.n731 0.362676
R5214 VGND.n1854 VGND.n1670 0.362676
R5215 VGND.n1854 VGND.n1853 0.362676
R5216 VGND.n1853 VGND.n582 0.362676
R5217 VGND.n2132 VGND.n582 0.362676
R5218 VGND.n2133 VGND.n2132 0.362676
R5219 VGND.n2133 VGND.n421 0.362676
R5220 VGND.n2506 VGND.n421 0.362676
R5221 VGND.n2507 VGND.n2506 0.362676
R5222 VGND.n2507 VGND.n301 0.362676
R5223 VGND.n2760 VGND.n301 0.362676
R5224 VGND.n1290 VGND.n923 0.362676
R5225 VGND.n923 VGND.n241 0.362676
R5226 VGND.n2879 VGND.n241 0.362676
R5227 VGND.n2879 VGND.n2878 0.362676
R5228 VGND.n2878 VGND.n242 0.362676
R5229 VGND.n2854 VGND.n242 0.362676
R5230 VGND.n2854 VGND.n2853 0.362676
R5231 VGND.n2853 VGND.n254 0.362676
R5232 VGND.n2829 VGND.n254 0.362676
R5233 VGND.n2829 VGND.n2828 0.362676
R5234 VGND.n2828 VGND.n266 0.362676
R5235 VGND.n2804 VGND.n266 0.362676
R5236 VGND.n2804 VGND.n2803 0.362676
R5237 VGND.n2803 VGND.n278 0.362676
R5238 VGND.n2782 VGND.n278 0.362676
R5239 VGND.n2900 VGND.n229 0.362676
R5240 VGND.n2900 VGND.n2899 0.362676
R5241 VGND.n2899 VGND.n230 0.362676
R5242 VGND.n2875 VGND.n230 0.362676
R5243 VGND.n2875 VGND.n2874 0.362676
R5244 VGND.n2874 VGND.n245 0.362676
R5245 VGND.n2850 VGND.n245 0.362676
R5246 VGND.n2850 VGND.n2849 0.362676
R5247 VGND.n2849 VGND.n257 0.362676
R5248 VGND.n2825 VGND.n257 0.362676
R5249 VGND.n2825 VGND.n2824 0.362676
R5250 VGND.n2824 VGND.n269 0.362676
R5251 VGND.n2800 VGND.n269 0.362676
R5252 VGND.n2800 VGND.n2799 0.362676
R5253 VGND.n2799 VGND.n281 0.362676
R5254 VGND.n1286 VGND.n234 0.362676
R5255 VGND.n2896 VGND.n234 0.362676
R5256 VGND.n2896 VGND.n2895 0.362676
R5257 VGND.n2895 VGND.n235 0.362676
R5258 VGND.n2871 VGND.n235 0.362676
R5259 VGND.n2871 VGND.n2870 0.362676
R5260 VGND.n2870 VGND.n248 0.362676
R5261 VGND.n2846 VGND.n248 0.362676
R5262 VGND.n2846 VGND.n2845 0.362676
R5263 VGND.n2845 VGND.n260 0.362676
R5264 VGND.n2821 VGND.n260 0.362676
R5265 VGND.n2821 VGND.n2820 0.362676
R5266 VGND.n2820 VGND.n272 0.362676
R5267 VGND.n2796 VGND.n272 0.362676
R5268 VGND.n2796 VGND.n2795 0.362676
R5269 VGND.n1329 VGND.n792 0.362676
R5270 VGND.n1419 VGND.n792 0.362676
R5271 VGND.n1419 VGND.n1418 0.362676
R5272 VGND.n1418 VGND.n635 0.362676
R5273 VGND.n1893 VGND.n635 0.362676
R5274 VGND.n1894 VGND.n1893 0.362676
R5275 VGND.n1894 VGND.n551 0.362676
R5276 VGND.n2173 VGND.n551 0.362676
R5277 VGND.n2173 VGND.n2172 0.362676
R5278 VGND.n2172 VGND.n552 0.362676
R5279 VGND.n552 VGND.n461 0.362676
R5280 VGND.n2371 VGND.n461 0.362676
R5281 VGND.n2372 VGND.n2371 0.362676
R5282 VGND.n2372 VGND.n336 0.362676
R5283 VGND.n2694 VGND.n336 0.362676
R5284 VGND.n2769 VGND.n2768 0.349144
R5285 VGND.n2768 VGND.n2767 0.349144
R5286 VGND.n2767 VGND.n2764 0.349144
R5287 VGND.n2764 VGND.n298 0.349144
R5288 VGND.n2609 VGND.n298 0.349144
R5289 VGND.n2610 VGND.n2609 0.349144
R5290 VGND.n2613 VGND.n2610 0.349144
R5291 VGND.n2616 VGND.n2613 0.349144
R5292 VGND.n2619 VGND.n2616 0.349144
R5293 VGND.n2622 VGND.n2619 0.349144
R5294 VGND.n2625 VGND.n2622 0.349144
R5295 VGND.n2628 VGND.n2625 0.349144
R5296 VGND.n2629 VGND.n2628 0.349144
R5297 VGND.n1268 VGND.n1267 0.349144
R5298 VGND.n1268 VGND.n1264 0.349144
R5299 VGND.n1264 VGND.n1261 0.349144
R5300 VGND.n1261 VGND.n1258 0.349144
R5301 VGND.n1258 VGND.n1255 0.349144
R5302 VGND.n1255 VGND.n1252 0.349144
R5303 VGND.n1252 VGND.n999 0.349144
R5304 VGND.n1198 VGND.n999 0.349144
R5305 VGND.n1199 VGND.n1198 0.349144
R5306 VGND.n1199 VGND.n1194 0.349144
R5307 VGND.n1194 VGND.n1005 0.349144
R5308 VGND.n1017 VGND.n1005 0.349144
R5309 VGND.n1020 VGND.n1017 0.349144
R5310 VGND.n2700 VGND.n331 0.327628
R5311 VGND.n2697 VGND.n333 0.327628
R5312 VGND.n361 VGND.n358 0.327628
R5313 VGND.n369 VGND.n365 0.327628
R5314 VGND.n372 VGND.n354 0.327628
R5315 VGND.n380 VGND.n376 0.327628
R5316 VGND.n383 VGND.n353 0.327628
R5317 VGND.n389 VGND.n388 0.327628
R5318 VGND.n2707 VGND.n2706 0.327628
R5319 VGND.n2727 VGND.n2725 0.327628
R5320 VGND.n2740 VGND.n2739 0.327628
R5321 VGND.n2736 VGND.n300 0.327628
R5322 VGND.n2733 VGND.n2732 0.327628
R5323 VGND.n2778 VGND.n2777 0.327628
R5324 VGND.n2774 VGND.n2772 0.327628
R5325 VGND.n2793 VGND.n2792 0.327628
R5326 VGND.n2789 VGND.n2785 0.327628
R5327 VGND.n2754 VGND.n288 0.327628
R5328 VGND.n2758 VGND.n2757 0.327628
R5329 VGND.n2749 VGND.n2745 0.327628
R5330 VGND.n2720 VGND.n2719 0.327628
R5331 VGND.n2716 VGND.n2712 0.327628
R5332 VGND.n2674 VGND.n2673 0.327628
R5333 VGND.n2670 VGND.n350 0.327628
R5334 VGND.n2665 VGND.n349 0.327628
R5335 VGND.n2660 VGND.n344 0.327628
R5336 VGND.n2655 VGND.n343 0.327628
R5337 VGND.n2650 VGND.n338 0.327628
R5338 VGND.n2645 VGND.n337 0.327628
R5339 VGND.n2640 VGND.n2636 0.327628
R5340 VGND.n2537 VGND.n283 0.327628
R5341 VGND.n2542 VGND.n282 0.327628
R5342 VGND.n2546 VGND.n2545 0.327628
R5343 VGND.n2289 VGND.n412 0.327628
R5344 VGND.n2294 VGND.n411 0.327628
R5345 VGND.n2299 VGND.n410 0.327628
R5346 VGND.n2304 VGND.n409 0.327628
R5347 VGND.n2309 VGND.n408 0.327628
R5348 VGND.n2314 VGND.n407 0.327628
R5349 VGND.n2319 VGND.n406 0.327628
R5350 VGND.n2324 VGND.n405 0.327628
R5351 VGND.n2329 VGND.n404 0.327628
R5352 VGND.n2334 VGND.n403 0.327628
R5353 VGND.n2339 VGND.n402 0.327628
R5354 VGND.n2344 VGND.n401 0.327628
R5355 VGND.n2526 VGND.n420 0.327628
R5356 VGND.n2523 VGND.n280 0.327628
R5357 VGND.n2518 VGND.n279 0.327628
R5358 VGND.n2513 VGND.n2509 0.327628
R5359 VGND.n2486 VGND.n2485 0.327628
R5360 VGND.n2482 VGND.n2478 0.327628
R5361 VGND.n2460 VGND.n2459 0.327628
R5362 VGND.n2456 VGND.n2452 0.327628
R5363 VGND.n2434 VGND.n2433 0.327628
R5364 VGND.n2430 VGND.n2426 0.327628
R5365 VGND.n2408 VGND.n2407 0.327628
R5366 VGND.n2404 VGND.n2400 0.327628
R5367 VGND.n2382 VGND.n2381 0.327628
R5368 VGND.n2378 VGND.n2374 0.327628
R5369 VGND.n2356 VGND.n2355 0.327628
R5370 VGND.n2814 VGND.n273 0.327628
R5371 VGND.n2811 VGND.n2807 0.327628
R5372 VGND.n2500 VGND.n277 0.327628
R5373 VGND.n2504 VGND.n2503 0.327628
R5374 VGND.n2495 VGND.n2491 0.327628
R5375 VGND.n2473 VGND.n2472 0.327628
R5376 VGND.n2469 VGND.n2465 0.327628
R5377 VGND.n2447 VGND.n2446 0.327628
R5378 VGND.n2443 VGND.n2439 0.327628
R5379 VGND.n2421 VGND.n2420 0.327628
R5380 VGND.n2417 VGND.n2413 0.327628
R5381 VGND.n2395 VGND.n2394 0.327628
R5382 VGND.n2391 VGND.n2387 0.327628
R5383 VGND.n2369 VGND.n2368 0.327628
R5384 VGND.n2365 VGND.n2361 0.327628
R5385 VGND.n1986 VGND.n271 0.327628
R5386 VGND.n1983 VGND.n270 0.327628
R5387 VGND.n1978 VGND.n1974 0.327628
R5388 VGND.n1971 VGND.n1970 0.327628
R5389 VGND.n1967 VGND.n1963 0.327628
R5390 VGND.n1960 VGND.n1959 0.327628
R5391 VGND.n1956 VGND.n1952 0.327628
R5392 VGND.n1949 VGND.n1948 0.327628
R5393 VGND.n1945 VGND.n1941 0.327628
R5394 VGND.n1938 VGND.n1937 0.327628
R5395 VGND.n1934 VGND.n1930 0.327628
R5396 VGND.n1927 VGND.n1926 0.327628
R5397 VGND.n1923 VGND.n1919 0.327628
R5398 VGND.n1916 VGND.n1915 0.327628
R5399 VGND.n1912 VGND.n1908 0.327628
R5400 VGND.n1999 VGND.n602 0.327628
R5401 VGND.n2002 VGND.n268 0.327628
R5402 VGND.n2007 VGND.n267 0.327628
R5403 VGND.n2012 VGND.n581 0.327628
R5404 VGND.n2017 VGND.n580 0.327628
R5405 VGND.n2022 VGND.n575 0.327628
R5406 VGND.n2027 VGND.n574 0.327628
R5407 VGND.n2032 VGND.n569 0.327628
R5408 VGND.n2037 VGND.n568 0.327628
R5409 VGND.n2042 VGND.n563 0.327628
R5410 VGND.n2047 VGND.n562 0.327628
R5411 VGND.n2052 VGND.n557 0.327628
R5412 VGND.n2057 VGND.n556 0.327628
R5413 VGND.n2061 VGND.n2060 0.327628
R5414 VGND.n598 VGND.n591 0.327628
R5415 VGND.n2839 VGND.n261 0.327628
R5416 VGND.n2836 VGND.n2832 0.327628
R5417 VGND.n2126 VGND.n265 0.327628
R5418 VGND.n2130 VGND.n2129 0.327628
R5419 VGND.n2121 VGND.n578 0.327628
R5420 VGND.n2116 VGND.n577 0.327628
R5421 VGND.n2111 VGND.n572 0.327628
R5422 VGND.n2106 VGND.n571 0.327628
R5423 VGND.n2101 VGND.n566 0.327628
R5424 VGND.n2096 VGND.n565 0.327628
R5425 VGND.n2091 VGND.n560 0.327628
R5426 VGND.n2086 VGND.n559 0.327628
R5427 VGND.n2081 VGND.n554 0.327628
R5428 VGND.n2076 VGND.n553 0.327628
R5429 VGND.n2071 VGND.n2067 0.327628
R5430 VGND.n1826 VGND.n259 0.327628
R5431 VGND.n1823 VGND.n258 0.327628
R5432 VGND.n1818 VGND.n1814 0.327628
R5433 VGND.n1811 VGND.n1810 0.327628
R5434 VGND.n1807 VGND.n1803 0.327628
R5435 VGND.n1800 VGND.n1799 0.327628
R5436 VGND.n1796 VGND.n1792 0.327628
R5437 VGND.n1789 VGND.n1788 0.327628
R5438 VGND.n1785 VGND.n1781 0.327628
R5439 VGND.n1778 VGND.n1777 0.327628
R5440 VGND.n1774 VGND.n1770 0.327628
R5441 VGND.n1767 VGND.n1766 0.327628
R5442 VGND.n1763 VGND.n1759 0.327628
R5443 VGND.n2175 VGND.n550 0.327628
R5444 VGND.n2178 VGND.n548 0.327628
R5445 VGND.n1839 VGND.n1735 0.327628
R5446 VGND.n1842 VGND.n256 0.327628
R5447 VGND.n1847 VGND.n255 0.327628
R5448 VGND.n1851 VGND.n1850 0.327628
R5449 VGND.n1731 VGND.n662 0.327628
R5450 VGND.n1726 VGND.n661 0.327628
R5451 VGND.n1721 VGND.n656 0.327628
R5452 VGND.n1716 VGND.n655 0.327628
R5453 VGND.n1711 VGND.n650 0.327628
R5454 VGND.n1706 VGND.n649 0.327628
R5455 VGND.n1701 VGND.n644 0.327628
R5456 VGND.n1696 VGND.n643 0.327628
R5457 VGND.n1691 VGND.n1687 0.327628
R5458 VGND.n1684 VGND.n1683 0.327628
R5459 VGND.n1680 VGND.n629 0.327628
R5460 VGND.n2864 VGND.n249 0.327628
R5461 VGND.n2861 VGND.n2857 0.327628
R5462 VGND.n726 VGND.n253 0.327628
R5463 VGND.n730 VGND.n729 0.327628
R5464 VGND.n721 VGND.n664 0.327628
R5465 VGND.n716 VGND.n659 0.327628
R5466 VGND.n711 VGND.n658 0.327628
R5467 VGND.n706 VGND.n653 0.327628
R5468 VGND.n701 VGND.n652 0.327628
R5469 VGND.n696 VGND.n647 0.327628
R5470 VGND.n691 VGND.n646 0.327628
R5471 VGND.n686 VGND.n641 0.327628
R5472 VGND.n681 VGND.n640 0.327628
R5473 VGND.n676 VGND.n634 0.327628
R5474 VGND.n671 VGND.n633 0.327628
R5475 VGND.n1658 VGND.n247 0.327628
R5476 VGND.n1663 VGND.n246 0.327628
R5477 VGND.n1667 VGND.n1666 0.327628
R5478 VGND.n855 VGND.n732 0.327628
R5479 VGND.n859 VGND.n858 0.327628
R5480 VGND.n850 VGND.n817 0.327628
R5481 VGND.n845 VGND.n816 0.327628
R5482 VGND.n840 VGND.n815 0.327628
R5483 VGND.n835 VGND.n814 0.327628
R5484 VGND.n830 VGND.n813 0.327628
R5485 VGND.n825 VGND.n812 0.327628
R5486 VGND.n868 VGND.n808 0.327628
R5487 VGND.n871 VGND.n637 0.327628
R5488 VGND.n876 VGND.n636 0.327628
R5489 VGND.n1354 VGND.n1350 0.327628
R5490 VGND.n1647 VGND.n741 0.327628
R5491 VGND.n1644 VGND.n244 0.327628
R5492 VGND.n1639 VGND.n243 0.327628
R5493 VGND.n1634 VGND.n1630 0.327628
R5494 VGND.n1554 VGND.n742 0.327628
R5495 VGND.n1558 VGND.n1557 0.327628
R5496 VGND.n1549 VGND.n758 0.327628
R5497 VGND.n1544 VGND.n1540 0.327628
R5498 VGND.n1522 VGND.n1521 0.327628
R5499 VGND.n1518 VGND.n1514 0.327628
R5500 VGND.n1496 VGND.n1495 0.327628
R5501 VGND.n1492 VGND.n1488 0.327628
R5502 VGND.n1401 VGND.n1400 0.327628
R5503 VGND.n1397 VGND.n802 0.327628
R5504 VGND.n1392 VGND.n801 0.327628
R5505 VGND.n2889 VGND.n236 0.327628
R5506 VGND.n2886 VGND.n2882 0.327628
R5507 VGND.n1573 VGND.n240 0.327628
R5508 VGND.n1578 VGND.n745 0.327628
R5509 VGND.n1583 VGND.n744 0.327628
R5510 VGND.n1587 VGND.n1586 0.327628
R5511 VGND.n1568 VGND.n1564 0.327628
R5512 VGND.n1535 VGND.n1534 0.327628
R5513 VGND.n1531 VGND.n1527 0.327628
R5514 VGND.n1509 VGND.n1508 0.327628
R5515 VGND.n1505 VGND.n1501 0.327628
R5516 VGND.n1483 VGND.n1482 0.327628
R5517 VGND.n1479 VGND.n1475 0.327628
R5518 VGND.n1416 VGND.n1415 0.327628
R5519 VGND.n1412 VGND.n1408 0.327628
R5520 VGND.n1610 VGND.n232 0.327628
R5521 VGND.n1615 VGND.n231 0.327628
R5522 VGND.n1619 VGND.n1618 0.327628
R5523 VGND.n1602 VGND.n747 0.327628
R5524 VGND.n1597 VGND.n1593 0.327628
R5525 VGND.n1460 VGND.n751 0.327628
R5526 VGND.n1464 VGND.n1463 0.327628
R5527 VGND.n1455 VGND.n788 0.327628
R5528 VGND.n1450 VGND.n787 0.327628
R5529 VGND.n1445 VGND.n786 0.327628
R5530 VGND.n1440 VGND.n785 0.327628
R5531 VGND.n1435 VGND.n784 0.327628
R5532 VGND.n1430 VGND.n783 0.327628
R5533 VGND.n1425 VGND.n1421 0.327628
R5534 VGND.n1343 VGND.n1342 0.327628
R5535 VGND.n2909 VGND.n228 0.327628
R5536 VGND.n2906 VGND.n2902 0.327628
R5537 VGND.n1063 VGND.n1062 0.327628
R5538 VGND.n1059 VGND.n1046 0.327628
R5539 VGND.n1054 VGND.n1045 0.327628
R5540 VGND.n1068 VGND.n1041 0.327628
R5541 VGND.n1071 VGND.n912 0.327628
R5542 VGND.n1076 VGND.n911 0.327628
R5543 VGND.n1081 VGND.n906 0.327628
R5544 VGND.n1086 VGND.n905 0.327628
R5545 VGND.n1091 VGND.n900 0.327628
R5546 VGND.n1096 VGND.n899 0.327628
R5547 VGND.n1100 VGND.n1099 0.327628
R5548 VGND.n1038 VGND.n1026 0.327628
R5549 VGND.n1033 VGND.n1025 0.327628
R5550 VGND.n1167 VGND.n1165 0.327628
R5551 VGND.n1174 VGND.n1170 0.327628
R5552 VGND.n1177 VGND.n1011 0.327628
R5553 VGND.n1187 VGND.n1183 0.327628
R5554 VGND.n1191 VGND.n1190 0.327628
R5555 VGND.n1206 VGND.n1202 0.327628
R5556 VGND.n1209 VGND.n1003 0.327628
R5557 VGND.n1219 VGND.n1215 0.327628
R5558 VGND.n1249 VGND.n1248 0.327628
R5559 VGND.n1245 VGND.n1223 0.327628
R5560 VGND.n1242 VGND.n1241 0.327628
R5561 VGND.n1238 VGND.n1228 0.327628
R5562 VGND.n1235 VGND.n1234 0.327628
R5563 VGND.n1276 VGND.n1272 0.327628
R5564 VGND.n1279 VGND.n997 0.327628
R5565 VGND.n992 VGND.n991 0.327628
R5566 VGND.n988 VGND.n925 0.327628
R5567 VGND.n983 VGND.n924 0.327628
R5568 VGND.n978 VGND.n920 0.327628
R5569 VGND.n973 VGND.n919 0.327628
R5570 VGND.n968 VGND.n915 0.327628
R5571 VGND.n963 VGND.n914 0.327628
R5572 VGND.n958 VGND.n909 0.327628
R5573 VGND.n953 VGND.n908 0.327628
R5574 VGND.n948 VGND.n903 0.327628
R5575 VGND.n943 VGND.n902 0.327628
R5576 VGND.n938 VGND.n897 0.327628
R5577 VGND.n933 VGND.n896 0.327628
R5578 VGND.n1331 VGND.n890 0.327628
R5579 VGND.n1334 VGND.n888 0.327628
R5580 VGND.n126 VGND.n125 0.213567
R5581 VGND.n125 VGND.n32 0.213567
R5582 VGND.n3002 VGND.n32 0.213567
R5583 VGND.n3002 VGND.n3001 0.213567
R5584 VGND.n1157 VGND.n1134 0.213567
R5585 VGND.n1134 VGND.n543 0.213567
R5586 VGND.n2219 VGND.n543 0.213567
R5587 VGND.n2219 VGND.n2218 0.213567
R5588 VGND.n2218 VGND.n0 0.213567
R5589 VGND.n3001 VGND.n33 0.2073
R5590 VGND.n3024 VGND.n2 0.18968
R5591 VGND.n1159 VGND.n1158 0.175967
R5592 VGND.n2633 VGND 0.169807
R5593 VGND.n2695 VGND 0.169807
R5594 VGND.n2690 VGND 0.169807
R5595 VGND.n2689 VGND 0.169807
R5596 VGND.n2684 VGND 0.169807
R5597 VGND.n2683 VGND 0.169807
R5598 VGND.n2678 VGND 0.169807
R5599 VGND.n2677 VGND 0.169807
R5600 VGND.n2709 VGND 0.169807
R5601 VGND.n2723 VGND 0.169807
R5602 VGND.n2742 VGND 0.169807
R5603 VGND.n2761 VGND 0.169807
R5604 VGND.n2781 VGND 0.169807
R5605 VGND.n2780 VGND 0.169807
R5606 VGND.n284 VGND 0.169807
R5607 VGND.n2635 VGND 0.169807
R5608 VGND.n2693 VGND 0.169807
R5609 VGND.n2692 VGND 0.169807
R5610 VGND.n2687 VGND 0.169807
R5611 VGND.n2686 VGND 0.169807
R5612 VGND.n2681 VGND 0.169807
R5613 VGND.n2680 VGND 0.169807
R5614 VGND.n2675 VGND 0.169807
R5615 VGND.n2711 VGND 0.169807
R5616 VGND.n2721 VGND 0.169807
R5617 VGND.n2744 VGND 0.169807
R5618 VGND.n2759 VGND 0.169807
R5619 VGND VGND.n2783 0.169807
R5620 VGND.n2784 VGND 0.169807
R5621 VGND.n2794 VGND 0.169807
R5622 VGND.n2559 VGND 0.169807
R5623 VGND.n2558 VGND 0.169807
R5624 VGND.n2557 VGND 0.169807
R5625 VGND.n2556 VGND 0.169807
R5626 VGND.n2555 VGND 0.169807
R5627 VGND.n2554 VGND 0.169807
R5628 VGND.n2553 VGND 0.169807
R5629 VGND.n2552 VGND 0.169807
R5630 VGND.n2551 VGND 0.169807
R5631 VGND.n2550 VGND 0.169807
R5632 VGND.n2549 VGND 0.169807
R5633 VGND.n2548 VGND 0.169807
R5634 VGND.n2547 VGND 0.169807
R5635 VGND.n2798 VGND 0.169807
R5636 VGND.n2797 VGND 0.169807
R5637 VGND.n2357 VGND 0.169807
R5638 VGND.n2373 VGND 0.169807
R5639 VGND.n2383 VGND 0.169807
R5640 VGND.n2399 VGND 0.169807
R5641 VGND.n2409 VGND 0.169807
R5642 VGND.n2425 VGND 0.169807
R5643 VGND.n2435 VGND 0.169807
R5644 VGND.n2451 VGND 0.169807
R5645 VGND.n2461 VGND 0.169807
R5646 VGND.n2477 VGND 0.169807
R5647 VGND.n2487 VGND 0.169807
R5648 VGND.n2508 VGND 0.169807
R5649 VGND.n2802 VGND 0.169807
R5650 VGND.n2801 VGND 0.169807
R5651 VGND.n419 VGND 0.169807
R5652 VGND.n2360 VGND 0.169807
R5653 VGND.n2370 VGND 0.169807
R5654 VGND.n2386 VGND 0.169807
R5655 VGND.n2396 VGND 0.169807
R5656 VGND.n2412 VGND 0.169807
R5657 VGND.n2422 VGND 0.169807
R5658 VGND.n2438 VGND 0.169807
R5659 VGND.n2448 VGND 0.169807
R5660 VGND.n2464 VGND 0.169807
R5661 VGND.n2474 VGND 0.169807
R5662 VGND.n2490 VGND 0.169807
R5663 VGND.n2505 VGND 0.169807
R5664 VGND VGND.n2805 0.169807
R5665 VGND.n2806 VGND 0.169807
R5666 VGND.n2819 VGND 0.169807
R5667 VGND.n1907 VGND 0.169807
R5668 VGND VGND.n1917 0.169807
R5669 VGND.n1918 VGND 0.169807
R5670 VGND VGND.n1928 0.169807
R5671 VGND.n1929 VGND 0.169807
R5672 VGND VGND.n1939 0.169807
R5673 VGND.n1940 VGND 0.169807
R5674 VGND VGND.n1950 0.169807
R5675 VGND.n1951 VGND 0.169807
R5676 VGND VGND.n1961 0.169807
R5677 VGND.n1962 VGND 0.169807
R5678 VGND VGND.n1972 0.169807
R5679 VGND.n1973 VGND 0.169807
R5680 VGND.n2823 VGND 0.169807
R5681 VGND.n2822 VGND 0.169807
R5682 VGND.n2063 VGND 0.169807
R5683 VGND.n2062 VGND 0.169807
R5684 VGND.n2167 VGND 0.169807
R5685 VGND.n2166 VGND 0.169807
R5686 VGND.n2159 VGND 0.169807
R5687 VGND.n2158 VGND 0.169807
R5688 VGND.n2151 VGND 0.169807
R5689 VGND.n2150 VGND 0.169807
R5690 VGND.n2143 VGND 0.169807
R5691 VGND.n2142 VGND 0.169807
R5692 VGND.n2135 VGND 0.169807
R5693 VGND.n2134 VGND 0.169807
R5694 VGND.n2827 VGND 0.169807
R5695 VGND.n2826 VGND 0.169807
R5696 VGND.n1998 VGND 0.169807
R5697 VGND.n2066 VGND 0.169807
R5698 VGND.n2171 VGND 0.169807
R5699 VGND.n2170 VGND 0.169807
R5700 VGND.n2163 VGND 0.169807
R5701 VGND.n2162 VGND 0.169807
R5702 VGND.n2155 VGND 0.169807
R5703 VGND.n2154 VGND 0.169807
R5704 VGND.n2147 VGND 0.169807
R5705 VGND.n2146 VGND 0.169807
R5706 VGND.n2139 VGND 0.169807
R5707 VGND.n2138 VGND 0.169807
R5708 VGND.n2131 VGND 0.169807
R5709 VGND VGND.n2830 0.169807
R5710 VGND.n2831 VGND 0.169807
R5711 VGND.n2844 VGND 0.169807
R5712 VGND.n1901 VGND 0.169807
R5713 VGND.n2174 VGND 0.169807
R5714 VGND.n1758 VGND 0.169807
R5715 VGND VGND.n1768 0.169807
R5716 VGND.n1769 VGND 0.169807
R5717 VGND VGND.n1779 0.169807
R5718 VGND.n1780 VGND 0.169807
R5719 VGND VGND.n1790 0.169807
R5720 VGND.n1791 VGND 0.169807
R5721 VGND VGND.n1801 0.169807
R5722 VGND.n1802 VGND 0.169807
R5723 VGND VGND.n1812 0.169807
R5724 VGND.n1813 VGND 0.169807
R5725 VGND.n2848 VGND 0.169807
R5726 VGND.n2847 VGND 0.169807
R5727 VGND.n1899 VGND 0.169807
R5728 VGND VGND.n1685 0.169807
R5729 VGND.n1686 VGND 0.169807
R5730 VGND.n1884 VGND 0.169807
R5731 VGND.n1883 VGND 0.169807
R5732 VGND.n1876 VGND 0.169807
R5733 VGND.n1875 VGND 0.169807
R5734 VGND.n1868 VGND 0.169807
R5735 VGND.n1867 VGND 0.169807
R5736 VGND.n1860 VGND 0.169807
R5737 VGND.n1859 VGND 0.169807
R5738 VGND.n1852 VGND 0.169807
R5739 VGND.n2852 VGND 0.169807
R5740 VGND.n2851 VGND 0.169807
R5741 VGND.n1838 VGND 0.169807
R5742 VGND.n1896 VGND 0.169807
R5743 VGND.n1895 VGND 0.169807
R5744 VGND.n1888 VGND 0.169807
R5745 VGND.n1887 VGND 0.169807
R5746 VGND.n1880 VGND 0.169807
R5747 VGND.n1879 VGND 0.169807
R5748 VGND.n1872 VGND 0.169807
R5749 VGND.n1871 VGND 0.169807
R5750 VGND.n1864 VGND 0.169807
R5751 VGND.n1863 VGND 0.169807
R5752 VGND.n1856 VGND 0.169807
R5753 VGND.n1855 VGND 0.169807
R5754 VGND VGND.n2855 0.169807
R5755 VGND.n2856 VGND 0.169807
R5756 VGND.n2869 VGND 0.169807
R5757 VGND.n1349 VGND 0.169807
R5758 VGND.n1892 VGND 0.169807
R5759 VGND.n1891 VGND 0.169807
R5760 VGND.n867 VGND 0.169807
R5761 VGND.n866 VGND 0.169807
R5762 VGND.n865 VGND 0.169807
R5763 VGND.n864 VGND 0.169807
R5764 VGND.n863 VGND 0.169807
R5765 VGND.n862 VGND 0.169807
R5766 VGND.n861 VGND 0.169807
R5767 VGND.n860 VGND 0.169807
R5768 VGND.n1669 VGND 0.169807
R5769 VGND.n1668 VGND 0.169807
R5770 VGND.n2873 VGND 0.169807
R5771 VGND.n2872 VGND 0.169807
R5772 VGND.n1404 VGND 0.169807
R5773 VGND.n1403 VGND 0.169807
R5774 VGND.n1402 VGND 0.169807
R5775 VGND.n1487 VGND 0.169807
R5776 VGND.n1497 VGND 0.169807
R5777 VGND.n1513 VGND 0.169807
R5778 VGND.n1523 VGND 0.169807
R5779 VGND.n1539 VGND 0.169807
R5780 VGND.n1560 VGND 0.169807
R5781 VGND.n1559 VGND 0.169807
R5782 VGND VGND.n1628 0.169807
R5783 VGND.n1629 VGND 0.169807
R5784 VGND.n2877 VGND 0.169807
R5785 VGND.n2876 VGND 0.169807
R5786 VGND.n740 VGND 0.169807
R5787 VGND.n1407 VGND 0.169807
R5788 VGND.n1417 VGND 0.169807
R5789 VGND.n1474 VGND 0.169807
R5790 VGND.n1484 VGND 0.169807
R5791 VGND.n1500 VGND 0.169807
R5792 VGND.n1510 VGND 0.169807
R5793 VGND.n1526 VGND 0.169807
R5794 VGND.n1536 VGND 0.169807
R5795 VGND.n1563 VGND 0.169807
R5796 VGND.n1588 VGND 0.169807
R5797 VGND.n1625 VGND 0.169807
R5798 VGND.n1624 VGND 0.169807
R5799 VGND VGND.n2880 0.169807
R5800 VGND.n2881 VGND 0.169807
R5801 VGND.n2894 VGND 0.169807
R5802 VGND.n1344 VGND 0.169807
R5803 VGND.n1420 VGND 0.169807
R5804 VGND.n1471 VGND 0.169807
R5805 VGND.n1470 VGND 0.169807
R5806 VGND.n1469 VGND 0.169807
R5807 VGND.n1468 VGND 0.169807
R5808 VGND.n1467 VGND 0.169807
R5809 VGND.n1466 VGND 0.169807
R5810 VGND.n1465 VGND 0.169807
R5811 VGND VGND.n1591 0.169807
R5812 VGND.n1592 VGND 0.169807
R5813 VGND.n1621 VGND 0.169807
R5814 VGND.n1620 VGND 0.169807
R5815 VGND.n2898 VGND 0.169807
R5816 VGND.n2897 VGND 0.169807
R5817 VGND.n1103 VGND 0.169807
R5818 VGND.n1102 VGND 0.169807
R5819 VGND.n1101 VGND 0.169807
R5820 VGND.n1321 VGND 0.169807
R5821 VGND.n1320 VGND 0.169807
R5822 VGND.n1313 VGND 0.169807
R5823 VGND.n1312 VGND 0.169807
R5824 VGND.n1305 VGND 0.169807
R5825 VGND.n1304 VGND 0.169807
R5826 VGND.n1067 VGND 0.169807
R5827 VGND.n1066 VGND 0.169807
R5828 VGND.n1065 VGND 0.169807
R5829 VGND.n1064 VGND 0.169807
R5830 VGND.n2901 VGND 0.169807
R5831 VGND.n233 VGND 0.169807
R5832 VGND.n1163 VGND 0.169807
R5833 VGND.n1328 VGND 0.169807
R5834 VGND.n1327 VGND 0.169807
R5835 VGND VGND.n898 0.169807
R5836 VGND VGND.n901 0.169807
R5837 VGND VGND.n904 0.169807
R5838 VGND VGND.n907 0.169807
R5839 VGND VGND.n910 0.169807
R5840 VGND VGND.n913 0.169807
R5841 VGND.n1298 VGND 0.169807
R5842 VGND.n1297 VGND 0.169807
R5843 VGND.n1292 VGND 0.169807
R5844 VGND.n1291 VGND 0.169807
R5845 VGND.n1270 VGND 0.169807
R5846 VGND.n1285 VGND 0.169807
R5847 VGND.n1161 VGND 0.169807
R5848 VGND.n1330 VGND 0.169807
R5849 VGND.n1325 VGND 0.169807
R5850 VGND.n1324 VGND 0.169807
R5851 VGND.n1317 VGND 0.169807
R5852 VGND.n1316 VGND 0.169807
R5853 VGND.n1309 VGND 0.169807
R5854 VGND.n1308 VGND 0.169807
R5855 VGND.n1301 VGND 0.169807
R5856 VGND.n1300 VGND 0.169807
R5857 VGND.n1295 VGND 0.169807
R5858 VGND.n1294 VGND 0.169807
R5859 VGND.n1289 VGND 0.169807
R5860 VGND.n1288 VGND 0.169807
R5861 VGND.n1287 VGND 0.169807
R5862 VGND.n190 VGND 0.159538
R5863 VGND.n161 VGND 0.159538
R5864 VGND.n2915 VGND.n224 0.154425
R5865 VGND.n2915 VGND.n2914 0.154425
R5866 VGND.n2914 VGND.n225 0.154425
R5867 VGND.n238 VGND.n225 0.154425
R5868 VGND.n1652 VGND.n238 0.154425
R5869 VGND.n1653 VGND.n1652 0.154425
R5870 VGND.n1653 VGND.n251 0.154425
R5871 VGND.n1832 VGND.n251 0.154425
R5872 VGND.n1832 VGND.n1831 0.154425
R5873 VGND.n1831 VGND.n263 0.154425
R5874 VGND.n1992 VGND.n263 0.154425
R5875 VGND.n1992 VGND.n1991 0.154425
R5876 VGND.n1991 VGND.n275 0.154425
R5877 VGND.n417 VGND.n275 0.154425
R5878 VGND.n417 VGND.n207 0.154425
R5879 VGND.n2938 VGND.n207 0.154425
R5880 VGND.n2939 VGND.n2938 0.154425
R5881 VGND.n1160 VGND.n1159 0.154425
R5882 VGND.n1160 VGND.n880 0.154425
R5883 VGND.n1345 VGND.n880 0.154425
R5884 VGND.n1346 VGND.n1345 0.154425
R5885 VGND.n1347 VGND.n1346 0.154425
R5886 VGND.n1348 VGND.n1347 0.154425
R5887 VGND.n1348 VGND.n626 0.154425
R5888 VGND.n1900 VGND.n626 0.154425
R5889 VGND.n1902 VGND.n1900 0.154425
R5890 VGND.n1903 VGND.n1902 0.154425
R5891 VGND.n1904 VGND.n1903 0.154425
R5892 VGND.n1906 VGND.n1904 0.154425
R5893 VGND.n1906 VGND.n1905 0.154425
R5894 VGND.n1905 VGND.n398 0.154425
R5895 VGND.n2560 VGND.n398 0.154425
R5896 VGND.n2561 VGND.n2560 0.154425
R5897 VGND.n2562 VGND.n2561 0.154425
R5898 VGND.n1144 VGND.n1138 0.144904
R5899 VGND.n1117 VGND.n1109 0.144904
R5900 VGND.n2232 VGND.n2228 0.144904
R5901 VGND.n1370 VGND.n1366 0.144904
R5902 VGND.n2632 VGND.n2608 0.138284
R5903 VGND.n2700 VGND.n2699 0.13638
R5904 VGND.n355 VGND.n333 0.13638
R5905 VGND.n362 VGND.n361 0.13638
R5906 VGND.n369 VGND.n368 0.13638
R5907 VGND.n373 VGND.n372 0.13638
R5908 VGND.n380 VGND.n379 0.13638
R5909 VGND.n384 VGND.n383 0.13638
R5910 VGND.n388 VGND.n387 0.13638
R5911 VGND.n2706 VGND.n326 0.13638
R5912 VGND.n2727 VGND.n2726 0.13638
R5913 VGND.n2739 VGND.n312 0.13638
R5914 VGND.n2736 VGND.n2735 0.13638
R5915 VGND.n2732 VGND.n2730 0.13638
R5916 VGND.n2777 VGND.n294 0.13638
R5917 VGND.n2774 VGND.n2773 0.13638
R5918 VGND.n2792 VGND.n287 0.13638
R5919 VGND.n2789 VGND.n2788 0.13638
R5920 VGND.n2754 VGND.n2753 0.13638
R5921 VGND.n2757 VGND.n304 0.13638
R5922 VGND.n2749 VGND.n2748 0.13638
R5923 VGND.n2719 VGND.n320 0.13638
R5924 VGND.n2716 VGND.n2715 0.13638
R5925 VGND.n2673 VGND.n394 0.13638
R5926 VGND.n2670 VGND.n2669 0.13638
R5927 VGND.n2665 VGND.n2664 0.13638
R5928 VGND.n2660 VGND.n2659 0.13638
R5929 VGND.n2655 VGND.n2654 0.13638
R5930 VGND.n2650 VGND.n2649 0.13638
R5931 VGND.n2645 VGND.n2644 0.13638
R5932 VGND.n2640 VGND.n2639 0.13638
R5933 VGND.n2537 VGND.n2536 0.13638
R5934 VGND.n2542 VGND.n2541 0.13638
R5935 VGND.n2545 VGND.n415 0.13638
R5936 VGND.n2289 VGND.n2288 0.13638
R5937 VGND.n2294 VGND.n2293 0.13638
R5938 VGND.n2299 VGND.n2298 0.13638
R5939 VGND.n2304 VGND.n2303 0.13638
R5940 VGND.n2309 VGND.n2308 0.13638
R5941 VGND.n2314 VGND.n2313 0.13638
R5942 VGND.n2319 VGND.n2318 0.13638
R5943 VGND.n2324 VGND.n2323 0.13638
R5944 VGND.n2329 VGND.n2328 0.13638
R5945 VGND.n2334 VGND.n2333 0.13638
R5946 VGND.n2339 VGND.n2338 0.13638
R5947 VGND.n2344 VGND.n2343 0.13638
R5948 VGND.n2527 VGND.n2526 0.13638
R5949 VGND.n2523 VGND.n2522 0.13638
R5950 VGND.n2518 VGND.n2517 0.13638
R5951 VGND.n2513 VGND.n2512 0.13638
R5952 VGND.n2485 VGND.n428 0.13638
R5953 VGND.n2482 VGND.n2481 0.13638
R5954 VGND.n2459 VGND.n436 0.13638
R5955 VGND.n2456 VGND.n2455 0.13638
R5956 VGND.n2433 VGND.n444 0.13638
R5957 VGND.n2430 VGND.n2429 0.13638
R5958 VGND.n2407 VGND.n452 0.13638
R5959 VGND.n2404 VGND.n2403 0.13638
R5960 VGND.n2381 VGND.n460 0.13638
R5961 VGND.n2378 VGND.n2377 0.13638
R5962 VGND.n2355 VGND.n472 0.13638
R5963 VGND.n2815 VGND.n2814 0.13638
R5964 VGND.n2811 VGND.n2810 0.13638
R5965 VGND.n2500 VGND.n2499 0.13638
R5966 VGND.n2503 VGND.n424 0.13638
R5967 VGND.n2495 VGND.n2494 0.13638
R5968 VGND.n2472 VGND.n432 0.13638
R5969 VGND.n2469 VGND.n2468 0.13638
R5970 VGND.n2446 VGND.n440 0.13638
R5971 VGND.n2443 VGND.n2442 0.13638
R5972 VGND.n2420 VGND.n448 0.13638
R5973 VGND.n2417 VGND.n2416 0.13638
R5974 VGND.n2394 VGND.n456 0.13638
R5975 VGND.n2391 VGND.n2390 0.13638
R5976 VGND.n2368 VGND.n464 0.13638
R5977 VGND.n2365 VGND.n2364 0.13638
R5978 VGND.n1987 VGND.n1986 0.13638
R5979 VGND.n1983 VGND.n1982 0.13638
R5980 VGND.n1978 VGND.n1977 0.13638
R5981 VGND.n1970 VGND.n608 0.13638
R5982 VGND.n1967 VGND.n1966 0.13638
R5983 VGND.n1959 VGND.n611 0.13638
R5984 VGND.n1956 VGND.n1955 0.13638
R5985 VGND.n1948 VGND.n614 0.13638
R5986 VGND.n1945 VGND.n1944 0.13638
R5987 VGND.n1937 VGND.n617 0.13638
R5988 VGND.n1934 VGND.n1933 0.13638
R5989 VGND.n1926 VGND.n620 0.13638
R5990 VGND.n1923 VGND.n1922 0.13638
R5991 VGND.n1915 VGND.n623 0.13638
R5992 VGND.n1912 VGND.n1911 0.13638
R5993 VGND.n1994 VGND.n602 0.13638
R5994 VGND.n2002 VGND.n2001 0.13638
R5995 VGND.n2007 VGND.n2006 0.13638
R5996 VGND.n2012 VGND.n2011 0.13638
R5997 VGND.n2017 VGND.n2016 0.13638
R5998 VGND.n2022 VGND.n2021 0.13638
R5999 VGND.n2027 VGND.n2026 0.13638
R6000 VGND.n2032 VGND.n2031 0.13638
R6001 VGND.n2037 VGND.n2036 0.13638
R6002 VGND.n2042 VGND.n2041 0.13638
R6003 VGND.n2047 VGND.n2046 0.13638
R6004 VGND.n2052 VGND.n2051 0.13638
R6005 VGND.n2057 VGND.n2056 0.13638
R6006 VGND.n2060 VGND.n594 0.13638
R6007 VGND.n598 VGND.n597 0.13638
R6008 VGND.n2840 VGND.n2839 0.13638
R6009 VGND.n2836 VGND.n2835 0.13638
R6010 VGND.n2126 VGND.n2125 0.13638
R6011 VGND.n2129 VGND.n585 0.13638
R6012 VGND.n2121 VGND.n2120 0.13638
R6013 VGND.n2116 VGND.n2115 0.13638
R6014 VGND.n2111 VGND.n2110 0.13638
R6015 VGND.n2106 VGND.n2105 0.13638
R6016 VGND.n2101 VGND.n2100 0.13638
R6017 VGND.n2096 VGND.n2095 0.13638
R6018 VGND.n2091 VGND.n2090 0.13638
R6019 VGND.n2086 VGND.n2085 0.13638
R6020 VGND.n2081 VGND.n2080 0.13638
R6021 VGND.n2076 VGND.n2075 0.13638
R6022 VGND.n2071 VGND.n2070 0.13638
R6023 VGND.n1827 VGND.n1826 0.13638
R6024 VGND.n1823 VGND.n1822 0.13638
R6025 VGND.n1818 VGND.n1817 0.13638
R6026 VGND.n1810 VGND.n1741 0.13638
R6027 VGND.n1807 VGND.n1806 0.13638
R6028 VGND.n1799 VGND.n1744 0.13638
R6029 VGND.n1796 VGND.n1795 0.13638
R6030 VGND.n1788 VGND.n1747 0.13638
R6031 VGND.n1785 VGND.n1784 0.13638
R6032 VGND.n1777 VGND.n1750 0.13638
R6033 VGND.n1774 VGND.n1773 0.13638
R6034 VGND.n1766 VGND.n1753 0.13638
R6035 VGND.n1763 VGND.n1762 0.13638
R6036 VGND.n1756 VGND.n550 0.13638
R6037 VGND.n2178 VGND.n2177 0.13638
R6038 VGND.n1834 VGND.n1735 0.13638
R6039 VGND.n1842 VGND.n1841 0.13638
R6040 VGND.n1847 VGND.n1846 0.13638
R6041 VGND.n1850 VGND.n1673 0.13638
R6042 VGND.n1731 VGND.n1730 0.13638
R6043 VGND.n1726 VGND.n1725 0.13638
R6044 VGND.n1721 VGND.n1720 0.13638
R6045 VGND.n1716 VGND.n1715 0.13638
R6046 VGND.n1711 VGND.n1710 0.13638
R6047 VGND.n1706 VGND.n1705 0.13638
R6048 VGND.n1701 VGND.n1700 0.13638
R6049 VGND.n1696 VGND.n1695 0.13638
R6050 VGND.n1691 VGND.n1690 0.13638
R6051 VGND.n1683 VGND.n1676 0.13638
R6052 VGND.n1680 VGND.n1679 0.13638
R6053 VGND.n2865 VGND.n2864 0.13638
R6054 VGND.n2861 VGND.n2860 0.13638
R6055 VGND.n726 VGND.n725 0.13638
R6056 VGND.n729 VGND.n667 0.13638
R6057 VGND.n721 VGND.n720 0.13638
R6058 VGND.n716 VGND.n715 0.13638
R6059 VGND.n711 VGND.n710 0.13638
R6060 VGND.n706 VGND.n705 0.13638
R6061 VGND.n701 VGND.n700 0.13638
R6062 VGND.n696 VGND.n695 0.13638
R6063 VGND.n691 VGND.n690 0.13638
R6064 VGND.n686 VGND.n685 0.13638
R6065 VGND.n681 VGND.n680 0.13638
R6066 VGND.n676 VGND.n675 0.13638
R6067 VGND.n671 VGND.n670 0.13638
R6068 VGND.n1658 VGND.n1657 0.13638
R6069 VGND.n1663 VGND.n1662 0.13638
R6070 VGND.n1666 VGND.n735 0.13638
R6071 VGND.n855 VGND.n854 0.13638
R6072 VGND.n858 VGND.n820 0.13638
R6073 VGND.n850 VGND.n849 0.13638
R6074 VGND.n845 VGND.n844 0.13638
R6075 VGND.n840 VGND.n839 0.13638
R6076 VGND.n835 VGND.n834 0.13638
R6077 VGND.n830 VGND.n829 0.13638
R6078 VGND.n825 VGND.n824 0.13638
R6079 VGND.n810 VGND.n808 0.13638
R6080 VGND.n871 VGND.n870 0.13638
R6081 VGND.n876 VGND.n875 0.13638
R6082 VGND.n1354 VGND.n1353 0.13638
R6083 VGND.n1648 VGND.n1647 0.13638
R6084 VGND.n1644 VGND.n1643 0.13638
R6085 VGND.n1639 VGND.n1638 0.13638
R6086 VGND.n1634 VGND.n1633 0.13638
R6087 VGND.n1554 VGND.n1553 0.13638
R6088 VGND.n1557 VGND.n761 0.13638
R6089 VGND.n1549 VGND.n1548 0.13638
R6090 VGND.n1544 VGND.n1543 0.13638
R6091 VGND.n1521 VGND.n769 0.13638
R6092 VGND.n1518 VGND.n1517 0.13638
R6093 VGND.n1495 VGND.n777 0.13638
R6094 VGND.n1492 VGND.n1491 0.13638
R6095 VGND.n1400 VGND.n805 0.13638
R6096 VGND.n1397 VGND.n1396 0.13638
R6097 VGND.n1392 VGND.n1391 0.13638
R6098 VGND.n2890 VGND.n2889 0.13638
R6099 VGND.n2886 VGND.n2885 0.13638
R6100 VGND.n1573 VGND.n1572 0.13638
R6101 VGND.n1578 VGND.n1577 0.13638
R6102 VGND.n1583 VGND.n1582 0.13638
R6103 VGND.n1586 VGND.n756 0.13638
R6104 VGND.n1568 VGND.n1567 0.13638
R6105 VGND.n1534 VGND.n765 0.13638
R6106 VGND.n1531 VGND.n1530 0.13638
R6107 VGND.n1508 VGND.n773 0.13638
R6108 VGND.n1505 VGND.n1504 0.13638
R6109 VGND.n1482 VGND.n781 0.13638
R6110 VGND.n1479 VGND.n1478 0.13638
R6111 VGND.n1415 VGND.n795 0.13638
R6112 VGND.n1412 VGND.n1411 0.13638
R6113 VGND.n1610 VGND.n1609 0.13638
R6114 VGND.n1615 VGND.n1614 0.13638
R6115 VGND.n1618 VGND.n750 0.13638
R6116 VGND.n1602 VGND.n1601 0.13638
R6117 VGND.n1597 VGND.n1596 0.13638
R6118 VGND.n1460 VGND.n1459 0.13638
R6119 VGND.n1463 VGND.n791 0.13638
R6120 VGND.n1455 VGND.n1454 0.13638
R6121 VGND.n1450 VGND.n1449 0.13638
R6122 VGND.n1445 VGND.n1444 0.13638
R6123 VGND.n1440 VGND.n1439 0.13638
R6124 VGND.n1435 VGND.n1434 0.13638
R6125 VGND.n1430 VGND.n1429 0.13638
R6126 VGND.n1425 VGND.n1424 0.13638
R6127 VGND.n1342 VGND.n885 0.13638
R6128 VGND.n2910 VGND.n2909 0.13638
R6129 VGND.n2906 VGND.n2905 0.13638
R6130 VGND.n1062 VGND.n1049 0.13638
R6131 VGND.n1059 VGND.n1058 0.13638
R6132 VGND.n1054 VGND.n1053 0.13638
R6133 VGND.n1043 VGND.n1041 0.13638
R6134 VGND.n1071 VGND.n1070 0.13638
R6135 VGND.n1076 VGND.n1075 0.13638
R6136 VGND.n1081 VGND.n1080 0.13638
R6137 VGND.n1086 VGND.n1085 0.13638
R6138 VGND.n1091 VGND.n1090 0.13638
R6139 VGND.n1096 VGND.n1095 0.13638
R6140 VGND.n1099 VGND.n1029 0.13638
R6141 VGND.n1038 VGND.n1037 0.13638
R6142 VGND.n1033 VGND.n1032 0.13638
R6143 VGND.n1168 VGND.n1167 0.13638
R6144 VGND.n1174 VGND.n1173 0.13638
R6145 VGND.n1178 VGND.n1177 0.13638
R6146 VGND.n1187 VGND.n1186 0.13638
R6147 VGND.n1190 VGND.n1009 0.13638
R6148 VGND.n1206 VGND.n1205 0.13638
R6149 VGND.n1210 VGND.n1209 0.13638
R6150 VGND.n1219 VGND.n1218 0.13638
R6151 VGND.n1248 VGND.n1001 0.13638
R6152 VGND.n1245 VGND.n1244 0.13638
R6153 VGND.n1241 VGND.n1225 0.13638
R6154 VGND.n1238 VGND.n1237 0.13638
R6155 VGND.n1234 VGND.n1232 0.13638
R6156 VGND.n1276 VGND.n1275 0.13638
R6157 VGND.n1280 VGND.n1279 0.13638
R6158 VGND.n991 VGND.n928 0.13638
R6159 VGND.n988 VGND.n987 0.13638
R6160 VGND.n983 VGND.n982 0.13638
R6161 VGND.n978 VGND.n977 0.13638
R6162 VGND.n973 VGND.n972 0.13638
R6163 VGND.n968 VGND.n967 0.13638
R6164 VGND.n963 VGND.n962 0.13638
R6165 VGND.n958 VGND.n957 0.13638
R6166 VGND.n953 VGND.n952 0.13638
R6167 VGND.n948 VGND.n947 0.13638
R6168 VGND.n943 VGND.n942 0.13638
R6169 VGND.n938 VGND.n937 0.13638
R6170 VGND.n933 VGND.n932 0.13638
R6171 VGND.n894 VGND.n890 0.13638
R6172 VGND.n1334 VGND.n1333 0.13638
R6173 VGND VGND.n190 0.120838
R6174 VGND.n19 VGND.n13 0.120292
R6175 VGND.n24 VGND.n13 0.120292
R6176 VGND.n25 VGND.n24 0.120292
R6177 VGND.n26 VGND.n25 0.120292
R6178 VGND.n26 VGND.n11 0.120292
R6179 VGND.n30 VGND.n11 0.120292
R6180 VGND.n31 VGND.n30 0.120292
R6181 VGND.n3008 VGND.n3007 0.120292
R6182 VGND.n3007 VGND.n3003 0.120292
R6183 VGND.n182 VGND.n174 0.120292
R6184 VGND.n183 VGND.n182 0.120292
R6185 VGND.n183 VGND.n168 0.120292
R6186 VGND.n188 VGND.n168 0.120292
R6187 VGND.n189 VGND.n188 0.120292
R6188 VGND.n2952 VGND.n2948 0.120292
R6189 VGND.n2957 VGND.n2948 0.120292
R6190 VGND.n2958 VGND.n2957 0.120292
R6191 VGND.n2959 VGND.n2958 0.120292
R6192 VGND.n2959 VGND.n2946 0.120292
R6193 VGND.n2963 VGND.n2946 0.120292
R6194 VGND.n2964 VGND.n2963 0.120292
R6195 VGND.n45 VGND.n39 0.120292
R6196 VGND.n50 VGND.n39 0.120292
R6197 VGND.n51 VGND.n50 0.120292
R6198 VGND.n52 VGND.n51 0.120292
R6199 VGND.n52 VGND.n37 0.120292
R6200 VGND.n56 VGND.n37 0.120292
R6201 VGND.n57 VGND.n56 0.120292
R6202 VGND.n63 VGND.n62 0.120292
R6203 VGND.n62 VGND.n58 0.120292
R6204 VGND.n106 VGND.n99 0.120292
R6205 VGND.n107 VGND.n106 0.120292
R6206 VGND.n107 VGND.n94 0.120292
R6207 VGND.n112 VGND.n94 0.120292
R6208 VGND.n113 VGND.n112 0.120292
R6209 VGND.n124 VGND.n91 0.120292
R6210 VGND.n83 VGND.n75 0.120292
R6211 VGND.n84 VGND.n83 0.120292
R6212 VGND.n84 VGND.n69 0.120292
R6213 VGND.n89 VGND.n69 0.120292
R6214 VGND.n90 VGND.n89 0.120292
R6215 VGND.n130 VGND.n127 0.120292
R6216 VGND.n151 VGND.n143 0.120292
R6217 VGND.n152 VGND.n151 0.120292
R6218 VGND.n152 VGND.n137 0.120292
R6219 VGND.n157 VGND.n137 0.120292
R6220 VGND.n158 VGND.n157 0.120292
R6221 VGND.n1152 VGND.n1151 0.120292
R6222 VGND.n1151 VGND.n1150 0.120292
R6223 VGND.n1150 VGND.n1136 0.120292
R6224 VGND.n1146 VGND.n1136 0.120292
R6225 VGND.n1146 VGND.n1145 0.120292
R6226 VGND.n1145 VGND.n1144 0.120292
R6227 VGND.n1130 VGND.n1129 0.120292
R6228 VGND.n1125 VGND.n1124 0.120292
R6229 VGND.n1124 VGND.n1123 0.120292
R6230 VGND.n1123 VGND.n1107 0.120292
R6231 VGND.n1119 VGND.n1107 0.120292
R6232 VGND.n1119 VGND.n1118 0.120292
R6233 VGND.n1118 VGND.n1117 0.120292
R6234 VGND.n499 VGND.n476 0.120292
R6235 VGND.n493 VGND.n476 0.120292
R6236 VGND.n493 VGND.n492 0.120292
R6237 VGND.n492 VGND.n480 0.120292
R6238 VGND.n485 VGND.n480 0.120292
R6239 VGND.n485 VGND.n484 0.120292
R6240 VGND.n484 VGND.n483 0.120292
R6241 VGND.n2280 VGND.n2257 0.120292
R6242 VGND.n2274 VGND.n2257 0.120292
R6243 VGND.n2274 VGND.n2273 0.120292
R6244 VGND.n2273 VGND.n2261 0.120292
R6245 VGND.n2266 VGND.n2261 0.120292
R6246 VGND.n2266 VGND.n2265 0.120292
R6247 VGND.n2265 VGND.n2264 0.120292
R6248 VGND.n510 VGND.n507 0.120292
R6249 VGND.n511 VGND.n510 0.120292
R6250 VGND.n535 VGND.n512 0.120292
R6251 VGND.n529 VGND.n512 0.120292
R6252 VGND.n529 VGND.n528 0.120292
R6253 VGND.n528 VGND.n516 0.120292
R6254 VGND.n521 VGND.n516 0.120292
R6255 VGND.n521 VGND.n520 0.120292
R6256 VGND.n520 VGND.n519 0.120292
R6257 VGND.n2214 VGND.n2213 0.120292
R6258 VGND.n2207 VGND.n2183 0.120292
R6259 VGND.n2202 VGND.n2183 0.120292
R6260 VGND.n2202 VGND.n2201 0.120292
R6261 VGND.n2198 VGND.n2197 0.120292
R6262 VGND.n2197 VGND.n2192 0.120292
R6263 VGND.n2193 VGND.n2192 0.120292
R6264 VGND.n2225 VGND.n2224 0.120292
R6265 VGND.n2245 VGND.n2244 0.120292
R6266 VGND.n2244 VGND.n2226 0.120292
R6267 VGND.n2240 VGND.n2226 0.120292
R6268 VGND.n2240 VGND.n2239 0.120292
R6269 VGND.n2239 VGND.n2238 0.120292
R6270 VGND.n2238 VGND.n2228 0.120292
R6271 VGND.n1363 VGND.n1362 0.120292
R6272 VGND.n1383 VGND.n1382 0.120292
R6273 VGND.n1382 VGND.n1364 0.120292
R6274 VGND.n1378 VGND.n1364 0.120292
R6275 VGND.n1378 VGND.n1377 0.120292
R6276 VGND.n1377 VGND.n1376 0.120292
R6277 VGND.n1376 VGND.n1366 0.120292
R6278 VGND.n2983 VGND.n2982 0.120292
R6279 VGND.n2983 VGND.n2975 0.120292
R6280 VGND.n2988 VGND.n2975 0.120292
R6281 VGND.n2989 VGND.n2988 0.120292
R6282 VGND.n2990 VGND.n2989 0.120292
R6283 VGND.n2990 VGND.n2973 0.120292
R6284 VGND.n2994 VGND.n2973 0.120292
R6285 VGND.n2996 VGND.n34 0.120292
R6286 VGND.n3000 VGND.n34 0.120292
R6287 VGND VGND.n161 0.119536
R6288 VGND.n1138 VGND 0.117202
R6289 VGND.n1109 VGND 0.117202
R6290 VGND.n2232 VGND 0.117202
R6291 VGND.n1370 VGND 0.117202
R6292 VGND.n287 VGND.n286 0.110872
R6293 VGND.n2788 VGND.n2787 0.110872
R6294 VGND.n2753 VGND.n2752 0.110872
R6295 VGND.n304 VGND.n303 0.110872
R6296 VGND.n2748 VGND.n2747 0.110872
R6297 VGND.n320 VGND.n319 0.110872
R6298 VGND.n2715 VGND.n2714 0.110872
R6299 VGND.n394 VGND.n393 0.110872
R6300 VGND.n2669 VGND.n2668 0.110872
R6301 VGND.n2664 VGND.n2663 0.110872
R6302 VGND.n2659 VGND.n2658 0.110872
R6303 VGND.n2654 VGND.n2653 0.110872
R6304 VGND.n2649 VGND.n2648 0.110872
R6305 VGND.n2644 VGND.n2643 0.110872
R6306 VGND.n2639 VGND.n2638 0.110872
R6307 VGND.n2536 VGND.n2535 0.110872
R6308 VGND.n2541 VGND.n2540 0.110872
R6309 VGND.n415 VGND.n414 0.110872
R6310 VGND.n2288 VGND.n2287 0.110872
R6311 VGND.n2293 VGND.n2292 0.110872
R6312 VGND.n2298 VGND.n2297 0.110872
R6313 VGND.n2303 VGND.n2302 0.110872
R6314 VGND.n2308 VGND.n2307 0.110872
R6315 VGND.n2313 VGND.n2312 0.110872
R6316 VGND.n2318 VGND.n2317 0.110872
R6317 VGND.n2323 VGND.n2322 0.110872
R6318 VGND.n2328 VGND.n2327 0.110872
R6319 VGND.n2333 VGND.n2332 0.110872
R6320 VGND.n2338 VGND.n2337 0.110872
R6321 VGND.n2343 VGND.n2342 0.110872
R6322 VGND.n2528 VGND.n2527 0.110872
R6323 VGND.n2522 VGND.n2521 0.110872
R6324 VGND.n2517 VGND.n2516 0.110872
R6325 VGND.n2512 VGND.n2511 0.110872
R6326 VGND.n428 VGND.n427 0.110872
R6327 VGND.n2481 VGND.n2480 0.110872
R6328 VGND.n436 VGND.n435 0.110872
R6329 VGND.n2455 VGND.n2454 0.110872
R6330 VGND.n444 VGND.n443 0.110872
R6331 VGND.n2429 VGND.n2428 0.110872
R6332 VGND.n452 VGND.n451 0.110872
R6333 VGND.n2403 VGND.n2402 0.110872
R6334 VGND.n460 VGND.n459 0.110872
R6335 VGND.n2377 VGND.n2376 0.110872
R6336 VGND.n472 VGND.n471 0.110872
R6337 VGND.n2816 VGND.n2815 0.110872
R6338 VGND.n2810 VGND.n2809 0.110872
R6339 VGND.n2499 VGND.n2498 0.110872
R6340 VGND.n424 VGND.n423 0.110872
R6341 VGND.n2494 VGND.n2493 0.110872
R6342 VGND.n432 VGND.n431 0.110872
R6343 VGND.n2468 VGND.n2467 0.110872
R6344 VGND.n440 VGND.n439 0.110872
R6345 VGND.n2442 VGND.n2441 0.110872
R6346 VGND.n448 VGND.n447 0.110872
R6347 VGND.n2416 VGND.n2415 0.110872
R6348 VGND.n456 VGND.n455 0.110872
R6349 VGND.n2390 VGND.n2389 0.110872
R6350 VGND.n464 VGND.n463 0.110872
R6351 VGND.n2364 VGND.n2363 0.110872
R6352 VGND.n1988 VGND.n1987 0.110872
R6353 VGND.n1982 VGND.n1981 0.110872
R6354 VGND.n1977 VGND.n1976 0.110872
R6355 VGND.n608 VGND.n607 0.110872
R6356 VGND.n1966 VGND.n1965 0.110872
R6357 VGND.n611 VGND.n610 0.110872
R6358 VGND.n1955 VGND.n1954 0.110872
R6359 VGND.n614 VGND.n613 0.110872
R6360 VGND.n1944 VGND.n1943 0.110872
R6361 VGND.n617 VGND.n616 0.110872
R6362 VGND.n1933 VGND.n1932 0.110872
R6363 VGND.n620 VGND.n619 0.110872
R6364 VGND.n1922 VGND.n1921 0.110872
R6365 VGND.n623 VGND.n622 0.110872
R6366 VGND.n1911 VGND.n1910 0.110872
R6367 VGND.n1995 VGND.n1994 0.110872
R6368 VGND.n2001 VGND.n2000 0.110872
R6369 VGND.n2006 VGND.n2005 0.110872
R6370 VGND.n2011 VGND.n2010 0.110872
R6371 VGND.n2016 VGND.n2015 0.110872
R6372 VGND.n2021 VGND.n2020 0.110872
R6373 VGND.n2026 VGND.n2025 0.110872
R6374 VGND.n2031 VGND.n2030 0.110872
R6375 VGND.n2036 VGND.n2035 0.110872
R6376 VGND.n2041 VGND.n2040 0.110872
R6377 VGND.n2046 VGND.n2045 0.110872
R6378 VGND.n2051 VGND.n2050 0.110872
R6379 VGND.n2056 VGND.n2055 0.110872
R6380 VGND.n594 VGND.n593 0.110872
R6381 VGND.n597 VGND.n596 0.110872
R6382 VGND.n2841 VGND.n2840 0.110872
R6383 VGND.n2835 VGND.n2834 0.110872
R6384 VGND.n2125 VGND.n2124 0.110872
R6385 VGND.n585 VGND.n584 0.110872
R6386 VGND.n2120 VGND.n2119 0.110872
R6387 VGND.n2115 VGND.n2114 0.110872
R6388 VGND.n2110 VGND.n2109 0.110872
R6389 VGND.n2105 VGND.n2104 0.110872
R6390 VGND.n2100 VGND.n2099 0.110872
R6391 VGND.n2095 VGND.n2094 0.110872
R6392 VGND.n2090 VGND.n2089 0.110872
R6393 VGND.n2085 VGND.n2084 0.110872
R6394 VGND.n2080 VGND.n2079 0.110872
R6395 VGND.n2075 VGND.n2074 0.110872
R6396 VGND.n2070 VGND.n2069 0.110872
R6397 VGND.n1828 VGND.n1827 0.110872
R6398 VGND.n1822 VGND.n1821 0.110872
R6399 VGND.n1817 VGND.n1816 0.110872
R6400 VGND.n1741 VGND.n1740 0.110872
R6401 VGND.n1806 VGND.n1805 0.110872
R6402 VGND.n1744 VGND.n1743 0.110872
R6403 VGND.n1795 VGND.n1794 0.110872
R6404 VGND.n1747 VGND.n1746 0.110872
R6405 VGND.n1784 VGND.n1783 0.110872
R6406 VGND.n1750 VGND.n1749 0.110872
R6407 VGND.n1773 VGND.n1772 0.110872
R6408 VGND.n1753 VGND.n1752 0.110872
R6409 VGND.n1762 VGND.n1761 0.110872
R6410 VGND.n1757 VGND.n1756 0.110872
R6411 VGND.n2177 VGND.n2176 0.110872
R6412 VGND.n1835 VGND.n1834 0.110872
R6413 VGND.n1841 VGND.n1840 0.110872
R6414 VGND.n1846 VGND.n1845 0.110872
R6415 VGND.n1673 VGND.n1672 0.110872
R6416 VGND.n1730 VGND.n1729 0.110872
R6417 VGND.n1725 VGND.n1724 0.110872
R6418 VGND.n1720 VGND.n1719 0.110872
R6419 VGND.n1715 VGND.n1714 0.110872
R6420 VGND.n1710 VGND.n1709 0.110872
R6421 VGND.n1705 VGND.n1704 0.110872
R6422 VGND.n1700 VGND.n1699 0.110872
R6423 VGND.n1695 VGND.n1694 0.110872
R6424 VGND.n1690 VGND.n1689 0.110872
R6425 VGND.n1676 VGND.n1675 0.110872
R6426 VGND.n1679 VGND.n1678 0.110872
R6427 VGND.n2866 VGND.n2865 0.110872
R6428 VGND.n2860 VGND.n2859 0.110872
R6429 VGND.n725 VGND.n724 0.110872
R6430 VGND.n667 VGND.n666 0.110872
R6431 VGND.n720 VGND.n719 0.110872
R6432 VGND.n715 VGND.n714 0.110872
R6433 VGND.n710 VGND.n709 0.110872
R6434 VGND.n705 VGND.n704 0.110872
R6435 VGND.n700 VGND.n699 0.110872
R6436 VGND.n695 VGND.n694 0.110872
R6437 VGND.n690 VGND.n689 0.110872
R6438 VGND.n685 VGND.n684 0.110872
R6439 VGND.n680 VGND.n679 0.110872
R6440 VGND.n675 VGND.n674 0.110872
R6441 VGND.n670 VGND.n669 0.110872
R6442 VGND.n1657 VGND.n1656 0.110872
R6443 VGND.n1662 VGND.n1661 0.110872
R6444 VGND.n735 VGND.n734 0.110872
R6445 VGND.n854 VGND.n853 0.110872
R6446 VGND.n820 VGND.n819 0.110872
R6447 VGND.n849 VGND.n848 0.110872
R6448 VGND.n844 VGND.n843 0.110872
R6449 VGND.n839 VGND.n838 0.110872
R6450 VGND.n834 VGND.n833 0.110872
R6451 VGND.n829 VGND.n828 0.110872
R6452 VGND.n824 VGND.n823 0.110872
R6453 VGND.n811 VGND.n810 0.110872
R6454 VGND.n870 VGND.n869 0.110872
R6455 VGND.n875 VGND.n874 0.110872
R6456 VGND.n1353 VGND.n1352 0.110872
R6457 VGND.n1649 VGND.n1648 0.110872
R6458 VGND.n1643 VGND.n1642 0.110872
R6459 VGND.n1638 VGND.n1637 0.110872
R6460 VGND.n1633 VGND.n1632 0.110872
R6461 VGND.n1553 VGND.n1552 0.110872
R6462 VGND.n761 VGND.n760 0.110872
R6463 VGND.n1548 VGND.n1547 0.110872
R6464 VGND.n1543 VGND.n1542 0.110872
R6465 VGND.n769 VGND.n768 0.110872
R6466 VGND.n1517 VGND.n1516 0.110872
R6467 VGND.n777 VGND.n776 0.110872
R6468 VGND.n1491 VGND.n1490 0.110872
R6469 VGND.n805 VGND.n804 0.110872
R6470 VGND.n1396 VGND.n1395 0.110872
R6471 VGND.n1391 VGND.n1390 0.110872
R6472 VGND.n2891 VGND.n2890 0.110872
R6473 VGND.n2885 VGND.n2884 0.110872
R6474 VGND.n1572 VGND.n1571 0.110872
R6475 VGND.n1577 VGND.n1576 0.110872
R6476 VGND.n1582 VGND.n1581 0.110872
R6477 VGND.n756 VGND.n755 0.110872
R6478 VGND.n1567 VGND.n1566 0.110872
R6479 VGND.n765 VGND.n764 0.110872
R6480 VGND.n1530 VGND.n1529 0.110872
R6481 VGND.n773 VGND.n772 0.110872
R6482 VGND.n1504 VGND.n1503 0.110872
R6483 VGND.n781 VGND.n780 0.110872
R6484 VGND.n1478 VGND.n1477 0.110872
R6485 VGND.n795 VGND.n794 0.110872
R6486 VGND.n1411 VGND.n1410 0.110872
R6487 VGND.n1609 VGND.n1608 0.110872
R6488 VGND.n1614 VGND.n1613 0.110872
R6489 VGND.n750 VGND.n749 0.110872
R6490 VGND.n1601 VGND.n1600 0.110872
R6491 VGND.n1596 VGND.n1595 0.110872
R6492 VGND.n1459 VGND.n1458 0.110872
R6493 VGND.n791 VGND.n790 0.110872
R6494 VGND.n1454 VGND.n1453 0.110872
R6495 VGND.n1449 VGND.n1448 0.110872
R6496 VGND.n1444 VGND.n1443 0.110872
R6497 VGND.n1439 VGND.n1438 0.110872
R6498 VGND.n1434 VGND.n1433 0.110872
R6499 VGND.n1429 VGND.n1428 0.110872
R6500 VGND.n1424 VGND.n1423 0.110872
R6501 VGND.n885 VGND.n884 0.110872
R6502 VGND.n2911 VGND.n2910 0.110872
R6503 VGND.n2905 VGND.n2904 0.110872
R6504 VGND.n1049 VGND.n1048 0.110872
R6505 VGND.n1058 VGND.n1057 0.110872
R6506 VGND.n1053 VGND.n1052 0.110872
R6507 VGND.n1044 VGND.n1043 0.110872
R6508 VGND.n1070 VGND.n1069 0.110872
R6509 VGND.n1075 VGND.n1074 0.110872
R6510 VGND.n1080 VGND.n1079 0.110872
R6511 VGND.n1085 VGND.n1084 0.110872
R6512 VGND.n1090 VGND.n1089 0.110872
R6513 VGND.n1095 VGND.n1094 0.110872
R6514 VGND.n1029 VGND.n1028 0.110872
R6515 VGND.n1037 VGND.n1036 0.110872
R6516 VGND.n1032 VGND.n1031 0.110872
R6517 VGND.n1169 VGND.n1168 0.110872
R6518 VGND.n1173 VGND.n1172 0.110872
R6519 VGND.n1179 VGND.n1178 0.110872
R6520 VGND.n1186 VGND.n1185 0.110872
R6521 VGND.n1009 VGND.n1008 0.110872
R6522 VGND.n1205 VGND.n1204 0.110872
R6523 VGND.n1211 VGND.n1210 0.110872
R6524 VGND.n1218 VGND.n1217 0.110872
R6525 VGND.n1222 VGND.n1001 0.110872
R6526 VGND.n1244 VGND.n1243 0.110872
R6527 VGND.n1227 VGND.n1225 0.110872
R6528 VGND.n1237 VGND.n1236 0.110872
R6529 VGND.n1232 VGND.n1231 0.110872
R6530 VGND.n1275 VGND.n1274 0.110872
R6531 VGND.n1281 VGND.n1280 0.110872
R6532 VGND.n928 VGND.n927 0.110872
R6533 VGND.n987 VGND.n986 0.110872
R6534 VGND.n982 VGND.n981 0.110872
R6535 VGND.n977 VGND.n976 0.110872
R6536 VGND.n972 VGND.n971 0.110872
R6537 VGND.n967 VGND.n966 0.110872
R6538 VGND.n962 VGND.n961 0.110872
R6539 VGND.n957 VGND.n956 0.110872
R6540 VGND.n952 VGND.n951 0.110872
R6541 VGND.n947 VGND.n946 0.110872
R6542 VGND.n942 VGND.n941 0.110872
R6543 VGND.n937 VGND.n936 0.110872
R6544 VGND.n932 VGND.n931 0.110872
R6545 VGND.n895 VGND.n894 0.110872
R6546 VGND.n1333 VGND.n1332 0.110872
R6547 VGND.n1130 VGND 0.0981562
R6548 VGND.n2214 VGND 0.0981562
R6549 VGND.n1362 VGND 0.0981562
R6550 VGND.n19 VGND 0.0968542
R6551 VGND.n2952 VGND 0.0968542
R6552 VGND.n45 VGND 0.0968542
R6553 VGND VGND.n91 0.0968542
R6554 VGND VGND.n130 0.0968542
R6555 VGND VGND.n499 0.0968542
R6556 VGND VGND.n2280 0.0968542
R6557 VGND VGND.n535 0.0968542
R6558 VGND VGND.n2207 0.0968542
R6559 VGND.n2224 VGND 0.0968542
R6560 VGND.n2982 VGND 0.0968542
R6561 VGND.n2562 VGND 0.088625
R6562 VGND.n2633 VGND 0.0790114
R6563 VGND.n2695 VGND 0.0790114
R6564 VGND.n2690 VGND 0.0790114
R6565 VGND VGND.n2689 0.0790114
R6566 VGND.n2684 VGND 0.0790114
R6567 VGND VGND.n2683 0.0790114
R6568 VGND.n2678 VGND 0.0790114
R6569 VGND VGND.n2677 0.0790114
R6570 VGND.n2709 VGND 0.0790114
R6571 VGND.n2723 VGND 0.0790114
R6572 VGND.n2742 VGND 0.0790114
R6573 VGND.n2761 VGND 0.0790114
R6574 VGND.n2781 VGND 0.0790114
R6575 VGND VGND.n2780 0.0790114
R6576 VGND VGND.n284 0.0790114
R6577 VGND.n2940 VGND 0.0790114
R6578 VGND.n2635 VGND 0.0790114
R6579 VGND.n2693 VGND 0.0790114
R6580 VGND VGND.n2692 0.0790114
R6581 VGND.n2687 VGND 0.0790114
R6582 VGND VGND.n2686 0.0790114
R6583 VGND.n2681 VGND 0.0790114
R6584 VGND VGND.n2680 0.0790114
R6585 VGND.n2675 VGND 0.0790114
R6586 VGND.n2711 VGND 0.0790114
R6587 VGND.n2721 VGND 0.0790114
R6588 VGND.n2744 VGND 0.0790114
R6589 VGND.n2759 VGND 0.0790114
R6590 VGND.n2783 VGND 0.0790114
R6591 VGND.n2784 VGND 0.0790114
R6592 VGND.n2794 VGND 0.0790114
R6593 VGND.n2937 VGND 0.0790114
R6594 VGND VGND.n2559 0.0790114
R6595 VGND VGND.n2558 0.0790114
R6596 VGND VGND.n2557 0.0790114
R6597 VGND VGND.n2556 0.0790114
R6598 VGND VGND.n2555 0.0790114
R6599 VGND VGND.n2554 0.0790114
R6600 VGND VGND.n2553 0.0790114
R6601 VGND VGND.n2552 0.0790114
R6602 VGND VGND.n2551 0.0790114
R6603 VGND VGND.n2550 0.0790114
R6604 VGND VGND.n2549 0.0790114
R6605 VGND VGND.n2548 0.0790114
R6606 VGND VGND.n2547 0.0790114
R6607 VGND.n2798 VGND 0.0790114
R6608 VGND VGND.n2797 0.0790114
R6609 VGND.n2533 VGND 0.0790114
R6610 VGND.n2357 VGND 0.0790114
R6611 VGND.n2373 VGND 0.0790114
R6612 VGND.n2383 VGND 0.0790114
R6613 VGND.n2399 VGND 0.0790114
R6614 VGND.n2409 VGND 0.0790114
R6615 VGND.n2425 VGND 0.0790114
R6616 VGND.n2435 VGND 0.0790114
R6617 VGND.n2451 VGND 0.0790114
R6618 VGND.n2461 VGND 0.0790114
R6619 VGND.n2477 VGND 0.0790114
R6620 VGND.n2487 VGND 0.0790114
R6621 VGND.n2508 VGND 0.0790114
R6622 VGND.n2802 VGND 0.0790114
R6623 VGND VGND.n2801 0.0790114
R6624 VGND.n419 VGND 0.0790114
R6625 VGND.n2530 VGND 0.0790114
R6626 VGND.n2360 VGND 0.0790114
R6627 VGND.n2370 VGND 0.0790114
R6628 VGND.n2386 VGND 0.0790114
R6629 VGND.n2396 VGND 0.0790114
R6630 VGND.n2412 VGND 0.0790114
R6631 VGND.n2422 VGND 0.0790114
R6632 VGND.n2438 VGND 0.0790114
R6633 VGND.n2448 VGND 0.0790114
R6634 VGND.n2464 VGND 0.0790114
R6635 VGND.n2474 VGND 0.0790114
R6636 VGND.n2490 VGND 0.0790114
R6637 VGND.n2505 VGND 0.0790114
R6638 VGND.n2805 VGND 0.0790114
R6639 VGND.n2806 VGND 0.0790114
R6640 VGND.n2819 VGND 0.0790114
R6641 VGND VGND.n2818 0.0790114
R6642 VGND.n1907 VGND 0.0790114
R6643 VGND.n1917 VGND 0.0790114
R6644 VGND.n1918 VGND 0.0790114
R6645 VGND.n1928 VGND 0.0790114
R6646 VGND.n1929 VGND 0.0790114
R6647 VGND.n1939 VGND 0.0790114
R6648 VGND.n1940 VGND 0.0790114
R6649 VGND.n1950 VGND 0.0790114
R6650 VGND.n1951 VGND 0.0790114
R6651 VGND.n1961 VGND 0.0790114
R6652 VGND.n1962 VGND 0.0790114
R6653 VGND.n1972 VGND 0.0790114
R6654 VGND.n1973 VGND 0.0790114
R6655 VGND.n2823 VGND 0.0790114
R6656 VGND VGND.n2822 0.0790114
R6657 VGND.n1990 VGND 0.0790114
R6658 VGND.n2063 VGND 0.0790114
R6659 VGND VGND.n2062 0.0790114
R6660 VGND.n2167 VGND 0.0790114
R6661 VGND VGND.n2166 0.0790114
R6662 VGND.n2159 VGND 0.0790114
R6663 VGND VGND.n2158 0.0790114
R6664 VGND.n2151 VGND 0.0790114
R6665 VGND VGND.n2150 0.0790114
R6666 VGND.n2143 VGND 0.0790114
R6667 VGND VGND.n2142 0.0790114
R6668 VGND.n2135 VGND 0.0790114
R6669 VGND VGND.n2134 0.0790114
R6670 VGND.n2827 VGND 0.0790114
R6671 VGND VGND.n2826 0.0790114
R6672 VGND.n1998 VGND 0.0790114
R6673 VGND VGND.n1997 0.0790114
R6674 VGND.n2066 VGND 0.0790114
R6675 VGND.n2171 VGND 0.0790114
R6676 VGND VGND.n2170 0.0790114
R6677 VGND.n2163 VGND 0.0790114
R6678 VGND VGND.n2162 0.0790114
R6679 VGND.n2155 VGND 0.0790114
R6680 VGND VGND.n2154 0.0790114
R6681 VGND.n2147 VGND 0.0790114
R6682 VGND VGND.n2146 0.0790114
R6683 VGND.n2139 VGND 0.0790114
R6684 VGND VGND.n2138 0.0790114
R6685 VGND.n2131 VGND 0.0790114
R6686 VGND.n2830 VGND 0.0790114
R6687 VGND.n2831 VGND 0.0790114
R6688 VGND.n2844 VGND 0.0790114
R6689 VGND VGND.n2843 0.0790114
R6690 VGND VGND.n1901 0.0790114
R6691 VGND.n2174 VGND 0.0790114
R6692 VGND.n1758 VGND 0.0790114
R6693 VGND.n1768 VGND 0.0790114
R6694 VGND.n1769 VGND 0.0790114
R6695 VGND.n1779 VGND 0.0790114
R6696 VGND.n1780 VGND 0.0790114
R6697 VGND.n1790 VGND 0.0790114
R6698 VGND.n1791 VGND 0.0790114
R6699 VGND.n1801 VGND 0.0790114
R6700 VGND.n1802 VGND 0.0790114
R6701 VGND.n1812 VGND 0.0790114
R6702 VGND.n1813 VGND 0.0790114
R6703 VGND.n2848 VGND 0.0790114
R6704 VGND VGND.n2847 0.0790114
R6705 VGND.n1830 VGND 0.0790114
R6706 VGND VGND.n1899 0.0790114
R6707 VGND.n1685 VGND 0.0790114
R6708 VGND.n1686 VGND 0.0790114
R6709 VGND.n1884 VGND 0.0790114
R6710 VGND VGND.n1883 0.0790114
R6711 VGND.n1876 VGND 0.0790114
R6712 VGND VGND.n1875 0.0790114
R6713 VGND.n1868 VGND 0.0790114
R6714 VGND VGND.n1867 0.0790114
R6715 VGND.n1860 VGND 0.0790114
R6716 VGND VGND.n1859 0.0790114
R6717 VGND.n1852 VGND 0.0790114
R6718 VGND.n2852 VGND 0.0790114
R6719 VGND VGND.n2851 0.0790114
R6720 VGND.n1838 VGND 0.0790114
R6721 VGND VGND.n1837 0.0790114
R6722 VGND.n1896 VGND 0.0790114
R6723 VGND VGND.n1895 0.0790114
R6724 VGND.n1888 VGND 0.0790114
R6725 VGND VGND.n1887 0.0790114
R6726 VGND.n1880 VGND 0.0790114
R6727 VGND VGND.n1879 0.0790114
R6728 VGND.n1872 VGND 0.0790114
R6729 VGND VGND.n1871 0.0790114
R6730 VGND.n1864 VGND 0.0790114
R6731 VGND VGND.n1863 0.0790114
R6732 VGND.n1856 VGND 0.0790114
R6733 VGND VGND.n1855 0.0790114
R6734 VGND.n2855 VGND 0.0790114
R6735 VGND.n2856 VGND 0.0790114
R6736 VGND.n2869 VGND 0.0790114
R6737 VGND VGND.n2868 0.0790114
R6738 VGND.n1349 VGND 0.0790114
R6739 VGND.n1892 VGND 0.0790114
R6740 VGND VGND.n1891 0.0790114
R6741 VGND.n867 VGND 0.0790114
R6742 VGND VGND.n866 0.0790114
R6743 VGND VGND.n865 0.0790114
R6744 VGND VGND.n864 0.0790114
R6745 VGND VGND.n863 0.0790114
R6746 VGND VGND.n862 0.0790114
R6747 VGND VGND.n861 0.0790114
R6748 VGND VGND.n860 0.0790114
R6749 VGND.n1669 VGND 0.0790114
R6750 VGND VGND.n1668 0.0790114
R6751 VGND.n2873 VGND 0.0790114
R6752 VGND VGND.n2872 0.0790114
R6753 VGND.n1654 VGND 0.0790114
R6754 VGND.n1404 VGND 0.0790114
R6755 VGND VGND.n1403 0.0790114
R6756 VGND VGND.n1402 0.0790114
R6757 VGND.n1487 VGND 0.0790114
R6758 VGND.n1497 VGND 0.0790114
R6759 VGND.n1513 VGND 0.0790114
R6760 VGND.n1523 VGND 0.0790114
R6761 VGND.n1539 VGND 0.0790114
R6762 VGND.n1560 VGND 0.0790114
R6763 VGND VGND.n1559 0.0790114
R6764 VGND.n1628 VGND 0.0790114
R6765 VGND.n1629 VGND 0.0790114
R6766 VGND.n2877 VGND 0.0790114
R6767 VGND VGND.n2876 0.0790114
R6768 VGND.n740 VGND 0.0790114
R6769 VGND.n1651 VGND 0.0790114
R6770 VGND.n1407 VGND 0.0790114
R6771 VGND.n1417 VGND 0.0790114
R6772 VGND.n1474 VGND 0.0790114
R6773 VGND.n1484 VGND 0.0790114
R6774 VGND.n1500 VGND 0.0790114
R6775 VGND.n1510 VGND 0.0790114
R6776 VGND.n1526 VGND 0.0790114
R6777 VGND.n1536 VGND 0.0790114
R6778 VGND.n1563 VGND 0.0790114
R6779 VGND.n1588 VGND 0.0790114
R6780 VGND.n1625 VGND 0.0790114
R6781 VGND VGND.n1624 0.0790114
R6782 VGND.n2880 VGND 0.0790114
R6783 VGND.n2881 VGND 0.0790114
R6784 VGND.n2894 VGND 0.0790114
R6785 VGND VGND.n2893 0.0790114
R6786 VGND VGND.n1344 0.0790114
R6787 VGND.n1420 VGND 0.0790114
R6788 VGND.n1471 VGND 0.0790114
R6789 VGND VGND.n1470 0.0790114
R6790 VGND VGND.n1469 0.0790114
R6791 VGND VGND.n1468 0.0790114
R6792 VGND VGND.n1467 0.0790114
R6793 VGND VGND.n1466 0.0790114
R6794 VGND VGND.n1465 0.0790114
R6795 VGND.n1591 VGND 0.0790114
R6796 VGND.n1592 VGND 0.0790114
R6797 VGND.n1621 VGND 0.0790114
R6798 VGND VGND.n1620 0.0790114
R6799 VGND.n2898 VGND 0.0790114
R6800 VGND VGND.n2897 0.0790114
R6801 VGND.n1606 VGND 0.0790114
R6802 VGND.n1103 VGND 0.0790114
R6803 VGND VGND.n1102 0.0790114
R6804 VGND VGND.n1101 0.0790114
R6805 VGND.n1321 VGND 0.0790114
R6806 VGND VGND.n1320 0.0790114
R6807 VGND.n1313 VGND 0.0790114
R6808 VGND VGND.n1312 0.0790114
R6809 VGND.n1305 VGND 0.0790114
R6810 VGND VGND.n1304 0.0790114
R6811 VGND.n1067 VGND 0.0790114
R6812 VGND VGND.n1066 0.0790114
R6813 VGND VGND.n1065 0.0790114
R6814 VGND VGND.n1064 0.0790114
R6815 VGND.n2901 VGND 0.0790114
R6816 VGND.n233 VGND 0.0790114
R6817 VGND.n2913 VGND 0.0790114
R6818 VGND.n1163 VGND 0.0790114
R6819 VGND.n1328 VGND 0.0790114
R6820 VGND VGND.n1327 0.0790114
R6821 VGND.n898 VGND 0.0790114
R6822 VGND.n901 VGND 0.0790114
R6823 VGND.n904 VGND 0.0790114
R6824 VGND.n907 VGND 0.0790114
R6825 VGND.n910 VGND 0.0790114
R6826 VGND.n913 VGND 0.0790114
R6827 VGND.n1298 VGND 0.0790114
R6828 VGND VGND.n1297 0.0790114
R6829 VGND.n1292 VGND 0.0790114
R6830 VGND VGND.n1291 0.0790114
R6831 VGND.n1270 VGND 0.0790114
R6832 VGND.n1285 VGND 0.0790114
R6833 VGND VGND.n1284 0.0790114
R6834 VGND.n1161 VGND 0.0790114
R6835 VGND.n1330 VGND 0.0790114
R6836 VGND.n1325 VGND 0.0790114
R6837 VGND VGND.n1324 0.0790114
R6838 VGND.n1317 VGND 0.0790114
R6839 VGND VGND.n1316 0.0790114
R6840 VGND.n1309 VGND 0.0790114
R6841 VGND VGND.n1308 0.0790114
R6842 VGND.n1301 VGND 0.0790114
R6843 VGND VGND.n1300 0.0790114
R6844 VGND.n1295 VGND 0.0790114
R6845 VGND VGND.n1294 0.0790114
R6846 VGND.n1289 VGND 0.0790114
R6847 VGND VGND.n1288 0.0790114
R6848 VGND VGND.n1287 0.0790114
R6849 VGND.n2916 VGND 0.0790114
R6850 VGND.n2699 VGND.n2698 0.0656596
R6851 VGND.n357 VGND.n355 0.0656596
R6852 VGND.n364 VGND.n362 0.0656596
R6853 VGND.n368 VGND.n367 0.0656596
R6854 VGND.n375 VGND.n373 0.0656596
R6855 VGND.n379 VGND.n378 0.0656596
R6856 VGND.n386 VGND.n384 0.0656596
R6857 VGND.n387 VGND.n325 0.0656596
R6858 VGND.n326 VGND.n314 0.0656596
R6859 VGND.n2726 VGND.n309 0.0656596
R6860 VGND.n312 VGND.n311 0.0656596
R6861 VGND.n2735 VGND.n2734 0.0656596
R6862 VGND.n2730 VGND.n293 0.0656596
R6863 VGND.n296 VGND.n294 0.0656596
R6864 VGND.n2773 VGND.n203 0.0656596
R6865 VGND.n2606 VGND 0.063
R6866 VGND.n2603 VGND 0.063
R6867 VGND.n2600 VGND 0.063
R6868 VGND.n2597 VGND 0.063
R6869 VGND.n2594 VGND 0.063
R6870 VGND.n2591 VGND 0.063
R6871 VGND.n2588 VGND 0.063
R6872 VGND.n2585 VGND 0.063
R6873 VGND.n2582 VGND 0.063
R6874 VGND.n2579 VGND 0.063
R6875 VGND.n2576 VGND 0.063
R6876 VGND.n2573 VGND 0.063
R6877 VGND.n2570 VGND 0.063
R6878 VGND.n2567 VGND 0.063
R6879 VGND.n2564 VGND 0.063
R6880 VGND VGND.n31 0.0603958
R6881 VGND.n3009 VGND 0.0603958
R6882 VGND VGND.n3008 0.0603958
R6883 VGND.n192 VGND 0.0603958
R6884 VGND VGND.n191 0.0603958
R6885 VGND VGND.n2964 0.0603958
R6886 VGND.n2965 VGND 0.0603958
R6887 VGND VGND.n57 0.0603958
R6888 VGND.n64 VGND 0.0603958
R6889 VGND VGND.n63 0.0603958
R6890 VGND.n118 VGND 0.0603958
R6891 VGND.n119 VGND 0.0603958
R6892 VGND.n132 VGND 0.0603958
R6893 VGND VGND.n131 0.0603958
R6894 VGND.n127 VGND 0.0603958
R6895 VGND.n163 VGND 0.0603958
R6896 VGND VGND.n162 0.0603958
R6897 VGND.n1152 VGND 0.0603958
R6898 VGND.n1129 VGND 0.0603958
R6899 VGND VGND.n1128 0.0603958
R6900 VGND.n1125 VGND 0.0603958
R6901 VGND.n501 VGND 0.0603958
R6902 VGND VGND.n500 0.0603958
R6903 VGND.n483 VGND 0.0603958
R6904 VGND.n2282 VGND 0.0603958
R6905 VGND VGND.n2281 0.0603958
R6906 VGND.n2264 VGND 0.0603958
R6907 VGND.n537 VGND 0.0603958
R6908 VGND VGND.n536 0.0603958
R6909 VGND.n519 VGND 0.0603958
R6910 VGND.n2209 VGND 0.0603958
R6911 VGND VGND.n2208 0.0603958
R6912 VGND.n2201 VGND 0.0603958
R6913 VGND.n2198 VGND 0.0603958
R6914 VGND.n2193 VGND 0.0603958
R6915 VGND VGND.n2225 0.0603958
R6916 VGND.n2246 VGND 0.0603958
R6917 VGND VGND.n2245 0.0603958
R6918 VGND VGND.n1363 0.0603958
R6919 VGND.n1384 VGND 0.0603958
R6920 VGND VGND.n1383 0.0603958
R6921 VGND VGND.n2994 0.0603958
R6922 VGND.n2995 VGND 0.0603958
R6923 VGND.n2996 VGND 0.0603958
R6924 VGND.n2698 VGND 0.0574853
R6925 VGND.n357 VGND 0.0574853
R6926 VGND.n364 VGND 0.0574853
R6927 VGND.n367 VGND 0.0574853
R6928 VGND.n375 VGND 0.0574853
R6929 VGND.n378 VGND 0.0574853
R6930 VGND.n386 VGND 0.0574853
R6931 VGND.n325 VGND 0.0574853
R6932 VGND.n314 VGND 0.0574853
R6933 VGND.n309 VGND 0.0574853
R6934 VGND.n311 VGND 0.0574853
R6935 VGND.n2734 VGND 0.0574853
R6936 VGND.n293 VGND 0.0574853
R6937 VGND.n296 VGND 0.0574853
R6938 VGND.n203 VGND 0.0574853
R6939 VGND.n1021 VGND 0.0489375
R6940 VGND.n994 VGND 0.0489375
R6941 VGND.n2630 VGND 0.0489375
R6942 VGND.n204 VGND 0.0489375
R6943 VGND.n334 VGND 0.0489375
R6944 VGND.n2626 VGND 0.0489375
R6945 VGND.n2623 VGND 0.0489375
R6946 VGND.n2620 VGND 0.0489375
R6947 VGND.n2617 VGND 0.0489375
R6948 VGND.n2614 VGND 0.0489375
R6949 VGND.n2611 VGND 0.0489375
R6950 VGND.n322 VGND 0.0489375
R6951 VGND.n315 VGND 0.0489375
R6952 VGND.n306 VGND 0.0489375
R6953 VGND.n299 VGND 0.0489375
R6954 VGND.n2765 VGND 0.0489375
R6955 VGND.n290 VGND 0.0489375
R6956 VGND.n297 VGND 0.0489375
R6957 VGND.n1018 VGND 0.0489375
R6958 VGND.n1015 VGND 0.0489375
R6959 VGND.n1180 VGND 0.0489375
R6960 VGND.n1006 VGND 0.0489375
R6961 VGND.n1004 VGND 0.0489375
R6962 VGND.n1195 VGND 0.0489375
R6963 VGND.n1212 VGND 0.0489375
R6964 VGND.n1000 VGND 0.0489375
R6965 VGND.n1253 VGND 0.0489375
R6966 VGND.n1256 VGND 0.0489375
R6967 VGND.n1259 VGND 0.0489375
R6968 VGND.n1262 VGND 0.0489375
R6969 VGND.n998 VGND 0.0489375
R6970 VGND.n1265 VGND 0.0489375
R6971 VGND VGND.n330 0.037734
R6972 VGND.n286 VGND 0.037734
R6973 VGND.n2787 VGND 0.037734
R6974 VGND.n2752 VGND 0.037734
R6975 VGND.n303 VGND 0.037734
R6976 VGND.n2747 VGND 0.037734
R6977 VGND.n319 VGND 0.037734
R6978 VGND.n2714 VGND 0.037734
R6979 VGND.n393 VGND 0.037734
R6980 VGND.n2668 VGND 0.037734
R6981 VGND.n2663 VGND 0.037734
R6982 VGND.n2658 VGND 0.037734
R6983 VGND.n2653 VGND 0.037734
R6984 VGND.n2648 VGND 0.037734
R6985 VGND.n2643 VGND 0.037734
R6986 VGND.n2638 VGND 0.037734
R6987 VGND VGND.n396 0.037734
R6988 VGND.n2535 VGND 0.037734
R6989 VGND.n2540 VGND 0.037734
R6990 VGND.n414 VGND 0.037734
R6991 VGND.n2287 VGND 0.037734
R6992 VGND.n2292 VGND 0.037734
R6993 VGND.n2297 VGND 0.037734
R6994 VGND.n2302 VGND 0.037734
R6995 VGND.n2307 VGND 0.037734
R6996 VGND.n2312 VGND 0.037734
R6997 VGND.n2317 VGND 0.037734
R6998 VGND.n2322 VGND 0.037734
R6999 VGND.n2327 VGND 0.037734
R7000 VGND.n2332 VGND 0.037734
R7001 VGND.n2337 VGND 0.037734
R7002 VGND.n2342 VGND 0.037734
R7003 VGND VGND.n400 0.037734
R7004 VGND VGND.n2528 0.037734
R7005 VGND.n2521 VGND 0.037734
R7006 VGND.n2516 VGND 0.037734
R7007 VGND.n2511 VGND 0.037734
R7008 VGND.n427 VGND 0.037734
R7009 VGND.n2480 VGND 0.037734
R7010 VGND.n435 VGND 0.037734
R7011 VGND.n2454 VGND 0.037734
R7012 VGND.n443 VGND 0.037734
R7013 VGND.n2428 VGND 0.037734
R7014 VGND.n451 VGND 0.037734
R7015 VGND.n2402 VGND 0.037734
R7016 VGND.n459 VGND 0.037734
R7017 VGND.n2376 VGND 0.037734
R7018 VGND.n471 VGND 0.037734
R7019 VGND VGND.n469 0.037734
R7020 VGND VGND.n2816 0.037734
R7021 VGND.n2809 VGND 0.037734
R7022 VGND.n2498 VGND 0.037734
R7023 VGND.n423 VGND 0.037734
R7024 VGND.n2493 VGND 0.037734
R7025 VGND.n431 VGND 0.037734
R7026 VGND.n2467 VGND 0.037734
R7027 VGND.n439 VGND 0.037734
R7028 VGND.n2441 VGND 0.037734
R7029 VGND.n447 VGND 0.037734
R7030 VGND.n2415 VGND 0.037734
R7031 VGND.n455 VGND 0.037734
R7032 VGND.n2389 VGND 0.037734
R7033 VGND.n463 VGND 0.037734
R7034 VGND.n2363 VGND 0.037734
R7035 VGND VGND.n466 0.037734
R7036 VGND VGND.n1988 0.037734
R7037 VGND.n1981 VGND 0.037734
R7038 VGND.n1976 VGND 0.037734
R7039 VGND.n607 VGND 0.037734
R7040 VGND.n1965 VGND 0.037734
R7041 VGND.n610 VGND 0.037734
R7042 VGND.n1954 VGND 0.037734
R7043 VGND.n613 VGND 0.037734
R7044 VGND.n1943 VGND 0.037734
R7045 VGND.n616 VGND 0.037734
R7046 VGND.n1932 VGND 0.037734
R7047 VGND.n619 VGND 0.037734
R7048 VGND.n1921 VGND 0.037734
R7049 VGND.n622 VGND 0.037734
R7050 VGND.n1910 VGND 0.037734
R7051 VGND VGND.n625 0.037734
R7052 VGND VGND.n1995 0.037734
R7053 VGND.n2000 VGND 0.037734
R7054 VGND.n2005 VGND 0.037734
R7055 VGND.n2010 VGND 0.037734
R7056 VGND.n2015 VGND 0.037734
R7057 VGND.n2020 VGND 0.037734
R7058 VGND.n2025 VGND 0.037734
R7059 VGND.n2030 VGND 0.037734
R7060 VGND.n2035 VGND 0.037734
R7061 VGND.n2040 VGND 0.037734
R7062 VGND.n2045 VGND 0.037734
R7063 VGND.n2050 VGND 0.037734
R7064 VGND.n2055 VGND 0.037734
R7065 VGND.n593 VGND 0.037734
R7066 VGND.n596 VGND 0.037734
R7067 VGND VGND.n590 0.037734
R7068 VGND VGND.n2841 0.037734
R7069 VGND.n2834 VGND 0.037734
R7070 VGND.n2124 VGND 0.037734
R7071 VGND.n584 VGND 0.037734
R7072 VGND.n2119 VGND 0.037734
R7073 VGND.n2114 VGND 0.037734
R7074 VGND.n2109 VGND 0.037734
R7075 VGND.n2104 VGND 0.037734
R7076 VGND.n2099 VGND 0.037734
R7077 VGND.n2094 VGND 0.037734
R7078 VGND.n2089 VGND 0.037734
R7079 VGND.n2084 VGND 0.037734
R7080 VGND.n2079 VGND 0.037734
R7081 VGND.n2074 VGND 0.037734
R7082 VGND.n2069 VGND 0.037734
R7083 VGND VGND.n587 0.037734
R7084 VGND VGND.n1828 0.037734
R7085 VGND.n1821 VGND 0.037734
R7086 VGND.n1816 VGND 0.037734
R7087 VGND.n1740 VGND 0.037734
R7088 VGND.n1805 VGND 0.037734
R7089 VGND.n1743 VGND 0.037734
R7090 VGND.n1794 VGND 0.037734
R7091 VGND.n1746 VGND 0.037734
R7092 VGND.n1783 VGND 0.037734
R7093 VGND.n1749 VGND 0.037734
R7094 VGND.n1772 VGND 0.037734
R7095 VGND.n1752 VGND 0.037734
R7096 VGND.n1761 VGND 0.037734
R7097 VGND VGND.n1757 0.037734
R7098 VGND.n2176 VGND 0.037734
R7099 VGND VGND.n547 0.037734
R7100 VGND VGND.n1835 0.037734
R7101 VGND.n1840 VGND 0.037734
R7102 VGND.n1845 VGND 0.037734
R7103 VGND.n1672 VGND 0.037734
R7104 VGND.n1729 VGND 0.037734
R7105 VGND.n1724 VGND 0.037734
R7106 VGND.n1719 VGND 0.037734
R7107 VGND.n1714 VGND 0.037734
R7108 VGND.n1709 VGND 0.037734
R7109 VGND.n1704 VGND 0.037734
R7110 VGND.n1699 VGND 0.037734
R7111 VGND.n1694 VGND 0.037734
R7112 VGND.n1689 VGND 0.037734
R7113 VGND.n1675 VGND 0.037734
R7114 VGND.n1678 VGND 0.037734
R7115 VGND VGND.n628 0.037734
R7116 VGND VGND.n2866 0.037734
R7117 VGND.n2859 VGND 0.037734
R7118 VGND.n724 VGND 0.037734
R7119 VGND.n666 VGND 0.037734
R7120 VGND.n719 VGND 0.037734
R7121 VGND.n714 VGND 0.037734
R7122 VGND.n709 VGND 0.037734
R7123 VGND.n704 VGND 0.037734
R7124 VGND.n699 VGND 0.037734
R7125 VGND.n694 VGND 0.037734
R7126 VGND.n689 VGND 0.037734
R7127 VGND.n684 VGND 0.037734
R7128 VGND.n679 VGND 0.037734
R7129 VGND.n674 VGND 0.037734
R7130 VGND.n669 VGND 0.037734
R7131 VGND VGND.n632 0.037734
R7132 VGND.n1656 VGND 0.037734
R7133 VGND.n1661 VGND 0.037734
R7134 VGND.n734 VGND 0.037734
R7135 VGND.n853 VGND 0.037734
R7136 VGND.n819 VGND 0.037734
R7137 VGND.n848 VGND 0.037734
R7138 VGND.n843 VGND 0.037734
R7139 VGND.n838 VGND 0.037734
R7140 VGND.n833 VGND 0.037734
R7141 VGND.n828 VGND 0.037734
R7142 VGND.n823 VGND 0.037734
R7143 VGND VGND.n811 0.037734
R7144 VGND.n869 VGND 0.037734
R7145 VGND.n874 VGND 0.037734
R7146 VGND.n1352 VGND 0.037734
R7147 VGND VGND.n879 0.037734
R7148 VGND VGND.n1649 0.037734
R7149 VGND.n1642 VGND 0.037734
R7150 VGND.n1637 VGND 0.037734
R7151 VGND.n1632 VGND 0.037734
R7152 VGND.n1552 VGND 0.037734
R7153 VGND.n760 VGND 0.037734
R7154 VGND.n1547 VGND 0.037734
R7155 VGND.n1542 VGND 0.037734
R7156 VGND.n768 VGND 0.037734
R7157 VGND.n1516 VGND 0.037734
R7158 VGND.n776 VGND 0.037734
R7159 VGND.n1490 VGND 0.037734
R7160 VGND.n804 VGND 0.037734
R7161 VGND.n1395 VGND 0.037734
R7162 VGND.n1390 VGND 0.037734
R7163 VGND VGND.n800 0.037734
R7164 VGND VGND.n2891 0.037734
R7165 VGND.n2884 VGND 0.037734
R7166 VGND.n1571 VGND 0.037734
R7167 VGND.n1576 VGND 0.037734
R7168 VGND.n1581 VGND 0.037734
R7169 VGND.n755 VGND 0.037734
R7170 VGND.n1566 VGND 0.037734
R7171 VGND.n764 VGND 0.037734
R7172 VGND.n1529 VGND 0.037734
R7173 VGND.n772 VGND 0.037734
R7174 VGND.n1503 VGND 0.037734
R7175 VGND.n780 VGND 0.037734
R7176 VGND.n1477 VGND 0.037734
R7177 VGND.n794 VGND 0.037734
R7178 VGND.n1410 VGND 0.037734
R7179 VGND VGND.n797 0.037734
R7180 VGND.n1608 VGND 0.037734
R7181 VGND.n1613 VGND 0.037734
R7182 VGND.n749 VGND 0.037734
R7183 VGND.n1600 VGND 0.037734
R7184 VGND.n1595 VGND 0.037734
R7185 VGND.n1458 VGND 0.037734
R7186 VGND.n790 VGND 0.037734
R7187 VGND.n1453 VGND 0.037734
R7188 VGND.n1448 VGND 0.037734
R7189 VGND.n1443 VGND 0.037734
R7190 VGND.n1438 VGND 0.037734
R7191 VGND.n1433 VGND 0.037734
R7192 VGND.n1428 VGND 0.037734
R7193 VGND.n1423 VGND 0.037734
R7194 VGND.n884 VGND 0.037734
R7195 VGND VGND.n882 0.037734
R7196 VGND VGND.n2911 0.037734
R7197 VGND.n2904 VGND 0.037734
R7198 VGND.n1048 VGND 0.037734
R7199 VGND.n1057 VGND 0.037734
R7200 VGND.n1052 VGND 0.037734
R7201 VGND VGND.n1044 0.037734
R7202 VGND.n1069 VGND 0.037734
R7203 VGND.n1074 VGND 0.037734
R7204 VGND.n1079 VGND 0.037734
R7205 VGND.n1084 VGND 0.037734
R7206 VGND.n1089 VGND 0.037734
R7207 VGND.n1094 VGND 0.037734
R7208 VGND.n1028 VGND 0.037734
R7209 VGND.n1036 VGND 0.037734
R7210 VGND.n1031 VGND 0.037734
R7211 VGND VGND.n1024 0.037734
R7212 VGND VGND.n1014 0.037734
R7213 VGND VGND.n1169 0.037734
R7214 VGND.n1172 VGND 0.037734
R7215 VGND VGND.n1179 0.037734
R7216 VGND.n1185 VGND 0.037734
R7217 VGND.n1008 VGND 0.037734
R7218 VGND.n1204 VGND 0.037734
R7219 VGND VGND.n1211 0.037734
R7220 VGND.n1217 VGND 0.037734
R7221 VGND VGND.n1222 0.037734
R7222 VGND.n1243 VGND 0.037734
R7223 VGND VGND.n1227 0.037734
R7224 VGND.n1236 VGND 0.037734
R7225 VGND.n1231 VGND 0.037734
R7226 VGND.n1274 VGND 0.037734
R7227 VGND VGND.n1281 0.037734
R7228 VGND.n927 VGND 0.037734
R7229 VGND.n986 VGND 0.037734
R7230 VGND.n981 VGND 0.037734
R7231 VGND.n976 VGND 0.037734
R7232 VGND.n971 VGND 0.037734
R7233 VGND.n966 VGND 0.037734
R7234 VGND.n961 VGND 0.037734
R7235 VGND.n956 VGND 0.037734
R7236 VGND.n951 VGND 0.037734
R7237 VGND.n946 VGND 0.037734
R7238 VGND.n941 VGND 0.037734
R7239 VGND.n936 VGND 0.037734
R7240 VGND.n931 VGND 0.037734
R7241 VGND VGND.n895 0.037734
R7242 VGND.n1332 VGND 0.037734
R7243 VGND VGND.n887 0.037734
R7244 VGND.n1156 VGND 0.0343542
R7245 VGND.n1128 VGND 0.0343542
R7246 VGND.n501 VGND 0.0343542
R7247 VGND.n2282 VGND 0.0343542
R7248 VGND.n537 VGND 0.0343542
R7249 VGND.n2209 VGND 0.0343542
R7250 VGND.n2246 VGND 0.0343542
R7251 VGND.n1384 VGND 0.0343542
R7252 VGND.n3009 VGND 0.0330521
R7253 VGND.n192 VGND 0.0330521
R7254 VGND.n2965 VGND 0.0330521
R7255 VGND.n64 VGND 0.0330521
R7256 VGND VGND.n118 0.0330521
R7257 VGND.n132 VGND 0.0330521
R7258 VGND.n163 VGND 0.0330521
R7259 VGND VGND.n2995 0.0330521
R7260 VGND.n33 VGND 0.024
R7261 VGND.n1 VGND 0.024
R7262 VGND.n119 VGND 0.0239375
R7263 VGND.n131 VGND 0.0239375
R7264 VGND.n500 VGND 0.0239375
R7265 VGND.n2281 VGND 0.0239375
R7266 VGND.n536 VGND 0.0239375
R7267 VGND.n3003 VGND 0.0226354
R7268 VGND VGND.n124 0.0226354
R7269 VGND.n1133 VGND 0.0226354
R7270 VGND VGND.n2256 0.0226354
R7271 VGND.n2217 VGND 0.0226354
R7272 VGND.n2208 VGND 0.0226354
R7273 VGND.n2220 VGND 0.0226354
R7274 VGND VGND.n3000 0.0226354
R7275 VGND VGND.n189 0.0213333
R7276 VGND.n191 VGND 0.0213333
R7277 VGND.n58 VGND 0.0213333
R7278 VGND.n113 VGND 0.0213333
R7279 VGND VGND.n90 0.0213333
R7280 VGND VGND.n158 0.0213333
R7281 VGND.n162 VGND 0.0213333
R7282 VGND VGND.n511 0.0213333
R7283 VGND.n2213 VGND 0.0213333
R7284 VGND.n1358 VGND 0.0213333
R7285 VGND VGND.n3024 0.0193356
R7286 VGND.n33 VGND 0.0161667
R7287 VGND.n331 VGND 0.00980851
R7288 VGND.n2936 VGND 0.00980851
R7289 VGND.n2793 VGND 0.00980851
R7290 VGND.n2785 VGND 0.00980851
R7291 VGND VGND.n288 0.00980851
R7292 VGND.n2758 VGND 0.00980851
R7293 VGND.n2745 VGND 0.00980851
R7294 VGND.n2720 VGND 0.00980851
R7295 VGND.n2712 VGND 0.00980851
R7296 VGND.n2674 VGND 0.00980851
R7297 VGND VGND.n350 0.00980851
R7298 VGND VGND.n349 0.00980851
R7299 VGND VGND.n344 0.00980851
R7300 VGND VGND.n343 0.00980851
R7301 VGND VGND.n338 0.00980851
R7302 VGND VGND.n337 0.00980851
R7303 VGND.n2636 VGND 0.00980851
R7304 VGND VGND.n2534 0.00980851
R7305 VGND VGND.n283 0.00980851
R7306 VGND VGND.n282 0.00980851
R7307 VGND.n2546 VGND 0.00980851
R7308 VGND VGND.n412 0.00980851
R7309 VGND VGND.n411 0.00980851
R7310 VGND VGND.n410 0.00980851
R7311 VGND VGND.n409 0.00980851
R7312 VGND VGND.n408 0.00980851
R7313 VGND VGND.n407 0.00980851
R7314 VGND VGND.n406 0.00980851
R7315 VGND VGND.n405 0.00980851
R7316 VGND VGND.n404 0.00980851
R7317 VGND VGND.n403 0.00980851
R7318 VGND VGND.n402 0.00980851
R7319 VGND.n401 VGND 0.00980851
R7320 VGND.n2529 VGND 0.00980851
R7321 VGND VGND.n420 0.00980851
R7322 VGND VGND.n280 0.00980851
R7323 VGND VGND.n279 0.00980851
R7324 VGND.n2509 VGND 0.00980851
R7325 VGND.n2486 VGND 0.00980851
R7326 VGND.n2478 VGND 0.00980851
R7327 VGND.n2460 VGND 0.00980851
R7328 VGND.n2452 VGND 0.00980851
R7329 VGND.n2434 VGND 0.00980851
R7330 VGND.n2426 VGND 0.00980851
R7331 VGND.n2408 VGND 0.00980851
R7332 VGND.n2400 VGND 0.00980851
R7333 VGND.n2382 VGND 0.00980851
R7334 VGND.n2374 VGND 0.00980851
R7335 VGND.n2356 VGND 0.00980851
R7336 VGND.n2817 VGND 0.00980851
R7337 VGND VGND.n273 0.00980851
R7338 VGND.n2807 VGND 0.00980851
R7339 VGND VGND.n277 0.00980851
R7340 VGND.n2504 VGND 0.00980851
R7341 VGND.n2491 VGND 0.00980851
R7342 VGND.n2473 VGND 0.00980851
R7343 VGND.n2465 VGND 0.00980851
R7344 VGND.n2447 VGND 0.00980851
R7345 VGND.n2439 VGND 0.00980851
R7346 VGND.n2421 VGND 0.00980851
R7347 VGND.n2413 VGND 0.00980851
R7348 VGND.n2395 VGND 0.00980851
R7349 VGND.n2387 VGND 0.00980851
R7350 VGND.n2369 VGND 0.00980851
R7351 VGND.n2361 VGND 0.00980851
R7352 VGND.n1989 VGND 0.00980851
R7353 VGND VGND.n271 0.00980851
R7354 VGND VGND.n270 0.00980851
R7355 VGND.n1974 VGND 0.00980851
R7356 VGND.n1971 VGND 0.00980851
R7357 VGND.n1963 VGND 0.00980851
R7358 VGND.n1960 VGND 0.00980851
R7359 VGND.n1952 VGND 0.00980851
R7360 VGND.n1949 VGND 0.00980851
R7361 VGND.n1941 VGND 0.00980851
R7362 VGND.n1938 VGND 0.00980851
R7363 VGND.n1930 VGND 0.00980851
R7364 VGND.n1927 VGND 0.00980851
R7365 VGND.n1919 VGND 0.00980851
R7366 VGND.n1916 VGND 0.00980851
R7367 VGND.n1908 VGND 0.00980851
R7368 VGND.n1996 VGND 0.00980851
R7369 VGND VGND.n1999 0.00980851
R7370 VGND VGND.n268 0.00980851
R7371 VGND VGND.n267 0.00980851
R7372 VGND VGND.n581 0.00980851
R7373 VGND VGND.n580 0.00980851
R7374 VGND VGND.n575 0.00980851
R7375 VGND VGND.n574 0.00980851
R7376 VGND VGND.n569 0.00980851
R7377 VGND VGND.n568 0.00980851
R7378 VGND VGND.n563 0.00980851
R7379 VGND VGND.n562 0.00980851
R7380 VGND VGND.n557 0.00980851
R7381 VGND VGND.n556 0.00980851
R7382 VGND.n2061 VGND 0.00980851
R7383 VGND.n591 VGND 0.00980851
R7384 VGND.n2842 VGND 0.00980851
R7385 VGND VGND.n261 0.00980851
R7386 VGND.n2832 VGND 0.00980851
R7387 VGND VGND.n265 0.00980851
R7388 VGND.n2130 VGND 0.00980851
R7389 VGND VGND.n578 0.00980851
R7390 VGND VGND.n577 0.00980851
R7391 VGND VGND.n572 0.00980851
R7392 VGND VGND.n571 0.00980851
R7393 VGND VGND.n566 0.00980851
R7394 VGND VGND.n565 0.00980851
R7395 VGND VGND.n560 0.00980851
R7396 VGND VGND.n559 0.00980851
R7397 VGND VGND.n554 0.00980851
R7398 VGND VGND.n553 0.00980851
R7399 VGND.n2067 VGND 0.00980851
R7400 VGND.n1829 VGND 0.00980851
R7401 VGND VGND.n259 0.00980851
R7402 VGND VGND.n258 0.00980851
R7403 VGND.n1814 VGND 0.00980851
R7404 VGND.n1811 VGND 0.00980851
R7405 VGND.n1803 VGND 0.00980851
R7406 VGND.n1800 VGND 0.00980851
R7407 VGND.n1792 VGND 0.00980851
R7408 VGND.n1789 VGND 0.00980851
R7409 VGND.n1781 VGND 0.00980851
R7410 VGND.n1778 VGND 0.00980851
R7411 VGND.n1770 VGND 0.00980851
R7412 VGND.n1767 VGND 0.00980851
R7413 VGND.n1759 VGND 0.00980851
R7414 VGND VGND.n2175 0.00980851
R7415 VGND.n548 VGND 0.00980851
R7416 VGND.n1836 VGND 0.00980851
R7417 VGND VGND.n1839 0.00980851
R7418 VGND VGND.n256 0.00980851
R7419 VGND VGND.n255 0.00980851
R7420 VGND.n1851 VGND 0.00980851
R7421 VGND VGND.n662 0.00980851
R7422 VGND VGND.n661 0.00980851
R7423 VGND VGND.n656 0.00980851
R7424 VGND VGND.n655 0.00980851
R7425 VGND VGND.n650 0.00980851
R7426 VGND VGND.n649 0.00980851
R7427 VGND VGND.n644 0.00980851
R7428 VGND VGND.n643 0.00980851
R7429 VGND.n1687 VGND 0.00980851
R7430 VGND.n1684 VGND 0.00980851
R7431 VGND.n629 VGND 0.00980851
R7432 VGND.n2867 VGND 0.00980851
R7433 VGND VGND.n249 0.00980851
R7434 VGND.n2857 VGND 0.00980851
R7435 VGND VGND.n253 0.00980851
R7436 VGND.n730 VGND 0.00980851
R7437 VGND VGND.n664 0.00980851
R7438 VGND VGND.n659 0.00980851
R7439 VGND VGND.n658 0.00980851
R7440 VGND VGND.n653 0.00980851
R7441 VGND VGND.n652 0.00980851
R7442 VGND VGND.n647 0.00980851
R7443 VGND VGND.n646 0.00980851
R7444 VGND VGND.n641 0.00980851
R7445 VGND VGND.n640 0.00980851
R7446 VGND VGND.n634 0.00980851
R7447 VGND.n633 VGND 0.00980851
R7448 VGND VGND.n1655 0.00980851
R7449 VGND VGND.n247 0.00980851
R7450 VGND VGND.n246 0.00980851
R7451 VGND.n1667 VGND 0.00980851
R7452 VGND VGND.n732 0.00980851
R7453 VGND.n859 VGND 0.00980851
R7454 VGND VGND.n817 0.00980851
R7455 VGND VGND.n816 0.00980851
R7456 VGND VGND.n815 0.00980851
R7457 VGND VGND.n814 0.00980851
R7458 VGND VGND.n813 0.00980851
R7459 VGND.n812 VGND 0.00980851
R7460 VGND VGND.n868 0.00980851
R7461 VGND VGND.n637 0.00980851
R7462 VGND VGND.n636 0.00980851
R7463 VGND.n1350 VGND 0.00980851
R7464 VGND.n1650 VGND 0.00980851
R7465 VGND VGND.n741 0.00980851
R7466 VGND VGND.n244 0.00980851
R7467 VGND VGND.n243 0.00980851
R7468 VGND.n1630 VGND 0.00980851
R7469 VGND VGND.n742 0.00980851
R7470 VGND.n1558 VGND 0.00980851
R7471 VGND VGND.n758 0.00980851
R7472 VGND.n1540 VGND 0.00980851
R7473 VGND.n1522 VGND 0.00980851
R7474 VGND.n1514 VGND 0.00980851
R7475 VGND.n1496 VGND 0.00980851
R7476 VGND.n1488 VGND 0.00980851
R7477 VGND.n1401 VGND 0.00980851
R7478 VGND VGND.n802 0.00980851
R7479 VGND.n801 VGND 0.00980851
R7480 VGND.n2892 VGND 0.00980851
R7481 VGND VGND.n236 0.00980851
R7482 VGND.n2882 VGND 0.00980851
R7483 VGND VGND.n240 0.00980851
R7484 VGND VGND.n745 0.00980851
R7485 VGND VGND.n744 0.00980851
R7486 VGND.n1587 VGND 0.00980851
R7487 VGND.n1564 VGND 0.00980851
R7488 VGND.n1535 VGND 0.00980851
R7489 VGND.n1527 VGND 0.00980851
R7490 VGND.n1509 VGND 0.00980851
R7491 VGND.n1501 VGND 0.00980851
R7492 VGND.n1483 VGND 0.00980851
R7493 VGND.n1475 VGND 0.00980851
R7494 VGND.n1416 VGND 0.00980851
R7495 VGND.n1408 VGND 0.00980851
R7496 VGND VGND.n1607 0.00980851
R7497 VGND VGND.n232 0.00980851
R7498 VGND VGND.n231 0.00980851
R7499 VGND.n1619 VGND 0.00980851
R7500 VGND VGND.n747 0.00980851
R7501 VGND.n1593 VGND 0.00980851
R7502 VGND VGND.n751 0.00980851
R7503 VGND.n1464 VGND 0.00980851
R7504 VGND VGND.n788 0.00980851
R7505 VGND VGND.n787 0.00980851
R7506 VGND VGND.n786 0.00980851
R7507 VGND VGND.n785 0.00980851
R7508 VGND VGND.n784 0.00980851
R7509 VGND VGND.n783 0.00980851
R7510 VGND.n1421 VGND 0.00980851
R7511 VGND.n1343 VGND 0.00980851
R7512 VGND.n2912 VGND 0.00980851
R7513 VGND VGND.n228 0.00980851
R7514 VGND.n2902 VGND 0.00980851
R7515 VGND.n1063 VGND 0.00980851
R7516 VGND VGND.n1046 0.00980851
R7517 VGND.n1045 VGND 0.00980851
R7518 VGND VGND.n1068 0.00980851
R7519 VGND VGND.n912 0.00980851
R7520 VGND VGND.n911 0.00980851
R7521 VGND VGND.n906 0.00980851
R7522 VGND VGND.n905 0.00980851
R7523 VGND VGND.n900 0.00980851
R7524 VGND VGND.n899 0.00980851
R7525 VGND.n1100 VGND 0.00980851
R7526 VGND VGND.n1026 0.00980851
R7527 VGND.n1025 VGND 0.00980851
R7528 VGND.n1165 VGND 0.00980851
R7529 VGND.n1170 VGND 0.00980851
R7530 VGND VGND.n1011 0.00980851
R7531 VGND.n1183 VGND 0.00980851
R7532 VGND.n1191 VGND 0.00980851
R7533 VGND.n1202 VGND 0.00980851
R7534 VGND VGND.n1003 0.00980851
R7535 VGND.n1215 VGND 0.00980851
R7536 VGND.n1249 VGND 0.00980851
R7537 VGND.n1223 VGND 0.00980851
R7538 VGND VGND.n1242 0.00980851
R7539 VGND.n1228 VGND 0.00980851
R7540 VGND VGND.n1235 0.00980851
R7541 VGND.n1272 VGND 0.00980851
R7542 VGND VGND.n997 0.00980851
R7543 VGND.n1282 VGND 0.00980851
R7544 VGND.n2917 VGND 0.00980851
R7545 VGND.n992 VGND 0.00980851
R7546 VGND VGND.n925 0.00980851
R7547 VGND VGND.n924 0.00980851
R7548 VGND VGND.n920 0.00980851
R7549 VGND VGND.n919 0.00980851
R7550 VGND VGND.n915 0.00980851
R7551 VGND VGND.n914 0.00980851
R7552 VGND VGND.n909 0.00980851
R7553 VGND VGND.n908 0.00980851
R7554 VGND VGND.n903 0.00980851
R7555 VGND VGND.n902 0.00980851
R7556 VGND VGND.n897 0.00980851
R7557 VGND.n896 VGND 0.00980851
R7558 VGND VGND.n1331 0.00980851
R7559 VGND.n888 VGND 0.00980851
R7560 VGND.n2698 VGND.n2697 0.00182979
R7561 VGND.n358 VGND.n357 0.00182979
R7562 VGND.n365 VGND.n364 0.00182979
R7563 VGND.n367 VGND.n354 0.00182979
R7564 VGND.n376 VGND.n375 0.00182979
R7565 VGND.n378 VGND.n353 0.00182979
R7566 VGND.n389 VGND.n386 0.00182979
R7567 VGND.n2707 VGND.n325 0.00182979
R7568 VGND.n2725 VGND.n314 0.00182979
R7569 VGND.n2740 VGND.n309 0.00182979
R7570 VGND.n311 VGND.n300 0.00182979
R7571 VGND.n2734 VGND.n2733 0.00182979
R7572 VGND.n2778 VGND.n293 0.00182979
R7573 VGND.n2772 VGND.n296 0.00182979
R7574 VGND.n2942 VGND.n203 0.00182979
R7575 XThR.Tn[2].n2 XThR.Tn[2].n1 332.332
R7576 XThR.Tn[2].n2 XThR.Tn[2].n0 296.493
R7577 XThR.Tn[2] XThR.Tn[2].n82 161.363
R7578 XThR.Tn[2] XThR.Tn[2].n77 161.363
R7579 XThR.Tn[2] XThR.Tn[2].n72 161.363
R7580 XThR.Tn[2] XThR.Tn[2].n67 161.363
R7581 XThR.Tn[2] XThR.Tn[2].n62 161.363
R7582 XThR.Tn[2] XThR.Tn[2].n57 161.363
R7583 XThR.Tn[2] XThR.Tn[2].n52 161.363
R7584 XThR.Tn[2] XThR.Tn[2].n47 161.363
R7585 XThR.Tn[2] XThR.Tn[2].n42 161.363
R7586 XThR.Tn[2] XThR.Tn[2].n37 161.363
R7587 XThR.Tn[2] XThR.Tn[2].n32 161.363
R7588 XThR.Tn[2] XThR.Tn[2].n27 161.363
R7589 XThR.Tn[2] XThR.Tn[2].n22 161.363
R7590 XThR.Tn[2] XThR.Tn[2].n17 161.363
R7591 XThR.Tn[2] XThR.Tn[2].n12 161.363
R7592 XThR.Tn[2] XThR.Tn[2].n10 161.363
R7593 XThR.Tn[2].n84 XThR.Tn[2].n83 161.3
R7594 XThR.Tn[2].n79 XThR.Tn[2].n78 161.3
R7595 XThR.Tn[2].n74 XThR.Tn[2].n73 161.3
R7596 XThR.Tn[2].n69 XThR.Tn[2].n68 161.3
R7597 XThR.Tn[2].n64 XThR.Tn[2].n63 161.3
R7598 XThR.Tn[2].n59 XThR.Tn[2].n58 161.3
R7599 XThR.Tn[2].n54 XThR.Tn[2].n53 161.3
R7600 XThR.Tn[2].n49 XThR.Tn[2].n48 161.3
R7601 XThR.Tn[2].n44 XThR.Tn[2].n43 161.3
R7602 XThR.Tn[2].n39 XThR.Tn[2].n38 161.3
R7603 XThR.Tn[2].n34 XThR.Tn[2].n33 161.3
R7604 XThR.Tn[2].n29 XThR.Tn[2].n28 161.3
R7605 XThR.Tn[2].n24 XThR.Tn[2].n23 161.3
R7606 XThR.Tn[2].n19 XThR.Tn[2].n18 161.3
R7607 XThR.Tn[2].n14 XThR.Tn[2].n13 161.3
R7608 XThR.Tn[2].n82 XThR.Tn[2].t65 161.106
R7609 XThR.Tn[2].n77 XThR.Tn[2].t72 161.106
R7610 XThR.Tn[2].n72 XThR.Tn[2].t51 161.106
R7611 XThR.Tn[2].n67 XThR.Tn[2].t36 161.106
R7612 XThR.Tn[2].n62 XThR.Tn[2].t64 161.106
R7613 XThR.Tn[2].n57 XThR.Tn[2].t26 161.106
R7614 XThR.Tn[2].n52 XThR.Tn[2].t69 161.106
R7615 XThR.Tn[2].n47 XThR.Tn[2].t49 161.106
R7616 XThR.Tn[2].n42 XThR.Tn[2].t35 161.106
R7617 XThR.Tn[2].n37 XThR.Tn[2].t41 161.106
R7618 XThR.Tn[2].n32 XThR.Tn[2].t25 161.106
R7619 XThR.Tn[2].n27 XThR.Tn[2].t50 161.106
R7620 XThR.Tn[2].n22 XThR.Tn[2].t23 161.106
R7621 XThR.Tn[2].n17 XThR.Tn[2].t67 161.106
R7622 XThR.Tn[2].n12 XThR.Tn[2].t31 161.106
R7623 XThR.Tn[2].n10 XThR.Tn[2].t14 161.106
R7624 XThR.Tn[2].n83 XThR.Tn[2].t38 159.978
R7625 XThR.Tn[2].n78 XThR.Tn[2].t46 159.978
R7626 XThR.Tn[2].n73 XThR.Tn[2].t29 159.978
R7627 XThR.Tn[2].n68 XThR.Tn[2].t13 159.978
R7628 XThR.Tn[2].n63 XThR.Tn[2].t37 159.978
R7629 XThR.Tn[2].n58 XThR.Tn[2].t63 159.978
R7630 XThR.Tn[2].n53 XThR.Tn[2].t45 159.978
R7631 XThR.Tn[2].n48 XThR.Tn[2].t27 159.978
R7632 XThR.Tn[2].n43 XThR.Tn[2].t12 159.978
R7633 XThR.Tn[2].n38 XThR.Tn[2].t20 159.978
R7634 XThR.Tn[2].n33 XThR.Tn[2].t62 159.978
R7635 XThR.Tn[2].n28 XThR.Tn[2].t28 159.978
R7636 XThR.Tn[2].n23 XThR.Tn[2].t60 159.978
R7637 XThR.Tn[2].n18 XThR.Tn[2].t43 159.978
R7638 XThR.Tn[2].n13 XThR.Tn[2].t66 159.978
R7639 XThR.Tn[2].n82 XThR.Tn[2].t53 145.038
R7640 XThR.Tn[2].n77 XThR.Tn[2].t19 145.038
R7641 XThR.Tn[2].n72 XThR.Tn[2].t59 145.038
R7642 XThR.Tn[2].n67 XThR.Tn[2].t42 145.038
R7643 XThR.Tn[2].n62 XThR.Tn[2].t73 145.038
R7644 XThR.Tn[2].n57 XThR.Tn[2].t52 145.038
R7645 XThR.Tn[2].n52 XThR.Tn[2].t61 145.038
R7646 XThR.Tn[2].n47 XThR.Tn[2].t44 145.038
R7647 XThR.Tn[2].n42 XThR.Tn[2].t39 145.038
R7648 XThR.Tn[2].n37 XThR.Tn[2].t70 145.038
R7649 XThR.Tn[2].n32 XThR.Tn[2].t34 145.038
R7650 XThR.Tn[2].n27 XThR.Tn[2].t58 145.038
R7651 XThR.Tn[2].n22 XThR.Tn[2].t32 145.038
R7652 XThR.Tn[2].n17 XThR.Tn[2].t15 145.038
R7653 XThR.Tn[2].n12 XThR.Tn[2].t40 145.038
R7654 XThR.Tn[2].n10 XThR.Tn[2].t21 145.038
R7655 XThR.Tn[2].n83 XThR.Tn[2].t71 143.911
R7656 XThR.Tn[2].n78 XThR.Tn[2].t33 143.911
R7657 XThR.Tn[2].n73 XThR.Tn[2].t17 143.911
R7658 XThR.Tn[2].n68 XThR.Tn[2].t56 143.911
R7659 XThR.Tn[2].n63 XThR.Tn[2].t24 143.911
R7660 XThR.Tn[2].n58 XThR.Tn[2].t68 143.911
R7661 XThR.Tn[2].n53 XThR.Tn[2].t18 143.911
R7662 XThR.Tn[2].n48 XThR.Tn[2].t57 143.911
R7663 XThR.Tn[2].n43 XThR.Tn[2].t54 143.911
R7664 XThR.Tn[2].n38 XThR.Tn[2].t22 143.911
R7665 XThR.Tn[2].n33 XThR.Tn[2].t48 143.911
R7666 XThR.Tn[2].n28 XThR.Tn[2].t16 143.911
R7667 XThR.Tn[2].n23 XThR.Tn[2].t47 143.911
R7668 XThR.Tn[2].n18 XThR.Tn[2].t30 143.911
R7669 XThR.Tn[2].n13 XThR.Tn[2].t55 143.911
R7670 XThR.Tn[2].n7 XThR.Tn[2].n5 135.249
R7671 XThR.Tn[2].n9 XThR.Tn[2].n3 98.982
R7672 XThR.Tn[2].n8 XThR.Tn[2].n4 98.982
R7673 XThR.Tn[2].n7 XThR.Tn[2].n6 98.982
R7674 XThR.Tn[2].n9 XThR.Tn[2].n8 36.2672
R7675 XThR.Tn[2].n8 XThR.Tn[2].n7 36.2672
R7676 XThR.Tn[2].n88 XThR.Tn[2].n9 32.6405
R7677 XThR.Tn[2].n1 XThR.Tn[2].t6 26.5955
R7678 XThR.Tn[2].n1 XThR.Tn[2].t5 26.5955
R7679 XThR.Tn[2].n0 XThR.Tn[2].t7 26.5955
R7680 XThR.Tn[2].n0 XThR.Tn[2].t4 26.5955
R7681 XThR.Tn[2].n3 XThR.Tn[2].t10 24.9236
R7682 XThR.Tn[2].n3 XThR.Tn[2].t11 24.9236
R7683 XThR.Tn[2].n4 XThR.Tn[2].t9 24.9236
R7684 XThR.Tn[2].n4 XThR.Tn[2].t8 24.9236
R7685 XThR.Tn[2].n5 XThR.Tn[2].t1 24.9236
R7686 XThR.Tn[2].n5 XThR.Tn[2].t2 24.9236
R7687 XThR.Tn[2].n6 XThR.Tn[2].t0 24.9236
R7688 XThR.Tn[2].n6 XThR.Tn[2].t3 24.9236
R7689 XThR.Tn[2] XThR.Tn[2].n2 23.3605
R7690 XThR.Tn[2] XThR.Tn[2].n88 6.7205
R7691 XThR.Tn[2].n88 XThR.Tn[2] 6.30883
R7692 XThR.Tn[2] XThR.Tn[2].n11 5.34038
R7693 XThR.Tn[2].n16 XThR.Tn[2].n15 4.5005
R7694 XThR.Tn[2].n21 XThR.Tn[2].n20 4.5005
R7695 XThR.Tn[2].n26 XThR.Tn[2].n25 4.5005
R7696 XThR.Tn[2].n31 XThR.Tn[2].n30 4.5005
R7697 XThR.Tn[2].n36 XThR.Tn[2].n35 4.5005
R7698 XThR.Tn[2].n41 XThR.Tn[2].n40 4.5005
R7699 XThR.Tn[2].n46 XThR.Tn[2].n45 4.5005
R7700 XThR.Tn[2].n51 XThR.Tn[2].n50 4.5005
R7701 XThR.Tn[2].n56 XThR.Tn[2].n55 4.5005
R7702 XThR.Tn[2].n61 XThR.Tn[2].n60 4.5005
R7703 XThR.Tn[2].n66 XThR.Tn[2].n65 4.5005
R7704 XThR.Tn[2].n71 XThR.Tn[2].n70 4.5005
R7705 XThR.Tn[2].n76 XThR.Tn[2].n75 4.5005
R7706 XThR.Tn[2].n81 XThR.Tn[2].n80 4.5005
R7707 XThR.Tn[2].n86 XThR.Tn[2].n85 4.5005
R7708 XThR.Tn[2].n87 XThR.Tn[2] 3.70586
R7709 XThR.Tn[2].n16 XThR.Tn[2] 2.52282
R7710 XThR.Tn[2].n21 XThR.Tn[2] 2.52282
R7711 XThR.Tn[2].n26 XThR.Tn[2] 2.52282
R7712 XThR.Tn[2].n31 XThR.Tn[2] 2.52282
R7713 XThR.Tn[2].n36 XThR.Tn[2] 2.52282
R7714 XThR.Tn[2].n41 XThR.Tn[2] 2.52282
R7715 XThR.Tn[2].n46 XThR.Tn[2] 2.52282
R7716 XThR.Tn[2].n51 XThR.Tn[2] 2.52282
R7717 XThR.Tn[2].n56 XThR.Tn[2] 2.52282
R7718 XThR.Tn[2].n61 XThR.Tn[2] 2.52282
R7719 XThR.Tn[2].n66 XThR.Tn[2] 2.52282
R7720 XThR.Tn[2].n71 XThR.Tn[2] 2.52282
R7721 XThR.Tn[2].n76 XThR.Tn[2] 2.52282
R7722 XThR.Tn[2].n81 XThR.Tn[2] 2.52282
R7723 XThR.Tn[2].n86 XThR.Tn[2] 2.52282
R7724 XThR.Tn[2].n84 XThR.Tn[2] 1.08677
R7725 XThR.Tn[2].n79 XThR.Tn[2] 1.08677
R7726 XThR.Tn[2].n74 XThR.Tn[2] 1.08677
R7727 XThR.Tn[2].n69 XThR.Tn[2] 1.08677
R7728 XThR.Tn[2].n64 XThR.Tn[2] 1.08677
R7729 XThR.Tn[2].n59 XThR.Tn[2] 1.08677
R7730 XThR.Tn[2].n54 XThR.Tn[2] 1.08677
R7731 XThR.Tn[2].n49 XThR.Tn[2] 1.08677
R7732 XThR.Tn[2].n44 XThR.Tn[2] 1.08677
R7733 XThR.Tn[2].n39 XThR.Tn[2] 1.08677
R7734 XThR.Tn[2].n34 XThR.Tn[2] 1.08677
R7735 XThR.Tn[2].n29 XThR.Tn[2] 1.08677
R7736 XThR.Tn[2].n24 XThR.Tn[2] 1.08677
R7737 XThR.Tn[2].n19 XThR.Tn[2] 1.08677
R7738 XThR.Tn[2].n14 XThR.Tn[2] 1.08677
R7739 XThR.Tn[2] XThR.Tn[2].n16 0.839786
R7740 XThR.Tn[2] XThR.Tn[2].n21 0.839786
R7741 XThR.Tn[2] XThR.Tn[2].n26 0.839786
R7742 XThR.Tn[2] XThR.Tn[2].n31 0.839786
R7743 XThR.Tn[2] XThR.Tn[2].n36 0.839786
R7744 XThR.Tn[2] XThR.Tn[2].n41 0.839786
R7745 XThR.Tn[2] XThR.Tn[2].n46 0.839786
R7746 XThR.Tn[2] XThR.Tn[2].n51 0.839786
R7747 XThR.Tn[2] XThR.Tn[2].n56 0.839786
R7748 XThR.Tn[2] XThR.Tn[2].n61 0.839786
R7749 XThR.Tn[2] XThR.Tn[2].n66 0.839786
R7750 XThR.Tn[2] XThR.Tn[2].n71 0.839786
R7751 XThR.Tn[2] XThR.Tn[2].n76 0.839786
R7752 XThR.Tn[2] XThR.Tn[2].n81 0.839786
R7753 XThR.Tn[2] XThR.Tn[2].n86 0.839786
R7754 XThR.Tn[2].n11 XThR.Tn[2] 0.499542
R7755 XThR.Tn[2].n85 XThR.Tn[2] 0.063
R7756 XThR.Tn[2].n80 XThR.Tn[2] 0.063
R7757 XThR.Tn[2].n75 XThR.Tn[2] 0.063
R7758 XThR.Tn[2].n70 XThR.Tn[2] 0.063
R7759 XThR.Tn[2].n65 XThR.Tn[2] 0.063
R7760 XThR.Tn[2].n60 XThR.Tn[2] 0.063
R7761 XThR.Tn[2].n55 XThR.Tn[2] 0.063
R7762 XThR.Tn[2].n50 XThR.Tn[2] 0.063
R7763 XThR.Tn[2].n45 XThR.Tn[2] 0.063
R7764 XThR.Tn[2].n40 XThR.Tn[2] 0.063
R7765 XThR.Tn[2].n35 XThR.Tn[2] 0.063
R7766 XThR.Tn[2].n30 XThR.Tn[2] 0.063
R7767 XThR.Tn[2].n25 XThR.Tn[2] 0.063
R7768 XThR.Tn[2].n20 XThR.Tn[2] 0.063
R7769 XThR.Tn[2].n15 XThR.Tn[2] 0.063
R7770 XThR.Tn[2].n87 XThR.Tn[2] 0.0540714
R7771 XThR.Tn[2] XThR.Tn[2].n87 0.038
R7772 XThR.Tn[2].n11 XThR.Tn[2] 0.0143889
R7773 XThR.Tn[2].n85 XThR.Tn[2].n84 0.00771154
R7774 XThR.Tn[2].n80 XThR.Tn[2].n79 0.00771154
R7775 XThR.Tn[2].n75 XThR.Tn[2].n74 0.00771154
R7776 XThR.Tn[2].n70 XThR.Tn[2].n69 0.00771154
R7777 XThR.Tn[2].n65 XThR.Tn[2].n64 0.00771154
R7778 XThR.Tn[2].n60 XThR.Tn[2].n59 0.00771154
R7779 XThR.Tn[2].n55 XThR.Tn[2].n54 0.00771154
R7780 XThR.Tn[2].n50 XThR.Tn[2].n49 0.00771154
R7781 XThR.Tn[2].n45 XThR.Tn[2].n44 0.00771154
R7782 XThR.Tn[2].n40 XThR.Tn[2].n39 0.00771154
R7783 XThR.Tn[2].n35 XThR.Tn[2].n34 0.00771154
R7784 XThR.Tn[2].n30 XThR.Tn[2].n29 0.00771154
R7785 XThR.Tn[2].n25 XThR.Tn[2].n24 0.00771154
R7786 XThR.Tn[2].n20 XThR.Tn[2].n19 0.00771154
R7787 XThR.Tn[2].n15 XThR.Tn[2].n14 0.00771154
R7788 VPWR.n2837 VPWR.n2823 2618.82
R7789 VPWR.n2835 VPWR.n2829 2618.82
R7790 VPWR.n2853 VPWR.n2823 1916.47
R7791 VPWR.n2828 VPWR.n2827 1916.47
R7792 VPWR.n2827 VPWR.n2821 1916.47
R7793 VPWR.n2829 VPWR.n2822 1916.47
R7794 VPWR.n2852 VPWR.n2824 1912.94
R7795 VPWR.n2849 VPWR.n2843 1560
R7796 VPWR.n2850 VPWR.n2824 1408.24
R7797 VPWR.n2853 VPWR.n2852 1210.59
R7798 VPWR.n2851 VPWR.n2821 1210.59
R7799 VPWR.n2380 VPWR.t713 1005.7
R7800 VPWR.t931 VPWR.n485 1005.7
R7801 VPWR.t780 VPWR.n2210 1005.7
R7802 VPWR.n639 VPWR.t888 1005.7
R7803 VPWR.n2184 VPWR.t614 1005.7
R7804 VPWR.t721 VPWR.n677 1005.7
R7805 VPWR.t681 VPWR.n2014 1005.7
R7806 VPWR.n831 VPWR.t786 1005.7
R7807 VPWR.n1988 VPWR.t609 1005.7
R7808 VPWR.t793 VPWR.n869 1005.7
R7809 VPWR.n447 VPWR.t601 1005.7
R7810 VPWR.t901 VPWR.n1818 1005.7
R7811 VPWR.t880 VPWR.n2406 1005.7
R7812 VPWR.n1023 VPWR.t753 1005.7
R7813 VPWR.t923 VPWR.n293 1005.7
R7814 VPWR.n1792 VPWR.t864 1005.7
R7815 VPWR.n2591 VPWR.t815 1005.7
R7816 VPWR.n1062 VPWR.t699 1005.7
R7817 VPWR.t85 VPWR.n2309 983.14
R7818 VPWR.n2310 VPWR.t128 983.14
R7819 VPWR.t1189 VPWR.n2319 983.14
R7820 VPWR.n2320 VPWR.t146 983.14
R7821 VPWR.t1579 VPWR.n2329 983.14
R7822 VPWR.n2330 VPWR.t1289 983.14
R7823 VPWR.t220 VPWR.n2339 983.14
R7824 VPWR.n2340 VPWR.t1384 983.14
R7825 VPWR.t561 VPWR.n2349 983.14
R7826 VPWR.n2350 VPWR.t447 983.14
R7827 VPWR.t1735 VPWR.n2359 983.14
R7828 VPWR.n2360 VPWR.t1899 983.14
R7829 VPWR.t182 VPWR.n2369 983.14
R7830 VPWR.n2370 VPWR.t1206 983.14
R7831 VPWR.t4 VPWR.n2379 983.14
R7832 VPWR.n542 VPWR.t1619 983.14
R7833 VPWR.n541 VPWR.t1712 983.14
R7834 VPWR.n537 VPWR.t1165 983.14
R7835 VPWR.n533 VPWR.t1044 983.14
R7836 VPWR.n529 VPWR.t1526 983.14
R7837 VPWR.n525 VPWR.t1480 983.14
R7838 VPWR.n521 VPWR.t1859 983.14
R7839 VPWR.n517 VPWR.t499 983.14
R7840 VPWR.n513 VPWR.t1038 983.14
R7841 VPWR.n509 VPWR.t380 983.14
R7842 VPWR.n505 VPWR.t1512 983.14
R7843 VPWR.n501 VPWR.t35 983.14
R7844 VPWR.n497 VPWR.t282 983.14
R7845 VPWR.n493 VPWR.t527 983.14
R7846 VPWR.n489 VPWR.t192 983.14
R7847 VPWR.n2281 VPWR.t557 983.14
R7848 VPWR.n2280 VPWR.t1647 983.14
R7849 VPWR.n2271 VPWR.t1143 983.14
R7850 VPWR.n2270 VPWR.t1068 983.14
R7851 VPWR.n2261 VPWR.t1554 983.14
R7852 VPWR.n2260 VPWR.t1496 983.14
R7853 VPWR.n2251 VPWR.t1697 983.14
R7854 VPWR.n2250 VPWR.t250 983.14
R7855 VPWR.n2241 VPWR.t522 983.14
R7856 VPWR.n2240 VPWR.t435 983.14
R7857 VPWR.n2231 VPWR.t475 983.14
R7858 VPWR.n2230 VPWR.t1441 983.14
R7859 VPWR.n2221 VPWR.t166 983.14
R7860 VPWR.n2220 VPWR.t1568 983.14
R7861 VPWR.n2211 VPWR.t1635 983.14
R7862 VPWR.t983 VPWR.n582 983.14
R7863 VPWR.t1546 VPWR.n586 983.14
R7864 VPWR.t1157 VPWR.n590 983.14
R7865 VPWR.t1050 VPWR.n594 983.14
R7866 VPWR.t113 VPWR.n598 983.14
R7867 VPWR.t1259 VPWR.n602 983.14
R7868 VPWR.t1869 VPWR.n606 983.14
R7869 VPWR.t276 VPWR.n610 983.14
R7870 VPWR.t320 VPWR.n614 983.14
R7871 VPWR.t401 VPWR.n618 983.14
R7872 VPWR.t1749 VPWR.n622 983.14
R7873 VPWR.t962 VPWR.n626 983.14
R7874 VPWR.t290 VPWR.n630 983.14
R7875 VPWR.t1420 VPWR.n634 983.14
R7876 VPWR.t389 VPWR.n638 983.14
R7877 VPWR.t308 VPWR.n2113 983.14
R7878 VPWR.n2114 VPWR.t1607 983.14
R7879 VPWR.t1179 VPWR.n2123 983.14
R7880 VPWR.n2124 VPWR.t1027 983.14
R7881 VPWR.t1520 VPWR.n2133 983.14
R7882 VPWR.n2134 VPWR.t1271 983.14
R7883 VPWR.t230 VPWR.n2143 983.14
R7884 VPWR.n2144 VPWR.t1405 983.14
R7885 VPWR.t130 VPWR.n2153 983.14
R7886 VPWR.n2154 VPWR.t356 983.14
R7887 VPWR.t1118 VPWR.n2163 983.14
R7888 VPWR.n2164 VPWR.t1536 983.14
R7889 VPWR.t49 VPWR.n2173 983.14
R7890 VPWR.n2174 VPWR.t485 983.14
R7891 VPWR.t206 VPWR.n2183 983.14
R7892 VPWR.n734 VPWR.t1109 983.14
R7893 VPWR.n733 VPWR.t126 983.14
R7894 VPWR.n729 VPWR.t1191 983.14
R7895 VPWR.n725 VPWR.t144 983.14
R7896 VPWR.n721 VPWR.t1577 983.14
R7897 VPWR.n717 VPWR.t1287 983.14
R7898 VPWR.n713 VPWR.t952 983.14
R7899 VPWR.n709 VPWR.t958 983.14
R7900 VPWR.n705 VPWR.t559 983.14
R7901 VPWR.n701 VPWR.t445 983.14
R7902 VPWR.n697 VPWR.t1733 983.14
R7903 VPWR.n693 VPWR.t1897 983.14
R7904 VPWR.n689 VPWR.t180 983.14
R7905 VPWR.n685 VPWR.t1204 983.14
R7906 VPWR.n681 VPWR.t1645 983.14
R7907 VPWR.n2085 VPWR.t459 983.14
R7908 VPWR.n2084 VPWR.t510 983.14
R7909 VPWR.n2075 VPWR.t1185 983.14
R7910 VPWR.n2074 VPWR.t148 983.14
R7911 VPWR.n2065 VPWR.t1306 983.14
R7912 VPWR.n2064 VPWR.t1343 983.14
R7913 VPWR.n2055 VPWR.t226 983.14
R7914 VPWR.n2054 VPWR.t1386 983.14
R7915 VPWR.n2045 VPWR.t1221 983.14
R7916 VPWR.n2044 VPWR.t350 983.14
R7917 VPWR.n2035 VPWR.t1848 983.14
R7918 VPWR.n2034 VPWR.t1884 983.14
R7919 VPWR.n2025 VPWR.t39 983.14
R7920 VPWR.n2024 VPWR.t1585 983.14
R7921 VPWR.n2015 VPWR.t6 983.14
R7922 VPWR.t555 VPWR.n774 983.14
R7923 VPWR.t516 VPWR.n778 983.14
R7924 VPWR.t1145 VPWR.n782 983.14
R7925 VPWR.t1064 VPWR.n786 983.14
R7926 VPWR.t1552 VPWR.n790 983.14
R7927 VPWR.t1494 VPWR.n794 983.14
R7928 VPWR.t1695 VPWR.n798 983.14
R7929 VPWR.t246 VPWR.n802 983.14
R7930 VPWR.t520 VPWR.n806 983.14
R7931 VPWR.t374 VPWR.n810 983.14
R7932 VPWR.t473 VPWR.n814 983.14
R7933 VPWR.t1359 VPWR.n818 983.14
R7934 VPWR.t162 VPWR.n822 983.14
R7935 VPWR.t1566 VPWR.n826 983.14
R7936 VPWR.t1631 VPWR.n830 983.14
R7937 VPWR.t310 VPWR.n1917 983.14
R7938 VPWR.n1918 VPWR.t1609 983.14
R7939 VPWR.t1177 VPWR.n1927 983.14
R7940 VPWR.n1928 VPWR.t1060 983.14
R7941 VPWR.t1522 VPWR.n1937 983.14
R7942 VPWR.n1938 VPWR.t1273 983.14
R7943 VPWR.t232 VPWR.n1947 983.14
R7944 VPWR.n1948 VPWR.t240 983.14
R7945 VPWR.t132 VPWR.n1957 983.14
R7946 VPWR.n1958 VPWR.t358 983.14
R7947 VPWR.t1120 VPWR.n1967 983.14
R7948 VPWR.n1968 VPWR.t1538 983.14
R7949 VPWR.t51 VPWR.n1977 983.14
R7950 VPWR.n1978 VPWR.t487 983.14
R7951 VPWR.t208 VPWR.n1987 983.14
R7952 VPWR.n926 VPWR.t553 983.14
R7953 VPWR.n925 VPWR.t514 983.14
R7954 VPWR.n921 VPWR.t1147 983.14
R7955 VPWR.n917 VPWR.t1062 983.14
R7956 VPWR.n913 VPWR.t1699 983.14
R7957 VPWR.n909 VPWR.t1492 983.14
R7958 VPWR.n905 VPWR.t1693 983.14
R7959 VPWR.n901 VPWR.t268 983.14
R7960 VPWR.n897 VPWR.t518 983.14
R7961 VPWR.n893 VPWR.t372 983.14
R7962 VPWR.n889 VPWR.t471 983.14
R7963 VPWR.n885 VPWR.t1357 983.14
R7964 VPWR.n881 VPWR.t158 983.14
R7965 VPWR.n877 VPWR.t1564 983.14
R7966 VPWR.n873 VPWR.t1629 983.14
R7967 VPWR.t312 VPWR.n390 983.14
R7968 VPWR.t1611 VPWR.n394 983.14
R7969 VPWR.t1173 VPWR.n398 983.14
R7970 VPWR.t1410 VPWR.n402 983.14
R7971 VPWR.t1524 VPWR.n406 983.14
R7972 VPWR.t1275 VPWR.n410 983.14
R7973 VPWR.t234 VPWR.n414 983.14
R7974 VPWR.t242 VPWR.n418 983.14
R7975 VPWR.t134 VPWR.n422 983.14
R7976 VPWR.t360 VPWR.n426 983.14
R7977 VPWR.t1122 VPWR.n430 983.14
R7978 VPWR.t1540 VPWR.n434 983.14
R7979 VPWR.t53 VPWR.n438 983.14
R7980 VPWR.t489 VPWR.n442 983.14
R7981 VPWR.t186 VPWR.n446 983.14
R7982 VPWR.n1889 VPWR.t16 983.14
R7983 VPWR.n1888 VPWR.t1542 983.14
R7984 VPWR.n1879 VPWR.t1159 983.14
R7985 VPWR.n1878 VPWR.t1048 983.14
R7986 VPWR.n1869 VPWR.t109 983.14
R7987 VPWR.n1868 VPWR.t1486 983.14
R7988 VPWR.n1859 VPWR.t1865 983.14
R7989 VPWR.n1858 VPWR.t274 983.14
R7990 VPWR.n1849 VPWR.t316 983.14
R7991 VPWR.n1848 VPWR.t384 983.14
R7992 VPWR.n1839 VPWR.t1745 983.14
R7993 VPWR.n1838 VPWR.t960 983.14
R7994 VPWR.n1829 VPWR.t288 983.14
R7995 VPWR.n1828 VPWR.t1418 983.14
R7996 VPWR.n1819 VPWR.t196 983.14
R7997 VPWR.n2477 VPWR.t985 983.14
R7998 VPWR.n2476 VPWR.t1548 983.14
R7999 VPWR.n2467 VPWR.t1155 983.14
R8000 VPWR.n2466 VPWR.t1054 983.14
R8001 VPWR.n2457 VPWR.t115 983.14
R8002 VPWR.n2456 VPWR.t1261 983.14
R8003 VPWR.n2447 VPWR.t1871 983.14
R8004 VPWR.n2446 VPWR.t278 983.14
R8005 VPWR.n2437 VPWR.t322 983.14
R8006 VPWR.n2436 VPWR.t403 983.14
R8007 VPWR.n2427 VPWR.t1751 983.14
R8008 VPWR.n2426 VPWR.t964 983.14
R8009 VPWR.n2417 VPWR.t292 983.14
R8010 VPWR.n2416 VPWR.t1422 983.14
R8011 VPWR.n2407 VPWR.t393 983.14
R8012 VPWR.t1101 VPWR.n966 983.14
R8013 VPWR.t1653 VPWR.n970 983.14
R8014 VPWR.t1137 VPWR.n974 983.14
R8015 VPWR.t1074 VPWR.n978 983.14
R8016 VPWR.t1560 VPWR.n982 983.14
R8017 VPWR.t1502 VPWR.n986 983.14
R8018 VPWR.t214 VPWR.n990 983.14
R8019 VPWR.t254 VPWR.n994 983.14
R8020 VPWR.t71 VPWR.n998 983.14
R8021 VPWR.t437 VPWR.n1002 983.14
R8022 VPWR.t481 VPWR.n1006 983.14
R8023 VPWR.t1443 VPWR.n1010 983.14
R8024 VPWR.t172 VPWR.n1014 983.14
R8025 VPWR.t103 VPWR.n1018 983.14
R8026 VPWR.t1641 VPWR.n1022 983.14
R8027 VPWR.n350 VPWR.t1621 983.14
R8028 VPWR.n349 VPWR.t1714 983.14
R8029 VPWR.n345 VPWR.t1163 983.14
R8030 VPWR.n341 VPWR.t1046 983.14
R8031 VPWR.n337 VPWR.t1528 983.14
R8032 VPWR.n333 VPWR.t1482 983.14
R8033 VPWR.n329 VPWR.t1861 983.14
R8034 VPWR.n325 VPWR.t272 983.14
R8035 VPWR.n321 VPWR.t1040 983.14
R8036 VPWR.n317 VPWR.t382 983.14
R8037 VPWR.n313 VPWR.t1514 983.14
R8038 VPWR.n309 VPWR.t37 983.14
R8039 VPWR.n305 VPWR.t286 983.14
R8040 VPWR.n301 VPWR.t529 983.14
R8041 VPWR.n297 VPWR.t194 983.14
R8042 VPWR.t834 VPWR.n1468 983.14
R8043 VPWR.t936 VPWR.n1475 983.14
R8044 VPWR.t707 VPWR.n1481 983.14
R8045 VPWR.t809 VPWR.n1492 983.14
R8046 VPWR.n1493 VPWR.t831 983.14
R8047 VPWR.t582 VPWR.n1506 983.14
R8048 VPWR.n1507 VPWR.t704 983.14
R8049 VPWR.t845 VPWR.n1520 983.14
R8050 VPWR.n1521 VPWR.t861 983.14
R8051 VPWR.n1536 VPWR.t604 983.14
R8052 VPWR.n1535 VPWR.t734 983.14
R8053 VPWR.n1761 VPWR.t775 983.14
R8054 VPWR.n1760 VPWR.t598 983.14
R8055 VPWR.n1749 VPWR.t648 983.14
R8056 VPWR.t756 VPWR.n1791 983.14
R8057 VPWR.t762 VPWR.n2506 983.14
R8058 VPWR.n2507 VPWR.t874 983.14
R8059 VPWR.t639 VPWR.n2518 983.14
R8060 VPWR.n2519 VPWR.t750 983.14
R8061 VPWR.t759 VPWR.n2530 983.14
R8062 VPWR.n2531 VPWR.t915 983.14
R8063 VPWR.t636 VPWR.n2542 983.14
R8064 VPWR.n2543 VPWR.t796 983.14
R8065 VPWR.t812 VPWR.n2554 983.14
R8066 VPWR.n2555 VPWR.t942 983.14
R8067 VPWR.t686 VPWR.n2566 983.14
R8068 VPWR.n2567 VPWR.t716 983.14
R8069 VPWR.t566 VPWR.n2578 983.14
R8070 VPWR.n2579 VPWR.t585 983.14
R8071 VPWR.t710 VPWR.n2590 983.14
R8072 VPWR.n1594 VPWR.t645 983.14
R8073 VPWR.n1593 VPWR.t747 983.14
R8074 VPWR.t912 VPWR.n1182 983.14
R8075 VPWR.t630 VPWR.n1185 983.14
R8076 VPWR.n1220 VPWR.t642 983.14
R8077 VPWR.n1219 VPWR.t801 983.14
R8078 VPWR.n1216 VPWR.t909 983.14
R8079 VPWR.n1213 VPWR.t670 983.14
R8080 VPWR.n1205 VPWR.t696 983.14
R8081 VPWR.n1202 VPWR.t823 983.14
R8082 VPWR.n1199 VPWR.t569 983.14
R8083 VPWR.n1191 VPWR.t590 983.14
R8084 VPWR.n1188 VPWR.t828 983.14
R8085 VPWR.n1740 VPWR.t856 983.14
R8086 VPWR.n1739 VPWR.t576 983.14
R8087 VPWR.n1308 VPWR.t1758 877.144
R8088 VPWR.n2723 VPWR.t1807 877.144
R8089 VPWR.n2843 VPWR.n2822 857.648
R8090 VPWR.n1122 VPWR.t878 738.074
R8091 VPWR.n99 VPWR.t618 738.074
R8092 VPWR.n290 VPWR.t1464 738.074
R8093 VPWR.n68 VPWR.t687 738.074
R8094 VPWR.n346 VPWR.t1622 738.074
R8095 VPWR.n98 VPWR.t763 738.074
R8096 VPWR.n963 VPWR.t1450 738.074
R8097 VPWR.n356 VPWR.t1458 738.074
R8098 VPWR.n357 VPWR.t986 738.074
R8099 VPWR.n318 VPWR.t273 738.074
R8100 VPWR.n75 VPWR.t797 738.074
R8101 VPWR.n971 VPWR.t1654 738.074
R8102 VPWR.n369 VPWR.t1872 738.074
R8103 VPWR.n322 VPWR.t1862 738.074
R8104 VPWR.n80 VPWR.t637 738.074
R8105 VPWR.n932 VPWR.t1462 738.074
R8106 VPWR.n933 VPWR.t17 738.074
R8107 VPWR.n936 VPWR.t1543 738.074
R8108 VPWR.n387 VPWR.t1468 738.074
R8109 VPWR.n391 VPWR.t313 738.074
R8110 VPWR.n395 VPWR.t1612 738.074
R8111 VPWR.n365 VPWR.t116 738.074
R8112 VPWR.n330 VPWR.t1529 738.074
R8113 VPWR.n86 VPWR.t760 738.074
R8114 VPWR.n937 VPWR.t1160 738.074
R8115 VPWR.n403 VPWR.t1411 738.074
R8116 VPWR.n364 VPWR.t1055 738.074
R8117 VPWR.n334 VPWR.t1047 738.074
R8118 VPWR.n87 VPWR.t751 738.074
R8119 VPWR.n481 VPWR.t1477 738.074
R8120 VPWR.n480 VPWR.t86 738.074
R8121 VPWR.n477 VPWR.t129 738.074
R8122 VPWR.n476 VPWR.t1190 738.074
R8123 VPWR.n472 VPWR.t1580 738.074
R8124 VPWR.n469 VPWR.t1290 738.074
R8125 VPWR.n468 VPWR.t221 738.074
R8126 VPWR.n465 VPWR.t1385 738.074
R8127 VPWR.n464 VPWR.t562 738.074
R8128 VPWR.n461 VPWR.t448 738.074
R8129 VPWR.n460 VPWR.t1736 738.074
R8130 VPWR.n457 VPWR.t1900 738.074
R8131 VPWR.n456 VPWR.t183 738.074
R8132 VPWR.n453 VPWR.t1207 738.074
R8133 VPWR.n452 VPWR.t5 738.074
R8134 VPWR.n473 VPWR.t147 738.074
R8135 VPWR.n482 VPWR.t1466 738.074
R8136 VPWR.n538 VPWR.t1620 738.074
R8137 VPWR.n534 VPWR.t1713 738.074
R8138 VPWR.n530 VPWR.t1166 738.074
R8139 VPWR.n522 VPWR.t1527 738.074
R8140 VPWR.n518 VPWR.t1481 738.074
R8141 VPWR.n514 VPWR.t1860 738.074
R8142 VPWR.n510 VPWR.t500 738.074
R8143 VPWR.n506 VPWR.t1039 738.074
R8144 VPWR.n502 VPWR.t381 738.074
R8145 VPWR.n498 VPWR.t1513 738.074
R8146 VPWR.n494 VPWR.t36 738.074
R8147 VPWR.n490 VPWR.t283 738.074
R8148 VPWR.n486 VPWR.t528 738.074
R8149 VPWR.n483 VPWR.t193 738.074
R8150 VPWR.n526 VPWR.t1045 738.074
R8151 VPWR.n548 VPWR.t1452 738.074
R8152 VPWR.n549 VPWR.t558 738.074
R8153 VPWR.n552 VPWR.t1648 738.074
R8154 VPWR.n553 VPWR.t1144 738.074
R8155 VPWR.n557 VPWR.t1555 738.074
R8156 VPWR.n560 VPWR.t1497 738.074
R8157 VPWR.n561 VPWR.t1698 738.074
R8158 VPWR.n564 VPWR.t251 738.074
R8159 VPWR.n565 VPWR.t523 738.074
R8160 VPWR.n568 VPWR.t436 738.074
R8161 VPWR.n569 VPWR.t476 738.074
R8162 VPWR.n572 VPWR.t1442 738.074
R8163 VPWR.n573 VPWR.t167 738.074
R8164 VPWR.n576 VPWR.t1569 738.074
R8165 VPWR.n577 VPWR.t1636 738.074
R8166 VPWR.n556 VPWR.t1069 738.074
R8167 VPWR.n579 VPWR.t1460 738.074
R8168 VPWR.n583 VPWR.t984 738.074
R8169 VPWR.n587 VPWR.t1547 738.074
R8170 VPWR.n591 VPWR.t1158 738.074
R8171 VPWR.n599 VPWR.t114 738.074
R8172 VPWR.n603 VPWR.t1260 738.074
R8173 VPWR.n607 VPWR.t1870 738.074
R8174 VPWR.n611 VPWR.t277 738.074
R8175 VPWR.n615 VPWR.t321 738.074
R8176 VPWR.n619 VPWR.t402 738.074
R8177 VPWR.n623 VPWR.t1750 738.074
R8178 VPWR.n627 VPWR.t963 738.074
R8179 VPWR.n631 VPWR.t291 738.074
R8180 VPWR.n635 VPWR.t1421 738.074
R8181 VPWR.n578 VPWR.t390 738.074
R8182 VPWR.n595 VPWR.t1051 738.074
R8183 VPWR.n673 VPWR.t1472 738.074
R8184 VPWR.n672 VPWR.t309 738.074
R8185 VPWR.n669 VPWR.t1608 738.074
R8186 VPWR.n668 VPWR.t1180 738.074
R8187 VPWR.n664 VPWR.t1521 738.074
R8188 VPWR.n661 VPWR.t1272 738.074
R8189 VPWR.n660 VPWR.t231 738.074
R8190 VPWR.n657 VPWR.t1406 738.074
R8191 VPWR.n656 VPWR.t131 738.074
R8192 VPWR.n653 VPWR.t357 738.074
R8193 VPWR.n652 VPWR.t1119 738.074
R8194 VPWR.n649 VPWR.t1537 738.074
R8195 VPWR.n648 VPWR.t50 738.074
R8196 VPWR.n645 VPWR.t486 738.074
R8197 VPWR.n644 VPWR.t207 738.074
R8198 VPWR.n665 VPWR.t1028 738.074
R8199 VPWR.n674 VPWR.t1479 738.074
R8200 VPWR.n730 VPWR.t1110 738.074
R8201 VPWR.n726 VPWR.t127 738.074
R8202 VPWR.n722 VPWR.t1192 738.074
R8203 VPWR.n714 VPWR.t1578 738.074
R8204 VPWR.n710 VPWR.t1288 738.074
R8205 VPWR.n706 VPWR.t953 738.074
R8206 VPWR.n702 VPWR.t959 738.074
R8207 VPWR.n698 VPWR.t560 738.074
R8208 VPWR.n694 VPWR.t446 738.074
R8209 VPWR.n690 VPWR.t1734 738.074
R8210 VPWR.n686 VPWR.t1898 738.074
R8211 VPWR.n682 VPWR.t181 738.074
R8212 VPWR.n678 VPWR.t1205 738.074
R8213 VPWR.n675 VPWR.t1646 738.074
R8214 VPWR.n718 VPWR.t145 738.074
R8215 VPWR.n740 VPWR.t1475 738.074
R8216 VPWR.n741 VPWR.t460 738.074
R8217 VPWR.n744 VPWR.t511 738.074
R8218 VPWR.n745 VPWR.t1186 738.074
R8219 VPWR.n749 VPWR.t1307 738.074
R8220 VPWR.n752 VPWR.t1344 738.074
R8221 VPWR.n753 VPWR.t227 738.074
R8222 VPWR.n756 VPWR.t1387 738.074
R8223 VPWR.n757 VPWR.t1222 738.074
R8224 VPWR.n760 VPWR.t351 738.074
R8225 VPWR.n761 VPWR.t1849 738.074
R8226 VPWR.n764 VPWR.t1885 738.074
R8227 VPWR.n765 VPWR.t40 738.074
R8228 VPWR.n768 VPWR.t1586 738.074
R8229 VPWR.n769 VPWR.t7 738.074
R8230 VPWR.n748 VPWR.t149 738.074
R8231 VPWR.n771 VPWR.t1454 738.074
R8232 VPWR.n775 VPWR.t556 738.074
R8233 VPWR.n779 VPWR.t517 738.074
R8234 VPWR.n783 VPWR.t1146 738.074
R8235 VPWR.n791 VPWR.t1553 738.074
R8236 VPWR.n795 VPWR.t1495 738.074
R8237 VPWR.n799 VPWR.t1696 738.074
R8238 VPWR.n803 VPWR.t247 738.074
R8239 VPWR.n807 VPWR.t521 738.074
R8240 VPWR.n811 VPWR.t375 738.074
R8241 VPWR.n815 VPWR.t474 738.074
R8242 VPWR.n819 VPWR.t1360 738.074
R8243 VPWR.n823 VPWR.t163 738.074
R8244 VPWR.n827 VPWR.t1567 738.074
R8245 VPWR.n770 VPWR.t1632 738.074
R8246 VPWR.n787 VPWR.t1065 738.074
R8247 VPWR.n865 VPWR.t1470 738.074
R8248 VPWR.n864 VPWR.t311 738.074
R8249 VPWR.n861 VPWR.t1610 738.074
R8250 VPWR.n860 VPWR.t1178 738.074
R8251 VPWR.n856 VPWR.t1523 738.074
R8252 VPWR.n853 VPWR.t1274 738.074
R8253 VPWR.n852 VPWR.t233 738.074
R8254 VPWR.n849 VPWR.t241 738.074
R8255 VPWR.n848 VPWR.t133 738.074
R8256 VPWR.n845 VPWR.t359 738.074
R8257 VPWR.n844 VPWR.t1121 738.074
R8258 VPWR.n841 VPWR.t1539 738.074
R8259 VPWR.n840 VPWR.t52 738.074
R8260 VPWR.n837 VPWR.t488 738.074
R8261 VPWR.n836 VPWR.t209 738.074
R8262 VPWR.n857 VPWR.t1061 738.074
R8263 VPWR.n866 VPWR.t1456 738.074
R8264 VPWR.n922 VPWR.t554 738.074
R8265 VPWR.n918 VPWR.t515 738.074
R8266 VPWR.n914 VPWR.t1148 738.074
R8267 VPWR.n906 VPWR.t1700 738.074
R8268 VPWR.n902 VPWR.t1493 738.074
R8269 VPWR.n898 VPWR.t1694 738.074
R8270 VPWR.n894 VPWR.t269 738.074
R8271 VPWR.n890 VPWR.t519 738.074
R8272 VPWR.n886 VPWR.t373 738.074
R8273 VPWR.n882 VPWR.t472 738.074
R8274 VPWR.n878 VPWR.t1358 738.074
R8275 VPWR.n874 VPWR.t159 738.074
R8276 VPWR.n870 VPWR.t1565 738.074
R8277 VPWR.n867 VPWR.t1630 738.074
R8278 VPWR.n910 VPWR.t1063 738.074
R8279 VPWR.n940 VPWR.t1049 738.074
R8280 VPWR.n979 VPWR.t1075 738.074
R8281 VPWR.n1179 VPWR.t631 738.074
R8282 VPWR.n399 VPWR.t1174 738.074
R8283 VPWR.n361 VPWR.t1156 738.074
R8284 VPWR.n338 VPWR.t1164 738.074
R8285 VPWR.n92 VPWR.t640 738.074
R8286 VPWR.n975 VPWR.t1138 738.074
R8287 VPWR.n1183 VPWR.t913 738.074
R8288 VPWR.n941 VPWR.t110 738.074
R8289 VPWR.n983 VPWR.t1561 738.074
R8290 VPWR.n1217 VPWR.t643 738.074
R8291 VPWR.n407 VPWR.t1525 738.074
R8292 VPWR.n415 VPWR.t235 738.074
R8293 VPWR.n419 VPWR.t243 738.074
R8294 VPWR.n423 VPWR.t135 738.074
R8295 VPWR.n427 VPWR.t361 738.074
R8296 VPWR.n431 VPWR.t1123 738.074
R8297 VPWR.n435 VPWR.t1541 738.074
R8298 VPWR.n439 VPWR.t54 738.074
R8299 VPWR.n443 VPWR.t490 738.074
R8300 VPWR.n386 VPWR.t187 738.074
R8301 VPWR.n411 VPWR.t1276 738.074
R8302 VPWR.n368 VPWR.t1262 738.074
R8303 VPWR.n326 VPWR.t1483 738.074
R8304 VPWR.n81 VPWR.t916 738.074
R8305 VPWR.n987 VPWR.t1503 738.074
R8306 VPWR.n1214 VPWR.t802 738.074
R8307 VPWR.n944 VPWR.t1487 738.074
R8308 VPWR.n948 VPWR.t275 738.074
R8309 VPWR.n949 VPWR.t317 738.074
R8310 VPWR.n952 VPWR.t385 738.074
R8311 VPWR.n953 VPWR.t1746 738.074
R8312 VPWR.n956 VPWR.t961 738.074
R8313 VPWR.n957 VPWR.t289 738.074
R8314 VPWR.n960 VPWR.t1419 738.074
R8315 VPWR.n961 VPWR.t197 738.074
R8316 VPWR.n945 VPWR.t1866 738.074
R8317 VPWR.n991 VPWR.t215 738.074
R8318 VPWR.n1206 VPWR.t910 738.074
R8319 VPWR.n360 VPWR.t1549 738.074
R8320 VPWR.n342 VPWR.t1715 738.074
R8321 VPWR.n93 VPWR.t875 738.074
R8322 VPWR.n1180 VPWR.t748 738.074
R8323 VPWR.n995 VPWR.t255 738.074
R8324 VPWR.n1203 VPWR.t671 738.074
R8325 VPWR.n372 VPWR.t279 738.074
R8326 VPWR.n376 VPWR.t404 738.074
R8327 VPWR.n377 VPWR.t1752 738.074
R8328 VPWR.n380 VPWR.t965 738.074
R8329 VPWR.n381 VPWR.t293 738.074
R8330 VPWR.n384 VPWR.t1423 738.074
R8331 VPWR.n385 VPWR.t394 738.074
R8332 VPWR.n373 VPWR.t323 738.074
R8333 VPWR.n314 VPWR.t1041 738.074
R8334 VPWR.n74 VPWR.t813 738.074
R8335 VPWR.n1200 VPWR.t697 738.074
R8336 VPWR.n999 VPWR.t72 738.074
R8337 VPWR.n1003 VPWR.t438 738.074
R8338 VPWR.n1007 VPWR.t482 738.074
R8339 VPWR.n1011 VPWR.t1444 738.074
R8340 VPWR.n1015 VPWR.t173 738.074
R8341 VPWR.n1019 VPWR.t104 738.074
R8342 VPWR.n962 VPWR.t1642 738.074
R8343 VPWR.n967 VPWR.t1102 738.074
R8344 VPWR.n1123 VPWR.t646 738.074
R8345 VPWR.n310 VPWR.t383 738.074
R8346 VPWR.n69 VPWR.t943 738.074
R8347 VPWR.n1192 VPWR.t824 738.074
R8348 VPWR.n1189 VPWR.t570 738.074
R8349 VPWR.n306 VPWR.t1515 738.074
R8350 VPWR.n302 VPWR.t38 738.074
R8351 VPWR.n294 VPWR.t530 738.074
R8352 VPWR.n291 VPWR.t195 738.074
R8353 VPWR.n298 VPWR.t287 738.074
R8354 VPWR.n1058 VPWR.t829 738.074
R8355 VPWR.n1186 VPWR.t591 738.074
R8356 VPWR.n63 VPWR.t717 738.074
R8357 VPWR.n62 VPWR.t567 738.074
R8358 VPWR.n57 VPWR.t586 738.074
R8359 VPWR.n56 VPWR.t711 738.074
R8360 VPWR.n1059 VPWR.t857 738.074
R8361 VPWR.n1061 VPWR.t577 738.074
R8362 VPWR.n2856 VPWR.n2821 702.354
R8363 VPWR.n2856 VPWR.n2822 702.354
R8364 VPWR.n2854 VPWR.n2853 702.354
R8365 VPWR.n2854 VPWR.n2821 702.354
R8366 VPWR.n2837 VPWR.n2828 702.354
R8367 VPWR.n2850 VPWR.n2849 702.354
R8368 VPWR.n2835 VPWR.n2828 702.354
R8369 VPWR.n2815 VPWR.t267 651.634
R8370 VPWR.n2831 VPWR.t1473 651.505
R8371 VPWR.n2825 VPWR.t94 651.505
R8372 VPWR.n2862 VPWR.t1095 651.431
R8373 VPWR.n1061 VPWR.t700 646.071
R8374 VPWR.n1122 VPWR.t596 646.071
R8375 VPWR.n1059 VPWR.t849 646.071
R8376 VPWR.n56 VPWR.t816 646.071
R8377 VPWR.n62 VPWR.t940 646.071
R8378 VPWR.n99 VPWR.t725 646.071
R8379 VPWR.n1053 VPWR.t179 646.071
R8380 VPWR.n1231 VPWR.t66 646.071
R8381 VPWR.n298 VPWR.t1427 646.071
R8382 VPWR.n290 VPWR.t990 646.071
R8383 VPWR.n306 VPWR.t969 646.071
R8384 VPWR.n68 VPWR.t679 646.071
R8385 VPWR.n1153 VPWR.t201 646.071
R8386 VPWR.n346 VPWR.t1545 646.071
R8387 VPWR.n98 VPWR.t854 646.071
R8388 VPWR.n967 VPWR.t125 646.071
R8389 VPWR.n963 VPWR.t88 646.071
R8390 VPWR.n999 VPWR.t450 646.071
R8391 VPWR.n373 VPWR.t414 646.071
R8392 VPWR.n356 VPWR.t64 646.071
R8393 VPWR.n357 VPWR.t1531 646.071
R8394 VPWR.n372 VPWR.t1112 646.071
R8395 VPWR.n318 VPWR.t319 646.071
R8396 VPWR.n75 VPWR.t784 646.071
R8397 VPWR.n971 VPWR.t1172 646.071
R8398 VPWR.n369 VPWR.t955 646.071
R8399 VPWR.n322 VPWR.t249 646.071
R8400 VPWR.n80 VPWR.t656 646.071
R8401 VPWR.n945 VPWR.t253 646.071
R8402 VPWR.n932 VPWR.t992 646.071
R8403 VPWR.n933 VPWR.t1551 646.071
R8404 VPWR.n936 VPWR.t1136 646.071
R8405 VPWR.n944 VPWR.t1686 646.071
R8406 VPWR.n411 VPWR.t1858 646.071
R8407 VPWR.n387 VPWR.t1618 646.071
R8408 VPWR.n391 VPWR.t1709 646.071
R8409 VPWR.n395 VPWR.t1150 646.071
R8410 VPWR.n407 VPWR.t1282 646.071
R8411 VPWR.n365 VPWR.t1268 646.071
R8412 VPWR.n330 VPWR.t1258 646.071
R8413 VPWR.n86 VPWR.t897 646.071
R8414 VPWR.n937 VPWR.t1067 646.071
R8415 VPWR.n403 VPWR.t1319 646.071
R8416 VPWR.n364 VPWR.t1604 646.071
R8417 VPWR.n334 VPWR.t112 646.071
R8418 VPWR.n87 VPWR.t742 646.071
R8419 VPWR.n473 VPWR.t1305 646.071
R8420 VPWR.n481 VPWR.t462 646.071
R8421 VPWR.n480 VPWR.t509 646.071
R8422 VPWR.n477 VPWR.t1168 646.071
R8423 VPWR.n476 VPWR.t1413 646.071
R8424 VPWR.n472 VPWR.t1342 646.071
R8425 VPWR.n469 VPWR.t225 646.071
R8426 VPWR.n468 VPWR.t169 646.071
R8427 VPWR.n465 VPWR.t1220 646.071
R8428 VPWR.n464 VPWR.t353 646.071
R8429 VPWR.n461 VPWR.t452 646.071
R8430 VPWR.n460 VPWR.t1887 646.071
R8431 VPWR.n457 VPWR.t281 646.071
R8432 VPWR.n456 VPWR.t1083 646.071
R8433 VPWR.n453 VPWR.t189 646.071
R8434 VPWR.n452 VPWR.t714 646.071
R8435 VPWR.n526 VPWR.t108 646.071
R8436 VPWR.n482 VPWR.t988 646.071
R8437 VPWR.n538 VPWR.t1717 646.071
R8438 VPWR.n534 VPWR.t1142 646.071
R8439 VPWR.n530 VPWR.t1079 646.071
R8440 VPWR.n522 VPWR.t1485 646.071
R8441 VPWR.n518 VPWR.t1864 646.071
R8442 VPWR.n514 VPWR.t271 646.071
R8443 VPWR.n510 VPWR.t1043 646.071
R8444 VPWR.n506 VPWR.t406 646.071
R8445 VPWR.n502 VPWR.t1744 646.071
R8446 VPWR.n498 VPWR.t967 646.071
R8447 VPWR.n494 VPWR.t161 646.071
R8448 VPWR.n490 VPWR.t1425 646.071
R8449 VPWR.n486 VPWR.t400 646.071
R8450 VPWR.n483 VPWR.t932 646.071
R8451 VPWR.n556 VPWR.t1563 646.071
R8452 VPWR.n548 VPWR.t1108 646.071
R8453 VPWR.n549 VPWR.t1656 646.071
R8454 VPWR.n552 VPWR.t1182 646.071
R8455 VPWR.n553 VPWR.t1024 646.071
R8456 VPWR.n557 VPWR.t1505 646.071
R8457 VPWR.n560 VPWR.t217 646.071
R8458 VPWR.n561 VPWR.t1402 646.071
R8459 VPWR.n564 VPWR.t74 646.071
R8460 VPWR.n565 VPWR.t444 646.071
R8461 VPWR.n568 VPWR.t484 646.071
R8462 VPWR.n569 VPWR.t1896 646.071
R8463 VPWR.n572 VPWR.t46 646.071
R8464 VPWR.n573 VPWR.t1203 646.071
R8465 VPWR.n576 VPWR.t203 646.071
R8466 VPWR.n577 VPWR.t781 646.071
R8467 VPWR.n595 VPWR.t1602 646.071
R8468 VPWR.n579 VPWR.t994 646.071
R8469 VPWR.n583 VPWR.t315 646.071
R8470 VPWR.n587 VPWR.t1134 646.071
R8471 VPWR.n591 VPWR.t1071 646.071
R8472 VPWR.n599 VPWR.t1266 646.071
R8473 VPWR.n603 VPWR.t1688 646.071
R8474 VPWR.n607 VPWR.t257 646.071
R8475 VPWR.n611 VPWR.t327 646.071
R8476 VPWR.n615 VPWR.t412 646.071
R8477 VPWR.n619 VPWR.t1756 646.071
R8478 VPWR.n623 VPWR.t494 646.071
R8479 VPWR.n627 VPWR.t175 646.071
R8480 VPWR.n631 VPWR.t1431 646.071
R8481 VPWR.n635 VPWR.t1638 646.071
R8482 VPWR.n578 VPWR.t889 646.071
R8483 VPWR.n665 VPWR.t1315 646.071
R8484 VPWR.n673 VPWR.t996 646.071
R8485 VPWR.n672 VPWR.t1614 646.071
R8486 VPWR.n669 VPWR.t1154 646.071
R8487 VPWR.n668 VPWR.t1053 646.071
R8488 VPWR.n664 VPWR.t1278 646.071
R8489 VPWR.n661 VPWR.t237 646.071
R8490 VPWR.n660 VPWR.t532 646.071
R8491 VPWR.n657 VPWR.t137 646.071
R8492 VPWR.n656 VPWR.t363 646.071
R8493 VPWR.n653 VPWR.t1125 646.071
R8494 VPWR.n652 VPWR.t1840 646.071
R8495 VPWR.n649 VPWR.t295 646.071
R8496 VPWR.n648 VPWR.t492 646.071
R8497 VPWR.n645 VPWR.t392 646.071
R8498 VPWR.n644 VPWR.t615 646.071
R8499 VPWR.n718 VPWR.t1303 646.071
R8500 VPWR.n674 VPWR.t90 646.071
R8501 VPWR.n730 VPWR.t507 646.071
R8502 VPWR.n726 VPWR.t1170 646.071
R8503 VPWR.n722 VPWR.t1409 646.071
R8504 VPWR.n714 VPWR.t1292 646.071
R8505 VPWR.n710 VPWR.t223 646.071
R8506 VPWR.n706 VPWR.t245 646.071
R8507 VPWR.n702 VPWR.t564 646.071
R8508 VPWR.n698 VPWR.t349 646.071
R8509 VPWR.n694 VPWR.t1738 646.071
R8510 VPWR.n690 VPWR.t1883 646.071
R8511 VPWR.n686 VPWR.t56 646.071
R8512 VPWR.n682 VPWR.t1584 646.071
R8513 VPWR.n678 VPWR.t185 646.071
R8514 VPWR.n675 VPWR.t722 646.071
R8515 VPWR.n748 VPWR.t1309 646.071
R8516 VPWR.n740 VPWR.t464 646.071
R8517 VPWR.n741 VPWR.t513 646.071
R8518 VPWR.n744 VPWR.t1162 646.071
R8519 VPWR.n745 VPWR.t1415 646.071
R8520 VPWR.n749 VPWR.t1346 646.071
R8521 VPWR.n752 VPWR.t229 646.071
R8522 VPWR.n753 VPWR.t502 646.071
R8523 VPWR.n756 VPWR.t1224 646.071
R8524 VPWR.n757 VPWR.t355 646.071
R8525 VPWR.n760 VPWR.t1851 646.071
R8526 VPWR.n761 VPWR.t1535 646.071
R8527 VPWR.n764 VPWR.t285 646.071
R8528 VPWR.n765 VPWR.t1085 646.071
R8529 VPWR.n768 VPWR.t191 646.071
R8530 VPWR.n769 VPWR.t682 646.071
R8531 VPWR.n787 VPWR.t1559 646.071
R8532 VPWR.n771 VPWR.t1106 646.071
R8533 VPWR.n775 VPWR.t1652 646.071
R8534 VPWR.n779 VPWR.t1176 646.071
R8535 VPWR.n783 VPWR.t153 646.071
R8536 VPWR.n791 VPWR.t1501 646.071
R8537 VPWR.n795 VPWR.t213 646.071
R8538 VPWR.n799 VPWR.t1400 646.071
R8539 VPWR.n803 VPWR.t70 646.071
R8540 VPWR.n807 VPWR.t442 646.071
R8541 VPWR.n811 VPWR.t480 646.071
R8542 VPWR.n815 VPWR.t1448 646.071
R8543 VPWR.n819 VPWR.t44 646.071
R8544 VPWR.n823 VPWR.t1201 646.071
R8545 VPWR.n827 VPWR.t11 646.071
R8546 VPWR.n770 VPWR.t787 646.071
R8547 VPWR.n857 VPWR.t1317 646.071
R8548 VPWR.n865 VPWR.t1616 646.071
R8549 VPWR.n864 VPWR.t1707 646.071
R8550 VPWR.n861 VPWR.t1152 646.071
R8551 VPWR.n860 VPWR.t1057 646.071
R8552 VPWR.n856 VPWR.t1280 646.071
R8553 VPWR.n853 VPWR.t239 646.071
R8554 VPWR.n852 VPWR.t534 646.071
R8555 VPWR.n849 VPWR.t139 646.071
R8556 VPWR.n848 VPWR.t377 646.071
R8557 VPWR.n845 VPWR.t1509 646.071
R8558 VPWR.n844 VPWR.t1842 646.071
R8559 VPWR.n841 VPWR.t297 646.071
R8560 VPWR.n840 VPWR.t973 646.071
R8561 VPWR.n837 VPWR.t396 646.071
R8562 VPWR.n836 VPWR.t610 646.071
R8563 VPWR.n910 VPWR.t1557 646.071
R8564 VPWR.n866 VPWR.t1104 646.071
R8565 VPWR.n922 VPWR.t1650 646.071
R8566 VPWR.n918 VPWR.t1184 646.071
R8567 VPWR.n914 VPWR.t151 646.071
R8568 VPWR.n906 VPWR.t1499 646.071
R8569 VPWR.n902 VPWR.t211 646.071
R8570 VPWR.n898 VPWR.t1398 646.071
R8571 VPWR.n894 VPWR.t68 646.071
R8572 VPWR.n890 VPWR.t440 646.071
R8573 VPWR.n886 VPWR.t478 646.071
R8574 VPWR.n882 VPWR.t1446 646.071
R8575 VPWR.n878 VPWR.t42 646.071
R8576 VPWR.n874 VPWR.t106 646.071
R8577 VPWR.n870 VPWR.t9 646.071
R8578 VPWR.n867 VPWR.t794 646.071
R8579 VPWR.n940 VPWR.t118 646.071
R8580 VPWR.n979 VPWR.t1576 646.071
R8581 VPWR.n1227 VPWR.t1606 646.071
R8582 VPWR.n1179 VPWR.t626 646.071
R8583 VPWR.n399 VPWR.t1059 646.071
R8584 VPWR.n361 VPWR.t1073 646.071
R8585 VPWR.n338 VPWR.t1081 646.071
R8586 VPWR.n92 VPWR.t634 646.071
R8587 VPWR.n975 VPWR.t1026 646.071
R8588 VPWR.n1485 VPWR.t1077 646.071
R8589 VPWR.n1183 VPWR.t905 646.071
R8590 VPWR.n941 VPWR.t1264 646.071
R8591 VPWR.n983 VPWR.t1286 646.071
R8592 VPWR.n1173 VPWR.t1763 646.071
R8593 VPWR.n1217 VPWR.t773 646.071
R8594 VPWR.n415 VPWR.t536 646.071
R8595 VPWR.n419 VPWR.t982 646.071
R8596 VPWR.n423 VPWR.t379 646.071
R8597 VPWR.n427 VPWR.t1511 646.071
R8598 VPWR.n431 VPWR.t1844 646.071
R8599 VPWR.n435 VPWR.t299 646.071
R8600 VPWR.n439 VPWR.t975 646.071
R8601 VPWR.n443 VPWR.t398 646.071
R8602 VPWR.n386 VPWR.t602 646.071
R8603 VPWR.n368 VPWR.t1690 646.071
R8604 VPWR.n326 VPWR.t1868 646.071
R8605 VPWR.n81 VPWR.t621 646.071
R8606 VPWR.n987 VPWR.t219 646.071
R8607 VPWR.n1169 VPWR.t1692 646.071
R8608 VPWR.n1214 VPWR.t884 646.071
R8609 VPWR.n948 VPWR.t325 646.071
R8610 VPWR.n949 VPWR.t410 646.071
R8611 VPWR.n952 VPWR.t1754 646.071
R8612 VPWR.n953 VPWR.t971 646.071
R8613 VPWR.n956 VPWR.t171 646.071
R8614 VPWR.n957 VPWR.t1429 646.071
R8615 VPWR.n960 VPWR.t1634 646.071
R8616 VPWR.n961 VPWR.t902 646.071
R8617 VPWR.n991 VPWR.t1404 646.071
R8618 VPWR.n1163 VPWR.t957 646.071
R8619 VPWR.n1206 VPWR.t921 646.071
R8620 VPWR.n360 VPWR.t1132 646.071
R8621 VPWR.n342 VPWR.t1140 646.071
R8622 VPWR.n93 VPWR.t872 646.071
R8623 VPWR.n1479 VPWR.t1188 646.071
R8624 VPWR.n1180 VPWR.t745 646.071
R8625 VPWR.n995 VPWR.t76 646.071
R8626 VPWR.n1159 VPWR.t1114 646.071
R8627 VPWR.n1203 VPWR.t666 646.071
R8628 VPWR.n376 VPWR.t199 646.071
R8629 VPWR.n377 VPWR.t496 646.071
R8630 VPWR.n380 VPWR.t177 646.071
R8631 VPWR.n381 VPWR.t1433 646.071
R8632 VPWR.n384 VPWR.t1640 646.071
R8633 VPWR.n385 VPWR.t881 646.071
R8634 VPWR.n314 VPWR.t408 646.071
R8635 VPWR.n74 VPWR.t894 646.071
R8636 VPWR.n1149 VPWR.t416 646.071
R8637 VPWR.n1200 VPWR.t770 646.071
R8638 VPWR.n1003 VPWR.t1732 646.071
R8639 VPWR.n1007 VPWR.t1902 646.071
R8640 VPWR.n1011 VPWR.t48 646.071
R8641 VPWR.n1015 VPWR.t1582 646.071
R8642 VPWR.n1019 VPWR.t205 646.071
R8643 VPWR.n962 VPWR.t754 646.071
R8644 VPWR.n1472 VPWR.t1533 646.071
R8645 VPWR.n1123 VPWR.t732 646.071
R8646 VPWR.n310 VPWR.t1748 646.071
R8647 VPWR.n69 VPWR.t661 646.071
R8648 VPWR.n1192 VPWR.t929 646.071
R8649 VPWR.n1049 VPWR.t498 646.071
R8650 VPWR.n1189 VPWR.t948 646.071
R8651 VPWR.n302 VPWR.t165 646.071
R8652 VPWR.n294 VPWR.t1628 646.071
R8653 VPWR.n291 VPWR.t924 646.071
R8654 VPWR.n1058 VPWR.t821 646.071
R8655 VPWR.n1748 VPWR.t1417 646.071
R8656 VPWR.n1036 VPWR.t1644 646.071
R8657 VPWR.n1032 VPWR.t865 646.071
R8658 VPWR.n1186 VPWR.t692 646.071
R8659 VPWR.n63 VPWR.t807 646.071
R8660 VPWR.n57 VPWR.t580 646.071
R8661 VPWR.n1230 VPWR.t674 642.13
R8662 VPWR.n1152 VPWR.t605 642.13
R8663 VPWR.n1226 VPWR.t810 642.13
R8664 VPWR.n1484 VPWR.t708 642.13
R8665 VPWR.n1172 VPWR.t832 642.13
R8666 VPWR.n1168 VPWR.t583 642.13
R8667 VPWR.n1162 VPWR.t705 642.13
R8668 VPWR.n1478 VPWR.t937 642.13
R8669 VPWR.n1158 VPWR.t846 642.13
R8670 VPWR.n1148 VPWR.t862 642.13
R8671 VPWR.n1471 VPWR.t835 642.13
R8672 VPWR.n1048 VPWR.t735 642.13
R8673 VPWR.n1747 VPWR.t599 642.13
R8674 VPWR.n1035 VPWR.t649 642.13
R8675 VPWR.n1031 VPWR.t757 642.13
R8676 VPWR.n1052 VPWR.t776 642.13
R8677 VPWR.n2309 VPWR.t461 629.652
R8678 VPWR.n2310 VPWR.t508 629.652
R8679 VPWR.n2319 VPWR.t1167 629.652
R8680 VPWR.n2320 VPWR.t1412 629.652
R8681 VPWR.n2329 VPWR.t1304 629.652
R8682 VPWR.n2330 VPWR.t1341 629.652
R8683 VPWR.n2339 VPWR.t224 629.652
R8684 VPWR.n2340 VPWR.t168 629.652
R8685 VPWR.n2349 VPWR.t1219 629.652
R8686 VPWR.n2350 VPWR.t352 629.652
R8687 VPWR.n2359 VPWR.t451 629.652
R8688 VPWR.n2360 VPWR.t1886 629.652
R8689 VPWR.n2369 VPWR.t280 629.652
R8690 VPWR.n2370 VPWR.t1082 629.652
R8691 VPWR.n2379 VPWR.t188 629.652
R8692 VPWR.n542 VPWR.t987 629.652
R8693 VPWR.t1716 VPWR.n541 629.652
R8694 VPWR.t1141 VPWR.n537 629.652
R8695 VPWR.t1078 VPWR.n533 629.652
R8696 VPWR.t107 VPWR.n529 629.652
R8697 VPWR.t1484 VPWR.n525 629.652
R8698 VPWR.t1863 VPWR.n521 629.652
R8699 VPWR.t270 VPWR.n517 629.652
R8700 VPWR.t1042 VPWR.n513 629.652
R8701 VPWR.t405 VPWR.n509 629.652
R8702 VPWR.t1743 VPWR.n505 629.652
R8703 VPWR.t966 VPWR.n501 629.652
R8704 VPWR.t160 VPWR.n497 629.652
R8705 VPWR.t1424 VPWR.n493 629.652
R8706 VPWR.t399 VPWR.n489 629.652
R8707 VPWR.n2281 VPWR.t1107 629.652
R8708 VPWR.t1655 VPWR.n2280 629.652
R8709 VPWR.n2271 VPWR.t1181 629.652
R8710 VPWR.t1023 VPWR.n2270 629.652
R8711 VPWR.n2261 VPWR.t1562 629.652
R8712 VPWR.t1504 VPWR.n2260 629.652
R8713 VPWR.n2251 VPWR.t216 629.652
R8714 VPWR.t1401 VPWR.n2250 629.652
R8715 VPWR.n2241 VPWR.t73 629.652
R8716 VPWR.t443 VPWR.n2240 629.652
R8717 VPWR.n2231 VPWR.t483 629.652
R8718 VPWR.t1895 VPWR.n2230 629.652
R8719 VPWR.n2221 VPWR.t45 629.652
R8720 VPWR.t1202 VPWR.n2220 629.652
R8721 VPWR.n2211 VPWR.t202 629.652
R8722 VPWR.n582 VPWR.t993 629.652
R8723 VPWR.n586 VPWR.t314 629.652
R8724 VPWR.n590 VPWR.t1133 629.652
R8725 VPWR.n594 VPWR.t1070 629.652
R8726 VPWR.n598 VPWR.t1601 629.652
R8727 VPWR.n602 VPWR.t1265 629.652
R8728 VPWR.n606 VPWR.t1687 629.652
R8729 VPWR.n610 VPWR.t256 629.652
R8730 VPWR.n614 VPWR.t326 629.652
R8731 VPWR.n618 VPWR.t411 629.652
R8732 VPWR.n622 VPWR.t1755 629.652
R8733 VPWR.n626 VPWR.t493 629.652
R8734 VPWR.n630 VPWR.t174 629.652
R8735 VPWR.n634 VPWR.t1430 629.652
R8736 VPWR.n638 VPWR.t1637 629.652
R8737 VPWR.n2113 VPWR.t995 629.652
R8738 VPWR.n2114 VPWR.t1613 629.652
R8739 VPWR.n2123 VPWR.t1153 629.652
R8740 VPWR.n2124 VPWR.t1052 629.652
R8741 VPWR.n2133 VPWR.t1314 629.652
R8742 VPWR.n2134 VPWR.t1277 629.652
R8743 VPWR.n2143 VPWR.t236 629.652
R8744 VPWR.n2144 VPWR.t531 629.652
R8745 VPWR.n2153 VPWR.t136 629.652
R8746 VPWR.n2154 VPWR.t362 629.652
R8747 VPWR.n2163 VPWR.t1124 629.652
R8748 VPWR.n2164 VPWR.t1839 629.652
R8749 VPWR.n2173 VPWR.t294 629.652
R8750 VPWR.n2174 VPWR.t491 629.652
R8751 VPWR.n2183 VPWR.t391 629.652
R8752 VPWR.n734 VPWR.t89 629.652
R8753 VPWR.t506 VPWR.n733 629.652
R8754 VPWR.t1169 VPWR.n729 629.652
R8755 VPWR.t1408 VPWR.n725 629.652
R8756 VPWR.t1302 VPWR.n721 629.652
R8757 VPWR.t1291 VPWR.n717 629.652
R8758 VPWR.t222 VPWR.n713 629.652
R8759 VPWR.t244 VPWR.n709 629.652
R8760 VPWR.t563 VPWR.n705 629.652
R8761 VPWR.t348 VPWR.n701 629.652
R8762 VPWR.t1737 VPWR.n697 629.652
R8763 VPWR.t1882 VPWR.n693 629.652
R8764 VPWR.t55 VPWR.n689 629.652
R8765 VPWR.t1583 VPWR.n685 629.652
R8766 VPWR.t184 VPWR.n681 629.652
R8767 VPWR.n2085 VPWR.t463 629.652
R8768 VPWR.t512 VPWR.n2084 629.652
R8769 VPWR.n2075 VPWR.t1161 629.652
R8770 VPWR.t1414 VPWR.n2074 629.652
R8771 VPWR.n2065 VPWR.t1308 629.652
R8772 VPWR.t1345 VPWR.n2064 629.652
R8773 VPWR.n2055 VPWR.t228 629.652
R8774 VPWR.t501 VPWR.n2054 629.652
R8775 VPWR.n2045 VPWR.t1223 629.652
R8776 VPWR.t354 VPWR.n2044 629.652
R8777 VPWR.n2035 VPWR.t1850 629.652
R8778 VPWR.t1534 VPWR.n2034 629.652
R8779 VPWR.n2025 VPWR.t284 629.652
R8780 VPWR.t1084 VPWR.n2024 629.652
R8781 VPWR.n2015 VPWR.t190 629.652
R8782 VPWR.n774 VPWR.t1105 629.652
R8783 VPWR.n778 VPWR.t1651 629.652
R8784 VPWR.n782 VPWR.t1175 629.652
R8785 VPWR.n786 VPWR.t152 629.652
R8786 VPWR.n790 VPWR.t1558 629.652
R8787 VPWR.n794 VPWR.t1500 629.652
R8788 VPWR.n798 VPWR.t212 629.652
R8789 VPWR.n802 VPWR.t1399 629.652
R8790 VPWR.n806 VPWR.t69 629.652
R8791 VPWR.n810 VPWR.t441 629.652
R8792 VPWR.n814 VPWR.t479 629.652
R8793 VPWR.n818 VPWR.t1447 629.652
R8794 VPWR.n822 VPWR.t43 629.652
R8795 VPWR.n826 VPWR.t1200 629.652
R8796 VPWR.n830 VPWR.t10 629.652
R8797 VPWR.n1917 VPWR.t1615 629.652
R8798 VPWR.n1918 VPWR.t1706 629.652
R8799 VPWR.n1927 VPWR.t1151 629.652
R8800 VPWR.n1928 VPWR.t1056 629.652
R8801 VPWR.n1937 VPWR.t1316 629.652
R8802 VPWR.n1938 VPWR.t1279 629.652
R8803 VPWR.n1947 VPWR.t238 629.652
R8804 VPWR.n1948 VPWR.t533 629.652
R8805 VPWR.n1957 VPWR.t138 629.652
R8806 VPWR.n1958 VPWR.t376 629.652
R8807 VPWR.n1967 VPWR.t1508 629.652
R8808 VPWR.n1968 VPWR.t1841 629.652
R8809 VPWR.n1977 VPWR.t296 629.652
R8810 VPWR.n1978 VPWR.t972 629.652
R8811 VPWR.n1987 VPWR.t395 629.652
R8812 VPWR.n926 VPWR.t1103 629.652
R8813 VPWR.t1649 VPWR.n925 629.652
R8814 VPWR.t1183 VPWR.n921 629.652
R8815 VPWR.t150 VPWR.n917 629.652
R8816 VPWR.t1556 VPWR.n913 629.652
R8817 VPWR.t1498 VPWR.n909 629.652
R8818 VPWR.t210 VPWR.n905 629.652
R8819 VPWR.t1397 VPWR.n901 629.652
R8820 VPWR.t67 VPWR.n897 629.652
R8821 VPWR.t439 VPWR.n893 629.652
R8822 VPWR.t477 VPWR.n889 629.652
R8823 VPWR.t1445 VPWR.n885 629.652
R8824 VPWR.t41 VPWR.n881 629.652
R8825 VPWR.t105 VPWR.n877 629.652
R8826 VPWR.t8 VPWR.n873 629.652
R8827 VPWR.n390 VPWR.t1617 629.652
R8828 VPWR.n394 VPWR.t1708 629.652
R8829 VPWR.n398 VPWR.t1149 629.652
R8830 VPWR.n402 VPWR.t1058 629.652
R8831 VPWR.n406 VPWR.t1318 629.652
R8832 VPWR.n410 VPWR.t1281 629.652
R8833 VPWR.n414 VPWR.t1857 629.652
R8834 VPWR.n418 VPWR.t535 629.652
R8835 VPWR.n422 VPWR.t981 629.652
R8836 VPWR.n426 VPWR.t378 629.652
R8837 VPWR.n430 VPWR.t1510 629.652
R8838 VPWR.n434 VPWR.t1843 629.652
R8839 VPWR.n438 VPWR.t298 629.652
R8840 VPWR.n442 VPWR.t974 629.652
R8841 VPWR.n446 VPWR.t397 629.652
R8842 VPWR.n1889 VPWR.t991 629.652
R8843 VPWR.t1550 VPWR.n1888 629.652
R8844 VPWR.n1879 VPWR.t1135 629.652
R8845 VPWR.t1066 VPWR.n1878 629.652
R8846 VPWR.n1869 VPWR.t117 629.652
R8847 VPWR.t1263 VPWR.n1868 629.652
R8848 VPWR.n1859 VPWR.t1685 629.652
R8849 VPWR.t252 VPWR.n1858 629.652
R8850 VPWR.n1849 VPWR.t324 629.652
R8851 VPWR.t409 VPWR.n1848 629.652
R8852 VPWR.n1839 VPWR.t1753 629.652
R8853 VPWR.t970 VPWR.n1838 629.652
R8854 VPWR.n1829 VPWR.t170 629.652
R8855 VPWR.t1428 VPWR.n1828 629.652
R8856 VPWR.n1819 VPWR.t1633 629.652
R8857 VPWR.n2477 VPWR.t63 629.652
R8858 VPWR.t1530 VPWR.n2476 629.652
R8859 VPWR.n2467 VPWR.t1131 629.652
R8860 VPWR.t1072 VPWR.n2466 629.652
R8861 VPWR.n2457 VPWR.t1603 629.652
R8862 VPWR.t1267 VPWR.n2456 629.652
R8863 VPWR.n2447 VPWR.t1689 629.652
R8864 VPWR.t954 VPWR.n2446 629.652
R8865 VPWR.n2437 VPWR.t1111 629.652
R8866 VPWR.t413 VPWR.n2436 629.652
R8867 VPWR.n2427 VPWR.t198 629.652
R8868 VPWR.t495 VPWR.n2426 629.652
R8869 VPWR.n2417 VPWR.t176 629.652
R8870 VPWR.t1432 VPWR.n2416 629.652
R8871 VPWR.n2407 VPWR.t1639 629.652
R8872 VPWR.n966 VPWR.t87 629.652
R8873 VPWR.n970 VPWR.t124 629.652
R8874 VPWR.n974 VPWR.t1171 629.652
R8875 VPWR.n978 VPWR.t1025 629.652
R8876 VPWR.n982 VPWR.t1575 629.652
R8877 VPWR.n986 VPWR.t1285 629.652
R8878 VPWR.n990 VPWR.t218 629.652
R8879 VPWR.n994 VPWR.t1403 629.652
R8880 VPWR.n998 VPWR.t75 629.652
R8881 VPWR.n1002 VPWR.t449 629.652
R8882 VPWR.n1006 VPWR.t1731 629.652
R8883 VPWR.n1010 VPWR.t1901 629.652
R8884 VPWR.n1014 VPWR.t47 629.652
R8885 VPWR.n1018 VPWR.t1581 629.652
R8886 VPWR.n1022 VPWR.t204 629.652
R8887 VPWR.n350 VPWR.t989 629.652
R8888 VPWR.t1544 VPWR.n349 629.652
R8889 VPWR.t1139 VPWR.n345 629.652
R8890 VPWR.t1080 VPWR.n341 629.652
R8891 VPWR.t111 VPWR.n337 629.652
R8892 VPWR.t1257 VPWR.n333 629.652
R8893 VPWR.t1867 VPWR.n329 629.652
R8894 VPWR.t248 VPWR.n325 629.652
R8895 VPWR.t318 VPWR.n321 629.652
R8896 VPWR.t407 VPWR.n317 629.652
R8897 VPWR.t1747 VPWR.n313 629.652
R8898 VPWR.t968 VPWR.n309 629.652
R8899 VPWR.t164 VPWR.n305 629.652
R8900 VPWR.t1426 VPWR.n301 629.652
R8901 VPWR.t1627 VPWR.n297 629.652
R8902 VPWR.n1468 VPWR.t65 629.652
R8903 VPWR.n1475 VPWR.t1532 629.652
R8904 VPWR.n1481 VPWR.t1187 629.652
R8905 VPWR.n1492 VPWR.t1076 629.652
R8906 VPWR.n1493 VPWR.t1605 629.652
R8907 VPWR.n1506 VPWR.t1762 629.652
R8908 VPWR.n1507 VPWR.t1691 629.652
R8909 VPWR.n1520 VPWR.t956 629.652
R8910 VPWR.n1521 VPWR.t1113 629.652
R8911 VPWR.n1536 VPWR.t415 629.652
R8912 VPWR.t200 VPWR.n1535 629.652
R8913 VPWR.n1761 VPWR.t497 629.652
R8914 VPWR.t178 VPWR.n1760 629.652
R8915 VPWR.n1749 VPWR.t1416 629.652
R8916 VPWR.n1791 VPWR.t1643 629.652
R8917 VPWR.n2506 VPWR.t724 629.652
R8918 VPWR.n2507 VPWR.t853 629.652
R8919 VPWR.n2518 VPWR.t871 629.652
R8920 VPWR.n2519 VPWR.t633 629.652
R8921 VPWR.n2530 VPWR.t741 629.652
R8922 VPWR.n2531 VPWR.t896 629.652
R8923 VPWR.n2542 VPWR.t620 629.652
R8924 VPWR.n2543 VPWR.t655 629.652
R8925 VPWR.n2554 VPWR.t783 629.652
R8926 VPWR.n2555 VPWR.t893 629.652
R8927 VPWR.n2566 VPWR.t660 629.652
R8928 VPWR.n2567 VPWR.t678 629.652
R8929 VPWR.n2578 VPWR.t806 629.652
R8930 VPWR.n2579 VPWR.t939 629.652
R8931 VPWR.n2590 VPWR.t579 629.652
R8932 VPWR.n1594 VPWR.t595 629.652
R8933 VPWR.t731 VPWR.n1593 629.652
R8934 VPWR.n1182 VPWR.t744 629.652
R8935 VPWR.n1185 VPWR.t904 629.652
R8936 VPWR.n1220 VPWR.t625 629.652
R8937 VPWR.t772 VPWR.n1219 629.652
R8938 VPWR.t883 VPWR.n1216 629.652
R8939 VPWR.t920 VPWR.n1213 629.652
R8940 VPWR.t665 VPWR.n1205 629.652
R8941 VPWR.t769 VPWR.n1202 629.652
R8942 VPWR.t928 VPWR.n1199 629.652
R8943 VPWR.t947 VPWR.n1191 629.652
R8944 VPWR.t691 VPWR.n1188 629.652
R8945 VPWR.n1740 VPWR.t820 629.652
R8946 VPWR.t848 VPWR.n1739 629.652
R8947 VPWR.n2836 VPWR.t93 531.804
R8948 VPWR.n2855 VPWR.t93 531.804
R8949 VPWR.n2851 VPWR.n2850 504.707
R8950 VPWR.t461 VPWR.t1677 486.048
R8951 VPWR.t508 VPWR.t1572 486.048
R8952 VPWR.t1855 VPWR.t1167 486.048
R8953 VPWR.t1412 VPWR.t1854 486.048
R8954 VPWR.t1676 VPWR.t1304 486.048
R8955 VPWR.t1341 VPWR.t1725 486.048
R8956 VPWR.t1724 VPWR.t224 486.048
R8957 VPWR.t168 VPWR.t1675 486.048
R8958 VPWR.t1574 VPWR.t1219 486.048
R8959 VPWR.t352 VPWR.t1726 486.048
R8960 VPWR.t1853 VPWR.t451 486.048
R8961 VPWR.t1886 VPWR.t1852 486.048
R8962 VPWR.t1723 VPWR.t280 486.048
R8963 VPWR.t1082 VPWR.t1722 486.048
R8964 VPWR.t1856 VPWR.t188 486.048
R8965 VPWR.t713 VPWR.t1573 486.048
R8966 VPWR.t987 VPWR.t1911 486.048
R8967 VPWR.t18 VPWR.t1716 486.048
R8968 VPWR.t1846 VPWR.t1141 486.048
R8969 VPWR.t1845 VPWR.t1078 486.048
R8970 VPWR.t1910 VPWR.t107 486.048
R8971 VPWR.t33 VPWR.t1484 486.048
R8972 VPWR.t32 VPWR.t1863 486.048
R8973 VPWR.t1909 VPWR.t270 486.048
R8974 VPWR.t20 VPWR.t1042 486.048
R8975 VPWR.t34 VPWR.t405 486.048
R8976 VPWR.t1913 VPWR.t1743 486.048
R8977 VPWR.t1912 VPWR.t966 486.048
R8978 VPWR.t31 VPWR.t160 486.048
R8979 VPWR.t30 VPWR.t1424 486.048
R8980 VPWR.t1847 VPWR.t399 486.048
R8981 VPWR.t19 VPWR.t931 486.048
R8982 VPWR.t1107 VPWR.t347 486.048
R8983 VPWR.t1683 VPWR.t1655 486.048
R8984 VPWR.t1181 VPWR.t1439 486.048
R8985 VPWR.t1438 VPWR.t1023 486.048
R8986 VPWR.t1562 VPWR.t346 486.048
R8987 VPWR.t1681 VPWR.t1504 486.048
R8988 VPWR.t216 VPWR.t1680 486.048
R8989 VPWR.t345 VPWR.t1401 486.048
R8990 VPWR.t73 VPWR.t344 486.048
R8991 VPWR.t1682 VPWR.t443 486.048
R8992 VPWR.t483 VPWR.t1437 486.048
R8993 VPWR.t1436 VPWR.t1895 486.048
R8994 VPWR.t45 VPWR.t1679 486.048
R8995 VPWR.t1678 VPWR.t1202 486.048
R8996 VPWR.t202 VPWR.t1440 486.048
R8997 VPWR.t1684 VPWR.t780 486.048
R8998 VPWR.t993 VPWR.t433 486.048
R8999 VPWR.t314 VPWR.t428 486.048
R9000 VPWR.t1133 VPWR.t470 486.048
R9001 VPWR.t1070 VPWR.t469 486.048
R9002 VPWR.t1601 VPWR.t432 486.048
R9003 VPWR.t1265 VPWR.t426 486.048
R9004 VPWR.t1687 VPWR.t425 486.048
R9005 VPWR.t256 VPWR.t431 486.048
R9006 VPWR.t326 VPWR.t430 486.048
R9007 VPWR.t411 VPWR.t427 486.048
R9008 VPWR.t1755 VPWR.t468 486.048
R9009 VPWR.t493 VPWR.t434 486.048
R9010 VPWR.t174 VPWR.t424 486.048
R9011 VPWR.t1430 VPWR.t423 486.048
R9012 VPWR.t1637 VPWR.t422 486.048
R9013 VPWR.t888 VPWR.t429 486.048
R9014 VPWR.t995 VPWR.t1089 486.048
R9015 VPWR.t1613 VPWR.t1090 486.048
R9016 VPWR.t1517 VPWR.t1153 486.048
R9017 VPWR.t1052 VPWR.t505 486.048
R9018 VPWR.t1088 VPWR.t1314 486.048
R9019 VPWR.t1277 VPWR.t97 486.048
R9020 VPWR.t96 VPWR.t236 486.048
R9021 VPWR.t531 VPWR.t1087 486.048
R9022 VPWR.t1086 VPWR.t136 486.048
R9023 VPWR.t362 VPWR.t98 486.048
R9024 VPWR.t504 VPWR.t1124 486.048
R9025 VPWR.t1839 VPWR.t503 486.048
R9026 VPWR.t95 VPWR.t294 486.048
R9027 VPWR.t491 VPWR.t1519 486.048
R9028 VPWR.t1518 VPWR.t391 486.048
R9029 VPWR.t614 VPWR.t1091 486.048
R9030 VPWR.t89 VPWR.t467 486.048
R9031 VPWR.t1674 VPWR.t506 486.048
R9032 VPWR.t1196 VPWR.t1169 486.048
R9033 VPWR.t1100 VPWR.t1408 486.048
R9034 VPWR.t466 VPWR.t1302 486.048
R9035 VPWR.t1672 VPWR.t1291 486.048
R9036 VPWR.t1671 VPWR.t222 486.048
R9037 VPWR.t465 VPWR.t244 486.048
R9038 VPWR.t1097 VPWR.t563 486.048
R9039 VPWR.t1673 VPWR.t348 486.048
R9040 VPWR.t1099 VPWR.t1737 486.048
R9041 VPWR.t1098 VPWR.t1882 486.048
R9042 VPWR.t1199 VPWR.t55 486.048
R9043 VPWR.t1198 VPWR.t1583 486.048
R9044 VPWR.t1197 VPWR.t184 486.048
R9045 VPWR.t1096 VPWR.t721 486.048
R9046 VPWR.t463 VPWR.t1250 486.048
R9047 VPWR.t1571 VPWR.t512 486.048
R9048 VPWR.t1161 VPWR.t1006 486.048
R9049 VPWR.t1005 VPWR.t1414 486.048
R9050 VPWR.t1308 VPWR.t1249 486.048
R9051 VPWR.t1011 VPWR.t1345 486.048
R9052 VPWR.t228 VPWR.t1010 486.048
R9053 VPWR.t1248 VPWR.t501 486.048
R9054 VPWR.t1223 VPWR.t1247 486.048
R9055 VPWR.t1570 VPWR.t354 486.048
R9056 VPWR.t1850 VPWR.t1004 486.048
R9057 VPWR.t1003 VPWR.t1534 486.048
R9058 VPWR.t284 VPWR.t1009 486.048
R9059 VPWR.t1008 VPWR.t1084 486.048
R9060 VPWR.t190 VPWR.t1007 486.048
R9061 VPWR.t1246 VPWR.t681 486.048
R9062 VPWR.t1105 VPWR.t1340 486.048
R9063 VPWR.t1651 VPWR.t1335 486.048
R9064 VPWR.t1175 VPWR.t1380 486.048
R9065 VPWR.t152 VPWR.t1379 486.048
R9066 VPWR.t1558 VPWR.t1339 486.048
R9067 VPWR.t1500 VPWR.t1333 486.048
R9068 VPWR.t212 VPWR.t1332 486.048
R9069 VPWR.t1399 VPWR.t1338 486.048
R9070 VPWR.t69 VPWR.t1337 486.048
R9071 VPWR.t441 VPWR.t1334 486.048
R9072 VPWR.t479 VPWR.t1378 486.048
R9073 VPWR.t1447 VPWR.t1377 486.048
R9074 VPWR.t43 VPWR.t1383 486.048
R9075 VPWR.t1200 VPWR.t1382 486.048
R9076 VPWR.t10 VPWR.t1381 486.048
R9077 VPWR.t786 VPWR.t1336 486.048
R9078 VPWR.t1615 VPWR.t1002 486.048
R9079 VPWR.t1706 VPWR.t997 486.048
R9080 VPWR.t331 VPWR.t1151 486.048
R9081 VPWR.t1056 VPWR.t330 486.048
R9082 VPWR.t1001 VPWR.t1316 486.048
R9083 VPWR.t1279 VPWR.t1904 486.048
R9084 VPWR.t1903 VPWR.t238 486.048
R9085 VPWR.t533 VPWR.t1000 486.048
R9086 VPWR.t999 VPWR.t138 486.048
R9087 VPWR.t376 VPWR.t1905 486.048
R9088 VPWR.t329 VPWR.t1508 486.048
R9089 VPWR.t1841 VPWR.t328 486.048
R9090 VPWR.t334 VPWR.t296 486.048
R9091 VPWR.t972 VPWR.t333 486.048
R9092 VPWR.t332 VPWR.t395 486.048
R9093 VPWR.t609 VPWR.t998 486.048
R9094 VPWR.t1103 VPWR.t1396 486.048
R9095 VPWR.t62 VPWR.t1649 486.048
R9096 VPWR.t1919 VPWR.t1183 486.048
R9097 VPWR.t1918 VPWR.t150 486.048
R9098 VPWR.t1395 VPWR.t1556 486.048
R9099 VPWR.t60 VPWR.t1498 486.048
R9100 VPWR.t59 VPWR.t210 486.048
R9101 VPWR.t1394 VPWR.t1397 486.048
R9102 VPWR.t1393 VPWR.t67 486.048
R9103 VPWR.t61 VPWR.t439 486.048
R9104 VPWR.t1917 VPWR.t477 486.048
R9105 VPWR.t1916 VPWR.t1445 486.048
R9106 VPWR.t58 VPWR.t41 486.048
R9107 VPWR.t57 VPWR.t105 486.048
R9108 VPWR.t1920 VPWR.t8 486.048
R9109 VPWR.t1392 VPWR.t793 486.048
R9110 VPWR.t1617 VPWR.t123 486.048
R9111 VPWR.t1708 VPWR.t980 486.048
R9112 VPWR.t1149 VPWR.t1323 486.048
R9113 VPWR.t1058 VPWR.t1322 486.048
R9114 VPWR.t1318 VPWR.t122 486.048
R9115 VPWR.t1281 VPWR.t1704 486.048
R9116 VPWR.t1857 VPWR.t1703 486.048
R9117 VPWR.t535 VPWR.t121 486.048
R9118 VPWR.t981 VPWR.t120 486.048
R9119 VPWR.t378 VPWR.t1705 486.048
R9120 VPWR.t1510 VPWR.t1321 486.048
R9121 VPWR.t1843 VPWR.t1320 486.048
R9122 VPWR.t298 VPWR.t1702 486.048
R9123 VPWR.t974 VPWR.t1701 486.048
R9124 VPWR.t397 VPWR.t1324 486.048
R9125 VPWR.t601 VPWR.t119 486.048
R9126 VPWR.t991 VPWR.t1921 486.048
R9127 VPWR.t25 VPWR.t1550 486.048
R9128 VPWR.t1135 VPWR.t1925 486.048
R9129 VPWR.t1924 VPWR.t1066 486.048
R9130 VPWR.t117 VPWR.t29 486.048
R9131 VPWR.t1330 VPWR.t1263 486.048
R9132 VPWR.t1685 VPWR.t1329 486.048
R9133 VPWR.t28 VPWR.t252 486.048
R9134 VPWR.t324 VPWR.t27 486.048
R9135 VPWR.t1331 VPWR.t409 486.048
R9136 VPWR.t1753 VPWR.t1923 486.048
R9137 VPWR.t1922 VPWR.t970 486.048
R9138 VPWR.t170 VPWR.t1328 486.048
R9139 VPWR.t1327 VPWR.t1428 486.048
R9140 VPWR.t1633 VPWR.t1326 486.048
R9141 VPWR.t26 VPWR.t901 486.048
R9142 VPWR.t63 VPWR.t1877 486.048
R9143 VPWR.t1881 VPWR.t1530 486.048
R9144 VPWR.t1131 VPWR.t99 486.048
R9145 VPWR.t1721 VPWR.t1072 486.048
R9146 VPWR.t1603 VPWR.t1876 486.048
R9147 VPWR.t1879 VPWR.t1267 486.048
R9148 VPWR.t1689 VPWR.t1878 486.048
R9149 VPWR.t1875 VPWR.t954 486.048
R9150 VPWR.t1111 VPWR.t1874 486.048
R9151 VPWR.t1880 VPWR.t413 486.048
R9152 VPWR.t198 VPWR.t1720 486.048
R9153 VPWR.t1719 VPWR.t495 486.048
R9154 VPWR.t176 VPWR.t102 486.048
R9155 VPWR.t101 VPWR.t1432 486.048
R9156 VPWR.t1639 VPWR.t100 486.048
R9157 VPWR.t1873 VPWR.t880 486.048
R9158 VPWR.t87 VPWR.t1626 486.048
R9159 VPWR.t124 VPWR.t1625 486.048
R9160 VPWR.t1171 VPWR.t84 486.048
R9161 VPWR.t1025 VPWR.t83 486.048
R9162 VPWR.t1575 VPWR.t80 486.048
R9163 VPWR.t1285 VPWR.t1623 486.048
R9164 VPWR.t218 VPWR.t1660 486.048
R9165 VPWR.t1403 VPWR.t79 486.048
R9166 VPWR.t75 VPWR.t78 486.048
R9167 VPWR.t449 VPWR.t1624 486.048
R9168 VPWR.t1731 VPWR.t82 486.048
R9169 VPWR.t1901 VPWR.t81 486.048
R9170 VPWR.t47 VPWR.t1659 486.048
R9171 VPWR.t1581 VPWR.t1658 486.048
R9172 VPWR.t204 VPWR.t1657 486.048
R9173 VPWR.t753 VPWR.t77 486.048
R9174 VPWR.t989 VPWR.t1253 486.048
R9175 VPWR.t1590 VPWR.t1544 486.048
R9176 VPWR.t1914 VPWR.t1139 486.048
R9177 VPWR.t1256 VPWR.t1080 486.048
R9178 VPWR.t1252 VPWR.t111 486.048
R9179 VPWR.t1588 VPWR.t1257 486.048
R9180 VPWR.t1587 VPWR.t1867 486.048
R9181 VPWR.t1251 VPWR.t248 486.048
R9182 VPWR.t1592 VPWR.t318 486.048
R9183 VPWR.t1589 VPWR.t407 486.048
R9184 VPWR.t1255 VPWR.t1747 486.048
R9185 VPWR.t1254 VPWR.t968 486.048
R9186 VPWR.t1711 VPWR.t164 486.048
R9187 VPWR.t1710 VPWR.t1426 486.048
R9188 VPWR.t1915 VPWR.t1627 486.048
R9189 VPWR.t1591 VPWR.t923 486.048
R9190 VPWR.t65 VPWR.t658 486.048
R9191 VPWR.t1532 VPWR.t789 486.048
R9192 VPWR.t1187 VPWR.t918 486.048
R9193 VPWR.t1076 VPWR.t574 486.048
R9194 VPWR.t1605 VPWR.t684 486.048
R9195 VPWR.t839 VPWR.t1762 486.048
R9196 VPWR.t1691 VPWR.t841 486.048
R9197 VPWR.t689 VPWR.t956 486.048
R9198 VPWR.t1113 VPWR.t719 486.048
R9199 VPWR.t837 VPWR.t415 486.048
R9200 VPWR.t588 VPWR.t200 486.048
R9201 VPWR.t607 VPWR.t497 486.048
R9202 VPWR.t851 VPWR.t178 486.048
R9203 VPWR.t1416 VPWR.t869 486.048
R9204 VPWR.t907 VPWR.t1643 486.048
R9205 VPWR.t864 VPWR.t739 486.048
R9206 VPWR.t724 VPWR.t593 486.048
R9207 VPWR.t853 VPWR.t729 486.048
R9208 VPWR.t859 VPWR.t871 486.048
R9209 VPWR.t633 VPWR.t899 486.048
R9210 VPWR.t623 VPWR.t741 486.048
R9211 VPWR.t896 VPWR.t767 486.048
R9212 VPWR.t791 VPWR.t620 486.048
R9213 VPWR.t655 VPWR.t628 486.048
R9214 VPWR.t663 VPWR.t783 486.048
R9215 VPWR.t893 VPWR.t765 486.048
R9216 VPWR.t926 VPWR.t660 486.048
R9217 VPWR.t678 VPWR.t945 486.048
R9218 VPWR.t799 VPWR.t806 486.048
R9219 VPWR.t939 VPWR.t818 486.048
R9220 VPWR.t843 VPWR.t579 486.048
R9221 VPWR.t815 VPWR.t694 486.048
R9222 VPWR.t595 VPWR.t867 486.048
R9223 VPWR.t612 VPWR.t731 486.048
R9224 VPWR.t744 VPWR.t737 486.048
R9225 VPWR.t904 VPWR.t778 486.048
R9226 VPWR.t625 VPWR.t886 486.048
R9227 VPWR.t653 VPWR.t772 486.048
R9228 VPWR.t668 VPWR.t883 486.048
R9229 VPWR.t891 VPWR.t920 486.048
R9230 VPWR.t934 VPWR.t665 486.048
R9231 VPWR.t651 VPWR.t769 486.048
R9232 VPWR.t804 VPWR.t928 486.048
R9233 VPWR.t826 VPWR.t947 486.048
R9234 VPWR.t676 VPWR.t691 486.048
R9235 VPWR.t702 VPWR.t820 486.048
R9236 VPWR.t727 VPWR.t848 486.048
R9237 VPWR.t699 VPWR.t572 486.048
R9238 VPWR.t1677 VPWR.t1476 463.954
R9239 VPWR.t1572 VPWR.t85 463.954
R9240 VPWR.t128 VPWR.t1855 463.954
R9241 VPWR.t1854 VPWR.t1189 463.954
R9242 VPWR.t146 VPWR.t1676 463.954
R9243 VPWR.t1725 VPWR.t1579 463.954
R9244 VPWR.t1289 VPWR.t1724 463.954
R9245 VPWR.t1675 VPWR.t220 463.954
R9246 VPWR.t1384 VPWR.t1574 463.954
R9247 VPWR.t1726 VPWR.t561 463.954
R9248 VPWR.t447 VPWR.t1853 463.954
R9249 VPWR.t1852 VPWR.t1735 463.954
R9250 VPWR.t1899 VPWR.t1723 463.954
R9251 VPWR.t1722 VPWR.t182 463.954
R9252 VPWR.t1206 VPWR.t1856 463.954
R9253 VPWR.t1573 VPWR.t4 463.954
R9254 VPWR.t1911 VPWR.t1465 463.954
R9255 VPWR.t1619 VPWR.t18 463.954
R9256 VPWR.t1712 VPWR.t1846 463.954
R9257 VPWR.t1165 VPWR.t1845 463.954
R9258 VPWR.t1044 VPWR.t1910 463.954
R9259 VPWR.t1526 VPWR.t33 463.954
R9260 VPWR.t1480 VPWR.t32 463.954
R9261 VPWR.t1859 VPWR.t1909 463.954
R9262 VPWR.t499 VPWR.t20 463.954
R9263 VPWR.t1038 VPWR.t34 463.954
R9264 VPWR.t380 VPWR.t1913 463.954
R9265 VPWR.t1512 VPWR.t1912 463.954
R9266 VPWR.t35 VPWR.t31 463.954
R9267 VPWR.t282 VPWR.t30 463.954
R9268 VPWR.t527 VPWR.t1847 463.954
R9269 VPWR.t192 VPWR.t19 463.954
R9270 VPWR.t347 VPWR.t1451 463.954
R9271 VPWR.t557 VPWR.t1683 463.954
R9272 VPWR.t1439 VPWR.t1647 463.954
R9273 VPWR.t1143 VPWR.t1438 463.954
R9274 VPWR.t346 VPWR.t1068 463.954
R9275 VPWR.t1554 VPWR.t1681 463.954
R9276 VPWR.t1680 VPWR.t1496 463.954
R9277 VPWR.t1697 VPWR.t345 463.954
R9278 VPWR.t344 VPWR.t250 463.954
R9279 VPWR.t522 VPWR.t1682 463.954
R9280 VPWR.t1437 VPWR.t435 463.954
R9281 VPWR.t475 VPWR.t1436 463.954
R9282 VPWR.t1679 VPWR.t1441 463.954
R9283 VPWR.t166 VPWR.t1678 463.954
R9284 VPWR.t1440 VPWR.t1568 463.954
R9285 VPWR.t1635 VPWR.t1684 463.954
R9286 VPWR.t433 VPWR.t1459 463.954
R9287 VPWR.t428 VPWR.t983 463.954
R9288 VPWR.t470 VPWR.t1546 463.954
R9289 VPWR.t469 VPWR.t1157 463.954
R9290 VPWR.t432 VPWR.t1050 463.954
R9291 VPWR.t426 VPWR.t113 463.954
R9292 VPWR.t425 VPWR.t1259 463.954
R9293 VPWR.t431 VPWR.t1869 463.954
R9294 VPWR.t430 VPWR.t276 463.954
R9295 VPWR.t427 VPWR.t320 463.954
R9296 VPWR.t468 VPWR.t401 463.954
R9297 VPWR.t434 VPWR.t1749 463.954
R9298 VPWR.t424 VPWR.t962 463.954
R9299 VPWR.t423 VPWR.t290 463.954
R9300 VPWR.t422 VPWR.t1420 463.954
R9301 VPWR.t429 VPWR.t389 463.954
R9302 VPWR.t1089 VPWR.t1471 463.954
R9303 VPWR.t1090 VPWR.t308 463.954
R9304 VPWR.t1607 VPWR.t1517 463.954
R9305 VPWR.t505 VPWR.t1179 463.954
R9306 VPWR.t1027 VPWR.t1088 463.954
R9307 VPWR.t97 VPWR.t1520 463.954
R9308 VPWR.t1271 VPWR.t96 463.954
R9309 VPWR.t1087 VPWR.t230 463.954
R9310 VPWR.t1405 VPWR.t1086 463.954
R9311 VPWR.t98 VPWR.t130 463.954
R9312 VPWR.t356 VPWR.t504 463.954
R9313 VPWR.t503 VPWR.t1118 463.954
R9314 VPWR.t1536 VPWR.t95 463.954
R9315 VPWR.t1519 VPWR.t49 463.954
R9316 VPWR.t485 VPWR.t1518 463.954
R9317 VPWR.t1091 VPWR.t206 463.954
R9318 VPWR.t467 VPWR.t1478 463.954
R9319 VPWR.t1109 VPWR.t1674 463.954
R9320 VPWR.t126 VPWR.t1196 463.954
R9321 VPWR.t1191 VPWR.t1100 463.954
R9322 VPWR.t144 VPWR.t466 463.954
R9323 VPWR.t1577 VPWR.t1672 463.954
R9324 VPWR.t1287 VPWR.t1671 463.954
R9325 VPWR.t952 VPWR.t465 463.954
R9326 VPWR.t958 VPWR.t1097 463.954
R9327 VPWR.t559 VPWR.t1673 463.954
R9328 VPWR.t445 VPWR.t1099 463.954
R9329 VPWR.t1733 VPWR.t1098 463.954
R9330 VPWR.t1897 VPWR.t1199 463.954
R9331 VPWR.t180 VPWR.t1198 463.954
R9332 VPWR.t1204 VPWR.t1197 463.954
R9333 VPWR.t1645 VPWR.t1096 463.954
R9334 VPWR.t1250 VPWR.t1474 463.954
R9335 VPWR.t459 VPWR.t1571 463.954
R9336 VPWR.t1006 VPWR.t510 463.954
R9337 VPWR.t1185 VPWR.t1005 463.954
R9338 VPWR.t1249 VPWR.t148 463.954
R9339 VPWR.t1306 VPWR.t1011 463.954
R9340 VPWR.t1010 VPWR.t1343 463.954
R9341 VPWR.t226 VPWR.t1248 463.954
R9342 VPWR.t1247 VPWR.t1386 463.954
R9343 VPWR.t1221 VPWR.t1570 463.954
R9344 VPWR.t1004 VPWR.t350 463.954
R9345 VPWR.t1848 VPWR.t1003 463.954
R9346 VPWR.t1009 VPWR.t1884 463.954
R9347 VPWR.t39 VPWR.t1008 463.954
R9348 VPWR.t1007 VPWR.t1585 463.954
R9349 VPWR.t6 VPWR.t1246 463.954
R9350 VPWR.t1340 VPWR.t1453 463.954
R9351 VPWR.t1335 VPWR.t555 463.954
R9352 VPWR.t1380 VPWR.t516 463.954
R9353 VPWR.t1379 VPWR.t1145 463.954
R9354 VPWR.t1339 VPWR.t1064 463.954
R9355 VPWR.t1333 VPWR.t1552 463.954
R9356 VPWR.t1332 VPWR.t1494 463.954
R9357 VPWR.t1338 VPWR.t1695 463.954
R9358 VPWR.t1337 VPWR.t246 463.954
R9359 VPWR.t1334 VPWR.t520 463.954
R9360 VPWR.t1378 VPWR.t374 463.954
R9361 VPWR.t1377 VPWR.t473 463.954
R9362 VPWR.t1383 VPWR.t1359 463.954
R9363 VPWR.t1382 VPWR.t162 463.954
R9364 VPWR.t1381 VPWR.t1566 463.954
R9365 VPWR.t1336 VPWR.t1631 463.954
R9366 VPWR.t1002 VPWR.t1469 463.954
R9367 VPWR.t997 VPWR.t310 463.954
R9368 VPWR.t1609 VPWR.t331 463.954
R9369 VPWR.t330 VPWR.t1177 463.954
R9370 VPWR.t1060 VPWR.t1001 463.954
R9371 VPWR.t1904 VPWR.t1522 463.954
R9372 VPWR.t1273 VPWR.t1903 463.954
R9373 VPWR.t1000 VPWR.t232 463.954
R9374 VPWR.t240 VPWR.t999 463.954
R9375 VPWR.t1905 VPWR.t132 463.954
R9376 VPWR.t358 VPWR.t329 463.954
R9377 VPWR.t328 VPWR.t1120 463.954
R9378 VPWR.t1538 VPWR.t334 463.954
R9379 VPWR.t333 VPWR.t51 463.954
R9380 VPWR.t487 VPWR.t332 463.954
R9381 VPWR.t998 VPWR.t208 463.954
R9382 VPWR.t1396 VPWR.t1455 463.954
R9383 VPWR.t553 VPWR.t62 463.954
R9384 VPWR.t514 VPWR.t1919 463.954
R9385 VPWR.t1147 VPWR.t1918 463.954
R9386 VPWR.t1062 VPWR.t1395 463.954
R9387 VPWR.t1699 VPWR.t60 463.954
R9388 VPWR.t1492 VPWR.t59 463.954
R9389 VPWR.t1693 VPWR.t1394 463.954
R9390 VPWR.t268 VPWR.t1393 463.954
R9391 VPWR.t518 VPWR.t61 463.954
R9392 VPWR.t372 VPWR.t1917 463.954
R9393 VPWR.t471 VPWR.t1916 463.954
R9394 VPWR.t1357 VPWR.t58 463.954
R9395 VPWR.t158 VPWR.t57 463.954
R9396 VPWR.t1564 VPWR.t1920 463.954
R9397 VPWR.t1629 VPWR.t1392 463.954
R9398 VPWR.t123 VPWR.t1467 463.954
R9399 VPWR.t980 VPWR.t312 463.954
R9400 VPWR.t1323 VPWR.t1611 463.954
R9401 VPWR.t1322 VPWR.t1173 463.954
R9402 VPWR.t122 VPWR.t1410 463.954
R9403 VPWR.t1704 VPWR.t1524 463.954
R9404 VPWR.t1703 VPWR.t1275 463.954
R9405 VPWR.t121 VPWR.t234 463.954
R9406 VPWR.t120 VPWR.t242 463.954
R9407 VPWR.t1705 VPWR.t134 463.954
R9408 VPWR.t1321 VPWR.t360 463.954
R9409 VPWR.t1320 VPWR.t1122 463.954
R9410 VPWR.t1702 VPWR.t1540 463.954
R9411 VPWR.t1701 VPWR.t53 463.954
R9412 VPWR.t1324 VPWR.t489 463.954
R9413 VPWR.t119 VPWR.t186 463.954
R9414 VPWR.t1921 VPWR.t1461 463.954
R9415 VPWR.t16 VPWR.t25 463.954
R9416 VPWR.t1925 VPWR.t1542 463.954
R9417 VPWR.t1159 VPWR.t1924 463.954
R9418 VPWR.t29 VPWR.t1048 463.954
R9419 VPWR.t109 VPWR.t1330 463.954
R9420 VPWR.t1329 VPWR.t1486 463.954
R9421 VPWR.t1865 VPWR.t28 463.954
R9422 VPWR.t27 VPWR.t274 463.954
R9423 VPWR.t316 VPWR.t1331 463.954
R9424 VPWR.t1923 VPWR.t384 463.954
R9425 VPWR.t1745 VPWR.t1922 463.954
R9426 VPWR.t1328 VPWR.t960 463.954
R9427 VPWR.t288 VPWR.t1327 463.954
R9428 VPWR.t1326 VPWR.t1418 463.954
R9429 VPWR.t196 VPWR.t26 463.954
R9430 VPWR.t1877 VPWR.t1457 463.954
R9431 VPWR.t985 VPWR.t1881 463.954
R9432 VPWR.t99 VPWR.t1548 463.954
R9433 VPWR.t1155 VPWR.t1721 463.954
R9434 VPWR.t1876 VPWR.t1054 463.954
R9435 VPWR.t115 VPWR.t1879 463.954
R9436 VPWR.t1878 VPWR.t1261 463.954
R9437 VPWR.t1871 VPWR.t1875 463.954
R9438 VPWR.t1874 VPWR.t278 463.954
R9439 VPWR.t322 VPWR.t1880 463.954
R9440 VPWR.t1720 VPWR.t403 463.954
R9441 VPWR.t1751 VPWR.t1719 463.954
R9442 VPWR.t102 VPWR.t964 463.954
R9443 VPWR.t292 VPWR.t101 463.954
R9444 VPWR.t100 VPWR.t1422 463.954
R9445 VPWR.t393 VPWR.t1873 463.954
R9446 VPWR.t1626 VPWR.t1449 463.954
R9447 VPWR.t1625 VPWR.t1101 463.954
R9448 VPWR.t84 VPWR.t1653 463.954
R9449 VPWR.t83 VPWR.t1137 463.954
R9450 VPWR.t80 VPWR.t1074 463.954
R9451 VPWR.t1623 VPWR.t1560 463.954
R9452 VPWR.t1660 VPWR.t1502 463.954
R9453 VPWR.t79 VPWR.t214 463.954
R9454 VPWR.t78 VPWR.t254 463.954
R9455 VPWR.t1624 VPWR.t71 463.954
R9456 VPWR.t82 VPWR.t437 463.954
R9457 VPWR.t81 VPWR.t481 463.954
R9458 VPWR.t1659 VPWR.t1443 463.954
R9459 VPWR.t1658 VPWR.t172 463.954
R9460 VPWR.t1657 VPWR.t103 463.954
R9461 VPWR.t77 VPWR.t1641 463.954
R9462 VPWR.t1253 VPWR.t1463 463.954
R9463 VPWR.t1621 VPWR.t1590 463.954
R9464 VPWR.t1714 VPWR.t1914 463.954
R9465 VPWR.t1163 VPWR.t1256 463.954
R9466 VPWR.t1046 VPWR.t1252 463.954
R9467 VPWR.t1528 VPWR.t1588 463.954
R9468 VPWR.t1482 VPWR.t1587 463.954
R9469 VPWR.t1861 VPWR.t1251 463.954
R9470 VPWR.t272 VPWR.t1592 463.954
R9471 VPWR.t1040 VPWR.t1589 463.954
R9472 VPWR.t382 VPWR.t1255 463.954
R9473 VPWR.t1514 VPWR.t1254 463.954
R9474 VPWR.t37 VPWR.t1711 463.954
R9475 VPWR.t286 VPWR.t1710 463.954
R9476 VPWR.t529 VPWR.t1915 463.954
R9477 VPWR.t194 VPWR.t1591 463.954
R9478 VPWR.t658 VPWR.t673 463.954
R9479 VPWR.t789 VPWR.t834 463.954
R9480 VPWR.t918 VPWR.t936 463.954
R9481 VPWR.t574 VPWR.t707 463.954
R9482 VPWR.t684 VPWR.t809 463.954
R9483 VPWR.t831 VPWR.t839 463.954
R9484 VPWR.t841 VPWR.t582 463.954
R9485 VPWR.t704 VPWR.t689 463.954
R9486 VPWR.t719 VPWR.t845 463.954
R9487 VPWR.t861 VPWR.t837 463.954
R9488 VPWR.t604 VPWR.t588 463.954
R9489 VPWR.t734 VPWR.t607 463.954
R9490 VPWR.t775 VPWR.t851 463.954
R9491 VPWR.t869 VPWR.t598 463.954
R9492 VPWR.t648 VPWR.t907 463.954
R9493 VPWR.t739 VPWR.t756 463.954
R9494 VPWR.t593 VPWR.t617 463.954
R9495 VPWR.t729 VPWR.t762 463.954
R9496 VPWR.t874 VPWR.t859 463.954
R9497 VPWR.t899 VPWR.t639 463.954
R9498 VPWR.t750 VPWR.t623 463.954
R9499 VPWR.t767 VPWR.t759 463.954
R9500 VPWR.t915 VPWR.t791 463.954
R9501 VPWR.t628 VPWR.t636 463.954
R9502 VPWR.t796 VPWR.t663 463.954
R9503 VPWR.t765 VPWR.t812 463.954
R9504 VPWR.t942 VPWR.t926 463.954
R9505 VPWR.t945 VPWR.t686 463.954
R9506 VPWR.t716 VPWR.t799 463.954
R9507 VPWR.t818 VPWR.t566 463.954
R9508 VPWR.t585 VPWR.t843 463.954
R9509 VPWR.t694 VPWR.t710 463.954
R9510 VPWR.t867 VPWR.t877 463.954
R9511 VPWR.t645 VPWR.t612 463.954
R9512 VPWR.t737 VPWR.t747 463.954
R9513 VPWR.t778 VPWR.t912 463.954
R9514 VPWR.t886 VPWR.t630 463.954
R9515 VPWR.t642 VPWR.t653 463.954
R9516 VPWR.t801 VPWR.t668 463.954
R9517 VPWR.t909 VPWR.t891 463.954
R9518 VPWR.t670 VPWR.t934 463.954
R9519 VPWR.t696 VPWR.t651 463.954
R9520 VPWR.t823 VPWR.t804 463.954
R9521 VPWR.t569 VPWR.t826 463.954
R9522 VPWR.t590 VPWR.t676 463.954
R9523 VPWR.t828 VPWR.t702 463.954
R9524 VPWR.t856 VPWR.t727 463.954
R9525 VPWR.t572 VPWR.t576 463.954
R9526 VPWR.n2626 VPWR.t539 428.822
R9527 VPWR.n1595 VPWR.n1594 376.045
R9528 VPWR.n2506 VPWR.n2505 376.045
R9529 VPWR.n1468 VPWR.n1467 376.045
R9530 VPWR.n351 VPWR.n350 376.045
R9531 VPWR.n2568 VPWR.n2567 376.045
R9532 VPWR.n1535 VPWR.n1534 376.045
R9533 VPWR.n349 VPWR.n348 376.045
R9534 VPWR.n2508 VPWR.n2507 376.045
R9535 VPWR.n966 VPWR.n965 376.045
R9536 VPWR.n2478 VPWR.n2477 376.045
R9537 VPWR.n2476 VPWR.n2475 376.045
R9538 VPWR.n321 VPWR.n320 376.045
R9539 VPWR.n2554 VPWR.n2553 376.045
R9540 VPWR.n974 VPWR.n973 376.045
R9541 VPWR.n2446 VPWR.n2445 376.045
R9542 VPWR.n325 VPWR.n324 376.045
R9543 VPWR.n2544 VPWR.n2543 376.045
R9544 VPWR.n1890 VPWR.n1889 376.045
R9545 VPWR.n1888 VPWR.n1887 376.045
R9546 VPWR.n1880 VPWR.n1879 376.045
R9547 VPWR.n390 VPWR.n389 376.045
R9548 VPWR.n394 VPWR.n393 376.045
R9549 VPWR.n398 VPWR.n397 376.045
R9550 VPWR.n2456 VPWR.n2455 376.045
R9551 VPWR.n333 VPWR.n332 376.045
R9552 VPWR.n2532 VPWR.n2531 376.045
R9553 VPWR.n1878 VPWR.n1877 376.045
R9554 VPWR.n406 VPWR.n405 376.045
R9555 VPWR.n2458 VPWR.n2457 376.045
R9556 VPWR.n337 VPWR.n336 376.045
R9557 VPWR.n2530 VPWR.n2529 376.045
R9558 VPWR.n2309 VPWR.n2308 376.045
R9559 VPWR.n2311 VPWR.n2310 376.045
R9560 VPWR.n2319 VPWR.n2318 376.045
R9561 VPWR.n2321 VPWR.n2320 376.045
R9562 VPWR.n2331 VPWR.n2330 376.045
R9563 VPWR.n2339 VPWR.n2338 376.045
R9564 VPWR.n2341 VPWR.n2340 376.045
R9565 VPWR.n2349 VPWR.n2348 376.045
R9566 VPWR.n2351 VPWR.n2350 376.045
R9567 VPWR.n2359 VPWR.n2358 376.045
R9568 VPWR.n2361 VPWR.n2360 376.045
R9569 VPWR.n2369 VPWR.n2368 376.045
R9570 VPWR.n2371 VPWR.n2370 376.045
R9571 VPWR.n2379 VPWR.n2378 376.045
R9572 VPWR.n2329 VPWR.n2328 376.045
R9573 VPWR.n543 VPWR.n542 376.045
R9574 VPWR.n541 VPWR.n540 376.045
R9575 VPWR.n537 VPWR.n536 376.045
R9576 VPWR.n533 VPWR.n532 376.045
R9577 VPWR.n525 VPWR.n524 376.045
R9578 VPWR.n521 VPWR.n520 376.045
R9579 VPWR.n517 VPWR.n516 376.045
R9580 VPWR.n513 VPWR.n512 376.045
R9581 VPWR.n509 VPWR.n508 376.045
R9582 VPWR.n505 VPWR.n504 376.045
R9583 VPWR.n501 VPWR.n500 376.045
R9584 VPWR.n497 VPWR.n496 376.045
R9585 VPWR.n493 VPWR.n492 376.045
R9586 VPWR.n489 VPWR.n488 376.045
R9587 VPWR.n529 VPWR.n528 376.045
R9588 VPWR.n2282 VPWR.n2281 376.045
R9589 VPWR.n2280 VPWR.n2279 376.045
R9590 VPWR.n2272 VPWR.n2271 376.045
R9591 VPWR.n2270 VPWR.n2269 376.045
R9592 VPWR.n2260 VPWR.n2259 376.045
R9593 VPWR.n2252 VPWR.n2251 376.045
R9594 VPWR.n2250 VPWR.n2249 376.045
R9595 VPWR.n2242 VPWR.n2241 376.045
R9596 VPWR.n2240 VPWR.n2239 376.045
R9597 VPWR.n2232 VPWR.n2231 376.045
R9598 VPWR.n2230 VPWR.n2229 376.045
R9599 VPWR.n2222 VPWR.n2221 376.045
R9600 VPWR.n2220 VPWR.n2219 376.045
R9601 VPWR.n2212 VPWR.n2211 376.045
R9602 VPWR.n2262 VPWR.n2261 376.045
R9603 VPWR.n582 VPWR.n581 376.045
R9604 VPWR.n586 VPWR.n585 376.045
R9605 VPWR.n590 VPWR.n589 376.045
R9606 VPWR.n594 VPWR.n593 376.045
R9607 VPWR.n602 VPWR.n601 376.045
R9608 VPWR.n606 VPWR.n605 376.045
R9609 VPWR.n610 VPWR.n609 376.045
R9610 VPWR.n614 VPWR.n613 376.045
R9611 VPWR.n618 VPWR.n617 376.045
R9612 VPWR.n622 VPWR.n621 376.045
R9613 VPWR.n626 VPWR.n625 376.045
R9614 VPWR.n630 VPWR.n629 376.045
R9615 VPWR.n634 VPWR.n633 376.045
R9616 VPWR.n638 VPWR.n637 376.045
R9617 VPWR.n598 VPWR.n597 376.045
R9618 VPWR.n2113 VPWR.n2112 376.045
R9619 VPWR.n2115 VPWR.n2114 376.045
R9620 VPWR.n2123 VPWR.n2122 376.045
R9621 VPWR.n2125 VPWR.n2124 376.045
R9622 VPWR.n2135 VPWR.n2134 376.045
R9623 VPWR.n2143 VPWR.n2142 376.045
R9624 VPWR.n2145 VPWR.n2144 376.045
R9625 VPWR.n2153 VPWR.n2152 376.045
R9626 VPWR.n2155 VPWR.n2154 376.045
R9627 VPWR.n2163 VPWR.n2162 376.045
R9628 VPWR.n2165 VPWR.n2164 376.045
R9629 VPWR.n2173 VPWR.n2172 376.045
R9630 VPWR.n2175 VPWR.n2174 376.045
R9631 VPWR.n2183 VPWR.n2182 376.045
R9632 VPWR.n2133 VPWR.n2132 376.045
R9633 VPWR.n735 VPWR.n734 376.045
R9634 VPWR.n733 VPWR.n732 376.045
R9635 VPWR.n729 VPWR.n728 376.045
R9636 VPWR.n725 VPWR.n724 376.045
R9637 VPWR.n717 VPWR.n716 376.045
R9638 VPWR.n713 VPWR.n712 376.045
R9639 VPWR.n709 VPWR.n708 376.045
R9640 VPWR.n705 VPWR.n704 376.045
R9641 VPWR.n701 VPWR.n700 376.045
R9642 VPWR.n697 VPWR.n696 376.045
R9643 VPWR.n693 VPWR.n692 376.045
R9644 VPWR.n689 VPWR.n688 376.045
R9645 VPWR.n685 VPWR.n684 376.045
R9646 VPWR.n681 VPWR.n680 376.045
R9647 VPWR.n721 VPWR.n720 376.045
R9648 VPWR.n2086 VPWR.n2085 376.045
R9649 VPWR.n2084 VPWR.n2083 376.045
R9650 VPWR.n2076 VPWR.n2075 376.045
R9651 VPWR.n2074 VPWR.n2073 376.045
R9652 VPWR.n2064 VPWR.n2063 376.045
R9653 VPWR.n2056 VPWR.n2055 376.045
R9654 VPWR.n2054 VPWR.n2053 376.045
R9655 VPWR.n2046 VPWR.n2045 376.045
R9656 VPWR.n2044 VPWR.n2043 376.045
R9657 VPWR.n2036 VPWR.n2035 376.045
R9658 VPWR.n2034 VPWR.n2033 376.045
R9659 VPWR.n2026 VPWR.n2025 376.045
R9660 VPWR.n2024 VPWR.n2023 376.045
R9661 VPWR.n2016 VPWR.n2015 376.045
R9662 VPWR.n2066 VPWR.n2065 376.045
R9663 VPWR.n774 VPWR.n773 376.045
R9664 VPWR.n778 VPWR.n777 376.045
R9665 VPWR.n782 VPWR.n781 376.045
R9666 VPWR.n786 VPWR.n785 376.045
R9667 VPWR.n794 VPWR.n793 376.045
R9668 VPWR.n798 VPWR.n797 376.045
R9669 VPWR.n802 VPWR.n801 376.045
R9670 VPWR.n806 VPWR.n805 376.045
R9671 VPWR.n810 VPWR.n809 376.045
R9672 VPWR.n814 VPWR.n813 376.045
R9673 VPWR.n818 VPWR.n817 376.045
R9674 VPWR.n822 VPWR.n821 376.045
R9675 VPWR.n826 VPWR.n825 376.045
R9676 VPWR.n830 VPWR.n829 376.045
R9677 VPWR.n790 VPWR.n789 376.045
R9678 VPWR.n1917 VPWR.n1916 376.045
R9679 VPWR.n1919 VPWR.n1918 376.045
R9680 VPWR.n1927 VPWR.n1926 376.045
R9681 VPWR.n1929 VPWR.n1928 376.045
R9682 VPWR.n1939 VPWR.n1938 376.045
R9683 VPWR.n1947 VPWR.n1946 376.045
R9684 VPWR.n1949 VPWR.n1948 376.045
R9685 VPWR.n1957 VPWR.n1956 376.045
R9686 VPWR.n1959 VPWR.n1958 376.045
R9687 VPWR.n1967 VPWR.n1966 376.045
R9688 VPWR.n1969 VPWR.n1968 376.045
R9689 VPWR.n1977 VPWR.n1976 376.045
R9690 VPWR.n1979 VPWR.n1978 376.045
R9691 VPWR.n1987 VPWR.n1986 376.045
R9692 VPWR.n1937 VPWR.n1936 376.045
R9693 VPWR.n927 VPWR.n926 376.045
R9694 VPWR.n925 VPWR.n924 376.045
R9695 VPWR.n921 VPWR.n920 376.045
R9696 VPWR.n917 VPWR.n916 376.045
R9697 VPWR.n909 VPWR.n908 376.045
R9698 VPWR.n905 VPWR.n904 376.045
R9699 VPWR.n901 VPWR.n900 376.045
R9700 VPWR.n897 VPWR.n896 376.045
R9701 VPWR.n893 VPWR.n892 376.045
R9702 VPWR.n889 VPWR.n888 376.045
R9703 VPWR.n885 VPWR.n884 376.045
R9704 VPWR.n881 VPWR.n880 376.045
R9705 VPWR.n877 VPWR.n876 376.045
R9706 VPWR.n873 VPWR.n872 376.045
R9707 VPWR.n913 VPWR.n912 376.045
R9708 VPWR.n1870 VPWR.n1869 376.045
R9709 VPWR.n982 VPWR.n981 376.045
R9710 VPWR.n1494 VPWR.n1493 376.045
R9711 VPWR.n1221 VPWR.n1220 376.045
R9712 VPWR.n402 VPWR.n401 376.045
R9713 VPWR.n2466 VPWR.n2465 376.045
R9714 VPWR.n341 VPWR.n340 376.045
R9715 VPWR.n2520 VPWR.n2519 376.045
R9716 VPWR.n978 VPWR.n977 376.045
R9717 VPWR.n1492 VPWR.n1491 376.045
R9718 VPWR.n1185 VPWR.n1184 376.045
R9719 VPWR.n1868 VPWR.n1867 376.045
R9720 VPWR.n986 VPWR.n985 376.045
R9721 VPWR.n1506 VPWR.n1505 376.045
R9722 VPWR.n1219 VPWR.n1218 376.045
R9723 VPWR.n410 VPWR.n409 376.045
R9724 VPWR.n418 VPWR.n417 376.045
R9725 VPWR.n422 VPWR.n421 376.045
R9726 VPWR.n426 VPWR.n425 376.045
R9727 VPWR.n430 VPWR.n429 376.045
R9728 VPWR.n434 VPWR.n433 376.045
R9729 VPWR.n438 VPWR.n437 376.045
R9730 VPWR.n442 VPWR.n441 376.045
R9731 VPWR.n446 VPWR.n445 376.045
R9732 VPWR.n414 VPWR.n413 376.045
R9733 VPWR.n2448 VPWR.n2447 376.045
R9734 VPWR.n329 VPWR.n328 376.045
R9735 VPWR.n2542 VPWR.n2541 376.045
R9736 VPWR.n990 VPWR.n989 376.045
R9737 VPWR.n1508 VPWR.n1507 376.045
R9738 VPWR.n1216 VPWR.n1215 376.045
R9739 VPWR.n1860 VPWR.n1859 376.045
R9740 VPWR.n1850 VPWR.n1849 376.045
R9741 VPWR.n1848 VPWR.n1847 376.045
R9742 VPWR.n1840 VPWR.n1839 376.045
R9743 VPWR.n1838 VPWR.n1837 376.045
R9744 VPWR.n1830 VPWR.n1829 376.045
R9745 VPWR.n1828 VPWR.n1827 376.045
R9746 VPWR.n1820 VPWR.n1819 376.045
R9747 VPWR.n1858 VPWR.n1857 376.045
R9748 VPWR.n994 VPWR.n993 376.045
R9749 VPWR.n1520 VPWR.n1519 376.045
R9750 VPWR.n1213 VPWR.n1212 376.045
R9751 VPWR.n2468 VPWR.n2467 376.045
R9752 VPWR.n345 VPWR.n344 376.045
R9753 VPWR.n2518 VPWR.n2517 376.045
R9754 VPWR.n1481 VPWR.n1480 376.045
R9755 VPWR.n1182 VPWR.n1181 376.045
R9756 VPWR.n998 VPWR.n997 376.045
R9757 VPWR.n1522 VPWR.n1521 376.045
R9758 VPWR.n1205 VPWR.n1204 376.045
R9759 VPWR.n2438 VPWR.n2437 376.045
R9760 VPWR.n2428 VPWR.n2427 376.045
R9761 VPWR.n2426 VPWR.n2425 376.045
R9762 VPWR.n2418 VPWR.n2417 376.045
R9763 VPWR.n2416 VPWR.n2415 376.045
R9764 VPWR.n2408 VPWR.n2407 376.045
R9765 VPWR.n2436 VPWR.n2435 376.045
R9766 VPWR.n317 VPWR.n316 376.045
R9767 VPWR.n2556 VPWR.n2555 376.045
R9768 VPWR.n1537 VPWR.n1536 376.045
R9769 VPWR.n1202 VPWR.n1201 376.045
R9770 VPWR.n1002 VPWR.n1001 376.045
R9771 VPWR.n1006 VPWR.n1005 376.045
R9772 VPWR.n1010 VPWR.n1009 376.045
R9773 VPWR.n1014 VPWR.n1013 376.045
R9774 VPWR.n1018 VPWR.n1017 376.045
R9775 VPWR.n1022 VPWR.n1021 376.045
R9776 VPWR.n970 VPWR.n969 376.045
R9777 VPWR.n1475 VPWR.n1474 376.045
R9778 VPWR.n1593 VPWR.n1592 376.045
R9779 VPWR.n313 VPWR.n312 376.045
R9780 VPWR.n2566 VPWR.n2565 376.045
R9781 VPWR.n1199 VPWR.n1198 376.045
R9782 VPWR.n1762 VPWR.n1761 376.045
R9783 VPWR.n1191 VPWR.n1190 376.045
R9784 VPWR.n309 VPWR.n308 376.045
R9785 VPWR.n305 VPWR.n304 376.045
R9786 VPWR.n297 VPWR.n296 376.045
R9787 VPWR.n301 VPWR.n300 376.045
R9788 VPWR.n1741 VPWR.n1740 376.045
R9789 VPWR.n1750 VPWR.n1749 376.045
R9790 VPWR.n1791 VPWR.n1790 376.045
R9791 VPWR.n1760 VPWR.n1759 376.045
R9792 VPWR.n1188 VPWR.n1187 376.045
R9793 VPWR.n2578 VPWR.n2577 376.045
R9794 VPWR.n2580 VPWR.n2579 376.045
R9795 VPWR.n2590 VPWR.n2589 376.045
R9796 VPWR.n1739 VPWR.n1738 376.045
R9797 VPWR.n1339 VPWR.t1718 342.841
R9798 VPWR.n1378 VPWR.t337 342.841
R9799 VPWR.n1415 VPWR.t1353 342.841
R9800 VPWR.n2693 VPWR.t1227 342.841
R9801 VPWR.n2656 VPWR.t1235 342.841
R9802 VPWR.n2599 VPWR.t1017 342.841
R9803 VPWR.n1339 VPWR.t1599 342.839
R9804 VPWR.n1378 VPWR.t156 342.839
R9805 VPWR.n1415 VPWR.t1032 342.839
R9806 VPWR.n2693 VPWR.t1666 342.839
R9807 VPWR.n2656 VPWR.t1489 342.839
R9808 VPWR.n2599 VPWR.t540 342.839
R9809 VPWR.n2842 VPWR.n2824 339.212
R9810 VPWR.n1306 VPWR.t1730 338.488
R9811 VPWR.n2729 VPWR.t1366 338.488
R9812 VPWR.n1315 VPWR.n1314 327.377
R9813 VPWR.n1308 VPWR.n1307 327.377
R9814 VPWR.n1322 VPWR.n1321 327.377
R9815 VPWR.n1352 VPWR.n1350 327.377
R9816 VPWR.n1345 VPWR.n1343 327.377
R9817 VPWR.n1360 VPWR.n1358 327.377
R9818 VPWR.n1391 VPWR.n1389 327.377
R9819 VPWR.n1384 VPWR.n1382 327.377
R9820 VPWR.n1399 VPWR.n1397 327.377
R9821 VPWR.n1428 VPWR.n1426 327.377
R9822 VPWR.n1421 VPWR.n1419 327.377
R9823 VPWR.n1436 VPWR.n1434 327.377
R9824 VPWR.n1324 VPWR.n1323 327.375
R9825 VPWR.n1352 VPWR.n1351 327.375
R9826 VPWR.n1345 VPWR.n1344 327.375
R9827 VPWR.n1360 VPWR.n1359 327.375
R9828 VPWR.n1391 VPWR.n1390 327.375
R9829 VPWR.n1384 VPWR.n1383 327.375
R9830 VPWR.n1399 VPWR.n1398 327.375
R9831 VPWR.n1428 VPWR.n1427 327.375
R9832 VPWR.n1421 VPWR.n1420 327.375
R9833 VPWR.n1436 VPWR.n1435 327.375
R9834 VPWR.n1 VPWR 325.546
R9835 VPWR.n2667 VPWR.t1226 322.262
R9836 VPWR.n2630 VPWR.t1234 322.262
R9837 VPWR.n2805 VPWR.n2804 321.642
R9838 VPWR.n2722 VPWR.n2712 320.976
R9839 VPWR.n2716 VPWR.n2715 320.976
R9840 VPWR.n2710 VPWR.n2709 320.976
R9841 VPWR.n2680 VPWR.n2679 320.976
R9842 VPWR.n2686 VPWR.n2675 320.976
R9843 VPWR.n2672 VPWR.n2671 320.976
R9844 VPWR.n2643 VPWR.n2642 320.976
R9845 VPWR.n2649 VPWR.n2638 320.976
R9846 VPWR.n2635 VPWR.n2634 320.976
R9847 VPWR.n2610 VPWR.n2606 320.976
R9848 VPWR.n2614 VPWR.n2613 320.976
R9849 VPWR.n2620 VPWR.n2602 320.976
R9850 VPWR.n2727 VPWR.n2708 320.976
R9851 VPWR.n2680 VPWR.n2678 320.976
R9852 VPWR.n2686 VPWR.n2674 320.976
R9853 VPWR.n2672 VPWR.n2670 320.976
R9854 VPWR.n2643 VPWR.n2641 320.976
R9855 VPWR.n2649 VPWR.n2637 320.976
R9856 VPWR.n2635 VPWR.n2633 320.976
R9857 VPWR.n2610 VPWR.n2605 320.976
R9858 VPWR.n2614 VPWR.n2612 320.976
R9859 VPWR.n2620 VPWR.n2601 320.976
R9860 VPWR.n2801 VPWR 319.627
R9861 VPWR.n6 VPWR.n5 316.245
R9862 VPWR.n1241 VPWR.n1239 316.245
R9863 VPWR.n1264 VPWR.n1262 316.245
R9864 VPWR.n1288 VPWR.n1286 316.245
R9865 VPWR.n2784 VPWR.n2783 316.245
R9866 VPWR.n2764 VPWR.n2763 316.245
R9867 VPWR.n2745 VPWR.n2744 316.245
R9868 VPWR.n1241 VPWR.n1240 316.245
R9869 VPWR.n1264 VPWR.n1263 316.245
R9870 VPWR.n1288 VPWR.n1287 316.245
R9871 VPWR.n2784 VPWR.n2782 316.245
R9872 VPWR.n2764 VPWR.n2762 316.245
R9873 VPWR.n2745 VPWR.n2743 316.245
R9874 VPWR.n2630 VPWR.t525 313.87
R9875 VPWR.n10 VPWR.n4 310.502
R9876 VPWR.n1246 VPWR.n1238 310.502
R9877 VPWR.n1269 VPWR.n1261 310.502
R9878 VPWR.n1293 VPWR.n1285 310.502
R9879 VPWR.n2803 VPWR.n2802 310.502
R9880 VPWR.n2788 VPWR.n2787 310.502
R9881 VPWR.n2768 VPWR.n2767 310.502
R9882 VPWR.n2749 VPWR.n2748 310.502
R9883 VPWR.n1246 VPWR.n1245 310.5
R9884 VPWR.n1269 VPWR.n1268 310.5
R9885 VPWR.n1293 VPWR.n1292 310.5
R9886 VPWR.n2788 VPWR.n2786 310.5
R9887 VPWR.n2768 VPWR.n2766 310.5
R9888 VPWR.n2749 VPWR.n2747 310.5
R9889 VPWR.n2834 VPWR.n2833 279.341
R9890 VPWR.n2839 VPWR.n2838 279.341
R9891 VPWR.n1412 VPWR.t1225 255.905
R9892 VPWR.n2663 VPWR.t526 255.905
R9893 VPWR.n1275 VPWR.t1130 255.904
R9894 VPWR.n1412 VPWR.t1 255.904
R9895 VPWR.n2774 VPWR.t1215 255.904
R9896 VPWR.n2663 VPWR.t1012 255.904
R9897 VPWR.n1303 VPWR.t979 254.019
R9898 VPWR.n2735 VPWR.t1894 254.019
R9899 VPWR.n1335 VPWR.t977 252.948
R9900 VPWR.n2737 VPWR.t1892 252.948
R9901 VPWR.n1373 VPWR.t1906 250.722
R9902 VPWR.n2700 VPWR.t1742 250.722
R9903 VPWR.n1310 VPWR.t304 249.901
R9904 VPWR.n1346 VPWR.t368 249.901
R9905 VPWR.n1385 VPWR.t1310 249.901
R9906 VPWR.n1422 VPWR.t371 249.901
R9907 VPWR.n2714 VPWR.t1819 249.901
R9908 VPWR.n2677 VPWR.t1816 249.901
R9909 VPWR.n2640 VPWR.t1830 249.901
R9910 VPWR.n2607 VPWR.t1784 249.901
R9911 VPWR.n1346 VPWR.t1295 249.901
R9912 VPWR.n1385 VPWR.t421 249.901
R9913 VPWR.n1422 VPWR.t1117 249.901
R9914 VPWR.n2677 VPWR.t1829 249.901
R9915 VPWR.n2640 VPWR.t1782 249.901
R9916 VPWR.n2607 VPWR.t1805 249.901
R9917 VPWR.n1253 VPWR.t1739 249.363
R9918 VPWR.n1338 VPWR.t949 249.363
R9919 VPWR.n2811 VPWR.t13 249.363
R9920 VPWR.n2795 VPWR.t1389 249.363
R9921 VPWR.n2698 VPWR.t458 249.363
R9922 VPWR.n17 VPWR.t1838 249.362
R9923 VPWR.n1253 VPWR.t1208 249.362
R9924 VPWR.n2795 VPWR.t1662 249.362
R9925 VPWR.t1126 VPWR.t1837 248.599
R9926 VPWR.t1727 VPWR.t258 248.599
R9927 VPWR.t258 VPWR.t262 248.599
R9928 VPWR.t262 VPWR.t140 248.599
R9929 VPWR.t140 VPWR.t1325 248.599
R9930 VPWR.t1325 VPWR.t1759 248.599
R9931 VPWR.t1759 VPWR.t366 248.599
R9932 VPWR.t366 VPWR.t387 248.599
R9933 VPWR.t1766 VPWR.t1293 248.599
R9934 VPWR.t1293 VPWR.t303 248.599
R9935 VPWR.t1832 VPWR.t1808 248.599
R9936 VPWR.t1796 VPWR.t1832 248.599
R9937 VPWR.t1770 VPWR.t1796 248.599
R9938 VPWR.t1367 VPWR.t1770 248.599
R9939 VPWR.t1361 VPWR.t1367 248.599
R9940 VPWR.t1373 VPWR.t1361 248.599
R9941 VPWR.t1375 VPWR.t1373 248.599
R9942 VPWR.t1216 VPWR.t12 248.599
R9943 VPWR.t1776 VPWR.t1818 248.599
R9944 VPWR.t1824 VPWR.t1776 248.599
R9945 VPWR.n15 VPWR.t1127 247.394
R9946 VPWR.n1251 VPWR.t1129 247.394
R9947 VPWR.n2809 VPWR.t1217 247.394
R9948 VPWR.n2793 VPWR.t1211 247.394
R9949 VPWR.n1251 VPWR.t1128 247.394
R9950 VPWR.n2793 VPWR.t1213 247.394
R9951 VPWR.n1304 VPWR.t307 244.737
R9952 VPWR.n2730 VPWR.t1834 244.737
R9953 VPWR.n1374 VPWR.t1516 243.886
R9954 VPWR.n2701 VPWR.t1908 243.886
R9955 VPWR.n1277 VPWR.t1836 243.512
R9956 VPWR.n1300 VPWR.t1740 243.512
R9957 VPWR.n1303 VPWR.t951 243.512
R9958 VPWR.n2776 VPWR.t15 243.512
R9959 VPWR.n2756 VPWR.t1391 243.512
R9960 VPWR.n2735 VPWR.t456 243.512
R9961 VPWR.n1300 VPWR.t1209 243.512
R9962 VPWR.n2756 VPWR.t1661 243.512
R9963 VPWR.n1329 VPWR.t978 238.339
R9964 VPWR.n2705 VPWR.t1893 238.339
R9965 VPWR.n2855 VPWR.t266 237.99
R9966 VPWR.n2667 VPWR.t457 234.982
R9967 VPWR.t1764 VPWR.t1766 228.101
R9968 VPWR.t1802 VPWR.t1824 228.101
R9969 VPWR.n2801 VPWR 224.923
R9970 VPWR.n1 VPWR 219.004
R9971 VPWR.n1444 VPWR.n1443 214.613
R9972 VPWR.n1444 VPWR.n1442 214.613
R9973 VPWR.n1236 VPWR.n1235 214.326
R9974 VPWR.n1259 VPWR.n1258 214.326
R9975 VPWR.n1283 VPWR.n1282 214.326
R9976 VPWR.n1368 VPWR.n1367 214.326
R9977 VPWR.n1407 VPWR.n1406 214.326
R9978 VPWR.n1236 VPWR.n1234 214.326
R9979 VPWR.n1259 VPWR.n1257 214.326
R9980 VPWR.n1283 VPWR.n1281 214.326
R9981 VPWR.n1368 VPWR.n1366 214.326
R9982 VPWR.n1407 VPWR.n1405 214.326
R9983 VPWR.n2 VPWR.n1 213.119
R9984 VPWR.n2808 VPWR.n2801 213.119
R9985 VPWR VPWR.t1126 207.166
R9986 VPWR.n2840 VPWR.n2839 204.424
R9987 VPWR.n2830 VPWR.n2817 204.424
R9988 VPWR.n2833 VPWR.n2820 204.424
R9989 VPWR.n2844 VPWR.n2841 204.048
R9990 VPWR VPWR.t1375 201.246
R9991 VPWR.t303 VPWR 189.409
R9992 VPWR.n2741 VPWR 184.63
R9993 VPWR.n1329 VPWR 182.952
R9994 VPWR.n2760 VPWR 182.952
R9995 VPWR.n2780 VPWR 181.273
R9996 VPWR.t525 VPWR 177.916
R9997 VPWR.n2848 VPWR.n2847 166.4
R9998 VPWR.n1770 VPWR.n1768 161.365
R9999 VPWR.n1041 VPWR.n1039 161.365
R10000 VPWR.n1545 VPWR.n1543 161.365
R10001 VPWR.n1550 VPWR.n1548 161.365
R10002 VPWR.n1555 VPWR.n1553 161.365
R10003 VPWR.n1560 VPWR.n1558 161.365
R10004 VPWR.n1565 VPWR.n1563 161.365
R10005 VPWR.n1570 VPWR.n1568 161.365
R10006 VPWR.n1575 VPWR.n1573 161.365
R10007 VPWR.n1580 VPWR.n1578 161.365
R10008 VPWR.n1135 VPWR.n1133 161.365
R10009 VPWR.n1460 VPWR.n1458 161.365
R10010 VPWR.n1455 VPWR.n1453 161.365
R10011 VPWR.n1775 VPWR.n1773 161.365
R10012 VPWR.n1783 VPWR.n1781 161.365
R10013 VPWR.n1779 VPWR.n1777 161.365
R10014 VPWR VPWR.n53 161.363
R10015 VPWR VPWR.n51 161.363
R10016 VPWR VPWR.n49 161.363
R10017 VPWR VPWR.n47 161.363
R10018 VPWR VPWR.n45 161.363
R10019 VPWR VPWR.n43 161.363
R10020 VPWR VPWR.n41 161.363
R10021 VPWR VPWR.n39 161.363
R10022 VPWR VPWR.n37 161.363
R10023 VPWR VPWR.n35 161.363
R10024 VPWR VPWR.n33 161.363
R10025 VPWR VPWR.n31 161.363
R10026 VPWR VPWR.n29 161.363
R10027 VPWR VPWR.n27 161.363
R10028 VPWR VPWR.n25 161.363
R10029 VPWR VPWR.n23 161.363
R10030 VPWR.n1115 VPWR.n1114 161.303
R10031 VPWR.n107 VPWR.n106 161.303
R10032 VPWR.n1120 VPWR.n1119 161.3
R10033 VPWR.n1599 VPWR.n1598 161.3
R10034 VPWR.n1602 VPWR.n1601 161.3
R10035 VPWR.n1111 VPWR.n1110 161.3
R10036 VPWR.n1126 VPWR.n1125 161.3
R10037 VPWR.n1107 VPWR.n1106 161.3
R10038 VPWR.n1612 VPWR.n1611 161.3
R10039 VPWR.n1615 VPWR.n1614 161.3
R10040 VPWR.n1618 VPWR.n1617 161.3
R10041 VPWR.n1623 VPWR.n1622 161.3
R10042 VPWR.n1626 VPWR.n1625 161.3
R10043 VPWR.n1629 VPWR.n1628 161.3
R10044 VPWR.n1101 VPWR.n1100 161.3
R10045 VPWR.n1177 VPWR.n1176 161.3
R10046 VPWR.n1097 VPWR.n1096 161.3
R10047 VPWR.n1639 VPWR.n1638 161.3
R10048 VPWR.n1642 VPWR.n1641 161.3
R10049 VPWR.n1645 VPWR.n1644 161.3
R10050 VPWR.n1650 VPWR.n1649 161.3
R10051 VPWR.n1653 VPWR.n1652 161.3
R10052 VPWR.n1656 VPWR.n1655 161.3
R10053 VPWR.n1091 VPWR.n1090 161.3
R10054 VPWR.n1209 VPWR.n1208 161.3
R10055 VPWR.n1087 VPWR.n1086 161.3
R10056 VPWR.n1666 VPWR.n1665 161.3
R10057 VPWR.n1669 VPWR.n1668 161.3
R10058 VPWR.n1672 VPWR.n1671 161.3
R10059 VPWR.n1677 VPWR.n1676 161.3
R10060 VPWR.n1680 VPWR.n1679 161.3
R10061 VPWR.n1683 VPWR.n1682 161.3
R10062 VPWR.n1081 VPWR.n1080 161.3
R10063 VPWR.n1195 VPWR.n1194 161.3
R10064 VPWR.n1077 VPWR.n1076 161.3
R10065 VPWR.n1693 VPWR.n1692 161.3
R10066 VPWR.n1696 VPWR.n1695 161.3
R10067 VPWR.n1699 VPWR.n1698 161.3
R10068 VPWR.n1704 VPWR.n1703 161.3
R10069 VPWR.n1707 VPWR.n1706 161.3
R10070 VPWR.n1710 VPWR.n1709 161.3
R10071 VPWR.n1070 VPWR.n1069 161.3
R10072 VPWR.n1719 VPWR.n1718 161.3
R10073 VPWR.n1722 VPWR.n1721 161.3
R10074 VPWR.n1717 VPWR.n1716 161.3
R10075 VPWR.n1734 VPWR.n1733 161.3
R10076 VPWR.n1117 VPWR.n1116 161.3
R10077 VPWR.n1731 VPWR.n1730 161.3
R10078 VPWR.n1065 VPWR.n1064 161.3
R10079 VPWR.n126 VPWR.n125 161.3
R10080 VPWR.n117 VPWR.n116 161.3
R10081 VPWR.n120 VPWR.n119 161.3
R10082 VPWR.n115 VPWR.n114 161.3
R10083 VPWR.n138 VPWR.n137 161.3
R10084 VPWR.n128 VPWR.n127 161.3
R10085 VPWR.n109 VPWR.n108 161.3
R10086 VPWR.n105 VPWR.n104 161.3
R10087 VPWR.n288 VPWR.n287 161.3
R10088 VPWR.n285 VPWR.n284 161.3
R10089 VPWR.n101 VPWR.n100 161.3
R10090 VPWR.n272 VPWR.n271 161.3
R10091 VPWR.n275 VPWR.n274 161.3
R10092 VPWR.n270 VPWR.n269 161.3
R10093 VPWR.n260 VPWR.n259 161.3
R10094 VPWR.n263 VPWR.n262 161.3
R10095 VPWR.n258 VPWR.n257 161.3
R10096 VPWR.n248 VPWR.n247 161.3
R10097 VPWR.n251 VPWR.n250 161.3
R10098 VPWR.n246 VPWR.n245 161.3
R10099 VPWR.n236 VPWR.n235 161.3
R10100 VPWR.n239 VPWR.n238 161.3
R10101 VPWR.n234 VPWR.n233 161.3
R10102 VPWR.n224 VPWR.n223 161.3
R10103 VPWR.n227 VPWR.n226 161.3
R10104 VPWR.n222 VPWR.n221 161.3
R10105 VPWR.n212 VPWR.n211 161.3
R10106 VPWR.n215 VPWR.n214 161.3
R10107 VPWR.n210 VPWR.n209 161.3
R10108 VPWR.n200 VPWR.n199 161.3
R10109 VPWR.n203 VPWR.n202 161.3
R10110 VPWR.n198 VPWR.n197 161.3
R10111 VPWR.n188 VPWR.n187 161.3
R10112 VPWR.n191 VPWR.n190 161.3
R10113 VPWR.n186 VPWR.n185 161.3
R10114 VPWR.n176 VPWR.n175 161.3
R10115 VPWR.n179 VPWR.n178 161.3
R10116 VPWR.n174 VPWR.n173 161.3
R10117 VPWR.n164 VPWR.n163 161.3
R10118 VPWR.n167 VPWR.n166 161.3
R10119 VPWR.n162 VPWR.n161 161.3
R10120 VPWR.n152 VPWR.n151 161.3
R10121 VPWR.n155 VPWR.n154 161.3
R10122 VPWR.n150 VPWR.n149 161.3
R10123 VPWR.n140 VPWR.n139 161.3
R10124 VPWR.n143 VPWR.n142 161.3
R10125 VPWR.n131 VPWR.n130 161.3
R10126 VPWR.n1601 VPWR.t611 161.202
R10127 VPWR.n1106 VPWR.t736 161.202
R10128 VPWR.n1617 VPWR.t777 161.202
R10129 VPWR.n1628 VPWR.t885 161.202
R10130 VPWR.n1096 VPWR.t652 161.202
R10131 VPWR.n1644 VPWR.t667 161.202
R10132 VPWR.n1655 VPWR.t890 161.202
R10133 VPWR.n1086 VPWR.t933 161.202
R10134 VPWR.n1671 VPWR.t650 161.202
R10135 VPWR.n1682 VPWR.t803 161.202
R10136 VPWR.n1076 VPWR.t825 161.202
R10137 VPWR.n1698 VPWR.t675 161.202
R10138 VPWR.n1709 VPWR.t701 161.202
R10139 VPWR.n1721 VPWR.t726 161.202
R10140 VPWR.n1116 VPWR.t866 161.202
R10141 VPWR.n1730 VPWR.t571 161.202
R10142 VPWR.n119 VPWR.t693 161.202
R10143 VPWR.n108 VPWR.t592 161.202
R10144 VPWR.n284 VPWR.t728 161.202
R10145 VPWR.n274 VPWR.t858 161.202
R10146 VPWR.n262 VPWR.t898 161.202
R10147 VPWR.n250 VPWR.t622 161.202
R10148 VPWR.n238 VPWR.t766 161.202
R10149 VPWR.n226 VPWR.t790 161.202
R10150 VPWR.n214 VPWR.t627 161.202
R10151 VPWR.n202 VPWR.t662 161.202
R10152 VPWR.n190 VPWR.t764 161.202
R10153 VPWR.n178 VPWR.t925 161.202
R10154 VPWR.n166 VPWR.t944 161.202
R10155 VPWR.n154 VPWR.t798 161.202
R10156 VPWR.n1768 VPWR.t850 161.202
R10157 VPWR.n1039 VPWR.t606 161.202
R10158 VPWR.n1543 VPWR.t587 161.202
R10159 VPWR.n1548 VPWR.t836 161.202
R10160 VPWR.n1553 VPWR.t718 161.202
R10161 VPWR.n1558 VPWR.t688 161.202
R10162 VPWR.n1563 VPWR.t840 161.202
R10163 VPWR.n1568 VPWR.t838 161.202
R10164 VPWR.n1573 VPWR.t683 161.202
R10165 VPWR.n1578 VPWR.t573 161.202
R10166 VPWR.n1133 VPWR.t917 161.202
R10167 VPWR.n1458 VPWR.t788 161.202
R10168 VPWR.n1453 VPWR.t657 161.202
R10169 VPWR.n1773 VPWR.t868 161.202
R10170 VPWR.n1781 VPWR.t906 161.202
R10171 VPWR.n1777 VPWR.t738 161.202
R10172 VPWR.n142 VPWR.t817 161.202
R10173 VPWR.n130 VPWR.t842 161.202
R10174 VPWR.n1119 VPWR.t594 161.106
R10175 VPWR.n1110 VPWR.t730 161.106
R10176 VPWR.n1611 VPWR.t743 161.106
R10177 VPWR.n1622 VPWR.t903 161.106
R10178 VPWR.n1100 VPWR.t624 161.106
R10179 VPWR.n1638 VPWR.t771 161.106
R10180 VPWR.n1649 VPWR.t882 161.106
R10181 VPWR.n1090 VPWR.t919 161.106
R10182 VPWR.n1665 VPWR.t664 161.106
R10183 VPWR.n1676 VPWR.t768 161.106
R10184 VPWR.n1080 VPWR.t927 161.106
R10185 VPWR.n1692 VPWR.t946 161.106
R10186 VPWR.n1703 VPWR.t690 161.106
R10187 VPWR.n1069 VPWR.t819 161.106
R10188 VPWR.n1716 VPWR.t847 161.106
R10189 VPWR.n1064 VPWR.t698 161.106
R10190 VPWR.n125 VPWR.t578 161.106
R10191 VPWR.n114 VPWR.t814 161.106
R10192 VPWR.n137 VPWR.t938 161.106
R10193 VPWR.n104 VPWR.t723 161.106
R10194 VPWR.n100 VPWR.t852 161.106
R10195 VPWR.n269 VPWR.t870 161.106
R10196 VPWR.n257 VPWR.t632 161.106
R10197 VPWR.n245 VPWR.t740 161.106
R10198 VPWR.n233 VPWR.t895 161.106
R10199 VPWR.n221 VPWR.t619 161.106
R10200 VPWR.n209 VPWR.t654 161.106
R10201 VPWR.n197 VPWR.t782 161.106
R10202 VPWR.n185 VPWR.t892 161.106
R10203 VPWR.n173 VPWR.t659 161.106
R10204 VPWR.n161 VPWR.t677 161.106
R10205 VPWR.n149 VPWR.t805 161.106
R10206 VPWR.n53 VPWR.t922 161.106
R10207 VPWR.n51 VPWR.t879 161.106
R10208 VPWR.n49 VPWR.t600 161.106
R10209 VPWR.n47 VPWR.t712 161.106
R10210 VPWR.n45 VPWR.t930 161.106
R10211 VPWR.n43 VPWR.t779 161.106
R10212 VPWR.n41 VPWR.t887 161.106
R10213 VPWR.n39 VPWR.t613 161.106
R10214 VPWR.n37 VPWR.t720 161.106
R10215 VPWR.n35 VPWR.t680 161.106
R10216 VPWR.n33 VPWR.t785 161.106
R10217 VPWR.n31 VPWR.t608 161.106
R10218 VPWR.n29 VPWR.t792 161.106
R10219 VPWR.n27 VPWR.t900 161.106
R10220 VPWR.n25 VPWR.t752 161.106
R10221 VPWR.n23 VPWR.t863 161.106
R10222 VPWR.n1598 VPWR.t644 159.978
R10223 VPWR.n1125 VPWR.t746 159.978
R10224 VPWR.n1614 VPWR.t911 159.978
R10225 VPWR.n1625 VPWR.t629 159.978
R10226 VPWR.n1176 VPWR.t641 159.978
R10227 VPWR.n1641 VPWR.t800 159.978
R10228 VPWR.n1652 VPWR.t908 159.978
R10229 VPWR.n1208 VPWR.t669 159.978
R10230 VPWR.n1668 VPWR.t695 159.978
R10231 VPWR.n1679 VPWR.t822 159.978
R10232 VPWR.n1194 VPWR.t568 159.978
R10233 VPWR.n1695 VPWR.t589 159.978
R10234 VPWR.n1706 VPWR.t827 159.978
R10235 VPWR.n1718 VPWR.t855 159.978
R10236 VPWR.n1733 VPWR.t575 159.978
R10237 VPWR.n1114 VPWR.t876 159.978
R10238 VPWR.n116 VPWR.t709 159.978
R10239 VPWR.n127 VPWR.t584 159.978
R10240 VPWR.n106 VPWR.t616 159.978
R10241 VPWR.n287 VPWR.t761 159.978
R10242 VPWR.n271 VPWR.t873 159.978
R10243 VPWR.n259 VPWR.t638 159.978
R10244 VPWR.n247 VPWR.t749 159.978
R10245 VPWR.n235 VPWR.t758 159.978
R10246 VPWR.n223 VPWR.t914 159.978
R10247 VPWR.n211 VPWR.t635 159.978
R10248 VPWR.n199 VPWR.t795 159.978
R10249 VPWR.n187 VPWR.t811 159.978
R10250 VPWR.n175 VPWR.t941 159.978
R10251 VPWR.n163 VPWR.t685 159.978
R10252 VPWR.n151 VPWR.t715 159.978
R10253 VPWR.n1228 VPWR.t672 159.978
R10254 VPWR.n1150 VPWR.t603 159.978
R10255 VPWR.n1224 VPWR.t808 159.978
R10256 VPWR.n1482 VPWR.t706 159.978
R10257 VPWR.n1170 VPWR.t830 159.978
R10258 VPWR.n1166 VPWR.t581 159.978
R10259 VPWR.n1160 VPWR.t703 159.978
R10260 VPWR.n1476 VPWR.t935 159.978
R10261 VPWR.n1156 VPWR.t844 159.978
R10262 VPWR.n1146 VPWR.t860 159.978
R10263 VPWR.n1469 VPWR.t833 159.978
R10264 VPWR.n1046 VPWR.t733 159.978
R10265 VPWR.n1745 VPWR.t597 159.978
R10266 VPWR.n1033 VPWR.t647 159.978
R10267 VPWR.n1029 VPWR.t755 159.978
R10268 VPWR.n1050 VPWR.t774 159.978
R10269 VPWR.n139 VPWR.t565 159.978
R10270 VPWR.n1229 VPWR.n1228 152
R10271 VPWR.n1151 VPWR.n1150 152
R10272 VPWR.n1225 VPWR.n1224 152
R10273 VPWR.n1483 VPWR.n1482 152
R10274 VPWR.n1171 VPWR.n1170 152
R10275 VPWR.n1167 VPWR.n1166 152
R10276 VPWR.n1161 VPWR.n1160 152
R10277 VPWR.n1477 VPWR.n1476 152
R10278 VPWR.n1157 VPWR.n1156 152
R10279 VPWR.n1147 VPWR.n1146 152
R10280 VPWR.n1470 VPWR.n1469 152
R10281 VPWR.n1047 VPWR.n1046 152
R10282 VPWR.n1746 VPWR.n1745 152
R10283 VPWR.n1034 VPWR.n1033 152
R10284 VPWR.n1030 VPWR.n1029 152
R10285 VPWR.n1051 VPWR.n1050 152
R10286 VPWR.n2845 VPWR.n2844 150.213
R10287 VPWR.n1601 VPWR.t2063 145.137
R10288 VPWR.n1106 VPWR.t2014 145.137
R10289 VPWR.n1617 VPWR.t2000 145.137
R10290 VPWR.n1628 VPWR.t1962 145.137
R10291 VPWR.n1096 VPWR.t2049 145.137
R10292 VPWR.n1644 VPWR.t2042 145.137
R10293 VPWR.n1655 VPWR.t1959 145.137
R10294 VPWR.n1086 VPWR.t1945 145.137
R10295 VPWR.n1671 VPWR.t2050 145.137
R10296 VPWR.n1682 VPWR.t1993 145.137
R10297 VPWR.n1076 VPWR.t1988 145.137
R10298 VPWR.n1698 VPWR.t2040 145.137
R10299 VPWR.n1709 VPWR.t2033 145.137
R10300 VPWR.n1721 VPWR.t2019 145.137
R10301 VPWR.n1116 VPWR.t1969 145.137
R10302 VPWR.n1730 VPWR.t1937 145.137
R10303 VPWR.n119 VPWR.t2048 145.137
R10304 VPWR.n108 VPWR.t1934 145.137
R10305 VPWR.n284 VPWR.t2030 145.137
R10306 VPWR.n274 VPWR.t1983 145.137
R10307 VPWR.n262 VPWR.t1971 145.137
R10308 VPWR.n250 VPWR.t1930 145.137
R10309 VPWR.n238 VPWR.t2016 145.137
R10310 VPWR.n226 VPWR.t2008 145.137
R10311 VPWR.n214 VPWR.t1928 145.137
R10312 VPWR.n202 VPWR.t2057 145.137
R10313 VPWR.n190 VPWR.t2017 145.137
R10314 VPWR.n178 VPWR.t1961 145.137
R10315 VPWR.n166 VPWR.t1952 145.137
R10316 VPWR.n154 VPWR.t2007 145.137
R10317 VPWR.n1768 VPWR.t1976 145.137
R10318 VPWR.n1039 VPWR.t2065 145.137
R10319 VPWR.n1543 VPWR.t1929 145.137
R10320 VPWR.n1548 VPWR.t1986 145.137
R10321 VPWR.n1553 VPWR.t2025 145.137
R10322 VPWR.n1558 VPWR.t2037 145.137
R10323 VPWR.n1563 VPWR.t1979 145.137
R10324 VPWR.n1568 VPWR.t1985 145.137
R10325 VPWR.n1573 VPWR.t2039 145.137
R10326 VPWR.n1578 VPWR.t1936 145.137
R10327 VPWR.n1133 VPWR.t1950 145.137
R10328 VPWR.n1458 VPWR.t1996 145.137
R10329 VPWR.n1453 VPWR.t2045 145.137
R10330 VPWR.n1773 VPWR.t1968 145.137
R10331 VPWR.n1781 VPWR.t1953 145.137
R10332 VPWR.n1777 VPWR.t2013 145.137
R10333 VPWR.n142 VPWR.t1999 145.137
R10334 VPWR.n130 VPWR.t1990 145.137
R10335 VPWR.n1119 VPWR.t2067 145.038
R10336 VPWR.n1110 VPWR.t2018 145.038
R10337 VPWR.n1611 VPWR.t2010 145.038
R10338 VPWR.n1622 VPWR.t1955 145.038
R10339 VPWR.n1100 VPWR.t2059 145.038
R10340 VPWR.n1638 VPWR.t2002 145.038
R10341 VPWR.n1649 VPWR.t1964 145.038
R10342 VPWR.n1090 VPWR.t1949 145.038
R10343 VPWR.n1665 VPWR.t2043 145.038
R10344 VPWR.n1676 VPWR.t2003 145.038
R10345 VPWR.n1080 VPWR.t1947 145.038
R10346 VPWR.n1692 VPWR.t1939 145.038
R10347 VPWR.n1703 VPWR.t2036 145.038
R10348 VPWR.n1069 VPWR.t1989 145.038
R10349 VPWR.n1716 VPWR.t1977 145.038
R10350 VPWR.n1064 VPWR.t2034 145.038
R10351 VPWR.n125 VPWR.t1940 145.038
R10352 VPWR.n114 VPWR.t2001 145.038
R10353 VPWR.n137 VPWR.t1954 145.038
R10354 VPWR.n104 VPWR.t2032 145.038
R10355 VPWR.n100 VPWR.t1987 145.038
R10356 VPWR.n269 VPWR.t1980 145.038
R10357 VPWR.n257 VPWR.t2068 145.038
R10358 VPWR.n245 VPWR.t2027 145.038
R10359 VPWR.n233 VPWR.t1972 145.038
R10360 VPWR.n221 VPWR.t1931 145.038
R10361 VPWR.n209 VPWR.t2060 145.038
R10362 VPWR.n197 VPWR.t2009 145.038
R10363 VPWR.n185 VPWR.t1973 145.038
R10364 VPWR.n173 VPWR.t2058 145.038
R10365 VPWR.n161 VPWR.t2052 145.038
R10366 VPWR.n149 VPWR.t2004 145.038
R10367 VPWR.n53 VPWR.t2053 145.038
R10368 VPWR.n51 VPWR.t1963 145.038
R10369 VPWR.n49 VPWR.t2066 145.038
R10370 VPWR.n47 VPWR.t2026 145.038
R10371 VPWR.n45 VPWR.t1946 145.038
R10372 VPWR.n43 VPWR.t2051 145.038
R10373 VPWR.n41 VPWR.t2069 145.038
R10374 VPWR.n39 VPWR.t2028 145.038
R10375 VPWR.n37 VPWR.t2022 145.038
R10376 VPWR.n35 VPWR.t1943 145.038
R10377 VPWR.n33 VPWR.t1997 145.038
R10378 VPWR.n31 VPWR.t2064 145.038
R10379 VPWR.n29 VPWR.t1995 145.038
R10380 VPWR.n27 VPWR.t1956 145.038
R10381 VPWR.n25 VPWR.t2021 145.038
R10382 VPWR.n23 VPWR.t1970 145.038
R10383 VPWR.n1598 VPWR.t1966 143.911
R10384 VPWR.n1125 VPWR.t2062 143.911
R10385 VPWR.n1614 VPWR.t2047 143.911
R10386 VPWR.n1625 VPWR.t1965 143.911
R10387 VPWR.n1176 VPWR.t1958 143.911
R10388 VPWR.n1641 VPWR.t1944 143.911
R10389 VPWR.n1652 VPWR.t2005 143.911
R10390 VPWR.n1208 VPWR.t1992 143.911
R10391 VPWR.n1668 VPWR.t1941 143.911
R10392 VPWR.n1679 VPWR.t2038 143.911
R10393 VPWR.n1194 VPWR.t2031 143.911
R10394 VPWR.n1695 VPWR.t1978 143.911
R10395 VPWR.n1706 VPWR.t1935 143.911
R10396 VPWR.n1718 VPWR.t2024 143.911
R10397 VPWR.n1733 VPWR.t1984 143.911
R10398 VPWR.n1114 VPWR.t2012 143.911
R10399 VPWR.n116 VPWR.t1951 143.911
R10400 VPWR.n127 VPWR.t1991 143.911
R10401 VPWR.n106 VPWR.t1981 143.911
R10402 VPWR.n287 VPWR.t1933 143.911
R10403 VPWR.n271 VPWR.t2029 143.911
R10404 VPWR.n259 VPWR.t2015 143.911
R10405 VPWR.n247 VPWR.t1932 143.911
R10406 VPWR.n235 VPWR.t1926 143.911
R10407 VPWR.n223 VPWR.t2056 143.911
R10408 VPWR.n211 VPWR.t1974 143.911
R10409 VPWR.n199 VPWR.t1960 143.911
R10410 VPWR.n187 VPWR.t2054 143.911
R10411 VPWR.n175 VPWR.t2006 143.911
R10412 VPWR.n163 VPWR.t1998 143.911
R10413 VPWR.n151 VPWR.t1942 143.911
R10414 VPWR.n1228 VPWR.t1948 143.911
R10415 VPWR.n1150 VPWR.t1975 143.911
R10416 VPWR.n1224 VPWR.t2041 143.911
R10417 VPWR.n1482 VPWR.t1982 143.911
R10418 VPWR.n1170 VPWR.t2035 143.911
R10419 VPWR.n1166 VPWR.t2023 143.911
R10420 VPWR.n1160 VPWR.t1938 143.911
R10421 VPWR.n1476 VPWR.t1994 143.911
R10422 VPWR.n1156 VPWR.t1927 143.911
R10423 VPWR.n1146 VPWR.t2020 143.911
R10424 VPWR.n1469 VPWR.t2044 143.911
R10425 VPWR.n1046 VPWR.t1967 143.911
R10426 VPWR.n1745 VPWR.t2011 143.911
R10427 VPWR.n1033 VPWR.t1957 143.911
R10428 VPWR.n1029 VPWR.t2061 143.911
R10429 VPWR.n1050 VPWR.t2055 143.911
R10430 VPWR.n139 VPWR.t2046 143.911
R10431 VPWR.t264 VPWR.t1764 140.989
R10432 VPWR.t1787 VPWR.t1774 140.989
R10433 VPWR.t1814 VPWR.t1787 140.989
R10434 VPWR.t1790 VPWR.t1814 140.989
R10435 VPWR.t1092 VPWR.t1790 140.989
R10436 VPWR.t1355 VPWR.t1092 140.989
R10437 VPWR.t91 VPWR.t1355 140.989
R10438 VPWR.t453 VPWR.t91 140.989
R10439 VPWR.t1210 VPWR.t1388 140.989
R10440 VPWR.t1826 VPWR.t1793 140.989
R10441 VPWR.t1780 VPWR.t1826 140.989
R10442 VPWR.t1827 VPWR.t1780 140.989
R10443 VPWR.t1228 VPWR.t1827 140.989
R10444 VPWR.t1240 VPWR.t1228 140.989
R10445 VPWR.t1232 VPWR.t1240 140.989
R10446 VPWR.t1236 VPWR.t1232 140.989
R10447 VPWR.t1771 VPWR.t1812 140.989
R10448 VPWR.t1801 VPWR.t1771 140.989
R10449 VPWR.t1775 VPWR.t1801 140.989
R10450 VPWR.t547 VPWR.t1775 140.989
R10451 VPWR.t541 VPWR.t547 140.989
R10452 VPWR.t549 VPWR.t541 140.989
R10453 VPWR.t551 VPWR.t549 140.989
R10454 VPWR.t1369 VPWR.t1802 140.989
R10455 VPWR.t1772 VPWR.t1815 140.989
R10456 VPWR.t1822 VPWR.t1772 140.989
R10457 VPWR.t1799 VPWR.t1822 140.989
R10458 VPWR.t2 VPWR.t1799 140.989
R10459 VPWR.t1506 VPWR.t2 140.989
R10460 VPWR.t1244 VPWR.t1506 140.989
R10461 VPWR.t1226 VPWR.t1244 140.989
R10462 VPWR.t1794 VPWR.t1781 140.989
R10463 VPWR.t1768 VPWR.t1794 140.989
R10464 VPWR.t1820 VPWR.t1768 140.989
R10465 VPWR.t1238 VPWR.t1820 140.989
R10466 VPWR.t1230 VPWR.t1238 140.989
R10467 VPWR.t1242 VPWR.t1230 140.989
R10468 VPWR.t1234 VPWR.t1242 140.989
R10469 VPWR.t1791 VPWR.t1783 140.989
R10470 VPWR.t1797 VPWR.t1791 140.989
R10471 VPWR.t1785 VPWR.t1797 140.989
R10472 VPWR.t543 VPWR.t1785 140.989
R10473 VPWR.t537 VPWR.t543 140.989
R10474 VPWR.t545 VPWR.t537 140.989
R10475 VPWR.t539 VPWR.t545 140.989
R10476 VPWR VPWR.n1442 133.312
R10477 VPWR.n2841 VPWR.n2840 129.13
R10478 VPWR.n2858 VPWR.n2819 129.13
R10479 VPWR.n2780 VPWR 127.562
R10480 VPWR.n2760 VPWR 127.562
R10481 VPWR.n2741 VPWR 127.562
R10482 VPWR VPWR.t1833 125.883
R10483 VPWR.n2705 VPWR 125.883
R10484 VPWR.t1212 VPWR.t1390 120.849
R10485 VPWR.t950 VPWR.t976 117.492
R10486 VPWR.t455 VPWR.t1891 117.492
R10487 VPWR.t1907 VPWR 115.814
R10488 VPWR VPWR.t453 114.135
R10489 VPWR VPWR.t1236 114.135
R10490 VPWR VPWR.t551 114.135
R10491 VPWR.n2859 VPWR.n2817 111.059
R10492 VPWR.t1407 VPWR 107.421
R10493 VPWR.n1330 VPWR.n1329 106.561
R10494 VPWR.n2781 VPWR.n2780 106.561
R10495 VPWR.n2761 VPWR.n2760 106.561
R10496 VPWR.n2742 VPWR.n2741 106.561
R10497 VPWR.n2706 VPWR.n2705 106.561
R10498 VPWR.n2668 VPWR.n2667 106.561
R10499 VPWR.n2631 VPWR.n2630 106.561
R10500 VPWR VPWR.t1216 106.543
R10501 VPWR VPWR.n1234 104.8
R10502 VPWR VPWR.n1257 104.8
R10503 VPWR VPWR.n1281 104.8
R10504 VPWR VPWR.n1366 104.8
R10505 VPWR VPWR.n1405 104.8
R10506 VPWR.n1443 VPWR 100.883
R10507 VPWR VPWR.t1727 100.624
R10508 VPWR.t1094 VPWR.t266 97.9386
R10509 VPWR.n2859 VPWR.n2858 93.3652
R10510 VPWR.n1231 VPWR.n1230 91.8492
R10511 VPWR.n1153 VPWR.n1152 91.8492
R10512 VPWR.n1227 VPWR.n1226 91.8492
R10513 VPWR.n1485 VPWR.n1484 91.8492
R10514 VPWR.n1173 VPWR.n1172 91.8492
R10515 VPWR.n1169 VPWR.n1168 91.8492
R10516 VPWR.n1163 VPWR.n1162 91.8492
R10517 VPWR.n1479 VPWR.n1478 91.8492
R10518 VPWR.n1159 VPWR.n1158 91.8492
R10519 VPWR.n1149 VPWR.n1148 91.8492
R10520 VPWR.n1472 VPWR.n1471 91.8492
R10521 VPWR.n1049 VPWR.n1048 91.8492
R10522 VPWR.n1748 VPWR.n1747 91.8492
R10523 VPWR.n1036 VPWR.n1035 91.8492
R10524 VPWR.n1032 VPWR.n1031 91.8492
R10525 VPWR.n1053 VPWR.n1052 91.8492
R10526 VPWR.n2847 VPWR.n2820 91.4829
R10527 VPWR.t1094 VPWR.n2842 90.0872
R10528 VPWR.t1818 VPWR 88.7855
R10529 VPWR.n1235 VPWR 79.407
R10530 VPWR.n1258 VPWR 79.407
R10531 VPWR.n1282 VPWR 79.407
R10532 VPWR.n1367 VPWR 79.407
R10533 VPWR.n1406 VPWR 79.407
R10534 VPWR.t457 VPWR.t1741 78.8874
R10535 VPWR.n2840 VPWR.n2818 74.9181
R10536 VPWR.n2858 VPWR.n2818 74.9181
R10537 VPWR.n2858 VPWR.n2857 74.9181
R10538 VPWR.n2857 VPWR.n2820 74.9181
R10539 VPWR.t306 VPWR.t1729 70.4952
R10540 VPWR.t1729 VPWR.t418 70.4952
R10541 VPWR.t418 VPWR.t260 70.4952
R10542 VPWR.t260 VPWR.t1115 70.4952
R10543 VPWR.t1115 VPWR.t142 70.4952
R10544 VPWR.t142 VPWR.t1757 70.4952
R10545 VPWR.t1757 VPWR.t264 70.4952
R10546 VPWR.t1806 VPWR.t1369 70.4952
R10547 VPWR.t1363 VPWR.t1806 70.4952
R10548 VPWR.t1778 VPWR.t1363 70.4952
R10549 VPWR.t1371 VPWR.t1778 70.4952
R10550 VPWR.t1810 VPWR.t1371 70.4952
R10551 VPWR.t1365 VPWR.t1810 70.4952
R10552 VPWR.t1833 VPWR.t1365 70.4952
R10553 VPWR VPWR.t306 68.8168
R10554 VPWR.t1218 VPWR.t1214 68.8168
R10555 VPWR.t1741 VPWR.t1907 62.103
R10556 VPWR VPWR.t1210 60.4245
R10557 VPWR.n2849 VPWR.n2842 59.762
R10558 VPWR.n2845 VPWR.n2819 53.8358
R10559 VPWR.t1214 VPWR.t14 52.0323
R10560 VPWR.t524 VPWR 50.3539
R10561 VPWR VPWR.t1218 50.3539
R10562 VPWR VPWR.t1212 50.3539
R10563 VPWR.t1815 VPWR 50.3539
R10564 VPWR.t1781 VPWR 50.3539
R10565 VPWR.t1783 VPWR 50.3539
R10566 VPWR.n2854 VPWR.n2818 46.2505
R10567 VPWR.n2855 VPWR.n2854 46.2505
R10568 VPWR.n2835 VPWR.n2834 46.2505
R10569 VPWR.n2836 VPWR.n2835 46.2505
R10570 VPWR.n2838 VPWR.n2837 46.2505
R10571 VPWR.n2837 VPWR.n2836 46.2505
R10572 VPWR.n2844 VPWR.n2824 46.2505
R10573 VPWR.n2857 VPWR.n2856 46.2505
R10574 VPWR.n2856 VPWR.n2855 46.2505
R10575 VPWR.n2849 VPWR.n2848 46.2505
R10576 VPWR.n2846 VPWR.n2845 45.9299
R10577 VPWR.n2832 VPWR.n2830 44.8005
R10578 VPWR.n2830 VPWR.n2826 44.8005
R10579 VPWR.n2847 VPWR.n2843 37.0005
R10580 VPWR.n2843 VPWR.t266 37.0005
R10581 VPWR.n1230 VPWR.n1229 34.7473
R10582 VPWR.n1152 VPWR.n1151 34.7473
R10583 VPWR.n1226 VPWR.n1225 34.7473
R10584 VPWR.n1484 VPWR.n1483 34.7473
R10585 VPWR.n1172 VPWR.n1171 34.7473
R10586 VPWR.n1168 VPWR.n1167 34.7473
R10587 VPWR.n1162 VPWR.n1161 34.7473
R10588 VPWR.n1478 VPWR.n1477 34.7473
R10589 VPWR.n1158 VPWR.n1157 34.7473
R10590 VPWR.n1148 VPWR.n1147 34.7473
R10591 VPWR.n1471 VPWR.n1470 34.7473
R10592 VPWR.n1048 VPWR.n1047 34.7473
R10593 VPWR.n1747 VPWR.n1746 34.7473
R10594 VPWR.n1035 VPWR.n1034 34.7473
R10595 VPWR.n1031 VPWR.n1030 34.7473
R10596 VPWR.n1052 VPWR.n1051 34.7473
R10597 VPWR.n1299 VPWR.n1298 34.6358
R10598 VPWR.n1357 VPWR.n1341 34.6358
R10599 VPWR.n1362 VPWR.n1361 34.6358
R10600 VPWR.n1396 VPWR.n1380 34.6358
R10601 VPWR.n1401 VPWR.n1400 34.6358
R10602 VPWR.n1411 VPWR.n1377 34.6358
R10603 VPWR.n1433 VPWR.n1417 34.6358
R10604 VPWR.n1438 VPWR.n1437 34.6358
R10605 VPWR.n2755 VPWR.n2754 34.6358
R10606 VPWR.n2721 VPWR.n2713 34.6358
R10607 VPWR.n2728 VPWR.n2727 34.6358
R10608 VPWR.n2685 VPWR.n2676 34.6358
R10609 VPWR.n2688 VPWR.n2687 34.6358
R10610 VPWR.n2692 VPWR.n2691 34.6358
R10611 VPWR.n2648 VPWR.n2639 34.6358
R10612 VPWR.n2651 VPWR.n2650 34.6358
R10613 VPWR.n2655 VPWR.n2654 34.6358
R10614 VPWR.n2662 VPWR.n2661 34.6358
R10615 VPWR.n2615 VPWR.n2611 34.6358
R10616 VPWR.n2619 VPWR.n2603 34.6358
R10617 VPWR.n2622 VPWR.n2621 34.6358
R10618 VPWR.n1316 VPWR.n1315 32.0005
R10619 VPWR.n1353 VPWR.n1352 32.0005
R10620 VPWR.n1392 VPWR.n1391 32.0005
R10621 VPWR.n1429 VPWR.n1428 32.0005
R10622 VPWR.n2717 VPWR.n2716 30.8711
R10623 VPWR.n2681 VPWR.n2680 30.8711
R10624 VPWR.n2644 VPWR.n2643 30.8711
R10625 VPWR.n2610 VPWR.n2609 30.8711
R10626 VPWR.n2834 VPWR.n2832 30.1181
R10627 VPWR.n2838 VPWR.n2826 30.1181
R10628 VPWR.n2848 VPWR.n2846 28.9887
R10629 VPWR.n1325 VPWR.n1324 28.2358
R10630 VPWR.n5 VPWR.t263 26.5955
R10631 VPWR.n5 VPWR.t141 26.5955
R10632 VPWR.n4 VPWR.t1728 26.5955
R10633 VPWR.n4 VPWR.t259 26.5955
R10634 VPWR.n1240 VPWR.t1597 26.5955
R10635 VPWR.n1240 VPWR.t1596 26.5955
R10636 VPWR.n1239 VPWR.t1195 26.5955
R10637 VPWR.n1239 VPWR.t1013 26.5955
R10638 VPWR.n1245 VPWR.t1593 26.5955
R10639 VPWR.n1245 VPWR.t1598 26.5955
R10640 VPWR.n1238 VPWR.t1434 26.5955
R10641 VPWR.n1238 VPWR.t1194 26.5955
R10642 VPWR.n1263 VPWR.t1300 26.5955
R10643 VPWR.n1263 VPWR.t1301 26.5955
R10644 VPWR.n1262 VPWR.t338 26.5955
R10645 VPWR.n1262 VPWR.t336 26.5955
R10646 VPWR.n1268 VPWR.t155 26.5955
R10647 VPWR.n1268 VPWR.t157 26.5955
R10648 VPWR.n1261 VPWR.t341 26.5955
R10649 VPWR.n1261 VPWR.t339 26.5955
R10650 VPWR.n1287 VPWR.t1030 26.5955
R10651 VPWR.n1287 VPWR.t1037 26.5955
R10652 VPWR.n1286 VPWR.t1351 26.5955
R10653 VPWR.n1286 VPWR.t1350 26.5955
R10654 VPWR.n1292 VPWR.t1034 26.5955
R10655 VPWR.n1292 VPWR.t1031 26.5955
R10656 VPWR.n1285 VPWR.t1354 26.5955
R10657 VPWR.n1285 VPWR.t1352 26.5955
R10658 VPWR.n1314 VPWR.t1767 26.5955
R10659 VPWR.n1314 VPWR.t1294 26.5955
R10660 VPWR.n1307 VPWR.t265 26.5955
R10661 VPWR.n1307 VPWR.t1765 26.5955
R10662 VPWR.n1321 VPWR.t261 26.5955
R10663 VPWR.n1321 VPWR.t143 26.5955
R10664 VPWR.n1323 VPWR.t419 26.5955
R10665 VPWR.n1323 VPWR.t1116 26.5955
R10666 VPWR.n1351 VPWR.t386 26.5955
R10667 VPWR.n1351 VPWR.t22 26.5955
R10668 VPWR.n1350 VPWR.t1297 26.5955
R10669 VPWR.n1350 VPWR.t1760 26.5955
R10670 VPWR.n1344 VPWR.t1600 26.5955
R10671 VPWR.n1344 VPWR.t365 26.5955
R10672 VPWR.n1343 VPWR.t1435 26.5955
R10673 VPWR.n1343 VPWR.t1312 26.5955
R10674 VPWR.n1359 VPWR.t1595 26.5955
R10675 VPWR.n1359 VPWR.t1594 26.5955
R10676 VPWR.n1358 VPWR.t1014 26.5955
R10677 VPWR.n1358 VPWR.t1193 26.5955
R10678 VPWR.n1390 VPWR.t1311 26.5955
R10679 VPWR.n1390 VPWR.t1299 26.5955
R10680 VPWR.n1389 VPWR.t388 26.5955
R10681 VPWR.n1389 VPWR.t24 26.5955
R10682 VPWR.n1383 VPWR.t1889 26.5955
R10683 VPWR.n1383 VPWR.t1296 26.5955
R10684 VPWR.n1382 VPWR.t342 26.5955
R10685 VPWR.n1382 VPWR.t369 26.5955
R10686 VPWR.n1398 VPWR.t1888 26.5955
R10687 VPWR.n1398 VPWR.t1890 26.5955
R10688 VPWR.n1397 VPWR.t343 26.5955
R10689 VPWR.n1397 VPWR.t340 26.5955
R10690 VPWR.n1427 VPWR.t305 26.5955
R10691 VPWR.n1427 VPWR.t420 26.5955
R10692 VPWR.n1426 VPWR.t1298 26.5955
R10693 VPWR.n1426 VPWR.t1761 26.5955
R10694 VPWR.n1420 VPWR.t1033 26.5955
R10695 VPWR.n1420 VPWR.t301 26.5955
R10696 VPWR.n1419 VPWR.t1348 26.5955
R10697 VPWR.n1419 VPWR.t1313 26.5955
R10698 VPWR.n1435 VPWR.t1036 26.5955
R10699 VPWR.n1435 VPWR.t1035 26.5955
R10700 VPWR.n1434 VPWR.t1349 26.5955
R10701 VPWR.n1434 VPWR.t1347 26.5955
R10702 VPWR.n2802 VPWR.t1374 26.5955
R10703 VPWR.n2802 VPWR.t1376 26.5955
R10704 VPWR.n2804 VPWR.t1368 26.5955
R10705 VPWR.n2804 VPWR.t1362 26.5955
R10706 VPWR.n2782 VPWR.t1670 26.5955
R10707 VPWR.n2782 VPWR.t1667 26.5955
R10708 VPWR.n2783 VPWR.t1093 26.5955
R10709 VPWR.n2783 VPWR.t1356 26.5955
R10710 VPWR.n2786 VPWR.t1663 26.5955
R10711 VPWR.n2786 VPWR.t1664 26.5955
R10712 VPWR.n2787 VPWR.t92 26.5955
R10713 VPWR.n2787 VPWR.t454 26.5955
R10714 VPWR.n2762 VPWR.t1284 26.5955
R10715 VPWR.n2762 VPWR.t1488 26.5955
R10716 VPWR.n2763 VPWR.t1229 26.5955
R10717 VPWR.n2763 VPWR.t1241 26.5955
R10718 VPWR.n2766 VPWR.t1283 26.5955
R10719 VPWR.n2766 VPWR.t1491 26.5955
R10720 VPWR.n2767 VPWR.t1233 26.5955
R10721 VPWR.n2767 VPWR.t1237 26.5955
R10722 VPWR.n2743 VPWR.t548 26.5955
R10723 VPWR.n2743 VPWR.t542 26.5955
R10724 VPWR.n2744 VPWR.t1019 26.5955
R10725 VPWR.n2744 VPWR.t1018 26.5955
R10726 VPWR.n2747 VPWR.t550 26.5955
R10727 VPWR.n2747 VPWR.t552 26.5955
R10728 VPWR.n2748 VPWR.t1021 26.5955
R10729 VPWR.n2748 VPWR.t1015 26.5955
R10730 VPWR.n2708 VPWR.t1779 26.5955
R10731 VPWR.n2708 VPWR.t1811 26.5955
R10732 VPWR.n2712 VPWR.t1803 26.5955
R10733 VPWR.n2712 VPWR.t1370 26.5955
R10734 VPWR.n2715 VPWR.t1777 26.5955
R10735 VPWR.n2715 VPWR.t1825 26.5955
R10736 VPWR.n2709 VPWR.t1364 26.5955
R10737 VPWR.n2709 VPWR.t1372 26.5955
R10738 VPWR.n2679 VPWR.t1773 26.5955
R10739 VPWR.n2679 VPWR.t1823 26.5955
R10740 VPWR.n2678 VPWR.t1789 26.5955
R10741 VPWR.n2678 VPWR.t1835 26.5955
R10742 VPWR.n2675 VPWR.t1800 26.5955
R10743 VPWR.n2675 VPWR.t3 26.5955
R10744 VPWR.n2674 VPWR.t1817 26.5955
R10745 VPWR.n2674 VPWR.t1668 26.5955
R10746 VPWR.n2671 VPWR.t1507 26.5955
R10747 VPWR.n2671 VPWR.t1245 26.5955
R10748 VPWR.n2670 VPWR.t1665 26.5955
R10749 VPWR.n2670 VPWR.t1669 26.5955
R10750 VPWR.n2642 VPWR.t1795 26.5955
R10751 VPWR.n2642 VPWR.t1769 26.5955
R10752 VPWR.n2641 VPWR.t1813 26.5955
R10753 VPWR.n2641 VPWR.t1788 26.5955
R10754 VPWR.n2638 VPWR.t1821 26.5955
R10755 VPWR.n2638 VPWR.t1239 26.5955
R10756 VPWR.n2637 VPWR.t1831 26.5955
R10757 VPWR.n2637 VPWR.t1270 26.5955
R10758 VPWR.n2634 VPWR.t1231 26.5955
R10759 VPWR.n2634 VPWR.t1243 26.5955
R10760 VPWR.n2633 VPWR.t1490 26.5955
R10761 VPWR.n2633 VPWR.t1269 26.5955
R10762 VPWR.n2606 VPWR.t1792 26.5955
R10763 VPWR.n2606 VPWR.t1798 26.5955
R10764 VPWR.n2605 VPWR.t1828 26.5955
R10765 VPWR.n2605 VPWR.t1809 26.5955
R10766 VPWR.n2613 VPWR.t1804 26.5955
R10767 VPWR.n2613 VPWR.t1020 26.5955
R10768 VPWR.n2612 VPWR.t1786 26.5955
R10769 VPWR.n2612 VPWR.t544 26.5955
R10770 VPWR.n2602 VPWR.t1022 26.5955
R10771 VPWR.n2602 VPWR.t1016 26.5955
R10772 VPWR.n2601 VPWR.t538 26.5955
R10773 VPWR.n2601 VPWR.t546 26.5955
R10774 VPWR.n17 VPWR.n16 25.977
R10775 VPWR.n1253 VPWR.n1252 25.977
R10776 VPWR.n1313 VPWR.n1310 25.977
R10777 VPWR.n1349 VPWR.n1346 25.977
R10778 VPWR.n1372 VPWR.n1338 25.977
R10779 VPWR.n1388 VPWR.n1385 25.977
R10780 VPWR.n1425 VPWR.n1422 25.977
R10781 VPWR.n2811 VPWR.n2810 25.977
R10782 VPWR.n2795 VPWR.n2794 25.977
R10783 VPWR.n2717 VPWR.n2714 25.977
R10784 VPWR.n2681 VPWR.n2677 25.977
R10785 VPWR.n2699 VPWR.n2698 25.977
R10786 VPWR.n2644 VPWR.n2640 25.977
R10787 VPWR.n2609 VPWR.n2607 25.977
R10788 VPWR.n1335 VPWR.n1334 25.224
R10789 VPWR.n2737 VPWR.n2736 25.224
R10790 VPWR.n2722 VPWR.n2721 24.8476
R10791 VPWR.n2686 VPWR.n2685 24.8476
R10792 VPWR.n2649 VPWR.n2648 24.8476
R10793 VPWR.n2615 VPWR.n2614 24.8476
R10794 VPWR.n16 VPWR.n15 24.4711
R10795 VPWR.n1252 VPWR.n1251 24.4711
R10796 VPWR.n1315 VPWR.n1313 24.4711
R10797 VPWR.n1352 VPWR.n1349 24.4711
R10798 VPWR.n1391 VPWR.n1388 24.4711
R10799 VPWR.n1428 VPWR.n1425 24.4711
R10800 VPWR.n2810 VPWR.n2809 24.4711
R10801 VPWR.n2794 VPWR.n2793 24.4711
R10802 VPWR.n11 VPWR.n2 23.7181
R10803 VPWR.n1247 VPWR.n1236 23.7181
R10804 VPWR.n1270 VPWR.n1259 23.7181
R10805 VPWR.n1274 VPWR.n1259 23.7181
R10806 VPWR.n1294 VPWR.n1283 23.7181
R10807 VPWR.n1298 VPWR.n1283 23.7181
R10808 VPWR.n1330 VPWR.n1328 23.7181
R10809 VPWR.n1368 VPWR.n1365 23.7181
R10810 VPWR.n1407 VPWR.n1404 23.7181
R10811 VPWR.n1407 VPWR.n1377 23.7181
R10812 VPWR.n1444 VPWR.n1441 23.7181
R10813 VPWR.n2808 VPWR.n2807 23.7181
R10814 VPWR.n2789 VPWR.n2781 23.7181
R10815 VPWR.n2769 VPWR.n2761 23.7181
R10816 VPWR.n2773 VPWR.n2761 23.7181
R10817 VPWR.n2750 VPWR.n2742 23.7181
R10818 VPWR.n2754 VPWR.n2742 23.7181
R10819 VPWR.n2731 VPWR.n2706 23.7181
R10820 VPWR.n2694 VPWR.n2668 23.7181
R10821 VPWR.n2657 VPWR.n2631 23.7181
R10822 VPWR.n2661 VPWR.n2631 23.7181
R10823 VPWR.n2626 VPWR.n2625 23.7181
R10824 VPWR.t978 VPWR.t950 23.4987
R10825 VPWR.t1893 VPWR.t455 23.4987
R10826 VPWR.n2852 VPWR.n2841 23.1255
R10827 VPWR.n2852 VPWR.t1094 23.1255
R10828 VPWR.n2851 VPWR.n2819 23.1255
R10829 VPWR.t1094 VPWR.n2851 23.1255
R10830 VPWR.n11 VPWR.n10 22.9652
R10831 VPWR.n1247 VPWR.n1246 22.9652
R10832 VPWR.n1270 VPWR.n1269 22.9652
R10833 VPWR.n1294 VPWR.n1293 22.9652
R10834 VPWR.n2807 VPWR.n2803 22.9652
R10835 VPWR.n2789 VPWR.n2788 22.9652
R10836 VPWR.n2769 VPWR.n2768 22.9652
R10837 VPWR.n2750 VPWR.n2749 22.9652
R10838 VPWR.n1320 VPWR.n1308 22.2123
R10839 VPWR.n2724 VPWR.n2723 22.2123
R10840 VPWR.n10 VPWR.n3 21.4593
R10841 VPWR.n1246 VPWR.n1237 21.4593
R10842 VPWR.n1269 VPWR.n1260 21.4593
R10843 VPWR.n1293 VPWR.n1284 21.4593
R10844 VPWR.n1442 VPWR.t370 20.5957
R10845 VPWR.n1443 VPWR.t300 20.5957
R10846 VPWR.n1277 VPWR.n1276 19.9534
R10847 VPWR.n1300 VPWR.n1299 19.9534
R10848 VPWR.n1334 VPWR.n1303 19.9534
R10849 VPWR.n2776 VPWR.n2775 19.9534
R10850 VPWR.n2756 VPWR.n2755 19.9534
R10851 VPWR.n2736 VPWR.n2735 19.9534
R10852 VPWR.n2724 VPWR.n2710 18.824
R10853 VPWR.n2688 VPWR.n2672 18.824
R10854 VPWR.n2651 VPWR.n2635 18.824
R10855 VPWR.n2620 VPWR.n2619 18.824
R10856 VPWR.n1316 VPWR.n1308 18.4476
R10857 VPWR.n1353 VPWR.n1345 18.4476
R10858 VPWR.n1373 VPWR.n1372 18.4476
R10859 VPWR.n1392 VPWR.n1384 18.4476
R10860 VPWR.n1429 VPWR.n1421 18.4476
R10861 VPWR.n2700 VPWR.n2699 18.4476
R10862 VPWR.n1413 VPWR.n1412 17.5829
R10863 VPWR.n2664 VPWR.n2663 17.5829
R10864 VPWR.n6 VPWR.n3 16.9417
R10865 VPWR.n1241 VPWR.n1237 16.9417
R10866 VPWR.n1264 VPWR.n1260 16.9417
R10867 VPWR.n1288 VPWR.n1284 16.9417
R10868 VPWR.n2730 VPWR.n2729 16.5652
R10869 VPWR.n1306 VPWR.n1304 16.1887
R10870 VPWR.n1374 VPWR.n1373 16.1887
R10871 VPWR.n2701 VPWR.n2700 16.1887
R10872 VPWR.n1235 VPWR.t364 16.0935
R10873 VPWR.n1258 VPWR.t154 16.0935
R10874 VPWR.n1282 VPWR.t1029 16.0935
R10875 VPWR.n1367 VPWR.t21 16.0935
R10876 VPWR.n1406 VPWR.t0 16.0935
R10877 VPWR.n1234 VPWR.t417 16.0935
R10878 VPWR.n1257 VPWR.t335 16.0935
R10879 VPWR.n1281 VPWR.t302 16.0935
R10880 VPWR.n1366 VPWR.t367 16.0935
R10881 VPWR.n1405 VPWR.t23 16.0935
R10882 VPWR.n1325 VPWR.n1306 15.8123
R10883 VPWR.n2727 VPWR.n2710 15.8123
R10884 VPWR.n2729 VPWR.n2728 15.8123
R10885 VPWR.n2691 VPWR.n2672 15.8123
R10886 VPWR.n2654 VPWR.n2635 15.8123
R10887 VPWR.n2621 VPWR.n2620 15.8123
R10888 VPWR.n1330 VPWR.n1303 13.5534
R10889 VPWR.n2735 VPWR.n2706 13.5534
R10890 VPWR.n2839 VPWR.n2823 13.2148
R10891 VPWR.n2823 VPWR.t93 13.2148
R10892 VPWR.n2827 VPWR.n2817 13.2148
R10893 VPWR.n2827 VPWR.t93 13.2148
R10894 VPWR.n2833 VPWR.n2829 13.2148
R10895 VPWR.n2829 VPWR.t93 13.2148
R10896 VPWR.n15 VPWR.n2 12.8005
R10897 VPWR.n1251 VPWR.n1236 12.8005
R10898 VPWR.n1368 VPWR.n1338 12.8005
R10899 VPWR.n2809 VPWR.n2808 12.8005
R10900 VPWR.n2793 VPWR.n2781 12.8005
R10901 VPWR.n2698 VPWR.n2668 12.8005
R10902 VPWR.n1322 VPWR.n1320 12.424
R10903 VPWR.n1360 VPWR.n1357 12.424
R10904 VPWR.n1399 VPWR.n1396 12.424
R10905 VPWR.n1436 VPWR.n1433 12.424
R10906 VPWR.n1276 VPWR.n1275 10.5417
R10907 VPWR.n1412 VPWR.n1411 10.5417
R10908 VPWR.n2775 VPWR.n2774 10.5417
R10909 VPWR.n2663 VPWR.n2662 10.5417
R10910 VPWR.n2687 VPWR.n2686 9.78874
R10911 VPWR.n2650 VPWR.n2649 9.78874
R10912 VPWR.n2614 VPWR.n2603 9.78874
R10913 VPWR.n1361 VPWR.n1360 9.41227
R10914 VPWR.n1365 VPWR.n1339 9.41227
R10915 VPWR.n1400 VPWR.n1399 9.41227
R10916 VPWR.n1404 VPWR.n1378 9.41227
R10917 VPWR.n1437 VPWR.n1436 9.41227
R10918 VPWR.n1441 VPWR.n1415 9.41227
R10919 VPWR.n2694 VPWR.n2693 9.41227
R10920 VPWR.n2657 VPWR.n2656 9.41227
R10921 VPWR.n2625 VPWR.n2599 9.41227
R10922 VPWR.n1229 VPWR 9.37021
R10923 VPWR.n1151 VPWR 9.37021
R10924 VPWR.n1225 VPWR 9.37021
R10925 VPWR.n1483 VPWR 9.37021
R10926 VPWR.n1171 VPWR 9.37021
R10927 VPWR.n1167 VPWR 9.37021
R10928 VPWR.n1161 VPWR 9.37021
R10929 VPWR.n1477 VPWR 9.37021
R10930 VPWR.n1157 VPWR 9.37021
R10931 VPWR.n1147 VPWR 9.37021
R10932 VPWR.n1470 VPWR 9.37021
R10933 VPWR.n1047 VPWR 9.37021
R10934 VPWR.n1746 VPWR 9.37021
R10935 VPWR.n1034 VPWR 9.37021
R10936 VPWR.n1030 VPWR 9.37021
R10937 VPWR.n1051 VPWR 9.37021
R10938 VPWR.n1467 VPWR.n1466 9.33404
R10939 VPWR.n352 VPWR.n351 9.33404
R10940 VPWR.n1534 VPWR.n1533 9.33404
R10941 VPWR.n348 VPWR.n347 9.33404
R10942 VPWR.n965 VPWR.n964 9.33404
R10943 VPWR.n2479 VPWR.n2478 9.33404
R10944 VPWR.n2475 VPWR.n2474 9.33404
R10945 VPWR.n320 VPWR.n319 9.33404
R10946 VPWR.n973 VPWR.n972 9.33404
R10947 VPWR.n2445 VPWR.n2444 9.33404
R10948 VPWR.n324 VPWR.n323 9.33404
R10949 VPWR.n1891 VPWR.n1890 9.33404
R10950 VPWR.n1887 VPWR.n1886 9.33404
R10951 VPWR.n1881 VPWR.n1880 9.33404
R10952 VPWR.n389 VPWR.n388 9.33404
R10953 VPWR.n393 VPWR.n392 9.33404
R10954 VPWR.n397 VPWR.n396 9.33404
R10955 VPWR.n2455 VPWR.n2454 9.33404
R10956 VPWR.n332 VPWR.n331 9.33404
R10957 VPWR.n1877 VPWR.n1876 9.33404
R10958 VPWR.n405 VPWR.n404 9.33404
R10959 VPWR.n2459 VPWR.n2458 9.33404
R10960 VPWR.n336 VPWR.n335 9.33404
R10961 VPWR.n2308 VPWR.n2307 9.33404
R10962 VPWR.n2312 VPWR.n2311 9.33404
R10963 VPWR.n2318 VPWR.n2317 9.33404
R10964 VPWR.n2322 VPWR.n2321 9.33404
R10965 VPWR.n2332 VPWR.n2331 9.33404
R10966 VPWR.n2338 VPWR.n2337 9.33404
R10967 VPWR.n2342 VPWR.n2341 9.33404
R10968 VPWR.n2348 VPWR.n2347 9.33404
R10969 VPWR.n2352 VPWR.n2351 9.33404
R10970 VPWR.n2358 VPWR.n2357 9.33404
R10971 VPWR.n2362 VPWR.n2361 9.33404
R10972 VPWR.n2368 VPWR.n2367 9.33404
R10973 VPWR.n2372 VPWR.n2371 9.33404
R10974 VPWR.n2378 VPWR.n2377 9.33404
R10975 VPWR.n2381 VPWR.n2380 9.33404
R10976 VPWR.n2328 VPWR.n2327 9.33404
R10977 VPWR.n544 VPWR.n543 9.33404
R10978 VPWR.n540 VPWR.n539 9.33404
R10979 VPWR.n536 VPWR.n535 9.33404
R10980 VPWR.n532 VPWR.n531 9.33404
R10981 VPWR.n524 VPWR.n523 9.33404
R10982 VPWR.n520 VPWR.n519 9.33404
R10983 VPWR.n516 VPWR.n515 9.33404
R10984 VPWR.n512 VPWR.n511 9.33404
R10985 VPWR.n508 VPWR.n507 9.33404
R10986 VPWR.n504 VPWR.n503 9.33404
R10987 VPWR.n500 VPWR.n499 9.33404
R10988 VPWR.n496 VPWR.n495 9.33404
R10989 VPWR.n492 VPWR.n491 9.33404
R10990 VPWR.n488 VPWR.n487 9.33404
R10991 VPWR.n485 VPWR.n484 9.33404
R10992 VPWR.n528 VPWR.n527 9.33404
R10993 VPWR.n2283 VPWR.n2282 9.33404
R10994 VPWR.n2279 VPWR.n2278 9.33404
R10995 VPWR.n2273 VPWR.n2272 9.33404
R10996 VPWR.n2269 VPWR.n2268 9.33404
R10997 VPWR.n2259 VPWR.n2258 9.33404
R10998 VPWR.n2253 VPWR.n2252 9.33404
R10999 VPWR.n2249 VPWR.n2248 9.33404
R11000 VPWR.n2243 VPWR.n2242 9.33404
R11001 VPWR.n2239 VPWR.n2238 9.33404
R11002 VPWR.n2233 VPWR.n2232 9.33404
R11003 VPWR.n2229 VPWR.n2228 9.33404
R11004 VPWR.n2223 VPWR.n2222 9.33404
R11005 VPWR.n2219 VPWR.n2218 9.33404
R11006 VPWR.n2213 VPWR.n2212 9.33404
R11007 VPWR.n2210 VPWR.n2209 9.33404
R11008 VPWR.n2263 VPWR.n2262 9.33404
R11009 VPWR.n581 VPWR.n580 9.33404
R11010 VPWR.n585 VPWR.n584 9.33404
R11011 VPWR.n589 VPWR.n588 9.33404
R11012 VPWR.n593 VPWR.n592 9.33404
R11013 VPWR.n601 VPWR.n600 9.33404
R11014 VPWR.n605 VPWR.n604 9.33404
R11015 VPWR.n609 VPWR.n608 9.33404
R11016 VPWR.n613 VPWR.n612 9.33404
R11017 VPWR.n617 VPWR.n616 9.33404
R11018 VPWR.n621 VPWR.n620 9.33404
R11019 VPWR.n625 VPWR.n624 9.33404
R11020 VPWR.n629 VPWR.n628 9.33404
R11021 VPWR.n633 VPWR.n632 9.33404
R11022 VPWR.n637 VPWR.n636 9.33404
R11023 VPWR.n640 VPWR.n639 9.33404
R11024 VPWR.n597 VPWR.n596 9.33404
R11025 VPWR.n2112 VPWR.n2111 9.33404
R11026 VPWR.n2116 VPWR.n2115 9.33404
R11027 VPWR.n2122 VPWR.n2121 9.33404
R11028 VPWR.n2126 VPWR.n2125 9.33404
R11029 VPWR.n2136 VPWR.n2135 9.33404
R11030 VPWR.n2142 VPWR.n2141 9.33404
R11031 VPWR.n2146 VPWR.n2145 9.33404
R11032 VPWR.n2152 VPWR.n2151 9.33404
R11033 VPWR.n2156 VPWR.n2155 9.33404
R11034 VPWR.n2162 VPWR.n2161 9.33404
R11035 VPWR.n2166 VPWR.n2165 9.33404
R11036 VPWR.n2172 VPWR.n2171 9.33404
R11037 VPWR.n2176 VPWR.n2175 9.33404
R11038 VPWR.n2182 VPWR.n2181 9.33404
R11039 VPWR.n2185 VPWR.n2184 9.33404
R11040 VPWR.n2132 VPWR.n2131 9.33404
R11041 VPWR.n736 VPWR.n735 9.33404
R11042 VPWR.n732 VPWR.n731 9.33404
R11043 VPWR.n728 VPWR.n727 9.33404
R11044 VPWR.n724 VPWR.n723 9.33404
R11045 VPWR.n716 VPWR.n715 9.33404
R11046 VPWR.n712 VPWR.n711 9.33404
R11047 VPWR.n708 VPWR.n707 9.33404
R11048 VPWR.n704 VPWR.n703 9.33404
R11049 VPWR.n700 VPWR.n699 9.33404
R11050 VPWR.n696 VPWR.n695 9.33404
R11051 VPWR.n692 VPWR.n691 9.33404
R11052 VPWR.n688 VPWR.n687 9.33404
R11053 VPWR.n684 VPWR.n683 9.33404
R11054 VPWR.n680 VPWR.n679 9.33404
R11055 VPWR.n677 VPWR.n676 9.33404
R11056 VPWR.n720 VPWR.n719 9.33404
R11057 VPWR.n2087 VPWR.n2086 9.33404
R11058 VPWR.n2083 VPWR.n2082 9.33404
R11059 VPWR.n2077 VPWR.n2076 9.33404
R11060 VPWR.n2073 VPWR.n2072 9.33404
R11061 VPWR.n2063 VPWR.n2062 9.33404
R11062 VPWR.n2057 VPWR.n2056 9.33404
R11063 VPWR.n2053 VPWR.n2052 9.33404
R11064 VPWR.n2047 VPWR.n2046 9.33404
R11065 VPWR.n2043 VPWR.n2042 9.33404
R11066 VPWR.n2037 VPWR.n2036 9.33404
R11067 VPWR.n2033 VPWR.n2032 9.33404
R11068 VPWR.n2027 VPWR.n2026 9.33404
R11069 VPWR.n2023 VPWR.n2022 9.33404
R11070 VPWR.n2017 VPWR.n2016 9.33404
R11071 VPWR.n2014 VPWR.n2013 9.33404
R11072 VPWR.n2067 VPWR.n2066 9.33404
R11073 VPWR.n773 VPWR.n772 9.33404
R11074 VPWR.n777 VPWR.n776 9.33404
R11075 VPWR.n781 VPWR.n780 9.33404
R11076 VPWR.n785 VPWR.n784 9.33404
R11077 VPWR.n793 VPWR.n792 9.33404
R11078 VPWR.n797 VPWR.n796 9.33404
R11079 VPWR.n801 VPWR.n800 9.33404
R11080 VPWR.n805 VPWR.n804 9.33404
R11081 VPWR.n809 VPWR.n808 9.33404
R11082 VPWR.n813 VPWR.n812 9.33404
R11083 VPWR.n817 VPWR.n816 9.33404
R11084 VPWR.n821 VPWR.n820 9.33404
R11085 VPWR.n825 VPWR.n824 9.33404
R11086 VPWR.n829 VPWR.n828 9.33404
R11087 VPWR.n832 VPWR.n831 9.33404
R11088 VPWR.n789 VPWR.n788 9.33404
R11089 VPWR.n1916 VPWR.n1915 9.33404
R11090 VPWR.n1920 VPWR.n1919 9.33404
R11091 VPWR.n1926 VPWR.n1925 9.33404
R11092 VPWR.n1930 VPWR.n1929 9.33404
R11093 VPWR.n1940 VPWR.n1939 9.33404
R11094 VPWR.n1946 VPWR.n1945 9.33404
R11095 VPWR.n1950 VPWR.n1949 9.33404
R11096 VPWR.n1956 VPWR.n1955 9.33404
R11097 VPWR.n1960 VPWR.n1959 9.33404
R11098 VPWR.n1966 VPWR.n1965 9.33404
R11099 VPWR.n1970 VPWR.n1969 9.33404
R11100 VPWR.n1976 VPWR.n1975 9.33404
R11101 VPWR.n1980 VPWR.n1979 9.33404
R11102 VPWR.n1986 VPWR.n1985 9.33404
R11103 VPWR.n1989 VPWR.n1988 9.33404
R11104 VPWR.n1936 VPWR.n1935 9.33404
R11105 VPWR.n928 VPWR.n927 9.33404
R11106 VPWR.n924 VPWR.n923 9.33404
R11107 VPWR.n920 VPWR.n919 9.33404
R11108 VPWR.n916 VPWR.n915 9.33404
R11109 VPWR.n908 VPWR.n907 9.33404
R11110 VPWR.n904 VPWR.n903 9.33404
R11111 VPWR.n900 VPWR.n899 9.33404
R11112 VPWR.n896 VPWR.n895 9.33404
R11113 VPWR.n892 VPWR.n891 9.33404
R11114 VPWR.n888 VPWR.n887 9.33404
R11115 VPWR.n884 VPWR.n883 9.33404
R11116 VPWR.n880 VPWR.n879 9.33404
R11117 VPWR.n876 VPWR.n875 9.33404
R11118 VPWR.n872 VPWR.n871 9.33404
R11119 VPWR.n869 VPWR.n868 9.33404
R11120 VPWR.n912 VPWR.n911 9.33404
R11121 VPWR.n1871 VPWR.n1870 9.33404
R11122 VPWR.n981 VPWR.n980 9.33404
R11123 VPWR.n1495 VPWR.n1494 9.33404
R11124 VPWR.n401 VPWR.n400 9.33404
R11125 VPWR.n2465 VPWR.n2464 9.33404
R11126 VPWR.n340 VPWR.n339 9.33404
R11127 VPWR.n977 VPWR.n976 9.33404
R11128 VPWR.n1491 VPWR.n1490 9.33404
R11129 VPWR.n1867 VPWR.n1866 9.33404
R11130 VPWR.n985 VPWR.n984 9.33404
R11131 VPWR.n1505 VPWR.n1504 9.33404
R11132 VPWR.n409 VPWR.n408 9.33404
R11133 VPWR.n417 VPWR.n416 9.33404
R11134 VPWR.n421 VPWR.n420 9.33404
R11135 VPWR.n425 VPWR.n424 9.33404
R11136 VPWR.n429 VPWR.n428 9.33404
R11137 VPWR.n433 VPWR.n432 9.33404
R11138 VPWR.n437 VPWR.n436 9.33404
R11139 VPWR.n441 VPWR.n440 9.33404
R11140 VPWR.n445 VPWR.n444 9.33404
R11141 VPWR.n448 VPWR.n447 9.33404
R11142 VPWR.n413 VPWR.n412 9.33404
R11143 VPWR.n2449 VPWR.n2448 9.33404
R11144 VPWR.n328 VPWR.n327 9.33404
R11145 VPWR.n989 VPWR.n988 9.33404
R11146 VPWR.n1509 VPWR.n1508 9.33404
R11147 VPWR.n1861 VPWR.n1860 9.33404
R11148 VPWR.n1851 VPWR.n1850 9.33404
R11149 VPWR.n1847 VPWR.n1846 9.33404
R11150 VPWR.n1841 VPWR.n1840 9.33404
R11151 VPWR.n1837 VPWR.n1836 9.33404
R11152 VPWR.n1831 VPWR.n1830 9.33404
R11153 VPWR.n1827 VPWR.n1826 9.33404
R11154 VPWR.n1821 VPWR.n1820 9.33404
R11155 VPWR.n1818 VPWR.n1817 9.33404
R11156 VPWR.n1857 VPWR.n1856 9.33404
R11157 VPWR.n993 VPWR.n992 9.33404
R11158 VPWR.n1519 VPWR.n1518 9.33404
R11159 VPWR.n2469 VPWR.n2468 9.33404
R11160 VPWR.n344 VPWR.n343 9.33404
R11161 VPWR.n1480 VPWR.n1130 9.33404
R11162 VPWR.n997 VPWR.n996 9.33404
R11163 VPWR.n1523 VPWR.n1522 9.33404
R11164 VPWR.n2439 VPWR.n2438 9.33404
R11165 VPWR.n2429 VPWR.n2428 9.33404
R11166 VPWR.n2425 VPWR.n2424 9.33404
R11167 VPWR.n2419 VPWR.n2418 9.33404
R11168 VPWR.n2415 VPWR.n2414 9.33404
R11169 VPWR.n2409 VPWR.n2408 9.33404
R11170 VPWR.n2406 VPWR.n2405 9.33404
R11171 VPWR.n2435 VPWR.n2434 9.33404
R11172 VPWR.n316 VPWR.n315 9.33404
R11173 VPWR.n1538 VPWR.n1537 9.33404
R11174 VPWR.n1001 VPWR.n1000 9.33404
R11175 VPWR.n1005 VPWR.n1004 9.33404
R11176 VPWR.n1009 VPWR.n1008 9.33404
R11177 VPWR.n1013 VPWR.n1012 9.33404
R11178 VPWR.n1017 VPWR.n1016 9.33404
R11179 VPWR.n1021 VPWR.n1020 9.33404
R11180 VPWR.n1024 VPWR.n1023 9.33404
R11181 VPWR.n969 VPWR.n968 9.33404
R11182 VPWR.n1474 VPWR.n1473 9.33404
R11183 VPWR.n312 VPWR.n311 9.33404
R11184 VPWR.n1763 VPWR.n1762 9.33404
R11185 VPWR.n308 VPWR.n307 9.33404
R11186 VPWR.n304 VPWR.n303 9.33404
R11187 VPWR.n296 VPWR.n295 9.33404
R11188 VPWR.n293 VPWR.n292 9.33404
R11189 VPWR.n300 VPWR.n299 9.33404
R11190 VPWR.n1751 VPWR.n1750 9.33404
R11191 VPWR.n1790 VPWR.n1789 9.33404
R11192 VPWR.n1793 VPWR.n1792 9.33404
R11193 VPWR.n1759 VPWR.n1758 9.33404
R11194 VPWR.n2714 VPWR 9.32394
R11195 VPWR.n2677 VPWR 9.32394
R11196 VPWR.n2640 VPWR 9.32394
R11197 VPWR VPWR.n2607 9.32394
R11198 VPWR.n18 VPWR.n17 9.3005
R11199 VPWR.n15 VPWR.n14 9.3005
R11200 VPWR.n13 VPWR.n2 9.3005
R11201 VPWR.n10 VPWR.n9 9.3005
R11202 VPWR.n8 VPWR.n3 9.3005
R11203 VPWR.n12 VPWR.n11 9.3005
R11204 VPWR.n16 VPWR.n0 9.3005
R11205 VPWR.n1254 VPWR.n1253 9.3005
R11206 VPWR.n1251 VPWR.n1250 9.3005
R11207 VPWR.n1249 VPWR.n1236 9.3005
R11208 VPWR.n1246 VPWR.n1244 9.3005
R11209 VPWR.n1243 VPWR.n1237 9.3005
R11210 VPWR.n1248 VPWR.n1247 9.3005
R11211 VPWR.n1252 VPWR.n1233 9.3005
R11212 VPWR.n1278 VPWR.n1277 9.3005
R11213 VPWR.n1272 VPWR.n1259 9.3005
R11214 VPWR.n1269 VPWR.n1267 9.3005
R11215 VPWR.n1266 VPWR.n1260 9.3005
R11216 VPWR.n1271 VPWR.n1270 9.3005
R11217 VPWR.n1274 VPWR.n1273 9.3005
R11218 VPWR.n1276 VPWR.n1256 9.3005
R11219 VPWR.n1301 VPWR.n1300 9.3005
R11220 VPWR.n1296 VPWR.n1283 9.3005
R11221 VPWR.n1293 VPWR.n1291 9.3005
R11222 VPWR.n1290 VPWR.n1284 9.3005
R11223 VPWR.n1295 VPWR.n1294 9.3005
R11224 VPWR.n1298 VPWR.n1297 9.3005
R11225 VPWR.n1299 VPWR.n1280 9.3005
R11226 VPWR.n1332 VPWR.n1303 9.3005
R11227 VPWR.n1331 VPWR.n1330 9.3005
R11228 VPWR.n1311 VPWR.n1310 9.3005
R11229 VPWR.n1313 VPWR.n1312 9.3005
R11230 VPWR.n1315 VPWR.n1309 9.3005
R11231 VPWR.n1317 VPWR.n1316 9.3005
R11232 VPWR.n1318 VPWR.n1308 9.3005
R11233 VPWR.n1320 VPWR.n1319 9.3005
R11234 VPWR.n1324 VPWR.n1305 9.3005
R11235 VPWR.n1326 VPWR.n1325 9.3005
R11236 VPWR.n1328 VPWR.n1327 9.3005
R11237 VPWR.n1334 VPWR.n1333 9.3005
R11238 VPWR.n1336 VPWR.n1335 9.3005
R11239 VPWR.n1375 VPWR.n1374 9.3005
R11240 VPWR.n1370 VPWR.n1338 9.3005
R11241 VPWR.n1369 VPWR.n1368 9.3005
R11242 VPWR.n1347 VPWR.n1346 9.3005
R11243 VPWR.n1349 VPWR.n1348 9.3005
R11244 VPWR.n1352 VPWR.n1342 9.3005
R11245 VPWR.n1354 VPWR.n1353 9.3005
R11246 VPWR.n1355 VPWR.n1341 9.3005
R11247 VPWR.n1357 VPWR.n1356 9.3005
R11248 VPWR.n1361 VPWR.n1340 9.3005
R11249 VPWR.n1363 VPWR.n1362 9.3005
R11250 VPWR.n1365 VPWR.n1364 9.3005
R11251 VPWR.n1372 VPWR.n1371 9.3005
R11252 VPWR.n1408 VPWR.n1407 9.3005
R11253 VPWR.n1386 VPWR.n1385 9.3005
R11254 VPWR.n1388 VPWR.n1387 9.3005
R11255 VPWR.n1391 VPWR.n1381 9.3005
R11256 VPWR.n1393 VPWR.n1392 9.3005
R11257 VPWR.n1394 VPWR.n1380 9.3005
R11258 VPWR.n1396 VPWR.n1395 9.3005
R11259 VPWR.n1400 VPWR.n1379 9.3005
R11260 VPWR.n1402 VPWR.n1401 9.3005
R11261 VPWR.n1404 VPWR.n1403 9.3005
R11262 VPWR.n1409 VPWR.n1377 9.3005
R11263 VPWR.n1411 VPWR.n1410 9.3005
R11264 VPWR.n1445 VPWR.n1444 9.3005
R11265 VPWR.n1423 VPWR.n1422 9.3005
R11266 VPWR.n1425 VPWR.n1424 9.3005
R11267 VPWR.n1428 VPWR.n1418 9.3005
R11268 VPWR.n1430 VPWR.n1429 9.3005
R11269 VPWR.n1431 VPWR.n1417 9.3005
R11270 VPWR.n1433 VPWR.n1432 9.3005
R11271 VPWR.n1437 VPWR.n1416 9.3005
R11272 VPWR.n1439 VPWR.n1438 9.3005
R11273 VPWR.n1441 VPWR.n1440 9.3005
R11274 VPWR.n2807 VPWR.n2806 9.3005
R11275 VPWR.n2808 VPWR.n2800 9.3005
R11276 VPWR.n2809 VPWR.n2799 9.3005
R11277 VPWR.n2810 VPWR.n2798 9.3005
R11278 VPWR.n2812 VPWR.n2811 9.3005
R11279 VPWR.n2796 VPWR.n2795 9.3005
R11280 VPWR.n2790 VPWR.n2789 9.3005
R11281 VPWR.n2791 VPWR.n2781 9.3005
R11282 VPWR.n2793 VPWR.n2792 9.3005
R11283 VPWR.n2794 VPWR.n2779 9.3005
R11284 VPWR.n2777 VPWR.n2776 9.3005
R11285 VPWR.n2775 VPWR.n2759 9.3005
R11286 VPWR.n2770 VPWR.n2769 9.3005
R11287 VPWR.n2771 VPWR.n2761 9.3005
R11288 VPWR.n2773 VPWR.n2772 9.3005
R11289 VPWR.n2757 VPWR.n2756 9.3005
R11290 VPWR.n2751 VPWR.n2750 9.3005
R11291 VPWR.n2752 VPWR.n2742 9.3005
R11292 VPWR.n2754 VPWR.n2753 9.3005
R11293 VPWR.n2755 VPWR.n2740 9.3005
R11294 VPWR.n2738 VPWR.n2737 9.3005
R11295 VPWR.n2718 VPWR.n2717 9.3005
R11296 VPWR.n2719 VPWR.n2713 9.3005
R11297 VPWR.n2721 VPWR.n2720 9.3005
R11298 VPWR.n2723 VPWR.n2711 9.3005
R11299 VPWR.n2725 VPWR.n2724 9.3005
R11300 VPWR.n2727 VPWR.n2726 9.3005
R11301 VPWR.n2728 VPWR.n2707 9.3005
R11302 VPWR.n2732 VPWR.n2731 9.3005
R11303 VPWR.n2733 VPWR.n2706 9.3005
R11304 VPWR.n2735 VPWR.n2734 9.3005
R11305 VPWR.n2736 VPWR.n2704 9.3005
R11306 VPWR.n2702 VPWR.n2701 9.3005
R11307 VPWR.n2682 VPWR.n2681 9.3005
R11308 VPWR.n2683 VPWR.n2676 9.3005
R11309 VPWR.n2685 VPWR.n2684 9.3005
R11310 VPWR.n2687 VPWR.n2673 9.3005
R11311 VPWR.n2689 VPWR.n2688 9.3005
R11312 VPWR.n2691 VPWR.n2690 9.3005
R11313 VPWR.n2692 VPWR.n2669 9.3005
R11314 VPWR.n2695 VPWR.n2694 9.3005
R11315 VPWR.n2696 VPWR.n2668 9.3005
R11316 VPWR.n2698 VPWR.n2697 9.3005
R11317 VPWR.n2699 VPWR.n2666 9.3005
R11318 VPWR.n2645 VPWR.n2644 9.3005
R11319 VPWR.n2646 VPWR.n2639 9.3005
R11320 VPWR.n2648 VPWR.n2647 9.3005
R11321 VPWR.n2650 VPWR.n2636 9.3005
R11322 VPWR.n2652 VPWR.n2651 9.3005
R11323 VPWR.n2654 VPWR.n2653 9.3005
R11324 VPWR.n2655 VPWR.n2632 9.3005
R11325 VPWR.n2658 VPWR.n2657 9.3005
R11326 VPWR.n2659 VPWR.n2631 9.3005
R11327 VPWR.n2661 VPWR.n2660 9.3005
R11328 VPWR.n2662 VPWR.n2629 9.3005
R11329 VPWR.n2627 VPWR.n2626 9.3005
R11330 VPWR.n2609 VPWR.n2608 9.3005
R11331 VPWR.n2611 VPWR.n2604 9.3005
R11332 VPWR.n2616 VPWR.n2615 9.3005
R11333 VPWR.n2617 VPWR.n2603 9.3005
R11334 VPWR.n2619 VPWR.n2618 9.3005
R11335 VPWR.n2621 VPWR.n2600 9.3005
R11336 VPWR.n2623 VPWR.n2622 9.3005
R11337 VPWR.n2625 VPWR.n2624 9.3005
R11338 VPWR.n2505 VPWR.n2504 9.3005
R11339 VPWR.n2569 VPWR.n2568 9.3005
R11340 VPWR.n2509 VPWR.n2508 9.3005
R11341 VPWR.n2553 VPWR.n2552 9.3005
R11342 VPWR.n2545 VPWR.n2544 9.3005
R11343 VPWR.n2533 VPWR.n2532 9.3005
R11344 VPWR.n2529 VPWR.n2528 9.3005
R11345 VPWR.n1222 VPWR.n1221 9.3005
R11346 VPWR.n2521 VPWR.n2520 9.3005
R11347 VPWR.n1184 VPWR.n1102 9.3005
R11348 VPWR.n1218 VPWR.n1094 9.3005
R11349 VPWR.n2541 VPWR.n2540 9.3005
R11350 VPWR.n1215 VPWR.n1092 9.3005
R11351 VPWR.n1212 VPWR.n1211 9.3005
R11352 VPWR.n2517 VPWR.n2516 9.3005
R11353 VPWR.n1181 VPWR.n1104 9.3005
R11354 VPWR.n1204 VPWR.n1084 9.3005
R11355 VPWR.n2557 VPWR.n2556 9.3005
R11356 VPWR.n1201 VPWR.n1082 9.3005
R11357 VPWR.n1592 VPWR.n1591 9.3005
R11358 VPWR.n2565 VPWR.n2564 9.3005
R11359 VPWR.n1198 VPWR.n1197 9.3005
R11360 VPWR.n1190 VPWR.n1074 9.3005
R11361 VPWR.n1742 VPWR.n1741 9.3005
R11362 VPWR.n1187 VPWR.n1071 9.3005
R11363 VPWR.n2577 VPWR.n2576 9.3005
R11364 VPWR.n2581 VPWR.n2580 9.3005
R11365 VPWR.n2592 VPWR.n2591 9.3005
R11366 VPWR.n2589 VPWR.n2588 9.3005
R11367 VPWR.n1738 VPWR.n1737 9.3005
R11368 VPWR.n1063 VPWR.n1062 9.3005
R11369 VPWR.n1596 VPWR.n1595 9.3005
R11370 VPWR.n1275 VPWR.n1274 8.28285
R11371 VPWR.n2774 VPWR.n2773 8.28285
R11372 VPWR.n1607 VPWR.n1109 8.25914
R11373 VPWR.n1728 VPWR.n1727 8.25914
R11374 VPWR.n281 VPWR.n113 8.25914
R11375 VPWR.n136 VPWR.n124 8.25914
R11376 VPWR.n1780 VPWR.n1779 7.91351
R11377 VPWR.n1771 VPWR.n1770 7.9105
R11378 VPWR.n1042 VPWR.n1041 7.9105
R11379 VPWR.n1546 VPWR.n1545 7.9105
R11380 VPWR.n1551 VPWR.n1550 7.9105
R11381 VPWR.n1556 VPWR.n1555 7.9105
R11382 VPWR.n1561 VPWR.n1560 7.9105
R11383 VPWR.n1566 VPWR.n1565 7.9105
R11384 VPWR.n1571 VPWR.n1570 7.9105
R11385 VPWR.n1576 VPWR.n1575 7.9105
R11386 VPWR.n1581 VPWR.n1580 7.9105
R11387 VPWR.n1136 VPWR.n1135 7.9105
R11388 VPWR.n1461 VPWR.n1460 7.9105
R11389 VPWR.n1456 VPWR.n1455 7.9105
R11390 VPWR.n1776 VPWR.n1775 7.9105
R11391 VPWR.n1784 VPWR.n1783 7.9105
R11392 VPWR.n282 VPWR.n281 7.9105
R11393 VPWR.n280 VPWR.n279 7.9105
R11394 VPWR.n268 VPWR.n267 7.9105
R11395 VPWR.n256 VPWR.n255 7.9105
R11396 VPWR.n244 VPWR.n243 7.9105
R11397 VPWR.n232 VPWR.n231 7.9105
R11398 VPWR.n220 VPWR.n219 7.9105
R11399 VPWR.n208 VPWR.n207 7.9105
R11400 VPWR.n196 VPWR.n195 7.9105
R11401 VPWR.n184 VPWR.n183 7.9105
R11402 VPWR.n172 VPWR.n171 7.9105
R11403 VPWR.n160 VPWR.n159 7.9105
R11404 VPWR.n148 VPWR.n147 7.9105
R11405 VPWR.n136 VPWR.n135 7.9105
R11406 VPWR.n1727 VPWR.n1726 7.9105
R11407 VPWR.n1715 VPWR.n1714 7.9105
R11408 VPWR.n1701 VPWR.n1068 7.9105
R11409 VPWR.n1690 VPWR.n1689 7.9105
R11410 VPWR.n1688 VPWR.n1687 7.9105
R11411 VPWR.n1674 VPWR.n1079 7.9105
R11412 VPWR.n1663 VPWR.n1662 7.9105
R11413 VPWR.n1661 VPWR.n1660 7.9105
R11414 VPWR.n1647 VPWR.n1089 7.9105
R11415 VPWR.n1636 VPWR.n1635 7.9105
R11416 VPWR.n1634 VPWR.n1633 7.9105
R11417 VPWR.n1620 VPWR.n1099 7.9105
R11418 VPWR.n1609 VPWR.n1608 7.9105
R11419 VPWR.n1607 VPWR.n1606 7.9105
R11420 VPWR.n26 VPWR.n24 7.8627
R11421 VPWR.n7 VPWR.n6 7.56315
R11422 VPWR.n1242 VPWR.n1241 7.56315
R11423 VPWR.n1265 VPWR.n1264 7.56315
R11424 VPWR.n1289 VPWR.n1288 7.56315
R11425 VPWR.n2805 VPWR.n2803 6.4511
R11426 VPWR.n2788 VPWR.n2785 6.4511
R11427 VPWR.n2768 VPWR.n2765 6.4511
R11428 VPWR.n2749 VPWR.n2746 6.4511
R11429 VPWR.n1362 VPWR.n1339 6.4005
R11430 VPWR.n1401 VPWR.n1378 6.4005
R11431 VPWR.n1438 VPWR.n1415 6.4005
R11432 VPWR.n2723 VPWR.n2722 6.4005
R11433 VPWR.n2693 VPWR.n2692 6.4005
R11434 VPWR.n2656 VPWR.n2655 6.4005
R11435 VPWR.n2622 VPWR.n2599 6.4005
R11436 VPWR.n1595 VPWR.n1122 6.04494
R11437 VPWR.n2505 VPWR.n99 6.04494
R11438 VPWR.n1467 VPWR.n1231 6.04494
R11439 VPWR.n351 VPWR.n290 6.04494
R11440 VPWR.n2568 VPWR.n68 6.04494
R11441 VPWR.n1534 VPWR.n1153 6.04494
R11442 VPWR.n348 VPWR.n346 6.04494
R11443 VPWR.n2508 VPWR.n98 6.04494
R11444 VPWR.n965 VPWR.n963 6.04494
R11445 VPWR.n2478 VPWR.n356 6.04494
R11446 VPWR.n2475 VPWR.n357 6.04494
R11447 VPWR.n320 VPWR.n318 6.04494
R11448 VPWR.n2553 VPWR.n75 6.04494
R11449 VPWR.n973 VPWR.n971 6.04494
R11450 VPWR.n2445 VPWR.n369 6.04494
R11451 VPWR.n324 VPWR.n322 6.04494
R11452 VPWR.n2544 VPWR.n80 6.04494
R11453 VPWR.n1890 VPWR.n932 6.04494
R11454 VPWR.n1887 VPWR.n933 6.04494
R11455 VPWR.n1880 VPWR.n936 6.04494
R11456 VPWR.n389 VPWR.n387 6.04494
R11457 VPWR.n393 VPWR.n391 6.04494
R11458 VPWR.n397 VPWR.n395 6.04494
R11459 VPWR.n2455 VPWR.n365 6.04494
R11460 VPWR.n332 VPWR.n330 6.04494
R11461 VPWR.n2532 VPWR.n86 6.04494
R11462 VPWR.n1877 VPWR.n937 6.04494
R11463 VPWR.n405 VPWR.n403 6.04494
R11464 VPWR.n2458 VPWR.n364 6.04494
R11465 VPWR.n336 VPWR.n334 6.04494
R11466 VPWR.n2529 VPWR.n87 6.04494
R11467 VPWR.n2308 VPWR.n481 6.04494
R11468 VPWR.n2311 VPWR.n480 6.04494
R11469 VPWR.n2318 VPWR.n477 6.04494
R11470 VPWR.n2321 VPWR.n476 6.04494
R11471 VPWR.n2331 VPWR.n472 6.04494
R11472 VPWR.n2338 VPWR.n469 6.04494
R11473 VPWR.n2341 VPWR.n468 6.04494
R11474 VPWR.n2348 VPWR.n465 6.04494
R11475 VPWR.n2351 VPWR.n464 6.04494
R11476 VPWR.n2358 VPWR.n461 6.04494
R11477 VPWR.n2361 VPWR.n460 6.04494
R11478 VPWR.n2368 VPWR.n457 6.04494
R11479 VPWR.n2371 VPWR.n456 6.04494
R11480 VPWR.n2378 VPWR.n453 6.04494
R11481 VPWR.n2380 VPWR.n452 6.04494
R11482 VPWR.n2328 VPWR.n473 6.04494
R11483 VPWR.n543 VPWR.n482 6.04494
R11484 VPWR.n540 VPWR.n538 6.04494
R11485 VPWR.n536 VPWR.n534 6.04494
R11486 VPWR.n532 VPWR.n530 6.04494
R11487 VPWR.n524 VPWR.n522 6.04494
R11488 VPWR.n520 VPWR.n518 6.04494
R11489 VPWR.n516 VPWR.n514 6.04494
R11490 VPWR.n512 VPWR.n510 6.04494
R11491 VPWR.n508 VPWR.n506 6.04494
R11492 VPWR.n504 VPWR.n502 6.04494
R11493 VPWR.n500 VPWR.n498 6.04494
R11494 VPWR.n496 VPWR.n494 6.04494
R11495 VPWR.n492 VPWR.n490 6.04494
R11496 VPWR.n488 VPWR.n486 6.04494
R11497 VPWR.n485 VPWR.n483 6.04494
R11498 VPWR.n528 VPWR.n526 6.04494
R11499 VPWR.n2282 VPWR.n548 6.04494
R11500 VPWR.n2279 VPWR.n549 6.04494
R11501 VPWR.n2272 VPWR.n552 6.04494
R11502 VPWR.n2269 VPWR.n553 6.04494
R11503 VPWR.n2259 VPWR.n557 6.04494
R11504 VPWR.n2252 VPWR.n560 6.04494
R11505 VPWR.n2249 VPWR.n561 6.04494
R11506 VPWR.n2242 VPWR.n564 6.04494
R11507 VPWR.n2239 VPWR.n565 6.04494
R11508 VPWR.n2232 VPWR.n568 6.04494
R11509 VPWR.n2229 VPWR.n569 6.04494
R11510 VPWR.n2222 VPWR.n572 6.04494
R11511 VPWR.n2219 VPWR.n573 6.04494
R11512 VPWR.n2212 VPWR.n576 6.04494
R11513 VPWR.n2210 VPWR.n577 6.04494
R11514 VPWR.n2262 VPWR.n556 6.04494
R11515 VPWR.n581 VPWR.n579 6.04494
R11516 VPWR.n585 VPWR.n583 6.04494
R11517 VPWR.n589 VPWR.n587 6.04494
R11518 VPWR.n593 VPWR.n591 6.04494
R11519 VPWR.n601 VPWR.n599 6.04494
R11520 VPWR.n605 VPWR.n603 6.04494
R11521 VPWR.n609 VPWR.n607 6.04494
R11522 VPWR.n613 VPWR.n611 6.04494
R11523 VPWR.n617 VPWR.n615 6.04494
R11524 VPWR.n621 VPWR.n619 6.04494
R11525 VPWR.n625 VPWR.n623 6.04494
R11526 VPWR.n629 VPWR.n627 6.04494
R11527 VPWR.n633 VPWR.n631 6.04494
R11528 VPWR.n637 VPWR.n635 6.04494
R11529 VPWR.n639 VPWR.n578 6.04494
R11530 VPWR.n597 VPWR.n595 6.04494
R11531 VPWR.n2112 VPWR.n673 6.04494
R11532 VPWR.n2115 VPWR.n672 6.04494
R11533 VPWR.n2122 VPWR.n669 6.04494
R11534 VPWR.n2125 VPWR.n668 6.04494
R11535 VPWR.n2135 VPWR.n664 6.04494
R11536 VPWR.n2142 VPWR.n661 6.04494
R11537 VPWR.n2145 VPWR.n660 6.04494
R11538 VPWR.n2152 VPWR.n657 6.04494
R11539 VPWR.n2155 VPWR.n656 6.04494
R11540 VPWR.n2162 VPWR.n653 6.04494
R11541 VPWR.n2165 VPWR.n652 6.04494
R11542 VPWR.n2172 VPWR.n649 6.04494
R11543 VPWR.n2175 VPWR.n648 6.04494
R11544 VPWR.n2182 VPWR.n645 6.04494
R11545 VPWR.n2184 VPWR.n644 6.04494
R11546 VPWR.n2132 VPWR.n665 6.04494
R11547 VPWR.n735 VPWR.n674 6.04494
R11548 VPWR.n732 VPWR.n730 6.04494
R11549 VPWR.n728 VPWR.n726 6.04494
R11550 VPWR.n724 VPWR.n722 6.04494
R11551 VPWR.n716 VPWR.n714 6.04494
R11552 VPWR.n712 VPWR.n710 6.04494
R11553 VPWR.n708 VPWR.n706 6.04494
R11554 VPWR.n704 VPWR.n702 6.04494
R11555 VPWR.n700 VPWR.n698 6.04494
R11556 VPWR.n696 VPWR.n694 6.04494
R11557 VPWR.n692 VPWR.n690 6.04494
R11558 VPWR.n688 VPWR.n686 6.04494
R11559 VPWR.n684 VPWR.n682 6.04494
R11560 VPWR.n680 VPWR.n678 6.04494
R11561 VPWR.n677 VPWR.n675 6.04494
R11562 VPWR.n720 VPWR.n718 6.04494
R11563 VPWR.n2086 VPWR.n740 6.04494
R11564 VPWR.n2083 VPWR.n741 6.04494
R11565 VPWR.n2076 VPWR.n744 6.04494
R11566 VPWR.n2073 VPWR.n745 6.04494
R11567 VPWR.n2063 VPWR.n749 6.04494
R11568 VPWR.n2056 VPWR.n752 6.04494
R11569 VPWR.n2053 VPWR.n753 6.04494
R11570 VPWR.n2046 VPWR.n756 6.04494
R11571 VPWR.n2043 VPWR.n757 6.04494
R11572 VPWR.n2036 VPWR.n760 6.04494
R11573 VPWR.n2033 VPWR.n761 6.04494
R11574 VPWR.n2026 VPWR.n764 6.04494
R11575 VPWR.n2023 VPWR.n765 6.04494
R11576 VPWR.n2016 VPWR.n768 6.04494
R11577 VPWR.n2014 VPWR.n769 6.04494
R11578 VPWR.n2066 VPWR.n748 6.04494
R11579 VPWR.n773 VPWR.n771 6.04494
R11580 VPWR.n777 VPWR.n775 6.04494
R11581 VPWR.n781 VPWR.n779 6.04494
R11582 VPWR.n785 VPWR.n783 6.04494
R11583 VPWR.n793 VPWR.n791 6.04494
R11584 VPWR.n797 VPWR.n795 6.04494
R11585 VPWR.n801 VPWR.n799 6.04494
R11586 VPWR.n805 VPWR.n803 6.04494
R11587 VPWR.n809 VPWR.n807 6.04494
R11588 VPWR.n813 VPWR.n811 6.04494
R11589 VPWR.n817 VPWR.n815 6.04494
R11590 VPWR.n821 VPWR.n819 6.04494
R11591 VPWR.n825 VPWR.n823 6.04494
R11592 VPWR.n829 VPWR.n827 6.04494
R11593 VPWR.n831 VPWR.n770 6.04494
R11594 VPWR.n789 VPWR.n787 6.04494
R11595 VPWR.n1916 VPWR.n865 6.04494
R11596 VPWR.n1919 VPWR.n864 6.04494
R11597 VPWR.n1926 VPWR.n861 6.04494
R11598 VPWR.n1929 VPWR.n860 6.04494
R11599 VPWR.n1939 VPWR.n856 6.04494
R11600 VPWR.n1946 VPWR.n853 6.04494
R11601 VPWR.n1949 VPWR.n852 6.04494
R11602 VPWR.n1956 VPWR.n849 6.04494
R11603 VPWR.n1959 VPWR.n848 6.04494
R11604 VPWR.n1966 VPWR.n845 6.04494
R11605 VPWR.n1969 VPWR.n844 6.04494
R11606 VPWR.n1976 VPWR.n841 6.04494
R11607 VPWR.n1979 VPWR.n840 6.04494
R11608 VPWR.n1986 VPWR.n837 6.04494
R11609 VPWR.n1988 VPWR.n836 6.04494
R11610 VPWR.n1936 VPWR.n857 6.04494
R11611 VPWR.n927 VPWR.n866 6.04494
R11612 VPWR.n924 VPWR.n922 6.04494
R11613 VPWR.n920 VPWR.n918 6.04494
R11614 VPWR.n916 VPWR.n914 6.04494
R11615 VPWR.n908 VPWR.n906 6.04494
R11616 VPWR.n904 VPWR.n902 6.04494
R11617 VPWR.n900 VPWR.n898 6.04494
R11618 VPWR.n896 VPWR.n894 6.04494
R11619 VPWR.n892 VPWR.n890 6.04494
R11620 VPWR.n888 VPWR.n886 6.04494
R11621 VPWR.n884 VPWR.n882 6.04494
R11622 VPWR.n880 VPWR.n878 6.04494
R11623 VPWR.n876 VPWR.n874 6.04494
R11624 VPWR.n872 VPWR.n870 6.04494
R11625 VPWR.n869 VPWR.n867 6.04494
R11626 VPWR.n912 VPWR.n910 6.04494
R11627 VPWR.n1870 VPWR.n940 6.04494
R11628 VPWR.n981 VPWR.n979 6.04494
R11629 VPWR.n1494 VPWR.n1227 6.04494
R11630 VPWR.n1221 VPWR.n1179 6.04494
R11631 VPWR.n401 VPWR.n399 6.04494
R11632 VPWR.n2465 VPWR.n361 6.04494
R11633 VPWR.n340 VPWR.n338 6.04494
R11634 VPWR.n2520 VPWR.n92 6.04494
R11635 VPWR.n977 VPWR.n975 6.04494
R11636 VPWR.n1491 VPWR.n1485 6.04494
R11637 VPWR.n1184 VPWR.n1183 6.04494
R11638 VPWR.n1867 VPWR.n941 6.04494
R11639 VPWR.n985 VPWR.n983 6.04494
R11640 VPWR.n1505 VPWR.n1173 6.04494
R11641 VPWR.n1218 VPWR.n1217 6.04494
R11642 VPWR.n409 VPWR.n407 6.04494
R11643 VPWR.n417 VPWR.n415 6.04494
R11644 VPWR.n421 VPWR.n419 6.04494
R11645 VPWR.n425 VPWR.n423 6.04494
R11646 VPWR.n429 VPWR.n427 6.04494
R11647 VPWR.n433 VPWR.n431 6.04494
R11648 VPWR.n437 VPWR.n435 6.04494
R11649 VPWR.n441 VPWR.n439 6.04494
R11650 VPWR.n445 VPWR.n443 6.04494
R11651 VPWR.n447 VPWR.n386 6.04494
R11652 VPWR.n413 VPWR.n411 6.04494
R11653 VPWR.n2448 VPWR.n368 6.04494
R11654 VPWR.n328 VPWR.n326 6.04494
R11655 VPWR.n2541 VPWR.n81 6.04494
R11656 VPWR.n989 VPWR.n987 6.04494
R11657 VPWR.n1508 VPWR.n1169 6.04494
R11658 VPWR.n1215 VPWR.n1214 6.04494
R11659 VPWR.n1860 VPWR.n944 6.04494
R11660 VPWR.n1850 VPWR.n948 6.04494
R11661 VPWR.n1847 VPWR.n949 6.04494
R11662 VPWR.n1840 VPWR.n952 6.04494
R11663 VPWR.n1837 VPWR.n953 6.04494
R11664 VPWR.n1830 VPWR.n956 6.04494
R11665 VPWR.n1827 VPWR.n957 6.04494
R11666 VPWR.n1820 VPWR.n960 6.04494
R11667 VPWR.n1818 VPWR.n961 6.04494
R11668 VPWR.n1857 VPWR.n945 6.04494
R11669 VPWR.n993 VPWR.n991 6.04494
R11670 VPWR.n1519 VPWR.n1163 6.04494
R11671 VPWR.n1212 VPWR.n1206 6.04494
R11672 VPWR.n2468 VPWR.n360 6.04494
R11673 VPWR.n344 VPWR.n342 6.04494
R11674 VPWR.n2517 VPWR.n93 6.04494
R11675 VPWR.n1480 VPWR.n1479 6.04494
R11676 VPWR.n1181 VPWR.n1180 6.04494
R11677 VPWR.n997 VPWR.n995 6.04494
R11678 VPWR.n1522 VPWR.n1159 6.04494
R11679 VPWR.n1204 VPWR.n1203 6.04494
R11680 VPWR.n2438 VPWR.n372 6.04494
R11681 VPWR.n2428 VPWR.n376 6.04494
R11682 VPWR.n2425 VPWR.n377 6.04494
R11683 VPWR.n2418 VPWR.n380 6.04494
R11684 VPWR.n2415 VPWR.n381 6.04494
R11685 VPWR.n2408 VPWR.n384 6.04494
R11686 VPWR.n2406 VPWR.n385 6.04494
R11687 VPWR.n2435 VPWR.n373 6.04494
R11688 VPWR.n316 VPWR.n314 6.04494
R11689 VPWR.n2556 VPWR.n74 6.04494
R11690 VPWR.n1537 VPWR.n1149 6.04494
R11691 VPWR.n1201 VPWR.n1200 6.04494
R11692 VPWR.n1001 VPWR.n999 6.04494
R11693 VPWR.n1005 VPWR.n1003 6.04494
R11694 VPWR.n1009 VPWR.n1007 6.04494
R11695 VPWR.n1013 VPWR.n1011 6.04494
R11696 VPWR.n1017 VPWR.n1015 6.04494
R11697 VPWR.n1021 VPWR.n1019 6.04494
R11698 VPWR.n1023 VPWR.n962 6.04494
R11699 VPWR.n969 VPWR.n967 6.04494
R11700 VPWR.n1474 VPWR.n1472 6.04494
R11701 VPWR.n1592 VPWR.n1123 6.04494
R11702 VPWR.n312 VPWR.n310 6.04494
R11703 VPWR.n2565 VPWR.n69 6.04494
R11704 VPWR.n1198 VPWR.n1192 6.04494
R11705 VPWR.n1762 VPWR.n1049 6.04494
R11706 VPWR.n1190 VPWR.n1189 6.04494
R11707 VPWR.n308 VPWR.n306 6.04494
R11708 VPWR.n304 VPWR.n302 6.04494
R11709 VPWR.n296 VPWR.n294 6.04494
R11710 VPWR.n293 VPWR.n291 6.04494
R11711 VPWR.n300 VPWR.n298 6.04494
R11712 VPWR.n1741 VPWR.n1058 6.04494
R11713 VPWR.n1750 VPWR.n1748 6.04494
R11714 VPWR.n1790 VPWR.n1036 6.04494
R11715 VPWR.n1792 VPWR.n1032 6.04494
R11716 VPWR.n1759 VPWR.n1053 6.04494
R11717 VPWR.n1187 VPWR.n1186 6.04494
R11718 VPWR.n2577 VPWR.n63 6.04494
R11719 VPWR.n2580 VPWR.n62 6.04494
R11720 VPWR.n2589 VPWR.n57 6.04494
R11721 VPWR.n2591 VPWR.n56 6.04494
R11722 VPWR.n1738 VPWR.n1059 6.04494
R11723 VPWR.n1062 VPWR.n1061 6.04494
R11724 VPWR.n2785 VPWR.n2784 5.39628
R11725 VPWR.n2765 VPWR.n2764 5.39628
R11726 VPWR.n2746 VPWR.n2745 5.39628
R11727 VPWR.n54 VPWR 4.72593
R11728 VPWR.n52 VPWR 4.72593
R11729 VPWR.n50 VPWR 4.72593
R11730 VPWR.n48 VPWR 4.72593
R11731 VPWR.n46 VPWR 4.72593
R11732 VPWR.n44 VPWR 4.72593
R11733 VPWR.n42 VPWR 4.72593
R11734 VPWR.n40 VPWR 4.72593
R11735 VPWR.n38 VPWR 4.72593
R11736 VPWR.n36 VPWR 4.72593
R11737 VPWR.n34 VPWR 4.72593
R11738 VPWR.n32 VPWR 4.72593
R11739 VPWR.n30 VPWR 4.72593
R11740 VPWR.n28 VPWR 4.72593
R11741 VPWR.n26 VPWR 4.72593
R11742 VPWR.n1446 VPWR.n1445 4.55954
R11743 VPWR.n2571 VPWR.n2570 4.5005
R11744 VPWR.n2511 VPWR.n2510 4.5005
R11745 VPWR.n2551 VPWR.n2550 4.5005
R11746 VPWR.n319 VPWR.n77 4.5005
R11747 VPWR.n2547 VPWR.n2546 4.5005
R11748 VPWR.n323 VPWR.n78 4.5005
R11749 VPWR.n2535 VPWR.n2534 4.5005
R11750 VPWR.n331 VPWR.n84 4.5005
R11751 VPWR.n2454 VPWR.n2453 4.5005
R11752 VPWR.n2527 VPWR.n2526 4.5005
R11753 VPWR.n335 VPWR.n89 4.5005
R11754 VPWR.n2460 VPWR.n2459 4.5005
R11755 VPWR.n1498 VPWR.n1223 4.5005
R11756 VPWR.n1497 VPWR.n1495 4.5005
R11757 VPWR.n980 VPWR.n939 4.5005
R11758 VPWR.n1872 VPWR.n1871 4.5005
R11759 VPWR.n911 VPWR.n858 4.5005
R11760 VPWR.n1935 VPWR.n1934 4.5005
R11761 VPWR.n788 VPWR.n747 4.5005
R11762 VPWR.n2068 VPWR.n2067 4.5005
R11763 VPWR.n719 VPWR.n666 4.5005
R11764 VPWR.n2131 VPWR.n2130 4.5005
R11765 VPWR.n596 VPWR.n555 4.5005
R11766 VPWR.n2264 VPWR.n2263 4.5005
R11767 VPWR.n527 VPWR.n474 4.5005
R11768 VPWR.n2327 VPWR.n2326 4.5005
R11769 VPWR.n404 VPWR.n363 4.5005
R11770 VPWR.n2523 VPWR.n2522 4.5005
R11771 VPWR.n339 VPWR.n90 4.5005
R11772 VPWR.n2464 VPWR.n2463 4.5005
R11773 VPWR.n400 VPWR.n362 4.5005
R11774 VPWR.n2323 VPWR.n2322 4.5005
R11775 VPWR.n531 VPWR.n475 4.5005
R11776 VPWR.n2268 VPWR.n2267 4.5005
R11777 VPWR.n592 VPWR.n554 4.5005
R11778 VPWR.n2127 VPWR.n2126 4.5005
R11779 VPWR.n723 VPWR.n667 4.5005
R11780 VPWR.n2072 VPWR.n2071 4.5005
R11781 VPWR.n784 VPWR.n746 4.5005
R11782 VPWR.n1931 VPWR.n1930 4.5005
R11783 VPWR.n915 VPWR.n859 4.5005
R11784 VPWR.n1488 VPWR.n1486 4.5005
R11785 VPWR.n1490 VPWR.n1489 4.5005
R11786 VPWR.n976 VPWR.n938 4.5005
R11787 VPWR.n1876 VPWR.n1875 4.5005
R11788 VPWR.n1501 VPWR.n1174 4.5005
R11789 VPWR.n1504 VPWR.n1503 4.5005
R11790 VPWR.n984 VPWR.n942 4.5005
R11791 VPWR.n1866 VPWR.n1865 4.5005
R11792 VPWR.n907 VPWR.n855 4.5005
R11793 VPWR.n1941 VPWR.n1940 4.5005
R11794 VPWR.n792 VPWR.n750 4.5005
R11795 VPWR.n2062 VPWR.n2061 4.5005
R11796 VPWR.n715 VPWR.n663 4.5005
R11797 VPWR.n2137 VPWR.n2136 4.5005
R11798 VPWR.n600 VPWR.n558 4.5005
R11799 VPWR.n2258 VPWR.n2257 4.5005
R11800 VPWR.n523 VPWR.n471 4.5005
R11801 VPWR.n2333 VPWR.n2332 4.5005
R11802 VPWR.n408 VPWR.n366 4.5005
R11803 VPWR.n2539 VPWR.n2538 4.5005
R11804 VPWR.n327 VPWR.n83 4.5005
R11805 VPWR.n2450 VPWR.n2449 4.5005
R11806 VPWR.n412 VPWR.n367 4.5005
R11807 VPWR.n2337 VPWR.n2336 4.5005
R11808 VPWR.n519 VPWR.n470 4.5005
R11809 VPWR.n2254 VPWR.n2253 4.5005
R11810 VPWR.n604 VPWR.n559 4.5005
R11811 VPWR.n2141 VPWR.n2140 4.5005
R11812 VPWR.n711 VPWR.n662 4.5005
R11813 VPWR.n2058 VPWR.n2057 4.5005
R11814 VPWR.n796 VPWR.n751 4.5005
R11815 VPWR.n1945 VPWR.n1944 4.5005
R11816 VPWR.n903 VPWR.n854 4.5005
R11817 VPWR.n1512 VPWR.n1165 4.5005
R11818 VPWR.n1511 VPWR.n1509 4.5005
R11819 VPWR.n988 VPWR.n943 4.5005
R11820 VPWR.n1862 VPWR.n1861 4.5005
R11821 VPWR.n1515 VPWR.n1164 4.5005
R11822 VPWR.n1518 VPWR.n1517 4.5005
R11823 VPWR.n992 VPWR.n946 4.5005
R11824 VPWR.n1856 VPWR.n1855 4.5005
R11825 VPWR.n899 VPWR.n851 4.5005
R11826 VPWR.n1951 VPWR.n1950 4.5005
R11827 VPWR.n800 VPWR.n754 4.5005
R11828 VPWR.n2052 VPWR.n2051 4.5005
R11829 VPWR.n707 VPWR.n659 4.5005
R11830 VPWR.n2147 VPWR.n2146 4.5005
R11831 VPWR.n608 VPWR.n562 4.5005
R11832 VPWR.n2248 VPWR.n2247 4.5005
R11833 VPWR.n515 VPWR.n467 4.5005
R11834 VPWR.n2343 VPWR.n2342 4.5005
R11835 VPWR.n416 VPWR.n370 4.5005
R11836 VPWR.n2444 VPWR.n2443 4.5005
R11837 VPWR.n2515 VPWR.n2514 4.5005
R11838 VPWR.n343 VPWR.n95 4.5005
R11839 VPWR.n2470 VPWR.n2469 4.5005
R11840 VPWR.n396 VPWR.n359 4.5005
R11841 VPWR.n2317 VPWR.n2316 4.5005
R11842 VPWR.n535 VPWR.n478 4.5005
R11843 VPWR.n2274 VPWR.n2273 4.5005
R11844 VPWR.n588 VPWR.n551 4.5005
R11845 VPWR.n2121 VPWR.n2120 4.5005
R11846 VPWR.n727 VPWR.n670 4.5005
R11847 VPWR.n2078 VPWR.n2077 4.5005
R11848 VPWR.n780 VPWR.n743 4.5005
R11849 VPWR.n1925 VPWR.n1924 4.5005
R11850 VPWR.n919 VPWR.n862 4.5005
R11851 VPWR.n1882 VPWR.n1881 4.5005
R11852 VPWR.n1586 VPWR.n1129 4.5005
R11853 VPWR.n1585 VPWR.n1130 4.5005
R11854 VPWR.n972 VPWR.n935 4.5005
R11855 VPWR.n1526 VPWR.n1155 4.5005
R11856 VPWR.n1525 VPWR.n1523 4.5005
R11857 VPWR.n996 VPWR.n947 4.5005
R11858 VPWR.n1852 VPWR.n1851 4.5005
R11859 VPWR.n895 VPWR.n850 4.5005
R11860 VPWR.n1955 VPWR.n1954 4.5005
R11861 VPWR.n804 VPWR.n755 4.5005
R11862 VPWR.n2048 VPWR.n2047 4.5005
R11863 VPWR.n703 VPWR.n658 4.5005
R11864 VPWR.n2151 VPWR.n2150 4.5005
R11865 VPWR.n612 VPWR.n563 4.5005
R11866 VPWR.n2244 VPWR.n2243 4.5005
R11867 VPWR.n511 VPWR.n466 4.5005
R11868 VPWR.n2347 VPWR.n2346 4.5005
R11869 VPWR.n420 VPWR.n371 4.5005
R11870 VPWR.n2440 VPWR.n2439 4.5005
R11871 VPWR.n2559 VPWR.n2558 4.5005
R11872 VPWR.n315 VPWR.n72 4.5005
R11873 VPWR.n2434 VPWR.n2433 4.5005
R11874 VPWR.n424 VPWR.n374 4.5005
R11875 VPWR.n2353 VPWR.n2352 4.5005
R11876 VPWR.n507 VPWR.n463 4.5005
R11877 VPWR.n2238 VPWR.n2237 4.5005
R11878 VPWR.n616 VPWR.n566 4.5005
R11879 VPWR.n2157 VPWR.n2156 4.5005
R11880 VPWR.n699 VPWR.n655 4.5005
R11881 VPWR.n2042 VPWR.n2041 4.5005
R11882 VPWR.n808 VPWR.n758 4.5005
R11883 VPWR.n1961 VPWR.n1960 4.5005
R11884 VPWR.n891 VPWR.n847 4.5005
R11885 VPWR.n1846 VPWR.n1845 4.5005
R11886 VPWR.n1145 VPWR.n1144 4.5005
R11887 VPWR.n1539 VPWR.n1538 4.5005
R11888 VPWR.n1000 VPWR.n950 4.5005
R11889 VPWR.n1590 VPWR.n1589 4.5005
R11890 VPWR.n1473 VPWR.n1128 4.5005
R11891 VPWR.n968 VPWR.n934 4.5005
R11892 VPWR.n1886 VPWR.n1885 4.5005
R11893 VPWR.n923 VPWR.n863 4.5005
R11894 VPWR.n1921 VPWR.n1920 4.5005
R11895 VPWR.n776 VPWR.n742 4.5005
R11896 VPWR.n2082 VPWR.n2081 4.5005
R11897 VPWR.n731 VPWR.n671 4.5005
R11898 VPWR.n2117 VPWR.n2116 4.5005
R11899 VPWR.n584 VPWR.n550 4.5005
R11900 VPWR.n2278 VPWR.n2277 4.5005
R11901 VPWR.n539 VPWR.n479 4.5005
R11902 VPWR.n2313 VPWR.n2312 4.5005
R11903 VPWR.n392 VPWR.n358 4.5005
R11904 VPWR.n2474 VPWR.n2473 4.5005
R11905 VPWR.n347 VPWR.n96 4.5005
R11906 VPWR.n2563 VPWR.n2562 4.5005
R11907 VPWR.n311 VPWR.n71 4.5005
R11908 VPWR.n2430 VPWR.n2429 4.5005
R11909 VPWR.n428 VPWR.n375 4.5005
R11910 VPWR.n2357 VPWR.n2356 4.5005
R11911 VPWR.n503 VPWR.n462 4.5005
R11912 VPWR.n2234 VPWR.n2233 4.5005
R11913 VPWR.n620 VPWR.n567 4.5005
R11914 VPWR.n2161 VPWR.n2160 4.5005
R11915 VPWR.n695 VPWR.n654 4.5005
R11916 VPWR.n2038 VPWR.n2037 4.5005
R11917 VPWR.n812 VPWR.n759 4.5005
R11918 VPWR.n1965 VPWR.n1964 4.5005
R11919 VPWR.n887 VPWR.n846 4.5005
R11920 VPWR.n1842 VPWR.n1841 4.5005
R11921 VPWR.n1004 VPWR.n951 4.5005
R11922 VPWR.n1531 VPWR.n1154 4.5005
R11923 VPWR.n1533 VPWR.n1532 4.5005
R11924 VPWR.n1073 VPWR.n1045 4.5005
R11925 VPWR.n1764 VPWR.n1763 4.5005
R11926 VPWR.n1008 VPWR.n954 4.5005
R11927 VPWR.n1836 VPWR.n1835 4.5005
R11928 VPWR.n883 VPWR.n843 4.5005
R11929 VPWR.n1971 VPWR.n1970 4.5005
R11930 VPWR.n816 VPWR.n762 4.5005
R11931 VPWR.n2032 VPWR.n2031 4.5005
R11932 VPWR.n691 VPWR.n651 4.5005
R11933 VPWR.n2167 VPWR.n2166 4.5005
R11934 VPWR.n624 VPWR.n570 4.5005
R11935 VPWR.n2228 VPWR.n2227 4.5005
R11936 VPWR.n499 VPWR.n459 4.5005
R11937 VPWR.n2363 VPWR.n2362 4.5005
R11938 VPWR.n432 VPWR.n378 4.5005
R11939 VPWR.n2424 VPWR.n2423 4.5005
R11940 VPWR.n307 VPWR.n66 4.5005
R11941 VPWR.n299 VPWR.n60 4.5005
R11942 VPWR.n2414 VPWR.n2413 4.5005
R11943 VPWR.n440 VPWR.n382 4.5005
R11944 VPWR.n2373 VPWR.n2372 4.5005
R11945 VPWR.n491 VPWR.n455 4.5005
R11946 VPWR.n2218 VPWR.n2217 4.5005
R11947 VPWR.n632 VPWR.n574 4.5005
R11948 VPWR.n2177 VPWR.n2176 4.5005
R11949 VPWR.n683 VPWR.n647 4.5005
R11950 VPWR.n2022 VPWR.n2021 4.5005
R11951 VPWR.n824 VPWR.n766 4.5005
R11952 VPWR.n1981 VPWR.n1980 4.5005
R11953 VPWR.n875 VPWR.n839 4.5005
R11954 VPWR.n1826 VPWR.n1825 4.5005
R11955 VPWR.n1016 VPWR.n958 4.5005
R11956 VPWR.n1753 VPWR.n1743 4.5005
R11957 VPWR.n1752 VPWR.n1751 4.5005
R11958 VPWR.n1756 VPWR.n1054 4.5005
R11959 VPWR.n1758 VPWR.n1757 4.5005
R11960 VPWR.n1012 VPWR.n955 4.5005
R11961 VPWR.n1832 VPWR.n1831 4.5005
R11962 VPWR.n879 VPWR.n842 4.5005
R11963 VPWR.n1975 VPWR.n1974 4.5005
R11964 VPWR.n820 VPWR.n763 4.5005
R11965 VPWR.n2028 VPWR.n2027 4.5005
R11966 VPWR.n687 VPWR.n650 4.5005
R11967 VPWR.n2171 VPWR.n2170 4.5005
R11968 VPWR.n628 VPWR.n571 4.5005
R11969 VPWR.n2224 VPWR.n2223 4.5005
R11970 VPWR.n495 VPWR.n458 4.5005
R11971 VPWR.n2367 VPWR.n2366 4.5005
R11972 VPWR.n436 VPWR.n379 4.5005
R11973 VPWR.n2420 VPWR.n2419 4.5005
R11974 VPWR.n303 VPWR.n65 4.5005
R11975 VPWR.n2575 VPWR.n2574 4.5005
R11976 VPWR.n2583 VPWR.n2582 4.5005
R11977 VPWR.n2587 VPWR.n2586 4.5005
R11978 VPWR.n295 VPWR.n59 4.5005
R11979 VPWR.n2410 VPWR.n2409 4.5005
R11980 VPWR.n444 VPWR.n383 4.5005
R11981 VPWR.n2377 VPWR.n2376 4.5005
R11982 VPWR.n487 VPWR.n454 4.5005
R11983 VPWR.n2214 VPWR.n2213 4.5005
R11984 VPWR.n636 VPWR.n575 4.5005
R11985 VPWR.n2181 VPWR.n2180 4.5005
R11986 VPWR.n679 VPWR.n646 4.5005
R11987 VPWR.n2018 VPWR.n2017 4.5005
R11988 VPWR.n828 VPWR.n767 4.5005
R11989 VPWR.n1985 VPWR.n1984 4.5005
R11990 VPWR.n871 VPWR.n838 4.5005
R11991 VPWR.n1822 VPWR.n1821 4.5005
R11992 VPWR.n1020 VPWR.n959 4.5005
R11993 VPWR.n1789 VPWR.n1788 4.5005
R11994 VPWR.n1736 VPWR.n1037 4.5005
R11995 VPWR.n1232 VPWR.n1121 4.5005
R11996 VPWR.n1466 VPWR.n1465 4.5005
R11997 VPWR.n964 VPWR.n931 4.5005
R11998 VPWR.n1892 VPWR.n1891 4.5005
R11999 VPWR.n929 VPWR.n928 4.5005
R12000 VPWR.n1915 VPWR.n1914 4.5005
R12001 VPWR.n772 VPWR.n739 4.5005
R12002 VPWR.n2088 VPWR.n2087 4.5005
R12003 VPWR.n737 VPWR.n736 4.5005
R12004 VPWR.n2111 VPWR.n2110 4.5005
R12005 VPWR.n580 VPWR.n547 4.5005
R12006 VPWR.n2284 VPWR.n2283 4.5005
R12007 VPWR.n545 VPWR.n544 4.5005
R12008 VPWR.n2307 VPWR.n2306 4.5005
R12009 VPWR.n388 VPWR.n355 4.5005
R12010 VPWR.n2480 VPWR.n2479 4.5005
R12011 VPWR.n353 VPWR.n352 4.5005
R12012 VPWR.n2503 VPWR.n2502 4.5005
R12013 VPWR.n2594 VPWR.n2593 4.5005
R12014 VPWR.n292 VPWR.n22 4.5005
R12015 VPWR.n2405 VPWR.n2404 4.5005
R12016 VPWR.n449 VPWR.n448 4.5005
R12017 VPWR.n2382 VPWR.n2381 4.5005
R12018 VPWR.n484 VPWR.n451 4.5005
R12019 VPWR.n2209 VPWR.n2208 4.5005
R12020 VPWR.n641 VPWR.n640 4.5005
R12021 VPWR.n2186 VPWR.n2185 4.5005
R12022 VPWR.n676 VPWR.n643 4.5005
R12023 VPWR.n2013 VPWR.n2012 4.5005
R12024 VPWR.n833 VPWR.n832 4.5005
R12025 VPWR.n1990 VPWR.n1989 4.5005
R12026 VPWR.n868 VPWR.n835 4.5005
R12027 VPWR.n1817 VPWR.n1816 4.5005
R12028 VPWR.n1025 VPWR.n1024 4.5005
R12029 VPWR.n1794 VPWR.n1793 4.5005
R12030 VPWR.n1060 VPWR.n1028 4.5005
R12031 VPWR.n2628 VPWR 4.49965
R12032 VPWR.n19 VPWR.n18 4.20017
R12033 VPWR.n1255 VPWR.n1254 4.20017
R12034 VPWR.n1279 VPWR.n1278 4.20017
R12035 VPWR.n1302 VPWR.n1301 4.20017
R12036 VPWR.n1337 VPWR.n1336 4.20017
R12037 VPWR.n1376 VPWR.n1375 4.20017
R12038 VPWR.n1414 VPWR.n1413 4.20017
R12039 VPWR.n2813 VPWR 4.14027
R12040 VPWR.n2797 VPWR 4.14027
R12041 VPWR.n2778 VPWR 4.14027
R12042 VPWR.n2758 VPWR 4.14027
R12043 VPWR.n2739 VPWR 4.14027
R12044 VPWR.n2703 VPWR 4.14027
R12045 VPWR.n2665 VPWR 4.14027
R12046 VPWR.n55 VPWR.n54 4.0005
R12047 VPWR.n2716 VPWR.n2713 3.76521
R12048 VPWR.n2680 VPWR.n2676 3.76521
R12049 VPWR.n2643 VPWR.n2639 3.76521
R12050 VPWR.n2611 VPWR.n2610 3.76521
R12051 VPWR.n1906 VPWR.n858 3.4105
R12052 VPWR.n1934 VPWR.n1933 3.4105
R12053 VPWR.n1997 VPWR.n747 3.4105
R12054 VPWR.n2069 VPWR.n2068 3.4105
R12055 VPWR.n2102 VPWR.n666 3.4105
R12056 VPWR.n2130 VPWR.n2129 3.4105
R12057 VPWR.n2193 VPWR.n555 3.4105
R12058 VPWR.n2265 VPWR.n2264 3.4105
R12059 VPWR.n2298 VPWR.n474 3.4105
R12060 VPWR.n2326 VPWR.n2325 3.4105
R12061 VPWR.n2389 VPWR.n363 3.4105
R12062 VPWR.n2388 VPWR.n362 3.4105
R12063 VPWR.n2324 VPWR.n2323 3.4105
R12064 VPWR.n2299 VPWR.n475 3.4105
R12065 VPWR.n2267 VPWR.n2266 3.4105
R12066 VPWR.n2192 VPWR.n554 3.4105
R12067 VPWR.n2128 VPWR.n2127 3.4105
R12068 VPWR.n2103 VPWR.n667 3.4105
R12069 VPWR.n2071 VPWR.n2070 3.4105
R12070 VPWR.n1996 VPWR.n746 3.4105
R12071 VPWR.n1932 VPWR.n1931 3.4105
R12072 VPWR.n1907 VPWR.n859 3.4105
R12073 VPWR.n1875 VPWR.n1874 3.4105
R12074 VPWR.n1873 VPWR.n1872 3.4105
R12075 VPWR.n1865 VPWR.n1864 3.4105
R12076 VPWR.n1905 VPWR.n855 3.4105
R12077 VPWR.n1942 VPWR.n1941 3.4105
R12078 VPWR.n1998 VPWR.n750 3.4105
R12079 VPWR.n2061 VPWR.n2060 3.4105
R12080 VPWR.n2101 VPWR.n663 3.4105
R12081 VPWR.n2138 VPWR.n2137 3.4105
R12082 VPWR.n2194 VPWR.n558 3.4105
R12083 VPWR.n2257 VPWR.n2256 3.4105
R12084 VPWR.n2297 VPWR.n471 3.4105
R12085 VPWR.n2334 VPWR.n2333 3.4105
R12086 VPWR.n2390 VPWR.n366 3.4105
R12087 VPWR.n2391 VPWR.n367 3.4105
R12088 VPWR.n2336 VPWR.n2335 3.4105
R12089 VPWR.n2296 VPWR.n470 3.4105
R12090 VPWR.n2255 VPWR.n2254 3.4105
R12091 VPWR.n2195 VPWR.n559 3.4105
R12092 VPWR.n2140 VPWR.n2139 3.4105
R12093 VPWR.n2100 VPWR.n662 3.4105
R12094 VPWR.n2059 VPWR.n2058 3.4105
R12095 VPWR.n1999 VPWR.n751 3.4105
R12096 VPWR.n1944 VPWR.n1943 3.4105
R12097 VPWR.n1904 VPWR.n854 3.4105
R12098 VPWR.n1863 VPWR.n1862 3.4105
R12099 VPWR.n1855 VPWR.n1854 3.4105
R12100 VPWR.n1903 VPWR.n851 3.4105
R12101 VPWR.n1952 VPWR.n1951 3.4105
R12102 VPWR.n2000 VPWR.n754 3.4105
R12103 VPWR.n2051 VPWR.n2050 3.4105
R12104 VPWR.n2099 VPWR.n659 3.4105
R12105 VPWR.n2148 VPWR.n2147 3.4105
R12106 VPWR.n2196 VPWR.n562 3.4105
R12107 VPWR.n2247 VPWR.n2246 3.4105
R12108 VPWR.n2295 VPWR.n467 3.4105
R12109 VPWR.n2344 VPWR.n2343 3.4105
R12110 VPWR.n2392 VPWR.n370 3.4105
R12111 VPWR.n2443 VPWR.n2442 3.4105
R12112 VPWR.n2451 VPWR.n2450 3.4105
R12113 VPWR.n2453 VPWR.n2452 3.4105
R12114 VPWR.n2461 VPWR.n2460 3.4105
R12115 VPWR.n2463 VPWR.n2462 3.4105
R12116 VPWR.n2471 VPWR.n2470 3.4105
R12117 VPWR.n2387 VPWR.n359 3.4105
R12118 VPWR.n2316 VPWR.n2315 3.4105
R12119 VPWR.n2300 VPWR.n478 3.4105
R12120 VPWR.n2275 VPWR.n2274 3.4105
R12121 VPWR.n2191 VPWR.n551 3.4105
R12122 VPWR.n2120 VPWR.n2119 3.4105
R12123 VPWR.n2104 VPWR.n670 3.4105
R12124 VPWR.n2079 VPWR.n2078 3.4105
R12125 VPWR.n1995 VPWR.n743 3.4105
R12126 VPWR.n1924 VPWR.n1923 3.4105
R12127 VPWR.n1908 VPWR.n862 3.4105
R12128 VPWR.n1883 VPWR.n1882 3.4105
R12129 VPWR.n1799 VPWR.n935 3.4105
R12130 VPWR.n1800 VPWR.n938 3.4105
R12131 VPWR.n1801 VPWR.n939 3.4105
R12132 VPWR.n1802 VPWR.n942 3.4105
R12133 VPWR.n1803 VPWR.n943 3.4105
R12134 VPWR.n1804 VPWR.n946 3.4105
R12135 VPWR.n1805 VPWR.n947 3.4105
R12136 VPWR.n1853 VPWR.n1852 3.4105
R12137 VPWR.n1902 VPWR.n850 3.4105
R12138 VPWR.n1954 VPWR.n1953 3.4105
R12139 VPWR.n2001 VPWR.n755 3.4105
R12140 VPWR.n2049 VPWR.n2048 3.4105
R12141 VPWR.n2098 VPWR.n658 3.4105
R12142 VPWR.n2150 VPWR.n2149 3.4105
R12143 VPWR.n2197 VPWR.n563 3.4105
R12144 VPWR.n2245 VPWR.n2244 3.4105
R12145 VPWR.n2294 VPWR.n466 3.4105
R12146 VPWR.n2346 VPWR.n2345 3.4105
R12147 VPWR.n2393 VPWR.n371 3.4105
R12148 VPWR.n2441 VPWR.n2440 3.4105
R12149 VPWR.n2433 VPWR.n2432 3.4105
R12150 VPWR.n2394 VPWR.n374 3.4105
R12151 VPWR.n2354 VPWR.n2353 3.4105
R12152 VPWR.n2293 VPWR.n463 3.4105
R12153 VPWR.n2237 VPWR.n2236 3.4105
R12154 VPWR.n2198 VPWR.n566 3.4105
R12155 VPWR.n2158 VPWR.n2157 3.4105
R12156 VPWR.n2097 VPWR.n655 3.4105
R12157 VPWR.n2041 VPWR.n2040 3.4105
R12158 VPWR.n2002 VPWR.n758 3.4105
R12159 VPWR.n1962 VPWR.n1961 3.4105
R12160 VPWR.n1901 VPWR.n847 3.4105
R12161 VPWR.n1845 VPWR.n1844 3.4105
R12162 VPWR.n1806 VPWR.n950 3.4105
R12163 VPWR.n1798 VPWR.n934 3.4105
R12164 VPWR.n1885 VPWR.n1884 3.4105
R12165 VPWR.n1909 VPWR.n863 3.4105
R12166 VPWR.n1922 VPWR.n1921 3.4105
R12167 VPWR.n1994 VPWR.n742 3.4105
R12168 VPWR.n2081 VPWR.n2080 3.4105
R12169 VPWR.n2105 VPWR.n671 3.4105
R12170 VPWR.n2118 VPWR.n2117 3.4105
R12171 VPWR.n2190 VPWR.n550 3.4105
R12172 VPWR.n2277 VPWR.n2276 3.4105
R12173 VPWR.n2301 VPWR.n479 3.4105
R12174 VPWR.n2314 VPWR.n2313 3.4105
R12175 VPWR.n2386 VPWR.n358 3.4105
R12176 VPWR.n2473 VPWR.n2472 3.4105
R12177 VPWR.n2497 VPWR.n96 3.4105
R12178 VPWR.n2496 VPWR.n95 3.4105
R12179 VPWR.n2495 VPWR.n90 3.4105
R12180 VPWR.n2494 VPWR.n89 3.4105
R12181 VPWR.n2493 VPWR.n84 3.4105
R12182 VPWR.n2492 VPWR.n83 3.4105
R12183 VPWR.n2491 VPWR.n78 3.4105
R12184 VPWR.n2490 VPWR.n77 3.4105
R12185 VPWR.n2489 VPWR.n72 3.4105
R12186 VPWR.n2488 VPWR.n71 3.4105
R12187 VPWR.n2431 VPWR.n2430 3.4105
R12188 VPWR.n2395 VPWR.n375 3.4105
R12189 VPWR.n2356 VPWR.n2355 3.4105
R12190 VPWR.n2292 VPWR.n462 3.4105
R12191 VPWR.n2235 VPWR.n2234 3.4105
R12192 VPWR.n2199 VPWR.n567 3.4105
R12193 VPWR.n2160 VPWR.n2159 3.4105
R12194 VPWR.n2096 VPWR.n654 3.4105
R12195 VPWR.n2039 VPWR.n2038 3.4105
R12196 VPWR.n2003 VPWR.n759 3.4105
R12197 VPWR.n1964 VPWR.n1963 3.4105
R12198 VPWR.n1900 VPWR.n846 3.4105
R12199 VPWR.n1843 VPWR.n1842 3.4105
R12200 VPWR.n1807 VPWR.n951 3.4105
R12201 VPWR.n1532 VPWR.n1143 3.4105
R12202 VPWR.n1540 VPWR.n1539 3.4105
R12203 VPWR.n1525 VPWR.n1524 3.4105
R12204 VPWR.n1517 VPWR.n1516 3.4105
R12205 VPWR.n1511 VPWR.n1510 3.4105
R12206 VPWR.n1503 VPWR.n1502 3.4105
R12207 VPWR.n1497 VPWR.n1496 3.4105
R12208 VPWR.n1489 VPWR.n1132 3.4105
R12209 VPWR.n1585 VPWR.n1584 3.4105
R12210 VPWR.n1452 VPWR.n1128 3.4105
R12211 VPWR.n1765 VPWR.n1764 3.4105
R12212 VPWR.n1808 VPWR.n954 3.4105
R12213 VPWR.n1835 VPWR.n1834 3.4105
R12214 VPWR.n1899 VPWR.n843 3.4105
R12215 VPWR.n1972 VPWR.n1971 3.4105
R12216 VPWR.n2004 VPWR.n762 3.4105
R12217 VPWR.n2031 VPWR.n2030 3.4105
R12218 VPWR.n2095 VPWR.n651 3.4105
R12219 VPWR.n2168 VPWR.n2167 3.4105
R12220 VPWR.n2200 VPWR.n570 3.4105
R12221 VPWR.n2227 VPWR.n2226 3.4105
R12222 VPWR.n2291 VPWR.n459 3.4105
R12223 VPWR.n2364 VPWR.n2363 3.4105
R12224 VPWR.n2396 VPWR.n378 3.4105
R12225 VPWR.n2423 VPWR.n2422 3.4105
R12226 VPWR.n2487 VPWR.n66 3.4105
R12227 VPWR.n2485 VPWR.n60 3.4105
R12228 VPWR.n2413 VPWR.n2412 3.4105
R12229 VPWR.n2398 VPWR.n382 3.4105
R12230 VPWR.n2374 VPWR.n2373 3.4105
R12231 VPWR.n2289 VPWR.n455 3.4105
R12232 VPWR.n2217 VPWR.n2216 3.4105
R12233 VPWR.n2202 VPWR.n574 3.4105
R12234 VPWR.n2178 VPWR.n2177 3.4105
R12235 VPWR.n2093 VPWR.n647 3.4105
R12236 VPWR.n2021 VPWR.n2020 3.4105
R12237 VPWR.n2006 VPWR.n766 3.4105
R12238 VPWR.n1982 VPWR.n1981 3.4105
R12239 VPWR.n1897 VPWR.n839 3.4105
R12240 VPWR.n1825 VPWR.n1824 3.4105
R12241 VPWR.n1810 VPWR.n958 3.4105
R12242 VPWR.n1752 VPWR.n1744 3.4105
R12243 VPWR.n1757 VPWR.n1043 3.4105
R12244 VPWR.n1809 VPWR.n955 3.4105
R12245 VPWR.n1833 VPWR.n1832 3.4105
R12246 VPWR.n1898 VPWR.n842 3.4105
R12247 VPWR.n1974 VPWR.n1973 3.4105
R12248 VPWR.n2005 VPWR.n763 3.4105
R12249 VPWR.n2029 VPWR.n2028 3.4105
R12250 VPWR.n2094 VPWR.n650 3.4105
R12251 VPWR.n2170 VPWR.n2169 3.4105
R12252 VPWR.n2201 VPWR.n571 3.4105
R12253 VPWR.n2225 VPWR.n2224 3.4105
R12254 VPWR.n2290 VPWR.n458 3.4105
R12255 VPWR.n2366 VPWR.n2365 3.4105
R12256 VPWR.n2397 VPWR.n379 3.4105
R12257 VPWR.n2421 VPWR.n2420 3.4105
R12258 VPWR.n2486 VPWR.n65 3.4105
R12259 VPWR.n2484 VPWR.n59 3.4105
R12260 VPWR.n2411 VPWR.n2410 3.4105
R12261 VPWR.n2399 VPWR.n383 3.4105
R12262 VPWR.n2376 VPWR.n2375 3.4105
R12263 VPWR.n2288 VPWR.n454 3.4105
R12264 VPWR.n2215 VPWR.n2214 3.4105
R12265 VPWR.n2203 VPWR.n575 3.4105
R12266 VPWR.n2180 VPWR.n2179 3.4105
R12267 VPWR.n2092 VPWR.n646 3.4105
R12268 VPWR.n2019 VPWR.n2018 3.4105
R12269 VPWR.n2007 VPWR.n767 3.4105
R12270 VPWR.n1984 VPWR.n1983 3.4105
R12271 VPWR.n1896 VPWR.n838 3.4105
R12272 VPWR.n1823 VPWR.n1822 3.4105
R12273 VPWR.n1811 VPWR.n959 3.4105
R12274 VPWR.n1788 VPWR.n1787 3.4105
R12275 VPWR.n1465 VPWR.n1464 3.4105
R12276 VPWR.n1797 VPWR.n931 3.4105
R12277 VPWR.n1893 VPWR.n1892 3.4105
R12278 VPWR.n1910 VPWR.n929 3.4105
R12279 VPWR.n1914 VPWR.n1913 3.4105
R12280 VPWR.n1993 VPWR.n739 3.4105
R12281 VPWR.n2089 VPWR.n2088 3.4105
R12282 VPWR.n2106 VPWR.n737 3.4105
R12283 VPWR.n2110 VPWR.n2109 3.4105
R12284 VPWR.n2189 VPWR.n547 3.4105
R12285 VPWR.n2285 VPWR.n2284 3.4105
R12286 VPWR.n2302 VPWR.n545 3.4105
R12287 VPWR.n2306 VPWR.n2305 3.4105
R12288 VPWR.n2385 VPWR.n355 3.4105
R12289 VPWR.n2481 VPWR.n2480 3.4105
R12290 VPWR.n2498 VPWR.n353 3.4105
R12291 VPWR.n2502 VPWR.n2501 3.4105
R12292 VPWR.n2512 VPWR.n2511 3.4105
R12293 VPWR.n2514 VPWR.n2513 3.4105
R12294 VPWR.n2524 VPWR.n2523 3.4105
R12295 VPWR.n2526 VPWR.n2525 3.4105
R12296 VPWR.n2536 VPWR.n2535 3.4105
R12297 VPWR.n2538 VPWR.n2537 3.4105
R12298 VPWR.n2548 VPWR.n2547 3.4105
R12299 VPWR.n2550 VPWR.n2549 3.4105
R12300 VPWR.n2560 VPWR.n2559 3.4105
R12301 VPWR.n2562 VPWR.n2561 3.4105
R12302 VPWR.n2572 VPWR.n2571 3.4105
R12303 VPWR.n2574 VPWR.n2573 3.4105
R12304 VPWR.n2584 VPWR.n2583 3.4105
R12305 VPWR.n2586 VPWR.n2585 3.4105
R12306 VPWR.n2595 VPWR.n2594 3.4105
R12307 VPWR.n2483 VPWR.n22 3.4105
R12308 VPWR.n2404 VPWR.n2403 3.4105
R12309 VPWR.n2400 VPWR.n449 3.4105
R12310 VPWR.n2383 VPWR.n2382 3.4105
R12311 VPWR.n2287 VPWR.n451 3.4105
R12312 VPWR.n2208 VPWR.n2207 3.4105
R12313 VPWR.n2204 VPWR.n641 3.4105
R12314 VPWR.n2187 VPWR.n2186 3.4105
R12315 VPWR.n2091 VPWR.n643 3.4105
R12316 VPWR.n2012 VPWR.n2011 3.4105
R12317 VPWR.n2008 VPWR.n833 3.4105
R12318 VPWR.n1991 VPWR.n1990 3.4105
R12319 VPWR.n1895 VPWR.n835 3.4105
R12320 VPWR.n1816 VPWR.n1815 3.4105
R12321 VPWR.n1812 VPWR.n1025 3.4105
R12322 VPWR.n1795 VPWR.n1794 3.4105
R12323 VPWR.n1055 VPWR.n1028 3.4105
R12324 VPWR.n1056 VPWR.n1037 3.4105
R12325 VPWR.n1754 VPWR.n1753 3.4105
R12326 VPWR.n1756 VPWR.n1755 3.4105
R12327 VPWR.n1529 VPWR.n1045 3.4105
R12328 VPWR.n1531 VPWR.n1530 3.4105
R12329 VPWR.n1528 VPWR.n1145 3.4105
R12330 VPWR.n1527 VPWR.n1526 3.4105
R12331 VPWR.n1515 VPWR.n1514 3.4105
R12332 VPWR.n1513 VPWR.n1512 3.4105
R12333 VPWR.n1501 VPWR.n1500 3.4105
R12334 VPWR.n1499 VPWR.n1498 3.4105
R12335 VPWR.n1488 VPWR.n1487 3.4105
R12336 VPWR.n1587 VPWR.n1586 3.4105
R12337 VPWR.n1589 VPWR.n1588 3.4105
R12338 VPWR.n1448 VPWR.n1232 3.4105
R12339 VPWR.n1345 VPWR.n1341 3.38874
R12340 VPWR.n1384 VPWR.n1380 3.38874
R12341 VPWR.n1421 VPWR.n1417 3.38874
R12342 VPWR.n28 VPWR.n26 3.36211
R12343 VPWR.n30 VPWR.n28 3.36211
R12344 VPWR.n32 VPWR.n30 3.36211
R12345 VPWR.n34 VPWR.n32 3.36211
R12346 VPWR.n36 VPWR.n34 3.36211
R12347 VPWR.n38 VPWR.n36 3.36211
R12348 VPWR.n40 VPWR.n38 3.36211
R12349 VPWR.n42 VPWR.n40 3.36211
R12350 VPWR.n44 VPWR.n42 3.36211
R12351 VPWR.n46 VPWR.n44 3.36211
R12352 VPWR.n48 VPWR.n46 3.36211
R12353 VPWR.n50 VPWR.n48 3.36211
R12354 VPWR.n52 VPWR.n50 3.36211
R12355 VPWR.n54 VPWR.n52 3.36211
R12356 VPWR.t976 VPWR.t524 3.35739
R12357 VPWR.t1891 VPWR.t1407 3.35739
R12358 VPWR.n2571 VPWR.n66 3.28012
R12359 VPWR.n2511 VPWR.n96 3.28012
R12360 VPWR.n2550 VPWR.n77 3.28012
R12361 VPWR.n2440 VPWR.n77 3.28012
R12362 VPWR.n2547 VPWR.n78 3.28012
R12363 VPWR.n2443 VPWR.n78 3.28012
R12364 VPWR.n2535 VPWR.n84 3.28012
R12365 VPWR.n2453 VPWR.n84 3.28012
R12366 VPWR.n2453 VPWR.n366 3.28012
R12367 VPWR.n2526 VPWR.n89 3.28012
R12368 VPWR.n2460 VPWR.n89 3.28012
R12369 VPWR.n2460 VPWR.n363 3.28012
R12370 VPWR.n1498 VPWR.n1497 3.28012
R12371 VPWR.n1497 VPWR.n939 3.28012
R12372 VPWR.n1872 VPWR.n939 3.28012
R12373 VPWR.n1872 VPWR.n858 3.28012
R12374 VPWR.n1934 VPWR.n858 3.28012
R12375 VPWR.n1934 VPWR.n747 3.28012
R12376 VPWR.n2068 VPWR.n747 3.28012
R12377 VPWR.n2068 VPWR.n666 3.28012
R12378 VPWR.n2130 VPWR.n666 3.28012
R12379 VPWR.n2130 VPWR.n555 3.28012
R12380 VPWR.n2264 VPWR.n555 3.28012
R12381 VPWR.n2264 VPWR.n474 3.28012
R12382 VPWR.n2326 VPWR.n474 3.28012
R12383 VPWR.n2326 VPWR.n363 3.28012
R12384 VPWR.n2523 VPWR.n90 3.28012
R12385 VPWR.n2463 VPWR.n90 3.28012
R12386 VPWR.n2463 VPWR.n362 3.28012
R12387 VPWR.n2323 VPWR.n362 3.28012
R12388 VPWR.n2323 VPWR.n475 3.28012
R12389 VPWR.n2267 VPWR.n475 3.28012
R12390 VPWR.n2267 VPWR.n554 3.28012
R12391 VPWR.n2127 VPWR.n554 3.28012
R12392 VPWR.n2127 VPWR.n667 3.28012
R12393 VPWR.n2071 VPWR.n667 3.28012
R12394 VPWR.n2071 VPWR.n746 3.28012
R12395 VPWR.n1931 VPWR.n746 3.28012
R12396 VPWR.n1931 VPWR.n859 3.28012
R12397 VPWR.n1875 VPWR.n859 3.28012
R12398 VPWR.n1489 VPWR.n1488 3.28012
R12399 VPWR.n1489 VPWR.n938 3.28012
R12400 VPWR.n1875 VPWR.n938 3.28012
R12401 VPWR.n1503 VPWR.n1501 3.28012
R12402 VPWR.n1503 VPWR.n942 3.28012
R12403 VPWR.n1865 VPWR.n942 3.28012
R12404 VPWR.n1865 VPWR.n855 3.28012
R12405 VPWR.n1941 VPWR.n855 3.28012
R12406 VPWR.n1941 VPWR.n750 3.28012
R12407 VPWR.n2061 VPWR.n750 3.28012
R12408 VPWR.n2061 VPWR.n663 3.28012
R12409 VPWR.n2137 VPWR.n663 3.28012
R12410 VPWR.n2137 VPWR.n558 3.28012
R12411 VPWR.n2257 VPWR.n558 3.28012
R12412 VPWR.n2257 VPWR.n471 3.28012
R12413 VPWR.n2333 VPWR.n471 3.28012
R12414 VPWR.n2333 VPWR.n366 3.28012
R12415 VPWR.n2538 VPWR.n83 3.28012
R12416 VPWR.n2450 VPWR.n83 3.28012
R12417 VPWR.n2450 VPWR.n367 3.28012
R12418 VPWR.n2336 VPWR.n367 3.28012
R12419 VPWR.n2336 VPWR.n470 3.28012
R12420 VPWR.n2254 VPWR.n470 3.28012
R12421 VPWR.n2254 VPWR.n559 3.28012
R12422 VPWR.n2140 VPWR.n559 3.28012
R12423 VPWR.n2140 VPWR.n662 3.28012
R12424 VPWR.n2058 VPWR.n662 3.28012
R12425 VPWR.n2058 VPWR.n751 3.28012
R12426 VPWR.n1944 VPWR.n751 3.28012
R12427 VPWR.n1944 VPWR.n854 3.28012
R12428 VPWR.n1862 VPWR.n854 3.28012
R12429 VPWR.n1512 VPWR.n1511 3.28012
R12430 VPWR.n1511 VPWR.n943 3.28012
R12431 VPWR.n1862 VPWR.n943 3.28012
R12432 VPWR.n1517 VPWR.n1515 3.28012
R12433 VPWR.n1517 VPWR.n946 3.28012
R12434 VPWR.n1855 VPWR.n946 3.28012
R12435 VPWR.n1855 VPWR.n851 3.28012
R12436 VPWR.n1951 VPWR.n851 3.28012
R12437 VPWR.n1951 VPWR.n754 3.28012
R12438 VPWR.n2051 VPWR.n754 3.28012
R12439 VPWR.n2051 VPWR.n659 3.28012
R12440 VPWR.n2147 VPWR.n659 3.28012
R12441 VPWR.n2147 VPWR.n562 3.28012
R12442 VPWR.n2247 VPWR.n562 3.28012
R12443 VPWR.n2247 VPWR.n467 3.28012
R12444 VPWR.n2343 VPWR.n467 3.28012
R12445 VPWR.n2343 VPWR.n370 3.28012
R12446 VPWR.n2443 VPWR.n370 3.28012
R12447 VPWR.n2514 VPWR.n95 3.28012
R12448 VPWR.n2470 VPWR.n95 3.28012
R12449 VPWR.n2470 VPWR.n359 3.28012
R12450 VPWR.n2316 VPWR.n359 3.28012
R12451 VPWR.n2316 VPWR.n478 3.28012
R12452 VPWR.n2274 VPWR.n478 3.28012
R12453 VPWR.n2274 VPWR.n551 3.28012
R12454 VPWR.n2120 VPWR.n551 3.28012
R12455 VPWR.n2120 VPWR.n670 3.28012
R12456 VPWR.n2078 VPWR.n670 3.28012
R12457 VPWR.n2078 VPWR.n743 3.28012
R12458 VPWR.n1924 VPWR.n743 3.28012
R12459 VPWR.n1924 VPWR.n862 3.28012
R12460 VPWR.n1882 VPWR.n862 3.28012
R12461 VPWR.n1882 VPWR.n935 3.28012
R12462 VPWR.n1586 VPWR.n1585 3.28012
R12463 VPWR.n1585 VPWR.n935 3.28012
R12464 VPWR.n1526 VPWR.n1525 3.28012
R12465 VPWR.n1525 VPWR.n947 3.28012
R12466 VPWR.n1852 VPWR.n947 3.28012
R12467 VPWR.n1852 VPWR.n850 3.28012
R12468 VPWR.n1954 VPWR.n850 3.28012
R12469 VPWR.n1954 VPWR.n755 3.28012
R12470 VPWR.n2048 VPWR.n755 3.28012
R12471 VPWR.n2048 VPWR.n658 3.28012
R12472 VPWR.n2150 VPWR.n658 3.28012
R12473 VPWR.n2150 VPWR.n563 3.28012
R12474 VPWR.n2244 VPWR.n563 3.28012
R12475 VPWR.n2244 VPWR.n466 3.28012
R12476 VPWR.n2346 VPWR.n466 3.28012
R12477 VPWR.n2346 VPWR.n371 3.28012
R12478 VPWR.n2440 VPWR.n371 3.28012
R12479 VPWR.n2559 VPWR.n72 3.28012
R12480 VPWR.n2433 VPWR.n72 3.28012
R12481 VPWR.n2433 VPWR.n374 3.28012
R12482 VPWR.n2353 VPWR.n374 3.28012
R12483 VPWR.n2353 VPWR.n463 3.28012
R12484 VPWR.n2237 VPWR.n463 3.28012
R12485 VPWR.n2237 VPWR.n566 3.28012
R12486 VPWR.n2157 VPWR.n566 3.28012
R12487 VPWR.n2157 VPWR.n655 3.28012
R12488 VPWR.n2041 VPWR.n655 3.28012
R12489 VPWR.n2041 VPWR.n758 3.28012
R12490 VPWR.n1961 VPWR.n758 3.28012
R12491 VPWR.n1961 VPWR.n847 3.28012
R12492 VPWR.n1845 VPWR.n847 3.28012
R12493 VPWR.n1845 VPWR.n950 3.28012
R12494 VPWR.n1539 VPWR.n1145 3.28012
R12495 VPWR.n1539 VPWR.n950 3.28012
R12496 VPWR.n1589 VPWR.n1128 3.28012
R12497 VPWR.n1128 VPWR.n934 3.28012
R12498 VPWR.n1885 VPWR.n934 3.28012
R12499 VPWR.n1885 VPWR.n863 3.28012
R12500 VPWR.n1921 VPWR.n863 3.28012
R12501 VPWR.n1921 VPWR.n742 3.28012
R12502 VPWR.n2081 VPWR.n742 3.28012
R12503 VPWR.n2081 VPWR.n671 3.28012
R12504 VPWR.n2117 VPWR.n671 3.28012
R12505 VPWR.n2117 VPWR.n550 3.28012
R12506 VPWR.n2277 VPWR.n550 3.28012
R12507 VPWR.n2277 VPWR.n479 3.28012
R12508 VPWR.n2313 VPWR.n479 3.28012
R12509 VPWR.n2313 VPWR.n358 3.28012
R12510 VPWR.n2473 VPWR.n358 3.28012
R12511 VPWR.n2473 VPWR.n96 3.28012
R12512 VPWR.n2562 VPWR.n71 3.28012
R12513 VPWR.n2430 VPWR.n71 3.28012
R12514 VPWR.n2430 VPWR.n375 3.28012
R12515 VPWR.n2356 VPWR.n375 3.28012
R12516 VPWR.n2356 VPWR.n462 3.28012
R12517 VPWR.n2234 VPWR.n462 3.28012
R12518 VPWR.n2234 VPWR.n567 3.28012
R12519 VPWR.n2160 VPWR.n567 3.28012
R12520 VPWR.n2160 VPWR.n654 3.28012
R12521 VPWR.n2038 VPWR.n654 3.28012
R12522 VPWR.n2038 VPWR.n759 3.28012
R12523 VPWR.n1964 VPWR.n759 3.28012
R12524 VPWR.n1964 VPWR.n846 3.28012
R12525 VPWR.n1842 VPWR.n846 3.28012
R12526 VPWR.n1842 VPWR.n951 3.28012
R12527 VPWR.n1532 VPWR.n951 3.28012
R12528 VPWR.n1532 VPWR.n1531 3.28012
R12529 VPWR.n1764 VPWR.n1045 3.28012
R12530 VPWR.n1764 VPWR.n954 3.28012
R12531 VPWR.n1835 VPWR.n954 3.28012
R12532 VPWR.n1835 VPWR.n843 3.28012
R12533 VPWR.n1971 VPWR.n843 3.28012
R12534 VPWR.n1971 VPWR.n762 3.28012
R12535 VPWR.n2031 VPWR.n762 3.28012
R12536 VPWR.n2031 VPWR.n651 3.28012
R12537 VPWR.n2167 VPWR.n651 3.28012
R12538 VPWR.n2167 VPWR.n570 3.28012
R12539 VPWR.n2227 VPWR.n570 3.28012
R12540 VPWR.n2227 VPWR.n459 3.28012
R12541 VPWR.n2363 VPWR.n459 3.28012
R12542 VPWR.n2363 VPWR.n378 3.28012
R12543 VPWR.n2423 VPWR.n378 3.28012
R12544 VPWR.n2423 VPWR.n66 3.28012
R12545 VPWR.n2583 VPWR.n60 3.28012
R12546 VPWR.n2413 VPWR.n60 3.28012
R12547 VPWR.n2413 VPWR.n382 3.28012
R12548 VPWR.n2373 VPWR.n382 3.28012
R12549 VPWR.n2373 VPWR.n455 3.28012
R12550 VPWR.n2217 VPWR.n455 3.28012
R12551 VPWR.n2217 VPWR.n574 3.28012
R12552 VPWR.n2177 VPWR.n574 3.28012
R12553 VPWR.n2177 VPWR.n647 3.28012
R12554 VPWR.n2021 VPWR.n647 3.28012
R12555 VPWR.n2021 VPWR.n766 3.28012
R12556 VPWR.n1981 VPWR.n766 3.28012
R12557 VPWR.n1981 VPWR.n839 3.28012
R12558 VPWR.n1825 VPWR.n839 3.28012
R12559 VPWR.n1825 VPWR.n958 3.28012
R12560 VPWR.n1752 VPWR.n958 3.28012
R12561 VPWR.n1753 VPWR.n1752 3.28012
R12562 VPWR.n1757 VPWR.n1756 3.28012
R12563 VPWR.n1757 VPWR.n955 3.28012
R12564 VPWR.n1832 VPWR.n955 3.28012
R12565 VPWR.n1832 VPWR.n842 3.28012
R12566 VPWR.n1974 VPWR.n842 3.28012
R12567 VPWR.n1974 VPWR.n763 3.28012
R12568 VPWR.n2028 VPWR.n763 3.28012
R12569 VPWR.n2028 VPWR.n650 3.28012
R12570 VPWR.n2170 VPWR.n650 3.28012
R12571 VPWR.n2170 VPWR.n571 3.28012
R12572 VPWR.n2224 VPWR.n571 3.28012
R12573 VPWR.n2224 VPWR.n458 3.28012
R12574 VPWR.n2366 VPWR.n458 3.28012
R12575 VPWR.n2366 VPWR.n379 3.28012
R12576 VPWR.n2420 VPWR.n379 3.28012
R12577 VPWR.n2420 VPWR.n65 3.28012
R12578 VPWR.n2574 VPWR.n65 3.28012
R12579 VPWR.n2586 VPWR.n59 3.28012
R12580 VPWR.n2410 VPWR.n59 3.28012
R12581 VPWR.n2410 VPWR.n383 3.28012
R12582 VPWR.n2376 VPWR.n383 3.28012
R12583 VPWR.n2376 VPWR.n454 3.28012
R12584 VPWR.n2214 VPWR.n454 3.28012
R12585 VPWR.n2214 VPWR.n575 3.28012
R12586 VPWR.n2180 VPWR.n575 3.28012
R12587 VPWR.n2180 VPWR.n646 3.28012
R12588 VPWR.n2018 VPWR.n646 3.28012
R12589 VPWR.n2018 VPWR.n767 3.28012
R12590 VPWR.n1984 VPWR.n767 3.28012
R12591 VPWR.n1984 VPWR.n838 3.28012
R12592 VPWR.n1822 VPWR.n838 3.28012
R12593 VPWR.n1822 VPWR.n959 3.28012
R12594 VPWR.n1788 VPWR.n959 3.28012
R12595 VPWR.n1788 VPWR.n1037 3.28012
R12596 VPWR.n1465 VPWR.n1232 3.28012
R12597 VPWR.n1465 VPWR.n931 3.28012
R12598 VPWR.n1892 VPWR.n931 3.28012
R12599 VPWR.n1892 VPWR.n929 3.28012
R12600 VPWR.n1914 VPWR.n929 3.28012
R12601 VPWR.n1914 VPWR.n739 3.28012
R12602 VPWR.n2088 VPWR.n739 3.28012
R12603 VPWR.n2088 VPWR.n737 3.28012
R12604 VPWR.n2110 VPWR.n737 3.28012
R12605 VPWR.n2110 VPWR.n547 3.28012
R12606 VPWR.n2284 VPWR.n547 3.28012
R12607 VPWR.n2284 VPWR.n545 3.28012
R12608 VPWR.n2306 VPWR.n545 3.28012
R12609 VPWR.n2306 VPWR.n355 3.28012
R12610 VPWR.n2480 VPWR.n355 3.28012
R12611 VPWR.n2480 VPWR.n353 3.28012
R12612 VPWR.n2502 VPWR.n353 3.28012
R12613 VPWR.n2404 VPWR.n22 3.28012
R12614 VPWR.n2404 VPWR.n449 3.28012
R12615 VPWR.n2382 VPWR.n449 3.28012
R12616 VPWR.n2382 VPWR.n451 3.28012
R12617 VPWR.n2208 VPWR.n451 3.28012
R12618 VPWR.n2208 VPWR.n641 3.28012
R12619 VPWR.n2186 VPWR.n641 3.28012
R12620 VPWR.n2186 VPWR.n643 3.28012
R12621 VPWR.n2012 VPWR.n643 3.28012
R12622 VPWR.n2012 VPWR.n833 3.28012
R12623 VPWR.n1990 VPWR.n833 3.28012
R12624 VPWR.n1990 VPWR.n835 3.28012
R12625 VPWR.n1816 VPWR.n835 3.28012
R12626 VPWR.n1816 VPWR.n1025 3.28012
R12627 VPWR.n1794 VPWR.n1025 3.28012
R12628 VPWR.n1794 VPWR.n1028 3.28012
R12629 VPWR.n2594 VPWR.n22 3.26393
R12630 VPWR.n2863 VPWR 3.18182
R12631 VPWR.n2832 VPWR.n2831 3.1005
R12632 VPWR.n2826 VPWR.n2825 3.1005
R12633 VPWR.n2846 VPWR.n2815 3.1005
R12634 VPWR.n1324 VPWR.n1322 3.01226
R12635 VPWR.n1328 VPWR.n1304 2.63579
R12636 VPWR.n2731 VPWR.n2730 2.25932
R12637 VPWR.n1447 VPWR.n1446 2.06026
R12638 VPWR.n1447 VPWR.n1026 1.78803
R12639 VPWR.n2384 VPWR.n2383 1.32852
R12640 VPWR.n2287 VPWR.n450 1.32852
R12641 VPWR.n2207 VPWR.n2206 1.32852
R12642 VPWR.n2205 VPWR.n2204 1.32852
R12643 VPWR.n2188 VPWR.n2187 1.32852
R12644 VPWR.n2091 VPWR.n642 1.32852
R12645 VPWR.n2011 VPWR.n2010 1.32852
R12646 VPWR.n2009 VPWR.n2008 1.32852
R12647 VPWR.n1992 VPWR.n1991 1.32852
R12648 VPWR.n1895 VPWR.n834 1.32852
R12649 VPWR.n2401 VPWR.n2400 1.32852
R12650 VPWR.n1815 VPWR.n1814 1.32852
R12651 VPWR.n2403 VPWR.n2402 1.32852
R12652 VPWR.n1813 VPWR.n1812 1.32852
R12653 VPWR.n2483 VPWR.n21 1.32852
R12654 VPWR.n1796 VPWR.n1795 1.32852
R12655 VPWR.n2596 VPWR.n2595 1.32852
R12656 VPWR.n1055 VPWR.n1026 1.32852
R12657 VPWR.n2482 VPWR 1.25994
R12658 VPWR VPWR.n354 1.25994
R12659 VPWR VPWR.n2304 1.25994
R12660 VPWR.n2303 VPWR 1.25994
R12661 VPWR.n2286 VPWR 1.25994
R12662 VPWR VPWR.n546 1.25994
R12663 VPWR VPWR.n2108 1.25994
R12664 VPWR.n2107 VPWR 1.25994
R12665 VPWR.n2090 VPWR 1.25994
R12666 VPWR VPWR.n738 1.25994
R12667 VPWR VPWR.n1912 1.25994
R12668 VPWR.n1911 VPWR 1.25994
R12669 VPWR.n1894 VPWR 1.25994
R12670 VPWR VPWR.n930 1.25994
R12671 VPWR.n2499 VPWR 1.25994
R12672 VPWR VPWR.n1450 1.25994
R12673 VPWR VPWR.n2500 1.25994
R12674 VPWR.n1449 VPWR 1.25994
R12675 VPWR.n2597 VPWR.n2596 1.144
R12676 VPWR.n2861 VPWR.n2860 0.936724
R12677 VPWR.n2592 VPWR 0.925943
R12678 VPWR VPWR.n1063 0.925943
R12679 VPWR.n2860 VPWR.n2816 0.925245
R12680 VPWR.n2569 VPWR.n67 0.904391
R12681 VPWR.n2509 VPWR.n97 0.904391
R12682 VPWR.n2552 VPWR.n76 0.904391
R12683 VPWR.n2545 VPWR.n79 0.904391
R12684 VPWR.n2533 VPWR.n85 0.904391
R12685 VPWR.n2528 VPWR.n88 0.904391
R12686 VPWR.n1222 VPWR.n1178 0.904391
R12687 VPWR.n2521 VPWR.n91 0.904391
R12688 VPWR.n1624 VPWR.n1102 0.904391
R12689 VPWR.n1640 VPWR.n1094 0.904391
R12690 VPWR.n2540 VPWR.n82 0.904391
R12691 VPWR.n1651 VPWR.n1092 0.904391
R12692 VPWR.n1211 VPWR.n1210 0.904391
R12693 VPWR.n2516 VPWR.n94 0.904391
R12694 VPWR.n1613 VPWR.n1104 0.904391
R12695 VPWR.n1667 VPWR.n1084 0.904391
R12696 VPWR.n2557 VPWR.n73 0.904391
R12697 VPWR.n1678 VPWR.n1082 0.904391
R12698 VPWR.n1591 VPWR.n1127 0.904391
R12699 VPWR.n2564 VPWR.n70 0.904391
R12700 VPWR.n1197 VPWR.n1196 0.904391
R12701 VPWR.n1694 VPWR.n1074 0.904391
R12702 VPWR.n1742 VPWR.n1057 0.904391
R12703 VPWR.n1705 VPWR.n1071 0.904391
R12704 VPWR.n2581 VPWR.n61 0.904391
R12705 VPWR.n2588 VPWR.n58 0.904391
R12706 VPWR.n1737 VPWR.n1735 0.904391
R12707 VPWR.n1597 VPWR.n1596 0.904391
R12708 VPWR.n2504 VPWR.n289 0.904391
R12709 VPWR.n2576 VPWR.n64 0.904391
R12710 VPWR VPWR.n2863 0.812229
R12711 VPWR.n140 VPWR.n64 0.675548
R12712 VPWR.n152 VPWR.n67 0.675548
R12713 VPWR.n164 VPWR.n70 0.675548
R12714 VPWR.n176 VPWR.n73 0.675548
R12715 VPWR.n188 VPWR.n76 0.675548
R12716 VPWR.n200 VPWR.n79 0.675548
R12717 VPWR.n212 VPWR.n82 0.675548
R12718 VPWR.n224 VPWR.n85 0.675548
R12719 VPWR.n236 VPWR.n88 0.675548
R12720 VPWR.n248 VPWR.n91 0.675548
R12721 VPWR.n260 VPWR.n94 0.675548
R12722 VPWR.n272 VPWR.n97 0.675548
R12723 VPWR.n289 VPWR.n288 0.675548
R12724 VPWR.n128 VPWR.n61 0.675548
R12725 VPWR.n117 VPWR.n58 0.675548
R12726 VPWR.n1735 VPWR.n1734 0.675548
R12727 VPWR.n1719 VPWR.n1057 0.675548
R12728 VPWR.n1707 VPWR.n1705 0.675548
R12729 VPWR.n1696 VPWR.n1694 0.675548
R12730 VPWR.n1196 VPWR.n1195 0.675548
R12731 VPWR.n1680 VPWR.n1678 0.675548
R12732 VPWR.n1669 VPWR.n1667 0.675548
R12733 VPWR.n1210 VPWR.n1209 0.675548
R12734 VPWR.n1653 VPWR.n1651 0.675548
R12735 VPWR.n1642 VPWR.n1640 0.675548
R12736 VPWR.n1178 VPWR.n1177 0.675548
R12737 VPWR.n1626 VPWR.n1624 0.675548
R12738 VPWR.n1615 VPWR.n1613 0.675548
R12739 VPWR.n1127 VPWR.n1126 0.675548
R12740 VPWR.n1599 VPWR.n1597 0.675548
R12741 VPWR.n2806 VPWR.n2805 0.672385
R12742 VPWR.n2790 VPWR.n2785 0.672385
R12743 VPWR.n2770 VPWR.n2765 0.672385
R12744 VPWR.n2751 VPWR.n2746 0.672385
R12745 VPWR.n7 VPWR 0.63497
R12746 VPWR.n1242 VPWR 0.63497
R12747 VPWR.n1265 VPWR 0.63497
R12748 VPWR.n1289 VPWR 0.63497
R12749 VPWR.n24 VPWR 0.499542
R12750 VPWR.n2814 VPWR.n2813 0.442692
R12751 VPWR.n1120 VPWR.n1118 0.404056
R12752 VPWR.n144 VPWR.n138 0.404056
R12753 VPWR.n156 VPWR.n150 0.404056
R12754 VPWR.n168 VPWR.n162 0.404056
R12755 VPWR.n180 VPWR.n174 0.404056
R12756 VPWR.n192 VPWR.n186 0.404056
R12757 VPWR.n204 VPWR.n198 0.404056
R12758 VPWR.n216 VPWR.n210 0.404056
R12759 VPWR.n228 VPWR.n222 0.404056
R12760 VPWR.n240 VPWR.n234 0.404056
R12761 VPWR.n252 VPWR.n246 0.404056
R12762 VPWR.n264 VPWR.n258 0.404056
R12763 VPWR.n276 VPWR.n270 0.404056
R12764 VPWR.n283 VPWR.n101 0.404056
R12765 VPWR.n110 VPWR.n105 0.404056
R12766 VPWR.n132 VPWR.n126 0.404056
R12767 VPWR.n121 VPWR.n115 0.404056
R12768 VPWR.n1729 VPWR.n1065 0.404056
R12769 VPWR.n1723 VPWR.n1717 0.404056
R12770 VPWR.n1711 VPWR.n1070 0.404056
R12771 VPWR.n1704 VPWR.n1702 0.404056
R12772 VPWR.n1693 VPWR.n1691 0.404056
R12773 VPWR.n1684 VPWR.n1081 0.404056
R12774 VPWR.n1677 VPWR.n1675 0.404056
R12775 VPWR.n1666 VPWR.n1664 0.404056
R12776 VPWR.n1657 VPWR.n1091 0.404056
R12777 VPWR.n1650 VPWR.n1648 0.404056
R12778 VPWR.n1639 VPWR.n1637 0.404056
R12779 VPWR.n1630 VPWR.n1101 0.404056
R12780 VPWR.n1623 VPWR.n1621 0.404056
R12781 VPWR.n1612 VPWR.n1610 0.404056
R12782 VPWR.n1603 VPWR.n1111 0.404056
R12783 VPWR.n2860 VPWR.n2859 0.388
R12784 VPWR.n1608 VPWR.n1607 0.349144
R12785 VPWR.n1608 VPWR.n1099 0.349144
R12786 VPWR.n1634 VPWR.n1099 0.349144
R12787 VPWR.n1635 VPWR.n1634 0.349144
R12788 VPWR.n1635 VPWR.n1089 0.349144
R12789 VPWR.n1661 VPWR.n1089 0.349144
R12790 VPWR.n1662 VPWR.n1661 0.349144
R12791 VPWR.n1662 VPWR.n1079 0.349144
R12792 VPWR.n1688 VPWR.n1079 0.349144
R12793 VPWR.n1689 VPWR.n1688 0.349144
R12794 VPWR.n1689 VPWR.n1068 0.349144
R12795 VPWR.n1715 VPWR.n1068 0.349144
R12796 VPWR.n1727 VPWR.n1715 0.349144
R12797 VPWR.n281 VPWR.n280 0.349144
R12798 VPWR.n280 VPWR.n268 0.349144
R12799 VPWR.n268 VPWR.n256 0.349144
R12800 VPWR.n256 VPWR.n244 0.349144
R12801 VPWR.n244 VPWR.n232 0.349144
R12802 VPWR.n232 VPWR.n220 0.349144
R12803 VPWR.n220 VPWR.n208 0.349144
R12804 VPWR.n208 VPWR.n196 0.349144
R12805 VPWR.n196 VPWR.n184 0.349144
R12806 VPWR.n184 VPWR.n172 0.349144
R12807 VPWR.n172 VPWR.n160 0.349144
R12808 VPWR.n160 VPWR.n148 0.349144
R12809 VPWR.n148 VPWR.n136 0.349144
R12810 VPWR.n1462 VPWR.n1456 0.346131
R12811 VPWR.n1461 VPWR.n1457 0.346131
R12812 VPWR.n1582 VPWR.n1136 0.346131
R12813 VPWR.n1581 VPWR.n1577 0.346131
R12814 VPWR.n1576 VPWR.n1572 0.346131
R12815 VPWR.n1571 VPWR.n1567 0.346131
R12816 VPWR.n1566 VPWR.n1562 0.346131
R12817 VPWR.n1561 VPWR.n1557 0.346131
R12818 VPWR.n1556 VPWR.n1552 0.346131
R12819 VPWR.n1551 VPWR.n1547 0.346131
R12820 VPWR.n1546 VPWR.n1542 0.346131
R12821 VPWR.n1767 VPWR.n1042 0.346131
R12822 VPWR.n1784 VPWR.n1780 0.346131
R12823 VPWR.n1785 VPWR.n1776 0.346131
R12824 VPWR.n1772 VPWR.n1771 0.346131
R12825 VPWR.n2862 VPWR.n2861 0.304571
R12826 VPWR.n2594 VPWR.n55 0.300179
R12827 VPWR.n1118 VPWR.n1113 0.286958
R12828 VPWR.n145 VPWR.n144 0.286958
R12829 VPWR.n157 VPWR.n156 0.286958
R12830 VPWR.n169 VPWR.n168 0.286958
R12831 VPWR.n181 VPWR.n180 0.286958
R12832 VPWR.n193 VPWR.n192 0.286958
R12833 VPWR.n205 VPWR.n204 0.286958
R12834 VPWR.n217 VPWR.n216 0.286958
R12835 VPWR.n229 VPWR.n228 0.286958
R12836 VPWR.n241 VPWR.n240 0.286958
R12837 VPWR.n253 VPWR.n252 0.286958
R12838 VPWR.n265 VPWR.n264 0.286958
R12839 VPWR.n277 VPWR.n276 0.286958
R12840 VPWR.n283 VPWR.n102 0.286958
R12841 VPWR.n111 VPWR.n110 0.286958
R12842 VPWR.n133 VPWR.n132 0.286958
R12843 VPWR.n122 VPWR.n121 0.286958
R12844 VPWR.n1729 VPWR.n1066 0.286958
R12845 VPWR.n1724 VPWR.n1723 0.286958
R12846 VPWR.n1712 VPWR.n1711 0.286958
R12847 VPWR.n1702 VPWR.n1072 0.286958
R12848 VPWR.n1691 VPWR.n1075 0.286958
R12849 VPWR.n1685 VPWR.n1684 0.286958
R12850 VPWR.n1675 VPWR.n1083 0.286958
R12851 VPWR.n1664 VPWR.n1085 0.286958
R12852 VPWR.n1658 VPWR.n1657 0.286958
R12853 VPWR.n1648 VPWR.n1093 0.286958
R12854 VPWR.n1637 VPWR.n1095 0.286958
R12855 VPWR.n1631 VPWR.n1630 0.286958
R12856 VPWR.n1621 VPWR.n1103 0.286958
R12857 VPWR.n1610 VPWR.n1105 0.286958
R12858 VPWR.n1604 VPWR.n1603 0.286958
R12859 VPWR.n55 VPWR 0.2505
R12860 VPWR VPWR.n2481 0.249238
R12861 VPWR.n2472 VPWR 0.249238
R12862 VPWR VPWR.n2471 0.249238
R12863 VPWR.n2385 VPWR 0.249238
R12864 VPWR.n2386 VPWR 0.249238
R12865 VPWR.n2387 VPWR 0.249238
R12866 VPWR.n2388 VPWR 0.249238
R12867 VPWR.n2305 VPWR 0.249238
R12868 VPWR.n2314 VPWR 0.249238
R12869 VPWR.n2315 VPWR 0.249238
R12870 VPWR.n2324 VPWR 0.249238
R12871 VPWR.n2325 VPWR 0.249238
R12872 VPWR.n2383 VPWR 0.249238
R12873 VPWR.n2375 VPWR 0.249238
R12874 VPWR.n2374 VPWR 0.249238
R12875 VPWR.n2365 VPWR 0.249238
R12876 VPWR.n2364 VPWR 0.249238
R12877 VPWR.n2355 VPWR 0.249238
R12878 VPWR.n2354 VPWR 0.249238
R12879 VPWR.n2345 VPWR 0.249238
R12880 VPWR.n2344 VPWR 0.249238
R12881 VPWR.n2335 VPWR 0.249238
R12882 VPWR.n2334 VPWR 0.249238
R12883 VPWR VPWR.n2302 0.249238
R12884 VPWR VPWR.n2301 0.249238
R12885 VPWR VPWR.n2300 0.249238
R12886 VPWR VPWR.n2299 0.249238
R12887 VPWR VPWR.n2298 0.249238
R12888 VPWR VPWR.n2287 0.249238
R12889 VPWR VPWR.n2288 0.249238
R12890 VPWR VPWR.n2289 0.249238
R12891 VPWR VPWR.n2290 0.249238
R12892 VPWR VPWR.n2291 0.249238
R12893 VPWR VPWR.n2292 0.249238
R12894 VPWR VPWR.n2293 0.249238
R12895 VPWR VPWR.n2294 0.249238
R12896 VPWR VPWR.n2295 0.249238
R12897 VPWR VPWR.n2296 0.249238
R12898 VPWR VPWR.n2297 0.249238
R12899 VPWR VPWR.n2285 0.249238
R12900 VPWR.n2276 VPWR 0.249238
R12901 VPWR VPWR.n2275 0.249238
R12902 VPWR.n2266 VPWR 0.249238
R12903 VPWR VPWR.n2265 0.249238
R12904 VPWR.n2207 VPWR 0.249238
R12905 VPWR VPWR.n2215 0.249238
R12906 VPWR.n2216 VPWR 0.249238
R12907 VPWR VPWR.n2225 0.249238
R12908 VPWR.n2226 VPWR 0.249238
R12909 VPWR VPWR.n2235 0.249238
R12910 VPWR.n2236 VPWR 0.249238
R12911 VPWR VPWR.n2245 0.249238
R12912 VPWR.n2246 VPWR 0.249238
R12913 VPWR VPWR.n2255 0.249238
R12914 VPWR.n2256 VPWR 0.249238
R12915 VPWR.n2189 VPWR 0.249238
R12916 VPWR.n2190 VPWR 0.249238
R12917 VPWR.n2191 VPWR 0.249238
R12918 VPWR.n2192 VPWR 0.249238
R12919 VPWR.n2193 VPWR 0.249238
R12920 VPWR.n2204 VPWR 0.249238
R12921 VPWR.n2203 VPWR 0.249238
R12922 VPWR.n2202 VPWR 0.249238
R12923 VPWR.n2201 VPWR 0.249238
R12924 VPWR.n2200 VPWR 0.249238
R12925 VPWR.n2199 VPWR 0.249238
R12926 VPWR.n2198 VPWR 0.249238
R12927 VPWR.n2197 VPWR 0.249238
R12928 VPWR.n2196 VPWR 0.249238
R12929 VPWR.n2195 VPWR 0.249238
R12930 VPWR.n2194 VPWR 0.249238
R12931 VPWR.n2109 VPWR 0.249238
R12932 VPWR.n2118 VPWR 0.249238
R12933 VPWR.n2119 VPWR 0.249238
R12934 VPWR.n2128 VPWR 0.249238
R12935 VPWR.n2129 VPWR 0.249238
R12936 VPWR.n2187 VPWR 0.249238
R12937 VPWR.n2179 VPWR 0.249238
R12938 VPWR.n2178 VPWR 0.249238
R12939 VPWR.n2169 VPWR 0.249238
R12940 VPWR.n2168 VPWR 0.249238
R12941 VPWR.n2159 VPWR 0.249238
R12942 VPWR.n2158 VPWR 0.249238
R12943 VPWR.n2149 VPWR 0.249238
R12944 VPWR.n2148 VPWR 0.249238
R12945 VPWR.n2139 VPWR 0.249238
R12946 VPWR.n2138 VPWR 0.249238
R12947 VPWR VPWR.n2106 0.249238
R12948 VPWR VPWR.n2105 0.249238
R12949 VPWR VPWR.n2104 0.249238
R12950 VPWR VPWR.n2103 0.249238
R12951 VPWR VPWR.n2102 0.249238
R12952 VPWR VPWR.n2091 0.249238
R12953 VPWR VPWR.n2092 0.249238
R12954 VPWR VPWR.n2093 0.249238
R12955 VPWR VPWR.n2094 0.249238
R12956 VPWR VPWR.n2095 0.249238
R12957 VPWR VPWR.n2096 0.249238
R12958 VPWR VPWR.n2097 0.249238
R12959 VPWR VPWR.n2098 0.249238
R12960 VPWR VPWR.n2099 0.249238
R12961 VPWR VPWR.n2100 0.249238
R12962 VPWR VPWR.n2101 0.249238
R12963 VPWR VPWR.n2089 0.249238
R12964 VPWR.n2080 VPWR 0.249238
R12965 VPWR VPWR.n2079 0.249238
R12966 VPWR.n2070 VPWR 0.249238
R12967 VPWR VPWR.n2069 0.249238
R12968 VPWR.n2011 VPWR 0.249238
R12969 VPWR VPWR.n2019 0.249238
R12970 VPWR.n2020 VPWR 0.249238
R12971 VPWR VPWR.n2029 0.249238
R12972 VPWR.n2030 VPWR 0.249238
R12973 VPWR VPWR.n2039 0.249238
R12974 VPWR.n2040 VPWR 0.249238
R12975 VPWR VPWR.n2049 0.249238
R12976 VPWR.n2050 VPWR 0.249238
R12977 VPWR VPWR.n2059 0.249238
R12978 VPWR.n2060 VPWR 0.249238
R12979 VPWR.n1993 VPWR 0.249238
R12980 VPWR.n1994 VPWR 0.249238
R12981 VPWR.n1995 VPWR 0.249238
R12982 VPWR.n1996 VPWR 0.249238
R12983 VPWR.n1997 VPWR 0.249238
R12984 VPWR.n2008 VPWR 0.249238
R12985 VPWR.n2007 VPWR 0.249238
R12986 VPWR.n2006 VPWR 0.249238
R12987 VPWR.n2005 VPWR 0.249238
R12988 VPWR.n2004 VPWR 0.249238
R12989 VPWR.n2003 VPWR 0.249238
R12990 VPWR.n2002 VPWR 0.249238
R12991 VPWR.n2001 VPWR 0.249238
R12992 VPWR.n2000 VPWR 0.249238
R12993 VPWR.n1999 VPWR 0.249238
R12994 VPWR.n1998 VPWR 0.249238
R12995 VPWR.n1913 VPWR 0.249238
R12996 VPWR.n1922 VPWR 0.249238
R12997 VPWR.n1923 VPWR 0.249238
R12998 VPWR.n1932 VPWR 0.249238
R12999 VPWR.n1933 VPWR 0.249238
R13000 VPWR.n1991 VPWR 0.249238
R13001 VPWR.n1983 VPWR 0.249238
R13002 VPWR.n1982 VPWR 0.249238
R13003 VPWR.n1973 VPWR 0.249238
R13004 VPWR.n1972 VPWR 0.249238
R13005 VPWR.n1963 VPWR 0.249238
R13006 VPWR.n1962 VPWR 0.249238
R13007 VPWR.n1953 VPWR 0.249238
R13008 VPWR.n1952 VPWR 0.249238
R13009 VPWR.n1943 VPWR 0.249238
R13010 VPWR.n1942 VPWR 0.249238
R13011 VPWR VPWR.n1910 0.249238
R13012 VPWR VPWR.n1909 0.249238
R13013 VPWR VPWR.n1908 0.249238
R13014 VPWR VPWR.n1907 0.249238
R13015 VPWR VPWR.n1906 0.249238
R13016 VPWR VPWR.n1895 0.249238
R13017 VPWR VPWR.n1896 0.249238
R13018 VPWR VPWR.n1897 0.249238
R13019 VPWR VPWR.n1898 0.249238
R13020 VPWR VPWR.n1899 0.249238
R13021 VPWR VPWR.n1900 0.249238
R13022 VPWR VPWR.n1901 0.249238
R13023 VPWR VPWR.n1902 0.249238
R13024 VPWR VPWR.n1903 0.249238
R13025 VPWR VPWR.n1904 0.249238
R13026 VPWR VPWR.n1905 0.249238
R13027 VPWR.n2400 VPWR 0.249238
R13028 VPWR.n2399 VPWR 0.249238
R13029 VPWR.n2398 VPWR 0.249238
R13030 VPWR.n2397 VPWR 0.249238
R13031 VPWR.n2396 VPWR 0.249238
R13032 VPWR.n2395 VPWR 0.249238
R13033 VPWR.n2394 VPWR 0.249238
R13034 VPWR.n2393 VPWR 0.249238
R13035 VPWR.n2392 VPWR 0.249238
R13036 VPWR.n2391 VPWR 0.249238
R13037 VPWR.n2390 VPWR 0.249238
R13038 VPWR.n2389 VPWR 0.249238
R13039 VPWR VPWR.n1893 0.249238
R13040 VPWR.n1884 VPWR 0.249238
R13041 VPWR VPWR.n1883 0.249238
R13042 VPWR.n1874 VPWR 0.249238
R13043 VPWR VPWR.n1873 0.249238
R13044 VPWR.n1864 VPWR 0.249238
R13045 VPWR.n1815 VPWR 0.249238
R13046 VPWR VPWR.n1823 0.249238
R13047 VPWR.n1824 VPWR 0.249238
R13048 VPWR VPWR.n1833 0.249238
R13049 VPWR.n1834 VPWR 0.249238
R13050 VPWR VPWR.n1843 0.249238
R13051 VPWR.n1844 VPWR 0.249238
R13052 VPWR VPWR.n1853 0.249238
R13053 VPWR.n1854 VPWR 0.249238
R13054 VPWR VPWR.n1863 0.249238
R13055 VPWR.n2403 VPWR 0.249238
R13056 VPWR VPWR.n2411 0.249238
R13057 VPWR.n2412 VPWR 0.249238
R13058 VPWR VPWR.n2421 0.249238
R13059 VPWR.n2422 VPWR 0.249238
R13060 VPWR VPWR.n2431 0.249238
R13061 VPWR.n2432 VPWR 0.249238
R13062 VPWR VPWR.n2441 0.249238
R13063 VPWR.n2442 VPWR 0.249238
R13064 VPWR VPWR.n2451 0.249238
R13065 VPWR.n2452 VPWR 0.249238
R13066 VPWR VPWR.n2461 0.249238
R13067 VPWR.n2462 VPWR 0.249238
R13068 VPWR.n1797 VPWR 0.249238
R13069 VPWR.n1798 VPWR 0.249238
R13070 VPWR.n1799 VPWR 0.249238
R13071 VPWR.n1800 VPWR 0.249238
R13072 VPWR.n1801 VPWR 0.249238
R13073 VPWR.n1802 VPWR 0.249238
R13074 VPWR.n1803 VPWR 0.249238
R13075 VPWR.n1804 VPWR 0.249238
R13076 VPWR.n1805 VPWR 0.249238
R13077 VPWR.n1812 VPWR 0.249238
R13078 VPWR.n1811 VPWR 0.249238
R13079 VPWR.n1810 VPWR 0.249238
R13080 VPWR.n1809 VPWR 0.249238
R13081 VPWR.n1808 VPWR 0.249238
R13082 VPWR.n1807 VPWR 0.249238
R13083 VPWR.n1806 VPWR 0.249238
R13084 VPWR VPWR.n2498 0.249238
R13085 VPWR VPWR.n2497 0.249238
R13086 VPWR VPWR.n2496 0.249238
R13087 VPWR VPWR.n2495 0.249238
R13088 VPWR VPWR.n2494 0.249238
R13089 VPWR VPWR.n2493 0.249238
R13090 VPWR VPWR.n2492 0.249238
R13091 VPWR VPWR.n2491 0.249238
R13092 VPWR VPWR.n2490 0.249238
R13093 VPWR VPWR.n2489 0.249238
R13094 VPWR VPWR.n2488 0.249238
R13095 VPWR VPWR.n2483 0.249238
R13096 VPWR VPWR.n2484 0.249238
R13097 VPWR VPWR.n2485 0.249238
R13098 VPWR VPWR.n2486 0.249238
R13099 VPWR VPWR.n2487 0.249238
R13100 VPWR.n2501 VPWR 0.249238
R13101 VPWR.n2512 VPWR 0.249238
R13102 VPWR.n2513 VPWR 0.249238
R13103 VPWR.n2524 VPWR 0.249238
R13104 VPWR.n2525 VPWR 0.249238
R13105 VPWR.n2536 VPWR 0.249238
R13106 VPWR.n2537 VPWR 0.249238
R13107 VPWR.n2548 VPWR 0.249238
R13108 VPWR.n2549 VPWR 0.249238
R13109 VPWR.n2560 VPWR 0.249238
R13110 VPWR.n2561 VPWR 0.249238
R13111 VPWR.n2572 VPWR 0.249238
R13112 VPWR.n2573 VPWR 0.249238
R13113 VPWR.n2584 VPWR 0.249238
R13114 VPWR.n2585 VPWR 0.249238
R13115 VPWR.n2595 VPWR 0.249238
R13116 VPWR VPWR.n1055 0.249238
R13117 VPWR VPWR.n1056 0.249238
R13118 VPWR VPWR.n1754 0.249238
R13119 VPWR.n1755 VPWR 0.249238
R13120 VPWR VPWR.n1529 0.249238
R13121 VPWR.n1530 VPWR 0.249238
R13122 VPWR.n1528 VPWR 0.249238
R13123 VPWR.n1527 VPWR 0.249238
R13124 VPWR.n1514 VPWR 0.249238
R13125 VPWR.n1513 VPWR 0.249238
R13126 VPWR.n1500 VPWR 0.249238
R13127 VPWR.n1499 VPWR 0.249238
R13128 VPWR.n1487 VPWR 0.249238
R13129 VPWR VPWR.n1587 0.249238
R13130 VPWR.n1588 VPWR 0.249238
R13131 VPWR VPWR.n1448 0.249238
R13132 VPWR.n2861 VPWR.n2815 0.245065
R13133 VPWR.n2813 VPWR.n2797 0.213567
R13134 VPWR.n2797 VPWR.n2778 0.213567
R13135 VPWR.n2778 VPWR.n2758 0.213567
R13136 VPWR.n2758 VPWR.n2739 0.213567
R13137 VPWR.n2739 VPWR.n2703 0.213567
R13138 VPWR.n2703 VPWR.n2665 0.213567
R13139 VPWR.n2665 VPWR.n2628 0.213567
R13140 VPWR.n1446 VPWR.n1414 0.213567
R13141 VPWR.n1414 VPWR.n1376 0.213567
R13142 VPWR.n1376 VPWR.n1337 0.213567
R13143 VPWR.n1337 VPWR.n1302 0.213567
R13144 VPWR.n1302 VPWR.n1279 0.213567
R13145 VPWR.n1279 VPWR.n1255 0.213567
R13146 VPWR.n1255 VPWR.n19 0.213567
R13147 VPWR VPWR.n2862 0.204304
R13148 VPWR.n1449 VPWR.n1447 0.179202
R13149 VPWR.n1450 VPWR.n1449 0.154425
R13150 VPWR.n1450 VPWR.n930 0.154425
R13151 VPWR.n1894 VPWR.n930 0.154425
R13152 VPWR.n1911 VPWR.n1894 0.154425
R13153 VPWR.n1912 VPWR.n1911 0.154425
R13154 VPWR.n1912 VPWR.n738 0.154425
R13155 VPWR.n2090 VPWR.n738 0.154425
R13156 VPWR.n2107 VPWR.n2090 0.154425
R13157 VPWR.n2108 VPWR.n2107 0.154425
R13158 VPWR.n2108 VPWR.n546 0.154425
R13159 VPWR.n2286 VPWR.n546 0.154425
R13160 VPWR.n2303 VPWR.n2286 0.154425
R13161 VPWR.n2304 VPWR.n2303 0.154425
R13162 VPWR.n2304 VPWR.n354 0.154425
R13163 VPWR.n2482 VPWR.n354 0.154425
R13164 VPWR.n2499 VPWR.n2482 0.154425
R13165 VPWR.n2500 VPWR.n2499 0.154425
R13166 VPWR.n1796 VPWR.n1026 0.154425
R13167 VPWR.n1813 VPWR.n1796 0.154425
R13168 VPWR.n1814 VPWR.n1813 0.154425
R13169 VPWR.n1814 VPWR.n834 0.154425
R13170 VPWR.n1992 VPWR.n834 0.154425
R13171 VPWR.n2009 VPWR.n1992 0.154425
R13172 VPWR.n2010 VPWR.n2009 0.154425
R13173 VPWR.n2010 VPWR.n642 0.154425
R13174 VPWR.n2188 VPWR.n642 0.154425
R13175 VPWR.n2205 VPWR.n2188 0.154425
R13176 VPWR.n2206 VPWR.n2205 0.154425
R13177 VPWR.n2206 VPWR.n450 0.154425
R13178 VPWR.n2384 VPWR.n450 0.154425
R13179 VPWR.n2401 VPWR.n2384 0.154425
R13180 VPWR.n2402 VPWR.n2401 0.154425
R13181 VPWR.n2402 VPWR.n21 0.154425
R13182 VPWR.n2596 VPWR.n21 0.154425
R13183 VPWR.n8 VPWR.n7 0.147771
R13184 VPWR.n1243 VPWR.n1242 0.147771
R13185 VPWR.n1266 VPWR.n1265 0.147771
R13186 VPWR.n1290 VPWR.n1289 0.147771
R13187 VPWR.n1113 VPWR 0.135917
R13188 VPWR.n145 VPWR 0.135917
R13189 VPWR.n157 VPWR 0.135917
R13190 VPWR.n169 VPWR 0.135917
R13191 VPWR.n181 VPWR 0.135917
R13192 VPWR.n193 VPWR 0.135917
R13193 VPWR.n205 VPWR 0.135917
R13194 VPWR.n217 VPWR 0.135917
R13195 VPWR.n229 VPWR 0.135917
R13196 VPWR.n241 VPWR 0.135917
R13197 VPWR.n253 VPWR 0.135917
R13198 VPWR.n265 VPWR 0.135917
R13199 VPWR.n277 VPWR 0.135917
R13200 VPWR.n102 VPWR 0.135917
R13201 VPWR.n111 VPWR 0.135917
R13202 VPWR.n133 VPWR 0.135917
R13203 VPWR.n122 VPWR 0.135917
R13204 VPWR.n1066 VPWR 0.135917
R13205 VPWR.n1724 VPWR 0.135917
R13206 VPWR.n1712 VPWR 0.135917
R13207 VPWR.n1072 VPWR 0.135917
R13208 VPWR.n1075 VPWR 0.135917
R13209 VPWR.n1685 VPWR 0.135917
R13210 VPWR.n1083 VPWR 0.135917
R13211 VPWR.n1085 VPWR 0.135917
R13212 VPWR.n1658 VPWR 0.135917
R13213 VPWR.n1093 VPWR 0.135917
R13214 VPWR.n1095 VPWR 0.135917
R13215 VPWR.n1631 VPWR 0.135917
R13216 VPWR.n1103 VPWR 0.135917
R13217 VPWR.n1105 VPWR 0.135917
R13218 VPWR.n1604 VPWR 0.135917
R13219 VPWR.n2863 VPWR.n2814 0.127988
R13220 VPWR.n2825 VPWR.n2816 0.1255
R13221 VPWR.n2831 VPWR.n2816 0.1255
R13222 VPWR.n18 VPWR.n0 0.120292
R13223 VPWR.n14 VPWR.n0 0.120292
R13224 VPWR.n9 VPWR.n8 0.120292
R13225 VPWR.n1254 VPWR.n1233 0.120292
R13226 VPWR.n1250 VPWR.n1233 0.120292
R13227 VPWR.n1244 VPWR.n1243 0.120292
R13228 VPWR.n1278 VPWR.n1256 0.120292
R13229 VPWR.n1273 VPWR.n1256 0.120292
R13230 VPWR.n1267 VPWR.n1266 0.120292
R13231 VPWR.n1301 VPWR.n1280 0.120292
R13232 VPWR.n1297 VPWR.n1280 0.120292
R13233 VPWR.n1291 VPWR.n1290 0.120292
R13234 VPWR.n1333 VPWR.n1332 0.120292
R13235 VPWR.n1326 VPWR.n1305 0.120292
R13236 VPWR.n1319 VPWR.n1305 0.120292
R13237 VPWR.n1319 VPWR.n1318 0.120292
R13238 VPWR.n1317 VPWR.n1309 0.120292
R13239 VPWR.n1312 VPWR.n1309 0.120292
R13240 VPWR.n1312 VPWR.n1311 0.120292
R13241 VPWR.n1371 VPWR.n1370 0.120292
R13242 VPWR.n1364 VPWR.n1363 0.120292
R13243 VPWR.n1363 VPWR.n1340 0.120292
R13244 VPWR.n1356 VPWR.n1340 0.120292
R13245 VPWR.n1356 VPWR.n1355 0.120292
R13246 VPWR.n1355 VPWR.n1354 0.120292
R13247 VPWR.n1354 VPWR.n1342 0.120292
R13248 VPWR.n1348 VPWR.n1342 0.120292
R13249 VPWR.n1348 VPWR.n1347 0.120292
R13250 VPWR.n1410 VPWR.n1409 0.120292
R13251 VPWR.n1403 VPWR.n1402 0.120292
R13252 VPWR.n1402 VPWR.n1379 0.120292
R13253 VPWR.n1395 VPWR.n1379 0.120292
R13254 VPWR.n1395 VPWR.n1394 0.120292
R13255 VPWR.n1394 VPWR.n1393 0.120292
R13256 VPWR.n1393 VPWR.n1381 0.120292
R13257 VPWR.n1387 VPWR.n1381 0.120292
R13258 VPWR.n1387 VPWR.n1386 0.120292
R13259 VPWR.n1440 VPWR.n1439 0.120292
R13260 VPWR.n1439 VPWR.n1416 0.120292
R13261 VPWR.n1432 VPWR.n1416 0.120292
R13262 VPWR.n1432 VPWR.n1431 0.120292
R13263 VPWR.n1431 VPWR.n1430 0.120292
R13264 VPWR.n1430 VPWR.n1418 0.120292
R13265 VPWR.n1424 VPWR.n1418 0.120292
R13266 VPWR.n1424 VPWR.n1423 0.120292
R13267 VPWR.n2812 VPWR.n2798 0.120292
R13268 VPWR.n2796 VPWR.n2779 0.120292
R13269 VPWR.n2777 VPWR.n2759 0.120292
R13270 VPWR.n2757 VPWR.n2740 0.120292
R13271 VPWR.n2719 VPWR.n2718 0.120292
R13272 VPWR.n2720 VPWR.n2719 0.120292
R13273 VPWR.n2720 VPWR.n2711 0.120292
R13274 VPWR.n2725 VPWR.n2711 0.120292
R13275 VPWR.n2726 VPWR.n2725 0.120292
R13276 VPWR.n2726 VPWR.n2707 0.120292
R13277 VPWR.n2732 VPWR.n2707 0.120292
R13278 VPWR.n2734 VPWR.n2704 0.120292
R13279 VPWR.n2738 VPWR.n2704 0.120292
R13280 VPWR.n2683 VPWR.n2682 0.120292
R13281 VPWR.n2684 VPWR.n2683 0.120292
R13282 VPWR.n2684 VPWR.n2673 0.120292
R13283 VPWR.n2689 VPWR.n2673 0.120292
R13284 VPWR.n2690 VPWR.n2689 0.120292
R13285 VPWR.n2690 VPWR.n2669 0.120292
R13286 VPWR.n2695 VPWR.n2669 0.120292
R13287 VPWR.n2697 VPWR.n2666 0.120292
R13288 VPWR.n2702 VPWR.n2666 0.120292
R13289 VPWR.n2646 VPWR.n2645 0.120292
R13290 VPWR.n2647 VPWR.n2646 0.120292
R13291 VPWR.n2647 VPWR.n2636 0.120292
R13292 VPWR.n2652 VPWR.n2636 0.120292
R13293 VPWR.n2653 VPWR.n2652 0.120292
R13294 VPWR.n2653 VPWR.n2632 0.120292
R13295 VPWR.n2658 VPWR.n2632 0.120292
R13296 VPWR.n2660 VPWR.n2629 0.120292
R13297 VPWR.n2664 VPWR.n2629 0.120292
R13298 VPWR.n2608 VPWR.n2604 0.120292
R13299 VPWR.n2616 VPWR.n2604 0.120292
R13300 VPWR.n2617 VPWR.n2616 0.120292
R13301 VPWR.n2618 VPWR.n2617 0.120292
R13302 VPWR.n2618 VPWR.n2600 0.120292
R13303 VPWR.n2623 VPWR.n2600 0.120292
R13304 VPWR.n2624 VPWR.n2623 0.120292
R13305 VPWR.n1605 VPWR 0.118556
R13306 VPWR.n1108 VPWR 0.118556
R13307 VPWR.n1619 VPWR 0.118556
R13308 VPWR.n1632 VPWR 0.118556
R13309 VPWR.n1098 VPWR 0.118556
R13310 VPWR.n1646 VPWR 0.118556
R13311 VPWR.n1659 VPWR 0.118556
R13312 VPWR.n1088 VPWR 0.118556
R13313 VPWR.n1673 VPWR 0.118556
R13314 VPWR.n1686 VPWR 0.118556
R13315 VPWR.n1078 VPWR 0.118556
R13316 VPWR.n1700 VPWR 0.118556
R13317 VPWR.n1713 VPWR 0.118556
R13318 VPWR.n1725 VPWR 0.118556
R13319 VPWR VPWR.n1112 0.118556
R13320 VPWR.n1067 VPWR 0.118556
R13321 VPWR.n123 VPWR 0.118556
R13322 VPWR.n112 VPWR 0.118556
R13323 VPWR.n103 VPWR 0.118556
R13324 VPWR.n278 VPWR 0.118556
R13325 VPWR.n266 VPWR 0.118556
R13326 VPWR.n254 VPWR 0.118556
R13327 VPWR.n242 VPWR 0.118556
R13328 VPWR.n230 VPWR 0.118556
R13329 VPWR.n218 VPWR 0.118556
R13330 VPWR.n206 VPWR 0.118556
R13331 VPWR.n194 VPWR 0.118556
R13332 VPWR.n182 VPWR 0.118556
R13333 VPWR.n170 VPWR 0.118556
R13334 VPWR.n158 VPWR 0.118556
R13335 VPWR.n146 VPWR 0.118556
R13336 VPWR.n134 VPWR 0.118556
R13337 VPWR.n1765 VPWR.n1044 0.108238
R13338 VPWR.n1541 VPWR.n1143 0.108238
R13339 VPWR.n1540 VPWR.n1142 0.108238
R13340 VPWR.n1524 VPWR.n1141 0.108238
R13341 VPWR.n1516 VPWR.n1140 0.108238
R13342 VPWR.n1510 VPWR.n1139 0.108238
R13343 VPWR.n1502 VPWR.n1138 0.108238
R13344 VPWR.n1496 VPWR.n1137 0.108238
R13345 VPWR.n1583 VPWR.n1132 0.108238
R13346 VPWR.n1584 VPWR.n1131 0.108238
R13347 VPWR.n1463 VPWR.n1452 0.108238
R13348 VPWR.n1464 VPWR.n1451 0.108238
R13349 VPWR.n1795 VPWR.n1027 0.108238
R13350 VPWR.n1766 VPWR.n1043 0.108238
R13351 VPWR.n1744 VPWR.n1038 0.108238
R13352 VPWR.n1787 VPWR.n1786 0.108238
R13353 VPWR.n2481 VPWR 0.100405
R13354 VPWR.n2472 VPWR 0.100405
R13355 VPWR VPWR.n2385 0.100405
R13356 VPWR VPWR.n2386 0.100405
R13357 VPWR VPWR.n2387 0.100405
R13358 VPWR.n2305 VPWR 0.100405
R13359 VPWR VPWR.n2314 0.100405
R13360 VPWR.n2315 VPWR 0.100405
R13361 VPWR VPWR.n2324 0.100405
R13362 VPWR.n2375 VPWR 0.100405
R13363 VPWR VPWR.n2374 0.100405
R13364 VPWR.n2365 VPWR 0.100405
R13365 VPWR VPWR.n2364 0.100405
R13366 VPWR.n2355 VPWR 0.100405
R13367 VPWR VPWR.n2354 0.100405
R13368 VPWR.n2345 VPWR 0.100405
R13369 VPWR VPWR.n2344 0.100405
R13370 VPWR.n2335 VPWR 0.100405
R13371 VPWR VPWR.n2334 0.100405
R13372 VPWR.n2325 VPWR 0.100405
R13373 VPWR.n2302 VPWR 0.100405
R13374 VPWR.n2301 VPWR 0.100405
R13375 VPWR.n2300 VPWR 0.100405
R13376 VPWR.n2299 VPWR 0.100405
R13377 VPWR.n2288 VPWR 0.100405
R13378 VPWR.n2289 VPWR 0.100405
R13379 VPWR.n2290 VPWR 0.100405
R13380 VPWR.n2291 VPWR 0.100405
R13381 VPWR.n2292 VPWR 0.100405
R13382 VPWR.n2293 VPWR 0.100405
R13383 VPWR.n2294 VPWR 0.100405
R13384 VPWR.n2295 VPWR 0.100405
R13385 VPWR.n2296 VPWR 0.100405
R13386 VPWR.n2297 VPWR 0.100405
R13387 VPWR.n2298 VPWR 0.100405
R13388 VPWR.n2285 VPWR 0.100405
R13389 VPWR.n2276 VPWR 0.100405
R13390 VPWR.n2275 VPWR 0.100405
R13391 VPWR.n2266 VPWR 0.100405
R13392 VPWR.n2215 VPWR 0.100405
R13393 VPWR.n2216 VPWR 0.100405
R13394 VPWR.n2225 VPWR 0.100405
R13395 VPWR.n2226 VPWR 0.100405
R13396 VPWR.n2235 VPWR 0.100405
R13397 VPWR.n2236 VPWR 0.100405
R13398 VPWR.n2245 VPWR 0.100405
R13399 VPWR.n2246 VPWR 0.100405
R13400 VPWR.n2255 VPWR 0.100405
R13401 VPWR.n2256 VPWR 0.100405
R13402 VPWR.n2265 VPWR 0.100405
R13403 VPWR VPWR.n2189 0.100405
R13404 VPWR VPWR.n2190 0.100405
R13405 VPWR VPWR.n2191 0.100405
R13406 VPWR VPWR.n2192 0.100405
R13407 VPWR VPWR.n2203 0.100405
R13408 VPWR VPWR.n2202 0.100405
R13409 VPWR VPWR.n2201 0.100405
R13410 VPWR VPWR.n2200 0.100405
R13411 VPWR VPWR.n2199 0.100405
R13412 VPWR VPWR.n2198 0.100405
R13413 VPWR VPWR.n2197 0.100405
R13414 VPWR VPWR.n2196 0.100405
R13415 VPWR VPWR.n2195 0.100405
R13416 VPWR VPWR.n2194 0.100405
R13417 VPWR VPWR.n2193 0.100405
R13418 VPWR.n2109 VPWR 0.100405
R13419 VPWR VPWR.n2118 0.100405
R13420 VPWR.n2119 VPWR 0.100405
R13421 VPWR VPWR.n2128 0.100405
R13422 VPWR.n2179 VPWR 0.100405
R13423 VPWR VPWR.n2178 0.100405
R13424 VPWR.n2169 VPWR 0.100405
R13425 VPWR VPWR.n2168 0.100405
R13426 VPWR.n2159 VPWR 0.100405
R13427 VPWR VPWR.n2158 0.100405
R13428 VPWR.n2149 VPWR 0.100405
R13429 VPWR VPWR.n2148 0.100405
R13430 VPWR.n2139 VPWR 0.100405
R13431 VPWR VPWR.n2138 0.100405
R13432 VPWR.n2129 VPWR 0.100405
R13433 VPWR.n2106 VPWR 0.100405
R13434 VPWR.n2105 VPWR 0.100405
R13435 VPWR.n2104 VPWR 0.100405
R13436 VPWR.n2103 VPWR 0.100405
R13437 VPWR.n2092 VPWR 0.100405
R13438 VPWR.n2093 VPWR 0.100405
R13439 VPWR.n2094 VPWR 0.100405
R13440 VPWR.n2095 VPWR 0.100405
R13441 VPWR.n2096 VPWR 0.100405
R13442 VPWR.n2097 VPWR 0.100405
R13443 VPWR.n2098 VPWR 0.100405
R13444 VPWR.n2099 VPWR 0.100405
R13445 VPWR.n2100 VPWR 0.100405
R13446 VPWR.n2101 VPWR 0.100405
R13447 VPWR.n2102 VPWR 0.100405
R13448 VPWR.n2089 VPWR 0.100405
R13449 VPWR.n2080 VPWR 0.100405
R13450 VPWR.n2079 VPWR 0.100405
R13451 VPWR.n2070 VPWR 0.100405
R13452 VPWR.n2019 VPWR 0.100405
R13453 VPWR.n2020 VPWR 0.100405
R13454 VPWR.n2029 VPWR 0.100405
R13455 VPWR.n2030 VPWR 0.100405
R13456 VPWR.n2039 VPWR 0.100405
R13457 VPWR.n2040 VPWR 0.100405
R13458 VPWR.n2049 VPWR 0.100405
R13459 VPWR.n2050 VPWR 0.100405
R13460 VPWR.n2059 VPWR 0.100405
R13461 VPWR.n2060 VPWR 0.100405
R13462 VPWR.n2069 VPWR 0.100405
R13463 VPWR VPWR.n1993 0.100405
R13464 VPWR VPWR.n1994 0.100405
R13465 VPWR VPWR.n1995 0.100405
R13466 VPWR VPWR.n1996 0.100405
R13467 VPWR VPWR.n2007 0.100405
R13468 VPWR VPWR.n2006 0.100405
R13469 VPWR VPWR.n2005 0.100405
R13470 VPWR VPWR.n2004 0.100405
R13471 VPWR VPWR.n2003 0.100405
R13472 VPWR VPWR.n2002 0.100405
R13473 VPWR VPWR.n2001 0.100405
R13474 VPWR VPWR.n2000 0.100405
R13475 VPWR VPWR.n1999 0.100405
R13476 VPWR VPWR.n1998 0.100405
R13477 VPWR VPWR.n1997 0.100405
R13478 VPWR.n1913 VPWR 0.100405
R13479 VPWR VPWR.n1922 0.100405
R13480 VPWR.n1923 VPWR 0.100405
R13481 VPWR VPWR.n1932 0.100405
R13482 VPWR.n1983 VPWR 0.100405
R13483 VPWR VPWR.n1982 0.100405
R13484 VPWR.n1973 VPWR 0.100405
R13485 VPWR VPWR.n1972 0.100405
R13486 VPWR.n1963 VPWR 0.100405
R13487 VPWR VPWR.n1962 0.100405
R13488 VPWR.n1953 VPWR 0.100405
R13489 VPWR VPWR.n1952 0.100405
R13490 VPWR.n1943 VPWR 0.100405
R13491 VPWR VPWR.n1942 0.100405
R13492 VPWR.n1933 VPWR 0.100405
R13493 VPWR.n1910 VPWR 0.100405
R13494 VPWR.n1909 VPWR 0.100405
R13495 VPWR.n1908 VPWR 0.100405
R13496 VPWR.n1907 VPWR 0.100405
R13497 VPWR.n1896 VPWR 0.100405
R13498 VPWR.n1897 VPWR 0.100405
R13499 VPWR.n1898 VPWR 0.100405
R13500 VPWR.n1899 VPWR 0.100405
R13501 VPWR.n1900 VPWR 0.100405
R13502 VPWR.n1901 VPWR 0.100405
R13503 VPWR.n1902 VPWR 0.100405
R13504 VPWR.n1903 VPWR 0.100405
R13505 VPWR.n1904 VPWR 0.100405
R13506 VPWR.n1905 VPWR 0.100405
R13507 VPWR.n1906 VPWR 0.100405
R13508 VPWR VPWR.n2399 0.100405
R13509 VPWR VPWR.n2398 0.100405
R13510 VPWR VPWR.n2397 0.100405
R13511 VPWR VPWR.n2396 0.100405
R13512 VPWR VPWR.n2395 0.100405
R13513 VPWR VPWR.n2394 0.100405
R13514 VPWR VPWR.n2393 0.100405
R13515 VPWR VPWR.n2392 0.100405
R13516 VPWR VPWR.n2391 0.100405
R13517 VPWR VPWR.n2390 0.100405
R13518 VPWR VPWR.n2389 0.100405
R13519 VPWR VPWR.n2388 0.100405
R13520 VPWR.n1893 VPWR 0.100405
R13521 VPWR.n1884 VPWR 0.100405
R13522 VPWR.n1883 VPWR 0.100405
R13523 VPWR.n1874 VPWR 0.100405
R13524 VPWR.n1873 VPWR 0.100405
R13525 VPWR.n1823 VPWR 0.100405
R13526 VPWR.n1824 VPWR 0.100405
R13527 VPWR.n1833 VPWR 0.100405
R13528 VPWR.n1834 VPWR 0.100405
R13529 VPWR.n1843 VPWR 0.100405
R13530 VPWR.n1844 VPWR 0.100405
R13531 VPWR.n1853 VPWR 0.100405
R13532 VPWR.n1854 VPWR 0.100405
R13533 VPWR.n1863 VPWR 0.100405
R13534 VPWR.n1864 VPWR 0.100405
R13535 VPWR.n2411 VPWR 0.100405
R13536 VPWR.n2412 VPWR 0.100405
R13537 VPWR.n2421 VPWR 0.100405
R13538 VPWR.n2422 VPWR 0.100405
R13539 VPWR.n2431 VPWR 0.100405
R13540 VPWR.n2432 VPWR 0.100405
R13541 VPWR.n2441 VPWR 0.100405
R13542 VPWR.n2442 VPWR 0.100405
R13543 VPWR.n2451 VPWR 0.100405
R13544 VPWR.n2452 VPWR 0.100405
R13545 VPWR.n2461 VPWR 0.100405
R13546 VPWR.n2462 VPWR 0.100405
R13547 VPWR.n2471 VPWR 0.100405
R13548 VPWR VPWR.n1797 0.100405
R13549 VPWR VPWR.n1798 0.100405
R13550 VPWR VPWR.n1799 0.100405
R13551 VPWR VPWR.n1800 0.100405
R13552 VPWR VPWR.n1801 0.100405
R13553 VPWR VPWR.n1802 0.100405
R13554 VPWR VPWR.n1803 0.100405
R13555 VPWR VPWR.n1804 0.100405
R13556 VPWR VPWR.n1811 0.100405
R13557 VPWR VPWR.n1810 0.100405
R13558 VPWR VPWR.n1809 0.100405
R13559 VPWR VPWR.n1808 0.100405
R13560 VPWR VPWR.n1807 0.100405
R13561 VPWR VPWR.n1806 0.100405
R13562 VPWR VPWR.n1805 0.100405
R13563 VPWR.n2498 VPWR 0.100405
R13564 VPWR.n2497 VPWR 0.100405
R13565 VPWR.n2496 VPWR 0.100405
R13566 VPWR.n2495 VPWR 0.100405
R13567 VPWR.n2494 VPWR 0.100405
R13568 VPWR.n2493 VPWR 0.100405
R13569 VPWR.n2492 VPWR 0.100405
R13570 VPWR.n2491 VPWR 0.100405
R13571 VPWR.n2490 VPWR 0.100405
R13572 VPWR.n2489 VPWR 0.100405
R13573 VPWR.n2484 VPWR 0.100405
R13574 VPWR.n2485 VPWR 0.100405
R13575 VPWR.n2486 VPWR 0.100405
R13576 VPWR.n2487 VPWR 0.100405
R13577 VPWR.n2488 VPWR 0.100405
R13578 VPWR.n1143 VPWR 0.100405
R13579 VPWR VPWR.n1540 0.100405
R13580 VPWR.n1524 VPWR 0.100405
R13581 VPWR.n1516 VPWR 0.100405
R13582 VPWR.n1510 VPWR 0.100405
R13583 VPWR.n1502 VPWR 0.100405
R13584 VPWR.n1496 VPWR 0.100405
R13585 VPWR VPWR.n1132 0.100405
R13586 VPWR.n1584 VPWR 0.100405
R13587 VPWR.n1452 VPWR 0.100405
R13588 VPWR.n1464 VPWR 0.100405
R13589 VPWR.n1043 VPWR 0.100405
R13590 VPWR.n1744 VPWR 0.100405
R13591 VPWR.n1787 VPWR 0.100405
R13592 VPWR VPWR.n1765 0.100405
R13593 VPWR.n2501 VPWR 0.100405
R13594 VPWR VPWR.n2512 0.100405
R13595 VPWR.n2513 VPWR 0.100405
R13596 VPWR VPWR.n2524 0.100405
R13597 VPWR.n2525 VPWR 0.100405
R13598 VPWR VPWR.n2536 0.100405
R13599 VPWR.n2537 VPWR 0.100405
R13600 VPWR VPWR.n2548 0.100405
R13601 VPWR.n2549 VPWR 0.100405
R13602 VPWR VPWR.n2560 0.100405
R13603 VPWR.n2561 VPWR 0.100405
R13604 VPWR VPWR.n2572 0.100405
R13605 VPWR.n2573 VPWR 0.100405
R13606 VPWR VPWR.n2584 0.100405
R13607 VPWR.n2585 VPWR 0.100405
R13608 VPWR.n1056 VPWR 0.100405
R13609 VPWR.n1754 VPWR 0.100405
R13610 VPWR.n1755 VPWR 0.100405
R13611 VPWR.n1529 VPWR 0.100405
R13612 VPWR.n1530 VPWR 0.100405
R13613 VPWR VPWR.n1528 0.100405
R13614 VPWR VPWR.n1527 0.100405
R13615 VPWR.n1514 VPWR 0.100405
R13616 VPWR VPWR.n1513 0.100405
R13617 VPWR.n1500 VPWR 0.100405
R13618 VPWR VPWR.n1499 0.100405
R13619 VPWR.n1487 VPWR 0.100405
R13620 VPWR.n1587 VPWR 0.100405
R13621 VPWR.n1588 VPWR 0.100405
R13622 VPWR.n1448 VPWR 0.100405
R13623 VPWR VPWR.n2798 0.0994583
R13624 VPWR VPWR.n2779 0.0994583
R13625 VPWR VPWR.n1326 0.0981562
R13626 VPWR.n1371 VPWR 0.0981562
R13627 VPWR.n1410 VPWR 0.0981562
R13628 VPWR.n9 VPWR 0.0968542
R13629 VPWR.n1244 VPWR 0.0968542
R13630 VPWR.n1267 VPWR 0.0968542
R13631 VPWR.n1291 VPWR 0.0968542
R13632 VPWR.n1333 VPWR 0.0968542
R13633 VPWR VPWR.n2759 0.0968542
R13634 VPWR VPWR.n2740 0.0968542
R13635 VPWR.n2718 VPWR 0.0968542
R13636 VPWR.n2682 VPWR 0.0968542
R13637 VPWR.n2645 VPWR 0.0968542
R13638 VPWR.n2608 VPWR 0.0968542
R13639 VPWR VPWR.n1044 0.0945
R13640 VPWR.n1541 VPWR 0.0945
R13641 VPWR VPWR.n1142 0.0945
R13642 VPWR VPWR.n1141 0.0945
R13643 VPWR VPWR.n1140 0.0945
R13644 VPWR VPWR.n1139 0.0945
R13645 VPWR VPWR.n1138 0.0945
R13646 VPWR.n1137 VPWR 0.0945
R13647 VPWR VPWR.n1583 0.0945
R13648 VPWR VPWR.n1131 0.0945
R13649 VPWR VPWR.n1463 0.0945
R13650 VPWR.n1451 VPWR 0.0945
R13651 VPWR VPWR.n1038 0.0945
R13652 VPWR.n1786 VPWR 0.0945
R13653 VPWR VPWR.n1027 0.0945
R13654 VPWR.n1766 VPWR 0.0945
R13655 VPWR.n1117 VPWR 0.093504
R13656 VPWR.n109 VPWR 0.093504
R13657 VPWR.n143 VPWR 0.093504
R13658 VPWR.n155 VPWR 0.093504
R13659 VPWR.n167 VPWR 0.093504
R13660 VPWR.n179 VPWR 0.093504
R13661 VPWR.n191 VPWR 0.093504
R13662 VPWR.n203 VPWR 0.093504
R13663 VPWR.n215 VPWR 0.093504
R13664 VPWR.n227 VPWR 0.093504
R13665 VPWR.n239 VPWR 0.093504
R13666 VPWR.n251 VPWR 0.093504
R13667 VPWR.n263 VPWR 0.093504
R13668 VPWR.n275 VPWR 0.093504
R13669 VPWR VPWR.n285 0.093504
R13670 VPWR.n131 VPWR 0.093504
R13671 VPWR.n120 VPWR 0.093504
R13672 VPWR VPWR.n1731 0.093504
R13673 VPWR.n1722 VPWR 0.093504
R13674 VPWR.n1710 VPWR 0.093504
R13675 VPWR.n1699 VPWR 0.093504
R13676 VPWR VPWR.n1077 0.093504
R13677 VPWR.n1683 VPWR 0.093504
R13678 VPWR.n1672 VPWR 0.093504
R13679 VPWR VPWR.n1087 0.093504
R13680 VPWR.n1656 VPWR 0.093504
R13681 VPWR.n1645 VPWR 0.093504
R13682 VPWR VPWR.n1097 0.093504
R13683 VPWR.n1629 VPWR 0.093504
R13684 VPWR.n1618 VPWR 0.093504
R13685 VPWR VPWR.n1107 0.093504
R13686 VPWR.n1602 VPWR 0.093504
R13687 VPWR.n2598 VPWR 0.0849042
R13688 VPWR.n1112 VPWR.n1109 0.0845517
R13689 VPWR.n147 VPWR.n146 0.0845517
R13690 VPWR.n159 VPWR.n158 0.0845517
R13691 VPWR.n171 VPWR.n170 0.0845517
R13692 VPWR.n183 VPWR.n182 0.0845517
R13693 VPWR.n195 VPWR.n194 0.0845517
R13694 VPWR.n207 VPWR.n206 0.0845517
R13695 VPWR.n219 VPWR.n218 0.0845517
R13696 VPWR.n231 VPWR.n230 0.0845517
R13697 VPWR.n243 VPWR.n242 0.0845517
R13698 VPWR.n255 VPWR.n254 0.0845517
R13699 VPWR.n267 VPWR.n266 0.0845517
R13700 VPWR.n279 VPWR.n278 0.0845517
R13701 VPWR.n282 VPWR.n103 0.0845517
R13702 VPWR.n113 VPWR.n112 0.0845517
R13703 VPWR.n135 VPWR.n134 0.0845517
R13704 VPWR.n124 VPWR.n123 0.0845517
R13705 VPWR.n1728 VPWR.n1067 0.0845517
R13706 VPWR.n1726 VPWR.n1725 0.0845517
R13707 VPWR.n1714 VPWR.n1713 0.0845517
R13708 VPWR.n1701 VPWR.n1700 0.0845517
R13709 VPWR.n1690 VPWR.n1078 0.0845517
R13710 VPWR.n1687 VPWR.n1686 0.0845517
R13711 VPWR.n1674 VPWR.n1673 0.0845517
R13712 VPWR.n1663 VPWR.n1088 0.0845517
R13713 VPWR.n1660 VPWR.n1659 0.0845517
R13714 VPWR.n1647 VPWR.n1646 0.0845517
R13715 VPWR.n1636 VPWR.n1098 0.0845517
R13716 VPWR.n1633 VPWR.n1632 0.0845517
R13717 VPWR.n1620 VPWR.n1619 0.0845517
R13718 VPWR.n1609 VPWR.n1108 0.0845517
R13719 VPWR.n1606 VPWR.n1605 0.0845517
R13720 VPWR.n1456 VPWR.n1451 0.0740128
R13721 VPWR.n1542 VPWR.n1044 0.071
R13722 VPWR.n1547 VPWR.n1541 0.071
R13723 VPWR.n1552 VPWR.n1142 0.071
R13724 VPWR.n1557 VPWR.n1141 0.071
R13725 VPWR.n1562 VPWR.n1140 0.071
R13726 VPWR.n1567 VPWR.n1139 0.071
R13727 VPWR.n1572 VPWR.n1138 0.071
R13728 VPWR.n1577 VPWR.n1137 0.071
R13729 VPWR.n1583 VPWR.n1582 0.071
R13730 VPWR.n1457 VPWR.n1131 0.071
R13731 VPWR.n1463 VPWR.n1462 0.071
R13732 VPWR.n1772 VPWR.n1038 0.071
R13733 VPWR.n1786 VPWR.n1785 0.071
R13734 VPWR.n1780 VPWR.n1027 0.071
R13735 VPWR.n1767 VPWR.n1766 0.071
R13736 VPWR VPWR.n1115 0.0678077
R13737 VPWR VPWR.n107 0.0678077
R13738 VPWR VPWR.n141 0.0678077
R13739 VPWR VPWR.n153 0.0678077
R13740 VPWR VPWR.n165 0.0678077
R13741 VPWR VPWR.n177 0.0678077
R13742 VPWR VPWR.n189 0.0678077
R13743 VPWR VPWR.n201 0.0678077
R13744 VPWR VPWR.n213 0.0678077
R13745 VPWR VPWR.n225 0.0678077
R13746 VPWR VPWR.n237 0.0678077
R13747 VPWR VPWR.n249 0.0678077
R13748 VPWR VPWR.n261 0.0678077
R13749 VPWR VPWR.n273 0.0678077
R13750 VPWR.n286 VPWR 0.0678077
R13751 VPWR VPWR.n129 0.0678077
R13752 VPWR VPWR.n118 0.0678077
R13753 VPWR.n1732 VPWR 0.0678077
R13754 VPWR VPWR.n1720 0.0678077
R13755 VPWR VPWR.n1708 0.0678077
R13756 VPWR VPWR.n1697 0.0678077
R13757 VPWR.n1193 VPWR 0.0678077
R13758 VPWR VPWR.n1681 0.0678077
R13759 VPWR VPWR.n1670 0.0678077
R13760 VPWR.n1207 VPWR 0.0678077
R13761 VPWR VPWR.n1654 0.0678077
R13762 VPWR VPWR.n1643 0.0678077
R13763 VPWR.n1175 VPWR 0.0678077
R13764 VPWR VPWR.n1627 0.0678077
R13765 VPWR VPWR.n1616 0.0678077
R13766 VPWR.n1124 VPWR 0.0678077
R13767 VPWR VPWR.n1600 0.0678077
R13768 VPWR.n150 VPWR 0.063
R13769 VPWR.n162 VPWR 0.063
R13770 VPWR.n174 VPWR 0.063
R13771 VPWR.n186 VPWR 0.063
R13772 VPWR.n198 VPWR 0.063
R13773 VPWR.n210 VPWR 0.063
R13774 VPWR.n222 VPWR 0.063
R13775 VPWR.n234 VPWR 0.063
R13776 VPWR.n246 VPWR 0.063
R13777 VPWR.n258 VPWR 0.063
R13778 VPWR.n270 VPWR 0.063
R13779 VPWR.n101 VPWR 0.063
R13780 VPWR.n105 VPWR 0.063
R13781 VPWR.n138 VPWR 0.063
R13782 VPWR.n115 VPWR 0.063
R13783 VPWR.n126 VPWR 0.063
R13784 VPWR.n1065 VPWR 0.063
R13785 VPWR.n1717 VPWR 0.063
R13786 VPWR.n1070 VPWR 0.063
R13787 VPWR VPWR.n1704 0.063
R13788 VPWR VPWR.n1693 0.063
R13789 VPWR VPWR.n1081 0.063
R13790 VPWR VPWR.n1677 0.063
R13791 VPWR VPWR.n1666 0.063
R13792 VPWR VPWR.n1091 0.063
R13793 VPWR VPWR.n1650 0.063
R13794 VPWR VPWR.n1639 0.063
R13795 VPWR VPWR.n1101 0.063
R13796 VPWR VPWR.n1623 0.063
R13797 VPWR VPWR.n1612 0.063
R13798 VPWR VPWR.n1111 0.063
R13799 VPWR VPWR.n1120 0.063
R13800 VPWR.n1115 VPWR 0.0608448
R13801 VPWR.n107 VPWR 0.0608448
R13802 VPWR.n141 VPWR 0.0608448
R13803 VPWR.n153 VPWR 0.0608448
R13804 VPWR.n165 VPWR 0.0608448
R13805 VPWR.n177 VPWR 0.0608448
R13806 VPWR.n189 VPWR 0.0608448
R13807 VPWR.n201 VPWR 0.0608448
R13808 VPWR.n213 VPWR 0.0608448
R13809 VPWR.n225 VPWR 0.0608448
R13810 VPWR.n237 VPWR 0.0608448
R13811 VPWR.n249 VPWR 0.0608448
R13812 VPWR.n261 VPWR 0.0608448
R13813 VPWR.n273 VPWR 0.0608448
R13814 VPWR.n286 VPWR 0.0608448
R13815 VPWR.n129 VPWR 0.0608448
R13816 VPWR.n118 VPWR 0.0608448
R13817 VPWR.n1732 VPWR 0.0608448
R13818 VPWR.n1720 VPWR 0.0608448
R13819 VPWR.n1708 VPWR 0.0608448
R13820 VPWR.n1697 VPWR 0.0608448
R13821 VPWR.n1193 VPWR 0.0608448
R13822 VPWR.n1681 VPWR 0.0608448
R13823 VPWR.n1670 VPWR 0.0608448
R13824 VPWR.n1207 VPWR 0.0608448
R13825 VPWR.n1654 VPWR 0.0608448
R13826 VPWR.n1643 VPWR 0.0608448
R13827 VPWR.n1175 VPWR 0.0608448
R13828 VPWR.n1627 VPWR 0.0608448
R13829 VPWR.n1616 VPWR 0.0608448
R13830 VPWR.n1124 VPWR 0.0608448
R13831 VPWR.n1600 VPWR 0.0608448
R13832 VPWR VPWR.n13 0.0603958
R13833 VPWR VPWR.n12 0.0603958
R13834 VPWR VPWR.n1249 0.0603958
R13835 VPWR VPWR.n1248 0.0603958
R13836 VPWR VPWR.n1272 0.0603958
R13837 VPWR VPWR.n1271 0.0603958
R13838 VPWR VPWR.n1296 0.0603958
R13839 VPWR VPWR.n1295 0.0603958
R13840 VPWR.n1332 VPWR 0.0603958
R13841 VPWR VPWR.n1331 0.0603958
R13842 VPWR.n1327 VPWR 0.0603958
R13843 VPWR.n1318 VPWR 0.0603958
R13844 VPWR VPWR.n1317 0.0603958
R13845 VPWR.n1370 VPWR 0.0603958
R13846 VPWR VPWR.n1369 0.0603958
R13847 VPWR.n1364 VPWR 0.0603958
R13848 VPWR.n1409 VPWR 0.0603958
R13849 VPWR VPWR.n1408 0.0603958
R13850 VPWR.n1403 VPWR 0.0603958
R13851 VPWR.n1440 VPWR 0.0603958
R13852 VPWR VPWR.n2800 0.0603958
R13853 VPWR VPWR.n2799 0.0603958
R13854 VPWR VPWR.n2812 0.0603958
R13855 VPWR.n2791 VPWR 0.0603958
R13856 VPWR.n2792 VPWR 0.0603958
R13857 VPWR VPWR.n2796 0.0603958
R13858 VPWR.n2771 VPWR 0.0603958
R13859 VPWR.n2772 VPWR 0.0603958
R13860 VPWR VPWR.n2777 0.0603958
R13861 VPWR.n2752 VPWR 0.0603958
R13862 VPWR.n2753 VPWR 0.0603958
R13863 VPWR VPWR.n2757 0.0603958
R13864 VPWR.n2733 VPWR 0.0603958
R13865 VPWR.n2734 VPWR 0.0603958
R13866 VPWR VPWR.n2695 0.0603958
R13867 VPWR.n2696 VPWR 0.0603958
R13868 VPWR.n2697 VPWR 0.0603958
R13869 VPWR VPWR.n2658 0.0603958
R13870 VPWR.n2659 VPWR 0.0603958
R13871 VPWR.n2660 VPWR 0.0603958
R13872 VPWR.n2624 VPWR 0.0603958
R13873 VPWR.n2627 VPWR 0.0603958
R13874 VPWR.n1770 VPWR.n1769 0.0599512
R13875 VPWR.n1041 VPWR.n1040 0.0599512
R13876 VPWR.n1545 VPWR.n1544 0.0599512
R13877 VPWR.n1550 VPWR.n1549 0.0599512
R13878 VPWR.n1555 VPWR.n1554 0.0599512
R13879 VPWR.n1560 VPWR.n1559 0.0599512
R13880 VPWR.n1565 VPWR.n1564 0.0599512
R13881 VPWR.n1570 VPWR.n1569 0.0599512
R13882 VPWR.n1575 VPWR.n1574 0.0599512
R13883 VPWR.n1580 VPWR.n1579 0.0599512
R13884 VPWR.n1135 VPWR.n1134 0.0599512
R13885 VPWR.n1460 VPWR.n1459 0.0599512
R13886 VPWR.n1455 VPWR.n1454 0.0599512
R13887 VPWR.n1775 VPWR.n1774 0.0599512
R13888 VPWR.n1783 VPWR.n1782 0.0599512
R13889 VPWR.n1779 VPWR.n1778 0.0599512
R13890 VPWR.n1118 VPWR.n1117 0.0565345
R13891 VPWR.n1112 VPWR 0.0565345
R13892 VPWR.n144 VPWR.n143 0.0565345
R13893 VPWR.n146 VPWR 0.0565345
R13894 VPWR.n156 VPWR.n155 0.0565345
R13895 VPWR.n158 VPWR 0.0565345
R13896 VPWR.n168 VPWR.n167 0.0565345
R13897 VPWR.n170 VPWR 0.0565345
R13898 VPWR.n180 VPWR.n179 0.0565345
R13899 VPWR.n182 VPWR 0.0565345
R13900 VPWR.n192 VPWR.n191 0.0565345
R13901 VPWR.n194 VPWR 0.0565345
R13902 VPWR.n204 VPWR.n203 0.0565345
R13903 VPWR.n206 VPWR 0.0565345
R13904 VPWR.n216 VPWR.n215 0.0565345
R13905 VPWR.n218 VPWR 0.0565345
R13906 VPWR.n228 VPWR.n227 0.0565345
R13907 VPWR.n230 VPWR 0.0565345
R13908 VPWR.n240 VPWR.n239 0.0565345
R13909 VPWR.n242 VPWR 0.0565345
R13910 VPWR.n252 VPWR.n251 0.0565345
R13911 VPWR.n254 VPWR 0.0565345
R13912 VPWR.n264 VPWR.n263 0.0565345
R13913 VPWR.n266 VPWR 0.0565345
R13914 VPWR.n276 VPWR.n275 0.0565345
R13915 VPWR.n278 VPWR 0.0565345
R13916 VPWR.n285 VPWR.n283 0.0565345
R13917 VPWR.n103 VPWR 0.0565345
R13918 VPWR.n110 VPWR.n109 0.0565345
R13919 VPWR.n112 VPWR 0.0565345
R13920 VPWR.n132 VPWR.n131 0.0565345
R13921 VPWR.n134 VPWR 0.0565345
R13922 VPWR.n121 VPWR.n120 0.0565345
R13923 VPWR.n123 VPWR 0.0565345
R13924 VPWR.n1731 VPWR.n1729 0.0565345
R13925 VPWR.n1067 VPWR 0.0565345
R13926 VPWR.n1723 VPWR.n1722 0.0565345
R13927 VPWR.n1725 VPWR 0.0565345
R13928 VPWR.n1711 VPWR.n1710 0.0565345
R13929 VPWR.n1713 VPWR 0.0565345
R13930 VPWR.n1702 VPWR.n1699 0.0565345
R13931 VPWR.n1700 VPWR 0.0565345
R13932 VPWR.n1691 VPWR.n1077 0.0565345
R13933 VPWR.n1078 VPWR 0.0565345
R13934 VPWR.n1684 VPWR.n1683 0.0565345
R13935 VPWR.n1686 VPWR 0.0565345
R13936 VPWR.n1675 VPWR.n1672 0.0565345
R13937 VPWR.n1673 VPWR 0.0565345
R13938 VPWR.n1664 VPWR.n1087 0.0565345
R13939 VPWR.n1088 VPWR 0.0565345
R13940 VPWR.n1657 VPWR.n1656 0.0565345
R13941 VPWR.n1659 VPWR 0.0565345
R13942 VPWR.n1648 VPWR.n1645 0.0565345
R13943 VPWR.n1646 VPWR 0.0565345
R13944 VPWR.n1637 VPWR.n1097 0.0565345
R13945 VPWR.n1098 VPWR 0.0565345
R13946 VPWR.n1630 VPWR.n1629 0.0565345
R13947 VPWR.n1632 VPWR 0.0565345
R13948 VPWR.n1621 VPWR.n1618 0.0565345
R13949 VPWR.n1619 VPWR 0.0565345
R13950 VPWR.n1610 VPWR.n1107 0.0565345
R13951 VPWR.n1108 VPWR 0.0565345
R13952 VPWR.n1603 VPWR.n1602 0.0565345
R13953 VPWR.n1605 VPWR 0.0565345
R13954 VPWR.n1769 VPWR 0.0469286
R13955 VPWR.n1040 VPWR 0.0469286
R13956 VPWR.n1544 VPWR 0.0469286
R13957 VPWR.n1549 VPWR 0.0469286
R13958 VPWR.n1554 VPWR 0.0469286
R13959 VPWR.n1559 VPWR 0.0469286
R13960 VPWR.n1564 VPWR 0.0469286
R13961 VPWR.n1569 VPWR 0.0469286
R13962 VPWR.n1574 VPWR 0.0469286
R13963 VPWR.n1579 VPWR 0.0469286
R13964 VPWR.n1134 VPWR 0.0469286
R13965 VPWR.n1459 VPWR 0.0469286
R13966 VPWR.n1454 VPWR 0.0469286
R13967 VPWR.n1774 VPWR 0.0469286
R13968 VPWR.n1782 VPWR 0.0469286
R13969 VPWR.n1778 VPWR 0.0469286
R13970 VPWR.n1769 VPWR 0.0401341
R13971 VPWR.n1040 VPWR 0.0401341
R13972 VPWR.n1544 VPWR 0.0401341
R13973 VPWR.n1549 VPWR 0.0401341
R13974 VPWR.n1554 VPWR 0.0401341
R13975 VPWR.n1559 VPWR 0.0401341
R13976 VPWR.n1564 VPWR 0.0401341
R13977 VPWR.n1569 VPWR 0.0401341
R13978 VPWR.n1574 VPWR 0.0401341
R13979 VPWR.n1579 VPWR 0.0401341
R13980 VPWR.n1134 VPWR 0.0401341
R13981 VPWR.n1459 VPWR 0.0401341
R13982 VPWR.n1454 VPWR 0.0401341
R13983 VPWR.n1774 VPWR 0.0401341
R13984 VPWR.n1782 VPWR 0.0401341
R13985 VPWR.n1778 VPWR 0.0401341
R13986 VPWR.n13 VPWR 0.0382604
R13987 VPWR.n1249 VPWR 0.0382604
R13988 VPWR.n1272 VPWR 0.0382604
R13989 VPWR.n1296 VPWR 0.0382604
R13990 VPWR.n1331 VPWR 0.0382604
R13991 VPWR.n1369 VPWR 0.0382604
R13992 VPWR.n1408 VPWR 0.0382604
R13993 VPWR.n1445 VPWR 0.0382604
R13994 VPWR.n20 VPWR 0.0375125
R13995 VPWR.n20 VPWR 0.0373589
R13996 VPWR.n1118 VPWR.n1109 0.0349828
R13997 VPWR.n147 VPWR.n144 0.0349828
R13998 VPWR.n159 VPWR.n156 0.0349828
R13999 VPWR.n171 VPWR.n168 0.0349828
R14000 VPWR.n183 VPWR.n180 0.0349828
R14001 VPWR.n195 VPWR.n192 0.0349828
R14002 VPWR.n207 VPWR.n204 0.0349828
R14003 VPWR.n219 VPWR.n216 0.0349828
R14004 VPWR.n231 VPWR.n228 0.0349828
R14005 VPWR.n243 VPWR.n240 0.0349828
R14006 VPWR.n255 VPWR.n252 0.0349828
R14007 VPWR.n267 VPWR.n264 0.0349828
R14008 VPWR.n279 VPWR.n276 0.0349828
R14009 VPWR.n283 VPWR.n282 0.0349828
R14010 VPWR.n113 VPWR.n110 0.0349828
R14011 VPWR.n135 VPWR.n132 0.0349828
R14012 VPWR.n124 VPWR.n121 0.0349828
R14013 VPWR.n1729 VPWR.n1728 0.0349828
R14014 VPWR.n1726 VPWR.n1723 0.0349828
R14015 VPWR.n1714 VPWR.n1711 0.0349828
R14016 VPWR.n1702 VPWR.n1701 0.0349828
R14017 VPWR.n1691 VPWR.n1690 0.0349828
R14018 VPWR.n1687 VPWR.n1684 0.0349828
R14019 VPWR.n1675 VPWR.n1674 0.0349828
R14020 VPWR.n1664 VPWR.n1663 0.0349828
R14021 VPWR.n1660 VPWR.n1657 0.0349828
R14022 VPWR.n1648 VPWR.n1647 0.0349828
R14023 VPWR.n1637 VPWR.n1636 0.0349828
R14024 VPWR.n1633 VPWR.n1630 0.0349828
R14025 VPWR.n1621 VPWR.n1620 0.0349828
R14026 VPWR.n1610 VPWR.n1609 0.0349828
R14027 VPWR.n1606 VPWR.n1603 0.0349828
R14028 VPWR.n2504 VPWR.n2503 0.0340366
R14029 VPWR.n2570 VPWR.n2569 0.0340366
R14030 VPWR.n2510 VPWR.n2509 0.0340366
R14031 VPWR.n2552 VPWR.n2551 0.0340366
R14032 VPWR.n2546 VPWR.n2545 0.0340366
R14033 VPWR.n2534 VPWR.n2533 0.0340366
R14034 VPWR.n2528 VPWR.n2527 0.0340366
R14035 VPWR.n1223 VPWR.n1222 0.0340366
R14036 VPWR.n2522 VPWR.n2521 0.0340366
R14037 VPWR.n1486 VPWR.n1102 0.0340366
R14038 VPWR.n1174 VPWR.n1094 0.0340366
R14039 VPWR.n2540 VPWR.n2539 0.0340366
R14040 VPWR.n1165 VPWR.n1092 0.0340366
R14041 VPWR.n1211 VPWR.n1164 0.0340366
R14042 VPWR.n2516 VPWR.n2515 0.0340366
R14043 VPWR.n1129 VPWR.n1104 0.0340366
R14044 VPWR.n1155 VPWR.n1084 0.0340366
R14045 VPWR.n2558 VPWR.n2557 0.0340366
R14046 VPWR.n1144 VPWR.n1082 0.0340366
R14047 VPWR.n1591 VPWR.n1590 0.0340366
R14048 VPWR.n2564 VPWR.n2563 0.0340366
R14049 VPWR.n1197 VPWR.n1154 0.0340366
R14050 VPWR.n1074 VPWR.n1073 0.0340366
R14051 VPWR.n1743 VPWR.n1742 0.0340366
R14052 VPWR.n1071 VPWR.n1054 0.0340366
R14053 VPWR.n2576 VPWR.n2575 0.0340366
R14054 VPWR.n2582 VPWR.n2581 0.0340366
R14055 VPWR.n2593 VPWR.n2592 0.0340366
R14056 VPWR.n2588 VPWR.n2587 0.0340366
R14057 VPWR.n1737 VPWR.n1736 0.0340366
R14058 VPWR.n1063 VPWR.n1060 0.0340366
R14059 VPWR.n1596 VPWR.n1121 0.0340366
R14060 VPWR.n2628 VPWR.n2598 0.0320292
R14061 VPWR.n2800 VPWR 0.03175
R14062 VPWR VPWR.n2791 0.03175
R14063 VPWR VPWR.n2771 0.03175
R14064 VPWR VPWR.n2752 0.03175
R14065 VPWR VPWR.n2733 0.03175
R14066 VPWR VPWR.n2696 0.03175
R14067 VPWR VPWR.n2659 0.03175
R14068 VPWR VPWR.n2627 0.03175
R14069 VPWR.n2598 VPWR.n2597 0.0240975
R14070 VPWR.n2597 VPWR.n20 0.0240975
R14071 VPWR.n2814 VPWR 0.024
R14072 VPWR.n14 VPWR 0.0239375
R14073 VPWR.n12 VPWR 0.0239375
R14074 VPWR.n1250 VPWR 0.0239375
R14075 VPWR.n1248 VPWR 0.0239375
R14076 VPWR.n1271 VPWR 0.0239375
R14077 VPWR.n1295 VPWR 0.0239375
R14078 VPWR.n2753 VPWR 0.0239375
R14079 VPWR.n2503 VPWR 0.0233659
R14080 VPWR.n1466 VPWR 0.0233659
R14081 VPWR.n352 VPWR 0.0233659
R14082 VPWR.n2570 VPWR 0.0233659
R14083 VPWR.n1533 VPWR 0.0233659
R14084 VPWR.n347 VPWR 0.0233659
R14085 VPWR.n2510 VPWR 0.0233659
R14086 VPWR.n964 VPWR 0.0233659
R14087 VPWR.n2479 VPWR 0.0233659
R14088 VPWR.n2474 VPWR 0.0233659
R14089 VPWR.n319 VPWR 0.0233659
R14090 VPWR.n2551 VPWR 0.0233659
R14091 VPWR.n972 VPWR 0.0233659
R14092 VPWR.n2444 VPWR 0.0233659
R14093 VPWR.n323 VPWR 0.0233659
R14094 VPWR.n2546 VPWR 0.0233659
R14095 VPWR.n1891 VPWR 0.0233659
R14096 VPWR.n1886 VPWR 0.0233659
R14097 VPWR.n1881 VPWR 0.0233659
R14098 VPWR.n388 VPWR 0.0233659
R14099 VPWR.n392 VPWR 0.0233659
R14100 VPWR.n396 VPWR 0.0233659
R14101 VPWR.n2454 VPWR 0.0233659
R14102 VPWR.n331 VPWR 0.0233659
R14103 VPWR.n2534 VPWR 0.0233659
R14104 VPWR.n1876 VPWR 0.0233659
R14105 VPWR.n404 VPWR 0.0233659
R14106 VPWR.n2459 VPWR 0.0233659
R14107 VPWR.n335 VPWR 0.0233659
R14108 VPWR.n2527 VPWR 0.0233659
R14109 VPWR.n2307 VPWR 0.0233659
R14110 VPWR.n2312 VPWR 0.0233659
R14111 VPWR.n2317 VPWR 0.0233659
R14112 VPWR.n2322 VPWR 0.0233659
R14113 VPWR.n2332 VPWR 0.0233659
R14114 VPWR.n2337 VPWR 0.0233659
R14115 VPWR.n2342 VPWR 0.0233659
R14116 VPWR.n2347 VPWR 0.0233659
R14117 VPWR.n2352 VPWR 0.0233659
R14118 VPWR.n2357 VPWR 0.0233659
R14119 VPWR.n2362 VPWR 0.0233659
R14120 VPWR.n2367 VPWR 0.0233659
R14121 VPWR.n2372 VPWR 0.0233659
R14122 VPWR.n2377 VPWR 0.0233659
R14123 VPWR.n2381 VPWR 0.0233659
R14124 VPWR.n2327 VPWR 0.0233659
R14125 VPWR.n544 VPWR 0.0233659
R14126 VPWR.n539 VPWR 0.0233659
R14127 VPWR.n535 VPWR 0.0233659
R14128 VPWR.n531 VPWR 0.0233659
R14129 VPWR.n523 VPWR 0.0233659
R14130 VPWR.n519 VPWR 0.0233659
R14131 VPWR.n515 VPWR 0.0233659
R14132 VPWR.n511 VPWR 0.0233659
R14133 VPWR.n507 VPWR 0.0233659
R14134 VPWR.n503 VPWR 0.0233659
R14135 VPWR.n499 VPWR 0.0233659
R14136 VPWR.n495 VPWR 0.0233659
R14137 VPWR.n491 VPWR 0.0233659
R14138 VPWR.n487 VPWR 0.0233659
R14139 VPWR.n484 VPWR 0.0233659
R14140 VPWR.n527 VPWR 0.0233659
R14141 VPWR.n2283 VPWR 0.0233659
R14142 VPWR.n2278 VPWR 0.0233659
R14143 VPWR.n2273 VPWR 0.0233659
R14144 VPWR.n2268 VPWR 0.0233659
R14145 VPWR.n2258 VPWR 0.0233659
R14146 VPWR.n2253 VPWR 0.0233659
R14147 VPWR.n2248 VPWR 0.0233659
R14148 VPWR.n2243 VPWR 0.0233659
R14149 VPWR.n2238 VPWR 0.0233659
R14150 VPWR.n2233 VPWR 0.0233659
R14151 VPWR.n2228 VPWR 0.0233659
R14152 VPWR.n2223 VPWR 0.0233659
R14153 VPWR.n2218 VPWR 0.0233659
R14154 VPWR.n2213 VPWR 0.0233659
R14155 VPWR.n2209 VPWR 0.0233659
R14156 VPWR.n2263 VPWR 0.0233659
R14157 VPWR.n580 VPWR 0.0233659
R14158 VPWR.n584 VPWR 0.0233659
R14159 VPWR.n588 VPWR 0.0233659
R14160 VPWR.n592 VPWR 0.0233659
R14161 VPWR.n600 VPWR 0.0233659
R14162 VPWR.n604 VPWR 0.0233659
R14163 VPWR.n608 VPWR 0.0233659
R14164 VPWR.n612 VPWR 0.0233659
R14165 VPWR.n616 VPWR 0.0233659
R14166 VPWR.n620 VPWR 0.0233659
R14167 VPWR.n624 VPWR 0.0233659
R14168 VPWR.n628 VPWR 0.0233659
R14169 VPWR.n632 VPWR 0.0233659
R14170 VPWR.n636 VPWR 0.0233659
R14171 VPWR.n640 VPWR 0.0233659
R14172 VPWR.n596 VPWR 0.0233659
R14173 VPWR.n2111 VPWR 0.0233659
R14174 VPWR.n2116 VPWR 0.0233659
R14175 VPWR.n2121 VPWR 0.0233659
R14176 VPWR.n2126 VPWR 0.0233659
R14177 VPWR.n2136 VPWR 0.0233659
R14178 VPWR.n2141 VPWR 0.0233659
R14179 VPWR.n2146 VPWR 0.0233659
R14180 VPWR.n2151 VPWR 0.0233659
R14181 VPWR.n2156 VPWR 0.0233659
R14182 VPWR.n2161 VPWR 0.0233659
R14183 VPWR.n2166 VPWR 0.0233659
R14184 VPWR.n2171 VPWR 0.0233659
R14185 VPWR.n2176 VPWR 0.0233659
R14186 VPWR.n2181 VPWR 0.0233659
R14187 VPWR.n2185 VPWR 0.0233659
R14188 VPWR.n2131 VPWR 0.0233659
R14189 VPWR.n736 VPWR 0.0233659
R14190 VPWR.n731 VPWR 0.0233659
R14191 VPWR.n727 VPWR 0.0233659
R14192 VPWR.n723 VPWR 0.0233659
R14193 VPWR.n715 VPWR 0.0233659
R14194 VPWR.n711 VPWR 0.0233659
R14195 VPWR.n707 VPWR 0.0233659
R14196 VPWR.n703 VPWR 0.0233659
R14197 VPWR.n699 VPWR 0.0233659
R14198 VPWR.n695 VPWR 0.0233659
R14199 VPWR.n691 VPWR 0.0233659
R14200 VPWR.n687 VPWR 0.0233659
R14201 VPWR.n683 VPWR 0.0233659
R14202 VPWR.n679 VPWR 0.0233659
R14203 VPWR.n676 VPWR 0.0233659
R14204 VPWR.n719 VPWR 0.0233659
R14205 VPWR.n2087 VPWR 0.0233659
R14206 VPWR.n2082 VPWR 0.0233659
R14207 VPWR.n2077 VPWR 0.0233659
R14208 VPWR.n2072 VPWR 0.0233659
R14209 VPWR.n2062 VPWR 0.0233659
R14210 VPWR.n2057 VPWR 0.0233659
R14211 VPWR.n2052 VPWR 0.0233659
R14212 VPWR.n2047 VPWR 0.0233659
R14213 VPWR.n2042 VPWR 0.0233659
R14214 VPWR.n2037 VPWR 0.0233659
R14215 VPWR.n2032 VPWR 0.0233659
R14216 VPWR.n2027 VPWR 0.0233659
R14217 VPWR.n2022 VPWR 0.0233659
R14218 VPWR.n2017 VPWR 0.0233659
R14219 VPWR.n2013 VPWR 0.0233659
R14220 VPWR.n2067 VPWR 0.0233659
R14221 VPWR.n772 VPWR 0.0233659
R14222 VPWR.n776 VPWR 0.0233659
R14223 VPWR.n780 VPWR 0.0233659
R14224 VPWR.n784 VPWR 0.0233659
R14225 VPWR.n792 VPWR 0.0233659
R14226 VPWR.n796 VPWR 0.0233659
R14227 VPWR.n800 VPWR 0.0233659
R14228 VPWR.n804 VPWR 0.0233659
R14229 VPWR.n808 VPWR 0.0233659
R14230 VPWR.n812 VPWR 0.0233659
R14231 VPWR.n816 VPWR 0.0233659
R14232 VPWR.n820 VPWR 0.0233659
R14233 VPWR.n824 VPWR 0.0233659
R14234 VPWR.n828 VPWR 0.0233659
R14235 VPWR.n832 VPWR 0.0233659
R14236 VPWR.n788 VPWR 0.0233659
R14237 VPWR.n1915 VPWR 0.0233659
R14238 VPWR.n1920 VPWR 0.0233659
R14239 VPWR.n1925 VPWR 0.0233659
R14240 VPWR.n1930 VPWR 0.0233659
R14241 VPWR.n1940 VPWR 0.0233659
R14242 VPWR.n1945 VPWR 0.0233659
R14243 VPWR.n1950 VPWR 0.0233659
R14244 VPWR.n1955 VPWR 0.0233659
R14245 VPWR.n1960 VPWR 0.0233659
R14246 VPWR.n1965 VPWR 0.0233659
R14247 VPWR.n1970 VPWR 0.0233659
R14248 VPWR.n1975 VPWR 0.0233659
R14249 VPWR.n1980 VPWR 0.0233659
R14250 VPWR.n1985 VPWR 0.0233659
R14251 VPWR.n1989 VPWR 0.0233659
R14252 VPWR.n1935 VPWR 0.0233659
R14253 VPWR.n928 VPWR 0.0233659
R14254 VPWR.n923 VPWR 0.0233659
R14255 VPWR.n919 VPWR 0.0233659
R14256 VPWR.n915 VPWR 0.0233659
R14257 VPWR.n907 VPWR 0.0233659
R14258 VPWR.n903 VPWR 0.0233659
R14259 VPWR.n899 VPWR 0.0233659
R14260 VPWR.n895 VPWR 0.0233659
R14261 VPWR.n891 VPWR 0.0233659
R14262 VPWR.n887 VPWR 0.0233659
R14263 VPWR.n883 VPWR 0.0233659
R14264 VPWR.n879 VPWR 0.0233659
R14265 VPWR.n875 VPWR 0.0233659
R14266 VPWR.n871 VPWR 0.0233659
R14267 VPWR.n868 VPWR 0.0233659
R14268 VPWR.n911 VPWR 0.0233659
R14269 VPWR.n1871 VPWR 0.0233659
R14270 VPWR.n980 VPWR 0.0233659
R14271 VPWR.n1495 VPWR 0.0233659
R14272 VPWR.n1223 VPWR 0.0233659
R14273 VPWR.n400 VPWR 0.0233659
R14274 VPWR.n2464 VPWR 0.0233659
R14275 VPWR.n339 VPWR 0.0233659
R14276 VPWR.n2522 VPWR 0.0233659
R14277 VPWR.n976 VPWR 0.0233659
R14278 VPWR.n1490 VPWR 0.0233659
R14279 VPWR.n1486 VPWR 0.0233659
R14280 VPWR.n1866 VPWR 0.0233659
R14281 VPWR.n984 VPWR 0.0233659
R14282 VPWR.n1504 VPWR 0.0233659
R14283 VPWR.n1174 VPWR 0.0233659
R14284 VPWR.n408 VPWR 0.0233659
R14285 VPWR.n416 VPWR 0.0233659
R14286 VPWR.n420 VPWR 0.0233659
R14287 VPWR.n424 VPWR 0.0233659
R14288 VPWR.n428 VPWR 0.0233659
R14289 VPWR.n432 VPWR 0.0233659
R14290 VPWR.n436 VPWR 0.0233659
R14291 VPWR.n440 VPWR 0.0233659
R14292 VPWR.n444 VPWR 0.0233659
R14293 VPWR.n448 VPWR 0.0233659
R14294 VPWR.n412 VPWR 0.0233659
R14295 VPWR.n2449 VPWR 0.0233659
R14296 VPWR.n327 VPWR 0.0233659
R14297 VPWR.n2539 VPWR 0.0233659
R14298 VPWR.n988 VPWR 0.0233659
R14299 VPWR.n1509 VPWR 0.0233659
R14300 VPWR.n1165 VPWR 0.0233659
R14301 VPWR.n1861 VPWR 0.0233659
R14302 VPWR.n1851 VPWR 0.0233659
R14303 VPWR.n1846 VPWR 0.0233659
R14304 VPWR.n1841 VPWR 0.0233659
R14305 VPWR.n1836 VPWR 0.0233659
R14306 VPWR.n1831 VPWR 0.0233659
R14307 VPWR.n1826 VPWR 0.0233659
R14308 VPWR.n1821 VPWR 0.0233659
R14309 VPWR.n1817 VPWR 0.0233659
R14310 VPWR.n1856 VPWR 0.0233659
R14311 VPWR.n992 VPWR 0.0233659
R14312 VPWR.n1518 VPWR 0.0233659
R14313 VPWR.n1164 VPWR 0.0233659
R14314 VPWR.n2469 VPWR 0.0233659
R14315 VPWR.n343 VPWR 0.0233659
R14316 VPWR.n2515 VPWR 0.0233659
R14317 VPWR.n1130 VPWR 0.0233659
R14318 VPWR.n1129 VPWR 0.0233659
R14319 VPWR.n996 VPWR 0.0233659
R14320 VPWR.n1523 VPWR 0.0233659
R14321 VPWR.n1155 VPWR 0.0233659
R14322 VPWR.n2439 VPWR 0.0233659
R14323 VPWR.n2429 VPWR 0.0233659
R14324 VPWR.n2424 VPWR 0.0233659
R14325 VPWR.n2419 VPWR 0.0233659
R14326 VPWR.n2414 VPWR 0.0233659
R14327 VPWR.n2409 VPWR 0.0233659
R14328 VPWR.n2405 VPWR 0.0233659
R14329 VPWR.n2434 VPWR 0.0233659
R14330 VPWR.n315 VPWR 0.0233659
R14331 VPWR.n2558 VPWR 0.0233659
R14332 VPWR.n1538 VPWR 0.0233659
R14333 VPWR.n1144 VPWR 0.0233659
R14334 VPWR.n1000 VPWR 0.0233659
R14335 VPWR.n1004 VPWR 0.0233659
R14336 VPWR.n1008 VPWR 0.0233659
R14337 VPWR.n1012 VPWR 0.0233659
R14338 VPWR.n1016 VPWR 0.0233659
R14339 VPWR.n1020 VPWR 0.0233659
R14340 VPWR.n1024 VPWR 0.0233659
R14341 VPWR.n968 VPWR 0.0233659
R14342 VPWR.n1473 VPWR 0.0233659
R14343 VPWR.n1590 VPWR 0.0233659
R14344 VPWR.n311 VPWR 0.0233659
R14345 VPWR.n2563 VPWR 0.0233659
R14346 VPWR.n1154 VPWR 0.0233659
R14347 VPWR.n1763 VPWR 0.0233659
R14348 VPWR.n1073 VPWR 0.0233659
R14349 VPWR.n307 VPWR 0.0233659
R14350 VPWR.n303 VPWR 0.0233659
R14351 VPWR.n295 VPWR 0.0233659
R14352 VPWR.n292 VPWR 0.0233659
R14353 VPWR.n299 VPWR 0.0233659
R14354 VPWR.n1743 VPWR 0.0233659
R14355 VPWR.n1751 VPWR 0.0233659
R14356 VPWR.n1789 VPWR 0.0233659
R14357 VPWR.n1793 VPWR 0.0233659
R14358 VPWR.n1758 VPWR 0.0233659
R14359 VPWR.n1054 VPWR 0.0233659
R14360 VPWR.n2575 VPWR 0.0233659
R14361 VPWR.n2582 VPWR 0.0233659
R14362 VPWR.n2593 VPWR 0.0233659
R14363 VPWR.n2587 VPWR 0.0233659
R14364 VPWR.n1736 VPWR 0.0233659
R14365 VPWR.n1060 VPWR 0.0233659
R14366 VPWR.n1121 VPWR 0.0233659
R14367 VPWR.n1336 VPWR 0.0226354
R14368 VPWR.n1327 VPWR 0.0226354
R14369 VPWR.n1413 VPWR 0.0226354
R14370 VPWR.n2772 VPWR 0.0226354
R14371 VPWR VPWR.n2732 0.0226354
R14372 VPWR VPWR.n2702 0.0226354
R14373 VPWR VPWR.n2664 0.0226354
R14374 VPWR VPWR.n64 0.0220517
R14375 VPWR VPWR.n67 0.0220517
R14376 VPWR VPWR.n70 0.0220517
R14377 VPWR VPWR.n73 0.0220517
R14378 VPWR VPWR.n76 0.0220517
R14379 VPWR VPWR.n79 0.0220517
R14380 VPWR VPWR.n82 0.0220517
R14381 VPWR VPWR.n85 0.0220517
R14382 VPWR VPWR.n88 0.0220517
R14383 VPWR VPWR.n91 0.0220517
R14384 VPWR VPWR.n94 0.0220517
R14385 VPWR VPWR.n97 0.0220517
R14386 VPWR.n289 VPWR 0.0220517
R14387 VPWR VPWR.n61 0.0220517
R14388 VPWR VPWR.n58 0.0220517
R14389 VPWR.n1735 VPWR 0.0220517
R14390 VPWR VPWR.n1057 0.0220517
R14391 VPWR.n1705 VPWR 0.0220517
R14392 VPWR.n1694 VPWR 0.0220517
R14393 VPWR.n1196 VPWR 0.0220517
R14394 VPWR.n1678 VPWR 0.0220517
R14395 VPWR.n1667 VPWR 0.0220517
R14396 VPWR.n1210 VPWR 0.0220517
R14397 VPWR.n1651 VPWR 0.0220517
R14398 VPWR.n1640 VPWR 0.0220517
R14399 VPWR.n1178 VPWR 0.0220517
R14400 VPWR.n1624 VPWR 0.0220517
R14401 VPWR.n1613 VPWR 0.0220517
R14402 VPWR.n1127 VPWR 0.0220517
R14403 VPWR.n1597 VPWR 0.0220517
R14404 VPWR.n1273 VPWR 0.0213333
R14405 VPWR.n1297 VPWR 0.0213333
R14406 VPWR.n1311 VPWR 0.0213333
R14407 VPWR.n1375 VPWR 0.0213333
R14408 VPWR.n1347 VPWR 0.0213333
R14409 VPWR.n1386 VPWR 0.0213333
R14410 VPWR.n1423 VPWR 0.0213333
R14411 VPWR.n2806 VPWR 0.0213333
R14412 VPWR.n2799 VPWR 0.0213333
R14413 VPWR VPWR.n2790 0.0213333
R14414 VPWR.n2792 VPWR 0.0213333
R14415 VPWR VPWR.n2770 0.0213333
R14416 VPWR VPWR.n2751 0.0213333
R14417 VPWR VPWR.n2738 0.0213333
R14418 VPWR.n2500 VPWR 0.0196917
R14419 VPWR.n24 VPWR 0.0143889
R14420 VPWR VPWR.n19 0.0099
R14421 VPWR VPWR.n1604 0.00397222
R14422 VPWR VPWR.n1105 0.00397222
R14423 VPWR VPWR.n1103 0.00397222
R14424 VPWR VPWR.n1631 0.00397222
R14425 VPWR VPWR.n1095 0.00397222
R14426 VPWR VPWR.n1093 0.00397222
R14427 VPWR VPWR.n1658 0.00397222
R14428 VPWR VPWR.n1085 0.00397222
R14429 VPWR VPWR.n1083 0.00397222
R14430 VPWR VPWR.n1685 0.00397222
R14431 VPWR VPWR.n1075 0.00397222
R14432 VPWR VPWR.n1072 0.00397222
R14433 VPWR VPWR.n1712 0.00397222
R14434 VPWR VPWR.n1724 0.00397222
R14435 VPWR.n1113 VPWR 0.00397222
R14436 VPWR VPWR.n1066 0.00397222
R14437 VPWR VPWR.n122 0.00397222
R14438 VPWR VPWR.n111 0.00397222
R14439 VPWR VPWR.n102 0.00397222
R14440 VPWR VPWR.n277 0.00397222
R14441 VPWR VPWR.n265 0.00397222
R14442 VPWR VPWR.n253 0.00397222
R14443 VPWR VPWR.n241 0.00397222
R14444 VPWR VPWR.n229 0.00397222
R14445 VPWR VPWR.n217 0.00397222
R14446 VPWR VPWR.n205 0.00397222
R14447 VPWR VPWR.n193 0.00397222
R14448 VPWR VPWR.n181 0.00397222
R14449 VPWR VPWR.n169 0.00397222
R14450 VPWR VPWR.n157 0.00397222
R14451 VPWR VPWR.n145 0.00397222
R14452 VPWR VPWR.n133 0.00397222
R14453 VPWR.n1462 VPWR.n1461 0.00351282
R14454 VPWR.n1457 VPWR.n1136 0.00351282
R14455 VPWR.n1582 VPWR.n1581 0.00351282
R14456 VPWR.n1577 VPWR.n1576 0.00351282
R14457 VPWR.n1572 VPWR.n1571 0.00351282
R14458 VPWR.n1567 VPWR.n1566 0.00351282
R14459 VPWR.n1562 VPWR.n1561 0.00351282
R14460 VPWR.n1557 VPWR.n1556 0.00351282
R14461 VPWR.n1552 VPWR.n1551 0.00351282
R14462 VPWR.n1547 VPWR.n1546 0.00351282
R14463 VPWR.n1542 VPWR.n1042 0.00351282
R14464 VPWR.n1785 VPWR.n1784 0.00351282
R14465 VPWR.n1776 VPWR.n1772 0.00351282
R14466 VPWR.n1771 VPWR.n1767 0.00351282
R14467 VPWR.n141 VPWR.n140 0.00265517
R14468 VPWR.n153 VPWR.n152 0.00265517
R14469 VPWR.n165 VPWR.n164 0.00265517
R14470 VPWR.n177 VPWR.n176 0.00265517
R14471 VPWR.n189 VPWR.n188 0.00265517
R14472 VPWR.n201 VPWR.n200 0.00265517
R14473 VPWR.n213 VPWR.n212 0.00265517
R14474 VPWR.n225 VPWR.n224 0.00265517
R14475 VPWR.n237 VPWR.n236 0.00265517
R14476 VPWR.n249 VPWR.n248 0.00265517
R14477 VPWR.n261 VPWR.n260 0.00265517
R14478 VPWR.n273 VPWR.n272 0.00265517
R14479 VPWR.n288 VPWR.n286 0.00265517
R14480 VPWR.n129 VPWR.n128 0.00265517
R14481 VPWR.n118 VPWR.n117 0.00265517
R14482 VPWR.n1734 VPWR.n1732 0.00265517
R14483 VPWR.n1720 VPWR.n1719 0.00265517
R14484 VPWR.n1708 VPWR.n1707 0.00265517
R14485 VPWR.n1697 VPWR.n1696 0.00265517
R14486 VPWR.n1195 VPWR.n1193 0.00265517
R14487 VPWR.n1681 VPWR.n1680 0.00265517
R14488 VPWR.n1670 VPWR.n1669 0.00265517
R14489 VPWR.n1209 VPWR.n1207 0.00265517
R14490 VPWR.n1654 VPWR.n1653 0.00265517
R14491 VPWR.n1643 VPWR.n1642 0.00265517
R14492 VPWR.n1177 VPWR.n1175 0.00265517
R14493 VPWR.n1627 VPWR.n1626 0.00265517
R14494 VPWR.n1616 VPWR.n1615 0.00265517
R14495 VPWR.n1126 VPWR.n1124 0.00265517
R14496 VPWR.n1600 VPWR.n1599 0.00265517
R14497 Iout.n1020 Iout.t222 239.927
R14498 Iout.n509 Iout.t138 239.927
R14499 Iout.n513 Iout.t4 239.927
R14500 Iout.n507 Iout.t76 239.927
R14501 Iout.n504 Iout.t246 239.927
R14502 Iout.n500 Iout.t98 239.927
R14503 Iout.n192 Iout.t175 239.927
R14504 Iout.n195 Iout.t234 239.927
R14505 Iout.n199 Iout.t143 239.927
R14506 Iout.n202 Iout.t75 239.927
R14507 Iout.n206 Iout.t187 239.927
R14508 Iout.n210 Iout.t44 239.927
R14509 Iout.n214 Iout.t6 239.927
R14510 Iout.n218 Iout.t52 239.927
R14511 Iout.n222 Iout.t115 239.927
R14512 Iout.n226 Iout.t116 239.927
R14513 Iout.n232 Iout.t199 239.927
R14514 Iout.n235 Iout.t196 239.927
R14515 Iout.n238 Iout.t89 239.927
R14516 Iout.n241 Iout.t88 239.927
R14517 Iout.n244 Iout.t254 239.927
R14518 Iout.n247 Iout.t20 239.927
R14519 Iout.n250 Iout.t19 239.927
R14520 Iout.n255 Iout.t5 239.927
R14521 Iout.n252 Iout.t72 239.927
R14522 Iout.n489 Iout.t30 239.927
R14523 Iout.n494 Iout.t207 239.927
R14524 Iout.n491 Iout.t91 239.927
R14525 Iout.n519 Iout.t27 239.927
R14526 Iout.n149 Iout.t102 239.927
R14527 Iout.n146 Iout.t217 239.927
R14528 Iout.n1010 Iout.t105 239.927
R14529 Iout.n1007 Iout.t67 239.927
R14530 Iout.n140 Iout.t253 239.927
R14531 Iout.n143 Iout.t9 239.927
R14532 Iout.n525 Iout.t112 239.927
R14533 Iout.n480 Iout.t156 239.927
R14534 Iout.n483 Iout.t57 239.927
R14535 Iout.n478 Iout.t247 239.927
R14536 Iout.n259 Iout.t169 239.927
R14537 Iout.n186 Iout.t51 239.927
R14538 Iout.n271 Iout.t93 239.927
R14539 Iout.n180 Iout.t84 239.927
R14540 Iout.n283 Iout.t3 239.927
R14541 Iout.n174 Iout.t188 239.927
R14542 Iout.n168 Iout.t251 239.927
R14543 Iout.n301 Iout.t55 239.927
R14544 Iout.n289 Iout.t165 239.927
R14545 Iout.n177 Iout.t129 239.927
R14546 Iout.n277 Iout.t62 239.927
R14547 Iout.n183 Iout.t14 239.927
R14548 Iout.n265 Iout.t41 239.927
R14549 Iout.n189 Iout.t18 239.927
R14550 Iout.n472 Iout.t221 239.927
R14551 Iout.n469 Iout.t153 239.927
R14552 Iout.n156 Iout.t94 239.927
R14553 Iout.n531 Iout.t50 239.927
R14554 Iout.n534 Iout.t46 239.927
R14555 Iout.n536 Iout.t140 239.927
R14556 Iout.n133 Iout.t47 239.927
R14557 Iout.n136 Iout.t230 239.927
R14558 Iout.n542 Iout.t209 239.927
R14559 Iout.n460 Iout.t177 239.927
R14560 Iout.n463 Iout.t232 239.927
R14561 Iout.n458 Iout.t126 239.927
R14562 Iout.n305 Iout.t121 239.927
R14563 Iout.n308 Iout.t136 239.927
R14564 Iout.n311 Iout.t168 239.927
R14565 Iout.n314 Iout.t239 239.927
R14566 Iout.n317 Iout.t109 239.927
R14567 Iout.n320 Iout.t139 239.927
R14568 Iout.n392 Iout.t111 239.927
R14569 Iout.n378 Iout.t235 239.927
R14570 Iout.n376 Iout.t43 239.927
R14571 Iout.n394 Iout.t154 239.927
R14572 Iout.n408 Iout.t8 239.927
R14573 Iout.n410 Iout.t180 239.927
R14574 Iout.n424 Iout.t206 239.927
R14575 Iout.n426 Iout.t203 239.927
R14576 Iout.n447 Iout.t218 239.927
R14577 Iout.n452 Iout.t65 239.927
R14578 Iout.n449 Iout.t63 239.927
R14579 Iout.n548 Iout.t242 239.927
R14580 Iout.n130 Iout.t210 239.927
R14581 Iout.n559 Iout.t220 239.927
R14582 Iout.n557 Iout.t119 239.927
R14583 Iout.n554 Iout.t53 239.927
R14584 Iout.n434 Iout.t189 239.927
R14585 Iout.n438 Iout.t233 239.927
R14586 Iout.n441 Iout.t176 239.927
R14587 Iout.n432 Iout.t164 239.927
R14588 Iout.n418 Iout.t70 239.927
R14589 Iout.n416 Iout.t45 239.927
R14590 Iout.n402 Iout.t7 239.927
R14591 Iout.n357 Iout.t192 239.927
R14592 Iout.n360 Iout.t110 239.927
R14593 Iout.n363 Iout.t229 239.927
R14594 Iout.n366 Iout.t90 239.927
R14595 Iout.n354 Iout.t131 239.927
R14596 Iout.n351 Iout.t78 239.927
R14597 Iout.n348 Iout.t191 239.927
R14598 Iout.n345 Iout.t123 239.927
R14599 Iout.n342 Iout.t194 239.927
R14600 Iout.n339 Iout.t157 239.927
R14601 Iout.n336 Iout.t117 239.927
R14602 Iout.n333 Iout.t227 239.927
R14603 Iout.n117 Iout.t82 239.927
R14604 Iout.n582 Iout.t181 239.927
R14605 Iout.n111 Iout.t122 239.927
R14606 Iout.n594 Iout.t127 239.927
R14607 Iout.n105 Iout.t104 239.927
R14608 Iout.n606 Iout.t147 239.927
R14609 Iout.n99 Iout.t141 239.927
R14610 Iout.n618 Iout.t99 239.927
R14611 Iout.n624 Iout.t255 239.927
R14612 Iout.n90 Iout.t215 239.927
R14613 Iout.n636 Iout.t64 239.927
R14614 Iout.n81 Iout.t118 239.927
R14615 Iout.n648 Iout.t34 239.927
R14616 Iout.n96 Iout.t74 239.927
R14617 Iout.n612 Iout.t173 239.927
R14618 Iout.n102 Iout.t149 239.927
R14619 Iout.n600 Iout.t172 239.927
R14620 Iout.n108 Iout.t29 239.927
R14621 Iout.n588 Iout.t40 239.927
R14622 Iout.n687 Iout.t36 239.927
R14623 Iout.n684 Iout.t10 239.927
R14624 Iout.n681 Iout.t15 239.927
R14625 Iout.n678 Iout.t213 239.927
R14626 Iout.n675 Iout.t151 239.927
R14627 Iout.n672 Iout.t160 239.927
R14628 Iout.n747 Iout.t66 239.927
R14629 Iout.n50 Iout.t77 239.927
R14630 Iout.n759 Iout.t33 239.927
R14631 Iout.n44 Iout.t241 239.927
R14632 Iout.n771 Iout.t219 239.927
R14633 Iout.n42 Iout.t103 239.927
R14634 Iout.n56 Iout.t39 239.927
R14635 Iout.n735 Iout.t48 239.927
R14636 Iout.n62 Iout.t240 239.927
R14637 Iout.n723 Iout.t13 239.927
R14638 Iout.n717 Iout.t132 239.927
R14639 Iout.n65 Iout.t202 239.927
R14640 Iout.n729 Iout.t204 239.927
R14641 Iout.n59 Iout.t101 239.927
R14642 Iout.n805 Iout.t183 239.927
R14643 Iout.n808 Iout.t195 239.927
R14644 Iout.n811 Iout.t162 239.927
R14645 Iout.n814 Iout.t73 239.927
R14646 Iout.n817 Iout.t49 239.927
R14647 Iout.n820 Iout.t69 239.927
R14648 Iout.n823 Iout.t174 239.927
R14649 Iout.n802 Iout.t26 239.927
R14650 Iout.n799 Iout.t100 239.927
R14651 Iout.n890 Iout.t225 239.927
R14652 Iout.n888 Iout.t243 239.927
R14653 Iout.n881 Iout.t238 239.927
R14654 Iout.n869 Iout.t35 239.927
R14655 Iout.n867 Iout.t252 239.927
R14656 Iout.n855 Iout.t158 239.927
R14657 Iout.n853 Iout.t135 239.927
R14658 Iout.n841 Iout.t197 239.927
R14659 Iout.n839 Iout.t128 239.927
R14660 Iout.n827 Iout.t182 239.927
R14661 Iout.n883 Iout.t2 239.927
R14662 Iout.n895 Iout.t216 239.927
R14663 Iout.n897 Iout.t113 239.927
R14664 Iout.n909 Iout.t244 239.927
R14665 Iout.n911 Iout.t68 239.927
R14666 Iout.n923 Iout.t80 239.927
R14667 Iout.n926 Iout.t124 239.927
R14668 Iout.n22 Iout.t223 239.927
R14669 Iout.n876 Iout.t108 239.927
R14670 Iout.n874 Iout.t249 239.927
R14671 Iout.n862 Iout.t107 239.927
R14672 Iout.n860 Iout.t31 239.927
R14673 Iout.n848 Iout.t166 239.927
R14674 Iout.n846 Iout.t96 239.927
R14675 Iout.n834 Iout.t60 239.927
R14676 Iout.n832 Iout.t205 239.927
R14677 Iout.n902 Iout.t86 239.927
R14678 Iout.n904 Iout.t148 239.927
R14679 Iout.n916 Iout.t167 239.927
R14680 Iout.n918 Iout.t12 239.927
R14681 Iout.n931 Iout.t1 239.927
R14682 Iout.n934 Iout.t17 239.927
R14683 Iout.n796 Iout.t155 239.927
R14684 Iout.n793 Iout.t231 239.927
R14685 Iout.n790 Iout.t146 239.927
R14686 Iout.n787 Iout.t245 239.927
R14687 Iout.n784 Iout.t142 239.927
R14688 Iout.n781 Iout.t228 239.927
R14689 Iout.n938 Iout.t79 239.927
R14690 Iout.n741 Iout.t114 239.927
R14691 Iout.n53 Iout.t159 239.927
R14692 Iout.n753 Iout.t184 239.927
R14693 Iout.n47 Iout.t185 239.927
R14694 Iout.n765 Iout.t71 239.927
R14695 Iout.n38 Iout.t61 239.927
R14696 Iout.n777 Iout.t201 239.927
R14697 Iout.n71 Iout.t59 239.927
R14698 Iout.n705 Iout.t190 239.927
R14699 Iout.n77 Iout.t171 239.927
R14700 Iout.n944 Iout.t54 239.927
R14701 Iout.n19 Iout.t56 239.927
R14702 Iout.n68 Iout.t250 239.927
R14703 Iout.n711 Iout.t161 239.927
R14704 Iout.n74 Iout.t32 239.927
R14705 Iout.n699 Iout.t226 239.927
R14706 Iout.n950 Iout.t198 239.927
R14707 Iout.n953 Iout.t224 239.927
R14708 Iout.n669 Iout.t214 239.927
R14709 Iout.n666 Iout.t83 239.927
R14710 Iout.n663 Iout.t23 239.927
R14711 Iout.n660 Iout.t95 239.927
R14712 Iout.n657 Iout.t87 239.927
R14713 Iout.n654 Iout.t211 239.927
R14714 Iout.n690 Iout.t25 239.927
R14715 Iout.n695 Iout.t163 239.927
R14716 Iout.n692 Iout.t179 239.927
R14717 Iout.n957 Iout.t42 239.927
R14718 Iout.n114 Iout.t130 239.927
R14719 Iout.n576 Iout.t193 239.927
R14720 Iout.n573 Iout.t16 239.927
R14721 Iout.n963 Iout.t97 239.927
R14722 Iout.n14 Iout.t11 239.927
R14723 Iout.n93 Iout.t134 239.927
R14724 Iout.n630 Iout.t248 239.927
R14725 Iout.n87 Iout.t208 239.927
R14726 Iout.n642 Iout.t237 239.927
R14727 Iout.n85 Iout.t81 239.927
R14728 Iout.n563 Iout.t92 239.927
R14729 Iout.n969 Iout.t236 239.927
R14730 Iout.n972 Iout.t145 239.927
R14731 Iout.n569 Iout.t24 239.927
R14732 Iout.n123 Iout.t150 239.927
R14733 Iout.n120 Iout.t0 239.927
R14734 Iout.n976 Iout.t106 239.927
R14735 Iout.n400 Iout.t120 239.927
R14736 Iout.n386 Iout.t38 239.927
R14737 Iout.n384 Iout.t178 239.927
R14738 Iout.n370 Iout.t28 239.927
R14739 Iout.n982 Iout.t137 239.927
R14740 Iout.n9 Iout.t170 239.927
R14741 Iout.n127 Iout.t152 239.927
R14742 Iout.n988 Iout.t85 239.927
R14743 Iout.n991 Iout.t125 239.927
R14744 Iout.n323 Iout.t200 239.927
R14745 Iout.n326 Iout.t133 239.927
R14746 Iout.n329 Iout.t22 239.927
R14747 Iout.n995 Iout.t21 239.927
R14748 Iout.n1001 Iout.t186 239.927
R14749 Iout.n4 Iout.t144 239.927
R14750 Iout.n295 Iout.t58 239.927
R14751 Iout.n172 Iout.t212 239.927
R14752 Iout.n1014 Iout.t37 239.927
R14753 Iout.n1021 Iout.n1020 7.9105
R14754 Iout.n510 Iout.n509 7.9105
R14755 Iout.n514 Iout.n513 7.9105
R14756 Iout.n508 Iout.n507 7.9105
R14757 Iout.n505 Iout.n504 7.9105
R14758 Iout.n501 Iout.n500 7.9105
R14759 Iout.n193 Iout.n192 7.9105
R14760 Iout.n196 Iout.n195 7.9105
R14761 Iout.n200 Iout.n199 7.9105
R14762 Iout.n203 Iout.n202 7.9105
R14763 Iout.n207 Iout.n206 7.9105
R14764 Iout.n211 Iout.n210 7.9105
R14765 Iout.n215 Iout.n214 7.9105
R14766 Iout.n219 Iout.n218 7.9105
R14767 Iout.n223 Iout.n222 7.9105
R14768 Iout.n227 Iout.n226 7.9105
R14769 Iout.n233 Iout.n232 7.9105
R14770 Iout.n236 Iout.n235 7.9105
R14771 Iout.n239 Iout.n238 7.9105
R14772 Iout.n242 Iout.n241 7.9105
R14773 Iout.n245 Iout.n244 7.9105
R14774 Iout.n248 Iout.n247 7.9105
R14775 Iout.n251 Iout.n250 7.9105
R14776 Iout.n256 Iout.n255 7.9105
R14777 Iout.n253 Iout.n252 7.9105
R14778 Iout.n490 Iout.n489 7.9105
R14779 Iout.n495 Iout.n494 7.9105
R14780 Iout.n492 Iout.n491 7.9105
R14781 Iout.n520 Iout.n519 7.9105
R14782 Iout.n150 Iout.n149 7.9105
R14783 Iout.n147 Iout.n146 7.9105
R14784 Iout.n1011 Iout.n1010 7.9105
R14785 Iout.n1008 Iout.n1007 7.9105
R14786 Iout.n141 Iout.n140 7.9105
R14787 Iout.n144 Iout.n143 7.9105
R14788 Iout.n526 Iout.n525 7.9105
R14789 Iout.n481 Iout.n480 7.9105
R14790 Iout.n484 Iout.n483 7.9105
R14791 Iout.n479 Iout.n478 7.9105
R14792 Iout.n260 Iout.n259 7.9105
R14793 Iout.n187 Iout.n186 7.9105
R14794 Iout.n272 Iout.n271 7.9105
R14795 Iout.n181 Iout.n180 7.9105
R14796 Iout.n284 Iout.n283 7.9105
R14797 Iout.n175 Iout.n174 7.9105
R14798 Iout.n169 Iout.n168 7.9105
R14799 Iout.n302 Iout.n301 7.9105
R14800 Iout.n290 Iout.n289 7.9105
R14801 Iout.n178 Iout.n177 7.9105
R14802 Iout.n278 Iout.n277 7.9105
R14803 Iout.n184 Iout.n183 7.9105
R14804 Iout.n266 Iout.n265 7.9105
R14805 Iout.n190 Iout.n189 7.9105
R14806 Iout.n473 Iout.n472 7.9105
R14807 Iout.n470 Iout.n469 7.9105
R14808 Iout.n157 Iout.n156 7.9105
R14809 Iout.n532 Iout.n531 7.9105
R14810 Iout.n535 Iout.n534 7.9105
R14811 Iout.n537 Iout.n536 7.9105
R14812 Iout.n134 Iout.n133 7.9105
R14813 Iout.n137 Iout.n136 7.9105
R14814 Iout.n543 Iout.n542 7.9105
R14815 Iout.n461 Iout.n460 7.9105
R14816 Iout.n464 Iout.n463 7.9105
R14817 Iout.n459 Iout.n458 7.9105
R14818 Iout.n306 Iout.n305 7.9105
R14819 Iout.n309 Iout.n308 7.9105
R14820 Iout.n312 Iout.n311 7.9105
R14821 Iout.n315 Iout.n314 7.9105
R14822 Iout.n318 Iout.n317 7.9105
R14823 Iout.n321 Iout.n320 7.9105
R14824 Iout.n393 Iout.n392 7.9105
R14825 Iout.n379 Iout.n378 7.9105
R14826 Iout.n377 Iout.n376 7.9105
R14827 Iout.n395 Iout.n394 7.9105
R14828 Iout.n409 Iout.n408 7.9105
R14829 Iout.n411 Iout.n410 7.9105
R14830 Iout.n425 Iout.n424 7.9105
R14831 Iout.n427 Iout.n426 7.9105
R14832 Iout.n448 Iout.n447 7.9105
R14833 Iout.n453 Iout.n452 7.9105
R14834 Iout.n450 Iout.n449 7.9105
R14835 Iout.n549 Iout.n548 7.9105
R14836 Iout.n131 Iout.n130 7.9105
R14837 Iout.n560 Iout.n559 7.9105
R14838 Iout.n558 Iout.n557 7.9105
R14839 Iout.n555 Iout.n554 7.9105
R14840 Iout.n435 Iout.n434 7.9105
R14841 Iout.n439 Iout.n438 7.9105
R14842 Iout.n442 Iout.n441 7.9105
R14843 Iout.n433 Iout.n432 7.9105
R14844 Iout.n419 Iout.n418 7.9105
R14845 Iout.n417 Iout.n416 7.9105
R14846 Iout.n403 Iout.n402 7.9105
R14847 Iout.n358 Iout.n357 7.9105
R14848 Iout.n361 Iout.n360 7.9105
R14849 Iout.n364 Iout.n363 7.9105
R14850 Iout.n367 Iout.n366 7.9105
R14851 Iout.n355 Iout.n354 7.9105
R14852 Iout.n352 Iout.n351 7.9105
R14853 Iout.n349 Iout.n348 7.9105
R14854 Iout.n346 Iout.n345 7.9105
R14855 Iout.n343 Iout.n342 7.9105
R14856 Iout.n340 Iout.n339 7.9105
R14857 Iout.n337 Iout.n336 7.9105
R14858 Iout.n334 Iout.n333 7.9105
R14859 Iout.n118 Iout.n117 7.9105
R14860 Iout.n583 Iout.n582 7.9105
R14861 Iout.n112 Iout.n111 7.9105
R14862 Iout.n595 Iout.n594 7.9105
R14863 Iout.n106 Iout.n105 7.9105
R14864 Iout.n607 Iout.n606 7.9105
R14865 Iout.n100 Iout.n99 7.9105
R14866 Iout.n619 Iout.n618 7.9105
R14867 Iout.n625 Iout.n624 7.9105
R14868 Iout.n91 Iout.n90 7.9105
R14869 Iout.n637 Iout.n636 7.9105
R14870 Iout.n82 Iout.n81 7.9105
R14871 Iout.n649 Iout.n648 7.9105
R14872 Iout.n97 Iout.n96 7.9105
R14873 Iout.n613 Iout.n612 7.9105
R14874 Iout.n103 Iout.n102 7.9105
R14875 Iout.n601 Iout.n600 7.9105
R14876 Iout.n109 Iout.n108 7.9105
R14877 Iout.n589 Iout.n588 7.9105
R14878 Iout.n688 Iout.n687 7.9105
R14879 Iout.n685 Iout.n684 7.9105
R14880 Iout.n682 Iout.n681 7.9105
R14881 Iout.n679 Iout.n678 7.9105
R14882 Iout.n676 Iout.n675 7.9105
R14883 Iout.n673 Iout.n672 7.9105
R14884 Iout.n748 Iout.n747 7.9105
R14885 Iout.n51 Iout.n50 7.9105
R14886 Iout.n760 Iout.n759 7.9105
R14887 Iout.n45 Iout.n44 7.9105
R14888 Iout.n772 Iout.n771 7.9105
R14889 Iout.n43 Iout.n42 7.9105
R14890 Iout.n57 Iout.n56 7.9105
R14891 Iout.n736 Iout.n735 7.9105
R14892 Iout.n63 Iout.n62 7.9105
R14893 Iout.n724 Iout.n723 7.9105
R14894 Iout.n718 Iout.n717 7.9105
R14895 Iout.n66 Iout.n65 7.9105
R14896 Iout.n730 Iout.n729 7.9105
R14897 Iout.n60 Iout.n59 7.9105
R14898 Iout.n806 Iout.n805 7.9105
R14899 Iout.n809 Iout.n808 7.9105
R14900 Iout.n812 Iout.n811 7.9105
R14901 Iout.n815 Iout.n814 7.9105
R14902 Iout.n818 Iout.n817 7.9105
R14903 Iout.n821 Iout.n820 7.9105
R14904 Iout.n824 Iout.n823 7.9105
R14905 Iout.n803 Iout.n802 7.9105
R14906 Iout.n800 Iout.n799 7.9105
R14907 Iout.n891 Iout.n890 7.9105
R14908 Iout.n889 Iout.n888 7.9105
R14909 Iout.n882 Iout.n881 7.9105
R14910 Iout.n870 Iout.n869 7.9105
R14911 Iout.n868 Iout.n867 7.9105
R14912 Iout.n856 Iout.n855 7.9105
R14913 Iout.n854 Iout.n853 7.9105
R14914 Iout.n842 Iout.n841 7.9105
R14915 Iout.n840 Iout.n839 7.9105
R14916 Iout.n828 Iout.n827 7.9105
R14917 Iout.n884 Iout.n883 7.9105
R14918 Iout.n896 Iout.n895 7.9105
R14919 Iout.n898 Iout.n897 7.9105
R14920 Iout.n910 Iout.n909 7.9105
R14921 Iout.n912 Iout.n911 7.9105
R14922 Iout.n924 Iout.n923 7.9105
R14923 Iout.n927 Iout.n926 7.9105
R14924 Iout.n23 Iout.n22 7.9105
R14925 Iout.n877 Iout.n876 7.9105
R14926 Iout.n875 Iout.n874 7.9105
R14927 Iout.n863 Iout.n862 7.9105
R14928 Iout.n861 Iout.n860 7.9105
R14929 Iout.n849 Iout.n848 7.9105
R14930 Iout.n847 Iout.n846 7.9105
R14931 Iout.n835 Iout.n834 7.9105
R14932 Iout.n833 Iout.n832 7.9105
R14933 Iout.n903 Iout.n902 7.9105
R14934 Iout.n905 Iout.n904 7.9105
R14935 Iout.n917 Iout.n916 7.9105
R14936 Iout.n919 Iout.n918 7.9105
R14937 Iout.n932 Iout.n931 7.9105
R14938 Iout.n935 Iout.n934 7.9105
R14939 Iout.n797 Iout.n796 7.9105
R14940 Iout.n794 Iout.n793 7.9105
R14941 Iout.n791 Iout.n790 7.9105
R14942 Iout.n788 Iout.n787 7.9105
R14943 Iout.n785 Iout.n784 7.9105
R14944 Iout.n782 Iout.n781 7.9105
R14945 Iout.n939 Iout.n938 7.9105
R14946 Iout.n742 Iout.n741 7.9105
R14947 Iout.n54 Iout.n53 7.9105
R14948 Iout.n754 Iout.n753 7.9105
R14949 Iout.n48 Iout.n47 7.9105
R14950 Iout.n766 Iout.n765 7.9105
R14951 Iout.n39 Iout.n38 7.9105
R14952 Iout.n778 Iout.n777 7.9105
R14953 Iout.n72 Iout.n71 7.9105
R14954 Iout.n706 Iout.n705 7.9105
R14955 Iout.n78 Iout.n77 7.9105
R14956 Iout.n945 Iout.n944 7.9105
R14957 Iout.n20 Iout.n19 7.9105
R14958 Iout.n69 Iout.n68 7.9105
R14959 Iout.n712 Iout.n711 7.9105
R14960 Iout.n75 Iout.n74 7.9105
R14961 Iout.n700 Iout.n699 7.9105
R14962 Iout.n951 Iout.n950 7.9105
R14963 Iout.n954 Iout.n953 7.9105
R14964 Iout.n670 Iout.n669 7.9105
R14965 Iout.n667 Iout.n666 7.9105
R14966 Iout.n664 Iout.n663 7.9105
R14967 Iout.n661 Iout.n660 7.9105
R14968 Iout.n658 Iout.n657 7.9105
R14969 Iout.n655 Iout.n654 7.9105
R14970 Iout.n691 Iout.n690 7.9105
R14971 Iout.n696 Iout.n695 7.9105
R14972 Iout.n693 Iout.n692 7.9105
R14973 Iout.n958 Iout.n957 7.9105
R14974 Iout.n115 Iout.n114 7.9105
R14975 Iout.n577 Iout.n576 7.9105
R14976 Iout.n574 Iout.n573 7.9105
R14977 Iout.n964 Iout.n963 7.9105
R14978 Iout.n15 Iout.n14 7.9105
R14979 Iout.n94 Iout.n93 7.9105
R14980 Iout.n631 Iout.n630 7.9105
R14981 Iout.n88 Iout.n87 7.9105
R14982 Iout.n643 Iout.n642 7.9105
R14983 Iout.n86 Iout.n85 7.9105
R14984 Iout.n564 Iout.n563 7.9105
R14985 Iout.n970 Iout.n969 7.9105
R14986 Iout.n973 Iout.n972 7.9105
R14987 Iout.n570 Iout.n569 7.9105
R14988 Iout.n124 Iout.n123 7.9105
R14989 Iout.n121 Iout.n120 7.9105
R14990 Iout.n977 Iout.n976 7.9105
R14991 Iout.n401 Iout.n400 7.9105
R14992 Iout.n387 Iout.n386 7.9105
R14993 Iout.n385 Iout.n384 7.9105
R14994 Iout.n371 Iout.n370 7.9105
R14995 Iout.n983 Iout.n982 7.9105
R14996 Iout.n10 Iout.n9 7.9105
R14997 Iout.n128 Iout.n127 7.9105
R14998 Iout.n989 Iout.n988 7.9105
R14999 Iout.n992 Iout.n991 7.9105
R15000 Iout.n324 Iout.n323 7.9105
R15001 Iout.n327 Iout.n326 7.9105
R15002 Iout.n330 Iout.n329 7.9105
R15003 Iout.n996 Iout.n995 7.9105
R15004 Iout.n1002 Iout.n1001 7.9105
R15005 Iout.n5 Iout.n4 7.9105
R15006 Iout.n296 Iout.n295 7.9105
R15007 Iout.n173 Iout.n172 7.9105
R15008 Iout.n1015 Iout.n1014 7.9105
R15009 Iout.n886 Iout.n885 3.86101
R15010 Iout.n880 Iout.n879 3.86101
R15011 Iout.n894 Iout.n893 3.86101
R15012 Iout.n872 Iout.n871 3.86101
R15013 Iout.n900 Iout.n899 3.86101
R15014 Iout.n866 Iout.n865 3.86101
R15015 Iout.n908 Iout.n907 3.86101
R15016 Iout.n858 Iout.n857 3.86101
R15017 Iout.n914 Iout.n913 3.86101
R15018 Iout.n852 Iout.n851 3.86101
R15019 Iout.n922 Iout.n921 3.86101
R15020 Iout.n844 Iout.n843 3.86101
R15021 Iout.n929 Iout.n928 3.86101
R15022 Iout.n838 Iout.n837 3.86101
R15023 Iout.n925 Iout.n21 3.86101
R15024 Iout.n830 Iout.n829 3.86101
R15025 Iout.n879 Iout.n878 3.4105
R15026 Iout.n887 Iout.n886 3.4105
R15027 Iout.n893 Iout.n892 3.4105
R15028 Iout.n798 Iout.n28 3.4105
R15029 Iout.n801 Iout.n29 3.4105
R15030 Iout.n804 Iout.n30 3.4105
R15031 Iout.n807 Iout.n31 3.4105
R15032 Iout.n873 Iout.n872 3.4105
R15033 Iout.n744 Iout.n743 3.4105
R15034 Iout.n740 Iout.n739 3.4105
R15035 Iout.n732 Iout.n731 3.4105
R15036 Iout.n728 Iout.n727 3.4105
R15037 Iout.n720 Iout.n719 3.4105
R15038 Iout.n795 Iout.n27 3.4105
R15039 Iout.n901 Iout.n900 3.4105
R15040 Iout.n722 Iout.n721 3.4105
R15041 Iout.n726 Iout.n725 3.4105
R15042 Iout.n734 Iout.n733 3.4105
R15043 Iout.n738 Iout.n737 3.4105
R15044 Iout.n746 Iout.n745 3.4105
R15045 Iout.n750 Iout.n749 3.4105
R15046 Iout.n752 Iout.n751 3.4105
R15047 Iout.n810 Iout.n32 3.4105
R15048 Iout.n865 Iout.n864 3.4105
R15049 Iout.n668 Iout.n55 3.4105
R15050 Iout.n671 Iout.n58 3.4105
R15051 Iout.n674 Iout.n61 3.4105
R15052 Iout.n677 Iout.n64 3.4105
R15053 Iout.n680 Iout.n67 3.4105
R15054 Iout.n683 Iout.n70 3.4105
R15055 Iout.n686 Iout.n73 3.4105
R15056 Iout.n714 Iout.n713 3.4105
R15057 Iout.n716 Iout.n715 3.4105
R15058 Iout.n792 Iout.n26 3.4105
R15059 Iout.n907 Iout.n906 3.4105
R15060 Iout.n587 Iout.n586 3.4105
R15061 Iout.n591 Iout.n590 3.4105
R15062 Iout.n599 Iout.n598 3.4105
R15063 Iout.n603 Iout.n602 3.4105
R15064 Iout.n611 Iout.n610 3.4105
R15065 Iout.n615 Iout.n614 3.4105
R15066 Iout.n623 Iout.n622 3.4105
R15067 Iout.n627 Iout.n626 3.4105
R15068 Iout.n665 Iout.n52 3.4105
R15069 Iout.n758 Iout.n757 3.4105
R15070 Iout.n756 Iout.n755 3.4105
R15071 Iout.n813 Iout.n33 3.4105
R15072 Iout.n859 Iout.n858 3.4105
R15073 Iout.n629 Iout.n628 3.4105
R15074 Iout.n621 Iout.n620 3.4105
R15075 Iout.n617 Iout.n616 3.4105
R15076 Iout.n609 Iout.n608 3.4105
R15077 Iout.n605 Iout.n604 3.4105
R15078 Iout.n597 Iout.n596 3.4105
R15079 Iout.n593 Iout.n592 3.4105
R15080 Iout.n585 Iout.n584 3.4105
R15081 Iout.n581 Iout.n580 3.4105
R15082 Iout.n579 Iout.n578 3.4105
R15083 Iout.n689 Iout.n76 3.4105
R15084 Iout.n710 Iout.n709 3.4105
R15085 Iout.n708 Iout.n707 3.4105
R15086 Iout.n789 Iout.n25 3.4105
R15087 Iout.n915 Iout.n914 3.4105
R15088 Iout.n572 Iout.n571 3.4105
R15089 Iout.n335 Iout.n116 3.4105
R15090 Iout.n338 Iout.n113 3.4105
R15091 Iout.n341 Iout.n110 3.4105
R15092 Iout.n344 Iout.n107 3.4105
R15093 Iout.n347 Iout.n104 3.4105
R15094 Iout.n350 Iout.n101 3.4105
R15095 Iout.n353 Iout.n98 3.4105
R15096 Iout.n356 Iout.n95 3.4105
R15097 Iout.n359 Iout.n92 3.4105
R15098 Iout.n633 Iout.n632 3.4105
R15099 Iout.n635 Iout.n634 3.4105
R15100 Iout.n662 Iout.n49 3.4105
R15101 Iout.n762 Iout.n761 3.4105
R15102 Iout.n764 Iout.n763 3.4105
R15103 Iout.n816 Iout.n34 3.4105
R15104 Iout.n851 Iout.n850 3.4105
R15105 Iout.n399 Iout.n398 3.4105
R15106 Iout.n405 Iout.n404 3.4105
R15107 Iout.n415 Iout.n414 3.4105
R15108 Iout.n421 Iout.n420 3.4105
R15109 Iout.n431 Iout.n430 3.4105
R15110 Iout.n444 Iout.n443 3.4105
R15111 Iout.n440 Iout.n159 3.4105
R15112 Iout.n437 Iout.n436 3.4105
R15113 Iout.n553 Iout.n552 3.4105
R15114 Iout.n556 Iout.n119 3.4105
R15115 Iout.n562 Iout.n561 3.4105
R15116 Iout.n568 Iout.n567 3.4105
R15117 Iout.n566 Iout.n565 3.4105
R15118 Iout.n575 Iout.n79 3.4105
R15119 Iout.n698 Iout.n697 3.4105
R15120 Iout.n702 Iout.n701 3.4105
R15121 Iout.n704 Iout.n703 3.4105
R15122 Iout.n786 Iout.n24 3.4105
R15123 Iout.n921 Iout.n920 3.4105
R15124 Iout.n129 Iout.n125 3.4105
R15125 Iout.n547 Iout.n546 3.4105
R15126 Iout.n551 Iout.n550 3.4105
R15127 Iout.n451 Iout.n158 3.4105
R15128 Iout.n455 Iout.n454 3.4105
R15129 Iout.n446 Iout.n445 3.4105
R15130 Iout.n429 Iout.n428 3.4105
R15131 Iout.n423 Iout.n422 3.4105
R15132 Iout.n413 Iout.n412 3.4105
R15133 Iout.n407 Iout.n406 3.4105
R15134 Iout.n397 Iout.n396 3.4105
R15135 Iout.n391 Iout.n390 3.4105
R15136 Iout.n389 Iout.n388 3.4105
R15137 Iout.n362 Iout.n89 3.4105
R15138 Iout.n641 Iout.n640 3.4105
R15139 Iout.n639 Iout.n638 3.4105
R15140 Iout.n659 Iout.n46 3.4105
R15141 Iout.n770 Iout.n769 3.4105
R15142 Iout.n768 Iout.n767 3.4105
R15143 Iout.n819 Iout.n35 3.4105
R15144 Iout.n845 Iout.n844 3.4105
R15145 Iout.n325 Iout.n165 3.4105
R15146 Iout.n322 Iout.n164 3.4105
R15147 Iout.n319 Iout.n163 3.4105
R15148 Iout.n316 Iout.n162 3.4105
R15149 Iout.n313 Iout.n161 3.4105
R15150 Iout.n310 Iout.n160 3.4105
R15151 Iout.n307 Iout.n155 3.4105
R15152 Iout.n457 Iout.n456 3.4105
R15153 Iout.n466 Iout.n465 3.4105
R15154 Iout.n462 Iout.n126 3.4105
R15155 Iout.n545 Iout.n544 3.4105
R15156 Iout.n541 Iout.n540 3.4105
R15157 Iout.n135 Iout.n3 3.4105
R15158 Iout.n987 Iout.n986 3.4105
R15159 Iout.n985 Iout.n984 3.4105
R15160 Iout.n122 Iout.n8 3.4105
R15161 Iout.n968 Iout.n967 3.4105
R15162 Iout.n966 Iout.n965 3.4105
R15163 Iout.n694 Iout.n13 3.4105
R15164 Iout.n949 Iout.n948 3.4105
R15165 Iout.n947 Iout.n946 3.4105
R15166 Iout.n783 Iout.n18 3.4105
R15167 Iout.n930 Iout.n929 3.4105
R15168 Iout.n1004 Iout.n1003 3.4105
R15169 Iout.n539 Iout.n538 3.4105
R15170 Iout.n533 Iout.n132 3.4105
R15171 Iout.n530 Iout.n529 3.4105
R15172 Iout.n468 Iout.n467 3.4105
R15173 Iout.n471 Iout.n153 3.4105
R15174 Iout.n475 Iout.n474 3.4105
R15175 Iout.n264 Iout.n263 3.4105
R15176 Iout.n268 Iout.n267 3.4105
R15177 Iout.n276 Iout.n275 3.4105
R15178 Iout.n280 Iout.n279 3.4105
R15179 Iout.n288 Iout.n287 3.4105
R15180 Iout.n292 Iout.n291 3.4105
R15181 Iout.n300 Iout.n299 3.4105
R15182 Iout.n328 Iout.n166 3.4105
R15183 Iout.n381 Iout.n380 3.4105
R15184 Iout.n383 Iout.n382 3.4105
R15185 Iout.n365 Iout.n83 3.4105
R15186 Iout.n645 Iout.n644 3.4105
R15187 Iout.n647 Iout.n646 3.4105
R15188 Iout.n656 Iout.n40 3.4105
R15189 Iout.n774 Iout.n773 3.4105
R15190 Iout.n776 Iout.n775 3.4105
R15191 Iout.n822 Iout.n36 3.4105
R15192 Iout.n837 Iout.n836 3.4105
R15193 Iout.n298 Iout.n297 3.4105
R15194 Iout.n294 Iout.n293 3.4105
R15195 Iout.n286 Iout.n285 3.4105
R15196 Iout.n282 Iout.n281 3.4105
R15197 Iout.n274 Iout.n273 3.4105
R15198 Iout.n270 Iout.n269 3.4105
R15199 Iout.n262 Iout.n261 3.4105
R15200 Iout.n477 Iout.n476 3.4105
R15201 Iout.n486 Iout.n485 3.4105
R15202 Iout.n482 Iout.n151 3.4105
R15203 Iout.n528 Iout.n527 3.4105
R15204 Iout.n524 Iout.n523 3.4105
R15205 Iout.n142 Iout.n138 3.4105
R15206 Iout.n1006 Iout.n1005 3.4105
R15207 Iout.n1009 Iout.n0 3.4105
R15208 Iout.n1000 Iout.n999 3.4105
R15209 Iout.n998 Iout.n997 3.4105
R15210 Iout.n990 Iout.n6 3.4105
R15211 Iout.n981 Iout.n980 3.4105
R15212 Iout.n979 Iout.n978 3.4105
R15213 Iout.n971 Iout.n11 3.4105
R15214 Iout.n962 Iout.n961 3.4105
R15215 Iout.n960 Iout.n959 3.4105
R15216 Iout.n952 Iout.n16 3.4105
R15217 Iout.n943 Iout.n942 3.4105
R15218 Iout.n941 Iout.n940 3.4105
R15219 Iout.n933 Iout.n21 3.4105
R15220 Iout.n1017 Iout.n1016 3.4105
R15221 Iout.n148 Iout.n2 3.4105
R15222 Iout.n518 Iout.n517 3.4105
R15223 Iout.n522 Iout.n521 3.4105
R15224 Iout.n493 Iout.n139 3.4105
R15225 Iout.n497 Iout.n496 3.4105
R15226 Iout.n488 Iout.n487 3.4105
R15227 Iout.n254 Iout.n154 3.4105
R15228 Iout.n258 Iout.n257 3.4105
R15229 Iout.n249 Iout.n188 3.4105
R15230 Iout.n246 Iout.n185 3.4105
R15231 Iout.n243 Iout.n182 3.4105
R15232 Iout.n240 Iout.n179 3.4105
R15233 Iout.n237 Iout.n176 3.4105
R15234 Iout.n234 Iout.n170 3.4105
R15235 Iout.n231 Iout.n230 3.4105
R15236 Iout.n171 Iout.n167 3.4105
R15237 Iout.n304 Iout.n303 3.4105
R15238 Iout.n332 Iout.n331 3.4105
R15239 Iout.n375 Iout.n374 3.4105
R15240 Iout.n373 Iout.n372 3.4105
R15241 Iout.n369 Iout.n368 3.4105
R15242 Iout.n84 Iout.n80 3.4105
R15243 Iout.n651 Iout.n650 3.4105
R15244 Iout.n653 Iout.n652 3.4105
R15245 Iout.n41 Iout.n37 3.4105
R15246 Iout.n780 Iout.n779 3.4105
R15247 Iout.n826 Iout.n825 3.4105
R15248 Iout.n831 Iout.n830 3.4105
R15249 Iout.n229 Iout.n228 3.4105
R15250 Iout.n225 Iout.n224 3.4105
R15251 Iout.n221 Iout.n220 3.4105
R15252 Iout.n217 Iout.n216 3.4105
R15253 Iout.n213 Iout.n212 3.4105
R15254 Iout.n209 Iout.n208 3.4105
R15255 Iout.n205 Iout.n204 3.4105
R15256 Iout.n201 Iout.n191 3.4105
R15257 Iout.n198 Iout.n197 3.4105
R15258 Iout.n194 Iout.n152 3.4105
R15259 Iout.n499 Iout.n498 3.4105
R15260 Iout.n503 Iout.n502 3.4105
R15261 Iout.n506 Iout.n145 3.4105
R15262 Iout.n516 Iout.n515 3.4105
R15263 Iout.n512 Iout.n511 3.4105
R15264 Iout.n1019 Iout.n1018 3.4105
R15265 Iout.n936 Iout.n23 1.43848
R15266 Iout.n936 Iout.n935 1.34612
R15267 Iout.n939 Iout.n937 1.34612
R15268 Iout.n20 Iout.n17 1.34612
R15269 Iout.n955 Iout.n954 1.34612
R15270 Iout.n958 Iout.n956 1.34612
R15271 Iout.n15 Iout.n12 1.34612
R15272 Iout.n974 Iout.n973 1.34612
R15273 Iout.n977 Iout.n975 1.34612
R15274 Iout.n10 Iout.n7 1.34612
R15275 Iout.n993 Iout.n992 1.34612
R15276 Iout.n996 Iout.n994 1.34612
R15277 Iout.n5 Iout.n1 1.34612
R15278 Iout.n1012 Iout.n1011 1.34612
R15279 Iout.n1015 Iout.n1013 1.34612
R15280 Iout.n1022 Iout.n1021 1.34612
R15281 Iout.n197 Iout.n154 0.451012
R15282 Iout.n476 Iout.n154 0.451012
R15283 Iout.n476 Iout.n475 0.451012
R15284 Iout.n475 Iout.n155 0.451012
R15285 Iout.n445 Iout.n155 0.451012
R15286 Iout.n445 Iout.n444 0.451012
R15287 Iout.n444 Iout.n107 0.451012
R15288 Iout.n604 Iout.n107 0.451012
R15289 Iout.n604 Iout.n603 0.451012
R15290 Iout.n603 Iout.n64 0.451012
R15291 Iout.n733 Iout.n64 0.451012
R15292 Iout.n733 Iout.n732 0.451012
R15293 Iout.n732 Iout.n29 0.451012
R15294 Iout.n886 Iout.n29 0.451012
R15295 Iout.n258 Iout.n191 0.451012
R15296 Iout.n262 Iout.n258 0.451012
R15297 Iout.n263 Iout.n262 0.451012
R15298 Iout.n263 Iout.n160 0.451012
R15299 Iout.n429 Iout.n160 0.451012
R15300 Iout.n430 Iout.n429 0.451012
R15301 Iout.n430 Iout.n104 0.451012
R15302 Iout.n609 Iout.n104 0.451012
R15303 Iout.n610 Iout.n609 0.451012
R15304 Iout.n610 Iout.n61 0.451012
R15305 Iout.n738 Iout.n61 0.451012
R15306 Iout.n739 Iout.n738 0.451012
R15307 Iout.n739 Iout.n30 0.451012
R15308 Iout.n879 Iout.n30 0.451012
R15309 Iout.n487 Iout.n152 0.451012
R15310 Iout.n487 Iout.n486 0.451012
R15311 Iout.n486 Iout.n153 0.451012
R15312 Iout.n456 Iout.n153 0.451012
R15313 Iout.n456 Iout.n455 0.451012
R15314 Iout.n455 Iout.n159 0.451012
R15315 Iout.n159 Iout.n110 0.451012
R15316 Iout.n597 Iout.n110 0.451012
R15317 Iout.n598 Iout.n597 0.451012
R15318 Iout.n598 Iout.n67 0.451012
R15319 Iout.n726 Iout.n67 0.451012
R15320 Iout.n727 Iout.n726 0.451012
R15321 Iout.n727 Iout.n28 0.451012
R15322 Iout.n893 Iout.n28 0.451012
R15323 Iout.n204 Iout.n188 0.451012
R15324 Iout.n269 Iout.n188 0.451012
R15325 Iout.n269 Iout.n268 0.451012
R15326 Iout.n268 Iout.n161 0.451012
R15327 Iout.n422 Iout.n161 0.451012
R15328 Iout.n422 Iout.n421 0.451012
R15329 Iout.n421 Iout.n101 0.451012
R15330 Iout.n616 Iout.n101 0.451012
R15331 Iout.n616 Iout.n615 0.451012
R15332 Iout.n615 Iout.n58 0.451012
R15333 Iout.n745 Iout.n58 0.451012
R15334 Iout.n745 Iout.n744 0.451012
R15335 Iout.n744 Iout.n31 0.451012
R15336 Iout.n872 Iout.n31 0.451012
R15337 Iout.n498 Iout.n497 0.451012
R15338 Iout.n497 Iout.n151 0.451012
R15339 Iout.n467 Iout.n151 0.451012
R15340 Iout.n467 Iout.n466 0.451012
R15341 Iout.n466 Iout.n158 0.451012
R15342 Iout.n436 Iout.n158 0.451012
R15343 Iout.n436 Iout.n113 0.451012
R15344 Iout.n592 Iout.n113 0.451012
R15345 Iout.n592 Iout.n591 0.451012
R15346 Iout.n591 Iout.n70 0.451012
R15347 Iout.n721 Iout.n70 0.451012
R15348 Iout.n721 Iout.n720 0.451012
R15349 Iout.n720 Iout.n27 0.451012
R15350 Iout.n900 Iout.n27 0.451012
R15351 Iout.n208 Iout.n185 0.451012
R15352 Iout.n274 Iout.n185 0.451012
R15353 Iout.n275 Iout.n274 0.451012
R15354 Iout.n275 Iout.n162 0.451012
R15355 Iout.n413 Iout.n162 0.451012
R15356 Iout.n414 Iout.n413 0.451012
R15357 Iout.n414 Iout.n98 0.451012
R15358 Iout.n621 Iout.n98 0.451012
R15359 Iout.n622 Iout.n621 0.451012
R15360 Iout.n622 Iout.n55 0.451012
R15361 Iout.n750 Iout.n55 0.451012
R15362 Iout.n751 Iout.n750 0.451012
R15363 Iout.n751 Iout.n32 0.451012
R15364 Iout.n865 Iout.n32 0.451012
R15365 Iout.n502 Iout.n139 0.451012
R15366 Iout.n528 Iout.n139 0.451012
R15367 Iout.n529 Iout.n528 0.451012
R15368 Iout.n529 Iout.n126 0.451012
R15369 Iout.n551 Iout.n126 0.451012
R15370 Iout.n552 Iout.n551 0.451012
R15371 Iout.n552 Iout.n116 0.451012
R15372 Iout.n585 Iout.n116 0.451012
R15373 Iout.n586 Iout.n585 0.451012
R15374 Iout.n586 Iout.n73 0.451012
R15375 Iout.n714 Iout.n73 0.451012
R15376 Iout.n715 Iout.n714 0.451012
R15377 Iout.n715 Iout.n26 0.451012
R15378 Iout.n907 Iout.n26 0.451012
R15379 Iout.n212 Iout.n182 0.451012
R15380 Iout.n281 Iout.n182 0.451012
R15381 Iout.n281 Iout.n280 0.451012
R15382 Iout.n280 Iout.n163 0.451012
R15383 Iout.n406 Iout.n163 0.451012
R15384 Iout.n406 Iout.n405 0.451012
R15385 Iout.n405 Iout.n95 0.451012
R15386 Iout.n628 Iout.n95 0.451012
R15387 Iout.n628 Iout.n627 0.451012
R15388 Iout.n627 Iout.n52 0.451012
R15389 Iout.n757 Iout.n52 0.451012
R15390 Iout.n757 Iout.n756 0.451012
R15391 Iout.n756 Iout.n33 0.451012
R15392 Iout.n858 Iout.n33 0.451012
R15393 Iout.n522 Iout.n145 0.451012
R15394 Iout.n523 Iout.n522 0.451012
R15395 Iout.n523 Iout.n132 0.451012
R15396 Iout.n545 Iout.n132 0.451012
R15397 Iout.n546 Iout.n545 0.451012
R15398 Iout.n546 Iout.n119 0.451012
R15399 Iout.n572 Iout.n119 0.451012
R15400 Iout.n580 Iout.n572 0.451012
R15401 Iout.n580 Iout.n579 0.451012
R15402 Iout.n579 Iout.n76 0.451012
R15403 Iout.n709 Iout.n76 0.451012
R15404 Iout.n709 Iout.n708 0.451012
R15405 Iout.n708 Iout.n25 0.451012
R15406 Iout.n914 Iout.n25 0.451012
R15407 Iout.n216 Iout.n179 0.451012
R15408 Iout.n286 Iout.n179 0.451012
R15409 Iout.n287 Iout.n286 0.451012
R15410 Iout.n287 Iout.n164 0.451012
R15411 Iout.n397 Iout.n164 0.451012
R15412 Iout.n398 Iout.n397 0.451012
R15413 Iout.n398 Iout.n92 0.451012
R15414 Iout.n633 Iout.n92 0.451012
R15415 Iout.n634 Iout.n633 0.451012
R15416 Iout.n634 Iout.n49 0.451012
R15417 Iout.n762 Iout.n49 0.451012
R15418 Iout.n763 Iout.n762 0.451012
R15419 Iout.n763 Iout.n34 0.451012
R15420 Iout.n851 Iout.n34 0.451012
R15421 Iout.n517 Iout.n516 0.451012
R15422 Iout.n517 Iout.n138 0.451012
R15423 Iout.n539 Iout.n138 0.451012
R15424 Iout.n540 Iout.n539 0.451012
R15425 Iout.n540 Iout.n125 0.451012
R15426 Iout.n562 Iout.n125 0.451012
R15427 Iout.n567 Iout.n562 0.451012
R15428 Iout.n567 Iout.n566 0.451012
R15429 Iout.n566 Iout.n79 0.451012
R15430 Iout.n698 Iout.n79 0.451012
R15431 Iout.n702 Iout.n698 0.451012
R15432 Iout.n703 Iout.n702 0.451012
R15433 Iout.n703 Iout.n24 0.451012
R15434 Iout.n921 Iout.n24 0.451012
R15435 Iout.n220 Iout.n176 0.451012
R15436 Iout.n293 Iout.n176 0.451012
R15437 Iout.n293 Iout.n292 0.451012
R15438 Iout.n292 Iout.n165 0.451012
R15439 Iout.n390 Iout.n165 0.451012
R15440 Iout.n390 Iout.n389 0.451012
R15441 Iout.n389 Iout.n89 0.451012
R15442 Iout.n640 Iout.n89 0.451012
R15443 Iout.n640 Iout.n639 0.451012
R15444 Iout.n639 Iout.n46 0.451012
R15445 Iout.n769 Iout.n46 0.451012
R15446 Iout.n769 Iout.n768 0.451012
R15447 Iout.n768 Iout.n35 0.451012
R15448 Iout.n844 Iout.n35 0.451012
R15449 Iout.n511 Iout.n2 0.451012
R15450 Iout.n1005 Iout.n2 0.451012
R15451 Iout.n1005 Iout.n1004 0.451012
R15452 Iout.n1004 Iout.n3 0.451012
R15453 Iout.n986 Iout.n3 0.451012
R15454 Iout.n986 Iout.n985 0.451012
R15455 Iout.n985 Iout.n8 0.451012
R15456 Iout.n967 Iout.n8 0.451012
R15457 Iout.n967 Iout.n966 0.451012
R15458 Iout.n966 Iout.n13 0.451012
R15459 Iout.n948 Iout.n13 0.451012
R15460 Iout.n948 Iout.n947 0.451012
R15461 Iout.n947 Iout.n18 0.451012
R15462 Iout.n929 Iout.n18 0.451012
R15463 Iout.n224 Iout.n170 0.451012
R15464 Iout.n298 Iout.n170 0.451012
R15465 Iout.n299 Iout.n298 0.451012
R15466 Iout.n299 Iout.n166 0.451012
R15467 Iout.n381 Iout.n166 0.451012
R15468 Iout.n382 Iout.n381 0.451012
R15469 Iout.n382 Iout.n83 0.451012
R15470 Iout.n645 Iout.n83 0.451012
R15471 Iout.n646 Iout.n645 0.451012
R15472 Iout.n646 Iout.n40 0.451012
R15473 Iout.n774 Iout.n40 0.451012
R15474 Iout.n775 Iout.n774 0.451012
R15475 Iout.n775 Iout.n36 0.451012
R15476 Iout.n837 Iout.n36 0.451012
R15477 Iout.n1018 Iout.n1017 0.451012
R15478 Iout.n1017 Iout.n0 0.451012
R15479 Iout.n999 Iout.n0 0.451012
R15480 Iout.n999 Iout.n998 0.451012
R15481 Iout.n998 Iout.n6 0.451012
R15482 Iout.n980 Iout.n6 0.451012
R15483 Iout.n980 Iout.n979 0.451012
R15484 Iout.n979 Iout.n11 0.451012
R15485 Iout.n961 Iout.n11 0.451012
R15486 Iout.n961 Iout.n960 0.451012
R15487 Iout.n960 Iout.n16 0.451012
R15488 Iout.n942 Iout.n16 0.451012
R15489 Iout.n942 Iout.n941 0.451012
R15490 Iout.n941 Iout.n21 0.451012
R15491 Iout.n230 Iout.n229 0.451012
R15492 Iout.n230 Iout.n167 0.451012
R15493 Iout.n304 Iout.n167 0.451012
R15494 Iout.n332 Iout.n304 0.451012
R15495 Iout.n374 Iout.n332 0.451012
R15496 Iout.n374 Iout.n373 0.451012
R15497 Iout.n373 Iout.n369 0.451012
R15498 Iout.n369 Iout.n80 0.451012
R15499 Iout.n651 Iout.n80 0.451012
R15500 Iout.n652 Iout.n651 0.451012
R15501 Iout.n652 Iout.n37 0.451012
R15502 Iout.n780 Iout.n37 0.451012
R15503 Iout.n826 Iout.n780 0.451012
R15504 Iout.n830 Iout.n826 0.451012
R15505 Iout.n231 Iout 0.2919
R15506 Iout.n303 Iout 0.2919
R15507 Iout Iout.n300 0.2919
R15508 Iout.n375 Iout 0.2919
R15509 Iout.n380 Iout 0.2919
R15510 Iout.n391 Iout 0.2919
R15511 Iout.n368 Iout 0.2919
R15512 Iout Iout.n365 0.2919
R15513 Iout Iout.n362 0.2919
R15514 Iout Iout.n359 0.2919
R15515 Iout.n650 Iout 0.2919
R15516 Iout Iout.n647 0.2919
R15517 Iout.n638 Iout 0.2919
R15518 Iout Iout.n635 0.2919
R15519 Iout.n626 Iout 0.2919
R15520 Iout.n41 Iout 0.2919
R15521 Iout.n773 Iout 0.2919
R15522 Iout Iout.n770 0.2919
R15523 Iout.n761 Iout 0.2919
R15524 Iout Iout.n758 0.2919
R15525 Iout.n749 Iout 0.2919
R15526 Iout.n825 Iout 0.2919
R15527 Iout Iout.n822 0.2919
R15528 Iout Iout.n819 0.2919
R15529 Iout Iout.n816 0.2919
R15530 Iout Iout.n813 0.2919
R15531 Iout Iout.n810 0.2919
R15532 Iout Iout.n807 0.2919
R15533 Iout.n829 Iout 0.2919
R15534 Iout.n838 Iout 0.2919
R15535 Iout.n843 Iout 0.2919
R15536 Iout.n852 Iout 0.2919
R15537 Iout.n857 Iout 0.2919
R15538 Iout.n866 Iout 0.2919
R15539 Iout.n871 Iout 0.2919
R15540 Iout.n880 Iout 0.2919
R15541 Iout Iout.n925 0.2919
R15542 Iout.n928 Iout 0.2919
R15543 Iout.n922 Iout 0.2919
R15544 Iout.n913 Iout 0.2919
R15545 Iout.n908 Iout 0.2919
R15546 Iout.n899 Iout 0.2919
R15547 Iout.n894 Iout 0.2919
R15548 Iout.n885 Iout 0.2919
R15549 Iout.n831 Iout 0.2919
R15550 Iout.n836 Iout 0.2919
R15551 Iout.n845 Iout 0.2919
R15552 Iout.n850 Iout 0.2919
R15553 Iout.n859 Iout 0.2919
R15554 Iout.n864 Iout 0.2919
R15555 Iout.n873 Iout 0.2919
R15556 Iout.n878 Iout 0.2919
R15557 Iout.n887 Iout 0.2919
R15558 Iout.n892 Iout 0.2919
R15559 Iout.n933 Iout 0.2919
R15560 Iout.n930 Iout 0.2919
R15561 Iout.n920 Iout 0.2919
R15562 Iout.n915 Iout 0.2919
R15563 Iout.n906 Iout 0.2919
R15564 Iout.n901 Iout 0.2919
R15565 Iout.n940 Iout 0.2919
R15566 Iout Iout.n783 0.2919
R15567 Iout Iout.n786 0.2919
R15568 Iout Iout.n789 0.2919
R15569 Iout Iout.n792 0.2919
R15570 Iout Iout.n795 0.2919
R15571 Iout Iout.n798 0.2919
R15572 Iout Iout.n801 0.2919
R15573 Iout Iout.n804 0.2919
R15574 Iout.n779 Iout 0.2919
R15575 Iout Iout.n776 0.2919
R15576 Iout.n767 Iout 0.2919
R15577 Iout Iout.n764 0.2919
R15578 Iout.n755 Iout 0.2919
R15579 Iout Iout.n752 0.2919
R15580 Iout.n743 Iout 0.2919
R15581 Iout Iout.n740 0.2919
R15582 Iout.n731 Iout 0.2919
R15583 Iout Iout.n728 0.2919
R15584 Iout.n719 Iout 0.2919
R15585 Iout Iout.n943 0.2919
R15586 Iout.n946 Iout 0.2919
R15587 Iout Iout.n704 0.2919
R15588 Iout.n707 Iout 0.2919
R15589 Iout Iout.n716 0.2919
R15590 Iout.n952 Iout 0.2919
R15591 Iout.n949 Iout 0.2919
R15592 Iout.n701 Iout 0.2919
R15593 Iout Iout.n710 0.2919
R15594 Iout.n713 Iout 0.2919
R15595 Iout Iout.n722 0.2919
R15596 Iout.n725 Iout 0.2919
R15597 Iout Iout.n734 0.2919
R15598 Iout.n737 Iout 0.2919
R15599 Iout Iout.n746 0.2919
R15600 Iout.n653 Iout 0.2919
R15601 Iout.n656 Iout 0.2919
R15602 Iout.n659 Iout 0.2919
R15603 Iout.n662 Iout 0.2919
R15604 Iout.n665 Iout 0.2919
R15605 Iout.n668 Iout 0.2919
R15606 Iout.n671 Iout 0.2919
R15607 Iout.n674 Iout 0.2919
R15608 Iout.n677 Iout 0.2919
R15609 Iout.n680 Iout 0.2919
R15610 Iout.n683 Iout 0.2919
R15611 Iout.n686 Iout 0.2919
R15612 Iout.n959 Iout 0.2919
R15613 Iout Iout.n694 0.2919
R15614 Iout.n697 Iout 0.2919
R15615 Iout.n689 Iout 0.2919
R15616 Iout Iout.n962 0.2919
R15617 Iout.n965 Iout 0.2919
R15618 Iout Iout.n575 0.2919
R15619 Iout.n578 Iout 0.2919
R15620 Iout Iout.n587 0.2919
R15621 Iout.n590 Iout 0.2919
R15622 Iout Iout.n599 0.2919
R15623 Iout.n602 Iout 0.2919
R15624 Iout Iout.n611 0.2919
R15625 Iout.n614 Iout 0.2919
R15626 Iout Iout.n623 0.2919
R15627 Iout.n84 Iout 0.2919
R15628 Iout.n644 Iout 0.2919
R15629 Iout Iout.n641 0.2919
R15630 Iout.n632 Iout 0.2919
R15631 Iout Iout.n629 0.2919
R15632 Iout.n620 Iout 0.2919
R15633 Iout Iout.n617 0.2919
R15634 Iout.n608 Iout 0.2919
R15635 Iout Iout.n605 0.2919
R15636 Iout.n596 Iout 0.2919
R15637 Iout Iout.n593 0.2919
R15638 Iout.n584 Iout 0.2919
R15639 Iout Iout.n581 0.2919
R15640 Iout.n971 Iout 0.2919
R15641 Iout.n968 Iout 0.2919
R15642 Iout.n565 Iout 0.2919
R15643 Iout.n978 Iout 0.2919
R15644 Iout Iout.n122 0.2919
R15645 Iout Iout.n568 0.2919
R15646 Iout.n571 Iout 0.2919
R15647 Iout Iout.n335 0.2919
R15648 Iout Iout.n338 0.2919
R15649 Iout Iout.n341 0.2919
R15650 Iout Iout.n344 0.2919
R15651 Iout Iout.n347 0.2919
R15652 Iout Iout.n350 0.2919
R15653 Iout Iout.n353 0.2919
R15654 Iout Iout.n356 0.2919
R15655 Iout.n372 Iout 0.2919
R15656 Iout.n383 Iout 0.2919
R15657 Iout.n388 Iout 0.2919
R15658 Iout.n399 Iout 0.2919
R15659 Iout.n404 Iout 0.2919
R15660 Iout.n415 Iout 0.2919
R15661 Iout.n420 Iout 0.2919
R15662 Iout.n431 Iout 0.2919
R15663 Iout.n443 Iout 0.2919
R15664 Iout Iout.n440 0.2919
R15665 Iout Iout.n437 0.2919
R15666 Iout.n553 Iout 0.2919
R15667 Iout.n556 Iout 0.2919
R15668 Iout.n561 Iout 0.2919
R15669 Iout Iout.n981 0.2919
R15670 Iout.n984 Iout 0.2919
R15671 Iout.n990 Iout 0.2919
R15672 Iout.n987 Iout 0.2919
R15673 Iout Iout.n129 0.2919
R15674 Iout Iout.n547 0.2919
R15675 Iout.n550 Iout 0.2919
R15676 Iout Iout.n451 0.2919
R15677 Iout.n454 Iout 0.2919
R15678 Iout.n446 Iout 0.2919
R15679 Iout.n428 Iout 0.2919
R15680 Iout.n423 Iout 0.2919
R15681 Iout.n412 Iout 0.2919
R15682 Iout.n407 Iout 0.2919
R15683 Iout.n396 Iout 0.2919
R15684 Iout.n331 Iout 0.2919
R15685 Iout Iout.n328 0.2919
R15686 Iout Iout.n325 0.2919
R15687 Iout Iout.n322 0.2919
R15688 Iout Iout.n319 0.2919
R15689 Iout Iout.n316 0.2919
R15690 Iout Iout.n313 0.2919
R15691 Iout Iout.n310 0.2919
R15692 Iout Iout.n307 0.2919
R15693 Iout.n457 Iout 0.2919
R15694 Iout.n465 Iout 0.2919
R15695 Iout Iout.n462 0.2919
R15696 Iout.n544 Iout 0.2919
R15697 Iout Iout.n541 0.2919
R15698 Iout Iout.n135 0.2919
R15699 Iout.n997 Iout 0.2919
R15700 Iout Iout.n1000 0.2919
R15701 Iout.n1003 Iout 0.2919
R15702 Iout.n538 Iout 0.2919
R15703 Iout.n533 Iout 0.2919
R15704 Iout.n530 Iout 0.2919
R15705 Iout Iout.n468 0.2919
R15706 Iout Iout.n471 0.2919
R15707 Iout.n474 Iout 0.2919
R15708 Iout Iout.n264 0.2919
R15709 Iout.n267 Iout 0.2919
R15710 Iout Iout.n276 0.2919
R15711 Iout.n279 Iout 0.2919
R15712 Iout Iout.n288 0.2919
R15713 Iout.n291 Iout 0.2919
R15714 Iout.n171 Iout 0.2919
R15715 Iout.n297 Iout 0.2919
R15716 Iout Iout.n294 0.2919
R15717 Iout.n285 Iout 0.2919
R15718 Iout Iout.n282 0.2919
R15719 Iout.n273 Iout 0.2919
R15720 Iout Iout.n270 0.2919
R15721 Iout.n261 Iout 0.2919
R15722 Iout.n477 Iout 0.2919
R15723 Iout.n485 Iout 0.2919
R15724 Iout Iout.n482 0.2919
R15725 Iout.n527 Iout 0.2919
R15726 Iout Iout.n524 0.2919
R15727 Iout Iout.n142 0.2919
R15728 Iout.n1006 Iout 0.2919
R15729 Iout.n1009 Iout 0.2919
R15730 Iout.n1016 Iout 0.2919
R15731 Iout Iout.n148 0.2919
R15732 Iout Iout.n518 0.2919
R15733 Iout.n521 Iout 0.2919
R15734 Iout Iout.n493 0.2919
R15735 Iout.n496 Iout 0.2919
R15736 Iout.n488 Iout 0.2919
R15737 Iout Iout.n254 0.2919
R15738 Iout.n257 Iout 0.2919
R15739 Iout.n249 Iout 0.2919
R15740 Iout.n246 Iout 0.2919
R15741 Iout.n243 Iout 0.2919
R15742 Iout.n240 Iout 0.2919
R15743 Iout.n237 Iout 0.2919
R15744 Iout.n234 Iout 0.2919
R15745 Iout.n228 Iout 0.2919
R15746 Iout Iout.n225 0.2919
R15747 Iout Iout.n221 0.2919
R15748 Iout Iout.n217 0.2919
R15749 Iout Iout.n213 0.2919
R15750 Iout Iout.n209 0.2919
R15751 Iout Iout.n205 0.2919
R15752 Iout Iout.n201 0.2919
R15753 Iout Iout.n198 0.2919
R15754 Iout Iout.n194 0.2919
R15755 Iout.n499 Iout 0.2919
R15756 Iout.n503 Iout 0.2919
R15757 Iout.n506 Iout 0.2919
R15758 Iout.n515 Iout 0.2919
R15759 Iout Iout.n512 0.2919
R15760 Iout.n1019 Iout 0.2919
R15761 Iout.n1013 Iout.n1012 0.092855
R15762 Iout.n1012 Iout.n1 0.092855
R15763 Iout.n994 Iout.n1 0.092855
R15764 Iout.n994 Iout.n993 0.092855
R15765 Iout.n993 Iout.n7 0.092855
R15766 Iout.n975 Iout.n7 0.092855
R15767 Iout.n975 Iout.n974 0.092855
R15768 Iout.n974 Iout.n12 0.092855
R15769 Iout.n956 Iout.n12 0.092855
R15770 Iout.n956 Iout.n955 0.092855
R15771 Iout.n955 Iout.n17 0.092855
R15772 Iout.n937 Iout.n17 0.092855
R15773 Iout.n937 Iout.n936 0.092855
R15774 Iout.n197 Iout 0.0818902
R15775 Iout.n191 Iout 0.0818902
R15776 Iout.n152 Iout 0.0818902
R15777 Iout.n204 Iout 0.0818902
R15778 Iout.n498 Iout 0.0818902
R15779 Iout.n208 Iout 0.0818902
R15780 Iout.n502 Iout 0.0818902
R15781 Iout.n212 Iout 0.0818902
R15782 Iout.n145 Iout 0.0818902
R15783 Iout.n216 Iout 0.0818902
R15784 Iout.n516 Iout 0.0818902
R15785 Iout.n220 Iout 0.0818902
R15786 Iout.n511 Iout 0.0818902
R15787 Iout.n224 Iout 0.0818902
R15788 Iout.n1018 Iout 0.0818902
R15789 Iout.n229 Iout 0.0818902
R15790 Iout.n1013 Iout 0.072645
R15791 Iout.n302 Iout 0.0532071
R15792 Iout Iout.n377 0.0532071
R15793 Iout.n379 Iout 0.0532071
R15794 Iout.n367 Iout 0.0532071
R15795 Iout.n364 Iout 0.0532071
R15796 Iout.n361 Iout 0.0532071
R15797 Iout.n649 Iout 0.0532071
R15798 Iout Iout.n82 0.0532071
R15799 Iout.n637 Iout 0.0532071
R15800 Iout Iout.n91 0.0532071
R15801 Iout Iout.n43 0.0532071
R15802 Iout.n772 Iout 0.0532071
R15803 Iout Iout.n45 0.0532071
R15804 Iout.n760 Iout 0.0532071
R15805 Iout Iout.n51 0.0532071
R15806 Iout.n824 Iout 0.0532071
R15807 Iout.n821 Iout 0.0532071
R15808 Iout.n818 Iout 0.0532071
R15809 Iout.n815 Iout 0.0532071
R15810 Iout.n812 Iout 0.0532071
R15811 Iout.n809 Iout 0.0532071
R15812 Iout.n828 Iout 0.0532071
R15813 Iout Iout.n840 0.0532071
R15814 Iout.n842 Iout 0.0532071
R15815 Iout Iout.n854 0.0532071
R15816 Iout.n856 Iout 0.0532071
R15817 Iout Iout.n868 0.0532071
R15818 Iout.n870 Iout 0.0532071
R15819 Iout.n927 Iout 0.0532071
R15820 Iout Iout.n924 0.0532071
R15821 Iout.n912 Iout 0.0532071
R15822 Iout Iout.n910 0.0532071
R15823 Iout.n898 Iout 0.0532071
R15824 Iout Iout.n896 0.0532071
R15825 Iout.n884 Iout 0.0532071
R15826 Iout Iout.n882 0.0532071
R15827 Iout Iout.n833 0.0532071
R15828 Iout.n835 Iout 0.0532071
R15829 Iout Iout.n847 0.0532071
R15830 Iout.n849 Iout 0.0532071
R15831 Iout Iout.n861 0.0532071
R15832 Iout.n863 Iout 0.0532071
R15833 Iout Iout.n875 0.0532071
R15834 Iout.n877 Iout 0.0532071
R15835 Iout Iout.n889 0.0532071
R15836 Iout Iout.n932 0.0532071
R15837 Iout.n919 Iout 0.0532071
R15838 Iout Iout.n917 0.0532071
R15839 Iout.n905 Iout 0.0532071
R15840 Iout Iout.n903 0.0532071
R15841 Iout.n891 Iout 0.0532071
R15842 Iout.n782 Iout 0.0532071
R15843 Iout.n785 Iout 0.0532071
R15844 Iout.n788 Iout 0.0532071
R15845 Iout.n791 Iout 0.0532071
R15846 Iout.n794 Iout 0.0532071
R15847 Iout.n797 Iout 0.0532071
R15848 Iout.n800 Iout 0.0532071
R15849 Iout.n803 Iout 0.0532071
R15850 Iout.n806 Iout 0.0532071
R15851 Iout.n778 Iout 0.0532071
R15852 Iout Iout.n39 0.0532071
R15853 Iout.n766 Iout 0.0532071
R15854 Iout Iout.n48 0.0532071
R15855 Iout.n754 Iout 0.0532071
R15856 Iout Iout.n54 0.0532071
R15857 Iout.n742 Iout 0.0532071
R15858 Iout Iout.n60 0.0532071
R15859 Iout.n730 Iout 0.0532071
R15860 Iout Iout.n66 0.0532071
R15861 Iout.n945 Iout 0.0532071
R15862 Iout.n78 Iout 0.0532071
R15863 Iout.n706 Iout 0.0532071
R15864 Iout Iout.n72 0.0532071
R15865 Iout.n718 Iout 0.0532071
R15866 Iout Iout.n951 0.0532071
R15867 Iout.n700 Iout 0.0532071
R15868 Iout Iout.n75 0.0532071
R15869 Iout.n712 Iout 0.0532071
R15870 Iout Iout.n69 0.0532071
R15871 Iout.n724 Iout 0.0532071
R15872 Iout Iout.n63 0.0532071
R15873 Iout.n736 Iout 0.0532071
R15874 Iout Iout.n57 0.0532071
R15875 Iout.n748 Iout 0.0532071
R15876 Iout Iout.n655 0.0532071
R15877 Iout Iout.n658 0.0532071
R15878 Iout Iout.n661 0.0532071
R15879 Iout Iout.n664 0.0532071
R15880 Iout Iout.n667 0.0532071
R15881 Iout Iout.n670 0.0532071
R15882 Iout Iout.n673 0.0532071
R15883 Iout Iout.n676 0.0532071
R15884 Iout Iout.n679 0.0532071
R15885 Iout Iout.n682 0.0532071
R15886 Iout Iout.n685 0.0532071
R15887 Iout.n693 Iout 0.0532071
R15888 Iout.n696 Iout 0.0532071
R15889 Iout Iout.n691 0.0532071
R15890 Iout Iout.n688 0.0532071
R15891 Iout.n964 Iout 0.0532071
R15892 Iout.n574 Iout 0.0532071
R15893 Iout.n577 Iout 0.0532071
R15894 Iout Iout.n115 0.0532071
R15895 Iout.n589 Iout 0.0532071
R15896 Iout Iout.n109 0.0532071
R15897 Iout.n601 Iout 0.0532071
R15898 Iout Iout.n103 0.0532071
R15899 Iout.n613 Iout 0.0532071
R15900 Iout Iout.n97 0.0532071
R15901 Iout.n625 Iout 0.0532071
R15902 Iout Iout.n86 0.0532071
R15903 Iout.n643 Iout 0.0532071
R15904 Iout Iout.n88 0.0532071
R15905 Iout.n631 Iout 0.0532071
R15906 Iout Iout.n94 0.0532071
R15907 Iout.n619 Iout 0.0532071
R15908 Iout Iout.n100 0.0532071
R15909 Iout.n607 Iout 0.0532071
R15910 Iout Iout.n106 0.0532071
R15911 Iout.n595 Iout 0.0532071
R15912 Iout Iout.n112 0.0532071
R15913 Iout.n583 Iout 0.0532071
R15914 Iout Iout.n970 0.0532071
R15915 Iout.n564 Iout 0.0532071
R15916 Iout Iout.n118 0.0532071
R15917 Iout.n121 Iout 0.0532071
R15918 Iout.n124 Iout 0.0532071
R15919 Iout.n570 Iout 0.0532071
R15920 Iout.n334 Iout 0.0532071
R15921 Iout.n337 Iout 0.0532071
R15922 Iout.n340 Iout 0.0532071
R15923 Iout.n343 Iout 0.0532071
R15924 Iout.n346 Iout 0.0532071
R15925 Iout.n349 Iout 0.0532071
R15926 Iout.n352 Iout 0.0532071
R15927 Iout.n355 Iout 0.0532071
R15928 Iout.n358 Iout 0.0532071
R15929 Iout.n371 Iout 0.0532071
R15930 Iout Iout.n385 0.0532071
R15931 Iout.n387 Iout 0.0532071
R15932 Iout Iout.n401 0.0532071
R15933 Iout.n403 Iout 0.0532071
R15934 Iout Iout.n417 0.0532071
R15935 Iout.n419 Iout 0.0532071
R15936 Iout Iout.n433 0.0532071
R15937 Iout.n442 Iout 0.0532071
R15938 Iout.n439 Iout 0.0532071
R15939 Iout.n435 Iout 0.0532071
R15940 Iout Iout.n555 0.0532071
R15941 Iout Iout.n558 0.0532071
R15942 Iout.n983 Iout 0.0532071
R15943 Iout.n560 Iout 0.0532071
R15944 Iout Iout.n989 0.0532071
R15945 Iout.n128 Iout 0.0532071
R15946 Iout.n131 Iout 0.0532071
R15947 Iout.n549 Iout 0.0532071
R15948 Iout.n450 Iout 0.0532071
R15949 Iout.n453 Iout 0.0532071
R15950 Iout Iout.n448 0.0532071
R15951 Iout.n427 Iout 0.0532071
R15952 Iout Iout.n425 0.0532071
R15953 Iout.n411 Iout 0.0532071
R15954 Iout Iout.n409 0.0532071
R15955 Iout.n395 Iout 0.0532071
R15956 Iout Iout.n393 0.0532071
R15957 Iout.n330 Iout 0.0532071
R15958 Iout.n327 Iout 0.0532071
R15959 Iout.n324 Iout 0.0532071
R15960 Iout.n321 Iout 0.0532071
R15961 Iout.n318 Iout 0.0532071
R15962 Iout.n315 Iout 0.0532071
R15963 Iout.n312 Iout 0.0532071
R15964 Iout.n309 Iout 0.0532071
R15965 Iout.n306 Iout 0.0532071
R15966 Iout Iout.n459 0.0532071
R15967 Iout.n464 Iout 0.0532071
R15968 Iout.n461 Iout 0.0532071
R15969 Iout.n543 Iout 0.0532071
R15970 Iout.n137 Iout 0.0532071
R15971 Iout.n134 Iout 0.0532071
R15972 Iout.n1002 Iout 0.0532071
R15973 Iout.n537 Iout 0.0532071
R15974 Iout Iout.n535 0.0532071
R15975 Iout Iout.n532 0.0532071
R15976 Iout.n157 Iout 0.0532071
R15977 Iout.n470 Iout 0.0532071
R15978 Iout.n473 Iout 0.0532071
R15979 Iout.n190 Iout 0.0532071
R15980 Iout.n266 Iout 0.0532071
R15981 Iout Iout.n184 0.0532071
R15982 Iout.n278 Iout 0.0532071
R15983 Iout Iout.n178 0.0532071
R15984 Iout.n290 Iout 0.0532071
R15985 Iout Iout.n169 0.0532071
R15986 Iout Iout.n173 0.0532071
R15987 Iout.n296 Iout 0.0532071
R15988 Iout Iout.n175 0.0532071
R15989 Iout.n284 Iout 0.0532071
R15990 Iout Iout.n181 0.0532071
R15991 Iout.n272 Iout 0.0532071
R15992 Iout Iout.n187 0.0532071
R15993 Iout.n260 Iout 0.0532071
R15994 Iout Iout.n479 0.0532071
R15995 Iout.n484 Iout 0.0532071
R15996 Iout.n481 Iout 0.0532071
R15997 Iout.n526 Iout 0.0532071
R15998 Iout.n144 Iout 0.0532071
R15999 Iout.n141 Iout 0.0532071
R16000 Iout Iout.n1008 0.0532071
R16001 Iout.n147 Iout 0.0532071
R16002 Iout.n150 Iout 0.0532071
R16003 Iout.n520 Iout 0.0532071
R16004 Iout.n492 Iout 0.0532071
R16005 Iout.n495 Iout 0.0532071
R16006 Iout Iout.n490 0.0532071
R16007 Iout.n253 Iout 0.0532071
R16008 Iout.n256 Iout 0.0532071
R16009 Iout Iout.n251 0.0532071
R16010 Iout Iout.n248 0.0532071
R16011 Iout Iout.n245 0.0532071
R16012 Iout Iout.n242 0.0532071
R16013 Iout Iout.n239 0.0532071
R16014 Iout Iout.n236 0.0532071
R16015 Iout Iout.n233 0.0532071
R16016 Iout.n227 Iout 0.0532071
R16017 Iout.n223 Iout 0.0532071
R16018 Iout.n219 Iout 0.0532071
R16019 Iout.n215 Iout 0.0532071
R16020 Iout.n211 Iout 0.0532071
R16021 Iout.n207 Iout 0.0532071
R16022 Iout.n203 Iout 0.0532071
R16023 Iout.n200 Iout 0.0532071
R16024 Iout.n196 Iout 0.0532071
R16025 Iout.n193 Iout 0.0532071
R16026 Iout Iout.n501 0.0532071
R16027 Iout Iout.n505 0.0532071
R16028 Iout Iout.n508 0.0532071
R16029 Iout.n514 Iout 0.0532071
R16030 Iout.n510 Iout 0.0532071
R16031 Iout.n1020 Iout 0.03925
R16032 Iout.n509 Iout 0.03925
R16033 Iout.n513 Iout 0.03925
R16034 Iout.n507 Iout 0.03925
R16035 Iout.n504 Iout 0.03925
R16036 Iout.n500 Iout 0.03925
R16037 Iout.n192 Iout 0.03925
R16038 Iout.n195 Iout 0.03925
R16039 Iout.n199 Iout 0.03925
R16040 Iout.n202 Iout 0.03925
R16041 Iout.n206 Iout 0.03925
R16042 Iout.n210 Iout 0.03925
R16043 Iout.n214 Iout 0.03925
R16044 Iout.n218 Iout 0.03925
R16045 Iout.n222 Iout 0.03925
R16046 Iout.n226 Iout 0.03925
R16047 Iout.n232 Iout 0.03925
R16048 Iout.n235 Iout 0.03925
R16049 Iout.n238 Iout 0.03925
R16050 Iout.n241 Iout 0.03925
R16051 Iout.n244 Iout 0.03925
R16052 Iout.n247 Iout 0.03925
R16053 Iout.n250 Iout 0.03925
R16054 Iout.n255 Iout 0.03925
R16055 Iout.n252 Iout 0.03925
R16056 Iout.n489 Iout 0.03925
R16057 Iout.n494 Iout 0.03925
R16058 Iout.n491 Iout 0.03925
R16059 Iout.n519 Iout 0.03925
R16060 Iout.n149 Iout 0.03925
R16061 Iout.n146 Iout 0.03925
R16062 Iout.n1010 Iout 0.03925
R16063 Iout.n1007 Iout 0.03925
R16064 Iout.n140 Iout 0.03925
R16065 Iout.n143 Iout 0.03925
R16066 Iout.n525 Iout 0.03925
R16067 Iout.n480 Iout 0.03925
R16068 Iout.n483 Iout 0.03925
R16069 Iout.n478 Iout 0.03925
R16070 Iout.n259 Iout 0.03925
R16071 Iout.n186 Iout 0.03925
R16072 Iout.n271 Iout 0.03925
R16073 Iout.n180 Iout 0.03925
R16074 Iout.n283 Iout 0.03925
R16075 Iout.n174 Iout 0.03925
R16076 Iout.n168 Iout 0.03925
R16077 Iout.n301 Iout 0.03925
R16078 Iout.n289 Iout 0.03925
R16079 Iout.n177 Iout 0.03925
R16080 Iout.n277 Iout 0.03925
R16081 Iout.n183 Iout 0.03925
R16082 Iout.n265 Iout 0.03925
R16083 Iout.n189 Iout 0.03925
R16084 Iout.n472 Iout 0.03925
R16085 Iout.n469 Iout 0.03925
R16086 Iout.n156 Iout 0.03925
R16087 Iout.n531 Iout 0.03925
R16088 Iout.n534 Iout 0.03925
R16089 Iout.n536 Iout 0.03925
R16090 Iout.n133 Iout 0.03925
R16091 Iout.n136 Iout 0.03925
R16092 Iout.n542 Iout 0.03925
R16093 Iout.n460 Iout 0.03925
R16094 Iout.n463 Iout 0.03925
R16095 Iout.n458 Iout 0.03925
R16096 Iout.n305 Iout 0.03925
R16097 Iout.n308 Iout 0.03925
R16098 Iout.n311 Iout 0.03925
R16099 Iout.n314 Iout 0.03925
R16100 Iout.n317 Iout 0.03925
R16101 Iout.n320 Iout 0.03925
R16102 Iout.n392 Iout 0.03925
R16103 Iout.n378 Iout 0.03925
R16104 Iout.n376 Iout 0.03925
R16105 Iout.n394 Iout 0.03925
R16106 Iout.n408 Iout 0.03925
R16107 Iout.n410 Iout 0.03925
R16108 Iout.n424 Iout 0.03925
R16109 Iout.n426 Iout 0.03925
R16110 Iout.n447 Iout 0.03925
R16111 Iout.n452 Iout 0.03925
R16112 Iout.n449 Iout 0.03925
R16113 Iout.n548 Iout 0.03925
R16114 Iout.n130 Iout 0.03925
R16115 Iout.n559 Iout 0.03925
R16116 Iout.n557 Iout 0.03925
R16117 Iout.n554 Iout 0.03925
R16118 Iout.n434 Iout 0.03925
R16119 Iout.n438 Iout 0.03925
R16120 Iout.n441 Iout 0.03925
R16121 Iout.n432 Iout 0.03925
R16122 Iout.n418 Iout 0.03925
R16123 Iout.n416 Iout 0.03925
R16124 Iout.n402 Iout 0.03925
R16125 Iout.n357 Iout 0.03925
R16126 Iout.n360 Iout 0.03925
R16127 Iout.n363 Iout 0.03925
R16128 Iout.n366 Iout 0.03925
R16129 Iout.n354 Iout 0.03925
R16130 Iout.n351 Iout 0.03925
R16131 Iout.n348 Iout 0.03925
R16132 Iout.n345 Iout 0.03925
R16133 Iout.n342 Iout 0.03925
R16134 Iout.n339 Iout 0.03925
R16135 Iout.n336 Iout 0.03925
R16136 Iout.n333 Iout 0.03925
R16137 Iout.n117 Iout 0.03925
R16138 Iout.n582 Iout 0.03925
R16139 Iout.n111 Iout 0.03925
R16140 Iout.n594 Iout 0.03925
R16141 Iout.n105 Iout 0.03925
R16142 Iout.n606 Iout 0.03925
R16143 Iout.n99 Iout 0.03925
R16144 Iout.n618 Iout 0.03925
R16145 Iout.n624 Iout 0.03925
R16146 Iout.n90 Iout 0.03925
R16147 Iout.n636 Iout 0.03925
R16148 Iout.n81 Iout 0.03925
R16149 Iout.n648 Iout 0.03925
R16150 Iout.n96 Iout 0.03925
R16151 Iout.n612 Iout 0.03925
R16152 Iout.n102 Iout 0.03925
R16153 Iout.n600 Iout 0.03925
R16154 Iout.n108 Iout 0.03925
R16155 Iout.n588 Iout 0.03925
R16156 Iout.n687 Iout 0.03925
R16157 Iout.n684 Iout 0.03925
R16158 Iout.n681 Iout 0.03925
R16159 Iout.n678 Iout 0.03925
R16160 Iout.n675 Iout 0.03925
R16161 Iout.n672 Iout 0.03925
R16162 Iout.n747 Iout 0.03925
R16163 Iout.n50 Iout 0.03925
R16164 Iout.n759 Iout 0.03925
R16165 Iout.n44 Iout 0.03925
R16166 Iout.n771 Iout 0.03925
R16167 Iout.n42 Iout 0.03925
R16168 Iout.n56 Iout 0.03925
R16169 Iout.n735 Iout 0.03925
R16170 Iout.n62 Iout 0.03925
R16171 Iout.n723 Iout 0.03925
R16172 Iout.n717 Iout 0.03925
R16173 Iout.n65 Iout 0.03925
R16174 Iout.n729 Iout 0.03925
R16175 Iout.n59 Iout 0.03925
R16176 Iout.n805 Iout 0.03925
R16177 Iout.n808 Iout 0.03925
R16178 Iout.n811 Iout 0.03925
R16179 Iout.n814 Iout 0.03925
R16180 Iout.n817 Iout 0.03925
R16181 Iout.n820 Iout 0.03925
R16182 Iout.n823 Iout 0.03925
R16183 Iout.n802 Iout 0.03925
R16184 Iout.n799 Iout 0.03925
R16185 Iout.n890 Iout 0.03925
R16186 Iout.n888 Iout 0.03925
R16187 Iout.n881 Iout 0.03925
R16188 Iout.n869 Iout 0.03925
R16189 Iout.n867 Iout 0.03925
R16190 Iout.n855 Iout 0.03925
R16191 Iout.n853 Iout 0.03925
R16192 Iout.n841 Iout 0.03925
R16193 Iout.n839 Iout 0.03925
R16194 Iout.n827 Iout 0.03925
R16195 Iout.n883 Iout 0.03925
R16196 Iout.n895 Iout 0.03925
R16197 Iout.n897 Iout 0.03925
R16198 Iout.n909 Iout 0.03925
R16199 Iout.n911 Iout 0.03925
R16200 Iout.n923 Iout 0.03925
R16201 Iout.n926 Iout 0.03925
R16202 Iout.n22 Iout 0.03925
R16203 Iout.n876 Iout 0.03925
R16204 Iout.n874 Iout 0.03925
R16205 Iout.n862 Iout 0.03925
R16206 Iout.n860 Iout 0.03925
R16207 Iout.n848 Iout 0.03925
R16208 Iout.n846 Iout 0.03925
R16209 Iout.n834 Iout 0.03925
R16210 Iout.n832 Iout 0.03925
R16211 Iout.n902 Iout 0.03925
R16212 Iout.n904 Iout 0.03925
R16213 Iout.n916 Iout 0.03925
R16214 Iout.n918 Iout 0.03925
R16215 Iout.n931 Iout 0.03925
R16216 Iout.n934 Iout 0.03925
R16217 Iout.n796 Iout 0.03925
R16218 Iout.n793 Iout 0.03925
R16219 Iout.n790 Iout 0.03925
R16220 Iout.n787 Iout 0.03925
R16221 Iout.n784 Iout 0.03925
R16222 Iout.n781 Iout 0.03925
R16223 Iout.n938 Iout 0.03925
R16224 Iout.n741 Iout 0.03925
R16225 Iout.n53 Iout 0.03925
R16226 Iout.n753 Iout 0.03925
R16227 Iout.n47 Iout 0.03925
R16228 Iout.n765 Iout 0.03925
R16229 Iout.n38 Iout 0.03925
R16230 Iout.n777 Iout 0.03925
R16231 Iout.n71 Iout 0.03925
R16232 Iout.n705 Iout 0.03925
R16233 Iout.n77 Iout 0.03925
R16234 Iout.n944 Iout 0.03925
R16235 Iout.n19 Iout 0.03925
R16236 Iout.n68 Iout 0.03925
R16237 Iout.n711 Iout 0.03925
R16238 Iout.n74 Iout 0.03925
R16239 Iout.n699 Iout 0.03925
R16240 Iout.n950 Iout 0.03925
R16241 Iout.n953 Iout 0.03925
R16242 Iout.n669 Iout 0.03925
R16243 Iout.n666 Iout 0.03925
R16244 Iout.n663 Iout 0.03925
R16245 Iout.n660 Iout 0.03925
R16246 Iout.n657 Iout 0.03925
R16247 Iout.n654 Iout 0.03925
R16248 Iout.n690 Iout 0.03925
R16249 Iout.n695 Iout 0.03925
R16250 Iout.n692 Iout 0.03925
R16251 Iout.n957 Iout 0.03925
R16252 Iout.n114 Iout 0.03925
R16253 Iout.n576 Iout 0.03925
R16254 Iout.n573 Iout 0.03925
R16255 Iout.n963 Iout 0.03925
R16256 Iout.n14 Iout 0.03925
R16257 Iout.n93 Iout 0.03925
R16258 Iout.n630 Iout 0.03925
R16259 Iout.n87 Iout 0.03925
R16260 Iout.n642 Iout 0.03925
R16261 Iout.n85 Iout 0.03925
R16262 Iout.n563 Iout 0.03925
R16263 Iout.n969 Iout 0.03925
R16264 Iout.n972 Iout 0.03925
R16265 Iout.n569 Iout 0.03925
R16266 Iout.n123 Iout 0.03925
R16267 Iout.n120 Iout 0.03925
R16268 Iout.n976 Iout 0.03925
R16269 Iout.n400 Iout 0.03925
R16270 Iout.n386 Iout 0.03925
R16271 Iout.n384 Iout 0.03925
R16272 Iout.n370 Iout 0.03925
R16273 Iout.n982 Iout 0.03925
R16274 Iout.n9 Iout 0.03925
R16275 Iout.n127 Iout 0.03925
R16276 Iout.n988 Iout 0.03925
R16277 Iout.n991 Iout 0.03925
R16278 Iout.n323 Iout 0.03925
R16279 Iout.n326 Iout 0.03925
R16280 Iout.n329 Iout 0.03925
R16281 Iout.n995 Iout 0.03925
R16282 Iout.n1001 Iout 0.03925
R16283 Iout.n4 Iout 0.03925
R16284 Iout.n295 Iout 0.03925
R16285 Iout.n172 Iout 0.03925
R16286 Iout.n1014 Iout 0.03925
R16287 Iout.n1022 Iout 0.02071
R16288 Iout Iout.n1022 0.00379
R16289 Iout.n303 Iout.n302 0.00105952
R16290 Iout.n377 Iout.n375 0.00105952
R16291 Iout.n380 Iout.n379 0.00105952
R16292 Iout.n368 Iout.n367 0.00105952
R16293 Iout.n365 Iout.n364 0.00105952
R16294 Iout.n362 Iout.n361 0.00105952
R16295 Iout.n650 Iout.n649 0.00105952
R16296 Iout.n647 Iout.n82 0.00105952
R16297 Iout.n638 Iout.n637 0.00105952
R16298 Iout.n635 Iout.n91 0.00105952
R16299 Iout.n43 Iout.n41 0.00105952
R16300 Iout.n773 Iout.n772 0.00105952
R16301 Iout.n770 Iout.n45 0.00105952
R16302 Iout.n761 Iout.n760 0.00105952
R16303 Iout.n758 Iout.n51 0.00105952
R16304 Iout.n825 Iout.n824 0.00105952
R16305 Iout.n822 Iout.n821 0.00105952
R16306 Iout.n819 Iout.n818 0.00105952
R16307 Iout.n816 Iout.n815 0.00105952
R16308 Iout.n813 Iout.n812 0.00105952
R16309 Iout.n810 Iout.n809 0.00105952
R16310 Iout.n829 Iout.n828 0.00105952
R16311 Iout.n840 Iout.n838 0.00105952
R16312 Iout.n843 Iout.n842 0.00105952
R16313 Iout.n854 Iout.n852 0.00105952
R16314 Iout.n857 Iout.n856 0.00105952
R16315 Iout.n868 Iout.n866 0.00105952
R16316 Iout.n871 Iout.n870 0.00105952
R16317 Iout.n925 Iout.n23 0.00105952
R16318 Iout.n928 Iout.n927 0.00105952
R16319 Iout.n924 Iout.n922 0.00105952
R16320 Iout.n913 Iout.n912 0.00105952
R16321 Iout.n910 Iout.n908 0.00105952
R16322 Iout.n899 Iout.n898 0.00105952
R16323 Iout.n896 Iout.n894 0.00105952
R16324 Iout.n885 Iout.n884 0.00105952
R16325 Iout.n882 Iout.n880 0.00105952
R16326 Iout.n833 Iout.n831 0.00105952
R16327 Iout.n836 Iout.n835 0.00105952
R16328 Iout.n847 Iout.n845 0.00105952
R16329 Iout.n850 Iout.n849 0.00105952
R16330 Iout.n861 Iout.n859 0.00105952
R16331 Iout.n864 Iout.n863 0.00105952
R16332 Iout.n875 Iout.n873 0.00105952
R16333 Iout.n878 Iout.n877 0.00105952
R16334 Iout.n889 Iout.n887 0.00105952
R16335 Iout.n935 Iout.n933 0.00105952
R16336 Iout.n932 Iout.n930 0.00105952
R16337 Iout.n920 Iout.n919 0.00105952
R16338 Iout.n917 Iout.n915 0.00105952
R16339 Iout.n906 Iout.n905 0.00105952
R16340 Iout.n903 Iout.n901 0.00105952
R16341 Iout.n892 Iout.n891 0.00105952
R16342 Iout.n940 Iout.n939 0.00105952
R16343 Iout.n783 Iout.n782 0.00105952
R16344 Iout.n786 Iout.n785 0.00105952
R16345 Iout.n789 Iout.n788 0.00105952
R16346 Iout.n792 Iout.n791 0.00105952
R16347 Iout.n795 Iout.n794 0.00105952
R16348 Iout.n798 Iout.n797 0.00105952
R16349 Iout.n801 Iout.n800 0.00105952
R16350 Iout.n804 Iout.n803 0.00105952
R16351 Iout.n807 Iout.n806 0.00105952
R16352 Iout.n779 Iout.n778 0.00105952
R16353 Iout.n776 Iout.n39 0.00105952
R16354 Iout.n767 Iout.n766 0.00105952
R16355 Iout.n764 Iout.n48 0.00105952
R16356 Iout.n755 Iout.n754 0.00105952
R16357 Iout.n752 Iout.n54 0.00105952
R16358 Iout.n743 Iout.n742 0.00105952
R16359 Iout.n740 Iout.n60 0.00105952
R16360 Iout.n731 Iout.n730 0.00105952
R16361 Iout.n728 Iout.n66 0.00105952
R16362 Iout.n943 Iout.n20 0.00105952
R16363 Iout.n946 Iout.n945 0.00105952
R16364 Iout.n704 Iout.n78 0.00105952
R16365 Iout.n707 Iout.n706 0.00105952
R16366 Iout.n716 Iout.n72 0.00105952
R16367 Iout.n719 Iout.n718 0.00105952
R16368 Iout.n954 Iout.n952 0.00105952
R16369 Iout.n951 Iout.n949 0.00105952
R16370 Iout.n701 Iout.n700 0.00105952
R16371 Iout.n710 Iout.n75 0.00105952
R16372 Iout.n713 Iout.n712 0.00105952
R16373 Iout.n722 Iout.n69 0.00105952
R16374 Iout.n725 Iout.n724 0.00105952
R16375 Iout.n734 Iout.n63 0.00105952
R16376 Iout.n737 Iout.n736 0.00105952
R16377 Iout.n746 Iout.n57 0.00105952
R16378 Iout.n749 Iout.n748 0.00105952
R16379 Iout.n655 Iout.n653 0.00105952
R16380 Iout.n658 Iout.n656 0.00105952
R16381 Iout.n661 Iout.n659 0.00105952
R16382 Iout.n664 Iout.n662 0.00105952
R16383 Iout.n667 Iout.n665 0.00105952
R16384 Iout.n670 Iout.n668 0.00105952
R16385 Iout.n673 Iout.n671 0.00105952
R16386 Iout.n676 Iout.n674 0.00105952
R16387 Iout.n679 Iout.n677 0.00105952
R16388 Iout.n682 Iout.n680 0.00105952
R16389 Iout.n685 Iout.n683 0.00105952
R16390 Iout.n959 Iout.n958 0.00105952
R16391 Iout.n694 Iout.n693 0.00105952
R16392 Iout.n697 Iout.n696 0.00105952
R16393 Iout.n691 Iout.n689 0.00105952
R16394 Iout.n688 Iout.n686 0.00105952
R16395 Iout.n962 Iout.n15 0.00105952
R16396 Iout.n965 Iout.n964 0.00105952
R16397 Iout.n575 Iout.n574 0.00105952
R16398 Iout.n578 Iout.n577 0.00105952
R16399 Iout.n587 Iout.n115 0.00105952
R16400 Iout.n590 Iout.n589 0.00105952
R16401 Iout.n599 Iout.n109 0.00105952
R16402 Iout.n602 Iout.n601 0.00105952
R16403 Iout.n611 Iout.n103 0.00105952
R16404 Iout.n614 Iout.n613 0.00105952
R16405 Iout.n623 Iout.n97 0.00105952
R16406 Iout.n626 Iout.n625 0.00105952
R16407 Iout.n86 Iout.n84 0.00105952
R16408 Iout.n644 Iout.n643 0.00105952
R16409 Iout.n641 Iout.n88 0.00105952
R16410 Iout.n632 Iout.n631 0.00105952
R16411 Iout.n629 Iout.n94 0.00105952
R16412 Iout.n620 Iout.n619 0.00105952
R16413 Iout.n617 Iout.n100 0.00105952
R16414 Iout.n608 Iout.n607 0.00105952
R16415 Iout.n605 Iout.n106 0.00105952
R16416 Iout.n596 Iout.n595 0.00105952
R16417 Iout.n593 Iout.n112 0.00105952
R16418 Iout.n584 Iout.n583 0.00105952
R16419 Iout.n973 Iout.n971 0.00105952
R16420 Iout.n970 Iout.n968 0.00105952
R16421 Iout.n565 Iout.n564 0.00105952
R16422 Iout.n581 Iout.n118 0.00105952
R16423 Iout.n978 Iout.n977 0.00105952
R16424 Iout.n122 Iout.n121 0.00105952
R16425 Iout.n568 Iout.n124 0.00105952
R16426 Iout.n571 Iout.n570 0.00105952
R16427 Iout.n335 Iout.n334 0.00105952
R16428 Iout.n338 Iout.n337 0.00105952
R16429 Iout.n341 Iout.n340 0.00105952
R16430 Iout.n344 Iout.n343 0.00105952
R16431 Iout.n347 Iout.n346 0.00105952
R16432 Iout.n350 Iout.n349 0.00105952
R16433 Iout.n353 Iout.n352 0.00105952
R16434 Iout.n356 Iout.n355 0.00105952
R16435 Iout.n359 Iout.n358 0.00105952
R16436 Iout.n372 Iout.n371 0.00105952
R16437 Iout.n385 Iout.n383 0.00105952
R16438 Iout.n388 Iout.n387 0.00105952
R16439 Iout.n401 Iout.n399 0.00105952
R16440 Iout.n404 Iout.n403 0.00105952
R16441 Iout.n417 Iout.n415 0.00105952
R16442 Iout.n420 Iout.n419 0.00105952
R16443 Iout.n433 Iout.n431 0.00105952
R16444 Iout.n443 Iout.n442 0.00105952
R16445 Iout.n440 Iout.n439 0.00105952
R16446 Iout.n437 Iout.n435 0.00105952
R16447 Iout.n555 Iout.n553 0.00105952
R16448 Iout.n558 Iout.n556 0.00105952
R16449 Iout.n981 Iout.n10 0.00105952
R16450 Iout.n984 Iout.n983 0.00105952
R16451 Iout.n561 Iout.n560 0.00105952
R16452 Iout.n992 Iout.n990 0.00105952
R16453 Iout.n989 Iout.n987 0.00105952
R16454 Iout.n129 Iout.n128 0.00105952
R16455 Iout.n547 Iout.n131 0.00105952
R16456 Iout.n550 Iout.n549 0.00105952
R16457 Iout.n451 Iout.n450 0.00105952
R16458 Iout.n454 Iout.n453 0.00105952
R16459 Iout.n448 Iout.n446 0.00105952
R16460 Iout.n428 Iout.n427 0.00105952
R16461 Iout.n425 Iout.n423 0.00105952
R16462 Iout.n412 Iout.n411 0.00105952
R16463 Iout.n409 Iout.n407 0.00105952
R16464 Iout.n396 Iout.n395 0.00105952
R16465 Iout.n393 Iout.n391 0.00105952
R16466 Iout.n331 Iout.n330 0.00105952
R16467 Iout.n328 Iout.n327 0.00105952
R16468 Iout.n325 Iout.n324 0.00105952
R16469 Iout.n322 Iout.n321 0.00105952
R16470 Iout.n319 Iout.n318 0.00105952
R16471 Iout.n316 Iout.n315 0.00105952
R16472 Iout.n313 Iout.n312 0.00105952
R16473 Iout.n310 Iout.n309 0.00105952
R16474 Iout.n307 Iout.n306 0.00105952
R16475 Iout.n459 Iout.n457 0.00105952
R16476 Iout.n465 Iout.n464 0.00105952
R16477 Iout.n462 Iout.n461 0.00105952
R16478 Iout.n544 Iout.n543 0.00105952
R16479 Iout.n541 Iout.n137 0.00105952
R16480 Iout.n997 Iout.n996 0.00105952
R16481 Iout.n135 Iout.n134 0.00105952
R16482 Iout.n1000 Iout.n5 0.00105952
R16483 Iout.n1003 Iout.n1002 0.00105952
R16484 Iout.n538 Iout.n537 0.00105952
R16485 Iout.n535 Iout.n533 0.00105952
R16486 Iout.n532 Iout.n530 0.00105952
R16487 Iout.n468 Iout.n157 0.00105952
R16488 Iout.n471 Iout.n470 0.00105952
R16489 Iout.n474 Iout.n473 0.00105952
R16490 Iout.n264 Iout.n190 0.00105952
R16491 Iout.n267 Iout.n266 0.00105952
R16492 Iout.n276 Iout.n184 0.00105952
R16493 Iout.n279 Iout.n278 0.00105952
R16494 Iout.n288 Iout.n178 0.00105952
R16495 Iout.n291 Iout.n290 0.00105952
R16496 Iout.n300 Iout.n169 0.00105952
R16497 Iout.n173 Iout.n171 0.00105952
R16498 Iout.n297 Iout.n296 0.00105952
R16499 Iout.n294 Iout.n175 0.00105952
R16500 Iout.n285 Iout.n284 0.00105952
R16501 Iout.n282 Iout.n181 0.00105952
R16502 Iout.n273 Iout.n272 0.00105952
R16503 Iout.n270 Iout.n187 0.00105952
R16504 Iout.n261 Iout.n260 0.00105952
R16505 Iout.n479 Iout.n477 0.00105952
R16506 Iout.n485 Iout.n484 0.00105952
R16507 Iout.n482 Iout.n481 0.00105952
R16508 Iout.n527 Iout.n526 0.00105952
R16509 Iout.n524 Iout.n144 0.00105952
R16510 Iout.n142 Iout.n141 0.00105952
R16511 Iout.n1008 Iout.n1006 0.00105952
R16512 Iout.n1011 Iout.n1009 0.00105952
R16513 Iout.n1016 Iout.n1015 0.00105952
R16514 Iout.n148 Iout.n147 0.00105952
R16515 Iout.n518 Iout.n150 0.00105952
R16516 Iout.n521 Iout.n520 0.00105952
R16517 Iout.n493 Iout.n492 0.00105952
R16518 Iout.n496 Iout.n495 0.00105952
R16519 Iout.n490 Iout.n488 0.00105952
R16520 Iout.n254 Iout.n253 0.00105952
R16521 Iout.n257 Iout.n256 0.00105952
R16522 Iout.n251 Iout.n249 0.00105952
R16523 Iout.n248 Iout.n246 0.00105952
R16524 Iout.n245 Iout.n243 0.00105952
R16525 Iout.n242 Iout.n240 0.00105952
R16526 Iout.n239 Iout.n237 0.00105952
R16527 Iout.n236 Iout.n234 0.00105952
R16528 Iout.n233 Iout.n231 0.00105952
R16529 Iout.n228 Iout.n227 0.00105952
R16530 Iout.n225 Iout.n223 0.00105952
R16531 Iout.n221 Iout.n219 0.00105952
R16532 Iout.n217 Iout.n215 0.00105952
R16533 Iout.n213 Iout.n211 0.00105952
R16534 Iout.n209 Iout.n207 0.00105952
R16535 Iout.n205 Iout.n203 0.00105952
R16536 Iout.n201 Iout.n200 0.00105952
R16537 Iout.n198 Iout.n196 0.00105952
R16538 Iout.n194 Iout.n193 0.00105952
R16539 Iout.n501 Iout.n499 0.00105952
R16540 Iout.n505 Iout.n503 0.00105952
R16541 Iout.n508 Iout.n506 0.00105952
R16542 Iout.n515 Iout.n514 0.00105952
R16543 Iout.n512 Iout.n510 0.00105952
R16544 Iout.n1021 Iout.n1019 0.00105952
R16545 XA.Cn[10].n55 XA.Cn[10].n54 256.104
R16546 XA.Cn[10].n59 XA.Cn[10].n58 243.679
R16547 XA.Cn[10].n2 XA.Cn[10].n0 241.847
R16548 XA.Cn[10].n59 XA.Cn[10].n57 205.28
R16549 XA.Cn[10].n55 XA.Cn[10].n53 202.095
R16550 XA.Cn[10].n2 XA.Cn[10].n1 185
R16551 XA.Cn[10].n5 XA.Cn[10].n3 161.406
R16552 XA.Cn[10].n8 XA.Cn[10].n6 161.406
R16553 XA.Cn[10].n11 XA.Cn[10].n9 161.406
R16554 XA.Cn[10].n14 XA.Cn[10].n12 161.406
R16555 XA.Cn[10].n17 XA.Cn[10].n15 161.406
R16556 XA.Cn[10].n20 XA.Cn[10].n18 161.406
R16557 XA.Cn[10].n23 XA.Cn[10].n21 161.406
R16558 XA.Cn[10].n26 XA.Cn[10].n24 161.406
R16559 XA.Cn[10].n29 XA.Cn[10].n27 161.406
R16560 XA.Cn[10].n32 XA.Cn[10].n30 161.406
R16561 XA.Cn[10].n35 XA.Cn[10].n33 161.406
R16562 XA.Cn[10].n38 XA.Cn[10].n36 161.406
R16563 XA.Cn[10].n41 XA.Cn[10].n39 161.406
R16564 XA.Cn[10].n44 XA.Cn[10].n42 161.406
R16565 XA.Cn[10].n47 XA.Cn[10].n45 161.406
R16566 XA.Cn[10].n50 XA.Cn[10].n48 161.406
R16567 XA.Cn[10].n3 XA.Cn[10].t36 161.202
R16568 XA.Cn[10].n6 XA.Cn[10].t21 161.202
R16569 XA.Cn[10].n9 XA.Cn[10].t23 161.202
R16570 XA.Cn[10].n12 XA.Cn[10].t25 161.202
R16571 XA.Cn[10].n15 XA.Cn[10].t14 161.202
R16572 XA.Cn[10].n18 XA.Cn[10].t15 161.202
R16573 XA.Cn[10].n21 XA.Cn[10].t28 161.202
R16574 XA.Cn[10].n24 XA.Cn[10].t37 161.202
R16575 XA.Cn[10].n27 XA.Cn[10].t39 161.202
R16576 XA.Cn[10].n30 XA.Cn[10].t26 161.202
R16577 XA.Cn[10].n33 XA.Cn[10].t27 161.202
R16578 XA.Cn[10].n36 XA.Cn[10].t40 161.202
R16579 XA.Cn[10].n39 XA.Cn[10].t16 161.202
R16580 XA.Cn[10].n42 XA.Cn[10].t19 161.202
R16581 XA.Cn[10].n45 XA.Cn[10].t32 161.202
R16582 XA.Cn[10].n48 XA.Cn[10].t42 161.202
R16583 XA.Cn[10].n3 XA.Cn[10].t38 145.137
R16584 XA.Cn[10].n6 XA.Cn[10].t24 145.137
R16585 XA.Cn[10].n9 XA.Cn[10].t29 145.137
R16586 XA.Cn[10].n12 XA.Cn[10].t30 145.137
R16587 XA.Cn[10].n15 XA.Cn[10].t17 145.137
R16588 XA.Cn[10].n18 XA.Cn[10].t18 145.137
R16589 XA.Cn[10].n21 XA.Cn[10].t34 145.137
R16590 XA.Cn[10].n24 XA.Cn[10].t41 145.137
R16591 XA.Cn[10].n27 XA.Cn[10].t43 145.137
R16592 XA.Cn[10].n30 XA.Cn[10].t31 145.137
R16593 XA.Cn[10].n33 XA.Cn[10].t33 145.137
R16594 XA.Cn[10].n36 XA.Cn[10].t12 145.137
R16595 XA.Cn[10].n39 XA.Cn[10].t20 145.137
R16596 XA.Cn[10].n42 XA.Cn[10].t22 145.137
R16597 XA.Cn[10].n45 XA.Cn[10].t35 145.137
R16598 XA.Cn[10].n48 XA.Cn[10].t13 145.137
R16599 XA.Cn[10].n53 XA.Cn[10].t2 26.5955
R16600 XA.Cn[10].n53 XA.Cn[10].t8 26.5955
R16601 XA.Cn[10].n54 XA.Cn[10].t9 26.5955
R16602 XA.Cn[10].n54 XA.Cn[10].t1 26.5955
R16603 XA.Cn[10].n57 XA.Cn[10].t5 26.5955
R16604 XA.Cn[10].n57 XA.Cn[10].t4 26.5955
R16605 XA.Cn[10].n58 XA.Cn[10].t11 26.5955
R16606 XA.Cn[10].n58 XA.Cn[10].t0 26.5955
R16607 XA.Cn[10].n1 XA.Cn[10].t10 24.9236
R16608 XA.Cn[10].n1 XA.Cn[10].t7 24.9236
R16609 XA.Cn[10].n0 XA.Cn[10].t6 24.9236
R16610 XA.Cn[10].n0 XA.Cn[10].t3 24.9236
R16611 XA.Cn[10] XA.Cn[10].n59 22.9652
R16612 XA.Cn[10] XA.Cn[10].n2 22.9615
R16613 XA.Cn[10].n56 XA.Cn[10].n55 13.9299
R16614 XA.Cn[10] XA.Cn[10].n56 13.9299
R16615 XA.Cn[10].n52 XA.Cn[10].n51 5.13256
R16616 XA.Cn[10].n56 XA.Cn[10].n52 2.99115
R16617 XA.Cn[10].n56 XA.Cn[10] 2.87153
R16618 XA.Cn[10].n52 XA.Cn[10] 2.2734
R16619 XA.Cn[10].n51 XA.Cn[10] 2.26343
R16620 XA.Cn[10].n8 XA.Cn[10] 0.931056
R16621 XA.Cn[10].n11 XA.Cn[10] 0.931056
R16622 XA.Cn[10].n14 XA.Cn[10] 0.931056
R16623 XA.Cn[10].n17 XA.Cn[10] 0.931056
R16624 XA.Cn[10].n20 XA.Cn[10] 0.931056
R16625 XA.Cn[10].n23 XA.Cn[10] 0.931056
R16626 XA.Cn[10].n26 XA.Cn[10] 0.931056
R16627 XA.Cn[10].n29 XA.Cn[10] 0.931056
R16628 XA.Cn[10].n32 XA.Cn[10] 0.931056
R16629 XA.Cn[10].n35 XA.Cn[10] 0.931056
R16630 XA.Cn[10].n38 XA.Cn[10] 0.931056
R16631 XA.Cn[10].n41 XA.Cn[10] 0.931056
R16632 XA.Cn[10].n44 XA.Cn[10] 0.931056
R16633 XA.Cn[10].n47 XA.Cn[10] 0.931056
R16634 XA.Cn[10].n50 XA.Cn[10] 0.931056
R16635 XA.Cn[10] XA.Cn[10].n5 0.396333
R16636 XA.Cn[10] XA.Cn[10].n8 0.396333
R16637 XA.Cn[10] XA.Cn[10].n11 0.396333
R16638 XA.Cn[10] XA.Cn[10].n14 0.396333
R16639 XA.Cn[10] XA.Cn[10].n17 0.396333
R16640 XA.Cn[10] XA.Cn[10].n20 0.396333
R16641 XA.Cn[10] XA.Cn[10].n23 0.396333
R16642 XA.Cn[10] XA.Cn[10].n26 0.396333
R16643 XA.Cn[10] XA.Cn[10].n29 0.396333
R16644 XA.Cn[10] XA.Cn[10].n32 0.396333
R16645 XA.Cn[10] XA.Cn[10].n35 0.396333
R16646 XA.Cn[10] XA.Cn[10].n38 0.396333
R16647 XA.Cn[10] XA.Cn[10].n41 0.396333
R16648 XA.Cn[10] XA.Cn[10].n44 0.396333
R16649 XA.Cn[10] XA.Cn[10].n47 0.396333
R16650 XA.Cn[10] XA.Cn[10].n50 0.396333
R16651 XA.Cn[10].n4 XA.Cn[10] 0.104667
R16652 XA.Cn[10].n7 XA.Cn[10] 0.104667
R16653 XA.Cn[10].n10 XA.Cn[10] 0.104667
R16654 XA.Cn[10].n13 XA.Cn[10] 0.104667
R16655 XA.Cn[10].n16 XA.Cn[10] 0.104667
R16656 XA.Cn[10].n19 XA.Cn[10] 0.104667
R16657 XA.Cn[10].n22 XA.Cn[10] 0.104667
R16658 XA.Cn[10].n25 XA.Cn[10] 0.104667
R16659 XA.Cn[10].n28 XA.Cn[10] 0.104667
R16660 XA.Cn[10].n31 XA.Cn[10] 0.104667
R16661 XA.Cn[10].n34 XA.Cn[10] 0.104667
R16662 XA.Cn[10].n37 XA.Cn[10] 0.104667
R16663 XA.Cn[10].n40 XA.Cn[10] 0.104667
R16664 XA.Cn[10].n43 XA.Cn[10] 0.104667
R16665 XA.Cn[10].n46 XA.Cn[10] 0.104667
R16666 XA.Cn[10].n49 XA.Cn[10] 0.104667
R16667 XA.Cn[10].n4 XA.Cn[10] 0.0309878
R16668 XA.Cn[10].n7 XA.Cn[10] 0.0309878
R16669 XA.Cn[10].n10 XA.Cn[10] 0.0309878
R16670 XA.Cn[10].n13 XA.Cn[10] 0.0309878
R16671 XA.Cn[10].n16 XA.Cn[10] 0.0309878
R16672 XA.Cn[10].n19 XA.Cn[10] 0.0309878
R16673 XA.Cn[10].n22 XA.Cn[10] 0.0309878
R16674 XA.Cn[10].n25 XA.Cn[10] 0.0309878
R16675 XA.Cn[10].n28 XA.Cn[10] 0.0309878
R16676 XA.Cn[10].n31 XA.Cn[10] 0.0309878
R16677 XA.Cn[10].n34 XA.Cn[10] 0.0309878
R16678 XA.Cn[10].n37 XA.Cn[10] 0.0309878
R16679 XA.Cn[10].n40 XA.Cn[10] 0.0309878
R16680 XA.Cn[10].n43 XA.Cn[10] 0.0309878
R16681 XA.Cn[10].n46 XA.Cn[10] 0.0309878
R16682 XA.Cn[10].n49 XA.Cn[10] 0.0309878
R16683 XA.Cn[10].n5 XA.Cn[10].n4 0.027939
R16684 XA.Cn[10].n8 XA.Cn[10].n7 0.027939
R16685 XA.Cn[10].n11 XA.Cn[10].n10 0.027939
R16686 XA.Cn[10].n14 XA.Cn[10].n13 0.027939
R16687 XA.Cn[10].n17 XA.Cn[10].n16 0.027939
R16688 XA.Cn[10].n20 XA.Cn[10].n19 0.027939
R16689 XA.Cn[10].n23 XA.Cn[10].n22 0.027939
R16690 XA.Cn[10].n26 XA.Cn[10].n25 0.027939
R16691 XA.Cn[10].n29 XA.Cn[10].n28 0.027939
R16692 XA.Cn[10].n32 XA.Cn[10].n31 0.027939
R16693 XA.Cn[10].n35 XA.Cn[10].n34 0.027939
R16694 XA.Cn[10].n38 XA.Cn[10].n37 0.027939
R16695 XA.Cn[10].n41 XA.Cn[10].n40 0.027939
R16696 XA.Cn[10].n44 XA.Cn[10].n43 0.027939
R16697 XA.Cn[10].n47 XA.Cn[10].n46 0.027939
R16698 XA.Cn[10].n50 XA.Cn[10].n49 0.027939
R16699 XA.Cn[10].n51 XA.Cn[10] 0.00285068
R16700 XThR.Tn[6].n2 XThR.Tn[6].n1 332.332
R16701 XThR.Tn[6].n2 XThR.Tn[6].n0 296.493
R16702 XThR.Tn[6] XThR.Tn[6].n82 161.363
R16703 XThR.Tn[6] XThR.Tn[6].n77 161.363
R16704 XThR.Tn[6] XThR.Tn[6].n72 161.363
R16705 XThR.Tn[6] XThR.Tn[6].n67 161.363
R16706 XThR.Tn[6] XThR.Tn[6].n62 161.363
R16707 XThR.Tn[6] XThR.Tn[6].n57 161.363
R16708 XThR.Tn[6] XThR.Tn[6].n52 161.363
R16709 XThR.Tn[6] XThR.Tn[6].n47 161.363
R16710 XThR.Tn[6] XThR.Tn[6].n42 161.363
R16711 XThR.Tn[6] XThR.Tn[6].n37 161.363
R16712 XThR.Tn[6] XThR.Tn[6].n32 161.363
R16713 XThR.Tn[6] XThR.Tn[6].n27 161.363
R16714 XThR.Tn[6] XThR.Tn[6].n22 161.363
R16715 XThR.Tn[6] XThR.Tn[6].n17 161.363
R16716 XThR.Tn[6] XThR.Tn[6].n12 161.363
R16717 XThR.Tn[6] XThR.Tn[6].n10 161.363
R16718 XThR.Tn[6].n84 XThR.Tn[6].n83 161.3
R16719 XThR.Tn[6].n79 XThR.Tn[6].n78 161.3
R16720 XThR.Tn[6].n74 XThR.Tn[6].n73 161.3
R16721 XThR.Tn[6].n69 XThR.Tn[6].n68 161.3
R16722 XThR.Tn[6].n64 XThR.Tn[6].n63 161.3
R16723 XThR.Tn[6].n59 XThR.Tn[6].n58 161.3
R16724 XThR.Tn[6].n54 XThR.Tn[6].n53 161.3
R16725 XThR.Tn[6].n49 XThR.Tn[6].n48 161.3
R16726 XThR.Tn[6].n44 XThR.Tn[6].n43 161.3
R16727 XThR.Tn[6].n39 XThR.Tn[6].n38 161.3
R16728 XThR.Tn[6].n34 XThR.Tn[6].n33 161.3
R16729 XThR.Tn[6].n29 XThR.Tn[6].n28 161.3
R16730 XThR.Tn[6].n24 XThR.Tn[6].n23 161.3
R16731 XThR.Tn[6].n19 XThR.Tn[6].n18 161.3
R16732 XThR.Tn[6].n14 XThR.Tn[6].n13 161.3
R16733 XThR.Tn[6].n82 XThR.Tn[6].t46 161.106
R16734 XThR.Tn[6].n77 XThR.Tn[6].t52 161.106
R16735 XThR.Tn[6].n72 XThR.Tn[6].t32 161.106
R16736 XThR.Tn[6].n67 XThR.Tn[6].t18 161.106
R16737 XThR.Tn[6].n62 XThR.Tn[6].t44 161.106
R16738 XThR.Tn[6].n57 XThR.Tn[6].t69 161.106
R16739 XThR.Tn[6].n52 XThR.Tn[6].t50 161.106
R16740 XThR.Tn[6].n47 XThR.Tn[6].t30 161.106
R16741 XThR.Tn[6].n42 XThR.Tn[6].t17 161.106
R16742 XThR.Tn[6].n37 XThR.Tn[6].t22 161.106
R16743 XThR.Tn[6].n32 XThR.Tn[6].t67 161.106
R16744 XThR.Tn[6].n27 XThR.Tn[6].t31 161.106
R16745 XThR.Tn[6].n22 XThR.Tn[6].t66 161.106
R16746 XThR.Tn[6].n17 XThR.Tn[6].t49 161.106
R16747 XThR.Tn[6].n12 XThR.Tn[6].t72 161.106
R16748 XThR.Tn[6].n10 XThR.Tn[6].t56 161.106
R16749 XThR.Tn[6].n83 XThR.Tn[6].t42 159.978
R16750 XThR.Tn[6].n78 XThR.Tn[6].t48 159.978
R16751 XThR.Tn[6].n73 XThR.Tn[6].t28 159.978
R16752 XThR.Tn[6].n68 XThR.Tn[6].t15 159.978
R16753 XThR.Tn[6].n63 XThR.Tn[6].t39 159.978
R16754 XThR.Tn[6].n58 XThR.Tn[6].t65 159.978
R16755 XThR.Tn[6].n53 XThR.Tn[6].t47 159.978
R16756 XThR.Tn[6].n48 XThR.Tn[6].t25 159.978
R16757 XThR.Tn[6].n43 XThR.Tn[6].t12 159.978
R16758 XThR.Tn[6].n38 XThR.Tn[6].t19 159.978
R16759 XThR.Tn[6].n33 XThR.Tn[6].t64 159.978
R16760 XThR.Tn[6].n28 XThR.Tn[6].t27 159.978
R16761 XThR.Tn[6].n23 XThR.Tn[6].t63 159.978
R16762 XThR.Tn[6].n18 XThR.Tn[6].t45 159.978
R16763 XThR.Tn[6].n13 XThR.Tn[6].t68 159.978
R16764 XThR.Tn[6].n82 XThR.Tn[6].t34 145.038
R16765 XThR.Tn[6].n77 XThR.Tn[6].t58 145.038
R16766 XThR.Tn[6].n72 XThR.Tn[6].t38 145.038
R16767 XThR.Tn[6].n67 XThR.Tn[6].t23 145.038
R16768 XThR.Tn[6].n62 XThR.Tn[6].t53 145.038
R16769 XThR.Tn[6].n57 XThR.Tn[6].t33 145.038
R16770 XThR.Tn[6].n52 XThR.Tn[6].t40 145.038
R16771 XThR.Tn[6].n47 XThR.Tn[6].t24 145.038
R16772 XThR.Tn[6].n42 XThR.Tn[6].t21 145.038
R16773 XThR.Tn[6].n37 XThR.Tn[6].t51 145.038
R16774 XThR.Tn[6].n32 XThR.Tn[6].t13 145.038
R16775 XThR.Tn[6].n27 XThR.Tn[6].t35 145.038
R16776 XThR.Tn[6].n22 XThR.Tn[6].t73 145.038
R16777 XThR.Tn[6].n17 XThR.Tn[6].t57 145.038
R16778 XThR.Tn[6].n12 XThR.Tn[6].t20 145.038
R16779 XThR.Tn[6].n10 XThR.Tn[6].t62 145.038
R16780 XThR.Tn[6].n83 XThR.Tn[6].t55 143.911
R16781 XThR.Tn[6].n78 XThR.Tn[6].t16 143.911
R16782 XThR.Tn[6].n73 XThR.Tn[6].t60 143.911
R16783 XThR.Tn[6].n68 XThR.Tn[6].t41 143.911
R16784 XThR.Tn[6].n63 XThR.Tn[6].t71 143.911
R16785 XThR.Tn[6].n58 XThR.Tn[6].t54 143.911
R16786 XThR.Tn[6].n53 XThR.Tn[6].t61 143.911
R16787 XThR.Tn[6].n48 XThR.Tn[6].t43 143.911
R16788 XThR.Tn[6].n43 XThR.Tn[6].t37 143.911
R16789 XThR.Tn[6].n38 XThR.Tn[6].t70 143.911
R16790 XThR.Tn[6].n33 XThR.Tn[6].t29 143.911
R16791 XThR.Tn[6].n28 XThR.Tn[6].t59 143.911
R16792 XThR.Tn[6].n23 XThR.Tn[6].t26 143.911
R16793 XThR.Tn[6].n18 XThR.Tn[6].t14 143.911
R16794 XThR.Tn[6].n13 XThR.Tn[6].t36 143.911
R16795 XThR.Tn[6].n7 XThR.Tn[6].n5 135.249
R16796 XThR.Tn[6].n9 XThR.Tn[6].n3 98.982
R16797 XThR.Tn[6].n8 XThR.Tn[6].n4 98.982
R16798 XThR.Tn[6].n7 XThR.Tn[6].n6 98.982
R16799 XThR.Tn[6].n9 XThR.Tn[6].n8 36.2672
R16800 XThR.Tn[6].n8 XThR.Tn[6].n7 36.2672
R16801 XThR.Tn[6].n88 XThR.Tn[6].n9 32.6405
R16802 XThR.Tn[6].n1 XThR.Tn[6].t6 26.5955
R16803 XThR.Tn[6].n1 XThR.Tn[6].t5 26.5955
R16804 XThR.Tn[6].n0 XThR.Tn[6].t7 26.5955
R16805 XThR.Tn[6].n0 XThR.Tn[6].t4 26.5955
R16806 XThR.Tn[6].n3 XThR.Tn[6].t8 24.9236
R16807 XThR.Tn[6].n3 XThR.Tn[6].t9 24.9236
R16808 XThR.Tn[6].n4 XThR.Tn[6].t11 24.9236
R16809 XThR.Tn[6].n4 XThR.Tn[6].t10 24.9236
R16810 XThR.Tn[6].n5 XThR.Tn[6].t0 24.9236
R16811 XThR.Tn[6].n5 XThR.Tn[6].t1 24.9236
R16812 XThR.Tn[6].n6 XThR.Tn[6].t3 24.9236
R16813 XThR.Tn[6].n6 XThR.Tn[6].t2 24.9236
R16814 XThR.Tn[6] XThR.Tn[6].n2 23.3605
R16815 XThR.Tn[6] XThR.Tn[6].n88 6.7205
R16816 XThR.Tn[6].n88 XThR.Tn[6] 5.37828
R16817 XThR.Tn[6] XThR.Tn[6].n11 5.34038
R16818 XThR.Tn[6].n16 XThR.Tn[6].n15 4.5005
R16819 XThR.Tn[6].n21 XThR.Tn[6].n20 4.5005
R16820 XThR.Tn[6].n26 XThR.Tn[6].n25 4.5005
R16821 XThR.Tn[6].n31 XThR.Tn[6].n30 4.5005
R16822 XThR.Tn[6].n36 XThR.Tn[6].n35 4.5005
R16823 XThR.Tn[6].n41 XThR.Tn[6].n40 4.5005
R16824 XThR.Tn[6].n46 XThR.Tn[6].n45 4.5005
R16825 XThR.Tn[6].n51 XThR.Tn[6].n50 4.5005
R16826 XThR.Tn[6].n56 XThR.Tn[6].n55 4.5005
R16827 XThR.Tn[6].n61 XThR.Tn[6].n60 4.5005
R16828 XThR.Tn[6].n66 XThR.Tn[6].n65 4.5005
R16829 XThR.Tn[6].n71 XThR.Tn[6].n70 4.5005
R16830 XThR.Tn[6].n76 XThR.Tn[6].n75 4.5005
R16831 XThR.Tn[6].n81 XThR.Tn[6].n80 4.5005
R16832 XThR.Tn[6].n86 XThR.Tn[6].n85 4.5005
R16833 XThR.Tn[6].n87 XThR.Tn[6] 3.70586
R16834 XThR.Tn[6].n16 XThR.Tn[6] 2.52282
R16835 XThR.Tn[6].n21 XThR.Tn[6] 2.52282
R16836 XThR.Tn[6].n26 XThR.Tn[6] 2.52282
R16837 XThR.Tn[6].n31 XThR.Tn[6] 2.52282
R16838 XThR.Tn[6].n36 XThR.Tn[6] 2.52282
R16839 XThR.Tn[6].n41 XThR.Tn[6] 2.52282
R16840 XThR.Tn[6].n46 XThR.Tn[6] 2.52282
R16841 XThR.Tn[6].n51 XThR.Tn[6] 2.52282
R16842 XThR.Tn[6].n56 XThR.Tn[6] 2.52282
R16843 XThR.Tn[6].n61 XThR.Tn[6] 2.52282
R16844 XThR.Tn[6].n66 XThR.Tn[6] 2.52282
R16845 XThR.Tn[6].n71 XThR.Tn[6] 2.52282
R16846 XThR.Tn[6].n76 XThR.Tn[6] 2.52282
R16847 XThR.Tn[6].n81 XThR.Tn[6] 2.52282
R16848 XThR.Tn[6].n86 XThR.Tn[6] 2.52282
R16849 XThR.Tn[6].n84 XThR.Tn[6] 1.08677
R16850 XThR.Tn[6].n79 XThR.Tn[6] 1.08677
R16851 XThR.Tn[6].n74 XThR.Tn[6] 1.08677
R16852 XThR.Tn[6].n69 XThR.Tn[6] 1.08677
R16853 XThR.Tn[6].n64 XThR.Tn[6] 1.08677
R16854 XThR.Tn[6].n59 XThR.Tn[6] 1.08677
R16855 XThR.Tn[6].n54 XThR.Tn[6] 1.08677
R16856 XThR.Tn[6].n49 XThR.Tn[6] 1.08677
R16857 XThR.Tn[6].n44 XThR.Tn[6] 1.08677
R16858 XThR.Tn[6].n39 XThR.Tn[6] 1.08677
R16859 XThR.Tn[6].n34 XThR.Tn[6] 1.08677
R16860 XThR.Tn[6].n29 XThR.Tn[6] 1.08677
R16861 XThR.Tn[6].n24 XThR.Tn[6] 1.08677
R16862 XThR.Tn[6].n19 XThR.Tn[6] 1.08677
R16863 XThR.Tn[6].n14 XThR.Tn[6] 1.08677
R16864 XThR.Tn[6] XThR.Tn[6].n16 0.839786
R16865 XThR.Tn[6] XThR.Tn[6].n21 0.839786
R16866 XThR.Tn[6] XThR.Tn[6].n26 0.839786
R16867 XThR.Tn[6] XThR.Tn[6].n31 0.839786
R16868 XThR.Tn[6] XThR.Tn[6].n36 0.839786
R16869 XThR.Tn[6] XThR.Tn[6].n41 0.839786
R16870 XThR.Tn[6] XThR.Tn[6].n46 0.839786
R16871 XThR.Tn[6] XThR.Tn[6].n51 0.839786
R16872 XThR.Tn[6] XThR.Tn[6].n56 0.839786
R16873 XThR.Tn[6] XThR.Tn[6].n61 0.839786
R16874 XThR.Tn[6] XThR.Tn[6].n66 0.839786
R16875 XThR.Tn[6] XThR.Tn[6].n71 0.839786
R16876 XThR.Tn[6] XThR.Tn[6].n76 0.839786
R16877 XThR.Tn[6] XThR.Tn[6].n81 0.839786
R16878 XThR.Tn[6] XThR.Tn[6].n86 0.839786
R16879 XThR.Tn[6].n11 XThR.Tn[6] 0.499542
R16880 XThR.Tn[6].n85 XThR.Tn[6] 0.063
R16881 XThR.Tn[6].n80 XThR.Tn[6] 0.063
R16882 XThR.Tn[6].n75 XThR.Tn[6] 0.063
R16883 XThR.Tn[6].n70 XThR.Tn[6] 0.063
R16884 XThR.Tn[6].n65 XThR.Tn[6] 0.063
R16885 XThR.Tn[6].n60 XThR.Tn[6] 0.063
R16886 XThR.Tn[6].n55 XThR.Tn[6] 0.063
R16887 XThR.Tn[6].n50 XThR.Tn[6] 0.063
R16888 XThR.Tn[6].n45 XThR.Tn[6] 0.063
R16889 XThR.Tn[6].n40 XThR.Tn[6] 0.063
R16890 XThR.Tn[6].n35 XThR.Tn[6] 0.063
R16891 XThR.Tn[6].n30 XThR.Tn[6] 0.063
R16892 XThR.Tn[6].n25 XThR.Tn[6] 0.063
R16893 XThR.Tn[6].n20 XThR.Tn[6] 0.063
R16894 XThR.Tn[6].n15 XThR.Tn[6] 0.063
R16895 XThR.Tn[6].n87 XThR.Tn[6] 0.0540714
R16896 XThR.Tn[6] XThR.Tn[6].n87 0.038
R16897 XThR.Tn[6].n11 XThR.Tn[6] 0.0143889
R16898 XThR.Tn[6].n85 XThR.Tn[6].n84 0.00771154
R16899 XThR.Tn[6].n80 XThR.Tn[6].n79 0.00771154
R16900 XThR.Tn[6].n75 XThR.Tn[6].n74 0.00771154
R16901 XThR.Tn[6].n70 XThR.Tn[6].n69 0.00771154
R16902 XThR.Tn[6].n65 XThR.Tn[6].n64 0.00771154
R16903 XThR.Tn[6].n60 XThR.Tn[6].n59 0.00771154
R16904 XThR.Tn[6].n55 XThR.Tn[6].n54 0.00771154
R16905 XThR.Tn[6].n50 XThR.Tn[6].n49 0.00771154
R16906 XThR.Tn[6].n45 XThR.Tn[6].n44 0.00771154
R16907 XThR.Tn[6].n40 XThR.Tn[6].n39 0.00771154
R16908 XThR.Tn[6].n35 XThR.Tn[6].n34 0.00771154
R16909 XThR.Tn[6].n30 XThR.Tn[6].n29 0.00771154
R16910 XThR.Tn[6].n25 XThR.Tn[6].n24 0.00771154
R16911 XThR.Tn[6].n20 XThR.Tn[6].n19 0.00771154
R16912 XThR.Tn[6].n15 XThR.Tn[6].n14 0.00771154
R16913 XThR.Tn[14].n87 XThR.Tn[14].n86 256.103
R16914 XThR.Tn[14].n2 XThR.Tn[14].n0 243.68
R16915 XThR.Tn[14].n5 XThR.Tn[14].n3 241.847
R16916 XThR.Tn[14].n2 XThR.Tn[14].n1 205.28
R16917 XThR.Tn[14].n87 XThR.Tn[14].n85 202.094
R16918 XThR.Tn[14].n5 XThR.Tn[14].n4 185
R16919 XThR.Tn[14] XThR.Tn[14].n78 161.363
R16920 XThR.Tn[14] XThR.Tn[14].n73 161.363
R16921 XThR.Tn[14] XThR.Tn[14].n68 161.363
R16922 XThR.Tn[14] XThR.Tn[14].n63 161.363
R16923 XThR.Tn[14] XThR.Tn[14].n58 161.363
R16924 XThR.Tn[14] XThR.Tn[14].n53 161.363
R16925 XThR.Tn[14] XThR.Tn[14].n48 161.363
R16926 XThR.Tn[14] XThR.Tn[14].n43 161.363
R16927 XThR.Tn[14] XThR.Tn[14].n38 161.363
R16928 XThR.Tn[14] XThR.Tn[14].n33 161.363
R16929 XThR.Tn[14] XThR.Tn[14].n28 161.363
R16930 XThR.Tn[14] XThR.Tn[14].n23 161.363
R16931 XThR.Tn[14] XThR.Tn[14].n18 161.363
R16932 XThR.Tn[14] XThR.Tn[14].n13 161.363
R16933 XThR.Tn[14] XThR.Tn[14].n8 161.363
R16934 XThR.Tn[14] XThR.Tn[14].n6 161.363
R16935 XThR.Tn[14].n80 XThR.Tn[14].n79 161.3
R16936 XThR.Tn[14].n75 XThR.Tn[14].n74 161.3
R16937 XThR.Tn[14].n70 XThR.Tn[14].n69 161.3
R16938 XThR.Tn[14].n65 XThR.Tn[14].n64 161.3
R16939 XThR.Tn[14].n60 XThR.Tn[14].n59 161.3
R16940 XThR.Tn[14].n55 XThR.Tn[14].n54 161.3
R16941 XThR.Tn[14].n50 XThR.Tn[14].n49 161.3
R16942 XThR.Tn[14].n45 XThR.Tn[14].n44 161.3
R16943 XThR.Tn[14].n40 XThR.Tn[14].n39 161.3
R16944 XThR.Tn[14].n35 XThR.Tn[14].n34 161.3
R16945 XThR.Tn[14].n30 XThR.Tn[14].n29 161.3
R16946 XThR.Tn[14].n25 XThR.Tn[14].n24 161.3
R16947 XThR.Tn[14].n20 XThR.Tn[14].n19 161.3
R16948 XThR.Tn[14].n15 XThR.Tn[14].n14 161.3
R16949 XThR.Tn[14].n10 XThR.Tn[14].n9 161.3
R16950 XThR.Tn[14].n78 XThR.Tn[14].t51 161.106
R16951 XThR.Tn[14].n73 XThR.Tn[14].t58 161.106
R16952 XThR.Tn[14].n68 XThR.Tn[14].t39 161.106
R16953 XThR.Tn[14].n63 XThR.Tn[14].t22 161.106
R16954 XThR.Tn[14].n58 XThR.Tn[14].t49 161.106
R16955 XThR.Tn[14].n53 XThR.Tn[14].t12 161.106
R16956 XThR.Tn[14].n48 XThR.Tn[14].t56 161.106
R16957 XThR.Tn[14].n43 XThR.Tn[14].t36 161.106
R16958 XThR.Tn[14].n38 XThR.Tn[14].t19 161.106
R16959 XThR.Tn[14].n33 XThR.Tn[14].t25 161.106
R16960 XThR.Tn[14].n28 XThR.Tn[14].t73 161.106
R16961 XThR.Tn[14].n23 XThR.Tn[14].t38 161.106
R16962 XThR.Tn[14].n18 XThR.Tn[14].t72 161.106
R16963 XThR.Tn[14].n13 XThR.Tn[14].t54 161.106
R16964 XThR.Tn[14].n8 XThR.Tn[14].t13 161.106
R16965 XThR.Tn[14].n6 XThR.Tn[14].t62 161.106
R16966 XThR.Tn[14].n79 XThR.Tn[14].t32 159.978
R16967 XThR.Tn[14].n74 XThR.Tn[14].t37 159.978
R16968 XThR.Tn[14].n69 XThR.Tn[14].t20 159.978
R16969 XThR.Tn[14].n64 XThR.Tn[14].t68 159.978
R16970 XThR.Tn[14].n59 XThR.Tn[14].t30 159.978
R16971 XThR.Tn[14].n54 XThR.Tn[14].t55 159.978
R16972 XThR.Tn[14].n49 XThR.Tn[14].t35 159.978
R16973 XThR.Tn[14].n44 XThR.Tn[14].t16 159.978
R16974 XThR.Tn[14].n39 XThR.Tn[14].t66 159.978
R16975 XThR.Tn[14].n34 XThR.Tn[14].t71 159.978
R16976 XThR.Tn[14].n29 XThR.Tn[14].t53 159.978
R16977 XThR.Tn[14].n24 XThR.Tn[14].t18 159.978
R16978 XThR.Tn[14].n19 XThR.Tn[14].t52 159.978
R16979 XThR.Tn[14].n14 XThR.Tn[14].t34 159.978
R16980 XThR.Tn[14].n9 XThR.Tn[14].t60 159.978
R16981 XThR.Tn[14].n78 XThR.Tn[14].t41 145.038
R16982 XThR.Tn[14].n73 XThR.Tn[14].t65 145.038
R16983 XThR.Tn[14].n68 XThR.Tn[14].t45 145.038
R16984 XThR.Tn[14].n63 XThR.Tn[14].t26 145.038
R16985 XThR.Tn[14].n58 XThR.Tn[14].t59 145.038
R16986 XThR.Tn[14].n53 XThR.Tn[14].t40 145.038
R16987 XThR.Tn[14].n48 XThR.Tn[14].t46 145.038
R16988 XThR.Tn[14].n43 XThR.Tn[14].t27 145.038
R16989 XThR.Tn[14].n38 XThR.Tn[14].t23 145.038
R16990 XThR.Tn[14].n33 XThR.Tn[14].t57 145.038
R16991 XThR.Tn[14].n28 XThR.Tn[14].t15 145.038
R16992 XThR.Tn[14].n23 XThR.Tn[14].t44 145.038
R16993 XThR.Tn[14].n18 XThR.Tn[14].t14 145.038
R16994 XThR.Tn[14].n13 XThR.Tn[14].t64 145.038
R16995 XThR.Tn[14].n8 XThR.Tn[14].t24 145.038
R16996 XThR.Tn[14].n6 XThR.Tn[14].t69 145.038
R16997 XThR.Tn[14].n79 XThR.Tn[14].t43 143.911
R16998 XThR.Tn[14].n74 XThR.Tn[14].t70 143.911
R16999 XThR.Tn[14].n69 XThR.Tn[14].t48 143.911
R17000 XThR.Tn[14].n64 XThR.Tn[14].t31 143.911
R17001 XThR.Tn[14].n59 XThR.Tn[14].t63 143.911
R17002 XThR.Tn[14].n54 XThR.Tn[14].t42 143.911
R17003 XThR.Tn[14].n49 XThR.Tn[14].t50 143.911
R17004 XThR.Tn[14].n44 XThR.Tn[14].t33 143.911
R17005 XThR.Tn[14].n39 XThR.Tn[14].t29 143.911
R17006 XThR.Tn[14].n34 XThR.Tn[14].t61 143.911
R17007 XThR.Tn[14].n29 XThR.Tn[14].t21 143.911
R17008 XThR.Tn[14].n24 XThR.Tn[14].t47 143.911
R17009 XThR.Tn[14].n19 XThR.Tn[14].t17 143.911
R17010 XThR.Tn[14].n14 XThR.Tn[14].t67 143.911
R17011 XThR.Tn[14].n9 XThR.Tn[14].t28 143.911
R17012 XThR.Tn[14] XThR.Tn[14].n2 35.7652
R17013 XThR.Tn[14].n86 XThR.Tn[14].t0 26.5955
R17014 XThR.Tn[14].n86 XThR.Tn[14].t1 26.5955
R17015 XThR.Tn[14].n0 XThR.Tn[14].t8 26.5955
R17016 XThR.Tn[14].n0 XThR.Tn[14].t9 26.5955
R17017 XThR.Tn[14].n1 XThR.Tn[14].t10 26.5955
R17018 XThR.Tn[14].n1 XThR.Tn[14].t11 26.5955
R17019 XThR.Tn[14].n85 XThR.Tn[14].t2 26.5955
R17020 XThR.Tn[14].n85 XThR.Tn[14].t3 26.5955
R17021 XThR.Tn[14].n4 XThR.Tn[14].t4 24.9236
R17022 XThR.Tn[14].n4 XThR.Tn[14].t5 24.9236
R17023 XThR.Tn[14].n3 XThR.Tn[14].t6 24.9236
R17024 XThR.Tn[14].n3 XThR.Tn[14].t7 24.9236
R17025 XThR.Tn[14] XThR.Tn[14].n5 18.8943
R17026 XThR.Tn[14].n88 XThR.Tn[14].n87 13.5534
R17027 XThR.Tn[14].n84 XThR.Tn[14] 8.47191
R17028 XThR.Tn[14].n84 XThR.Tn[14] 6.34069
R17029 XThR.Tn[14] XThR.Tn[14].n7 5.34038
R17030 XThR.Tn[14].n12 XThR.Tn[14].n11 4.5005
R17031 XThR.Tn[14].n17 XThR.Tn[14].n16 4.5005
R17032 XThR.Tn[14].n22 XThR.Tn[14].n21 4.5005
R17033 XThR.Tn[14].n27 XThR.Tn[14].n26 4.5005
R17034 XThR.Tn[14].n32 XThR.Tn[14].n31 4.5005
R17035 XThR.Tn[14].n37 XThR.Tn[14].n36 4.5005
R17036 XThR.Tn[14].n42 XThR.Tn[14].n41 4.5005
R17037 XThR.Tn[14].n47 XThR.Tn[14].n46 4.5005
R17038 XThR.Tn[14].n52 XThR.Tn[14].n51 4.5005
R17039 XThR.Tn[14].n57 XThR.Tn[14].n56 4.5005
R17040 XThR.Tn[14].n62 XThR.Tn[14].n61 4.5005
R17041 XThR.Tn[14].n67 XThR.Tn[14].n66 4.5005
R17042 XThR.Tn[14].n72 XThR.Tn[14].n71 4.5005
R17043 XThR.Tn[14].n77 XThR.Tn[14].n76 4.5005
R17044 XThR.Tn[14].n82 XThR.Tn[14].n81 4.5005
R17045 XThR.Tn[14].n83 XThR.Tn[14] 3.70586
R17046 XThR.Tn[14].n12 XThR.Tn[14] 2.52282
R17047 XThR.Tn[14].n17 XThR.Tn[14] 2.52282
R17048 XThR.Tn[14].n22 XThR.Tn[14] 2.52282
R17049 XThR.Tn[14].n27 XThR.Tn[14] 2.52282
R17050 XThR.Tn[14].n32 XThR.Tn[14] 2.52282
R17051 XThR.Tn[14].n37 XThR.Tn[14] 2.52282
R17052 XThR.Tn[14].n42 XThR.Tn[14] 2.52282
R17053 XThR.Tn[14].n47 XThR.Tn[14] 2.52282
R17054 XThR.Tn[14].n52 XThR.Tn[14] 2.52282
R17055 XThR.Tn[14].n57 XThR.Tn[14] 2.52282
R17056 XThR.Tn[14].n62 XThR.Tn[14] 2.52282
R17057 XThR.Tn[14].n67 XThR.Tn[14] 2.52282
R17058 XThR.Tn[14].n72 XThR.Tn[14] 2.52282
R17059 XThR.Tn[14].n77 XThR.Tn[14] 2.52282
R17060 XThR.Tn[14].n82 XThR.Tn[14] 2.52282
R17061 XThR.Tn[14] XThR.Tn[14].n84 1.79489
R17062 XThR.Tn[14] XThR.Tn[14].n88 1.50638
R17063 XThR.Tn[14].n88 XThR.Tn[14] 1.19676
R17064 XThR.Tn[14].n80 XThR.Tn[14] 1.08677
R17065 XThR.Tn[14].n75 XThR.Tn[14] 1.08677
R17066 XThR.Tn[14].n70 XThR.Tn[14] 1.08677
R17067 XThR.Tn[14].n65 XThR.Tn[14] 1.08677
R17068 XThR.Tn[14].n60 XThR.Tn[14] 1.08677
R17069 XThR.Tn[14].n55 XThR.Tn[14] 1.08677
R17070 XThR.Tn[14].n50 XThR.Tn[14] 1.08677
R17071 XThR.Tn[14].n45 XThR.Tn[14] 1.08677
R17072 XThR.Tn[14].n40 XThR.Tn[14] 1.08677
R17073 XThR.Tn[14].n35 XThR.Tn[14] 1.08677
R17074 XThR.Tn[14].n30 XThR.Tn[14] 1.08677
R17075 XThR.Tn[14].n25 XThR.Tn[14] 1.08677
R17076 XThR.Tn[14].n20 XThR.Tn[14] 1.08677
R17077 XThR.Tn[14].n15 XThR.Tn[14] 1.08677
R17078 XThR.Tn[14].n10 XThR.Tn[14] 1.08677
R17079 XThR.Tn[14] XThR.Tn[14].n12 0.839786
R17080 XThR.Tn[14] XThR.Tn[14].n17 0.839786
R17081 XThR.Tn[14] XThR.Tn[14].n22 0.839786
R17082 XThR.Tn[14] XThR.Tn[14].n27 0.839786
R17083 XThR.Tn[14] XThR.Tn[14].n32 0.839786
R17084 XThR.Tn[14] XThR.Tn[14].n37 0.839786
R17085 XThR.Tn[14] XThR.Tn[14].n42 0.839786
R17086 XThR.Tn[14] XThR.Tn[14].n47 0.839786
R17087 XThR.Tn[14] XThR.Tn[14].n52 0.839786
R17088 XThR.Tn[14] XThR.Tn[14].n57 0.839786
R17089 XThR.Tn[14] XThR.Tn[14].n62 0.839786
R17090 XThR.Tn[14] XThR.Tn[14].n67 0.839786
R17091 XThR.Tn[14] XThR.Tn[14].n72 0.839786
R17092 XThR.Tn[14] XThR.Tn[14].n77 0.839786
R17093 XThR.Tn[14] XThR.Tn[14].n82 0.839786
R17094 XThR.Tn[14].n7 XThR.Tn[14] 0.499542
R17095 XThR.Tn[14].n81 XThR.Tn[14] 0.063
R17096 XThR.Tn[14].n76 XThR.Tn[14] 0.063
R17097 XThR.Tn[14].n71 XThR.Tn[14] 0.063
R17098 XThR.Tn[14].n66 XThR.Tn[14] 0.063
R17099 XThR.Tn[14].n61 XThR.Tn[14] 0.063
R17100 XThR.Tn[14].n56 XThR.Tn[14] 0.063
R17101 XThR.Tn[14].n51 XThR.Tn[14] 0.063
R17102 XThR.Tn[14].n46 XThR.Tn[14] 0.063
R17103 XThR.Tn[14].n41 XThR.Tn[14] 0.063
R17104 XThR.Tn[14].n36 XThR.Tn[14] 0.063
R17105 XThR.Tn[14].n31 XThR.Tn[14] 0.063
R17106 XThR.Tn[14].n26 XThR.Tn[14] 0.063
R17107 XThR.Tn[14].n21 XThR.Tn[14] 0.063
R17108 XThR.Tn[14].n16 XThR.Tn[14] 0.063
R17109 XThR.Tn[14].n11 XThR.Tn[14] 0.063
R17110 XThR.Tn[14].n83 XThR.Tn[14] 0.0540714
R17111 XThR.Tn[14] XThR.Tn[14].n83 0.038
R17112 XThR.Tn[14].n7 XThR.Tn[14] 0.0143889
R17113 XThR.Tn[14].n81 XThR.Tn[14].n80 0.00771154
R17114 XThR.Tn[14].n76 XThR.Tn[14].n75 0.00771154
R17115 XThR.Tn[14].n71 XThR.Tn[14].n70 0.00771154
R17116 XThR.Tn[14].n66 XThR.Tn[14].n65 0.00771154
R17117 XThR.Tn[14].n61 XThR.Tn[14].n60 0.00771154
R17118 XThR.Tn[14].n56 XThR.Tn[14].n55 0.00771154
R17119 XThR.Tn[14].n51 XThR.Tn[14].n50 0.00771154
R17120 XThR.Tn[14].n46 XThR.Tn[14].n45 0.00771154
R17121 XThR.Tn[14].n41 XThR.Tn[14].n40 0.00771154
R17122 XThR.Tn[14].n36 XThR.Tn[14].n35 0.00771154
R17123 XThR.Tn[14].n31 XThR.Tn[14].n30 0.00771154
R17124 XThR.Tn[14].n26 XThR.Tn[14].n25 0.00771154
R17125 XThR.Tn[14].n21 XThR.Tn[14].n20 0.00771154
R17126 XThR.Tn[14].n16 XThR.Tn[14].n15 0.00771154
R17127 XThR.Tn[14].n11 XThR.Tn[14].n10 0.00771154
R17128 XThR.Tn[12].n5 XThR.Tn[12].n4 256.103
R17129 XThR.Tn[12].n2 XThR.Tn[12].n0 243.68
R17130 XThR.Tn[12].n88 XThR.Tn[12].n87 241.847
R17131 XThR.Tn[12].n2 XThR.Tn[12].n1 205.28
R17132 XThR.Tn[12].n5 XThR.Tn[12].n3 202.095
R17133 XThR.Tn[12].n88 XThR.Tn[12].n86 185
R17134 XThR.Tn[12] XThR.Tn[12].n79 161.363
R17135 XThR.Tn[12] XThR.Tn[12].n74 161.363
R17136 XThR.Tn[12] XThR.Tn[12].n69 161.363
R17137 XThR.Tn[12] XThR.Tn[12].n64 161.363
R17138 XThR.Tn[12] XThR.Tn[12].n59 161.363
R17139 XThR.Tn[12] XThR.Tn[12].n54 161.363
R17140 XThR.Tn[12] XThR.Tn[12].n49 161.363
R17141 XThR.Tn[12] XThR.Tn[12].n44 161.363
R17142 XThR.Tn[12] XThR.Tn[12].n39 161.363
R17143 XThR.Tn[12] XThR.Tn[12].n34 161.363
R17144 XThR.Tn[12] XThR.Tn[12].n29 161.363
R17145 XThR.Tn[12] XThR.Tn[12].n24 161.363
R17146 XThR.Tn[12] XThR.Tn[12].n19 161.363
R17147 XThR.Tn[12] XThR.Tn[12].n14 161.363
R17148 XThR.Tn[12] XThR.Tn[12].n9 161.363
R17149 XThR.Tn[12] XThR.Tn[12].n7 161.363
R17150 XThR.Tn[12].n81 XThR.Tn[12].n80 161.3
R17151 XThR.Tn[12].n76 XThR.Tn[12].n75 161.3
R17152 XThR.Tn[12].n71 XThR.Tn[12].n70 161.3
R17153 XThR.Tn[12].n66 XThR.Tn[12].n65 161.3
R17154 XThR.Tn[12].n61 XThR.Tn[12].n60 161.3
R17155 XThR.Tn[12].n56 XThR.Tn[12].n55 161.3
R17156 XThR.Tn[12].n51 XThR.Tn[12].n50 161.3
R17157 XThR.Tn[12].n46 XThR.Tn[12].n45 161.3
R17158 XThR.Tn[12].n41 XThR.Tn[12].n40 161.3
R17159 XThR.Tn[12].n36 XThR.Tn[12].n35 161.3
R17160 XThR.Tn[12].n31 XThR.Tn[12].n30 161.3
R17161 XThR.Tn[12].n26 XThR.Tn[12].n25 161.3
R17162 XThR.Tn[12].n21 XThR.Tn[12].n20 161.3
R17163 XThR.Tn[12].n16 XThR.Tn[12].n15 161.3
R17164 XThR.Tn[12].n11 XThR.Tn[12].n10 161.3
R17165 XThR.Tn[12].n79 XThR.Tn[12].t18 161.106
R17166 XThR.Tn[12].n74 XThR.Tn[12].t24 161.106
R17167 XThR.Tn[12].n69 XThR.Tn[12].t67 161.106
R17168 XThR.Tn[12].n64 XThR.Tn[12].t52 161.106
R17169 XThR.Tn[12].n59 XThR.Tn[12].t16 161.106
R17170 XThR.Tn[12].n54 XThR.Tn[12].t40 161.106
R17171 XThR.Tn[12].n49 XThR.Tn[12].t22 161.106
R17172 XThR.Tn[12].n44 XThR.Tn[12].t65 161.106
R17173 XThR.Tn[12].n39 XThR.Tn[12].t51 161.106
R17174 XThR.Tn[12].n34 XThR.Tn[12].t56 161.106
R17175 XThR.Tn[12].n29 XThR.Tn[12].t39 161.106
R17176 XThR.Tn[12].n24 XThR.Tn[12].t66 161.106
R17177 XThR.Tn[12].n19 XThR.Tn[12].t38 161.106
R17178 XThR.Tn[12].n14 XThR.Tn[12].t20 161.106
R17179 XThR.Tn[12].n9 XThR.Tn[12].t43 161.106
R17180 XThR.Tn[12].n7 XThR.Tn[12].t28 161.106
R17181 XThR.Tn[12].n80 XThR.Tn[12].t58 159.978
R17182 XThR.Tn[12].n75 XThR.Tn[12].t62 159.978
R17183 XThR.Tn[12].n70 XThR.Tn[12].t47 159.978
R17184 XThR.Tn[12].n65 XThR.Tn[12].t31 159.978
R17185 XThR.Tn[12].n60 XThR.Tn[12].t55 159.978
R17186 XThR.Tn[12].n55 XThR.Tn[12].t19 159.978
R17187 XThR.Tn[12].n50 XThR.Tn[12].t61 159.978
R17188 XThR.Tn[12].n45 XThR.Tn[12].t44 159.978
R17189 XThR.Tn[12].n40 XThR.Tn[12].t29 159.978
R17190 XThR.Tn[12].n35 XThR.Tn[12].t37 159.978
R17191 XThR.Tn[12].n30 XThR.Tn[12].t17 159.978
R17192 XThR.Tn[12].n25 XThR.Tn[12].t46 159.978
R17193 XThR.Tn[12].n20 XThR.Tn[12].t15 159.978
R17194 XThR.Tn[12].n15 XThR.Tn[12].t60 159.978
R17195 XThR.Tn[12].n10 XThR.Tn[12].t21 159.978
R17196 XThR.Tn[12].n79 XThR.Tn[12].t69 145.038
R17197 XThR.Tn[12].n74 XThR.Tn[12].t32 145.038
R17198 XThR.Tn[12].n69 XThR.Tn[12].t73 145.038
R17199 XThR.Tn[12].n64 XThR.Tn[12].t57 145.038
R17200 XThR.Tn[12].n59 XThR.Tn[12].t25 145.038
R17201 XThR.Tn[12].n54 XThR.Tn[12].t68 145.038
R17202 XThR.Tn[12].n49 XThR.Tn[12].t12 145.038
R17203 XThR.Tn[12].n44 XThR.Tn[12].t59 145.038
R17204 XThR.Tn[12].n39 XThR.Tn[12].t54 145.038
R17205 XThR.Tn[12].n34 XThR.Tn[12].t23 145.038
R17206 XThR.Tn[12].n29 XThR.Tn[12].t48 145.038
R17207 XThR.Tn[12].n24 XThR.Tn[12].t70 145.038
R17208 XThR.Tn[12].n19 XThR.Tn[12].t45 145.038
R17209 XThR.Tn[12].n14 XThR.Tn[12].t30 145.038
R17210 XThR.Tn[12].n9 XThR.Tn[12].t53 145.038
R17211 XThR.Tn[12].n7 XThR.Tn[12].t36 145.038
R17212 XThR.Tn[12].n80 XThR.Tn[12].t27 143.911
R17213 XThR.Tn[12].n75 XThR.Tn[12].t50 143.911
R17214 XThR.Tn[12].n70 XThR.Tn[12].t34 143.911
R17215 XThR.Tn[12].n65 XThR.Tn[12].t13 143.911
R17216 XThR.Tn[12].n60 XThR.Tn[12].t42 143.911
R17217 XThR.Tn[12].n55 XThR.Tn[12].t26 143.911
R17218 XThR.Tn[12].n50 XThR.Tn[12].t35 143.911
R17219 XThR.Tn[12].n45 XThR.Tn[12].t14 143.911
R17220 XThR.Tn[12].n40 XThR.Tn[12].t72 143.911
R17221 XThR.Tn[12].n35 XThR.Tn[12].t41 143.911
R17222 XThR.Tn[12].n30 XThR.Tn[12].t64 143.911
R17223 XThR.Tn[12].n25 XThR.Tn[12].t33 143.911
R17224 XThR.Tn[12].n20 XThR.Tn[12].t63 143.911
R17225 XThR.Tn[12].n15 XThR.Tn[12].t49 143.911
R17226 XThR.Tn[12].n10 XThR.Tn[12].t71 143.911
R17227 XThR.Tn[12] XThR.Tn[12].n2 35.7652
R17228 XThR.Tn[12].n3 XThR.Tn[12].t6 26.5955
R17229 XThR.Tn[12].n3 XThR.Tn[12].t4 26.5955
R17230 XThR.Tn[12].n4 XThR.Tn[12].t7 26.5955
R17231 XThR.Tn[12].n4 XThR.Tn[12].t5 26.5955
R17232 XThR.Tn[12].n0 XThR.Tn[12].t11 26.5955
R17233 XThR.Tn[12].n0 XThR.Tn[12].t9 26.5955
R17234 XThR.Tn[12].n1 XThR.Tn[12].t8 26.5955
R17235 XThR.Tn[12].n1 XThR.Tn[12].t10 26.5955
R17236 XThR.Tn[12].n86 XThR.Tn[12].t2 24.9236
R17237 XThR.Tn[12].n86 XThR.Tn[12].t0 24.9236
R17238 XThR.Tn[12].n87 XThR.Tn[12].t3 24.9236
R17239 XThR.Tn[12].n87 XThR.Tn[12].t1 24.9236
R17240 XThR.Tn[12] XThR.Tn[12].n88 18.8943
R17241 XThR.Tn[12].n6 XThR.Tn[12].n5 13.5534
R17242 XThR.Tn[12].n85 XThR.Tn[12] 8.18715
R17243 XThR.Tn[12] XThR.Tn[12].n85 6.34069
R17244 XThR.Tn[12] XThR.Tn[12].n8 5.34038
R17245 XThR.Tn[12].n13 XThR.Tn[12].n12 4.5005
R17246 XThR.Tn[12].n18 XThR.Tn[12].n17 4.5005
R17247 XThR.Tn[12].n23 XThR.Tn[12].n22 4.5005
R17248 XThR.Tn[12].n28 XThR.Tn[12].n27 4.5005
R17249 XThR.Tn[12].n33 XThR.Tn[12].n32 4.5005
R17250 XThR.Tn[12].n38 XThR.Tn[12].n37 4.5005
R17251 XThR.Tn[12].n43 XThR.Tn[12].n42 4.5005
R17252 XThR.Tn[12].n48 XThR.Tn[12].n47 4.5005
R17253 XThR.Tn[12].n53 XThR.Tn[12].n52 4.5005
R17254 XThR.Tn[12].n58 XThR.Tn[12].n57 4.5005
R17255 XThR.Tn[12].n63 XThR.Tn[12].n62 4.5005
R17256 XThR.Tn[12].n68 XThR.Tn[12].n67 4.5005
R17257 XThR.Tn[12].n73 XThR.Tn[12].n72 4.5005
R17258 XThR.Tn[12].n78 XThR.Tn[12].n77 4.5005
R17259 XThR.Tn[12].n83 XThR.Tn[12].n82 4.5005
R17260 XThR.Tn[12].n84 XThR.Tn[12] 3.70586
R17261 XThR.Tn[12].n13 XThR.Tn[12] 2.52282
R17262 XThR.Tn[12].n18 XThR.Tn[12] 2.52282
R17263 XThR.Tn[12].n23 XThR.Tn[12] 2.52282
R17264 XThR.Tn[12].n28 XThR.Tn[12] 2.52282
R17265 XThR.Tn[12].n33 XThR.Tn[12] 2.52282
R17266 XThR.Tn[12].n38 XThR.Tn[12] 2.52282
R17267 XThR.Tn[12].n43 XThR.Tn[12] 2.52282
R17268 XThR.Tn[12].n48 XThR.Tn[12] 2.52282
R17269 XThR.Tn[12].n53 XThR.Tn[12] 2.52282
R17270 XThR.Tn[12].n58 XThR.Tn[12] 2.52282
R17271 XThR.Tn[12].n63 XThR.Tn[12] 2.52282
R17272 XThR.Tn[12].n68 XThR.Tn[12] 2.52282
R17273 XThR.Tn[12].n73 XThR.Tn[12] 2.52282
R17274 XThR.Tn[12].n78 XThR.Tn[12] 2.52282
R17275 XThR.Tn[12].n83 XThR.Tn[12] 2.52282
R17276 XThR.Tn[12].n85 XThR.Tn[12] 1.79489
R17277 XThR.Tn[12].n6 XThR.Tn[12] 1.50638
R17278 XThR.Tn[12] XThR.Tn[12].n6 1.19676
R17279 XThR.Tn[12].n81 XThR.Tn[12] 1.08677
R17280 XThR.Tn[12].n76 XThR.Tn[12] 1.08677
R17281 XThR.Tn[12].n71 XThR.Tn[12] 1.08677
R17282 XThR.Tn[12].n66 XThR.Tn[12] 1.08677
R17283 XThR.Tn[12].n61 XThR.Tn[12] 1.08677
R17284 XThR.Tn[12].n56 XThR.Tn[12] 1.08677
R17285 XThR.Tn[12].n51 XThR.Tn[12] 1.08677
R17286 XThR.Tn[12].n46 XThR.Tn[12] 1.08677
R17287 XThR.Tn[12].n41 XThR.Tn[12] 1.08677
R17288 XThR.Tn[12].n36 XThR.Tn[12] 1.08677
R17289 XThR.Tn[12].n31 XThR.Tn[12] 1.08677
R17290 XThR.Tn[12].n26 XThR.Tn[12] 1.08677
R17291 XThR.Tn[12].n21 XThR.Tn[12] 1.08677
R17292 XThR.Tn[12].n16 XThR.Tn[12] 1.08677
R17293 XThR.Tn[12].n11 XThR.Tn[12] 1.08677
R17294 XThR.Tn[12] XThR.Tn[12].n13 0.839786
R17295 XThR.Tn[12] XThR.Tn[12].n18 0.839786
R17296 XThR.Tn[12] XThR.Tn[12].n23 0.839786
R17297 XThR.Tn[12] XThR.Tn[12].n28 0.839786
R17298 XThR.Tn[12] XThR.Tn[12].n33 0.839786
R17299 XThR.Tn[12] XThR.Tn[12].n38 0.839786
R17300 XThR.Tn[12] XThR.Tn[12].n43 0.839786
R17301 XThR.Tn[12] XThR.Tn[12].n48 0.839786
R17302 XThR.Tn[12] XThR.Tn[12].n53 0.839786
R17303 XThR.Tn[12] XThR.Tn[12].n58 0.839786
R17304 XThR.Tn[12] XThR.Tn[12].n63 0.839786
R17305 XThR.Tn[12] XThR.Tn[12].n68 0.839786
R17306 XThR.Tn[12] XThR.Tn[12].n73 0.839786
R17307 XThR.Tn[12] XThR.Tn[12].n78 0.839786
R17308 XThR.Tn[12] XThR.Tn[12].n83 0.839786
R17309 XThR.Tn[12].n8 XThR.Tn[12] 0.499542
R17310 XThR.Tn[12].n82 XThR.Tn[12] 0.063
R17311 XThR.Tn[12].n77 XThR.Tn[12] 0.063
R17312 XThR.Tn[12].n72 XThR.Tn[12] 0.063
R17313 XThR.Tn[12].n67 XThR.Tn[12] 0.063
R17314 XThR.Tn[12].n62 XThR.Tn[12] 0.063
R17315 XThR.Tn[12].n57 XThR.Tn[12] 0.063
R17316 XThR.Tn[12].n52 XThR.Tn[12] 0.063
R17317 XThR.Tn[12].n47 XThR.Tn[12] 0.063
R17318 XThR.Tn[12].n42 XThR.Tn[12] 0.063
R17319 XThR.Tn[12].n37 XThR.Tn[12] 0.063
R17320 XThR.Tn[12].n32 XThR.Tn[12] 0.063
R17321 XThR.Tn[12].n27 XThR.Tn[12] 0.063
R17322 XThR.Tn[12].n22 XThR.Tn[12] 0.063
R17323 XThR.Tn[12].n17 XThR.Tn[12] 0.063
R17324 XThR.Tn[12].n12 XThR.Tn[12] 0.063
R17325 XThR.Tn[12].n84 XThR.Tn[12] 0.0540714
R17326 XThR.Tn[12] XThR.Tn[12].n84 0.038
R17327 XThR.Tn[12].n8 XThR.Tn[12] 0.0143889
R17328 XThR.Tn[12].n82 XThR.Tn[12].n81 0.00771154
R17329 XThR.Tn[12].n77 XThR.Tn[12].n76 0.00771154
R17330 XThR.Tn[12].n72 XThR.Tn[12].n71 0.00771154
R17331 XThR.Tn[12].n67 XThR.Tn[12].n66 0.00771154
R17332 XThR.Tn[12].n62 XThR.Tn[12].n61 0.00771154
R17333 XThR.Tn[12].n57 XThR.Tn[12].n56 0.00771154
R17334 XThR.Tn[12].n52 XThR.Tn[12].n51 0.00771154
R17335 XThR.Tn[12].n47 XThR.Tn[12].n46 0.00771154
R17336 XThR.Tn[12].n42 XThR.Tn[12].n41 0.00771154
R17337 XThR.Tn[12].n37 XThR.Tn[12].n36 0.00771154
R17338 XThR.Tn[12].n32 XThR.Tn[12].n31 0.00771154
R17339 XThR.Tn[12].n27 XThR.Tn[12].n26 0.00771154
R17340 XThR.Tn[12].n22 XThR.Tn[12].n21 0.00771154
R17341 XThR.Tn[12].n17 XThR.Tn[12].n16 0.00771154
R17342 XThR.Tn[12].n12 XThR.Tn[12].n11 0.00771154
R17343 thermo15c_0.XTBN.Y.n182 thermo15c_0.XTBN.Y.t9 212.081
R17344 thermo15c_0.XTBN.Y.n181 thermo15c_0.XTBN.Y.t75 212.081
R17345 thermo15c_0.XTBN.Y.n175 thermo15c_0.XTBN.Y.t33 212.081
R17346 thermo15c_0.XTBN.Y.n176 thermo15c_0.XTBN.Y.t27 212.081
R17347 thermo15c_0.XTBN.Y.n87 thermo15c_0.XTBN.Y.t25 212.081
R17348 thermo15c_0.XTBN.Y.n78 thermo15c_0.XTBN.Y.t100 212.081
R17349 thermo15c_0.XTBN.Y.n82 thermo15c_0.XTBN.Y.t93 212.081
R17350 thermo15c_0.XTBN.Y.n80 thermo15c_0.XTBN.Y.t90 212.081
R17351 thermo15c_0.XTBN.Y.n61 thermo15c_0.XTBN.Y.t47 212.081
R17352 thermo15c_0.XTBN.Y.n52 thermo15c_0.XTBN.Y.t17 212.081
R17353 thermo15c_0.XTBN.Y.n56 thermo15c_0.XTBN.Y.t116 212.081
R17354 thermo15c_0.XTBN.Y.n54 thermo15c_0.XTBN.Y.t111 212.081
R17355 thermo15c_0.XTBN.Y.n35 thermo15c_0.XTBN.Y.t106 212.081
R17356 thermo15c_0.XTBN.Y.n26 thermo15c_0.XTBN.Y.t70 212.081
R17357 thermo15c_0.XTBN.Y.n30 thermo15c_0.XTBN.Y.t56 212.081
R17358 thermo15c_0.XTBN.Y.n28 thermo15c_0.XTBN.Y.t48 212.081
R17359 thermo15c_0.XTBN.Y.n10 thermo15c_0.XTBN.Y.t50 212.081
R17360 thermo15c_0.XTBN.Y.n1 thermo15c_0.XTBN.Y.t18 212.081
R17361 thermo15c_0.XTBN.Y.n5 thermo15c_0.XTBN.Y.t120 212.081
R17362 thermo15c_0.XTBN.Y.n3 thermo15c_0.XTBN.Y.t114 212.081
R17363 thermo15c_0.XTBN.Y.n74 thermo15c_0.XTBN.Y.t101 212.081
R17364 thermo15c_0.XTBN.Y.n65 thermo15c_0.XTBN.Y.t63 212.081
R17365 thermo15c_0.XTBN.Y.n69 thermo15c_0.XTBN.Y.t52 212.081
R17366 thermo15c_0.XTBN.Y.n67 thermo15c_0.XTBN.Y.t44 212.081
R17367 thermo15c_0.XTBN.Y.n48 thermo15c_0.XTBN.Y.t39 212.081
R17368 thermo15c_0.XTBN.Y.n39 thermo15c_0.XTBN.Y.t122 212.081
R17369 thermo15c_0.XTBN.Y.n43 thermo15c_0.XTBN.Y.t109 212.081
R17370 thermo15c_0.XTBN.Y.n41 thermo15c_0.XTBN.Y.t102 212.081
R17371 thermo15c_0.XTBN.Y.n22 thermo15c_0.XTBN.Y.t79 212.081
R17372 thermo15c_0.XTBN.Y.n13 thermo15c_0.XTBN.Y.t36 212.081
R17373 thermo15c_0.XTBN.Y.n17 thermo15c_0.XTBN.Y.t26 212.081
R17374 thermo15c_0.XTBN.Y.n15 thermo15c_0.XTBN.Y.t21 212.081
R17375 thermo15c_0.XTBN.Y.n99 thermo15c_0.XTBN.Y.t54 212.081
R17376 thermo15c_0.XTBN.Y.n98 thermo15c_0.XTBN.Y.t46 212.081
R17377 thermo15c_0.XTBN.Y.n93 thermo15c_0.XTBN.Y.t12 212.081
R17378 thermo15c_0.XTBN.Y.n92 thermo15c_0.XTBN.Y.t6 212.081
R17379 thermo15c_0.XTBN.Y.n122 thermo15c_0.XTBN.Y.t34 212.081
R17380 thermo15c_0.XTBN.Y.n121 thermo15c_0.XTBN.Y.t30 212.081
R17381 thermo15c_0.XTBN.Y.n116 thermo15c_0.XTBN.Y.t103 212.081
R17382 thermo15c_0.XTBN.Y.n115 thermo15c_0.XTBN.Y.t98 212.081
R17383 thermo15c_0.XTBN.Y.n146 thermo15c_0.XTBN.Y.t91 212.081
R17384 thermo15c_0.XTBN.Y.n145 thermo15c_0.XTBN.Y.t88 212.081
R17385 thermo15c_0.XTBN.Y.n140 thermo15c_0.XTBN.Y.t40 212.081
R17386 thermo15c_0.XTBN.Y.n139 thermo15c_0.XTBN.Y.t37 212.081
R17387 thermo15c_0.XTBN.Y.n170 thermo15c_0.XTBN.Y.t28 212.081
R17388 thermo15c_0.XTBN.Y.n169 thermo15c_0.XTBN.Y.t23 212.081
R17389 thermo15c_0.XTBN.Y.n164 thermo15c_0.XTBN.Y.t97 212.081
R17390 thermo15c_0.XTBN.Y.n163 thermo15c_0.XTBN.Y.t95 212.081
R17391 thermo15c_0.XTBN.Y.n110 thermo15c_0.XTBN.Y.t42 212.081
R17392 thermo15c_0.XTBN.Y.n109 thermo15c_0.XTBN.Y.t38 212.081
R17393 thermo15c_0.XTBN.Y.n104 thermo15c_0.XTBN.Y.t119 212.081
R17394 thermo15c_0.XTBN.Y.n103 thermo15c_0.XTBN.Y.t113 212.081
R17395 thermo15c_0.XTBN.Y.n134 thermo15c_0.XTBN.Y.t99 212.081
R17396 thermo15c_0.XTBN.Y.n133 thermo15c_0.XTBN.Y.t96 212.081
R17397 thermo15c_0.XTBN.Y.n128 thermo15c_0.XTBN.Y.t58 212.081
R17398 thermo15c_0.XTBN.Y.n127 thermo15c_0.XTBN.Y.t51 212.081
R17399 thermo15c_0.XTBN.Y.n158 thermo15c_0.XTBN.Y.t13 212.081
R17400 thermo15c_0.XTBN.Y.n157 thermo15c_0.XTBN.Y.t7 212.081
R17401 thermo15c_0.XTBN.Y.n152 thermo15c_0.XTBN.Y.t86 212.081
R17402 thermo15c_0.XTBN.Y.n151 thermo15c_0.XTBN.Y.t81 212.081
R17403 thermo15c_0.XTBN.Y.n192 thermo15c_0.XTBN.Y.n191 208.964
R17404 thermo15c_0.XTBN.Y.n176 thermo15c_0.XTBN.Y.n0 188.516
R17405 thermo15c_0.XTBN.Y.n88 thermo15c_0.XTBN.Y.n87 180.482
R17406 thermo15c_0.XTBN.Y.n62 thermo15c_0.XTBN.Y.n61 180.482
R17407 thermo15c_0.XTBN.Y.n36 thermo15c_0.XTBN.Y.n35 180.482
R17408 thermo15c_0.XTBN.Y.n11 thermo15c_0.XTBN.Y.n10 180.482
R17409 thermo15c_0.XTBN.Y.n75 thermo15c_0.XTBN.Y.n74 180.482
R17410 thermo15c_0.XTBN.Y.n49 thermo15c_0.XTBN.Y.n48 180.482
R17411 thermo15c_0.XTBN.Y.n23 thermo15c_0.XTBN.Y.n22 180.482
R17412 thermo15c_0.XTBN.Y.n95 thermo15c_0.XTBN.Y.n94 173.761
R17413 thermo15c_0.XTBN.Y.n118 thermo15c_0.XTBN.Y.n117 173.761
R17414 thermo15c_0.XTBN.Y.n142 thermo15c_0.XTBN.Y.n141 173.761
R17415 thermo15c_0.XTBN.Y.n166 thermo15c_0.XTBN.Y.n165 173.761
R17416 thermo15c_0.XTBN.Y.n106 thermo15c_0.XTBN.Y.n105 173.761
R17417 thermo15c_0.XTBN.Y.n130 thermo15c_0.XTBN.Y.n129 173.761
R17418 thermo15c_0.XTBN.Y.n154 thermo15c_0.XTBN.Y.n153 173.761
R17419 thermo15c_0.XTBN.Y.n81 thermo15c_0.XTBN.Y.n79 152
R17420 thermo15c_0.XTBN.Y.n84 thermo15c_0.XTBN.Y.n83 152
R17421 thermo15c_0.XTBN.Y.n86 thermo15c_0.XTBN.Y.n85 152
R17422 thermo15c_0.XTBN.Y.n55 thermo15c_0.XTBN.Y.n53 152
R17423 thermo15c_0.XTBN.Y.n58 thermo15c_0.XTBN.Y.n57 152
R17424 thermo15c_0.XTBN.Y.n60 thermo15c_0.XTBN.Y.n59 152
R17425 thermo15c_0.XTBN.Y.n29 thermo15c_0.XTBN.Y.n27 152
R17426 thermo15c_0.XTBN.Y.n32 thermo15c_0.XTBN.Y.n31 152
R17427 thermo15c_0.XTBN.Y.n34 thermo15c_0.XTBN.Y.n33 152
R17428 thermo15c_0.XTBN.Y.n4 thermo15c_0.XTBN.Y.n2 152
R17429 thermo15c_0.XTBN.Y.n7 thermo15c_0.XTBN.Y.n6 152
R17430 thermo15c_0.XTBN.Y.n9 thermo15c_0.XTBN.Y.n8 152
R17431 thermo15c_0.XTBN.Y.n68 thermo15c_0.XTBN.Y.n66 152
R17432 thermo15c_0.XTBN.Y.n71 thermo15c_0.XTBN.Y.n70 152
R17433 thermo15c_0.XTBN.Y.n73 thermo15c_0.XTBN.Y.n72 152
R17434 thermo15c_0.XTBN.Y.n42 thermo15c_0.XTBN.Y.n40 152
R17435 thermo15c_0.XTBN.Y.n45 thermo15c_0.XTBN.Y.n44 152
R17436 thermo15c_0.XTBN.Y.n47 thermo15c_0.XTBN.Y.n46 152
R17437 thermo15c_0.XTBN.Y.n16 thermo15c_0.XTBN.Y.n14 152
R17438 thermo15c_0.XTBN.Y.n19 thermo15c_0.XTBN.Y.n18 152
R17439 thermo15c_0.XTBN.Y.n21 thermo15c_0.XTBN.Y.n20 152
R17440 thermo15c_0.XTBN.Y.n95 thermo15c_0.XTBN.Y.n91 152
R17441 thermo15c_0.XTBN.Y.n97 thermo15c_0.XTBN.Y.n96 152
R17442 thermo15c_0.XTBN.Y.n101 thermo15c_0.XTBN.Y.n100 152
R17443 thermo15c_0.XTBN.Y.n118 thermo15c_0.XTBN.Y.n114 152
R17444 thermo15c_0.XTBN.Y.n120 thermo15c_0.XTBN.Y.n119 152
R17445 thermo15c_0.XTBN.Y.n124 thermo15c_0.XTBN.Y.n123 152
R17446 thermo15c_0.XTBN.Y.n142 thermo15c_0.XTBN.Y.n138 152
R17447 thermo15c_0.XTBN.Y.n144 thermo15c_0.XTBN.Y.n143 152
R17448 thermo15c_0.XTBN.Y.n148 thermo15c_0.XTBN.Y.n147 152
R17449 thermo15c_0.XTBN.Y.n166 thermo15c_0.XTBN.Y.n162 152
R17450 thermo15c_0.XTBN.Y.n168 thermo15c_0.XTBN.Y.n167 152
R17451 thermo15c_0.XTBN.Y.n172 thermo15c_0.XTBN.Y.n171 152
R17452 thermo15c_0.XTBN.Y.n106 thermo15c_0.XTBN.Y.n102 152
R17453 thermo15c_0.XTBN.Y.n108 thermo15c_0.XTBN.Y.n107 152
R17454 thermo15c_0.XTBN.Y.n112 thermo15c_0.XTBN.Y.n111 152
R17455 thermo15c_0.XTBN.Y.n130 thermo15c_0.XTBN.Y.n126 152
R17456 thermo15c_0.XTBN.Y.n132 thermo15c_0.XTBN.Y.n131 152
R17457 thermo15c_0.XTBN.Y.n136 thermo15c_0.XTBN.Y.n135 152
R17458 thermo15c_0.XTBN.Y.n154 thermo15c_0.XTBN.Y.n150 152
R17459 thermo15c_0.XTBN.Y.n156 thermo15c_0.XTBN.Y.n155 152
R17460 thermo15c_0.XTBN.Y.n160 thermo15c_0.XTBN.Y.n159 152
R17461 thermo15c_0.XTBN.Y.n178 thermo15c_0.XTBN.Y.n177 152
R17462 thermo15c_0.XTBN.Y.n180 thermo15c_0.XTBN.Y.n179 152
R17463 thermo15c_0.XTBN.Y.n184 thermo15c_0.XTBN.Y.n183 152
R17464 thermo15c_0.XTBN.Y.n182 thermo15c_0.XTBN.Y.t14 139.78
R17465 thermo15c_0.XTBN.Y.n181 thermo15c_0.XTBN.Y.t105 139.78
R17466 thermo15c_0.XTBN.Y.n175 thermo15c_0.XTBN.Y.t69 139.78
R17467 thermo15c_0.XTBN.Y.n176 thermo15c_0.XTBN.Y.t61 139.78
R17468 thermo15c_0.XTBN.Y.n87 thermo15c_0.XTBN.Y.t123 139.78
R17469 thermo15c_0.XTBN.Y.n78 thermo15c_0.XTBN.Y.t85 139.78
R17470 thermo15c_0.XTBN.Y.n82 thermo15c_0.XTBN.Y.t74 139.78
R17471 thermo15c_0.XTBN.Y.n80 thermo15c_0.XTBN.Y.t65 139.78
R17472 thermo15c_0.XTBN.Y.n61 thermo15c_0.XTBN.Y.t31 139.78
R17473 thermo15c_0.XTBN.Y.n52 thermo15c_0.XTBN.Y.t104 139.78
R17474 thermo15c_0.XTBN.Y.n56 thermo15c_0.XTBN.Y.t94 139.78
R17475 thermo15c_0.XTBN.Y.n54 thermo15c_0.XTBN.Y.t92 139.78
R17476 thermo15c_0.XTBN.Y.n35 thermo15c_0.XTBN.Y.t89 139.78
R17477 thermo15c_0.XTBN.Y.n26 thermo15c_0.XTBN.Y.t41 139.78
R17478 thermo15c_0.XTBN.Y.n30 thermo15c_0.XTBN.Y.t35 139.78
R17479 thermo15c_0.XTBN.Y.n28 thermo15c_0.XTBN.Y.t32 139.78
R17480 thermo15c_0.XTBN.Y.n10 thermo15c_0.XTBN.Y.t118 139.78
R17481 thermo15c_0.XTBN.Y.n1 thermo15c_0.XTBN.Y.t83 139.78
R17482 thermo15c_0.XTBN.Y.n5 thermo15c_0.XTBN.Y.t71 139.78
R17483 thermo15c_0.XTBN.Y.n3 thermo15c_0.XTBN.Y.t62 139.78
R17484 thermo15c_0.XTBN.Y.n74 thermo15c_0.XTBN.Y.t107 139.78
R17485 thermo15c_0.XTBN.Y.n65 thermo15c_0.XTBN.Y.t72 139.78
R17486 thermo15c_0.XTBN.Y.n69 thermo15c_0.XTBN.Y.t57 139.78
R17487 thermo15c_0.XTBN.Y.n67 thermo15c_0.XTBN.Y.t49 139.78
R17488 thermo15c_0.XTBN.Y.n48 thermo15c_0.XTBN.Y.t43 139.78
R17489 thermo15c_0.XTBN.Y.n39 thermo15c_0.XTBN.Y.t10 139.78
R17490 thermo15c_0.XTBN.Y.n43 thermo15c_0.XTBN.Y.t112 139.78
R17491 thermo15c_0.XTBN.Y.n41 thermo15c_0.XTBN.Y.t108 139.78
R17492 thermo15c_0.XTBN.Y.n22 thermo15c_0.XTBN.Y.t121 139.78
R17493 thermo15c_0.XTBN.Y.n13 thermo15c_0.XTBN.Y.t84 139.78
R17494 thermo15c_0.XTBN.Y.n17 thermo15c_0.XTBN.Y.t73 139.78
R17495 thermo15c_0.XTBN.Y.n15 thermo15c_0.XTBN.Y.t64 139.78
R17496 thermo15c_0.XTBN.Y.n99 thermo15c_0.XTBN.Y.t76 139.78
R17497 thermo15c_0.XTBN.Y.n98 thermo15c_0.XTBN.Y.t67 139.78
R17498 thermo15c_0.XTBN.Y.n93 thermo15c_0.XTBN.Y.t29 139.78
R17499 thermo15c_0.XTBN.Y.n92 thermo15c_0.XTBN.Y.t24 139.78
R17500 thermo15c_0.XTBN.Y.n122 thermo15c_0.XTBN.Y.t15 139.78
R17501 thermo15c_0.XTBN.Y.n121 thermo15c_0.XTBN.Y.t8 139.78
R17502 thermo15c_0.XTBN.Y.n116 thermo15c_0.XTBN.Y.t87 139.78
R17503 thermo15c_0.XTBN.Y.n115 thermo15c_0.XTBN.Y.t82 139.78
R17504 thermo15c_0.XTBN.Y.n146 thermo15c_0.XTBN.Y.t66 139.78
R17505 thermo15c_0.XTBN.Y.n145 thermo15c_0.XTBN.Y.t60 139.78
R17506 thermo15c_0.XTBN.Y.n140 thermo15c_0.XTBN.Y.t22 139.78
R17507 thermo15c_0.XTBN.Y.n139 thermo15c_0.XTBN.Y.t20 139.78
R17508 thermo15c_0.XTBN.Y.n170 thermo15c_0.XTBN.Y.t4 139.78
R17509 thermo15c_0.XTBN.Y.n169 thermo15c_0.XTBN.Y.t117 139.78
R17510 thermo15c_0.XTBN.Y.n164 thermo15c_0.XTBN.Y.t80 139.78
R17511 thermo15c_0.XTBN.Y.n163 thermo15c_0.XTBN.Y.t78 139.78
R17512 thermo15c_0.XTBN.Y.n110 thermo15c_0.XTBN.Y.t59 139.78
R17513 thermo15c_0.XTBN.Y.n109 thermo15c_0.XTBN.Y.t55 139.78
R17514 thermo15c_0.XTBN.Y.n104 thermo15c_0.XTBN.Y.t19 139.78
R17515 thermo15c_0.XTBN.Y.n103 thermo15c_0.XTBN.Y.t16 139.78
R17516 thermo15c_0.XTBN.Y.n134 thermo15c_0.XTBN.Y.t115 139.78
R17517 thermo15c_0.XTBN.Y.n133 thermo15c_0.XTBN.Y.t110 139.78
R17518 thermo15c_0.XTBN.Y.n128 thermo15c_0.XTBN.Y.t77 139.78
R17519 thermo15c_0.XTBN.Y.n127 thermo15c_0.XTBN.Y.t68 139.78
R17520 thermo15c_0.XTBN.Y.n158 thermo15c_0.XTBN.Y.t53 139.78
R17521 thermo15c_0.XTBN.Y.n157 thermo15c_0.XTBN.Y.t45 139.78
R17522 thermo15c_0.XTBN.Y.n152 thermo15c_0.XTBN.Y.t11 139.78
R17523 thermo15c_0.XTBN.Y.n151 thermo15c_0.XTBN.Y.t5 139.78
R17524 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n188 96.8352
R17525 thermo15c_0.XTBN.Y.n187 thermo15c_0.XTBN.Y.n0 64.6909
R17526 thermo15c_0.XTBN.Y.n97 thermo15c_0.XTBN.Y.n91 49.6611
R17527 thermo15c_0.XTBN.Y.n120 thermo15c_0.XTBN.Y.n114 49.6611
R17528 thermo15c_0.XTBN.Y.n144 thermo15c_0.XTBN.Y.n138 49.6611
R17529 thermo15c_0.XTBN.Y.n168 thermo15c_0.XTBN.Y.n162 49.6611
R17530 thermo15c_0.XTBN.Y.n108 thermo15c_0.XTBN.Y.n102 49.6611
R17531 thermo15c_0.XTBN.Y.n132 thermo15c_0.XTBN.Y.n126 49.6611
R17532 thermo15c_0.XTBN.Y.n156 thermo15c_0.XTBN.Y.n150 49.6611
R17533 thermo15c_0.XTBN.Y.n100 thermo15c_0.XTBN.Y.n98 44.549
R17534 thermo15c_0.XTBN.Y.n123 thermo15c_0.XTBN.Y.n121 44.549
R17535 thermo15c_0.XTBN.Y.n147 thermo15c_0.XTBN.Y.n145 44.549
R17536 thermo15c_0.XTBN.Y.n171 thermo15c_0.XTBN.Y.n169 44.549
R17537 thermo15c_0.XTBN.Y.n111 thermo15c_0.XTBN.Y.n109 44.549
R17538 thermo15c_0.XTBN.Y.n135 thermo15c_0.XTBN.Y.n133 44.549
R17539 thermo15c_0.XTBN.Y.n159 thermo15c_0.XTBN.Y.n157 44.549
R17540 thermo15c_0.XTBN.Y.n94 thermo15c_0.XTBN.Y.n93 43.0884
R17541 thermo15c_0.XTBN.Y.n117 thermo15c_0.XTBN.Y.n116 43.0884
R17542 thermo15c_0.XTBN.Y.n141 thermo15c_0.XTBN.Y.n140 43.0884
R17543 thermo15c_0.XTBN.Y.n165 thermo15c_0.XTBN.Y.n164 43.0884
R17544 thermo15c_0.XTBN.Y.n105 thermo15c_0.XTBN.Y.n104 43.0884
R17545 thermo15c_0.XTBN.Y.n129 thermo15c_0.XTBN.Y.n128 43.0884
R17546 thermo15c_0.XTBN.Y.n153 thermo15c_0.XTBN.Y.n152 43.0884
R17547 thermo15c_0.XTBN.Y.n177 thermo15c_0.XTBN.Y.n176 30.6732
R17548 thermo15c_0.XTBN.Y.n177 thermo15c_0.XTBN.Y.n175 30.6732
R17549 thermo15c_0.XTBN.Y.n180 thermo15c_0.XTBN.Y.n175 30.6732
R17550 thermo15c_0.XTBN.Y.n181 thermo15c_0.XTBN.Y.n180 30.6732
R17551 thermo15c_0.XTBN.Y.n183 thermo15c_0.XTBN.Y.n181 30.6732
R17552 thermo15c_0.XTBN.Y.n183 thermo15c_0.XTBN.Y.n182 30.6732
R17553 thermo15c_0.XTBN.Y.n81 thermo15c_0.XTBN.Y.n80 30.6732
R17554 thermo15c_0.XTBN.Y.n82 thermo15c_0.XTBN.Y.n81 30.6732
R17555 thermo15c_0.XTBN.Y.n83 thermo15c_0.XTBN.Y.n82 30.6732
R17556 thermo15c_0.XTBN.Y.n83 thermo15c_0.XTBN.Y.n78 30.6732
R17557 thermo15c_0.XTBN.Y.n86 thermo15c_0.XTBN.Y.n78 30.6732
R17558 thermo15c_0.XTBN.Y.n87 thermo15c_0.XTBN.Y.n86 30.6732
R17559 thermo15c_0.XTBN.Y.n55 thermo15c_0.XTBN.Y.n54 30.6732
R17560 thermo15c_0.XTBN.Y.n56 thermo15c_0.XTBN.Y.n55 30.6732
R17561 thermo15c_0.XTBN.Y.n57 thermo15c_0.XTBN.Y.n56 30.6732
R17562 thermo15c_0.XTBN.Y.n57 thermo15c_0.XTBN.Y.n52 30.6732
R17563 thermo15c_0.XTBN.Y.n60 thermo15c_0.XTBN.Y.n52 30.6732
R17564 thermo15c_0.XTBN.Y.n61 thermo15c_0.XTBN.Y.n60 30.6732
R17565 thermo15c_0.XTBN.Y.n29 thermo15c_0.XTBN.Y.n28 30.6732
R17566 thermo15c_0.XTBN.Y.n30 thermo15c_0.XTBN.Y.n29 30.6732
R17567 thermo15c_0.XTBN.Y.n31 thermo15c_0.XTBN.Y.n30 30.6732
R17568 thermo15c_0.XTBN.Y.n31 thermo15c_0.XTBN.Y.n26 30.6732
R17569 thermo15c_0.XTBN.Y.n34 thermo15c_0.XTBN.Y.n26 30.6732
R17570 thermo15c_0.XTBN.Y.n35 thermo15c_0.XTBN.Y.n34 30.6732
R17571 thermo15c_0.XTBN.Y.n4 thermo15c_0.XTBN.Y.n3 30.6732
R17572 thermo15c_0.XTBN.Y.n5 thermo15c_0.XTBN.Y.n4 30.6732
R17573 thermo15c_0.XTBN.Y.n6 thermo15c_0.XTBN.Y.n5 30.6732
R17574 thermo15c_0.XTBN.Y.n6 thermo15c_0.XTBN.Y.n1 30.6732
R17575 thermo15c_0.XTBN.Y.n9 thermo15c_0.XTBN.Y.n1 30.6732
R17576 thermo15c_0.XTBN.Y.n10 thermo15c_0.XTBN.Y.n9 30.6732
R17577 thermo15c_0.XTBN.Y.n68 thermo15c_0.XTBN.Y.n67 30.6732
R17578 thermo15c_0.XTBN.Y.n69 thermo15c_0.XTBN.Y.n68 30.6732
R17579 thermo15c_0.XTBN.Y.n70 thermo15c_0.XTBN.Y.n69 30.6732
R17580 thermo15c_0.XTBN.Y.n70 thermo15c_0.XTBN.Y.n65 30.6732
R17581 thermo15c_0.XTBN.Y.n73 thermo15c_0.XTBN.Y.n65 30.6732
R17582 thermo15c_0.XTBN.Y.n74 thermo15c_0.XTBN.Y.n73 30.6732
R17583 thermo15c_0.XTBN.Y.n42 thermo15c_0.XTBN.Y.n41 30.6732
R17584 thermo15c_0.XTBN.Y.n43 thermo15c_0.XTBN.Y.n42 30.6732
R17585 thermo15c_0.XTBN.Y.n44 thermo15c_0.XTBN.Y.n43 30.6732
R17586 thermo15c_0.XTBN.Y.n44 thermo15c_0.XTBN.Y.n39 30.6732
R17587 thermo15c_0.XTBN.Y.n47 thermo15c_0.XTBN.Y.n39 30.6732
R17588 thermo15c_0.XTBN.Y.n48 thermo15c_0.XTBN.Y.n47 30.6732
R17589 thermo15c_0.XTBN.Y.n16 thermo15c_0.XTBN.Y.n15 30.6732
R17590 thermo15c_0.XTBN.Y.n17 thermo15c_0.XTBN.Y.n16 30.6732
R17591 thermo15c_0.XTBN.Y.n18 thermo15c_0.XTBN.Y.n17 30.6732
R17592 thermo15c_0.XTBN.Y.n18 thermo15c_0.XTBN.Y.n13 30.6732
R17593 thermo15c_0.XTBN.Y.n21 thermo15c_0.XTBN.Y.n13 30.6732
R17594 thermo15c_0.XTBN.Y.n22 thermo15c_0.XTBN.Y.n21 30.6732
R17595 thermo15c_0.XTBN.Y.n191 thermo15c_0.XTBN.Y.t0 26.5955
R17596 thermo15c_0.XTBN.Y.n191 thermo15c_0.XTBN.Y.t1 26.5955
R17597 thermo15c_0.XTBN.Y.n188 thermo15c_0.XTBN.Y.t3 24.9236
R17598 thermo15c_0.XTBN.Y.n188 thermo15c_0.XTBN.Y.t2 24.9236
R17599 thermo15c_0.XTBN.Y.n96 thermo15c_0.XTBN.Y.n95 21.7605
R17600 thermo15c_0.XTBN.Y.n119 thermo15c_0.XTBN.Y.n118 21.7605
R17601 thermo15c_0.XTBN.Y.n143 thermo15c_0.XTBN.Y.n142 21.7605
R17602 thermo15c_0.XTBN.Y.n167 thermo15c_0.XTBN.Y.n166 21.7605
R17603 thermo15c_0.XTBN.Y.n107 thermo15c_0.XTBN.Y.n106 21.7605
R17604 thermo15c_0.XTBN.Y.n131 thermo15c_0.XTBN.Y.n130 21.7605
R17605 thermo15c_0.XTBN.Y.n155 thermo15c_0.XTBN.Y.n154 21.7605
R17606 thermo15c_0.XTBN.Y.n84 thermo15c_0.XTBN.Y.n79 21.5045
R17607 thermo15c_0.XTBN.Y.n58 thermo15c_0.XTBN.Y.n53 21.5045
R17608 thermo15c_0.XTBN.Y.n32 thermo15c_0.XTBN.Y.n27 21.5045
R17609 thermo15c_0.XTBN.Y.n7 thermo15c_0.XTBN.Y.n2 21.5045
R17610 thermo15c_0.XTBN.Y.n71 thermo15c_0.XTBN.Y.n66 21.5045
R17611 thermo15c_0.XTBN.Y.n45 thermo15c_0.XTBN.Y.n40 21.5045
R17612 thermo15c_0.XTBN.Y.n19 thermo15c_0.XTBN.Y.n14 21.5045
R17613 thermo15c_0.XTBN.Y.n178 thermo15c_0.XTBN.Y 21.2485
R17614 thermo15c_0.XTBN.Y.n85 thermo15c_0.XTBN.Y 19.9685
R17615 thermo15c_0.XTBN.Y.n59 thermo15c_0.XTBN.Y 19.9685
R17616 thermo15c_0.XTBN.Y.n33 thermo15c_0.XTBN.Y 19.9685
R17617 thermo15c_0.XTBN.Y.n8 thermo15c_0.XTBN.Y 19.9685
R17618 thermo15c_0.XTBN.Y.n72 thermo15c_0.XTBN.Y 19.9685
R17619 thermo15c_0.XTBN.Y.n46 thermo15c_0.XTBN.Y 19.9685
R17620 thermo15c_0.XTBN.Y.n20 thermo15c_0.XTBN.Y 19.9685
R17621 thermo15c_0.XTBN.Y.n179 thermo15c_0.XTBN.Y 19.2005
R17622 thermo15c_0.XTBN.Y.n94 thermo15c_0.XTBN.Y.n92 18.2581
R17623 thermo15c_0.XTBN.Y.n117 thermo15c_0.XTBN.Y.n115 18.2581
R17624 thermo15c_0.XTBN.Y.n141 thermo15c_0.XTBN.Y.n139 18.2581
R17625 thermo15c_0.XTBN.Y.n165 thermo15c_0.XTBN.Y.n163 18.2581
R17626 thermo15c_0.XTBN.Y.n105 thermo15c_0.XTBN.Y.n103 18.2581
R17627 thermo15c_0.XTBN.Y.n129 thermo15c_0.XTBN.Y.n127 18.2581
R17628 thermo15c_0.XTBN.Y.n153 thermo15c_0.XTBN.Y.n151 18.2581
R17629 thermo15c_0.XTBN.Y.n113 thermo15c_0.XTBN.Y.n101 17.1655
R17630 thermo15c_0.XTBN.Y.n88 thermo15c_0.XTBN.Y 17.1525
R17631 thermo15c_0.XTBN.Y.n62 thermo15c_0.XTBN.Y 17.1525
R17632 thermo15c_0.XTBN.Y.n36 thermo15c_0.XTBN.Y 17.1525
R17633 thermo15c_0.XTBN.Y.n11 thermo15c_0.XTBN.Y 17.1525
R17634 thermo15c_0.XTBN.Y.n75 thermo15c_0.XTBN.Y 17.1525
R17635 thermo15c_0.XTBN.Y.n49 thermo15c_0.XTBN.Y 17.1525
R17636 thermo15c_0.XTBN.Y.n23 thermo15c_0.XTBN.Y 17.1525
R17637 thermo15c_0.XTBN.Y.n100 thermo15c_0.XTBN.Y.n99 16.7975
R17638 thermo15c_0.XTBN.Y.n123 thermo15c_0.XTBN.Y.n122 16.7975
R17639 thermo15c_0.XTBN.Y.n147 thermo15c_0.XTBN.Y.n146 16.7975
R17640 thermo15c_0.XTBN.Y.n171 thermo15c_0.XTBN.Y.n170 16.7975
R17641 thermo15c_0.XTBN.Y.n111 thermo15c_0.XTBN.Y.n110 16.7975
R17642 thermo15c_0.XTBN.Y.n135 thermo15c_0.XTBN.Y.n134 16.7975
R17643 thermo15c_0.XTBN.Y.n159 thermo15c_0.XTBN.Y.n158 16.7975
R17644 thermo15c_0.XTBN.Y.n125 thermo15c_0.XTBN.Y.n124 16.0405
R17645 thermo15c_0.XTBN.Y.n149 thermo15c_0.XTBN.Y.n148 16.0405
R17646 thermo15c_0.XTBN.Y.n173 thermo15c_0.XTBN.Y.n172 16.0405
R17647 thermo15c_0.XTBN.Y.n113 thermo15c_0.XTBN.Y.n112 16.0405
R17648 thermo15c_0.XTBN.Y.n137 thermo15c_0.XTBN.Y.n136 16.0405
R17649 thermo15c_0.XTBN.Y.n161 thermo15c_0.XTBN.Y.n160 16.0405
R17650 thermo15c_0.XTBN.Y.n25 thermo15c_0.XTBN.Y.n12 15.262
R17651 thermo15c_0.XTBN.Y.n101 thermo15c_0.XTBN.Y 15.0405
R17652 thermo15c_0.XTBN.Y.n124 thermo15c_0.XTBN.Y 15.0405
R17653 thermo15c_0.XTBN.Y.n148 thermo15c_0.XTBN.Y 15.0405
R17654 thermo15c_0.XTBN.Y.n172 thermo15c_0.XTBN.Y 15.0405
R17655 thermo15c_0.XTBN.Y.n112 thermo15c_0.XTBN.Y 15.0405
R17656 thermo15c_0.XTBN.Y.n136 thermo15c_0.XTBN.Y 15.0405
R17657 thermo15c_0.XTBN.Y.n160 thermo15c_0.XTBN.Y 15.0405
R17658 thermo15c_0.XTBN.Y.n90 thermo15c_0.XTBN.Y.n89 13.8005
R17659 thermo15c_0.XTBN.Y.n64 thermo15c_0.XTBN.Y.n63 13.8005
R17660 thermo15c_0.XTBN.Y.n38 thermo15c_0.XTBN.Y.n37 13.8005
R17661 thermo15c_0.XTBN.Y.n77 thermo15c_0.XTBN.Y.n76 13.8005
R17662 thermo15c_0.XTBN.Y.n51 thermo15c_0.XTBN.Y.n50 13.8005
R17663 thermo15c_0.XTBN.Y.n25 thermo15c_0.XTBN.Y.n24 13.8005
R17664 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n190 12.5445
R17665 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n189 11.2645
R17666 thermo15c_0.XTBN.Y.n185 thermo15c_0.XTBN.Y.n184 9.2165
R17667 thermo15c_0.XTBN.Y.n185 thermo15c_0.XTBN.Y 7.9365
R17668 thermo15c_0.XTBN.Y.n96 thermo15c_0.XTBN.Y 6.7205
R17669 thermo15c_0.XTBN.Y.n119 thermo15c_0.XTBN.Y 6.7205
R17670 thermo15c_0.XTBN.Y.n143 thermo15c_0.XTBN.Y 6.7205
R17671 thermo15c_0.XTBN.Y.n167 thermo15c_0.XTBN.Y 6.7205
R17672 thermo15c_0.XTBN.Y.n107 thermo15c_0.XTBN.Y 6.7205
R17673 thermo15c_0.XTBN.Y.n131 thermo15c_0.XTBN.Y 6.7205
R17674 thermo15c_0.XTBN.Y.n155 thermo15c_0.XTBN.Y 6.7205
R17675 thermo15c_0.XTBN.Y.n93 thermo15c_0.XTBN.Y.n91 6.57323
R17676 thermo15c_0.XTBN.Y.n116 thermo15c_0.XTBN.Y.n114 6.57323
R17677 thermo15c_0.XTBN.Y.n140 thermo15c_0.XTBN.Y.n138 6.57323
R17678 thermo15c_0.XTBN.Y.n164 thermo15c_0.XTBN.Y.n162 6.57323
R17679 thermo15c_0.XTBN.Y.n104 thermo15c_0.XTBN.Y.n102 6.57323
R17680 thermo15c_0.XTBN.Y.n128 thermo15c_0.XTBN.Y.n126 6.57323
R17681 thermo15c_0.XTBN.Y.n152 thermo15c_0.XTBN.Y.n150 6.57323
R17682 thermo15c_0.XTBN.Y.n184 thermo15c_0.XTBN.Y 6.4005
R17683 thermo15c_0.XTBN.Y.n189 thermo15c_0.XTBN.Y 6.1445
R17684 thermo15c_0.XTBN.Y.n187 thermo15c_0.XTBN.Y.n186 5.74665
R17685 thermo15c_0.XTBN.Y.n186 thermo15c_0.XTBN.Y.n174 5.68319
R17686 thermo15c_0.XTBN.Y.n98 thermo15c_0.XTBN.Y.n97 5.11262
R17687 thermo15c_0.XTBN.Y.n121 thermo15c_0.XTBN.Y.n120 5.11262
R17688 thermo15c_0.XTBN.Y.n145 thermo15c_0.XTBN.Y.n144 5.11262
R17689 thermo15c_0.XTBN.Y.n169 thermo15c_0.XTBN.Y.n168 5.11262
R17690 thermo15c_0.XTBN.Y.n109 thermo15c_0.XTBN.Y.n108 5.11262
R17691 thermo15c_0.XTBN.Y.n133 thermo15c_0.XTBN.Y.n132 5.11262
R17692 thermo15c_0.XTBN.Y.n157 thermo15c_0.XTBN.Y.n156 5.11262
R17693 thermo15c_0.XTBN.Y.n190 thermo15c_0.XTBN.Y.n187 5.06717
R17694 thermo15c_0.XTBN.Y.n190 thermo15c_0.XTBN.Y 4.8645
R17695 thermo15c_0.XTBN.Y.n189 thermo15c_0.XTBN.Y 4.65505
R17696 thermo15c_0.XTBN.Y.n186 thermo15c_0.XTBN.Y.n185 4.6505
R17697 thermo15c_0.XTBN.Y.n89 thermo15c_0.XTBN.Y 4.6085
R17698 thermo15c_0.XTBN.Y.n63 thermo15c_0.XTBN.Y 4.6085
R17699 thermo15c_0.XTBN.Y.n37 thermo15c_0.XTBN.Y 4.6085
R17700 thermo15c_0.XTBN.Y.n12 thermo15c_0.XTBN.Y 4.6085
R17701 thermo15c_0.XTBN.Y.n76 thermo15c_0.XTBN.Y 4.6085
R17702 thermo15c_0.XTBN.Y.n50 thermo15c_0.XTBN.Y 4.6085
R17703 thermo15c_0.XTBN.Y.n24 thermo15c_0.XTBN.Y 4.6085
R17704 thermo15c_0.XTBN.Y.n179 thermo15c_0.XTBN.Y 4.3525
R17705 thermo15c_0.XTBN.Y.n85 thermo15c_0.XTBN.Y 3.5845
R17706 thermo15c_0.XTBN.Y.n59 thermo15c_0.XTBN.Y 3.5845
R17707 thermo15c_0.XTBN.Y.n33 thermo15c_0.XTBN.Y 3.5845
R17708 thermo15c_0.XTBN.Y.n8 thermo15c_0.XTBN.Y 3.5845
R17709 thermo15c_0.XTBN.Y.n72 thermo15c_0.XTBN.Y 3.5845
R17710 thermo15c_0.XTBN.Y.n46 thermo15c_0.XTBN.Y 3.5845
R17711 thermo15c_0.XTBN.Y.n20 thermo15c_0.XTBN.Y 3.5845
R17712 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n0 2.3045
R17713 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n178 2.3045
R17714 thermo15c_0.XTBN.Y.n192 thermo15c_0.XTBN.Y 2.0485
R17715 thermo15c_0.XTBN.Y.n89 thermo15c_0.XTBN.Y.n88 1.7925
R17716 thermo15c_0.XTBN.Y.n63 thermo15c_0.XTBN.Y.n62 1.7925
R17717 thermo15c_0.XTBN.Y.n37 thermo15c_0.XTBN.Y.n36 1.7925
R17718 thermo15c_0.XTBN.Y.n12 thermo15c_0.XTBN.Y.n11 1.7925
R17719 thermo15c_0.XTBN.Y.n76 thermo15c_0.XTBN.Y.n75 1.7925
R17720 thermo15c_0.XTBN.Y.n50 thermo15c_0.XTBN.Y.n49 1.7925
R17721 thermo15c_0.XTBN.Y.n24 thermo15c_0.XTBN.Y.n23 1.7925
R17722 thermo15c_0.XTBN.Y.n174 thermo15c_0.XTBN.Y.n173 1.59665
R17723 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n192 1.55202
R17724 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n84 1.5365
R17725 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n58 1.5365
R17726 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n32 1.5365
R17727 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n7 1.5365
R17728 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n71 1.5365
R17729 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n45 1.5365
R17730 thermo15c_0.XTBN.Y thermo15c_0.XTBN.Y.n19 1.5365
R17731 thermo15c_0.XTBN.Y.n149 thermo15c_0.XTBN.Y.n137 1.49088
R17732 thermo15c_0.XTBN.Y.n125 thermo15c_0.XTBN.Y.n113 1.49088
R17733 thermo15c_0.XTBN.Y.n173 thermo15c_0.XTBN.Y.n161 1.48608
R17734 thermo15c_0.XTBN.Y.n51 thermo15c_0.XTBN.Y.n38 1.46204
R17735 thermo15c_0.XTBN.Y.n77 thermo15c_0.XTBN.Y.n64 1.46204
R17736 thermo15c_0.XTBN.Y.n38 thermo15c_0.XTBN.Y.n25 1.15435
R17737 thermo15c_0.XTBN.Y.n64 thermo15c_0.XTBN.Y.n51 1.15435
R17738 thermo15c_0.XTBN.Y.n90 thermo15c_0.XTBN.Y.n77 1.15435
R17739 thermo15c_0.XTBN.Y.n174 thermo15c_0.XTBN.Y.n90 1.14473
R17740 thermo15c_0.XTBN.Y.n161 thermo15c_0.XTBN.Y.n149 1.13031
R17741 thermo15c_0.XTBN.Y.n137 thermo15c_0.XTBN.Y.n125 1.1255
R17742 thermo15c_0.XTBN.Y.n79 thermo15c_0.XTBN.Y 0.5125
R17743 thermo15c_0.XTBN.Y.n53 thermo15c_0.XTBN.Y 0.5125
R17744 thermo15c_0.XTBN.Y.n27 thermo15c_0.XTBN.Y 0.5125
R17745 thermo15c_0.XTBN.Y.n2 thermo15c_0.XTBN.Y 0.5125
R17746 thermo15c_0.XTBN.Y.n66 thermo15c_0.XTBN.Y 0.5125
R17747 thermo15c_0.XTBN.Y.n40 thermo15c_0.XTBN.Y 0.5125
R17748 thermo15c_0.XTBN.Y.n14 thermo15c_0.XTBN.Y 0.5125
R17749 XA.Cn[6].n59 XA.Cn[6].n57 332.332
R17750 XA.Cn[6].n59 XA.Cn[6].n58 296.493
R17751 XA.Cn[6].n9 XA.Cn[6].n7 161.406
R17752 XA.Cn[6].n12 XA.Cn[6].n10 161.406
R17753 XA.Cn[6].n15 XA.Cn[6].n13 161.406
R17754 XA.Cn[6].n18 XA.Cn[6].n16 161.406
R17755 XA.Cn[6].n21 XA.Cn[6].n19 161.406
R17756 XA.Cn[6].n24 XA.Cn[6].n22 161.406
R17757 XA.Cn[6].n27 XA.Cn[6].n25 161.406
R17758 XA.Cn[6].n30 XA.Cn[6].n28 161.406
R17759 XA.Cn[6].n33 XA.Cn[6].n31 161.406
R17760 XA.Cn[6].n36 XA.Cn[6].n34 161.406
R17761 XA.Cn[6].n39 XA.Cn[6].n37 161.406
R17762 XA.Cn[6].n42 XA.Cn[6].n40 161.406
R17763 XA.Cn[6].n45 XA.Cn[6].n43 161.406
R17764 XA.Cn[6].n48 XA.Cn[6].n46 161.406
R17765 XA.Cn[6].n51 XA.Cn[6].n49 161.406
R17766 XA.Cn[6].n54 XA.Cn[6].n52 161.406
R17767 XA.Cn[6].n7 XA.Cn[6].t26 161.202
R17768 XA.Cn[6].n10 XA.Cn[6].t13 161.202
R17769 XA.Cn[6].n13 XA.Cn[6].t17 161.202
R17770 XA.Cn[6].n16 XA.Cn[6].t18 161.202
R17771 XA.Cn[6].n19 XA.Cn[6].t37 161.202
R17772 XA.Cn[6].n22 XA.Cn[6].t38 161.202
R17773 XA.Cn[6].n25 XA.Cn[6].t22 161.202
R17774 XA.Cn[6].n28 XA.Cn[6].t29 161.202
R17775 XA.Cn[6].n31 XA.Cn[6].t31 161.202
R17776 XA.Cn[6].n34 XA.Cn[6].t19 161.202
R17777 XA.Cn[6].n37 XA.Cn[6].t21 161.202
R17778 XA.Cn[6].n40 XA.Cn[6].t32 161.202
R17779 XA.Cn[6].n43 XA.Cn[6].t41 161.202
R17780 XA.Cn[6].n46 XA.Cn[6].t43 161.202
R17781 XA.Cn[6].n49 XA.Cn[6].t24 161.202
R17782 XA.Cn[6].n52 XA.Cn[6].t34 161.202
R17783 XA.Cn[6].n7 XA.Cn[6].t23 145.137
R17784 XA.Cn[6].n10 XA.Cn[6].t40 145.137
R17785 XA.Cn[6].n13 XA.Cn[6].t42 145.137
R17786 XA.Cn[6].n16 XA.Cn[6].t12 145.137
R17787 XA.Cn[6].n19 XA.Cn[6].t33 145.137
R17788 XA.Cn[6].n22 XA.Cn[6].t35 145.137
R17789 XA.Cn[6].n25 XA.Cn[6].t16 145.137
R17790 XA.Cn[6].n28 XA.Cn[6].t25 145.137
R17791 XA.Cn[6].n31 XA.Cn[6].t27 145.137
R17792 XA.Cn[6].n34 XA.Cn[6].t14 145.137
R17793 XA.Cn[6].n37 XA.Cn[6].t15 145.137
R17794 XA.Cn[6].n40 XA.Cn[6].t28 145.137
R17795 XA.Cn[6].n43 XA.Cn[6].t36 145.137
R17796 XA.Cn[6].n46 XA.Cn[6].t39 145.137
R17797 XA.Cn[6].n49 XA.Cn[6].t20 145.137
R17798 XA.Cn[6].n52 XA.Cn[6].t30 145.137
R17799 XA.Cn[6].n2 XA.Cn[6].n0 135.248
R17800 XA.Cn[6].n2 XA.Cn[6].n1 98.982
R17801 XA.Cn[6].n4 XA.Cn[6].n3 98.982
R17802 XA.Cn[6].n6 XA.Cn[6].n5 98.982
R17803 XA.Cn[6].n4 XA.Cn[6].n2 36.2672
R17804 XA.Cn[6].n6 XA.Cn[6].n4 36.2672
R17805 XA.Cn[6].n56 XA.Cn[6].n6 32.6405
R17806 XA.Cn[6].n57 XA.Cn[6].t1 26.5955
R17807 XA.Cn[6].n57 XA.Cn[6].t0 26.5955
R17808 XA.Cn[6].n58 XA.Cn[6].t3 26.5955
R17809 XA.Cn[6].n58 XA.Cn[6].t2 26.5955
R17810 XA.Cn[6].n0 XA.Cn[6].t11 24.9236
R17811 XA.Cn[6].n0 XA.Cn[6].t10 24.9236
R17812 XA.Cn[6].n1 XA.Cn[6].t9 24.9236
R17813 XA.Cn[6].n1 XA.Cn[6].t8 24.9236
R17814 XA.Cn[6].n3 XA.Cn[6].t6 24.9236
R17815 XA.Cn[6].n3 XA.Cn[6].t5 24.9236
R17816 XA.Cn[6].n5 XA.Cn[6].t4 24.9236
R17817 XA.Cn[6].n5 XA.Cn[6].t7 24.9236
R17818 XA.Cn[6].n60 XA.Cn[6].n59 18.5605
R17819 XA.Cn[6].n60 XA.Cn[6].n56 11.5205
R17820 XA.Cn[6].n56 XA.Cn[6].n55 3.18344
R17821 XA.Cn[6].n55 XA.Cn[6] 3.09179
R17822 XA.Cn[6].n12 XA.Cn[6] 0.931056
R17823 XA.Cn[6].n15 XA.Cn[6] 0.931056
R17824 XA.Cn[6].n18 XA.Cn[6] 0.931056
R17825 XA.Cn[6].n21 XA.Cn[6] 0.931056
R17826 XA.Cn[6].n24 XA.Cn[6] 0.931056
R17827 XA.Cn[6].n27 XA.Cn[6] 0.931056
R17828 XA.Cn[6].n30 XA.Cn[6] 0.931056
R17829 XA.Cn[6].n33 XA.Cn[6] 0.931056
R17830 XA.Cn[6].n36 XA.Cn[6] 0.931056
R17831 XA.Cn[6].n39 XA.Cn[6] 0.931056
R17832 XA.Cn[6].n42 XA.Cn[6] 0.931056
R17833 XA.Cn[6].n45 XA.Cn[6] 0.931056
R17834 XA.Cn[6].n48 XA.Cn[6] 0.931056
R17835 XA.Cn[6].n51 XA.Cn[6] 0.931056
R17836 XA.Cn[6].n54 XA.Cn[6] 0.931056
R17837 XA.Cn[6] XA.Cn[6].n60 0.6405
R17838 XA.Cn[6] XA.Cn[6].n9 0.396333
R17839 XA.Cn[6] XA.Cn[6].n12 0.396333
R17840 XA.Cn[6] XA.Cn[6].n15 0.396333
R17841 XA.Cn[6] XA.Cn[6].n18 0.396333
R17842 XA.Cn[6] XA.Cn[6].n21 0.396333
R17843 XA.Cn[6] XA.Cn[6].n24 0.396333
R17844 XA.Cn[6] XA.Cn[6].n27 0.396333
R17845 XA.Cn[6] XA.Cn[6].n30 0.396333
R17846 XA.Cn[6] XA.Cn[6].n33 0.396333
R17847 XA.Cn[6] XA.Cn[6].n36 0.396333
R17848 XA.Cn[6] XA.Cn[6].n39 0.396333
R17849 XA.Cn[6] XA.Cn[6].n42 0.396333
R17850 XA.Cn[6] XA.Cn[6].n45 0.396333
R17851 XA.Cn[6] XA.Cn[6].n48 0.396333
R17852 XA.Cn[6] XA.Cn[6].n51 0.396333
R17853 XA.Cn[6] XA.Cn[6].n54 0.396333
R17854 XA.Cn[6].n8 XA.Cn[6] 0.104667
R17855 XA.Cn[6].n11 XA.Cn[6] 0.104667
R17856 XA.Cn[6].n14 XA.Cn[6] 0.104667
R17857 XA.Cn[6].n17 XA.Cn[6] 0.104667
R17858 XA.Cn[6].n20 XA.Cn[6] 0.104667
R17859 XA.Cn[6].n23 XA.Cn[6] 0.104667
R17860 XA.Cn[6].n26 XA.Cn[6] 0.104667
R17861 XA.Cn[6].n29 XA.Cn[6] 0.104667
R17862 XA.Cn[6].n32 XA.Cn[6] 0.104667
R17863 XA.Cn[6].n35 XA.Cn[6] 0.104667
R17864 XA.Cn[6].n38 XA.Cn[6] 0.104667
R17865 XA.Cn[6].n41 XA.Cn[6] 0.104667
R17866 XA.Cn[6].n44 XA.Cn[6] 0.104667
R17867 XA.Cn[6].n47 XA.Cn[6] 0.104667
R17868 XA.Cn[6].n50 XA.Cn[6] 0.104667
R17869 XA.Cn[6].n53 XA.Cn[6] 0.104667
R17870 XA.Cn[6].n8 XA.Cn[6] 0.0309878
R17871 XA.Cn[6].n11 XA.Cn[6] 0.0309878
R17872 XA.Cn[6].n14 XA.Cn[6] 0.0309878
R17873 XA.Cn[6].n17 XA.Cn[6] 0.0309878
R17874 XA.Cn[6].n20 XA.Cn[6] 0.0309878
R17875 XA.Cn[6].n23 XA.Cn[6] 0.0309878
R17876 XA.Cn[6].n26 XA.Cn[6] 0.0309878
R17877 XA.Cn[6].n29 XA.Cn[6] 0.0309878
R17878 XA.Cn[6].n32 XA.Cn[6] 0.0309878
R17879 XA.Cn[6].n35 XA.Cn[6] 0.0309878
R17880 XA.Cn[6].n38 XA.Cn[6] 0.0309878
R17881 XA.Cn[6].n41 XA.Cn[6] 0.0309878
R17882 XA.Cn[6].n44 XA.Cn[6] 0.0309878
R17883 XA.Cn[6].n47 XA.Cn[6] 0.0309878
R17884 XA.Cn[6].n50 XA.Cn[6] 0.0309878
R17885 XA.Cn[6].n53 XA.Cn[6] 0.0309878
R17886 XA.Cn[6].n9 XA.Cn[6].n8 0.027939
R17887 XA.Cn[6].n12 XA.Cn[6].n11 0.027939
R17888 XA.Cn[6].n15 XA.Cn[6].n14 0.027939
R17889 XA.Cn[6].n18 XA.Cn[6].n17 0.027939
R17890 XA.Cn[6].n21 XA.Cn[6].n20 0.027939
R17891 XA.Cn[6].n24 XA.Cn[6].n23 0.027939
R17892 XA.Cn[6].n27 XA.Cn[6].n26 0.027939
R17893 XA.Cn[6].n30 XA.Cn[6].n29 0.027939
R17894 XA.Cn[6].n33 XA.Cn[6].n32 0.027939
R17895 XA.Cn[6].n36 XA.Cn[6].n35 0.027939
R17896 XA.Cn[6].n39 XA.Cn[6].n38 0.027939
R17897 XA.Cn[6].n42 XA.Cn[6].n41 0.027939
R17898 XA.Cn[6].n45 XA.Cn[6].n44 0.027939
R17899 XA.Cn[6].n48 XA.Cn[6].n47 0.027939
R17900 XA.Cn[6].n51 XA.Cn[6].n50 0.027939
R17901 XA.Cn[6].n54 XA.Cn[6].n53 0.027939
R17902 XA.Cn[6].n55 XA.Cn[6] 0.0140108
R17903 XThR.Tn[9].n8 XThR.Tn[9].n7 256.104
R17904 XThR.Tn[9].n5 XThR.Tn[9].n3 243.68
R17905 XThR.Tn[9].n2 XThR.Tn[9].n1 241.847
R17906 XThR.Tn[9].n5 XThR.Tn[9].n4 205.28
R17907 XThR.Tn[9].n8 XThR.Tn[9].n6 202.094
R17908 XThR.Tn[9].n2 XThR.Tn[9].n0 185
R17909 XThR.Tn[9] XThR.Tn[9].n82 161.363
R17910 XThR.Tn[9] XThR.Tn[9].n77 161.363
R17911 XThR.Tn[9] XThR.Tn[9].n72 161.363
R17912 XThR.Tn[9] XThR.Tn[9].n67 161.363
R17913 XThR.Tn[9] XThR.Tn[9].n62 161.363
R17914 XThR.Tn[9] XThR.Tn[9].n57 161.363
R17915 XThR.Tn[9] XThR.Tn[9].n52 161.363
R17916 XThR.Tn[9] XThR.Tn[9].n47 161.363
R17917 XThR.Tn[9] XThR.Tn[9].n42 161.363
R17918 XThR.Tn[9] XThR.Tn[9].n37 161.363
R17919 XThR.Tn[9] XThR.Tn[9].n32 161.363
R17920 XThR.Tn[9] XThR.Tn[9].n27 161.363
R17921 XThR.Tn[9] XThR.Tn[9].n22 161.363
R17922 XThR.Tn[9] XThR.Tn[9].n17 161.363
R17923 XThR.Tn[9] XThR.Tn[9].n12 161.363
R17924 XThR.Tn[9] XThR.Tn[9].n10 161.363
R17925 XThR.Tn[9].n84 XThR.Tn[9].n83 161.3
R17926 XThR.Tn[9].n79 XThR.Tn[9].n78 161.3
R17927 XThR.Tn[9].n74 XThR.Tn[9].n73 161.3
R17928 XThR.Tn[9].n69 XThR.Tn[9].n68 161.3
R17929 XThR.Tn[9].n64 XThR.Tn[9].n63 161.3
R17930 XThR.Tn[9].n59 XThR.Tn[9].n58 161.3
R17931 XThR.Tn[9].n54 XThR.Tn[9].n53 161.3
R17932 XThR.Tn[9].n49 XThR.Tn[9].n48 161.3
R17933 XThR.Tn[9].n44 XThR.Tn[9].n43 161.3
R17934 XThR.Tn[9].n39 XThR.Tn[9].n38 161.3
R17935 XThR.Tn[9].n34 XThR.Tn[9].n33 161.3
R17936 XThR.Tn[9].n29 XThR.Tn[9].n28 161.3
R17937 XThR.Tn[9].n24 XThR.Tn[9].n23 161.3
R17938 XThR.Tn[9].n19 XThR.Tn[9].n18 161.3
R17939 XThR.Tn[9].n14 XThR.Tn[9].n13 161.3
R17940 XThR.Tn[9].n82 XThR.Tn[9].t63 161.106
R17941 XThR.Tn[9].n77 XThR.Tn[9].t69 161.106
R17942 XThR.Tn[9].n72 XThR.Tn[9].t47 161.106
R17943 XThR.Tn[9].n67 XThR.Tn[9].t34 161.106
R17944 XThR.Tn[9].n62 XThR.Tn[9].t62 161.106
R17945 XThR.Tn[9].n57 XThR.Tn[9].t24 161.106
R17946 XThR.Tn[9].n52 XThR.Tn[9].t66 161.106
R17947 XThR.Tn[9].n47 XThR.Tn[9].t45 161.106
R17948 XThR.Tn[9].n42 XThR.Tn[9].t32 161.106
R17949 XThR.Tn[9].n37 XThR.Tn[9].t37 161.106
R17950 XThR.Tn[9].n32 XThR.Tn[9].t23 161.106
R17951 XThR.Tn[9].n27 XThR.Tn[9].t46 161.106
R17952 XThR.Tn[9].n22 XThR.Tn[9].t21 161.106
R17953 XThR.Tn[9].n17 XThR.Tn[9].t64 161.106
R17954 XThR.Tn[9].n12 XThR.Tn[9].t28 161.106
R17955 XThR.Tn[9].n10 XThR.Tn[9].t71 161.106
R17956 XThR.Tn[9].n83 XThR.Tn[9].t54 159.978
R17957 XThR.Tn[9].n78 XThR.Tn[9].t61 159.978
R17958 XThR.Tn[9].n73 XThR.Tn[9].t43 159.978
R17959 XThR.Tn[9].n68 XThR.Tn[9].t27 159.978
R17960 XThR.Tn[9].n63 XThR.Tn[9].t52 159.978
R17961 XThR.Tn[9].n58 XThR.Tn[9].t18 159.978
R17962 XThR.Tn[9].n53 XThR.Tn[9].t60 159.978
R17963 XThR.Tn[9].n48 XThR.Tn[9].t40 159.978
R17964 XThR.Tn[9].n43 XThR.Tn[9].t25 159.978
R17965 XThR.Tn[9].n38 XThR.Tn[9].t33 159.978
R17966 XThR.Tn[9].n33 XThR.Tn[9].t16 159.978
R17967 XThR.Tn[9].n28 XThR.Tn[9].t42 159.978
R17968 XThR.Tn[9].n23 XThR.Tn[9].t15 159.978
R17969 XThR.Tn[9].n18 XThR.Tn[9].t59 159.978
R17970 XThR.Tn[9].n13 XThR.Tn[9].t19 159.978
R17971 XThR.Tn[9].n82 XThR.Tn[9].t49 145.038
R17972 XThR.Tn[9].n77 XThR.Tn[9].t14 145.038
R17973 XThR.Tn[9].n72 XThR.Tn[9].t57 145.038
R17974 XThR.Tn[9].n67 XThR.Tn[9].t38 145.038
R17975 XThR.Tn[9].n62 XThR.Tn[9].t70 145.038
R17976 XThR.Tn[9].n57 XThR.Tn[9].t48 145.038
R17977 XThR.Tn[9].n52 XThR.Tn[9].t58 145.038
R17978 XThR.Tn[9].n47 XThR.Tn[9].t39 145.038
R17979 XThR.Tn[9].n42 XThR.Tn[9].t36 145.038
R17980 XThR.Tn[9].n37 XThR.Tn[9].t67 145.038
R17981 XThR.Tn[9].n32 XThR.Tn[9].t31 145.038
R17982 XThR.Tn[9].n27 XThR.Tn[9].t56 145.038
R17983 XThR.Tn[9].n22 XThR.Tn[9].t29 145.038
R17984 XThR.Tn[9].n17 XThR.Tn[9].t72 145.038
R17985 XThR.Tn[9].n12 XThR.Tn[9].t35 145.038
R17986 XThR.Tn[9].n10 XThR.Tn[9].t17 145.038
R17987 XThR.Tn[9].n83 XThR.Tn[9].t68 143.911
R17988 XThR.Tn[9].n78 XThR.Tn[9].t30 143.911
R17989 XThR.Tn[9].n73 XThR.Tn[9].t12 143.911
R17990 XThR.Tn[9].n68 XThR.Tn[9].t53 143.911
R17991 XThR.Tn[9].n63 XThR.Tn[9].t22 143.911
R17992 XThR.Tn[9].n58 XThR.Tn[9].t65 143.911
R17993 XThR.Tn[9].n53 XThR.Tn[9].t13 143.911
R17994 XThR.Tn[9].n48 XThR.Tn[9].t55 143.911
R17995 XThR.Tn[9].n43 XThR.Tn[9].t51 143.911
R17996 XThR.Tn[9].n38 XThR.Tn[9].t20 143.911
R17997 XThR.Tn[9].n33 XThR.Tn[9].t44 143.911
R17998 XThR.Tn[9].n28 XThR.Tn[9].t73 143.911
R17999 XThR.Tn[9].n23 XThR.Tn[9].t41 143.911
R18000 XThR.Tn[9].n18 XThR.Tn[9].t26 143.911
R18001 XThR.Tn[9].n13 XThR.Tn[9].t50 143.911
R18002 XThR.Tn[9] XThR.Tn[9].n5 35.7652
R18003 XThR.Tn[9].n6 XThR.Tn[9].t6 26.5955
R18004 XThR.Tn[9].n6 XThR.Tn[9].t4 26.5955
R18005 XThR.Tn[9].n7 XThR.Tn[9].t7 26.5955
R18006 XThR.Tn[9].n7 XThR.Tn[9].t5 26.5955
R18007 XThR.Tn[9].n3 XThR.Tn[9].t10 26.5955
R18008 XThR.Tn[9].n3 XThR.Tn[9].t8 26.5955
R18009 XThR.Tn[9].n4 XThR.Tn[9].t11 26.5955
R18010 XThR.Tn[9].n4 XThR.Tn[9].t9 26.5955
R18011 XThR.Tn[9].n0 XThR.Tn[9].t0 24.9236
R18012 XThR.Tn[9].n0 XThR.Tn[9].t2 24.9236
R18013 XThR.Tn[9].n1 XThR.Tn[9].t1 24.9236
R18014 XThR.Tn[9].n1 XThR.Tn[9].t3 24.9236
R18015 XThR.Tn[9] XThR.Tn[9].n2 22.9615
R18016 XThR.Tn[9].n9 XThR.Tn[9].n8 13.5534
R18017 XThR.Tn[9].n88 XThR.Tn[9] 7.97984
R18018 XThR.Tn[9] XThR.Tn[9].n11 5.34038
R18019 XThR.Tn[9].n16 XThR.Tn[9].n15 4.5005
R18020 XThR.Tn[9].n21 XThR.Tn[9].n20 4.5005
R18021 XThR.Tn[9].n26 XThR.Tn[9].n25 4.5005
R18022 XThR.Tn[9].n31 XThR.Tn[9].n30 4.5005
R18023 XThR.Tn[9].n36 XThR.Tn[9].n35 4.5005
R18024 XThR.Tn[9].n41 XThR.Tn[9].n40 4.5005
R18025 XThR.Tn[9].n46 XThR.Tn[9].n45 4.5005
R18026 XThR.Tn[9].n51 XThR.Tn[9].n50 4.5005
R18027 XThR.Tn[9].n56 XThR.Tn[9].n55 4.5005
R18028 XThR.Tn[9].n61 XThR.Tn[9].n60 4.5005
R18029 XThR.Tn[9].n66 XThR.Tn[9].n65 4.5005
R18030 XThR.Tn[9].n71 XThR.Tn[9].n70 4.5005
R18031 XThR.Tn[9].n76 XThR.Tn[9].n75 4.5005
R18032 XThR.Tn[9].n81 XThR.Tn[9].n80 4.5005
R18033 XThR.Tn[9].n86 XThR.Tn[9].n85 4.5005
R18034 XThR.Tn[9].n87 XThR.Tn[9] 3.70586
R18035 XThR.Tn[9].n88 XThR.Tn[9].n9 2.99115
R18036 XThR.Tn[9].n9 XThR.Tn[9] 2.87153
R18037 XThR.Tn[9].n16 XThR.Tn[9] 2.52282
R18038 XThR.Tn[9].n21 XThR.Tn[9] 2.52282
R18039 XThR.Tn[9].n26 XThR.Tn[9] 2.52282
R18040 XThR.Tn[9].n31 XThR.Tn[9] 2.52282
R18041 XThR.Tn[9].n36 XThR.Tn[9] 2.52282
R18042 XThR.Tn[9].n41 XThR.Tn[9] 2.52282
R18043 XThR.Tn[9].n46 XThR.Tn[9] 2.52282
R18044 XThR.Tn[9].n51 XThR.Tn[9] 2.52282
R18045 XThR.Tn[9].n56 XThR.Tn[9] 2.52282
R18046 XThR.Tn[9].n61 XThR.Tn[9] 2.52282
R18047 XThR.Tn[9].n66 XThR.Tn[9] 2.52282
R18048 XThR.Tn[9].n71 XThR.Tn[9] 2.52282
R18049 XThR.Tn[9].n76 XThR.Tn[9] 2.52282
R18050 XThR.Tn[9].n81 XThR.Tn[9] 2.52282
R18051 XThR.Tn[9].n86 XThR.Tn[9] 2.52282
R18052 XThR.Tn[9] XThR.Tn[9].n88 2.2734
R18053 XThR.Tn[9].n9 XThR.Tn[9] 1.50638
R18054 XThR.Tn[9].n84 XThR.Tn[9] 1.08677
R18055 XThR.Tn[9].n79 XThR.Tn[9] 1.08677
R18056 XThR.Tn[9].n74 XThR.Tn[9] 1.08677
R18057 XThR.Tn[9].n69 XThR.Tn[9] 1.08677
R18058 XThR.Tn[9].n64 XThR.Tn[9] 1.08677
R18059 XThR.Tn[9].n59 XThR.Tn[9] 1.08677
R18060 XThR.Tn[9].n54 XThR.Tn[9] 1.08677
R18061 XThR.Tn[9].n49 XThR.Tn[9] 1.08677
R18062 XThR.Tn[9].n44 XThR.Tn[9] 1.08677
R18063 XThR.Tn[9].n39 XThR.Tn[9] 1.08677
R18064 XThR.Tn[9].n34 XThR.Tn[9] 1.08677
R18065 XThR.Tn[9].n29 XThR.Tn[9] 1.08677
R18066 XThR.Tn[9].n24 XThR.Tn[9] 1.08677
R18067 XThR.Tn[9].n19 XThR.Tn[9] 1.08677
R18068 XThR.Tn[9].n14 XThR.Tn[9] 1.08677
R18069 XThR.Tn[9] XThR.Tn[9].n16 0.839786
R18070 XThR.Tn[9] XThR.Tn[9].n21 0.839786
R18071 XThR.Tn[9] XThR.Tn[9].n26 0.839786
R18072 XThR.Tn[9] XThR.Tn[9].n31 0.839786
R18073 XThR.Tn[9] XThR.Tn[9].n36 0.839786
R18074 XThR.Tn[9] XThR.Tn[9].n41 0.839786
R18075 XThR.Tn[9] XThR.Tn[9].n46 0.839786
R18076 XThR.Tn[9] XThR.Tn[9].n51 0.839786
R18077 XThR.Tn[9] XThR.Tn[9].n56 0.839786
R18078 XThR.Tn[9] XThR.Tn[9].n61 0.839786
R18079 XThR.Tn[9] XThR.Tn[9].n66 0.839786
R18080 XThR.Tn[9] XThR.Tn[9].n71 0.839786
R18081 XThR.Tn[9] XThR.Tn[9].n76 0.839786
R18082 XThR.Tn[9] XThR.Tn[9].n81 0.839786
R18083 XThR.Tn[9] XThR.Tn[9].n86 0.839786
R18084 XThR.Tn[9].n11 XThR.Tn[9] 0.499542
R18085 XThR.Tn[9].n85 XThR.Tn[9] 0.063
R18086 XThR.Tn[9].n80 XThR.Tn[9] 0.063
R18087 XThR.Tn[9].n75 XThR.Tn[9] 0.063
R18088 XThR.Tn[9].n70 XThR.Tn[9] 0.063
R18089 XThR.Tn[9].n65 XThR.Tn[9] 0.063
R18090 XThR.Tn[9].n60 XThR.Tn[9] 0.063
R18091 XThR.Tn[9].n55 XThR.Tn[9] 0.063
R18092 XThR.Tn[9].n50 XThR.Tn[9] 0.063
R18093 XThR.Tn[9].n45 XThR.Tn[9] 0.063
R18094 XThR.Tn[9].n40 XThR.Tn[9] 0.063
R18095 XThR.Tn[9].n35 XThR.Tn[9] 0.063
R18096 XThR.Tn[9].n30 XThR.Tn[9] 0.063
R18097 XThR.Tn[9].n25 XThR.Tn[9] 0.063
R18098 XThR.Tn[9].n20 XThR.Tn[9] 0.063
R18099 XThR.Tn[9].n15 XThR.Tn[9] 0.063
R18100 XThR.Tn[9].n87 XThR.Tn[9] 0.0540714
R18101 XThR.Tn[9] XThR.Tn[9].n87 0.038
R18102 XThR.Tn[9].n11 XThR.Tn[9] 0.0143889
R18103 XThR.Tn[9].n85 XThR.Tn[9].n84 0.00771154
R18104 XThR.Tn[9].n80 XThR.Tn[9].n79 0.00771154
R18105 XThR.Tn[9].n75 XThR.Tn[9].n74 0.00771154
R18106 XThR.Tn[9].n70 XThR.Tn[9].n69 0.00771154
R18107 XThR.Tn[9].n65 XThR.Tn[9].n64 0.00771154
R18108 XThR.Tn[9].n60 XThR.Tn[9].n59 0.00771154
R18109 XThR.Tn[9].n55 XThR.Tn[9].n54 0.00771154
R18110 XThR.Tn[9].n50 XThR.Tn[9].n49 0.00771154
R18111 XThR.Tn[9].n45 XThR.Tn[9].n44 0.00771154
R18112 XThR.Tn[9].n40 XThR.Tn[9].n39 0.00771154
R18113 XThR.Tn[9].n35 XThR.Tn[9].n34 0.00771154
R18114 XThR.Tn[9].n30 XThR.Tn[9].n29 0.00771154
R18115 XThR.Tn[9].n25 XThR.Tn[9].n24 0.00771154
R18116 XThR.Tn[9].n20 XThR.Tn[9].n19 0.00771154
R18117 XThR.Tn[9].n15 XThR.Tn[9].n14 0.00771154
R18118 XA.Cn[5].n2 XA.Cn[5].n1 332.332
R18119 XA.Cn[5].n2 XA.Cn[5].n0 296.493
R18120 XA.Cn[5].n12 XA.Cn[5].n10 161.406
R18121 XA.Cn[5].n15 XA.Cn[5].n13 161.406
R18122 XA.Cn[5].n18 XA.Cn[5].n16 161.406
R18123 XA.Cn[5].n21 XA.Cn[5].n19 161.406
R18124 XA.Cn[5].n24 XA.Cn[5].n22 161.406
R18125 XA.Cn[5].n27 XA.Cn[5].n25 161.406
R18126 XA.Cn[5].n30 XA.Cn[5].n28 161.406
R18127 XA.Cn[5].n33 XA.Cn[5].n31 161.406
R18128 XA.Cn[5].n36 XA.Cn[5].n34 161.406
R18129 XA.Cn[5].n39 XA.Cn[5].n37 161.406
R18130 XA.Cn[5].n42 XA.Cn[5].n40 161.406
R18131 XA.Cn[5].n45 XA.Cn[5].n43 161.406
R18132 XA.Cn[5].n48 XA.Cn[5].n46 161.406
R18133 XA.Cn[5].n51 XA.Cn[5].n49 161.406
R18134 XA.Cn[5].n54 XA.Cn[5].n52 161.406
R18135 XA.Cn[5].n57 XA.Cn[5].n55 161.406
R18136 XA.Cn[5].n10 XA.Cn[5].t33 161.202
R18137 XA.Cn[5].n13 XA.Cn[5].t19 161.202
R18138 XA.Cn[5].n16 XA.Cn[5].t23 161.202
R18139 XA.Cn[5].n19 XA.Cn[5].t24 161.202
R18140 XA.Cn[5].n22 XA.Cn[5].t13 161.202
R18141 XA.Cn[5].n25 XA.Cn[5].t14 161.202
R18142 XA.Cn[5].n28 XA.Cn[5].t27 161.202
R18143 XA.Cn[5].n31 XA.Cn[5].t35 161.202
R18144 XA.Cn[5].n34 XA.Cn[5].t37 161.202
R18145 XA.Cn[5].n37 XA.Cn[5].t25 161.202
R18146 XA.Cn[5].n40 XA.Cn[5].t26 161.202
R18147 XA.Cn[5].n43 XA.Cn[5].t39 161.202
R18148 XA.Cn[5].n46 XA.Cn[5].t16 161.202
R18149 XA.Cn[5].n49 XA.Cn[5].t18 161.202
R18150 XA.Cn[5].n52 XA.Cn[5].t30 161.202
R18151 XA.Cn[5].n55 XA.Cn[5].t41 161.202
R18152 XA.Cn[5].n10 XA.Cn[5].t15 145.137
R18153 XA.Cn[5].n13 XA.Cn[5].t34 145.137
R18154 XA.Cn[5].n16 XA.Cn[5].t36 145.137
R18155 XA.Cn[5].n19 XA.Cn[5].t38 145.137
R18156 XA.Cn[5].n22 XA.Cn[5].t28 145.137
R18157 XA.Cn[5].n25 XA.Cn[5].t29 145.137
R18158 XA.Cn[5].n28 XA.Cn[5].t43 145.137
R18159 XA.Cn[5].n31 XA.Cn[5].t17 145.137
R18160 XA.Cn[5].n34 XA.Cn[5].t20 145.137
R18161 XA.Cn[5].n37 XA.Cn[5].t40 145.137
R18162 XA.Cn[5].n40 XA.Cn[5].t42 145.137
R18163 XA.Cn[5].n43 XA.Cn[5].t21 145.137
R18164 XA.Cn[5].n46 XA.Cn[5].t31 145.137
R18165 XA.Cn[5].n49 XA.Cn[5].t32 145.137
R18166 XA.Cn[5].n52 XA.Cn[5].t12 145.137
R18167 XA.Cn[5].n55 XA.Cn[5].t22 145.137
R18168 XA.Cn[5].n7 XA.Cn[5].n6 135.249
R18169 XA.Cn[5].n9 XA.Cn[5].n3 98.981
R18170 XA.Cn[5].n8 XA.Cn[5].n4 98.981
R18171 XA.Cn[5].n7 XA.Cn[5].n5 98.981
R18172 XA.Cn[5].n9 XA.Cn[5].n8 36.2672
R18173 XA.Cn[5].n8 XA.Cn[5].n7 36.2672
R18174 XA.Cn[5].n59 XA.Cn[5].n9 32.6405
R18175 XA.Cn[5].n1 XA.Cn[5].t5 26.5955
R18176 XA.Cn[5].n1 XA.Cn[5].t4 26.5955
R18177 XA.Cn[5].n0 XA.Cn[5].t7 26.5955
R18178 XA.Cn[5].n0 XA.Cn[5].t6 26.5955
R18179 XA.Cn[5].n3 XA.Cn[5].t9 24.9236
R18180 XA.Cn[5].n3 XA.Cn[5].t8 24.9236
R18181 XA.Cn[5].n4 XA.Cn[5].t11 24.9236
R18182 XA.Cn[5].n4 XA.Cn[5].t10 24.9236
R18183 XA.Cn[5].n5 XA.Cn[5].t2 24.9236
R18184 XA.Cn[5].n5 XA.Cn[5].t1 24.9236
R18185 XA.Cn[5].n6 XA.Cn[5].t0 24.9236
R18186 XA.Cn[5].n6 XA.Cn[5].t3 24.9236
R18187 XA.Cn[5] XA.Cn[5].n2 23.3605
R18188 XA.Cn[5] XA.Cn[5].n59 6.7205
R18189 XA.Cn[5].n58 XA.Cn[5] 3.62266
R18190 XA.Cn[5].n59 XA.Cn[5].n58 3.18437
R18191 XA.Cn[5].n15 XA.Cn[5] 0.931056
R18192 XA.Cn[5].n18 XA.Cn[5] 0.931056
R18193 XA.Cn[5].n21 XA.Cn[5] 0.931056
R18194 XA.Cn[5].n24 XA.Cn[5] 0.931056
R18195 XA.Cn[5].n27 XA.Cn[5] 0.931056
R18196 XA.Cn[5].n30 XA.Cn[5] 0.931056
R18197 XA.Cn[5].n33 XA.Cn[5] 0.931056
R18198 XA.Cn[5].n36 XA.Cn[5] 0.931056
R18199 XA.Cn[5].n39 XA.Cn[5] 0.931056
R18200 XA.Cn[5].n42 XA.Cn[5] 0.931056
R18201 XA.Cn[5].n45 XA.Cn[5] 0.931056
R18202 XA.Cn[5].n48 XA.Cn[5] 0.931056
R18203 XA.Cn[5].n51 XA.Cn[5] 0.931056
R18204 XA.Cn[5].n54 XA.Cn[5] 0.931056
R18205 XA.Cn[5].n57 XA.Cn[5] 0.931056
R18206 XA.Cn[5] XA.Cn[5].n12 0.396333
R18207 XA.Cn[5] XA.Cn[5].n15 0.396333
R18208 XA.Cn[5] XA.Cn[5].n18 0.396333
R18209 XA.Cn[5] XA.Cn[5].n21 0.396333
R18210 XA.Cn[5] XA.Cn[5].n24 0.396333
R18211 XA.Cn[5] XA.Cn[5].n27 0.396333
R18212 XA.Cn[5] XA.Cn[5].n30 0.396333
R18213 XA.Cn[5] XA.Cn[5].n33 0.396333
R18214 XA.Cn[5] XA.Cn[5].n36 0.396333
R18215 XA.Cn[5] XA.Cn[5].n39 0.396333
R18216 XA.Cn[5] XA.Cn[5].n42 0.396333
R18217 XA.Cn[5] XA.Cn[5].n45 0.396333
R18218 XA.Cn[5] XA.Cn[5].n48 0.396333
R18219 XA.Cn[5] XA.Cn[5].n51 0.396333
R18220 XA.Cn[5] XA.Cn[5].n54 0.396333
R18221 XA.Cn[5] XA.Cn[5].n57 0.396333
R18222 XA.Cn[5].n11 XA.Cn[5] 0.104667
R18223 XA.Cn[5].n14 XA.Cn[5] 0.104667
R18224 XA.Cn[5].n17 XA.Cn[5] 0.104667
R18225 XA.Cn[5].n20 XA.Cn[5] 0.104667
R18226 XA.Cn[5].n23 XA.Cn[5] 0.104667
R18227 XA.Cn[5].n26 XA.Cn[5] 0.104667
R18228 XA.Cn[5].n29 XA.Cn[5] 0.104667
R18229 XA.Cn[5].n32 XA.Cn[5] 0.104667
R18230 XA.Cn[5].n35 XA.Cn[5] 0.104667
R18231 XA.Cn[5].n38 XA.Cn[5] 0.104667
R18232 XA.Cn[5].n41 XA.Cn[5] 0.104667
R18233 XA.Cn[5].n44 XA.Cn[5] 0.104667
R18234 XA.Cn[5].n47 XA.Cn[5] 0.104667
R18235 XA.Cn[5].n50 XA.Cn[5] 0.104667
R18236 XA.Cn[5].n53 XA.Cn[5] 0.104667
R18237 XA.Cn[5].n56 XA.Cn[5] 0.104667
R18238 XA.Cn[5].n11 XA.Cn[5] 0.0309878
R18239 XA.Cn[5].n14 XA.Cn[5] 0.0309878
R18240 XA.Cn[5].n17 XA.Cn[5] 0.0309878
R18241 XA.Cn[5].n20 XA.Cn[5] 0.0309878
R18242 XA.Cn[5].n23 XA.Cn[5] 0.0309878
R18243 XA.Cn[5].n26 XA.Cn[5] 0.0309878
R18244 XA.Cn[5].n29 XA.Cn[5] 0.0309878
R18245 XA.Cn[5].n32 XA.Cn[5] 0.0309878
R18246 XA.Cn[5].n35 XA.Cn[5] 0.0309878
R18247 XA.Cn[5].n38 XA.Cn[5] 0.0309878
R18248 XA.Cn[5].n41 XA.Cn[5] 0.0309878
R18249 XA.Cn[5].n44 XA.Cn[5] 0.0309878
R18250 XA.Cn[5].n47 XA.Cn[5] 0.0309878
R18251 XA.Cn[5].n50 XA.Cn[5] 0.0309878
R18252 XA.Cn[5].n53 XA.Cn[5] 0.0309878
R18253 XA.Cn[5].n56 XA.Cn[5] 0.0309878
R18254 XA.Cn[5].n12 XA.Cn[5].n11 0.027939
R18255 XA.Cn[5].n15 XA.Cn[5].n14 0.027939
R18256 XA.Cn[5].n18 XA.Cn[5].n17 0.027939
R18257 XA.Cn[5].n21 XA.Cn[5].n20 0.027939
R18258 XA.Cn[5].n24 XA.Cn[5].n23 0.027939
R18259 XA.Cn[5].n27 XA.Cn[5].n26 0.027939
R18260 XA.Cn[5].n30 XA.Cn[5].n29 0.027939
R18261 XA.Cn[5].n33 XA.Cn[5].n32 0.027939
R18262 XA.Cn[5].n36 XA.Cn[5].n35 0.027939
R18263 XA.Cn[5].n39 XA.Cn[5].n38 0.027939
R18264 XA.Cn[5].n42 XA.Cn[5].n41 0.027939
R18265 XA.Cn[5].n45 XA.Cn[5].n44 0.027939
R18266 XA.Cn[5].n48 XA.Cn[5].n47 0.027939
R18267 XA.Cn[5].n51 XA.Cn[5].n50 0.027939
R18268 XA.Cn[5].n54 XA.Cn[5].n53 0.027939
R18269 XA.Cn[5].n57 XA.Cn[5].n56 0.027939
R18270 XA.Cn[5].n58 XA.Cn[5] 0.0129681
R18271 XA.Cn[9].n54 XA.Cn[9].n53 265.341
R18272 XA.Cn[9].n58 XA.Cn[9].n56 243.68
R18273 XA.Cn[9].n2 XA.Cn[9].n0 241.847
R18274 XA.Cn[9].n58 XA.Cn[9].n57 205.28
R18275 XA.Cn[9].n54 XA.Cn[9].n52 202.094
R18276 XA.Cn[9].n2 XA.Cn[9].n1 185
R18277 XA.Cn[9].n5 XA.Cn[9].n3 161.406
R18278 XA.Cn[9].n8 XA.Cn[9].n6 161.406
R18279 XA.Cn[9].n11 XA.Cn[9].n9 161.406
R18280 XA.Cn[9].n14 XA.Cn[9].n12 161.406
R18281 XA.Cn[9].n17 XA.Cn[9].n15 161.406
R18282 XA.Cn[9].n20 XA.Cn[9].n18 161.406
R18283 XA.Cn[9].n23 XA.Cn[9].n21 161.406
R18284 XA.Cn[9].n26 XA.Cn[9].n24 161.406
R18285 XA.Cn[9].n29 XA.Cn[9].n27 161.406
R18286 XA.Cn[9].n32 XA.Cn[9].n30 161.406
R18287 XA.Cn[9].n35 XA.Cn[9].n33 161.406
R18288 XA.Cn[9].n38 XA.Cn[9].n36 161.406
R18289 XA.Cn[9].n41 XA.Cn[9].n39 161.406
R18290 XA.Cn[9].n44 XA.Cn[9].n42 161.406
R18291 XA.Cn[9].n47 XA.Cn[9].n45 161.406
R18292 XA.Cn[9].n50 XA.Cn[9].n48 161.406
R18293 XA.Cn[9].n3 XA.Cn[9].t12 161.202
R18294 XA.Cn[9].n6 XA.Cn[9].t30 161.202
R18295 XA.Cn[9].n9 XA.Cn[9].t34 161.202
R18296 XA.Cn[9].n12 XA.Cn[9].t35 161.202
R18297 XA.Cn[9].n15 XA.Cn[9].t24 161.202
R18298 XA.Cn[9].n18 XA.Cn[9].t25 161.202
R18299 XA.Cn[9].n21 XA.Cn[9].t38 161.202
R18300 XA.Cn[9].n24 XA.Cn[9].t14 161.202
R18301 XA.Cn[9].n27 XA.Cn[9].t16 161.202
R18302 XA.Cn[9].n30 XA.Cn[9].t36 161.202
R18303 XA.Cn[9].n33 XA.Cn[9].t37 161.202
R18304 XA.Cn[9].n36 XA.Cn[9].t18 161.202
R18305 XA.Cn[9].n39 XA.Cn[9].t27 161.202
R18306 XA.Cn[9].n42 XA.Cn[9].t29 161.202
R18307 XA.Cn[9].n45 XA.Cn[9].t41 161.202
R18308 XA.Cn[9].n48 XA.Cn[9].t20 161.202
R18309 XA.Cn[9].n3 XA.Cn[9].t26 145.137
R18310 XA.Cn[9].n6 XA.Cn[9].t13 145.137
R18311 XA.Cn[9].n9 XA.Cn[9].t15 145.137
R18312 XA.Cn[9].n12 XA.Cn[9].t17 145.137
R18313 XA.Cn[9].n15 XA.Cn[9].t39 145.137
R18314 XA.Cn[9].n18 XA.Cn[9].t40 145.137
R18315 XA.Cn[9].n21 XA.Cn[9].t22 145.137
R18316 XA.Cn[9].n24 XA.Cn[9].t28 145.137
R18317 XA.Cn[9].n27 XA.Cn[9].t31 145.137
R18318 XA.Cn[9].n30 XA.Cn[9].t19 145.137
R18319 XA.Cn[9].n33 XA.Cn[9].t21 145.137
R18320 XA.Cn[9].n36 XA.Cn[9].t32 145.137
R18321 XA.Cn[9].n39 XA.Cn[9].t42 145.137
R18322 XA.Cn[9].n42 XA.Cn[9].t43 145.137
R18323 XA.Cn[9].n45 XA.Cn[9].t23 145.137
R18324 XA.Cn[9].n48 XA.Cn[9].t33 145.137
R18325 XA.Cn[9].n56 XA.Cn[9].t1 26.5955
R18326 XA.Cn[9].n56 XA.Cn[9].t0 26.5955
R18327 XA.Cn[9].n53 XA.Cn[9].t6 26.5955
R18328 XA.Cn[9].n53 XA.Cn[9].t5 26.5955
R18329 XA.Cn[9].n52 XA.Cn[9].t4 26.5955
R18330 XA.Cn[9].n52 XA.Cn[9].t7 26.5955
R18331 XA.Cn[9].n57 XA.Cn[9].t3 26.5955
R18332 XA.Cn[9].n57 XA.Cn[9].t2 26.5955
R18333 XA.Cn[9].n1 XA.Cn[9].t10 24.9236
R18334 XA.Cn[9].n1 XA.Cn[9].t11 24.9236
R18335 XA.Cn[9].n0 XA.Cn[9].t9 24.9236
R18336 XA.Cn[9].n0 XA.Cn[9].t8 24.9236
R18337 XA.Cn[9] XA.Cn[9].n58 22.9652
R18338 XA.Cn[9] XA.Cn[9].n2 18.8943
R18339 XA.Cn[9].n55 XA.Cn[9].n54 13.9299
R18340 XA.Cn[9] XA.Cn[9].n55 13.9299
R18341 XA.Cn[9].n51 XA.Cn[9] 6.34069
R18342 XA.Cn[9].n51 XA.Cn[9] 5.13485
R18343 XA.Cn[9] XA.Cn[9].n51 1.79489
R18344 XA.Cn[9].n55 XA.Cn[9] 1.19676
R18345 XA.Cn[9].n8 XA.Cn[9] 0.931056
R18346 XA.Cn[9].n11 XA.Cn[9] 0.931056
R18347 XA.Cn[9].n14 XA.Cn[9] 0.931056
R18348 XA.Cn[9].n17 XA.Cn[9] 0.931056
R18349 XA.Cn[9].n20 XA.Cn[9] 0.931056
R18350 XA.Cn[9].n23 XA.Cn[9] 0.931056
R18351 XA.Cn[9].n26 XA.Cn[9] 0.931056
R18352 XA.Cn[9].n29 XA.Cn[9] 0.931056
R18353 XA.Cn[9].n32 XA.Cn[9] 0.931056
R18354 XA.Cn[9].n35 XA.Cn[9] 0.931056
R18355 XA.Cn[9].n38 XA.Cn[9] 0.931056
R18356 XA.Cn[9].n41 XA.Cn[9] 0.931056
R18357 XA.Cn[9].n44 XA.Cn[9] 0.931056
R18358 XA.Cn[9].n47 XA.Cn[9] 0.931056
R18359 XA.Cn[9].n50 XA.Cn[9] 0.931056
R18360 XA.Cn[9] XA.Cn[9].n5 0.396333
R18361 XA.Cn[9] XA.Cn[9].n8 0.396333
R18362 XA.Cn[9] XA.Cn[9].n11 0.396333
R18363 XA.Cn[9] XA.Cn[9].n14 0.396333
R18364 XA.Cn[9] XA.Cn[9].n17 0.396333
R18365 XA.Cn[9] XA.Cn[9].n20 0.396333
R18366 XA.Cn[9] XA.Cn[9].n23 0.396333
R18367 XA.Cn[9] XA.Cn[9].n26 0.396333
R18368 XA.Cn[9] XA.Cn[9].n29 0.396333
R18369 XA.Cn[9] XA.Cn[9].n32 0.396333
R18370 XA.Cn[9] XA.Cn[9].n35 0.396333
R18371 XA.Cn[9] XA.Cn[9].n38 0.396333
R18372 XA.Cn[9] XA.Cn[9].n41 0.396333
R18373 XA.Cn[9] XA.Cn[9].n44 0.396333
R18374 XA.Cn[9] XA.Cn[9].n47 0.396333
R18375 XA.Cn[9] XA.Cn[9].n50 0.396333
R18376 XA.Cn[9].n4 XA.Cn[9] 0.104667
R18377 XA.Cn[9].n7 XA.Cn[9] 0.104667
R18378 XA.Cn[9].n10 XA.Cn[9] 0.104667
R18379 XA.Cn[9].n13 XA.Cn[9] 0.104667
R18380 XA.Cn[9].n16 XA.Cn[9] 0.104667
R18381 XA.Cn[9].n19 XA.Cn[9] 0.104667
R18382 XA.Cn[9].n22 XA.Cn[9] 0.104667
R18383 XA.Cn[9].n25 XA.Cn[9] 0.104667
R18384 XA.Cn[9].n28 XA.Cn[9] 0.104667
R18385 XA.Cn[9].n31 XA.Cn[9] 0.104667
R18386 XA.Cn[9].n34 XA.Cn[9] 0.104667
R18387 XA.Cn[9].n37 XA.Cn[9] 0.104667
R18388 XA.Cn[9].n40 XA.Cn[9] 0.104667
R18389 XA.Cn[9].n43 XA.Cn[9] 0.104667
R18390 XA.Cn[9].n46 XA.Cn[9] 0.104667
R18391 XA.Cn[9].n49 XA.Cn[9] 0.104667
R18392 XA.Cn[9].n4 XA.Cn[9] 0.0309878
R18393 XA.Cn[9].n7 XA.Cn[9] 0.0309878
R18394 XA.Cn[9].n10 XA.Cn[9] 0.0309878
R18395 XA.Cn[9].n13 XA.Cn[9] 0.0309878
R18396 XA.Cn[9].n16 XA.Cn[9] 0.0309878
R18397 XA.Cn[9].n19 XA.Cn[9] 0.0309878
R18398 XA.Cn[9].n22 XA.Cn[9] 0.0309878
R18399 XA.Cn[9].n25 XA.Cn[9] 0.0309878
R18400 XA.Cn[9].n28 XA.Cn[9] 0.0309878
R18401 XA.Cn[9].n31 XA.Cn[9] 0.0309878
R18402 XA.Cn[9].n34 XA.Cn[9] 0.0309878
R18403 XA.Cn[9].n37 XA.Cn[9] 0.0309878
R18404 XA.Cn[9].n40 XA.Cn[9] 0.0309878
R18405 XA.Cn[9].n43 XA.Cn[9] 0.0309878
R18406 XA.Cn[9].n46 XA.Cn[9] 0.0309878
R18407 XA.Cn[9].n49 XA.Cn[9] 0.0309878
R18408 XA.Cn[9].n5 XA.Cn[9].n4 0.027939
R18409 XA.Cn[9].n8 XA.Cn[9].n7 0.027939
R18410 XA.Cn[9].n11 XA.Cn[9].n10 0.027939
R18411 XA.Cn[9].n14 XA.Cn[9].n13 0.027939
R18412 XA.Cn[9].n17 XA.Cn[9].n16 0.027939
R18413 XA.Cn[9].n20 XA.Cn[9].n19 0.027939
R18414 XA.Cn[9].n23 XA.Cn[9].n22 0.027939
R18415 XA.Cn[9].n26 XA.Cn[9].n25 0.027939
R18416 XA.Cn[9].n29 XA.Cn[9].n28 0.027939
R18417 XA.Cn[9].n32 XA.Cn[9].n31 0.027939
R18418 XA.Cn[9].n35 XA.Cn[9].n34 0.027939
R18419 XA.Cn[9].n38 XA.Cn[9].n37 0.027939
R18420 XA.Cn[9].n41 XA.Cn[9].n40 0.027939
R18421 XA.Cn[9].n44 XA.Cn[9].n43 0.027939
R18422 XA.Cn[9].n47 XA.Cn[9].n46 0.027939
R18423 XA.Cn[9].n50 XA.Cn[9].n49 0.027939
R18424 XA.Cn[11].n2 XA.Cn[11].n1 265.341
R18425 XA.Cn[11].n5 XA.Cn[11].n3 243.68
R18426 XA.Cn[11].n58 XA.Cn[11].n56 241.847
R18427 XA.Cn[11].n5 XA.Cn[11].n4 205.28
R18428 XA.Cn[11].n2 XA.Cn[11].n0 202.094
R18429 XA.Cn[11].n58 XA.Cn[11].n57 185
R18430 XA.Cn[11].n9 XA.Cn[11].n7 161.406
R18431 XA.Cn[11].n12 XA.Cn[11].n10 161.406
R18432 XA.Cn[11].n15 XA.Cn[11].n13 161.406
R18433 XA.Cn[11].n18 XA.Cn[11].n16 161.406
R18434 XA.Cn[11].n21 XA.Cn[11].n19 161.406
R18435 XA.Cn[11].n24 XA.Cn[11].n22 161.406
R18436 XA.Cn[11].n27 XA.Cn[11].n25 161.406
R18437 XA.Cn[11].n30 XA.Cn[11].n28 161.406
R18438 XA.Cn[11].n33 XA.Cn[11].n31 161.406
R18439 XA.Cn[11].n36 XA.Cn[11].n34 161.406
R18440 XA.Cn[11].n39 XA.Cn[11].n37 161.406
R18441 XA.Cn[11].n42 XA.Cn[11].n40 161.406
R18442 XA.Cn[11].n45 XA.Cn[11].n43 161.406
R18443 XA.Cn[11].n48 XA.Cn[11].n46 161.406
R18444 XA.Cn[11].n51 XA.Cn[11].n49 161.406
R18445 XA.Cn[11].n54 XA.Cn[11].n52 161.406
R18446 XA.Cn[11].n7 XA.Cn[11].t18 161.202
R18447 XA.Cn[11].n10 XA.Cn[11].t35 161.202
R18448 XA.Cn[11].n13 XA.Cn[11].t37 161.202
R18449 XA.Cn[11].n16 XA.Cn[11].t39 161.202
R18450 XA.Cn[11].n19 XA.Cn[11].t28 161.202
R18451 XA.Cn[11].n22 XA.Cn[11].t29 161.202
R18452 XA.Cn[11].n25 XA.Cn[11].t42 161.202
R18453 XA.Cn[11].n28 XA.Cn[11].t19 161.202
R18454 XA.Cn[11].n31 XA.Cn[11].t21 161.202
R18455 XA.Cn[11].n34 XA.Cn[11].t40 161.202
R18456 XA.Cn[11].n37 XA.Cn[11].t41 161.202
R18457 XA.Cn[11].n40 XA.Cn[11].t22 161.202
R18458 XA.Cn[11].n43 XA.Cn[11].t30 161.202
R18459 XA.Cn[11].n46 XA.Cn[11].t33 161.202
R18460 XA.Cn[11].n49 XA.Cn[11].t14 161.202
R18461 XA.Cn[11].n52 XA.Cn[11].t24 161.202
R18462 XA.Cn[11].n7 XA.Cn[11].t20 145.137
R18463 XA.Cn[11].n10 XA.Cn[11].t38 145.137
R18464 XA.Cn[11].n13 XA.Cn[11].t43 145.137
R18465 XA.Cn[11].n16 XA.Cn[11].t12 145.137
R18466 XA.Cn[11].n19 XA.Cn[11].t31 145.137
R18467 XA.Cn[11].n22 XA.Cn[11].t32 145.137
R18468 XA.Cn[11].n25 XA.Cn[11].t16 145.137
R18469 XA.Cn[11].n28 XA.Cn[11].t23 145.137
R18470 XA.Cn[11].n31 XA.Cn[11].t25 145.137
R18471 XA.Cn[11].n34 XA.Cn[11].t13 145.137
R18472 XA.Cn[11].n37 XA.Cn[11].t15 145.137
R18473 XA.Cn[11].n40 XA.Cn[11].t26 145.137
R18474 XA.Cn[11].n43 XA.Cn[11].t34 145.137
R18475 XA.Cn[11].n46 XA.Cn[11].t36 145.137
R18476 XA.Cn[11].n49 XA.Cn[11].t17 145.137
R18477 XA.Cn[11].n52 XA.Cn[11].t27 145.137
R18478 XA.Cn[11].n1 XA.Cn[11].t1 26.5955
R18479 XA.Cn[11].n1 XA.Cn[11].t7 26.5955
R18480 XA.Cn[11].n0 XA.Cn[11].t11 26.5955
R18481 XA.Cn[11].n0 XA.Cn[11].t8 26.5955
R18482 XA.Cn[11].n3 XA.Cn[11].t2 26.5955
R18483 XA.Cn[11].n3 XA.Cn[11].t5 26.5955
R18484 XA.Cn[11].n4 XA.Cn[11].t4 26.5955
R18485 XA.Cn[11].n4 XA.Cn[11].t3 26.5955
R18486 XA.Cn[11].n56 XA.Cn[11].t6 24.9236
R18487 XA.Cn[11].n56 XA.Cn[11].t9 24.9236
R18488 XA.Cn[11].n57 XA.Cn[11].t0 24.9236
R18489 XA.Cn[11].n57 XA.Cn[11].t10 24.9236
R18490 XA.Cn[11] XA.Cn[11].n5 22.9652
R18491 XA.Cn[11] XA.Cn[11].n58 18.8943
R18492 XA.Cn[11].n6 XA.Cn[11].n2 13.9299
R18493 XA.Cn[11].n6 XA.Cn[11] 13.9299
R18494 XA.Cn[11] XA.Cn[11].n55 6.34069
R18495 XA.Cn[11].n55 XA.Cn[11] 5.13485
R18496 XA.Cn[11].n55 XA.Cn[11] 1.79489
R18497 XA.Cn[11] XA.Cn[11].n6 1.19676
R18498 XA.Cn[11].n12 XA.Cn[11] 0.931056
R18499 XA.Cn[11].n15 XA.Cn[11] 0.931056
R18500 XA.Cn[11].n18 XA.Cn[11] 0.931056
R18501 XA.Cn[11].n21 XA.Cn[11] 0.931056
R18502 XA.Cn[11].n24 XA.Cn[11] 0.931056
R18503 XA.Cn[11].n27 XA.Cn[11] 0.931056
R18504 XA.Cn[11].n30 XA.Cn[11] 0.931056
R18505 XA.Cn[11].n33 XA.Cn[11] 0.931056
R18506 XA.Cn[11].n36 XA.Cn[11] 0.931056
R18507 XA.Cn[11].n39 XA.Cn[11] 0.931056
R18508 XA.Cn[11].n42 XA.Cn[11] 0.931056
R18509 XA.Cn[11].n45 XA.Cn[11] 0.931056
R18510 XA.Cn[11].n48 XA.Cn[11] 0.931056
R18511 XA.Cn[11].n51 XA.Cn[11] 0.931056
R18512 XA.Cn[11].n54 XA.Cn[11] 0.931056
R18513 XA.Cn[11] XA.Cn[11].n9 0.396333
R18514 XA.Cn[11] XA.Cn[11].n12 0.396333
R18515 XA.Cn[11] XA.Cn[11].n15 0.396333
R18516 XA.Cn[11] XA.Cn[11].n18 0.396333
R18517 XA.Cn[11] XA.Cn[11].n21 0.396333
R18518 XA.Cn[11] XA.Cn[11].n24 0.396333
R18519 XA.Cn[11] XA.Cn[11].n27 0.396333
R18520 XA.Cn[11] XA.Cn[11].n30 0.396333
R18521 XA.Cn[11] XA.Cn[11].n33 0.396333
R18522 XA.Cn[11] XA.Cn[11].n36 0.396333
R18523 XA.Cn[11] XA.Cn[11].n39 0.396333
R18524 XA.Cn[11] XA.Cn[11].n42 0.396333
R18525 XA.Cn[11] XA.Cn[11].n45 0.396333
R18526 XA.Cn[11] XA.Cn[11].n48 0.396333
R18527 XA.Cn[11] XA.Cn[11].n51 0.396333
R18528 XA.Cn[11] XA.Cn[11].n54 0.396333
R18529 XA.Cn[11].n8 XA.Cn[11] 0.104667
R18530 XA.Cn[11].n11 XA.Cn[11] 0.104667
R18531 XA.Cn[11].n14 XA.Cn[11] 0.104667
R18532 XA.Cn[11].n17 XA.Cn[11] 0.104667
R18533 XA.Cn[11].n20 XA.Cn[11] 0.104667
R18534 XA.Cn[11].n23 XA.Cn[11] 0.104667
R18535 XA.Cn[11].n26 XA.Cn[11] 0.104667
R18536 XA.Cn[11].n29 XA.Cn[11] 0.104667
R18537 XA.Cn[11].n32 XA.Cn[11] 0.104667
R18538 XA.Cn[11].n35 XA.Cn[11] 0.104667
R18539 XA.Cn[11].n38 XA.Cn[11] 0.104667
R18540 XA.Cn[11].n41 XA.Cn[11] 0.104667
R18541 XA.Cn[11].n44 XA.Cn[11] 0.104667
R18542 XA.Cn[11].n47 XA.Cn[11] 0.104667
R18543 XA.Cn[11].n50 XA.Cn[11] 0.104667
R18544 XA.Cn[11].n53 XA.Cn[11] 0.104667
R18545 XA.Cn[11].n8 XA.Cn[11] 0.0309878
R18546 XA.Cn[11].n11 XA.Cn[11] 0.0309878
R18547 XA.Cn[11].n14 XA.Cn[11] 0.0309878
R18548 XA.Cn[11].n17 XA.Cn[11] 0.0309878
R18549 XA.Cn[11].n20 XA.Cn[11] 0.0309878
R18550 XA.Cn[11].n23 XA.Cn[11] 0.0309878
R18551 XA.Cn[11].n26 XA.Cn[11] 0.0309878
R18552 XA.Cn[11].n29 XA.Cn[11] 0.0309878
R18553 XA.Cn[11].n32 XA.Cn[11] 0.0309878
R18554 XA.Cn[11].n35 XA.Cn[11] 0.0309878
R18555 XA.Cn[11].n38 XA.Cn[11] 0.0309878
R18556 XA.Cn[11].n41 XA.Cn[11] 0.0309878
R18557 XA.Cn[11].n44 XA.Cn[11] 0.0309878
R18558 XA.Cn[11].n47 XA.Cn[11] 0.0309878
R18559 XA.Cn[11].n50 XA.Cn[11] 0.0309878
R18560 XA.Cn[11].n53 XA.Cn[11] 0.0309878
R18561 XA.Cn[11].n9 XA.Cn[11].n8 0.027939
R18562 XA.Cn[11].n12 XA.Cn[11].n11 0.027939
R18563 XA.Cn[11].n15 XA.Cn[11].n14 0.027939
R18564 XA.Cn[11].n18 XA.Cn[11].n17 0.027939
R18565 XA.Cn[11].n21 XA.Cn[11].n20 0.027939
R18566 XA.Cn[11].n24 XA.Cn[11].n23 0.027939
R18567 XA.Cn[11].n27 XA.Cn[11].n26 0.027939
R18568 XA.Cn[11].n30 XA.Cn[11].n29 0.027939
R18569 XA.Cn[11].n33 XA.Cn[11].n32 0.027939
R18570 XA.Cn[11].n36 XA.Cn[11].n35 0.027939
R18571 XA.Cn[11].n39 XA.Cn[11].n38 0.027939
R18572 XA.Cn[11].n42 XA.Cn[11].n41 0.027939
R18573 XA.Cn[11].n45 XA.Cn[11].n44 0.027939
R18574 XA.Cn[11].n48 XA.Cn[11].n47 0.027939
R18575 XA.Cn[11].n51 XA.Cn[11].n50 0.027939
R18576 XA.Cn[11].n54 XA.Cn[11].n53 0.027939
R18577 XA.Cn[12].n55 XA.Cn[12].n54 256.103
R18578 XA.Cn[12].n59 XA.Cn[12].n57 243.68
R18579 XA.Cn[12].n2 XA.Cn[12].n0 241.847
R18580 XA.Cn[12].n59 XA.Cn[12].n58 205.28
R18581 XA.Cn[12].n55 XA.Cn[12].n53 202.095
R18582 XA.Cn[12].n2 XA.Cn[12].n1 185
R18583 XA.Cn[12].n5 XA.Cn[12].n3 161.406
R18584 XA.Cn[12].n8 XA.Cn[12].n6 161.406
R18585 XA.Cn[12].n11 XA.Cn[12].n9 161.406
R18586 XA.Cn[12].n14 XA.Cn[12].n12 161.406
R18587 XA.Cn[12].n17 XA.Cn[12].n15 161.406
R18588 XA.Cn[12].n20 XA.Cn[12].n18 161.406
R18589 XA.Cn[12].n23 XA.Cn[12].n21 161.406
R18590 XA.Cn[12].n26 XA.Cn[12].n24 161.406
R18591 XA.Cn[12].n29 XA.Cn[12].n27 161.406
R18592 XA.Cn[12].n32 XA.Cn[12].n30 161.406
R18593 XA.Cn[12].n35 XA.Cn[12].n33 161.406
R18594 XA.Cn[12].n38 XA.Cn[12].n36 161.406
R18595 XA.Cn[12].n41 XA.Cn[12].n39 161.406
R18596 XA.Cn[12].n44 XA.Cn[12].n42 161.406
R18597 XA.Cn[12].n47 XA.Cn[12].n45 161.406
R18598 XA.Cn[12].n50 XA.Cn[12].n48 161.406
R18599 XA.Cn[12].n3 XA.Cn[12].t35 161.202
R18600 XA.Cn[12].n6 XA.Cn[12].t20 161.202
R18601 XA.Cn[12].n9 XA.Cn[12].t22 161.202
R18602 XA.Cn[12].n12 XA.Cn[12].t24 161.202
R18603 XA.Cn[12].n15 XA.Cn[12].t13 161.202
R18604 XA.Cn[12].n18 XA.Cn[12].t14 161.202
R18605 XA.Cn[12].n21 XA.Cn[12].t27 161.202
R18606 XA.Cn[12].n24 XA.Cn[12].t36 161.202
R18607 XA.Cn[12].n27 XA.Cn[12].t38 161.202
R18608 XA.Cn[12].n30 XA.Cn[12].t25 161.202
R18609 XA.Cn[12].n33 XA.Cn[12].t26 161.202
R18610 XA.Cn[12].n36 XA.Cn[12].t39 161.202
R18611 XA.Cn[12].n39 XA.Cn[12].t15 161.202
R18612 XA.Cn[12].n42 XA.Cn[12].t18 161.202
R18613 XA.Cn[12].n45 XA.Cn[12].t31 161.202
R18614 XA.Cn[12].n48 XA.Cn[12].t41 161.202
R18615 XA.Cn[12].n3 XA.Cn[12].t37 145.137
R18616 XA.Cn[12].n6 XA.Cn[12].t23 145.137
R18617 XA.Cn[12].n9 XA.Cn[12].t28 145.137
R18618 XA.Cn[12].n12 XA.Cn[12].t29 145.137
R18619 XA.Cn[12].n15 XA.Cn[12].t16 145.137
R18620 XA.Cn[12].n18 XA.Cn[12].t17 145.137
R18621 XA.Cn[12].n21 XA.Cn[12].t33 145.137
R18622 XA.Cn[12].n24 XA.Cn[12].t40 145.137
R18623 XA.Cn[12].n27 XA.Cn[12].t42 145.137
R18624 XA.Cn[12].n30 XA.Cn[12].t30 145.137
R18625 XA.Cn[12].n33 XA.Cn[12].t32 145.137
R18626 XA.Cn[12].n36 XA.Cn[12].t43 145.137
R18627 XA.Cn[12].n39 XA.Cn[12].t19 145.137
R18628 XA.Cn[12].n42 XA.Cn[12].t21 145.137
R18629 XA.Cn[12].n45 XA.Cn[12].t34 145.137
R18630 XA.Cn[12].n48 XA.Cn[12].t12 145.137
R18631 XA.Cn[12].n53 XA.Cn[12].t1 26.5955
R18632 XA.Cn[12].n53 XA.Cn[12].t2 26.5955
R18633 XA.Cn[12].n57 XA.Cn[12].t9 26.5955
R18634 XA.Cn[12].n57 XA.Cn[12].t8 26.5955
R18635 XA.Cn[12].n58 XA.Cn[12].t11 26.5955
R18636 XA.Cn[12].n58 XA.Cn[12].t10 26.5955
R18637 XA.Cn[12].n54 XA.Cn[12].t0 26.5955
R18638 XA.Cn[12].n54 XA.Cn[12].t3 26.5955
R18639 XA.Cn[12].n1 XA.Cn[12].t5 24.9236
R18640 XA.Cn[12].n1 XA.Cn[12].t4 24.9236
R18641 XA.Cn[12].n0 XA.Cn[12].t7 24.9236
R18642 XA.Cn[12].n0 XA.Cn[12].t6 24.9236
R18643 XA.Cn[12] XA.Cn[12].n59 22.9652
R18644 XA.Cn[12] XA.Cn[12].n2 22.9615
R18645 XA.Cn[12].n56 XA.Cn[12].n55 13.9299
R18646 XA.Cn[12] XA.Cn[12].n56 13.9299
R18647 XA.Cn[12].n52 XA.Cn[12].n51 5.13244
R18648 XA.Cn[12].n51 XA.Cn[12] 3.8444
R18649 XA.Cn[12].n56 XA.Cn[12].n52 2.99115
R18650 XA.Cn[12].n56 XA.Cn[12] 2.87153
R18651 XA.Cn[12].n52 XA.Cn[12] 2.2734
R18652 XA.Cn[12].n8 XA.Cn[12] 0.931056
R18653 XA.Cn[12].n11 XA.Cn[12] 0.931056
R18654 XA.Cn[12].n14 XA.Cn[12] 0.931056
R18655 XA.Cn[12].n17 XA.Cn[12] 0.931056
R18656 XA.Cn[12].n20 XA.Cn[12] 0.931056
R18657 XA.Cn[12].n23 XA.Cn[12] 0.931056
R18658 XA.Cn[12].n26 XA.Cn[12] 0.931056
R18659 XA.Cn[12].n29 XA.Cn[12] 0.931056
R18660 XA.Cn[12].n32 XA.Cn[12] 0.931056
R18661 XA.Cn[12].n35 XA.Cn[12] 0.931056
R18662 XA.Cn[12].n38 XA.Cn[12] 0.931056
R18663 XA.Cn[12].n41 XA.Cn[12] 0.931056
R18664 XA.Cn[12].n44 XA.Cn[12] 0.931056
R18665 XA.Cn[12].n47 XA.Cn[12] 0.931056
R18666 XA.Cn[12].n50 XA.Cn[12] 0.931056
R18667 XA.Cn[12] XA.Cn[12].n5 0.396333
R18668 XA.Cn[12] XA.Cn[12].n8 0.396333
R18669 XA.Cn[12] XA.Cn[12].n11 0.396333
R18670 XA.Cn[12] XA.Cn[12].n14 0.396333
R18671 XA.Cn[12] XA.Cn[12].n17 0.396333
R18672 XA.Cn[12] XA.Cn[12].n20 0.396333
R18673 XA.Cn[12] XA.Cn[12].n23 0.396333
R18674 XA.Cn[12] XA.Cn[12].n26 0.396333
R18675 XA.Cn[12] XA.Cn[12].n29 0.396333
R18676 XA.Cn[12] XA.Cn[12].n32 0.396333
R18677 XA.Cn[12] XA.Cn[12].n35 0.396333
R18678 XA.Cn[12] XA.Cn[12].n38 0.396333
R18679 XA.Cn[12] XA.Cn[12].n41 0.396333
R18680 XA.Cn[12] XA.Cn[12].n44 0.396333
R18681 XA.Cn[12] XA.Cn[12].n47 0.396333
R18682 XA.Cn[12] XA.Cn[12].n50 0.396333
R18683 XA.Cn[12].n4 XA.Cn[12] 0.104667
R18684 XA.Cn[12].n7 XA.Cn[12] 0.104667
R18685 XA.Cn[12].n10 XA.Cn[12] 0.104667
R18686 XA.Cn[12].n13 XA.Cn[12] 0.104667
R18687 XA.Cn[12].n16 XA.Cn[12] 0.104667
R18688 XA.Cn[12].n19 XA.Cn[12] 0.104667
R18689 XA.Cn[12].n22 XA.Cn[12] 0.104667
R18690 XA.Cn[12].n25 XA.Cn[12] 0.104667
R18691 XA.Cn[12].n28 XA.Cn[12] 0.104667
R18692 XA.Cn[12].n31 XA.Cn[12] 0.104667
R18693 XA.Cn[12].n34 XA.Cn[12] 0.104667
R18694 XA.Cn[12].n37 XA.Cn[12] 0.104667
R18695 XA.Cn[12].n40 XA.Cn[12] 0.104667
R18696 XA.Cn[12].n43 XA.Cn[12] 0.104667
R18697 XA.Cn[12].n46 XA.Cn[12] 0.104667
R18698 XA.Cn[12].n49 XA.Cn[12] 0.104667
R18699 XA.Cn[12].n4 XA.Cn[12] 0.0309878
R18700 XA.Cn[12].n7 XA.Cn[12] 0.0309878
R18701 XA.Cn[12].n10 XA.Cn[12] 0.0309878
R18702 XA.Cn[12].n13 XA.Cn[12] 0.0309878
R18703 XA.Cn[12].n16 XA.Cn[12] 0.0309878
R18704 XA.Cn[12].n19 XA.Cn[12] 0.0309878
R18705 XA.Cn[12].n22 XA.Cn[12] 0.0309878
R18706 XA.Cn[12].n25 XA.Cn[12] 0.0309878
R18707 XA.Cn[12].n28 XA.Cn[12] 0.0309878
R18708 XA.Cn[12].n31 XA.Cn[12] 0.0309878
R18709 XA.Cn[12].n34 XA.Cn[12] 0.0309878
R18710 XA.Cn[12].n37 XA.Cn[12] 0.0309878
R18711 XA.Cn[12].n40 XA.Cn[12] 0.0309878
R18712 XA.Cn[12].n43 XA.Cn[12] 0.0309878
R18713 XA.Cn[12].n46 XA.Cn[12] 0.0309878
R18714 XA.Cn[12].n49 XA.Cn[12] 0.0309878
R18715 XA.Cn[12].n5 XA.Cn[12].n4 0.027939
R18716 XA.Cn[12].n8 XA.Cn[12].n7 0.027939
R18717 XA.Cn[12].n11 XA.Cn[12].n10 0.027939
R18718 XA.Cn[12].n14 XA.Cn[12].n13 0.027939
R18719 XA.Cn[12].n17 XA.Cn[12].n16 0.027939
R18720 XA.Cn[12].n20 XA.Cn[12].n19 0.027939
R18721 XA.Cn[12].n23 XA.Cn[12].n22 0.027939
R18722 XA.Cn[12].n26 XA.Cn[12].n25 0.027939
R18723 XA.Cn[12].n29 XA.Cn[12].n28 0.027939
R18724 XA.Cn[12].n32 XA.Cn[12].n31 0.027939
R18725 XA.Cn[12].n35 XA.Cn[12].n34 0.027939
R18726 XA.Cn[12].n38 XA.Cn[12].n37 0.027939
R18727 XA.Cn[12].n41 XA.Cn[12].n40 0.027939
R18728 XA.Cn[12].n44 XA.Cn[12].n43 0.027939
R18729 XA.Cn[12].n47 XA.Cn[12].n46 0.027939
R18730 XA.Cn[12].n50 XA.Cn[12].n49 0.027939
R18731 XA.Cn[12].n51 XA.Cn[12] 0.00316553
R18732 XA.Cn[13].n55 XA.Cn[13].n54 265.341
R18733 XA.Cn[13].n59 XA.Cn[13].n57 243.68
R18734 XA.Cn[13].n2 XA.Cn[13].n0 241.847
R18735 XA.Cn[13].n59 XA.Cn[13].n58 205.28
R18736 XA.Cn[13].n55 XA.Cn[13].n53 202.094
R18737 XA.Cn[13].n2 XA.Cn[13].n1 185
R18738 XA.Cn[13].n5 XA.Cn[13].n3 161.406
R18739 XA.Cn[13].n8 XA.Cn[13].n6 161.406
R18740 XA.Cn[13].n11 XA.Cn[13].n9 161.406
R18741 XA.Cn[13].n14 XA.Cn[13].n12 161.406
R18742 XA.Cn[13].n17 XA.Cn[13].n15 161.406
R18743 XA.Cn[13].n20 XA.Cn[13].n18 161.406
R18744 XA.Cn[13].n23 XA.Cn[13].n21 161.406
R18745 XA.Cn[13].n26 XA.Cn[13].n24 161.406
R18746 XA.Cn[13].n29 XA.Cn[13].n27 161.406
R18747 XA.Cn[13].n32 XA.Cn[13].n30 161.406
R18748 XA.Cn[13].n35 XA.Cn[13].n33 161.406
R18749 XA.Cn[13].n38 XA.Cn[13].n36 161.406
R18750 XA.Cn[13].n41 XA.Cn[13].n39 161.406
R18751 XA.Cn[13].n44 XA.Cn[13].n42 161.406
R18752 XA.Cn[13].n47 XA.Cn[13].n45 161.406
R18753 XA.Cn[13].n50 XA.Cn[13].n48 161.406
R18754 XA.Cn[13].n3 XA.Cn[13].t27 161.202
R18755 XA.Cn[13].n6 XA.Cn[13].t12 161.202
R18756 XA.Cn[13].n9 XA.Cn[13].t14 161.202
R18757 XA.Cn[13].n12 XA.Cn[13].t16 161.202
R18758 XA.Cn[13].n15 XA.Cn[13].t37 161.202
R18759 XA.Cn[13].n18 XA.Cn[13].t38 161.202
R18760 XA.Cn[13].n21 XA.Cn[13].t19 161.202
R18761 XA.Cn[13].n24 XA.Cn[13].t28 161.202
R18762 XA.Cn[13].n27 XA.Cn[13].t30 161.202
R18763 XA.Cn[13].n30 XA.Cn[13].t17 161.202
R18764 XA.Cn[13].n33 XA.Cn[13].t18 161.202
R18765 XA.Cn[13].n36 XA.Cn[13].t31 161.202
R18766 XA.Cn[13].n39 XA.Cn[13].t39 161.202
R18767 XA.Cn[13].n42 XA.Cn[13].t42 161.202
R18768 XA.Cn[13].n45 XA.Cn[13].t23 161.202
R18769 XA.Cn[13].n48 XA.Cn[13].t33 161.202
R18770 XA.Cn[13].n3 XA.Cn[13].t29 145.137
R18771 XA.Cn[13].n6 XA.Cn[13].t15 145.137
R18772 XA.Cn[13].n9 XA.Cn[13].t20 145.137
R18773 XA.Cn[13].n12 XA.Cn[13].t21 145.137
R18774 XA.Cn[13].n15 XA.Cn[13].t40 145.137
R18775 XA.Cn[13].n18 XA.Cn[13].t41 145.137
R18776 XA.Cn[13].n21 XA.Cn[13].t25 145.137
R18777 XA.Cn[13].n24 XA.Cn[13].t32 145.137
R18778 XA.Cn[13].n27 XA.Cn[13].t34 145.137
R18779 XA.Cn[13].n30 XA.Cn[13].t22 145.137
R18780 XA.Cn[13].n33 XA.Cn[13].t24 145.137
R18781 XA.Cn[13].n36 XA.Cn[13].t35 145.137
R18782 XA.Cn[13].n39 XA.Cn[13].t43 145.137
R18783 XA.Cn[13].n42 XA.Cn[13].t13 145.137
R18784 XA.Cn[13].n45 XA.Cn[13].t26 145.137
R18785 XA.Cn[13].n48 XA.Cn[13].t36 145.137
R18786 XA.Cn[13].n53 XA.Cn[13].t2 26.5955
R18787 XA.Cn[13].n53 XA.Cn[13].t1 26.5955
R18788 XA.Cn[13].n57 XA.Cn[13].t9 26.5955
R18789 XA.Cn[13].n57 XA.Cn[13].t8 26.5955
R18790 XA.Cn[13].n58 XA.Cn[13].t11 26.5955
R18791 XA.Cn[13].n58 XA.Cn[13].t10 26.5955
R18792 XA.Cn[13].n54 XA.Cn[13].t0 26.5955
R18793 XA.Cn[13].n54 XA.Cn[13].t3 26.5955
R18794 XA.Cn[13].n1 XA.Cn[13].t4 24.9236
R18795 XA.Cn[13].n1 XA.Cn[13].t6 24.9236
R18796 XA.Cn[13].n0 XA.Cn[13].t7 24.9236
R18797 XA.Cn[13].n0 XA.Cn[13].t5 24.9236
R18798 XA.Cn[13] XA.Cn[13].n59 22.9652
R18799 XA.Cn[13] XA.Cn[13].n2 18.8943
R18800 XA.Cn[13].n56 XA.Cn[13].n55 13.9299
R18801 XA.Cn[13] XA.Cn[13].n56 13.9299
R18802 XA.Cn[13].n52 XA.Cn[13] 6.34069
R18803 XA.Cn[13].n52 XA.Cn[13].n51 5.13021
R18804 XA.Cn[13].n51 XA.Cn[13] 4.03795
R18805 XA.Cn[13] XA.Cn[13].n52 1.79489
R18806 XA.Cn[13].n56 XA.Cn[13] 1.19676
R18807 XA.Cn[13].n8 XA.Cn[13] 0.931056
R18808 XA.Cn[13].n11 XA.Cn[13] 0.931056
R18809 XA.Cn[13].n14 XA.Cn[13] 0.931056
R18810 XA.Cn[13].n17 XA.Cn[13] 0.931056
R18811 XA.Cn[13].n20 XA.Cn[13] 0.931056
R18812 XA.Cn[13].n23 XA.Cn[13] 0.931056
R18813 XA.Cn[13].n26 XA.Cn[13] 0.931056
R18814 XA.Cn[13].n29 XA.Cn[13] 0.931056
R18815 XA.Cn[13].n32 XA.Cn[13] 0.931056
R18816 XA.Cn[13].n35 XA.Cn[13] 0.931056
R18817 XA.Cn[13].n38 XA.Cn[13] 0.931056
R18818 XA.Cn[13].n41 XA.Cn[13] 0.931056
R18819 XA.Cn[13].n44 XA.Cn[13] 0.931056
R18820 XA.Cn[13].n47 XA.Cn[13] 0.931056
R18821 XA.Cn[13].n50 XA.Cn[13] 0.931056
R18822 XA.Cn[13] XA.Cn[13].n5 0.396333
R18823 XA.Cn[13] XA.Cn[13].n8 0.396333
R18824 XA.Cn[13] XA.Cn[13].n11 0.396333
R18825 XA.Cn[13] XA.Cn[13].n14 0.396333
R18826 XA.Cn[13] XA.Cn[13].n17 0.396333
R18827 XA.Cn[13] XA.Cn[13].n20 0.396333
R18828 XA.Cn[13] XA.Cn[13].n23 0.396333
R18829 XA.Cn[13] XA.Cn[13].n26 0.396333
R18830 XA.Cn[13] XA.Cn[13].n29 0.396333
R18831 XA.Cn[13] XA.Cn[13].n32 0.396333
R18832 XA.Cn[13] XA.Cn[13].n35 0.396333
R18833 XA.Cn[13] XA.Cn[13].n38 0.396333
R18834 XA.Cn[13] XA.Cn[13].n41 0.396333
R18835 XA.Cn[13] XA.Cn[13].n44 0.396333
R18836 XA.Cn[13] XA.Cn[13].n47 0.396333
R18837 XA.Cn[13] XA.Cn[13].n50 0.396333
R18838 XA.Cn[13].n4 XA.Cn[13] 0.104667
R18839 XA.Cn[13].n7 XA.Cn[13] 0.104667
R18840 XA.Cn[13].n10 XA.Cn[13] 0.104667
R18841 XA.Cn[13].n13 XA.Cn[13] 0.104667
R18842 XA.Cn[13].n16 XA.Cn[13] 0.104667
R18843 XA.Cn[13].n19 XA.Cn[13] 0.104667
R18844 XA.Cn[13].n22 XA.Cn[13] 0.104667
R18845 XA.Cn[13].n25 XA.Cn[13] 0.104667
R18846 XA.Cn[13].n28 XA.Cn[13] 0.104667
R18847 XA.Cn[13].n31 XA.Cn[13] 0.104667
R18848 XA.Cn[13].n34 XA.Cn[13] 0.104667
R18849 XA.Cn[13].n37 XA.Cn[13] 0.104667
R18850 XA.Cn[13].n40 XA.Cn[13] 0.104667
R18851 XA.Cn[13].n43 XA.Cn[13] 0.104667
R18852 XA.Cn[13].n46 XA.Cn[13] 0.104667
R18853 XA.Cn[13].n49 XA.Cn[13] 0.104667
R18854 XA.Cn[13].n4 XA.Cn[13] 0.0309878
R18855 XA.Cn[13].n7 XA.Cn[13] 0.0309878
R18856 XA.Cn[13].n10 XA.Cn[13] 0.0309878
R18857 XA.Cn[13].n13 XA.Cn[13] 0.0309878
R18858 XA.Cn[13].n16 XA.Cn[13] 0.0309878
R18859 XA.Cn[13].n19 XA.Cn[13] 0.0309878
R18860 XA.Cn[13].n22 XA.Cn[13] 0.0309878
R18861 XA.Cn[13].n25 XA.Cn[13] 0.0309878
R18862 XA.Cn[13].n28 XA.Cn[13] 0.0309878
R18863 XA.Cn[13].n31 XA.Cn[13] 0.0309878
R18864 XA.Cn[13].n34 XA.Cn[13] 0.0309878
R18865 XA.Cn[13].n37 XA.Cn[13] 0.0309878
R18866 XA.Cn[13].n40 XA.Cn[13] 0.0309878
R18867 XA.Cn[13].n43 XA.Cn[13] 0.0309878
R18868 XA.Cn[13].n46 XA.Cn[13] 0.0309878
R18869 XA.Cn[13].n49 XA.Cn[13] 0.0309878
R18870 XA.Cn[13].n5 XA.Cn[13].n4 0.027939
R18871 XA.Cn[13].n8 XA.Cn[13].n7 0.027939
R18872 XA.Cn[13].n11 XA.Cn[13].n10 0.027939
R18873 XA.Cn[13].n14 XA.Cn[13].n13 0.027939
R18874 XA.Cn[13].n17 XA.Cn[13].n16 0.027939
R18875 XA.Cn[13].n20 XA.Cn[13].n19 0.027939
R18876 XA.Cn[13].n23 XA.Cn[13].n22 0.027939
R18877 XA.Cn[13].n26 XA.Cn[13].n25 0.027939
R18878 XA.Cn[13].n29 XA.Cn[13].n28 0.027939
R18879 XA.Cn[13].n32 XA.Cn[13].n31 0.027939
R18880 XA.Cn[13].n35 XA.Cn[13].n34 0.027939
R18881 XA.Cn[13].n38 XA.Cn[13].n37 0.027939
R18882 XA.Cn[13].n41 XA.Cn[13].n40 0.027939
R18883 XA.Cn[13].n44 XA.Cn[13].n43 0.027939
R18884 XA.Cn[13].n47 XA.Cn[13].n46 0.027939
R18885 XA.Cn[13].n50 XA.Cn[13].n49 0.027939
R18886 XA.Cn[13].n51 XA.Cn[13] 0.00548355
R18887 XA.Cn[0].n2 XA.Cn[0].n1 332.332
R18888 XA.Cn[0].n2 XA.Cn[0].n0 296.493
R18889 XA.Cn[0].n12 XA.Cn[0].n10 161.406
R18890 XA.Cn[0].n15 XA.Cn[0].n13 161.406
R18891 XA.Cn[0].n18 XA.Cn[0].n16 161.406
R18892 XA.Cn[0].n21 XA.Cn[0].n19 161.406
R18893 XA.Cn[0].n24 XA.Cn[0].n22 161.406
R18894 XA.Cn[0].n27 XA.Cn[0].n25 161.406
R18895 XA.Cn[0].n30 XA.Cn[0].n28 161.406
R18896 XA.Cn[0].n33 XA.Cn[0].n31 161.406
R18897 XA.Cn[0].n36 XA.Cn[0].n34 161.406
R18898 XA.Cn[0].n39 XA.Cn[0].n37 161.406
R18899 XA.Cn[0].n42 XA.Cn[0].n40 161.406
R18900 XA.Cn[0].n45 XA.Cn[0].n43 161.406
R18901 XA.Cn[0].n48 XA.Cn[0].n46 161.406
R18902 XA.Cn[0].n51 XA.Cn[0].n49 161.406
R18903 XA.Cn[0].n54 XA.Cn[0].n52 161.406
R18904 XA.Cn[0].n57 XA.Cn[0].n55 161.406
R18905 XA.Cn[0].n10 XA.Cn[0].t22 161.202
R18906 XA.Cn[0].n13 XA.Cn[0].t41 161.202
R18907 XA.Cn[0].n16 XA.Cn[0].t12 161.202
R18908 XA.Cn[0].n19 XA.Cn[0].t13 161.202
R18909 XA.Cn[0].n22 XA.Cn[0].t32 161.202
R18910 XA.Cn[0].n25 XA.Cn[0].t34 161.202
R18911 XA.Cn[0].n28 XA.Cn[0].t17 161.202
R18912 XA.Cn[0].n31 XA.Cn[0].t25 161.202
R18913 XA.Cn[0].n34 XA.Cn[0].t26 161.202
R18914 XA.Cn[0].n37 XA.Cn[0].t15 161.202
R18915 XA.Cn[0].n40 XA.Cn[0].t16 161.202
R18916 XA.Cn[0].n43 XA.Cn[0].t27 161.202
R18917 XA.Cn[0].n46 XA.Cn[0].t36 161.202
R18918 XA.Cn[0].n49 XA.Cn[0].t38 161.202
R18919 XA.Cn[0].n52 XA.Cn[0].t19 161.202
R18920 XA.Cn[0].n55 XA.Cn[0].t29 161.202
R18921 XA.Cn[0].n10 XA.Cn[0].t18 145.137
R18922 XA.Cn[0].n13 XA.Cn[0].t35 145.137
R18923 XA.Cn[0].n16 XA.Cn[0].t37 145.137
R18924 XA.Cn[0].n19 XA.Cn[0].t39 145.137
R18925 XA.Cn[0].n22 XA.Cn[0].t28 145.137
R18926 XA.Cn[0].n25 XA.Cn[0].t30 145.137
R18927 XA.Cn[0].n28 XA.Cn[0].t43 145.137
R18928 XA.Cn[0].n31 XA.Cn[0].t20 145.137
R18929 XA.Cn[0].n34 XA.Cn[0].t21 145.137
R18930 XA.Cn[0].n37 XA.Cn[0].t40 145.137
R18931 XA.Cn[0].n40 XA.Cn[0].t42 145.137
R18932 XA.Cn[0].n43 XA.Cn[0].t23 145.137
R18933 XA.Cn[0].n46 XA.Cn[0].t31 145.137
R18934 XA.Cn[0].n49 XA.Cn[0].t33 145.137
R18935 XA.Cn[0].n52 XA.Cn[0].t14 145.137
R18936 XA.Cn[0].n55 XA.Cn[0].t24 145.137
R18937 XA.Cn[0].n7 XA.Cn[0].n6 135.248
R18938 XA.Cn[0].n9 XA.Cn[0].n3 98.982
R18939 XA.Cn[0].n8 XA.Cn[0].n4 98.982
R18940 XA.Cn[0].n7 XA.Cn[0].n5 98.982
R18941 XA.Cn[0].n9 XA.Cn[0].n8 36.2672
R18942 XA.Cn[0].n8 XA.Cn[0].n7 36.2672
R18943 XA.Cn[0].n59 XA.Cn[0].n9 32.6405
R18944 XA.Cn[0].n1 XA.Cn[0].t6 26.5955
R18945 XA.Cn[0].n1 XA.Cn[0].t5 26.5955
R18946 XA.Cn[0].n0 XA.Cn[0].t4 26.5955
R18947 XA.Cn[0].n0 XA.Cn[0].t3 26.5955
R18948 XA.Cn[0].n3 XA.Cn[0].t8 24.9236
R18949 XA.Cn[0].n3 XA.Cn[0].t7 24.9236
R18950 XA.Cn[0].n4 XA.Cn[0].t10 24.9236
R18951 XA.Cn[0].n4 XA.Cn[0].t9 24.9236
R18952 XA.Cn[0].n5 XA.Cn[0].t1 24.9236
R18953 XA.Cn[0].n5 XA.Cn[0].t11 24.9236
R18954 XA.Cn[0].n6 XA.Cn[0].t2 24.9236
R18955 XA.Cn[0].n6 XA.Cn[0].t0 24.9236
R18956 XA.Cn[0].n60 XA.Cn[0].n2 18.5605
R18957 XA.Cn[0].n60 XA.Cn[0].n59 11.5205
R18958 XA.Cn[0].n59 XA.Cn[0].n58 3.16389
R18959 XA.Cn[0].n15 XA.Cn[0] 0.931056
R18960 XA.Cn[0].n18 XA.Cn[0] 0.931056
R18961 XA.Cn[0].n21 XA.Cn[0] 0.931056
R18962 XA.Cn[0].n24 XA.Cn[0] 0.931056
R18963 XA.Cn[0].n27 XA.Cn[0] 0.931056
R18964 XA.Cn[0].n30 XA.Cn[0] 0.931056
R18965 XA.Cn[0].n33 XA.Cn[0] 0.931056
R18966 XA.Cn[0].n36 XA.Cn[0] 0.931056
R18967 XA.Cn[0].n39 XA.Cn[0] 0.931056
R18968 XA.Cn[0].n42 XA.Cn[0] 0.931056
R18969 XA.Cn[0].n45 XA.Cn[0] 0.931056
R18970 XA.Cn[0].n48 XA.Cn[0] 0.931056
R18971 XA.Cn[0].n51 XA.Cn[0] 0.931056
R18972 XA.Cn[0].n54 XA.Cn[0] 0.931056
R18973 XA.Cn[0].n57 XA.Cn[0] 0.931056
R18974 XA.Cn[0] XA.Cn[0].n60 0.6405
R18975 XA.Cn[0] XA.Cn[0].n12 0.396333
R18976 XA.Cn[0] XA.Cn[0].n15 0.396333
R18977 XA.Cn[0] XA.Cn[0].n18 0.396333
R18978 XA.Cn[0] XA.Cn[0].n21 0.396333
R18979 XA.Cn[0] XA.Cn[0].n24 0.396333
R18980 XA.Cn[0] XA.Cn[0].n27 0.396333
R18981 XA.Cn[0] XA.Cn[0].n30 0.396333
R18982 XA.Cn[0] XA.Cn[0].n33 0.396333
R18983 XA.Cn[0] XA.Cn[0].n36 0.396333
R18984 XA.Cn[0] XA.Cn[0].n39 0.396333
R18985 XA.Cn[0] XA.Cn[0].n42 0.396333
R18986 XA.Cn[0] XA.Cn[0].n45 0.396333
R18987 XA.Cn[0] XA.Cn[0].n48 0.396333
R18988 XA.Cn[0] XA.Cn[0].n51 0.396333
R18989 XA.Cn[0] XA.Cn[0].n54 0.396333
R18990 XA.Cn[0] XA.Cn[0].n57 0.396333
R18991 XA.Cn[0].n58 XA.Cn[0] 0.243556
R18992 XA.Cn[0].n11 XA.Cn[0] 0.104667
R18993 XA.Cn[0].n14 XA.Cn[0] 0.104667
R18994 XA.Cn[0].n17 XA.Cn[0] 0.104667
R18995 XA.Cn[0].n20 XA.Cn[0] 0.104667
R18996 XA.Cn[0].n23 XA.Cn[0] 0.104667
R18997 XA.Cn[0].n26 XA.Cn[0] 0.104667
R18998 XA.Cn[0].n29 XA.Cn[0] 0.104667
R18999 XA.Cn[0].n32 XA.Cn[0] 0.104667
R19000 XA.Cn[0].n35 XA.Cn[0] 0.104667
R19001 XA.Cn[0].n38 XA.Cn[0] 0.104667
R19002 XA.Cn[0].n41 XA.Cn[0] 0.104667
R19003 XA.Cn[0].n44 XA.Cn[0] 0.104667
R19004 XA.Cn[0].n47 XA.Cn[0] 0.104667
R19005 XA.Cn[0].n50 XA.Cn[0] 0.104667
R19006 XA.Cn[0].n53 XA.Cn[0] 0.104667
R19007 XA.Cn[0].n56 XA.Cn[0] 0.104667
R19008 XA.Cn[0].n58 XA.Cn[0] 0.0326429
R19009 XA.Cn[0].n11 XA.Cn[0] 0.0309878
R19010 XA.Cn[0].n14 XA.Cn[0] 0.0309878
R19011 XA.Cn[0].n17 XA.Cn[0] 0.0309878
R19012 XA.Cn[0].n20 XA.Cn[0] 0.0309878
R19013 XA.Cn[0].n23 XA.Cn[0] 0.0309878
R19014 XA.Cn[0].n26 XA.Cn[0] 0.0309878
R19015 XA.Cn[0].n29 XA.Cn[0] 0.0309878
R19016 XA.Cn[0].n32 XA.Cn[0] 0.0309878
R19017 XA.Cn[0].n35 XA.Cn[0] 0.0309878
R19018 XA.Cn[0].n38 XA.Cn[0] 0.0309878
R19019 XA.Cn[0].n41 XA.Cn[0] 0.0309878
R19020 XA.Cn[0].n44 XA.Cn[0] 0.0309878
R19021 XA.Cn[0].n47 XA.Cn[0] 0.0309878
R19022 XA.Cn[0].n50 XA.Cn[0] 0.0309878
R19023 XA.Cn[0].n53 XA.Cn[0] 0.0309878
R19024 XA.Cn[0].n56 XA.Cn[0] 0.0309878
R19025 XA.Cn[0].n12 XA.Cn[0].n11 0.027939
R19026 XA.Cn[0].n15 XA.Cn[0].n14 0.027939
R19027 XA.Cn[0].n18 XA.Cn[0].n17 0.027939
R19028 XA.Cn[0].n21 XA.Cn[0].n20 0.027939
R19029 XA.Cn[0].n24 XA.Cn[0].n23 0.027939
R19030 XA.Cn[0].n27 XA.Cn[0].n26 0.027939
R19031 XA.Cn[0].n30 XA.Cn[0].n29 0.027939
R19032 XA.Cn[0].n33 XA.Cn[0].n32 0.027939
R19033 XA.Cn[0].n36 XA.Cn[0].n35 0.027939
R19034 XA.Cn[0].n39 XA.Cn[0].n38 0.027939
R19035 XA.Cn[0].n42 XA.Cn[0].n41 0.027939
R19036 XA.Cn[0].n45 XA.Cn[0].n44 0.027939
R19037 XA.Cn[0].n48 XA.Cn[0].n47 0.027939
R19038 XA.Cn[0].n51 XA.Cn[0].n50 0.027939
R19039 XA.Cn[0].n54 XA.Cn[0].n53 0.027939
R19040 XA.Cn[0].n57 XA.Cn[0].n56 0.027939
R19041 thermo15c_0.XTB4.Y.n21 thermo15c_0.XTB4.Y.t0 235.56
R19042 thermo15c_0.XTB4.Y.n3 thermo15c_0.XTB4.Y.t3 212.081
R19043 thermo15c_0.XTB4.Y.n2 thermo15c_0.XTB4.Y.t2 212.081
R19044 thermo15c_0.XTB4.Y.n8 thermo15c_0.XTB4.Y.t17 212.081
R19045 thermo15c_0.XTB4.Y.n0 thermo15c_0.XTB4.Y.t13 212.081
R19046 thermo15c_0.XTB4.Y.n12 thermo15c_0.XTB4.Y.t8 212.081
R19047 thermo15c_0.XTB4.Y.n13 thermo15c_0.XTB4.Y.t12 212.081
R19048 thermo15c_0.XTB4.Y.n15 thermo15c_0.XTB4.Y.t6 212.081
R19049 thermo15c_0.XTB4.Y.n11 thermo15c_0.XTB4.Y.t16 212.081
R19050 thermo15c_0.XTB4.Y.n5 thermo15c_0.XTB4.Y.n4 173.761
R19051 thermo15c_0.XTB4.Y.n14 thermo15c_0.XTB4.Y 158.656
R19052 thermo15c_0.XTB4.Y.n7 thermo15c_0.XTB4.Y.n6 152
R19053 thermo15c_0.XTB4.Y.n5 thermo15c_0.XTB4.Y.n1 152
R19054 thermo15c_0.XTB4.Y.n10 thermo15c_0.XTB4.Y.n9 152
R19055 thermo15c_0.XTB4.Y.n17 thermo15c_0.XTB4.Y.n16 152
R19056 thermo15c_0.XTB4.Y.n3 thermo15c_0.XTB4.Y.t14 139.78
R19057 thermo15c_0.XTB4.Y.n2 thermo15c_0.XTB4.Y.t10 139.78
R19058 thermo15c_0.XTB4.Y.n8 thermo15c_0.XTB4.Y.t7 139.78
R19059 thermo15c_0.XTB4.Y.n0 thermo15c_0.XTB4.Y.t4 139.78
R19060 thermo15c_0.XTB4.Y.n12 thermo15c_0.XTB4.Y.t11 139.78
R19061 thermo15c_0.XTB4.Y.n13 thermo15c_0.XTB4.Y.t15 139.78
R19062 thermo15c_0.XTB4.Y.n15 thermo15c_0.XTB4.Y.t9 139.78
R19063 thermo15c_0.XTB4.Y.n11 thermo15c_0.XTB4.Y.t5 139.78
R19064 thermo15c_0.XTB4.Y.n20 thermo15c_0.XTB4.Y.t1 133.386
R19065 thermo15c_0.XTB4.Y.n19 thermo15c_0.XTB4.Y.n10 72.9296
R19066 thermo15c_0.XTB4.Y.n13 thermo15c_0.XTB4.Y.n12 61.346
R19067 thermo15c_0.XTB4.Y.n7 thermo15c_0.XTB4.Y.n1 49.6611
R19068 thermo15c_0.XTB4.Y.n9 thermo15c_0.XTB4.Y.n8 45.2793
R19069 thermo15c_0.XTB4.Y.n4 thermo15c_0.XTB4.Y.n2 42.3581
R19070 thermo15c_0.XTB4.Y.n19 thermo15c_0.XTB4.Y.n18 38.1854
R19071 thermo15c_0.XTB4.Y.n16 thermo15c_0.XTB4.Y.n11 30.6732
R19072 thermo15c_0.XTB4.Y.n16 thermo15c_0.XTB4.Y.n15 30.6732
R19073 thermo15c_0.XTB4.Y.n15 thermo15c_0.XTB4.Y.n14 30.6732
R19074 thermo15c_0.XTB4.Y.n14 thermo15c_0.XTB4.Y.n13 30.6732
R19075 thermo15c_0.XTB4.Y.n6 thermo15c_0.XTB4.Y.n5 21.7605
R19076 thermo15c_0.XTB4.Y thermo15c_0.XTB4.Y.n20 19.5051
R19077 thermo15c_0.XTB4.Y.n4 thermo15c_0.XTB4.Y.n3 18.9884
R19078 thermo15c_0.XTB4.Y.n9 thermo15c_0.XTB4.Y.n0 16.0672
R19079 thermo15c_0.XTB4.Y.n17 thermo15c_0.XTB4.Y 14.7905
R19080 thermo15c_0.XTB4.Y.n20 thermo15c_0.XTB4.Y.n19 11.994
R19081 thermo15c_0.XTB4.Y.n10 thermo15c_0.XTB4.Y 11.5205
R19082 thermo15c_0.XTB4.Y.n6 thermo15c_0.XTB4.Y 10.2405
R19083 thermo15c_0.XTB4.Y.n2 thermo15c_0.XTB4.Y.n1 7.30353
R19084 thermo15c_0.XTB4.Y.n18 thermo15c_0.XTB4.Y.n17 7.24578
R19085 thermo15c_0.XTB4.Y.n8 thermo15c_0.XTB4.Y.n7 4.38232
R19086 thermo15c_0.XTB4.Y.n21 thermo15c_0.XTB4.Y 2.22659
R19087 thermo15c_0.XTB4.Y thermo15c_0.XTB4.Y.n21 1.55202
R19088 thermo15c_0.XTB4.Y.n18 thermo15c_0.XTB4.Y 0.966538
R19089 XThR.Tn[3].n2 XThR.Tn[3].n1 332.332
R19090 XThR.Tn[3].n2 XThR.Tn[3].n0 296.493
R19091 XThR.Tn[3] XThR.Tn[3].n82 161.363
R19092 XThR.Tn[3] XThR.Tn[3].n77 161.363
R19093 XThR.Tn[3] XThR.Tn[3].n72 161.363
R19094 XThR.Tn[3] XThR.Tn[3].n67 161.363
R19095 XThR.Tn[3] XThR.Tn[3].n62 161.363
R19096 XThR.Tn[3] XThR.Tn[3].n57 161.363
R19097 XThR.Tn[3] XThR.Tn[3].n52 161.363
R19098 XThR.Tn[3] XThR.Tn[3].n47 161.363
R19099 XThR.Tn[3] XThR.Tn[3].n42 161.363
R19100 XThR.Tn[3] XThR.Tn[3].n37 161.363
R19101 XThR.Tn[3] XThR.Tn[3].n32 161.363
R19102 XThR.Tn[3] XThR.Tn[3].n27 161.363
R19103 XThR.Tn[3] XThR.Tn[3].n22 161.363
R19104 XThR.Tn[3] XThR.Tn[3].n17 161.363
R19105 XThR.Tn[3] XThR.Tn[3].n12 161.363
R19106 XThR.Tn[3] XThR.Tn[3].n10 161.363
R19107 XThR.Tn[3].n84 XThR.Tn[3].n83 161.3
R19108 XThR.Tn[3].n79 XThR.Tn[3].n78 161.3
R19109 XThR.Tn[3].n74 XThR.Tn[3].n73 161.3
R19110 XThR.Tn[3].n69 XThR.Tn[3].n68 161.3
R19111 XThR.Tn[3].n64 XThR.Tn[3].n63 161.3
R19112 XThR.Tn[3].n59 XThR.Tn[3].n58 161.3
R19113 XThR.Tn[3].n54 XThR.Tn[3].n53 161.3
R19114 XThR.Tn[3].n49 XThR.Tn[3].n48 161.3
R19115 XThR.Tn[3].n44 XThR.Tn[3].n43 161.3
R19116 XThR.Tn[3].n39 XThR.Tn[3].n38 161.3
R19117 XThR.Tn[3].n34 XThR.Tn[3].n33 161.3
R19118 XThR.Tn[3].n29 XThR.Tn[3].n28 161.3
R19119 XThR.Tn[3].n24 XThR.Tn[3].n23 161.3
R19120 XThR.Tn[3].n19 XThR.Tn[3].n18 161.3
R19121 XThR.Tn[3].n14 XThR.Tn[3].n13 161.3
R19122 XThR.Tn[3].n82 XThR.Tn[3].t46 161.106
R19123 XThR.Tn[3].n77 XThR.Tn[3].t53 161.106
R19124 XThR.Tn[3].n72 XThR.Tn[3].t34 161.106
R19125 XThR.Tn[3].n67 XThR.Tn[3].t17 161.106
R19126 XThR.Tn[3].n62 XThR.Tn[3].t44 161.106
R19127 XThR.Tn[3].n57 XThR.Tn[3].t69 161.106
R19128 XThR.Tn[3].n52 XThR.Tn[3].t51 161.106
R19129 XThR.Tn[3].n47 XThR.Tn[3].t31 161.106
R19130 XThR.Tn[3].n42 XThR.Tn[3].t14 161.106
R19131 XThR.Tn[3].n37 XThR.Tn[3].t20 161.106
R19132 XThR.Tn[3].n32 XThR.Tn[3].t68 161.106
R19133 XThR.Tn[3].n27 XThR.Tn[3].t33 161.106
R19134 XThR.Tn[3].n22 XThR.Tn[3].t67 161.106
R19135 XThR.Tn[3].n17 XThR.Tn[3].t49 161.106
R19136 XThR.Tn[3].n12 XThR.Tn[3].t70 161.106
R19137 XThR.Tn[3].n10 XThR.Tn[3].t57 161.106
R19138 XThR.Tn[3].n83 XThR.Tn[3].t27 159.978
R19139 XThR.Tn[3].n78 XThR.Tn[3].t32 159.978
R19140 XThR.Tn[3].n73 XThR.Tn[3].t15 159.978
R19141 XThR.Tn[3].n68 XThR.Tn[3].t63 159.978
R19142 XThR.Tn[3].n63 XThR.Tn[3].t25 159.978
R19143 XThR.Tn[3].n58 XThR.Tn[3].t50 159.978
R19144 XThR.Tn[3].n53 XThR.Tn[3].t30 159.978
R19145 XThR.Tn[3].n48 XThR.Tn[3].t73 159.978
R19146 XThR.Tn[3].n43 XThR.Tn[3].t61 159.978
R19147 XThR.Tn[3].n38 XThR.Tn[3].t66 159.978
R19148 XThR.Tn[3].n33 XThR.Tn[3].t48 159.978
R19149 XThR.Tn[3].n28 XThR.Tn[3].t13 159.978
R19150 XThR.Tn[3].n23 XThR.Tn[3].t47 159.978
R19151 XThR.Tn[3].n18 XThR.Tn[3].t29 159.978
R19152 XThR.Tn[3].n13 XThR.Tn[3].t55 159.978
R19153 XThR.Tn[3].n82 XThR.Tn[3].t36 145.038
R19154 XThR.Tn[3].n77 XThR.Tn[3].t60 145.038
R19155 XThR.Tn[3].n72 XThR.Tn[3].t40 145.038
R19156 XThR.Tn[3].n67 XThR.Tn[3].t21 145.038
R19157 XThR.Tn[3].n62 XThR.Tn[3].t54 145.038
R19158 XThR.Tn[3].n57 XThR.Tn[3].t35 145.038
R19159 XThR.Tn[3].n52 XThR.Tn[3].t41 145.038
R19160 XThR.Tn[3].n47 XThR.Tn[3].t22 145.038
R19161 XThR.Tn[3].n42 XThR.Tn[3].t19 145.038
R19162 XThR.Tn[3].n37 XThR.Tn[3].t52 145.038
R19163 XThR.Tn[3].n32 XThR.Tn[3].t72 145.038
R19164 XThR.Tn[3].n27 XThR.Tn[3].t39 145.038
R19165 XThR.Tn[3].n22 XThR.Tn[3].t71 145.038
R19166 XThR.Tn[3].n17 XThR.Tn[3].t59 145.038
R19167 XThR.Tn[3].n12 XThR.Tn[3].t18 145.038
R19168 XThR.Tn[3].n10 XThR.Tn[3].t64 145.038
R19169 XThR.Tn[3].n83 XThR.Tn[3].t38 143.911
R19170 XThR.Tn[3].n78 XThR.Tn[3].t65 143.911
R19171 XThR.Tn[3].n73 XThR.Tn[3].t43 143.911
R19172 XThR.Tn[3].n68 XThR.Tn[3].t26 143.911
R19173 XThR.Tn[3].n63 XThR.Tn[3].t58 143.911
R19174 XThR.Tn[3].n58 XThR.Tn[3].t37 143.911
R19175 XThR.Tn[3].n53 XThR.Tn[3].t45 143.911
R19176 XThR.Tn[3].n48 XThR.Tn[3].t28 143.911
R19177 XThR.Tn[3].n43 XThR.Tn[3].t23 143.911
R19178 XThR.Tn[3].n38 XThR.Tn[3].t56 143.911
R19179 XThR.Tn[3].n33 XThR.Tn[3].t16 143.911
R19180 XThR.Tn[3].n28 XThR.Tn[3].t42 143.911
R19181 XThR.Tn[3].n23 XThR.Tn[3].t12 143.911
R19182 XThR.Tn[3].n18 XThR.Tn[3].t62 143.911
R19183 XThR.Tn[3].n13 XThR.Tn[3].t24 143.911
R19184 XThR.Tn[3].n7 XThR.Tn[3].n6 135.249
R19185 XThR.Tn[3].n9 XThR.Tn[3].n3 98.981
R19186 XThR.Tn[3].n8 XThR.Tn[3].n4 98.981
R19187 XThR.Tn[3].n7 XThR.Tn[3].n5 98.981
R19188 XThR.Tn[3].n9 XThR.Tn[3].n8 36.2672
R19189 XThR.Tn[3].n8 XThR.Tn[3].n7 36.2672
R19190 XThR.Tn[3].n88 XThR.Tn[3].n9 32.6405
R19191 XThR.Tn[3].n1 XThR.Tn[3].t4 26.5955
R19192 XThR.Tn[3].n1 XThR.Tn[3].t7 26.5955
R19193 XThR.Tn[3].n0 XThR.Tn[3].t5 26.5955
R19194 XThR.Tn[3].n0 XThR.Tn[3].t6 26.5955
R19195 XThR.Tn[3].n3 XThR.Tn[3].t11 24.9236
R19196 XThR.Tn[3].n3 XThR.Tn[3].t8 24.9236
R19197 XThR.Tn[3].n4 XThR.Tn[3].t10 24.9236
R19198 XThR.Tn[3].n4 XThR.Tn[3].t9 24.9236
R19199 XThR.Tn[3].n5 XThR.Tn[3].t3 24.9236
R19200 XThR.Tn[3].n5 XThR.Tn[3].t1 24.9236
R19201 XThR.Tn[3].n6 XThR.Tn[3].t0 24.9236
R19202 XThR.Tn[3].n6 XThR.Tn[3].t2 24.9236
R19203 XThR.Tn[3].n89 XThR.Tn[3].n2 18.5605
R19204 XThR.Tn[3].n89 XThR.Tn[3].n88 11.5205
R19205 XThR.Tn[3].n88 XThR.Tn[3] 6.21508
R19206 XThR.Tn[3] XThR.Tn[3].n11 5.34038
R19207 XThR.Tn[3].n16 XThR.Tn[3].n15 4.5005
R19208 XThR.Tn[3].n21 XThR.Tn[3].n20 4.5005
R19209 XThR.Tn[3].n26 XThR.Tn[3].n25 4.5005
R19210 XThR.Tn[3].n31 XThR.Tn[3].n30 4.5005
R19211 XThR.Tn[3].n36 XThR.Tn[3].n35 4.5005
R19212 XThR.Tn[3].n41 XThR.Tn[3].n40 4.5005
R19213 XThR.Tn[3].n46 XThR.Tn[3].n45 4.5005
R19214 XThR.Tn[3].n51 XThR.Tn[3].n50 4.5005
R19215 XThR.Tn[3].n56 XThR.Tn[3].n55 4.5005
R19216 XThR.Tn[3].n61 XThR.Tn[3].n60 4.5005
R19217 XThR.Tn[3].n66 XThR.Tn[3].n65 4.5005
R19218 XThR.Tn[3].n71 XThR.Tn[3].n70 4.5005
R19219 XThR.Tn[3].n76 XThR.Tn[3].n75 4.5005
R19220 XThR.Tn[3].n81 XThR.Tn[3].n80 4.5005
R19221 XThR.Tn[3].n86 XThR.Tn[3].n85 4.5005
R19222 XThR.Tn[3].n87 XThR.Tn[3] 3.70586
R19223 XThR.Tn[3].n16 XThR.Tn[3] 2.52282
R19224 XThR.Tn[3].n21 XThR.Tn[3] 2.52282
R19225 XThR.Tn[3].n26 XThR.Tn[3] 2.52282
R19226 XThR.Tn[3].n31 XThR.Tn[3] 2.52282
R19227 XThR.Tn[3].n36 XThR.Tn[3] 2.52282
R19228 XThR.Tn[3].n41 XThR.Tn[3] 2.52282
R19229 XThR.Tn[3].n46 XThR.Tn[3] 2.52282
R19230 XThR.Tn[3].n51 XThR.Tn[3] 2.52282
R19231 XThR.Tn[3].n56 XThR.Tn[3] 2.52282
R19232 XThR.Tn[3].n61 XThR.Tn[3] 2.52282
R19233 XThR.Tn[3].n66 XThR.Tn[3] 2.52282
R19234 XThR.Tn[3].n71 XThR.Tn[3] 2.52282
R19235 XThR.Tn[3].n76 XThR.Tn[3] 2.52282
R19236 XThR.Tn[3].n81 XThR.Tn[3] 2.52282
R19237 XThR.Tn[3].n86 XThR.Tn[3] 2.52282
R19238 XThR.Tn[3].n84 XThR.Tn[3] 1.08677
R19239 XThR.Tn[3].n79 XThR.Tn[3] 1.08677
R19240 XThR.Tn[3].n74 XThR.Tn[3] 1.08677
R19241 XThR.Tn[3].n69 XThR.Tn[3] 1.08677
R19242 XThR.Tn[3].n64 XThR.Tn[3] 1.08677
R19243 XThR.Tn[3].n59 XThR.Tn[3] 1.08677
R19244 XThR.Tn[3].n54 XThR.Tn[3] 1.08677
R19245 XThR.Tn[3].n49 XThR.Tn[3] 1.08677
R19246 XThR.Tn[3].n44 XThR.Tn[3] 1.08677
R19247 XThR.Tn[3].n39 XThR.Tn[3] 1.08677
R19248 XThR.Tn[3].n34 XThR.Tn[3] 1.08677
R19249 XThR.Tn[3].n29 XThR.Tn[3] 1.08677
R19250 XThR.Tn[3].n24 XThR.Tn[3] 1.08677
R19251 XThR.Tn[3].n19 XThR.Tn[3] 1.08677
R19252 XThR.Tn[3].n14 XThR.Tn[3] 1.08677
R19253 XThR.Tn[3] XThR.Tn[3].n16 0.839786
R19254 XThR.Tn[3] XThR.Tn[3].n21 0.839786
R19255 XThR.Tn[3] XThR.Tn[3].n26 0.839786
R19256 XThR.Tn[3] XThR.Tn[3].n31 0.839786
R19257 XThR.Tn[3] XThR.Tn[3].n36 0.839786
R19258 XThR.Tn[3] XThR.Tn[3].n41 0.839786
R19259 XThR.Tn[3] XThR.Tn[3].n46 0.839786
R19260 XThR.Tn[3] XThR.Tn[3].n51 0.839786
R19261 XThR.Tn[3] XThR.Tn[3].n56 0.839786
R19262 XThR.Tn[3] XThR.Tn[3].n61 0.839786
R19263 XThR.Tn[3] XThR.Tn[3].n66 0.839786
R19264 XThR.Tn[3] XThR.Tn[3].n71 0.839786
R19265 XThR.Tn[3] XThR.Tn[3].n76 0.839786
R19266 XThR.Tn[3] XThR.Tn[3].n81 0.839786
R19267 XThR.Tn[3] XThR.Tn[3].n86 0.839786
R19268 XThR.Tn[3] XThR.Tn[3].n89 0.6405
R19269 XThR.Tn[3].n11 XThR.Tn[3] 0.499542
R19270 XThR.Tn[3].n85 XThR.Tn[3] 0.063
R19271 XThR.Tn[3].n80 XThR.Tn[3] 0.063
R19272 XThR.Tn[3].n75 XThR.Tn[3] 0.063
R19273 XThR.Tn[3].n70 XThR.Tn[3] 0.063
R19274 XThR.Tn[3].n65 XThR.Tn[3] 0.063
R19275 XThR.Tn[3].n60 XThR.Tn[3] 0.063
R19276 XThR.Tn[3].n55 XThR.Tn[3] 0.063
R19277 XThR.Tn[3].n50 XThR.Tn[3] 0.063
R19278 XThR.Tn[3].n45 XThR.Tn[3] 0.063
R19279 XThR.Tn[3].n40 XThR.Tn[3] 0.063
R19280 XThR.Tn[3].n35 XThR.Tn[3] 0.063
R19281 XThR.Tn[3].n30 XThR.Tn[3] 0.063
R19282 XThR.Tn[3].n25 XThR.Tn[3] 0.063
R19283 XThR.Tn[3].n20 XThR.Tn[3] 0.063
R19284 XThR.Tn[3].n15 XThR.Tn[3] 0.063
R19285 XThR.Tn[3].n87 XThR.Tn[3] 0.0540714
R19286 XThR.Tn[3] XThR.Tn[3].n87 0.038
R19287 XThR.Tn[3].n11 XThR.Tn[3] 0.0143889
R19288 XThR.Tn[3].n85 XThR.Tn[3].n84 0.00771154
R19289 XThR.Tn[3].n80 XThR.Tn[3].n79 0.00771154
R19290 XThR.Tn[3].n75 XThR.Tn[3].n74 0.00771154
R19291 XThR.Tn[3].n70 XThR.Tn[3].n69 0.00771154
R19292 XThR.Tn[3].n65 XThR.Tn[3].n64 0.00771154
R19293 XThR.Tn[3].n60 XThR.Tn[3].n59 0.00771154
R19294 XThR.Tn[3].n55 XThR.Tn[3].n54 0.00771154
R19295 XThR.Tn[3].n50 XThR.Tn[3].n49 0.00771154
R19296 XThR.Tn[3].n45 XThR.Tn[3].n44 0.00771154
R19297 XThR.Tn[3].n40 XThR.Tn[3].n39 0.00771154
R19298 XThR.Tn[3].n35 XThR.Tn[3].n34 0.00771154
R19299 XThR.Tn[3].n30 XThR.Tn[3].n29 0.00771154
R19300 XThR.Tn[3].n25 XThR.Tn[3].n24 0.00771154
R19301 XThR.Tn[3].n20 XThR.Tn[3].n19 0.00771154
R19302 XThR.Tn[3].n15 XThR.Tn[3].n14 0.00771154
R19303 XThR.Tn[5].n2 XThR.Tn[5].n1 332.332
R19304 XThR.Tn[5].n2 XThR.Tn[5].n0 296.493
R19305 XThR.Tn[5] XThR.Tn[5].n82 161.363
R19306 XThR.Tn[5] XThR.Tn[5].n77 161.363
R19307 XThR.Tn[5] XThR.Tn[5].n72 161.363
R19308 XThR.Tn[5] XThR.Tn[5].n67 161.363
R19309 XThR.Tn[5] XThR.Tn[5].n62 161.363
R19310 XThR.Tn[5] XThR.Tn[5].n57 161.363
R19311 XThR.Tn[5] XThR.Tn[5].n52 161.363
R19312 XThR.Tn[5] XThR.Tn[5].n47 161.363
R19313 XThR.Tn[5] XThR.Tn[5].n42 161.363
R19314 XThR.Tn[5] XThR.Tn[5].n37 161.363
R19315 XThR.Tn[5] XThR.Tn[5].n32 161.363
R19316 XThR.Tn[5] XThR.Tn[5].n27 161.363
R19317 XThR.Tn[5] XThR.Tn[5].n22 161.363
R19318 XThR.Tn[5] XThR.Tn[5].n17 161.363
R19319 XThR.Tn[5] XThR.Tn[5].n12 161.363
R19320 XThR.Tn[5] XThR.Tn[5].n10 161.363
R19321 XThR.Tn[5].n84 XThR.Tn[5].n83 161.3
R19322 XThR.Tn[5].n79 XThR.Tn[5].n78 161.3
R19323 XThR.Tn[5].n74 XThR.Tn[5].n73 161.3
R19324 XThR.Tn[5].n69 XThR.Tn[5].n68 161.3
R19325 XThR.Tn[5].n64 XThR.Tn[5].n63 161.3
R19326 XThR.Tn[5].n59 XThR.Tn[5].n58 161.3
R19327 XThR.Tn[5].n54 XThR.Tn[5].n53 161.3
R19328 XThR.Tn[5].n49 XThR.Tn[5].n48 161.3
R19329 XThR.Tn[5].n44 XThR.Tn[5].n43 161.3
R19330 XThR.Tn[5].n39 XThR.Tn[5].n38 161.3
R19331 XThR.Tn[5].n34 XThR.Tn[5].n33 161.3
R19332 XThR.Tn[5].n29 XThR.Tn[5].n28 161.3
R19333 XThR.Tn[5].n24 XThR.Tn[5].n23 161.3
R19334 XThR.Tn[5].n19 XThR.Tn[5].n18 161.3
R19335 XThR.Tn[5].n14 XThR.Tn[5].n13 161.3
R19336 XThR.Tn[5].n82 XThR.Tn[5].t62 161.106
R19337 XThR.Tn[5].n77 XThR.Tn[5].t70 161.106
R19338 XThR.Tn[5].n72 XThR.Tn[5].t52 161.106
R19339 XThR.Tn[5].n67 XThR.Tn[5].t35 161.106
R19340 XThR.Tn[5].n62 XThR.Tn[5].t60 161.106
R19341 XThR.Tn[5].n57 XThR.Tn[5].t24 161.106
R19342 XThR.Tn[5].n52 XThR.Tn[5].t68 161.106
R19343 XThR.Tn[5].n47 XThR.Tn[5].t49 161.106
R19344 XThR.Tn[5].n42 XThR.Tn[5].t32 161.106
R19345 XThR.Tn[5].n37 XThR.Tn[5].t40 161.106
R19346 XThR.Tn[5].n32 XThR.Tn[5].t22 161.106
R19347 XThR.Tn[5].n27 XThR.Tn[5].t51 161.106
R19348 XThR.Tn[5].n22 XThR.Tn[5].t21 161.106
R19349 XThR.Tn[5].n17 XThR.Tn[5].t66 161.106
R19350 XThR.Tn[5].n12 XThR.Tn[5].t26 161.106
R19351 XThR.Tn[5].n10 XThR.Tn[5].t72 161.106
R19352 XThR.Tn[5].n83 XThR.Tn[5].t59 159.978
R19353 XThR.Tn[5].n78 XThR.Tn[5].t64 159.978
R19354 XThR.Tn[5].n73 XThR.Tn[5].t47 159.978
R19355 XThR.Tn[5].n68 XThR.Tn[5].t31 159.978
R19356 XThR.Tn[5].n63 XThR.Tn[5].t57 159.978
R19357 XThR.Tn[5].n58 XThR.Tn[5].t20 159.978
R19358 XThR.Tn[5].n53 XThR.Tn[5].t63 159.978
R19359 XThR.Tn[5].n48 XThR.Tn[5].t45 159.978
R19360 XThR.Tn[5].n43 XThR.Tn[5].t29 159.978
R19361 XThR.Tn[5].n38 XThR.Tn[5].t37 159.978
R19362 XThR.Tn[5].n33 XThR.Tn[5].t19 159.978
R19363 XThR.Tn[5].n28 XThR.Tn[5].t46 159.978
R19364 XThR.Tn[5].n23 XThR.Tn[5].t18 159.978
R19365 XThR.Tn[5].n18 XThR.Tn[5].t61 159.978
R19366 XThR.Tn[5].n13 XThR.Tn[5].t23 159.978
R19367 XThR.Tn[5].n82 XThR.Tn[5].t54 145.038
R19368 XThR.Tn[5].n77 XThR.Tn[5].t12 145.038
R19369 XThR.Tn[5].n72 XThR.Tn[5].t56 145.038
R19370 XThR.Tn[5].n67 XThR.Tn[5].t41 145.038
R19371 XThR.Tn[5].n62 XThR.Tn[5].t71 145.038
R19372 XThR.Tn[5].n57 XThR.Tn[5].t53 145.038
R19373 XThR.Tn[5].n52 XThR.Tn[5].t58 145.038
R19374 XThR.Tn[5].n47 XThR.Tn[5].t42 145.038
R19375 XThR.Tn[5].n42 XThR.Tn[5].t38 145.038
R19376 XThR.Tn[5].n37 XThR.Tn[5].t69 145.038
R19377 XThR.Tn[5].n32 XThR.Tn[5].t30 145.038
R19378 XThR.Tn[5].n27 XThR.Tn[5].t55 145.038
R19379 XThR.Tn[5].n22 XThR.Tn[5].t28 145.038
R19380 XThR.Tn[5].n17 XThR.Tn[5].t73 145.038
R19381 XThR.Tn[5].n12 XThR.Tn[5].t39 145.038
R19382 XThR.Tn[5].n10 XThR.Tn[5].t17 145.038
R19383 XThR.Tn[5].n83 XThR.Tn[5].t27 143.911
R19384 XThR.Tn[5].n78 XThR.Tn[5].t50 143.911
R19385 XThR.Tn[5].n73 XThR.Tn[5].t34 143.911
R19386 XThR.Tn[5].n68 XThR.Tn[5].t15 143.911
R19387 XThR.Tn[5].n63 XThR.Tn[5].t44 143.911
R19388 XThR.Tn[5].n58 XThR.Tn[5].t25 143.911
R19389 XThR.Tn[5].n53 XThR.Tn[5].t36 143.911
R19390 XThR.Tn[5].n48 XThR.Tn[5].t16 143.911
R19391 XThR.Tn[5].n43 XThR.Tn[5].t14 143.911
R19392 XThR.Tn[5].n38 XThR.Tn[5].t43 143.911
R19393 XThR.Tn[5].n33 XThR.Tn[5].t67 143.911
R19394 XThR.Tn[5].n28 XThR.Tn[5].t33 143.911
R19395 XThR.Tn[5].n23 XThR.Tn[5].t65 143.911
R19396 XThR.Tn[5].n18 XThR.Tn[5].t48 143.911
R19397 XThR.Tn[5].n13 XThR.Tn[5].t13 143.911
R19398 XThR.Tn[5].n7 XThR.Tn[5].n5 135.249
R19399 XThR.Tn[5].n9 XThR.Tn[5].n3 98.981
R19400 XThR.Tn[5].n8 XThR.Tn[5].n4 98.981
R19401 XThR.Tn[5].n7 XThR.Tn[5].n6 98.981
R19402 XThR.Tn[5].n9 XThR.Tn[5].n8 36.2672
R19403 XThR.Tn[5].n8 XThR.Tn[5].n7 36.2672
R19404 XThR.Tn[5].n88 XThR.Tn[5].n9 32.6405
R19405 XThR.Tn[5].n1 XThR.Tn[5].t5 26.5955
R19406 XThR.Tn[5].n1 XThR.Tn[5].t4 26.5955
R19407 XThR.Tn[5].n0 XThR.Tn[5].t6 26.5955
R19408 XThR.Tn[5].n0 XThR.Tn[5].t7 26.5955
R19409 XThR.Tn[5].n3 XThR.Tn[5].t11 24.9236
R19410 XThR.Tn[5].n3 XThR.Tn[5].t8 24.9236
R19411 XThR.Tn[5].n4 XThR.Tn[5].t10 24.9236
R19412 XThR.Tn[5].n4 XThR.Tn[5].t9 24.9236
R19413 XThR.Tn[5].n5 XThR.Tn[5].t0 24.9236
R19414 XThR.Tn[5].n5 XThR.Tn[5].t1 24.9236
R19415 XThR.Tn[5].n6 XThR.Tn[5].t3 24.9236
R19416 XThR.Tn[5].n6 XThR.Tn[5].t2 24.9236
R19417 XThR.Tn[5].n89 XThR.Tn[5].n2 18.5605
R19418 XThR.Tn[5].n89 XThR.Tn[5].n88 11.5205
R19419 XThR.Tn[5].n88 XThR.Tn[5] 5.71508
R19420 XThR.Tn[5] XThR.Tn[5].n11 5.34038
R19421 XThR.Tn[5].n16 XThR.Tn[5].n15 4.5005
R19422 XThR.Tn[5].n21 XThR.Tn[5].n20 4.5005
R19423 XThR.Tn[5].n26 XThR.Tn[5].n25 4.5005
R19424 XThR.Tn[5].n31 XThR.Tn[5].n30 4.5005
R19425 XThR.Tn[5].n36 XThR.Tn[5].n35 4.5005
R19426 XThR.Tn[5].n41 XThR.Tn[5].n40 4.5005
R19427 XThR.Tn[5].n46 XThR.Tn[5].n45 4.5005
R19428 XThR.Tn[5].n51 XThR.Tn[5].n50 4.5005
R19429 XThR.Tn[5].n56 XThR.Tn[5].n55 4.5005
R19430 XThR.Tn[5].n61 XThR.Tn[5].n60 4.5005
R19431 XThR.Tn[5].n66 XThR.Tn[5].n65 4.5005
R19432 XThR.Tn[5].n71 XThR.Tn[5].n70 4.5005
R19433 XThR.Tn[5].n76 XThR.Tn[5].n75 4.5005
R19434 XThR.Tn[5].n81 XThR.Tn[5].n80 4.5005
R19435 XThR.Tn[5].n86 XThR.Tn[5].n85 4.5005
R19436 XThR.Tn[5].n87 XThR.Tn[5] 3.70586
R19437 XThR.Tn[5].n16 XThR.Tn[5] 2.52282
R19438 XThR.Tn[5].n21 XThR.Tn[5] 2.52282
R19439 XThR.Tn[5].n26 XThR.Tn[5] 2.52282
R19440 XThR.Tn[5].n31 XThR.Tn[5] 2.52282
R19441 XThR.Tn[5].n36 XThR.Tn[5] 2.52282
R19442 XThR.Tn[5].n41 XThR.Tn[5] 2.52282
R19443 XThR.Tn[5].n46 XThR.Tn[5] 2.52282
R19444 XThR.Tn[5].n51 XThR.Tn[5] 2.52282
R19445 XThR.Tn[5].n56 XThR.Tn[5] 2.52282
R19446 XThR.Tn[5].n61 XThR.Tn[5] 2.52282
R19447 XThR.Tn[5].n66 XThR.Tn[5] 2.52282
R19448 XThR.Tn[5].n71 XThR.Tn[5] 2.52282
R19449 XThR.Tn[5].n76 XThR.Tn[5] 2.52282
R19450 XThR.Tn[5].n81 XThR.Tn[5] 2.52282
R19451 XThR.Tn[5].n86 XThR.Tn[5] 2.52282
R19452 XThR.Tn[5].n84 XThR.Tn[5] 1.08677
R19453 XThR.Tn[5].n79 XThR.Tn[5] 1.08677
R19454 XThR.Tn[5].n74 XThR.Tn[5] 1.08677
R19455 XThR.Tn[5].n69 XThR.Tn[5] 1.08677
R19456 XThR.Tn[5].n64 XThR.Tn[5] 1.08677
R19457 XThR.Tn[5].n59 XThR.Tn[5] 1.08677
R19458 XThR.Tn[5].n54 XThR.Tn[5] 1.08677
R19459 XThR.Tn[5].n49 XThR.Tn[5] 1.08677
R19460 XThR.Tn[5].n44 XThR.Tn[5] 1.08677
R19461 XThR.Tn[5].n39 XThR.Tn[5] 1.08677
R19462 XThR.Tn[5].n34 XThR.Tn[5] 1.08677
R19463 XThR.Tn[5].n29 XThR.Tn[5] 1.08677
R19464 XThR.Tn[5].n24 XThR.Tn[5] 1.08677
R19465 XThR.Tn[5].n19 XThR.Tn[5] 1.08677
R19466 XThR.Tn[5].n14 XThR.Tn[5] 1.08677
R19467 XThR.Tn[5] XThR.Tn[5].n16 0.839786
R19468 XThR.Tn[5] XThR.Tn[5].n21 0.839786
R19469 XThR.Tn[5] XThR.Tn[5].n26 0.839786
R19470 XThR.Tn[5] XThR.Tn[5].n31 0.839786
R19471 XThR.Tn[5] XThR.Tn[5].n36 0.839786
R19472 XThR.Tn[5] XThR.Tn[5].n41 0.839786
R19473 XThR.Tn[5] XThR.Tn[5].n46 0.839786
R19474 XThR.Tn[5] XThR.Tn[5].n51 0.839786
R19475 XThR.Tn[5] XThR.Tn[5].n56 0.839786
R19476 XThR.Tn[5] XThR.Tn[5].n61 0.839786
R19477 XThR.Tn[5] XThR.Tn[5].n66 0.839786
R19478 XThR.Tn[5] XThR.Tn[5].n71 0.839786
R19479 XThR.Tn[5] XThR.Tn[5].n76 0.839786
R19480 XThR.Tn[5] XThR.Tn[5].n81 0.839786
R19481 XThR.Tn[5] XThR.Tn[5].n86 0.839786
R19482 XThR.Tn[5] XThR.Tn[5].n89 0.6405
R19483 XThR.Tn[5].n11 XThR.Tn[5] 0.499542
R19484 XThR.Tn[5].n85 XThR.Tn[5] 0.063
R19485 XThR.Tn[5].n80 XThR.Tn[5] 0.063
R19486 XThR.Tn[5].n75 XThR.Tn[5] 0.063
R19487 XThR.Tn[5].n70 XThR.Tn[5] 0.063
R19488 XThR.Tn[5].n65 XThR.Tn[5] 0.063
R19489 XThR.Tn[5].n60 XThR.Tn[5] 0.063
R19490 XThR.Tn[5].n55 XThR.Tn[5] 0.063
R19491 XThR.Tn[5].n50 XThR.Tn[5] 0.063
R19492 XThR.Tn[5].n45 XThR.Tn[5] 0.063
R19493 XThR.Tn[5].n40 XThR.Tn[5] 0.063
R19494 XThR.Tn[5].n35 XThR.Tn[5] 0.063
R19495 XThR.Tn[5].n30 XThR.Tn[5] 0.063
R19496 XThR.Tn[5].n25 XThR.Tn[5] 0.063
R19497 XThR.Tn[5].n20 XThR.Tn[5] 0.063
R19498 XThR.Tn[5].n15 XThR.Tn[5] 0.063
R19499 XThR.Tn[5].n87 XThR.Tn[5] 0.0540714
R19500 XThR.Tn[5] XThR.Tn[5].n87 0.038
R19501 XThR.Tn[5].n11 XThR.Tn[5] 0.0143889
R19502 XThR.Tn[5].n85 XThR.Tn[5].n84 0.00771154
R19503 XThR.Tn[5].n80 XThR.Tn[5].n79 0.00771154
R19504 XThR.Tn[5].n75 XThR.Tn[5].n74 0.00771154
R19505 XThR.Tn[5].n70 XThR.Tn[5].n69 0.00771154
R19506 XThR.Tn[5].n65 XThR.Tn[5].n64 0.00771154
R19507 XThR.Tn[5].n60 XThR.Tn[5].n59 0.00771154
R19508 XThR.Tn[5].n55 XThR.Tn[5].n54 0.00771154
R19509 XThR.Tn[5].n50 XThR.Tn[5].n49 0.00771154
R19510 XThR.Tn[5].n45 XThR.Tn[5].n44 0.00771154
R19511 XThR.Tn[5].n40 XThR.Tn[5].n39 0.00771154
R19512 XThR.Tn[5].n35 XThR.Tn[5].n34 0.00771154
R19513 XThR.Tn[5].n30 XThR.Tn[5].n29 0.00771154
R19514 XThR.Tn[5].n25 XThR.Tn[5].n24 0.00771154
R19515 XThR.Tn[5].n20 XThR.Tn[5].n19 0.00771154
R19516 XThR.Tn[5].n15 XThR.Tn[5].n14 0.00771154
R19517 XA.Cn[4].n2 XA.Cn[4].n1 332.332
R19518 XA.Cn[4].n2 XA.Cn[4].n0 296.493
R19519 XA.Cn[4].n12 XA.Cn[4].n10 161.406
R19520 XA.Cn[4].n15 XA.Cn[4].n13 161.406
R19521 XA.Cn[4].n18 XA.Cn[4].n16 161.406
R19522 XA.Cn[4].n21 XA.Cn[4].n19 161.406
R19523 XA.Cn[4].n24 XA.Cn[4].n22 161.406
R19524 XA.Cn[4].n27 XA.Cn[4].n25 161.406
R19525 XA.Cn[4].n30 XA.Cn[4].n28 161.406
R19526 XA.Cn[4].n33 XA.Cn[4].n31 161.406
R19527 XA.Cn[4].n36 XA.Cn[4].n34 161.406
R19528 XA.Cn[4].n39 XA.Cn[4].n37 161.406
R19529 XA.Cn[4].n42 XA.Cn[4].n40 161.406
R19530 XA.Cn[4].n45 XA.Cn[4].n43 161.406
R19531 XA.Cn[4].n48 XA.Cn[4].n46 161.406
R19532 XA.Cn[4].n51 XA.Cn[4].n49 161.406
R19533 XA.Cn[4].n54 XA.Cn[4].n52 161.406
R19534 XA.Cn[4].n57 XA.Cn[4].n55 161.406
R19535 XA.Cn[4].n10 XA.Cn[4].t26 161.202
R19536 XA.Cn[4].n13 XA.Cn[4].t43 161.202
R19537 XA.Cn[4].n16 XA.Cn[4].t13 161.202
R19538 XA.Cn[4].n19 XA.Cn[4].t15 161.202
R19539 XA.Cn[4].n22 XA.Cn[4].t36 161.202
R19540 XA.Cn[4].n25 XA.Cn[4].t37 161.202
R19541 XA.Cn[4].n28 XA.Cn[4].t18 161.202
R19542 XA.Cn[4].n31 XA.Cn[4].t27 161.202
R19543 XA.Cn[4].n34 XA.Cn[4].t29 161.202
R19544 XA.Cn[4].n37 XA.Cn[4].t16 161.202
R19545 XA.Cn[4].n40 XA.Cn[4].t17 161.202
R19546 XA.Cn[4].n43 XA.Cn[4].t30 161.202
R19547 XA.Cn[4].n46 XA.Cn[4].t38 161.202
R19548 XA.Cn[4].n49 XA.Cn[4].t41 161.202
R19549 XA.Cn[4].n52 XA.Cn[4].t22 161.202
R19550 XA.Cn[4].n55 XA.Cn[4].t32 161.202
R19551 XA.Cn[4].n10 XA.Cn[4].t28 145.137
R19552 XA.Cn[4].n13 XA.Cn[4].t14 145.137
R19553 XA.Cn[4].n16 XA.Cn[4].t19 145.137
R19554 XA.Cn[4].n19 XA.Cn[4].t20 145.137
R19555 XA.Cn[4].n22 XA.Cn[4].t39 145.137
R19556 XA.Cn[4].n25 XA.Cn[4].t40 145.137
R19557 XA.Cn[4].n28 XA.Cn[4].t24 145.137
R19558 XA.Cn[4].n31 XA.Cn[4].t31 145.137
R19559 XA.Cn[4].n34 XA.Cn[4].t33 145.137
R19560 XA.Cn[4].n37 XA.Cn[4].t21 145.137
R19561 XA.Cn[4].n40 XA.Cn[4].t23 145.137
R19562 XA.Cn[4].n43 XA.Cn[4].t34 145.137
R19563 XA.Cn[4].n46 XA.Cn[4].t42 145.137
R19564 XA.Cn[4].n49 XA.Cn[4].t12 145.137
R19565 XA.Cn[4].n52 XA.Cn[4].t25 145.137
R19566 XA.Cn[4].n55 XA.Cn[4].t35 145.137
R19567 XA.Cn[4].n7 XA.Cn[4].n6 135.248
R19568 XA.Cn[4].n9 XA.Cn[4].n3 98.982
R19569 XA.Cn[4].n8 XA.Cn[4].n4 98.982
R19570 XA.Cn[4].n7 XA.Cn[4].n5 98.982
R19571 XA.Cn[4].n9 XA.Cn[4].n8 36.2672
R19572 XA.Cn[4].n8 XA.Cn[4].n7 36.2672
R19573 XA.Cn[4].n59 XA.Cn[4].n9 32.6405
R19574 XA.Cn[4].n1 XA.Cn[4].t7 26.5955
R19575 XA.Cn[4].n1 XA.Cn[4].t6 26.5955
R19576 XA.Cn[4].n0 XA.Cn[4].t5 26.5955
R19577 XA.Cn[4].n0 XA.Cn[4].t4 26.5955
R19578 XA.Cn[4].n3 XA.Cn[4].t9 24.9236
R19579 XA.Cn[4].n3 XA.Cn[4].t8 24.9236
R19580 XA.Cn[4].n4 XA.Cn[4].t11 24.9236
R19581 XA.Cn[4].n4 XA.Cn[4].t10 24.9236
R19582 XA.Cn[4].n5 XA.Cn[4].t2 24.9236
R19583 XA.Cn[4].n5 XA.Cn[4].t1 24.9236
R19584 XA.Cn[4].n6 XA.Cn[4].t0 24.9236
R19585 XA.Cn[4].n6 XA.Cn[4].t3 24.9236
R19586 XA.Cn[4].n60 XA.Cn[4].n2 18.5605
R19587 XA.Cn[4].n60 XA.Cn[4].n59 11.5205
R19588 XA.Cn[4].n58 XA.Cn[4] 4.63701
R19589 XA.Cn[4].n59 XA.Cn[4].n58 3.1844
R19590 XA.Cn[4].n15 XA.Cn[4] 0.931056
R19591 XA.Cn[4].n18 XA.Cn[4] 0.931056
R19592 XA.Cn[4].n21 XA.Cn[4] 0.931056
R19593 XA.Cn[4].n24 XA.Cn[4] 0.931056
R19594 XA.Cn[4].n27 XA.Cn[4] 0.931056
R19595 XA.Cn[4].n30 XA.Cn[4] 0.931056
R19596 XA.Cn[4].n33 XA.Cn[4] 0.931056
R19597 XA.Cn[4].n36 XA.Cn[4] 0.931056
R19598 XA.Cn[4].n39 XA.Cn[4] 0.931056
R19599 XA.Cn[4].n42 XA.Cn[4] 0.931056
R19600 XA.Cn[4].n45 XA.Cn[4] 0.931056
R19601 XA.Cn[4].n48 XA.Cn[4] 0.931056
R19602 XA.Cn[4].n51 XA.Cn[4] 0.931056
R19603 XA.Cn[4].n54 XA.Cn[4] 0.931056
R19604 XA.Cn[4].n57 XA.Cn[4] 0.931056
R19605 XA.Cn[4] XA.Cn[4].n60 0.6405
R19606 XA.Cn[4] XA.Cn[4].n12 0.396333
R19607 XA.Cn[4] XA.Cn[4].n15 0.396333
R19608 XA.Cn[4] XA.Cn[4].n18 0.396333
R19609 XA.Cn[4] XA.Cn[4].n21 0.396333
R19610 XA.Cn[4] XA.Cn[4].n24 0.396333
R19611 XA.Cn[4] XA.Cn[4].n27 0.396333
R19612 XA.Cn[4] XA.Cn[4].n30 0.396333
R19613 XA.Cn[4] XA.Cn[4].n33 0.396333
R19614 XA.Cn[4] XA.Cn[4].n36 0.396333
R19615 XA.Cn[4] XA.Cn[4].n39 0.396333
R19616 XA.Cn[4] XA.Cn[4].n42 0.396333
R19617 XA.Cn[4] XA.Cn[4].n45 0.396333
R19618 XA.Cn[4] XA.Cn[4].n48 0.396333
R19619 XA.Cn[4] XA.Cn[4].n51 0.396333
R19620 XA.Cn[4] XA.Cn[4].n54 0.396333
R19621 XA.Cn[4] XA.Cn[4].n57 0.396333
R19622 XA.Cn[4].n11 XA.Cn[4] 0.104667
R19623 XA.Cn[4].n14 XA.Cn[4] 0.104667
R19624 XA.Cn[4].n17 XA.Cn[4] 0.104667
R19625 XA.Cn[4].n20 XA.Cn[4] 0.104667
R19626 XA.Cn[4].n23 XA.Cn[4] 0.104667
R19627 XA.Cn[4].n26 XA.Cn[4] 0.104667
R19628 XA.Cn[4].n29 XA.Cn[4] 0.104667
R19629 XA.Cn[4].n32 XA.Cn[4] 0.104667
R19630 XA.Cn[4].n35 XA.Cn[4] 0.104667
R19631 XA.Cn[4].n38 XA.Cn[4] 0.104667
R19632 XA.Cn[4].n41 XA.Cn[4] 0.104667
R19633 XA.Cn[4].n44 XA.Cn[4] 0.104667
R19634 XA.Cn[4].n47 XA.Cn[4] 0.104667
R19635 XA.Cn[4].n50 XA.Cn[4] 0.104667
R19636 XA.Cn[4].n53 XA.Cn[4] 0.104667
R19637 XA.Cn[4].n56 XA.Cn[4] 0.104667
R19638 XA.Cn[4].n11 XA.Cn[4] 0.0309878
R19639 XA.Cn[4].n14 XA.Cn[4] 0.0309878
R19640 XA.Cn[4].n17 XA.Cn[4] 0.0309878
R19641 XA.Cn[4].n20 XA.Cn[4] 0.0309878
R19642 XA.Cn[4].n23 XA.Cn[4] 0.0309878
R19643 XA.Cn[4].n26 XA.Cn[4] 0.0309878
R19644 XA.Cn[4].n29 XA.Cn[4] 0.0309878
R19645 XA.Cn[4].n32 XA.Cn[4] 0.0309878
R19646 XA.Cn[4].n35 XA.Cn[4] 0.0309878
R19647 XA.Cn[4].n38 XA.Cn[4] 0.0309878
R19648 XA.Cn[4].n41 XA.Cn[4] 0.0309878
R19649 XA.Cn[4].n44 XA.Cn[4] 0.0309878
R19650 XA.Cn[4].n47 XA.Cn[4] 0.0309878
R19651 XA.Cn[4].n50 XA.Cn[4] 0.0309878
R19652 XA.Cn[4].n53 XA.Cn[4] 0.0309878
R19653 XA.Cn[4].n56 XA.Cn[4] 0.0309878
R19654 XA.Cn[4].n12 XA.Cn[4].n11 0.027939
R19655 XA.Cn[4].n15 XA.Cn[4].n14 0.027939
R19656 XA.Cn[4].n18 XA.Cn[4].n17 0.027939
R19657 XA.Cn[4].n21 XA.Cn[4].n20 0.027939
R19658 XA.Cn[4].n24 XA.Cn[4].n23 0.027939
R19659 XA.Cn[4].n27 XA.Cn[4].n26 0.027939
R19660 XA.Cn[4].n30 XA.Cn[4].n29 0.027939
R19661 XA.Cn[4].n33 XA.Cn[4].n32 0.027939
R19662 XA.Cn[4].n36 XA.Cn[4].n35 0.027939
R19663 XA.Cn[4].n39 XA.Cn[4].n38 0.027939
R19664 XA.Cn[4].n42 XA.Cn[4].n41 0.027939
R19665 XA.Cn[4].n45 XA.Cn[4].n44 0.027939
R19666 XA.Cn[4].n48 XA.Cn[4].n47 0.027939
R19667 XA.Cn[4].n51 XA.Cn[4].n50 0.027939
R19668 XA.Cn[4].n54 XA.Cn[4].n53 0.027939
R19669 XA.Cn[4].n57 XA.Cn[4].n56 0.027939
R19670 XA.Cn[4].n58 XA.Cn[4] 0.0129465
R19671 XA.Cn[2].n2 XA.Cn[2].n1 332.332
R19672 XA.Cn[2].n2 XA.Cn[2].n0 296.493
R19673 XA.Cn[2].n12 XA.Cn[2].n10 161.406
R19674 XA.Cn[2].n15 XA.Cn[2].n13 161.406
R19675 XA.Cn[2].n18 XA.Cn[2].n16 161.406
R19676 XA.Cn[2].n21 XA.Cn[2].n19 161.406
R19677 XA.Cn[2].n24 XA.Cn[2].n22 161.406
R19678 XA.Cn[2].n27 XA.Cn[2].n25 161.406
R19679 XA.Cn[2].n30 XA.Cn[2].n28 161.406
R19680 XA.Cn[2].n33 XA.Cn[2].n31 161.406
R19681 XA.Cn[2].n36 XA.Cn[2].n34 161.406
R19682 XA.Cn[2].n39 XA.Cn[2].n37 161.406
R19683 XA.Cn[2].n42 XA.Cn[2].n40 161.406
R19684 XA.Cn[2].n45 XA.Cn[2].n43 161.406
R19685 XA.Cn[2].n48 XA.Cn[2].n46 161.406
R19686 XA.Cn[2].n51 XA.Cn[2].n49 161.406
R19687 XA.Cn[2].n54 XA.Cn[2].n52 161.406
R19688 XA.Cn[2].n57 XA.Cn[2].n55 161.406
R19689 XA.Cn[2].n10 XA.Cn[2].t18 161.202
R19690 XA.Cn[2].n13 XA.Cn[2].t35 161.202
R19691 XA.Cn[2].n16 XA.Cn[2].t37 161.202
R19692 XA.Cn[2].n19 XA.Cn[2].t39 161.202
R19693 XA.Cn[2].n22 XA.Cn[2].t28 161.202
R19694 XA.Cn[2].n25 XA.Cn[2].t29 161.202
R19695 XA.Cn[2].n28 XA.Cn[2].t42 161.202
R19696 XA.Cn[2].n31 XA.Cn[2].t19 161.202
R19697 XA.Cn[2].n34 XA.Cn[2].t21 161.202
R19698 XA.Cn[2].n37 XA.Cn[2].t40 161.202
R19699 XA.Cn[2].n40 XA.Cn[2].t41 161.202
R19700 XA.Cn[2].n43 XA.Cn[2].t22 161.202
R19701 XA.Cn[2].n46 XA.Cn[2].t30 161.202
R19702 XA.Cn[2].n49 XA.Cn[2].t33 161.202
R19703 XA.Cn[2].n52 XA.Cn[2].t14 161.202
R19704 XA.Cn[2].n55 XA.Cn[2].t24 161.202
R19705 XA.Cn[2].n10 XA.Cn[2].t20 145.137
R19706 XA.Cn[2].n13 XA.Cn[2].t38 145.137
R19707 XA.Cn[2].n16 XA.Cn[2].t43 145.137
R19708 XA.Cn[2].n19 XA.Cn[2].t12 145.137
R19709 XA.Cn[2].n22 XA.Cn[2].t31 145.137
R19710 XA.Cn[2].n25 XA.Cn[2].t32 145.137
R19711 XA.Cn[2].n28 XA.Cn[2].t16 145.137
R19712 XA.Cn[2].n31 XA.Cn[2].t23 145.137
R19713 XA.Cn[2].n34 XA.Cn[2].t25 145.137
R19714 XA.Cn[2].n37 XA.Cn[2].t13 145.137
R19715 XA.Cn[2].n40 XA.Cn[2].t15 145.137
R19716 XA.Cn[2].n43 XA.Cn[2].t26 145.137
R19717 XA.Cn[2].n46 XA.Cn[2].t34 145.137
R19718 XA.Cn[2].n49 XA.Cn[2].t36 145.137
R19719 XA.Cn[2].n52 XA.Cn[2].t17 145.137
R19720 XA.Cn[2].n55 XA.Cn[2].t27 145.137
R19721 XA.Cn[2].n7 XA.Cn[2].n6 135.248
R19722 XA.Cn[2].n9 XA.Cn[2].n3 98.982
R19723 XA.Cn[2].n8 XA.Cn[2].n4 98.982
R19724 XA.Cn[2].n7 XA.Cn[2].n5 98.982
R19725 XA.Cn[2].n9 XA.Cn[2].n8 36.2672
R19726 XA.Cn[2].n8 XA.Cn[2].n7 36.2672
R19727 XA.Cn[2].n59 XA.Cn[2].n9 32.6405
R19728 XA.Cn[2].n1 XA.Cn[2].t7 26.5955
R19729 XA.Cn[2].n1 XA.Cn[2].t6 26.5955
R19730 XA.Cn[2].n0 XA.Cn[2].t9 26.5955
R19731 XA.Cn[2].n0 XA.Cn[2].t8 26.5955
R19732 XA.Cn[2].n3 XA.Cn[2].t5 24.9236
R19733 XA.Cn[2].n3 XA.Cn[2].t4 24.9236
R19734 XA.Cn[2].n4 XA.Cn[2].t3 24.9236
R19735 XA.Cn[2].n4 XA.Cn[2].t2 24.9236
R19736 XA.Cn[2].n5 XA.Cn[2].t1 24.9236
R19737 XA.Cn[2].n5 XA.Cn[2].t10 24.9236
R19738 XA.Cn[2].n6 XA.Cn[2].t11 24.9236
R19739 XA.Cn[2].n6 XA.Cn[2].t0 24.9236
R19740 XA.Cn[2].n60 XA.Cn[2].n2 18.5605
R19741 XA.Cn[2].n60 XA.Cn[2].n59 11.5205
R19742 XA.Cn[2].n58 XA.Cn[2] 6.32799
R19743 XA.Cn[2].n59 XA.Cn[2].n58 3.18175
R19744 XA.Cn[2].n15 XA.Cn[2] 0.931056
R19745 XA.Cn[2].n18 XA.Cn[2] 0.931056
R19746 XA.Cn[2].n21 XA.Cn[2] 0.931056
R19747 XA.Cn[2].n24 XA.Cn[2] 0.931056
R19748 XA.Cn[2].n27 XA.Cn[2] 0.931056
R19749 XA.Cn[2].n30 XA.Cn[2] 0.931056
R19750 XA.Cn[2].n33 XA.Cn[2] 0.931056
R19751 XA.Cn[2].n36 XA.Cn[2] 0.931056
R19752 XA.Cn[2].n39 XA.Cn[2] 0.931056
R19753 XA.Cn[2].n42 XA.Cn[2] 0.931056
R19754 XA.Cn[2].n45 XA.Cn[2] 0.931056
R19755 XA.Cn[2].n48 XA.Cn[2] 0.931056
R19756 XA.Cn[2].n51 XA.Cn[2] 0.931056
R19757 XA.Cn[2].n54 XA.Cn[2] 0.931056
R19758 XA.Cn[2].n57 XA.Cn[2] 0.931056
R19759 XA.Cn[2] XA.Cn[2].n60 0.6405
R19760 XA.Cn[2] XA.Cn[2].n12 0.396333
R19761 XA.Cn[2] XA.Cn[2].n15 0.396333
R19762 XA.Cn[2] XA.Cn[2].n18 0.396333
R19763 XA.Cn[2] XA.Cn[2].n21 0.396333
R19764 XA.Cn[2] XA.Cn[2].n24 0.396333
R19765 XA.Cn[2] XA.Cn[2].n27 0.396333
R19766 XA.Cn[2] XA.Cn[2].n30 0.396333
R19767 XA.Cn[2] XA.Cn[2].n33 0.396333
R19768 XA.Cn[2] XA.Cn[2].n36 0.396333
R19769 XA.Cn[2] XA.Cn[2].n39 0.396333
R19770 XA.Cn[2] XA.Cn[2].n42 0.396333
R19771 XA.Cn[2] XA.Cn[2].n45 0.396333
R19772 XA.Cn[2] XA.Cn[2].n48 0.396333
R19773 XA.Cn[2] XA.Cn[2].n51 0.396333
R19774 XA.Cn[2] XA.Cn[2].n54 0.396333
R19775 XA.Cn[2] XA.Cn[2].n57 0.396333
R19776 XA.Cn[2].n11 XA.Cn[2] 0.104667
R19777 XA.Cn[2].n14 XA.Cn[2] 0.104667
R19778 XA.Cn[2].n17 XA.Cn[2] 0.104667
R19779 XA.Cn[2].n20 XA.Cn[2] 0.104667
R19780 XA.Cn[2].n23 XA.Cn[2] 0.104667
R19781 XA.Cn[2].n26 XA.Cn[2] 0.104667
R19782 XA.Cn[2].n29 XA.Cn[2] 0.104667
R19783 XA.Cn[2].n32 XA.Cn[2] 0.104667
R19784 XA.Cn[2].n35 XA.Cn[2] 0.104667
R19785 XA.Cn[2].n38 XA.Cn[2] 0.104667
R19786 XA.Cn[2].n41 XA.Cn[2] 0.104667
R19787 XA.Cn[2].n44 XA.Cn[2] 0.104667
R19788 XA.Cn[2].n47 XA.Cn[2] 0.104667
R19789 XA.Cn[2].n50 XA.Cn[2] 0.104667
R19790 XA.Cn[2].n53 XA.Cn[2] 0.104667
R19791 XA.Cn[2].n56 XA.Cn[2] 0.104667
R19792 XA.Cn[2].n11 XA.Cn[2] 0.0309878
R19793 XA.Cn[2].n14 XA.Cn[2] 0.0309878
R19794 XA.Cn[2].n17 XA.Cn[2] 0.0309878
R19795 XA.Cn[2].n20 XA.Cn[2] 0.0309878
R19796 XA.Cn[2].n23 XA.Cn[2] 0.0309878
R19797 XA.Cn[2].n26 XA.Cn[2] 0.0309878
R19798 XA.Cn[2].n29 XA.Cn[2] 0.0309878
R19799 XA.Cn[2].n32 XA.Cn[2] 0.0309878
R19800 XA.Cn[2].n35 XA.Cn[2] 0.0309878
R19801 XA.Cn[2].n38 XA.Cn[2] 0.0309878
R19802 XA.Cn[2].n41 XA.Cn[2] 0.0309878
R19803 XA.Cn[2].n44 XA.Cn[2] 0.0309878
R19804 XA.Cn[2].n47 XA.Cn[2] 0.0309878
R19805 XA.Cn[2].n50 XA.Cn[2] 0.0309878
R19806 XA.Cn[2].n53 XA.Cn[2] 0.0309878
R19807 XA.Cn[2].n56 XA.Cn[2] 0.0309878
R19808 XA.Cn[2].n12 XA.Cn[2].n11 0.027939
R19809 XA.Cn[2].n15 XA.Cn[2].n14 0.027939
R19810 XA.Cn[2].n18 XA.Cn[2].n17 0.027939
R19811 XA.Cn[2].n21 XA.Cn[2].n20 0.027939
R19812 XA.Cn[2].n24 XA.Cn[2].n23 0.027939
R19813 XA.Cn[2].n27 XA.Cn[2].n26 0.027939
R19814 XA.Cn[2].n30 XA.Cn[2].n29 0.027939
R19815 XA.Cn[2].n33 XA.Cn[2].n32 0.027939
R19816 XA.Cn[2].n36 XA.Cn[2].n35 0.027939
R19817 XA.Cn[2].n39 XA.Cn[2].n38 0.027939
R19818 XA.Cn[2].n42 XA.Cn[2].n41 0.027939
R19819 XA.Cn[2].n45 XA.Cn[2].n44 0.027939
R19820 XA.Cn[2].n48 XA.Cn[2].n47 0.027939
R19821 XA.Cn[2].n51 XA.Cn[2].n50 0.027939
R19822 XA.Cn[2].n54 XA.Cn[2].n53 0.027939
R19823 XA.Cn[2].n57 XA.Cn[2].n56 0.027939
R19824 XA.Cn[2].n58 XA.Cn[2] 0.0156819
R19825 Vbias.n512 Vbias.t2 651.571
R19826 Vbias.n512 Vbias.t0 651.571
R19827 Vbias.n513 Vbias.t1 651.571
R19828 Vbias.n513 Vbias.t5 651.571
R19829 Vbias.n509 Vbias.t181 119.309
R19830 Vbias.n507 Vbias.t24 119.309
R19831 Vbias.n505 Vbias.t12 119.309
R19832 Vbias.n503 Vbias.t248 119.309
R19833 Vbias.n501 Vbias.t95 119.309
R19834 Vbias.n499 Vbias.t75 119.309
R19835 Vbias.n497 Vbias.t246 119.309
R19836 Vbias.n495 Vbias.t169 119.309
R19837 Vbias.n493 Vbias.t147 119.309
R19838 Vbias.n491 Vbias.t60 119.309
R19839 Vbias.n489 Vbias.t227 119.309
R19840 Vbias.n487 Vbias.t141 119.309
R19841 Vbias.n485 Vbias.t56 119.309
R19842 Vbias.n483 Vbias.t41 119.309
R19843 Vbias.n481 Vbias.t201 119.309
R19844 Vbias.n480 Vbias.t129 119.309
R19845 Vbias.n477 Vbias.t110 119.309
R19846 Vbias.n475 Vbias.t210 119.309
R19847 Vbias.n473 Vbias.t193 119.309
R19848 Vbias.n471 Vbias.t173 119.309
R19849 Vbias.n469 Vbias.t25 119.309
R19850 Vbias.n467 Vbias.t258 119.309
R19851 Vbias.n465 Vbias.t171 119.309
R19852 Vbias.n463 Vbias.t96 119.309
R19853 Vbias.n461 Vbias.t76 119.309
R19854 Vbias.n459 Vbias.t247 119.309
R19855 Vbias.n457 Vbias.t156 119.309
R19856 Vbias.n455 Vbias.t69 119.309
R19857 Vbias.n453 Vbias.t242 119.309
R19858 Vbias.n451 Vbias.t229 119.309
R19859 Vbias.n449 Vbias.t130 119.309
R19860 Vbias.n448 Vbias.t57 119.309
R19861 Vbias.n445 Vbias.t146 119.309
R19862 Vbias.n443 Vbias.t238 119.309
R19863 Vbias.n441 Vbias.t225 119.309
R19864 Vbias.n439 Vbias.t205 119.309
R19865 Vbias.n437 Vbias.t52 119.309
R19866 Vbias.n435 Vbias.t32 119.309
R19867 Vbias.n433 Vbias.t199 119.309
R19868 Vbias.n431 Vbias.t125 119.309
R19869 Vbias.n429 Vbias.t102 119.309
R19870 Vbias.n427 Vbias.t18 119.309
R19871 Vbias.n425 Vbias.t183 119.309
R19872 Vbias.n423 Vbias.t99 119.309
R19873 Vbias.n421 Vbias.t14 119.309
R19874 Vbias.n419 Vbias.t261 119.309
R19875 Vbias.n417 Vbias.t160 119.309
R19876 Vbias.n416 Vbias.t87 119.309
R19877 Vbias.n413 Vbias.t73 119.309
R19878 Vbias.n411 Vbias.t165 119.309
R19879 Vbias.n409 Vbias.t153 119.309
R19880 Vbias.n407 Vbias.t133 119.309
R19881 Vbias.n405 Vbias.t239 119.309
R19882 Vbias.n403 Vbias.t217 119.309
R19883 Vbias.n401 Vbias.t126 119.309
R19884 Vbias.n399 Vbias.t53 119.309
R19885 Vbias.n397 Vbias.t33 119.309
R19886 Vbias.n395 Vbias.t200 119.309
R19887 Vbias.n393 Vbias.t112 119.309
R19888 Vbias.n391 Vbias.t29 119.309
R19889 Vbias.n389 Vbias.t196 119.309
R19890 Vbias.n387 Vbias.t185 119.309
R19891 Vbias.n385 Vbias.t88 119.309
R19892 Vbias.n384 Vbias.t16 119.309
R19893 Vbias.n381 Vbias.t255 119.309
R19894 Vbias.n379 Vbias.t92 119.309
R19895 Vbias.n377 Vbias.t81 119.309
R19896 Vbias.n375 Vbias.t62 119.309
R19897 Vbias.n373 Vbias.t166 119.309
R19898 Vbias.n371 Vbias.t144 119.309
R19899 Vbias.n369 Vbias.t54 119.309
R19900 Vbias.n367 Vbias.t240 119.309
R19901 Vbias.n365 Vbias.t219 119.309
R19902 Vbias.n363 Vbias.t127 119.309
R19903 Vbias.n361 Vbias.t40 119.309
R19904 Vbias.n359 Vbias.t213 119.309
R19905 Vbias.n357 Vbias.t124 119.309
R19906 Vbias.n355 Vbias.t113 119.309
R19907 Vbias.n353 Vbias.t17 119.309
R19908 Vbias.n352 Vbias.t198 119.309
R19909 Vbias.n349 Vbias.t176 119.309
R19910 Vbias.n347 Vbias.t20 119.309
R19911 Vbias.n345 Vbias.t7 119.309
R19912 Vbias.n343 Vbias.t243 119.309
R19913 Vbias.n341 Vbias.t90 119.309
R19914 Vbias.n339 Vbias.t65 119.309
R19915 Vbias.n337 Vbias.t236 119.309
R19916 Vbias.n335 Vbias.t163 119.309
R19917 Vbias.n333 Vbias.t138 119.309
R19918 Vbias.n331 Vbias.t50 119.309
R19919 Vbias.n329 Vbias.t221 119.309
R19920 Vbias.n327 Vbias.t135 119.309
R19921 Vbias.n325 Vbias.t48 119.309
R19922 Vbias.n323 Vbias.t37 119.309
R19923 Vbias.n321 Vbias.t195 119.309
R19924 Vbias.n320 Vbias.t121 119.309
R19925 Vbias.n317 Vbias.t105 119.309
R19926 Vbias.n315 Vbias.t204 119.309
R19927 Vbias.n313 Vbias.t187 119.309
R19928 Vbias.n311 Vbias.t168 119.309
R19929 Vbias.n309 Vbias.t21 119.309
R19930 Vbias.n307 Vbias.t251 119.309
R19931 Vbias.n305 Vbias.t164 119.309
R19932 Vbias.n303 Vbias.t91 119.309
R19933 Vbias.n301 Vbias.t68 119.309
R19934 Vbias.n299 Vbias.t237 119.309
R19935 Vbias.n297 Vbias.t150 119.309
R19936 Vbias.n295 Vbias.t63 119.309
R19937 Vbias.n293 Vbias.t235 119.309
R19938 Vbias.n291 Vbias.t222 119.309
R19939 Vbias.n289 Vbias.t122 119.309
R19940 Vbias.n288 Vbias.t49 119.309
R19941 Vbias.n285 Vbias.t137 119.309
R19942 Vbias.n283 Vbias.t232 119.309
R19943 Vbias.n281 Vbias.t220 119.309
R19944 Vbias.n279 Vbias.t197 119.309
R19945 Vbias.n277 Vbias.t44 119.309
R19946 Vbias.n275 Vbias.t27 119.309
R19947 Vbias.n273 Vbias.t190 119.309
R19948 Vbias.n271 Vbias.t118 119.309
R19949 Vbias.n269 Vbias.t98 119.309
R19950 Vbias.n267 Vbias.t11 119.309
R19951 Vbias.n265 Vbias.t179 119.309
R19952 Vbias.n263 Vbias.t93 119.309
R19953 Vbias.n261 Vbias.t8 119.309
R19954 Vbias.n259 Vbias.t257 119.309
R19955 Vbias.n257 Vbias.t154 119.309
R19956 Vbias.n256 Vbias.t82 119.309
R19957 Vbias.n253 Vbias.t64 119.309
R19958 Vbias.n251 Vbias.t161 119.309
R19959 Vbias.n249 Vbias.t149 119.309
R19960 Vbias.n247 Vbias.t123 119.309
R19961 Vbias.n245 Vbias.t233 119.309
R19962 Vbias.n243 Vbias.t211 119.309
R19963 Vbias.n241 Vbias.t119 119.309
R19964 Vbias.n239 Vbias.t45 119.309
R19965 Vbias.n237 Vbias.t28 119.309
R19966 Vbias.n235 Vbias.t192 119.309
R19967 Vbias.n233 Vbias.t107 119.309
R19968 Vbias.n231 Vbias.t23 119.309
R19969 Vbias.n229 Vbias.t188 119.309
R19970 Vbias.n227 Vbias.t180 119.309
R19971 Vbias.n225 Vbias.t83 119.309
R19972 Vbias.n224 Vbias.t9 119.309
R19973 Vbias.n221 Vbias.t250 119.309
R19974 Vbias.n219 Vbias.t89 119.309
R19975 Vbias.n217 Vbias.t80 119.309
R19976 Vbias.n215 Vbias.t51 119.309
R19977 Vbias.n213 Vbias.t162 119.309
R19978 Vbias.n211 Vbias.t136 119.309
R19979 Vbias.n209 Vbias.t46 119.309
R19980 Vbias.n207 Vbias.t234 119.309
R19981 Vbias.n205 Vbias.t212 119.309
R19982 Vbias.n203 Vbias.t120 119.309
R19983 Vbias.n201 Vbias.t36 119.309
R19984 Vbias.n199 Vbias.t208 119.309
R19985 Vbias.n197 Vbias.t117 119.309
R19986 Vbias.n195 Vbias.t108 119.309
R19987 Vbias.n193 Vbias.t10 119.309
R19988 Vbias.n192 Vbias.t189 119.309
R19989 Vbias.n189 Vbias.t109 119.309
R19990 Vbias.n187 Vbias.t207 119.309
R19991 Vbias.n185 Vbias.t191 119.309
R19992 Vbias.n183 Vbias.t172 119.309
R19993 Vbias.n181 Vbias.t22 119.309
R19994 Vbias.n179 Vbias.t256 119.309
R19995 Vbias.n177 Vbias.t167 119.309
R19996 Vbias.n175 Vbias.t94 119.309
R19997 Vbias.n173 Vbias.t74 119.309
R19998 Vbias.n171 Vbias.t244 119.309
R19999 Vbias.n169 Vbias.t155 119.309
R20000 Vbias.n167 Vbias.t66 119.309
R20001 Vbias.n165 Vbias.t241 119.309
R20002 Vbias.n163 Vbias.t226 119.309
R20003 Vbias.n161 Vbias.t128 119.309
R20004 Vbias.n160 Vbias.t55 119.309
R20005 Vbias.n157 Vbias.t249 119.309
R20006 Vbias.n155 Vbias.t85 119.309
R20007 Vbias.n153 Vbias.t78 119.309
R20008 Vbias.n151 Vbias.t47 119.309
R20009 Vbias.n149 Vbias.t159 119.309
R20010 Vbias.n147 Vbias.t134 119.309
R20011 Vbias.n145 Vbias.t43 119.309
R20012 Vbias.n143 Vbias.t231 119.309
R20013 Vbias.n141 Vbias.t209 119.309
R20014 Vbias.n139 Vbias.t116 119.309
R20015 Vbias.n137 Vbias.t34 119.309
R20016 Vbias.n135 Vbias.t206 119.309
R20017 Vbias.n133 Vbias.t115 119.309
R20018 Vbias.n131 Vbias.t103 119.309
R20019 Vbias.n129 Vbias.t6 119.309
R20020 Vbias.n128 Vbias.t186 119.309
R20021 Vbias.n125 Vbias.t86 119.309
R20022 Vbias.n123 Vbias.t175 119.309
R20023 Vbias.n121 Vbias.t170 119.309
R20024 Vbias.n119 Vbias.t148 119.309
R20025 Vbias.n117 Vbias.t252 119.309
R20026 Vbias.n115 Vbias.t228 119.309
R20027 Vbias.n113 Vbias.t143 119.309
R20028 Vbias.n111 Vbias.t70 119.309
R20029 Vbias.n109 Vbias.t42 119.309
R20030 Vbias.n107 Vbias.t218 119.309
R20031 Vbias.n105 Vbias.t131 119.309
R20032 Vbias.n103 Vbias.t38 119.309
R20033 Vbias.n101 Vbias.t214 119.309
R20034 Vbias.n99 Vbias.t203 119.309
R20035 Vbias.n97 Vbias.t100 119.309
R20036 Vbias.n96 Vbias.t30 119.309
R20037 Vbias.n93 Vbias.t13 119.309
R20038 Vbias.n91 Vbias.t104 119.309
R20039 Vbias.n89 Vbias.t97 119.309
R20040 Vbias.n87 Vbias.t77 119.309
R20041 Vbias.n85 Vbias.t177 119.309
R20042 Vbias.n83 Vbias.t157 119.309
R20043 Vbias.n81 Vbias.t71 119.309
R20044 Vbias.n79 Vbias.t253 119.309
R20045 Vbias.n77 Vbias.t230 119.309
R20046 Vbias.n75 Vbias.t145 119.309
R20047 Vbias.n73 Vbias.t58 119.309
R20048 Vbias.n71 Vbias.t224 119.309
R20049 Vbias.n69 Vbias.t139 119.309
R20050 Vbias.n67 Vbias.t132 119.309
R20051 Vbias.n65 Vbias.t31 119.309
R20052 Vbias.n64 Vbias.t215 119.309
R20053 Vbias.n61 Vbias.t194 119.309
R20054 Vbias.n59 Vbias.t35 119.309
R20055 Vbias.n57 Vbias.t26 119.309
R20056 Vbias.n55 Vbias.t259 119.309
R20057 Vbias.n53 Vbias.t106 119.309
R20058 Vbias.n51 Vbias.t84 119.309
R20059 Vbias.n49 Vbias.t254 119.309
R20060 Vbias.n47 Vbias.t178 119.309
R20061 Vbias.n45 Vbias.t158 119.309
R20062 Vbias.n43 Vbias.t72 119.309
R20063 Vbias.n41 Vbias.t245 119.309
R20064 Vbias.n39 Vbias.t152 119.309
R20065 Vbias.n37 Vbias.t67 119.309
R20066 Vbias.n35 Vbias.t59 119.309
R20067 Vbias.n33 Vbias.t216 119.309
R20068 Vbias.n32 Vbias.t140 119.309
R20069 Vbias.n29 Vbias.t61 119.309
R20070 Vbias.n27 Vbias.t151 119.309
R20071 Vbias.n25 Vbias.t142 119.309
R20072 Vbias.n23 Vbias.t114 119.309
R20073 Vbias.n21 Vbias.t223 119.309
R20074 Vbias.n19 Vbias.t202 119.309
R20075 Vbias.n17 Vbias.t111 119.309
R20076 Vbias.n15 Vbias.t39 119.309
R20077 Vbias.n13 Vbias.t19 119.309
R20078 Vbias.n11 Vbias.t184 119.309
R20079 Vbias.n9 Vbias.t101 119.309
R20080 Vbias.n7 Vbias.t15 119.309
R20081 Vbias.n5 Vbias.t182 119.309
R20082 Vbias.n3 Vbias.t174 119.309
R20083 Vbias.n1 Vbias.t79 119.309
R20084 Vbias.n0 Vbias.t260 119.309
R20085 Vbias.n515 Vbias.t3 77.1775
R20086 Vbias.n515 Vbias.t4 34.3847
R20087 Vbias Vbias.n480 8.00727
R20088 Vbias Vbias.n448 8.00727
R20089 Vbias Vbias.n416 8.00727
R20090 Vbias Vbias.n384 8.00727
R20091 Vbias Vbias.n352 8.00727
R20092 Vbias Vbias.n320 8.00727
R20093 Vbias Vbias.n288 8.00727
R20094 Vbias Vbias.n256 8.00727
R20095 Vbias Vbias.n224 8.00727
R20096 Vbias Vbias.n192 8.00727
R20097 Vbias Vbias.n160 8.00727
R20098 Vbias Vbias.n128 8.00727
R20099 Vbias Vbias.n96 8.00727
R20100 Vbias Vbias.n64 8.00727
R20101 Vbias Vbias.n32 8.00727
R20102 Vbias Vbias.n0 8.00727
R20103 Vbias.n510 Vbias.n509 7.9105
R20104 Vbias.n508 Vbias.n507 7.9105
R20105 Vbias.n506 Vbias.n505 7.9105
R20106 Vbias.n504 Vbias.n503 7.9105
R20107 Vbias.n502 Vbias.n501 7.9105
R20108 Vbias.n500 Vbias.n499 7.9105
R20109 Vbias.n498 Vbias.n497 7.9105
R20110 Vbias.n496 Vbias.n495 7.9105
R20111 Vbias.n494 Vbias.n493 7.9105
R20112 Vbias.n492 Vbias.n491 7.9105
R20113 Vbias.n490 Vbias.n489 7.9105
R20114 Vbias.n488 Vbias.n487 7.9105
R20115 Vbias.n486 Vbias.n485 7.9105
R20116 Vbias.n484 Vbias.n483 7.9105
R20117 Vbias.n482 Vbias.n481 7.9105
R20118 Vbias.n478 Vbias.n477 7.9105
R20119 Vbias.n476 Vbias.n475 7.9105
R20120 Vbias.n474 Vbias.n473 7.9105
R20121 Vbias.n472 Vbias.n471 7.9105
R20122 Vbias.n470 Vbias.n469 7.9105
R20123 Vbias.n468 Vbias.n467 7.9105
R20124 Vbias.n466 Vbias.n465 7.9105
R20125 Vbias.n464 Vbias.n463 7.9105
R20126 Vbias.n462 Vbias.n461 7.9105
R20127 Vbias.n460 Vbias.n459 7.9105
R20128 Vbias.n458 Vbias.n457 7.9105
R20129 Vbias.n456 Vbias.n455 7.9105
R20130 Vbias.n454 Vbias.n453 7.9105
R20131 Vbias.n452 Vbias.n451 7.9105
R20132 Vbias.n450 Vbias.n449 7.9105
R20133 Vbias.n446 Vbias.n445 7.9105
R20134 Vbias.n444 Vbias.n443 7.9105
R20135 Vbias.n442 Vbias.n441 7.9105
R20136 Vbias.n440 Vbias.n439 7.9105
R20137 Vbias.n438 Vbias.n437 7.9105
R20138 Vbias.n436 Vbias.n435 7.9105
R20139 Vbias.n434 Vbias.n433 7.9105
R20140 Vbias.n432 Vbias.n431 7.9105
R20141 Vbias.n430 Vbias.n429 7.9105
R20142 Vbias.n428 Vbias.n427 7.9105
R20143 Vbias.n426 Vbias.n425 7.9105
R20144 Vbias.n424 Vbias.n423 7.9105
R20145 Vbias.n422 Vbias.n421 7.9105
R20146 Vbias.n420 Vbias.n419 7.9105
R20147 Vbias.n418 Vbias.n417 7.9105
R20148 Vbias.n414 Vbias.n413 7.9105
R20149 Vbias.n412 Vbias.n411 7.9105
R20150 Vbias.n410 Vbias.n409 7.9105
R20151 Vbias.n408 Vbias.n407 7.9105
R20152 Vbias.n406 Vbias.n405 7.9105
R20153 Vbias.n404 Vbias.n403 7.9105
R20154 Vbias.n402 Vbias.n401 7.9105
R20155 Vbias.n400 Vbias.n399 7.9105
R20156 Vbias.n398 Vbias.n397 7.9105
R20157 Vbias.n396 Vbias.n395 7.9105
R20158 Vbias.n394 Vbias.n393 7.9105
R20159 Vbias.n392 Vbias.n391 7.9105
R20160 Vbias.n390 Vbias.n389 7.9105
R20161 Vbias.n388 Vbias.n387 7.9105
R20162 Vbias.n386 Vbias.n385 7.9105
R20163 Vbias.n382 Vbias.n381 7.9105
R20164 Vbias.n380 Vbias.n379 7.9105
R20165 Vbias.n378 Vbias.n377 7.9105
R20166 Vbias.n376 Vbias.n375 7.9105
R20167 Vbias.n374 Vbias.n373 7.9105
R20168 Vbias.n372 Vbias.n371 7.9105
R20169 Vbias.n370 Vbias.n369 7.9105
R20170 Vbias.n368 Vbias.n367 7.9105
R20171 Vbias.n366 Vbias.n365 7.9105
R20172 Vbias.n364 Vbias.n363 7.9105
R20173 Vbias.n362 Vbias.n361 7.9105
R20174 Vbias.n360 Vbias.n359 7.9105
R20175 Vbias.n358 Vbias.n357 7.9105
R20176 Vbias.n356 Vbias.n355 7.9105
R20177 Vbias.n354 Vbias.n353 7.9105
R20178 Vbias.n350 Vbias.n349 7.9105
R20179 Vbias.n348 Vbias.n347 7.9105
R20180 Vbias.n346 Vbias.n345 7.9105
R20181 Vbias.n344 Vbias.n343 7.9105
R20182 Vbias.n342 Vbias.n341 7.9105
R20183 Vbias.n340 Vbias.n339 7.9105
R20184 Vbias.n338 Vbias.n337 7.9105
R20185 Vbias.n336 Vbias.n335 7.9105
R20186 Vbias.n334 Vbias.n333 7.9105
R20187 Vbias.n332 Vbias.n331 7.9105
R20188 Vbias.n330 Vbias.n329 7.9105
R20189 Vbias.n328 Vbias.n327 7.9105
R20190 Vbias.n326 Vbias.n325 7.9105
R20191 Vbias.n324 Vbias.n323 7.9105
R20192 Vbias.n322 Vbias.n321 7.9105
R20193 Vbias.n318 Vbias.n317 7.9105
R20194 Vbias.n316 Vbias.n315 7.9105
R20195 Vbias.n314 Vbias.n313 7.9105
R20196 Vbias.n312 Vbias.n311 7.9105
R20197 Vbias.n310 Vbias.n309 7.9105
R20198 Vbias.n308 Vbias.n307 7.9105
R20199 Vbias.n306 Vbias.n305 7.9105
R20200 Vbias.n304 Vbias.n303 7.9105
R20201 Vbias.n302 Vbias.n301 7.9105
R20202 Vbias.n300 Vbias.n299 7.9105
R20203 Vbias.n298 Vbias.n297 7.9105
R20204 Vbias.n296 Vbias.n295 7.9105
R20205 Vbias.n294 Vbias.n293 7.9105
R20206 Vbias.n292 Vbias.n291 7.9105
R20207 Vbias.n290 Vbias.n289 7.9105
R20208 Vbias.n286 Vbias.n285 7.9105
R20209 Vbias.n284 Vbias.n283 7.9105
R20210 Vbias.n282 Vbias.n281 7.9105
R20211 Vbias.n280 Vbias.n279 7.9105
R20212 Vbias.n278 Vbias.n277 7.9105
R20213 Vbias.n276 Vbias.n275 7.9105
R20214 Vbias.n274 Vbias.n273 7.9105
R20215 Vbias.n272 Vbias.n271 7.9105
R20216 Vbias.n270 Vbias.n269 7.9105
R20217 Vbias.n268 Vbias.n267 7.9105
R20218 Vbias.n266 Vbias.n265 7.9105
R20219 Vbias.n264 Vbias.n263 7.9105
R20220 Vbias.n262 Vbias.n261 7.9105
R20221 Vbias.n260 Vbias.n259 7.9105
R20222 Vbias.n258 Vbias.n257 7.9105
R20223 Vbias.n254 Vbias.n253 7.9105
R20224 Vbias.n252 Vbias.n251 7.9105
R20225 Vbias.n250 Vbias.n249 7.9105
R20226 Vbias.n248 Vbias.n247 7.9105
R20227 Vbias.n246 Vbias.n245 7.9105
R20228 Vbias.n244 Vbias.n243 7.9105
R20229 Vbias.n242 Vbias.n241 7.9105
R20230 Vbias.n240 Vbias.n239 7.9105
R20231 Vbias.n238 Vbias.n237 7.9105
R20232 Vbias.n236 Vbias.n235 7.9105
R20233 Vbias.n234 Vbias.n233 7.9105
R20234 Vbias.n232 Vbias.n231 7.9105
R20235 Vbias.n230 Vbias.n229 7.9105
R20236 Vbias.n228 Vbias.n227 7.9105
R20237 Vbias.n226 Vbias.n225 7.9105
R20238 Vbias.n222 Vbias.n221 7.9105
R20239 Vbias.n220 Vbias.n219 7.9105
R20240 Vbias.n218 Vbias.n217 7.9105
R20241 Vbias.n216 Vbias.n215 7.9105
R20242 Vbias.n214 Vbias.n213 7.9105
R20243 Vbias.n212 Vbias.n211 7.9105
R20244 Vbias.n210 Vbias.n209 7.9105
R20245 Vbias.n208 Vbias.n207 7.9105
R20246 Vbias.n206 Vbias.n205 7.9105
R20247 Vbias.n204 Vbias.n203 7.9105
R20248 Vbias.n202 Vbias.n201 7.9105
R20249 Vbias.n200 Vbias.n199 7.9105
R20250 Vbias.n198 Vbias.n197 7.9105
R20251 Vbias.n196 Vbias.n195 7.9105
R20252 Vbias.n194 Vbias.n193 7.9105
R20253 Vbias.n190 Vbias.n189 7.9105
R20254 Vbias.n188 Vbias.n187 7.9105
R20255 Vbias.n186 Vbias.n185 7.9105
R20256 Vbias.n184 Vbias.n183 7.9105
R20257 Vbias.n182 Vbias.n181 7.9105
R20258 Vbias.n180 Vbias.n179 7.9105
R20259 Vbias.n178 Vbias.n177 7.9105
R20260 Vbias.n176 Vbias.n175 7.9105
R20261 Vbias.n174 Vbias.n173 7.9105
R20262 Vbias.n172 Vbias.n171 7.9105
R20263 Vbias.n170 Vbias.n169 7.9105
R20264 Vbias.n168 Vbias.n167 7.9105
R20265 Vbias.n166 Vbias.n165 7.9105
R20266 Vbias.n164 Vbias.n163 7.9105
R20267 Vbias.n162 Vbias.n161 7.9105
R20268 Vbias.n158 Vbias.n157 7.9105
R20269 Vbias.n156 Vbias.n155 7.9105
R20270 Vbias.n154 Vbias.n153 7.9105
R20271 Vbias.n152 Vbias.n151 7.9105
R20272 Vbias.n150 Vbias.n149 7.9105
R20273 Vbias.n148 Vbias.n147 7.9105
R20274 Vbias.n146 Vbias.n145 7.9105
R20275 Vbias.n144 Vbias.n143 7.9105
R20276 Vbias.n142 Vbias.n141 7.9105
R20277 Vbias.n140 Vbias.n139 7.9105
R20278 Vbias.n138 Vbias.n137 7.9105
R20279 Vbias.n136 Vbias.n135 7.9105
R20280 Vbias.n134 Vbias.n133 7.9105
R20281 Vbias.n132 Vbias.n131 7.9105
R20282 Vbias.n130 Vbias.n129 7.9105
R20283 Vbias.n126 Vbias.n125 7.9105
R20284 Vbias.n124 Vbias.n123 7.9105
R20285 Vbias.n122 Vbias.n121 7.9105
R20286 Vbias.n120 Vbias.n119 7.9105
R20287 Vbias.n118 Vbias.n117 7.9105
R20288 Vbias.n116 Vbias.n115 7.9105
R20289 Vbias.n114 Vbias.n113 7.9105
R20290 Vbias.n112 Vbias.n111 7.9105
R20291 Vbias.n110 Vbias.n109 7.9105
R20292 Vbias.n108 Vbias.n107 7.9105
R20293 Vbias.n106 Vbias.n105 7.9105
R20294 Vbias.n104 Vbias.n103 7.9105
R20295 Vbias.n102 Vbias.n101 7.9105
R20296 Vbias.n100 Vbias.n99 7.9105
R20297 Vbias.n98 Vbias.n97 7.9105
R20298 Vbias.n94 Vbias.n93 7.9105
R20299 Vbias.n92 Vbias.n91 7.9105
R20300 Vbias.n90 Vbias.n89 7.9105
R20301 Vbias.n88 Vbias.n87 7.9105
R20302 Vbias.n86 Vbias.n85 7.9105
R20303 Vbias.n84 Vbias.n83 7.9105
R20304 Vbias.n82 Vbias.n81 7.9105
R20305 Vbias.n80 Vbias.n79 7.9105
R20306 Vbias.n78 Vbias.n77 7.9105
R20307 Vbias.n76 Vbias.n75 7.9105
R20308 Vbias.n74 Vbias.n73 7.9105
R20309 Vbias.n72 Vbias.n71 7.9105
R20310 Vbias.n70 Vbias.n69 7.9105
R20311 Vbias.n68 Vbias.n67 7.9105
R20312 Vbias.n66 Vbias.n65 7.9105
R20313 Vbias.n62 Vbias.n61 7.9105
R20314 Vbias.n60 Vbias.n59 7.9105
R20315 Vbias.n58 Vbias.n57 7.9105
R20316 Vbias.n56 Vbias.n55 7.9105
R20317 Vbias.n54 Vbias.n53 7.9105
R20318 Vbias.n52 Vbias.n51 7.9105
R20319 Vbias.n50 Vbias.n49 7.9105
R20320 Vbias.n48 Vbias.n47 7.9105
R20321 Vbias.n46 Vbias.n45 7.9105
R20322 Vbias.n44 Vbias.n43 7.9105
R20323 Vbias.n42 Vbias.n41 7.9105
R20324 Vbias.n40 Vbias.n39 7.9105
R20325 Vbias.n38 Vbias.n37 7.9105
R20326 Vbias.n36 Vbias.n35 7.9105
R20327 Vbias.n34 Vbias.n33 7.9105
R20328 Vbias.n30 Vbias.n29 7.9105
R20329 Vbias.n28 Vbias.n27 7.9105
R20330 Vbias.n26 Vbias.n25 7.9105
R20331 Vbias.n24 Vbias.n23 7.9105
R20332 Vbias.n22 Vbias.n21 7.9105
R20333 Vbias.n20 Vbias.n19 7.9105
R20334 Vbias.n18 Vbias.n17 7.9105
R20335 Vbias.n16 Vbias.n15 7.9105
R20336 Vbias.n14 Vbias.n13 7.9105
R20337 Vbias.n12 Vbias.n11 7.9105
R20338 Vbias.n10 Vbias.n9 7.9105
R20339 Vbias.n8 Vbias.n7 7.9105
R20340 Vbias.n6 Vbias.n5 7.9105
R20341 Vbias.n4 Vbias.n3 7.9105
R20342 Vbias.n2 Vbias.n1 7.9105
R20343 Vbias.n514 Vbias.n512 4.78773
R20344 Vbias.n514 Vbias.n513 4.78773
R20345 Vbias.n516 Vbias.n514 2.09636
R20346 Vbias.n511 Vbias 1.6647
R20347 Vbias.n479 Vbias 1.6647
R20348 Vbias.n447 Vbias 1.6647
R20349 Vbias.n415 Vbias 1.6647
R20350 Vbias.n383 Vbias 1.6647
R20351 Vbias.n351 Vbias 1.6647
R20352 Vbias.n319 Vbias 1.6647
R20353 Vbias.n287 Vbias 1.6647
R20354 Vbias.n255 Vbias 1.6647
R20355 Vbias.n223 Vbias 1.6647
R20356 Vbias.n191 Vbias 1.6647
R20357 Vbias.n159 Vbias 1.6647
R20358 Vbias.n127 Vbias 1.6647
R20359 Vbias.n95 Vbias 1.6647
R20360 Vbias.n63 Vbias 1.6647
R20361 Vbias.n31 Vbias 1.6647
R20362 Vbias.n517 Vbias 1.34721
R20363 Vbias Vbias.n516 0.752103
R20364 Vbias.n517 Vbias.n511 0.5692
R20365 Vbias.n516 Vbias.n515 0.515506
R20366 Vbias.n63 Vbias.n31 0.410967
R20367 Vbias.n95 Vbias.n63 0.410967
R20368 Vbias.n127 Vbias.n95 0.410967
R20369 Vbias.n159 Vbias.n127 0.410967
R20370 Vbias.n191 Vbias.n159 0.410967
R20371 Vbias.n223 Vbias.n191 0.410967
R20372 Vbias.n255 Vbias.n223 0.410967
R20373 Vbias.n287 Vbias.n255 0.410967
R20374 Vbias.n319 Vbias.n287 0.410967
R20375 Vbias.n351 Vbias.n319 0.410967
R20376 Vbias.n383 Vbias.n351 0.410967
R20377 Vbias.n415 Vbias.n383 0.410967
R20378 Vbias.n447 Vbias.n415 0.410967
R20379 Vbias.n479 Vbias.n447 0.410967
R20380 Vbias.n511 Vbias.n479 0.410967
R20381 Vbias.n31 Vbias 0.383811
R20382 Vbias.n482 Vbias 0.252372
R20383 Vbias.n484 Vbias 0.252372
R20384 Vbias.n486 Vbias 0.252372
R20385 Vbias.n488 Vbias 0.252372
R20386 Vbias.n490 Vbias 0.252372
R20387 Vbias.n492 Vbias 0.252372
R20388 Vbias.n494 Vbias 0.252372
R20389 Vbias.n496 Vbias 0.252372
R20390 Vbias.n498 Vbias 0.252372
R20391 Vbias.n500 Vbias 0.252372
R20392 Vbias.n502 Vbias 0.252372
R20393 Vbias.n504 Vbias 0.252372
R20394 Vbias.n506 Vbias 0.252372
R20395 Vbias.n508 Vbias 0.252372
R20396 Vbias.n510 Vbias 0.252372
R20397 Vbias.n450 Vbias 0.252372
R20398 Vbias.n452 Vbias 0.252372
R20399 Vbias.n454 Vbias 0.252372
R20400 Vbias.n456 Vbias 0.252372
R20401 Vbias.n458 Vbias 0.252372
R20402 Vbias.n460 Vbias 0.252372
R20403 Vbias.n462 Vbias 0.252372
R20404 Vbias.n464 Vbias 0.252372
R20405 Vbias.n466 Vbias 0.252372
R20406 Vbias.n468 Vbias 0.252372
R20407 Vbias.n470 Vbias 0.252372
R20408 Vbias.n472 Vbias 0.252372
R20409 Vbias.n474 Vbias 0.252372
R20410 Vbias.n476 Vbias 0.252372
R20411 Vbias.n478 Vbias 0.252372
R20412 Vbias.n418 Vbias 0.252372
R20413 Vbias.n420 Vbias 0.252372
R20414 Vbias.n422 Vbias 0.252372
R20415 Vbias.n424 Vbias 0.252372
R20416 Vbias.n426 Vbias 0.252372
R20417 Vbias.n428 Vbias 0.252372
R20418 Vbias.n430 Vbias 0.252372
R20419 Vbias.n432 Vbias 0.252372
R20420 Vbias.n434 Vbias 0.252372
R20421 Vbias.n436 Vbias 0.252372
R20422 Vbias.n438 Vbias 0.252372
R20423 Vbias.n440 Vbias 0.252372
R20424 Vbias.n442 Vbias 0.252372
R20425 Vbias.n444 Vbias 0.252372
R20426 Vbias.n446 Vbias 0.252372
R20427 Vbias.n386 Vbias 0.252372
R20428 Vbias.n388 Vbias 0.252372
R20429 Vbias.n390 Vbias 0.252372
R20430 Vbias.n392 Vbias 0.252372
R20431 Vbias.n394 Vbias 0.252372
R20432 Vbias.n396 Vbias 0.252372
R20433 Vbias.n398 Vbias 0.252372
R20434 Vbias.n400 Vbias 0.252372
R20435 Vbias.n402 Vbias 0.252372
R20436 Vbias.n404 Vbias 0.252372
R20437 Vbias.n406 Vbias 0.252372
R20438 Vbias.n408 Vbias 0.252372
R20439 Vbias.n410 Vbias 0.252372
R20440 Vbias.n412 Vbias 0.252372
R20441 Vbias.n414 Vbias 0.252372
R20442 Vbias.n354 Vbias 0.252372
R20443 Vbias.n356 Vbias 0.252372
R20444 Vbias.n358 Vbias 0.252372
R20445 Vbias.n360 Vbias 0.252372
R20446 Vbias.n362 Vbias 0.252372
R20447 Vbias.n364 Vbias 0.252372
R20448 Vbias.n366 Vbias 0.252372
R20449 Vbias.n368 Vbias 0.252372
R20450 Vbias.n370 Vbias 0.252372
R20451 Vbias.n372 Vbias 0.252372
R20452 Vbias.n374 Vbias 0.252372
R20453 Vbias.n376 Vbias 0.252372
R20454 Vbias.n378 Vbias 0.252372
R20455 Vbias.n380 Vbias 0.252372
R20456 Vbias.n382 Vbias 0.252372
R20457 Vbias.n322 Vbias 0.252372
R20458 Vbias.n324 Vbias 0.252372
R20459 Vbias.n326 Vbias 0.252372
R20460 Vbias.n328 Vbias 0.252372
R20461 Vbias.n330 Vbias 0.252372
R20462 Vbias.n332 Vbias 0.252372
R20463 Vbias.n334 Vbias 0.252372
R20464 Vbias.n336 Vbias 0.252372
R20465 Vbias.n338 Vbias 0.252372
R20466 Vbias.n340 Vbias 0.252372
R20467 Vbias.n342 Vbias 0.252372
R20468 Vbias.n344 Vbias 0.252372
R20469 Vbias.n346 Vbias 0.252372
R20470 Vbias.n348 Vbias 0.252372
R20471 Vbias.n350 Vbias 0.252372
R20472 Vbias.n290 Vbias 0.252372
R20473 Vbias.n292 Vbias 0.252372
R20474 Vbias.n294 Vbias 0.252372
R20475 Vbias.n296 Vbias 0.252372
R20476 Vbias.n298 Vbias 0.252372
R20477 Vbias.n300 Vbias 0.252372
R20478 Vbias.n302 Vbias 0.252372
R20479 Vbias.n304 Vbias 0.252372
R20480 Vbias.n306 Vbias 0.252372
R20481 Vbias.n308 Vbias 0.252372
R20482 Vbias.n310 Vbias 0.252372
R20483 Vbias.n312 Vbias 0.252372
R20484 Vbias.n314 Vbias 0.252372
R20485 Vbias.n316 Vbias 0.252372
R20486 Vbias.n318 Vbias 0.252372
R20487 Vbias.n258 Vbias 0.252372
R20488 Vbias.n260 Vbias 0.252372
R20489 Vbias.n262 Vbias 0.252372
R20490 Vbias.n264 Vbias 0.252372
R20491 Vbias.n266 Vbias 0.252372
R20492 Vbias.n268 Vbias 0.252372
R20493 Vbias.n270 Vbias 0.252372
R20494 Vbias.n272 Vbias 0.252372
R20495 Vbias.n274 Vbias 0.252372
R20496 Vbias.n276 Vbias 0.252372
R20497 Vbias.n278 Vbias 0.252372
R20498 Vbias.n280 Vbias 0.252372
R20499 Vbias.n282 Vbias 0.252372
R20500 Vbias.n284 Vbias 0.252372
R20501 Vbias.n286 Vbias 0.252372
R20502 Vbias.n226 Vbias 0.252372
R20503 Vbias.n228 Vbias 0.252372
R20504 Vbias.n230 Vbias 0.252372
R20505 Vbias.n232 Vbias 0.252372
R20506 Vbias.n234 Vbias 0.252372
R20507 Vbias.n236 Vbias 0.252372
R20508 Vbias.n238 Vbias 0.252372
R20509 Vbias.n240 Vbias 0.252372
R20510 Vbias.n242 Vbias 0.252372
R20511 Vbias.n244 Vbias 0.252372
R20512 Vbias.n246 Vbias 0.252372
R20513 Vbias.n248 Vbias 0.252372
R20514 Vbias.n250 Vbias 0.252372
R20515 Vbias.n252 Vbias 0.252372
R20516 Vbias.n254 Vbias 0.252372
R20517 Vbias.n194 Vbias 0.252372
R20518 Vbias.n196 Vbias 0.252372
R20519 Vbias.n198 Vbias 0.252372
R20520 Vbias.n200 Vbias 0.252372
R20521 Vbias.n202 Vbias 0.252372
R20522 Vbias.n204 Vbias 0.252372
R20523 Vbias.n206 Vbias 0.252372
R20524 Vbias.n208 Vbias 0.252372
R20525 Vbias.n210 Vbias 0.252372
R20526 Vbias.n212 Vbias 0.252372
R20527 Vbias.n214 Vbias 0.252372
R20528 Vbias.n216 Vbias 0.252372
R20529 Vbias.n218 Vbias 0.252372
R20530 Vbias.n220 Vbias 0.252372
R20531 Vbias.n222 Vbias 0.252372
R20532 Vbias.n162 Vbias 0.252372
R20533 Vbias.n164 Vbias 0.252372
R20534 Vbias.n166 Vbias 0.252372
R20535 Vbias.n168 Vbias 0.252372
R20536 Vbias.n170 Vbias 0.252372
R20537 Vbias.n172 Vbias 0.252372
R20538 Vbias.n174 Vbias 0.252372
R20539 Vbias.n176 Vbias 0.252372
R20540 Vbias.n178 Vbias 0.252372
R20541 Vbias.n180 Vbias 0.252372
R20542 Vbias.n182 Vbias 0.252372
R20543 Vbias.n184 Vbias 0.252372
R20544 Vbias.n186 Vbias 0.252372
R20545 Vbias.n188 Vbias 0.252372
R20546 Vbias.n190 Vbias 0.252372
R20547 Vbias.n130 Vbias 0.252372
R20548 Vbias.n132 Vbias 0.252372
R20549 Vbias.n134 Vbias 0.252372
R20550 Vbias.n136 Vbias 0.252372
R20551 Vbias.n138 Vbias 0.252372
R20552 Vbias.n140 Vbias 0.252372
R20553 Vbias.n142 Vbias 0.252372
R20554 Vbias.n144 Vbias 0.252372
R20555 Vbias.n146 Vbias 0.252372
R20556 Vbias.n148 Vbias 0.252372
R20557 Vbias.n150 Vbias 0.252372
R20558 Vbias.n152 Vbias 0.252372
R20559 Vbias.n154 Vbias 0.252372
R20560 Vbias.n156 Vbias 0.252372
R20561 Vbias.n158 Vbias 0.252372
R20562 Vbias.n98 Vbias 0.252372
R20563 Vbias.n100 Vbias 0.252372
R20564 Vbias.n102 Vbias 0.252372
R20565 Vbias.n104 Vbias 0.252372
R20566 Vbias.n106 Vbias 0.252372
R20567 Vbias.n108 Vbias 0.252372
R20568 Vbias.n110 Vbias 0.252372
R20569 Vbias.n112 Vbias 0.252372
R20570 Vbias.n114 Vbias 0.252372
R20571 Vbias.n116 Vbias 0.252372
R20572 Vbias.n118 Vbias 0.252372
R20573 Vbias.n120 Vbias 0.252372
R20574 Vbias.n122 Vbias 0.252372
R20575 Vbias.n124 Vbias 0.252372
R20576 Vbias.n126 Vbias 0.252372
R20577 Vbias.n66 Vbias 0.252372
R20578 Vbias.n68 Vbias 0.252372
R20579 Vbias.n70 Vbias 0.252372
R20580 Vbias.n72 Vbias 0.252372
R20581 Vbias.n74 Vbias 0.252372
R20582 Vbias.n76 Vbias 0.252372
R20583 Vbias.n78 Vbias 0.252372
R20584 Vbias.n80 Vbias 0.252372
R20585 Vbias.n82 Vbias 0.252372
R20586 Vbias.n84 Vbias 0.252372
R20587 Vbias.n86 Vbias 0.252372
R20588 Vbias.n88 Vbias 0.252372
R20589 Vbias.n90 Vbias 0.252372
R20590 Vbias.n92 Vbias 0.252372
R20591 Vbias.n94 Vbias 0.252372
R20592 Vbias.n34 Vbias 0.252372
R20593 Vbias.n36 Vbias 0.252372
R20594 Vbias.n38 Vbias 0.252372
R20595 Vbias.n40 Vbias 0.252372
R20596 Vbias.n42 Vbias 0.252372
R20597 Vbias.n44 Vbias 0.252372
R20598 Vbias.n46 Vbias 0.252372
R20599 Vbias.n48 Vbias 0.252372
R20600 Vbias.n50 Vbias 0.252372
R20601 Vbias.n52 Vbias 0.252372
R20602 Vbias.n54 Vbias 0.252372
R20603 Vbias.n56 Vbias 0.252372
R20604 Vbias.n58 Vbias 0.252372
R20605 Vbias.n60 Vbias 0.252372
R20606 Vbias.n62 Vbias 0.252372
R20607 Vbias.n2 Vbias 0.252372
R20608 Vbias.n4 Vbias 0.252372
R20609 Vbias.n6 Vbias 0.252372
R20610 Vbias.n8 Vbias 0.252372
R20611 Vbias.n10 Vbias 0.252372
R20612 Vbias.n12 Vbias 0.252372
R20613 Vbias.n14 Vbias 0.252372
R20614 Vbias.n16 Vbias 0.252372
R20615 Vbias.n18 Vbias 0.252372
R20616 Vbias.n20 Vbias 0.252372
R20617 Vbias.n22 Vbias 0.252372
R20618 Vbias.n24 Vbias 0.252372
R20619 Vbias.n26 Vbias 0.252372
R20620 Vbias.n28 Vbias 0.252372
R20621 Vbias.n30 Vbias 0.252372
R20622 Vbias Vbias.n517 0.237067
R20623 Vbias Vbias.n482 0.0972718
R20624 Vbias Vbias.n484 0.0972718
R20625 Vbias Vbias.n486 0.0972718
R20626 Vbias Vbias.n488 0.0972718
R20627 Vbias Vbias.n490 0.0972718
R20628 Vbias Vbias.n492 0.0972718
R20629 Vbias Vbias.n494 0.0972718
R20630 Vbias Vbias.n496 0.0972718
R20631 Vbias Vbias.n498 0.0972718
R20632 Vbias Vbias.n500 0.0972718
R20633 Vbias Vbias.n502 0.0972718
R20634 Vbias Vbias.n504 0.0972718
R20635 Vbias Vbias.n506 0.0972718
R20636 Vbias Vbias.n508 0.0972718
R20637 Vbias Vbias.n510 0.0972718
R20638 Vbias Vbias.n450 0.0972718
R20639 Vbias Vbias.n452 0.0972718
R20640 Vbias Vbias.n454 0.0972718
R20641 Vbias Vbias.n456 0.0972718
R20642 Vbias Vbias.n458 0.0972718
R20643 Vbias Vbias.n460 0.0972718
R20644 Vbias Vbias.n462 0.0972718
R20645 Vbias Vbias.n464 0.0972718
R20646 Vbias Vbias.n466 0.0972718
R20647 Vbias Vbias.n468 0.0972718
R20648 Vbias Vbias.n470 0.0972718
R20649 Vbias Vbias.n472 0.0972718
R20650 Vbias Vbias.n474 0.0972718
R20651 Vbias Vbias.n476 0.0972718
R20652 Vbias Vbias.n478 0.0972718
R20653 Vbias Vbias.n418 0.0972718
R20654 Vbias Vbias.n420 0.0972718
R20655 Vbias Vbias.n422 0.0972718
R20656 Vbias Vbias.n424 0.0972718
R20657 Vbias Vbias.n426 0.0972718
R20658 Vbias Vbias.n428 0.0972718
R20659 Vbias Vbias.n430 0.0972718
R20660 Vbias Vbias.n432 0.0972718
R20661 Vbias Vbias.n434 0.0972718
R20662 Vbias Vbias.n436 0.0972718
R20663 Vbias Vbias.n438 0.0972718
R20664 Vbias Vbias.n440 0.0972718
R20665 Vbias Vbias.n442 0.0972718
R20666 Vbias Vbias.n444 0.0972718
R20667 Vbias Vbias.n446 0.0972718
R20668 Vbias Vbias.n386 0.0972718
R20669 Vbias Vbias.n388 0.0972718
R20670 Vbias Vbias.n390 0.0972718
R20671 Vbias Vbias.n392 0.0972718
R20672 Vbias Vbias.n394 0.0972718
R20673 Vbias Vbias.n396 0.0972718
R20674 Vbias Vbias.n398 0.0972718
R20675 Vbias Vbias.n400 0.0972718
R20676 Vbias Vbias.n402 0.0972718
R20677 Vbias Vbias.n404 0.0972718
R20678 Vbias Vbias.n406 0.0972718
R20679 Vbias Vbias.n408 0.0972718
R20680 Vbias Vbias.n410 0.0972718
R20681 Vbias Vbias.n412 0.0972718
R20682 Vbias Vbias.n414 0.0972718
R20683 Vbias Vbias.n354 0.0972718
R20684 Vbias Vbias.n356 0.0972718
R20685 Vbias Vbias.n358 0.0972718
R20686 Vbias Vbias.n360 0.0972718
R20687 Vbias Vbias.n362 0.0972718
R20688 Vbias Vbias.n364 0.0972718
R20689 Vbias Vbias.n366 0.0972718
R20690 Vbias Vbias.n368 0.0972718
R20691 Vbias Vbias.n370 0.0972718
R20692 Vbias Vbias.n372 0.0972718
R20693 Vbias Vbias.n374 0.0972718
R20694 Vbias Vbias.n376 0.0972718
R20695 Vbias Vbias.n378 0.0972718
R20696 Vbias Vbias.n380 0.0972718
R20697 Vbias Vbias.n382 0.0972718
R20698 Vbias Vbias.n322 0.0972718
R20699 Vbias Vbias.n324 0.0972718
R20700 Vbias Vbias.n326 0.0972718
R20701 Vbias Vbias.n328 0.0972718
R20702 Vbias Vbias.n330 0.0972718
R20703 Vbias Vbias.n332 0.0972718
R20704 Vbias Vbias.n334 0.0972718
R20705 Vbias Vbias.n336 0.0972718
R20706 Vbias Vbias.n338 0.0972718
R20707 Vbias Vbias.n340 0.0972718
R20708 Vbias Vbias.n342 0.0972718
R20709 Vbias Vbias.n344 0.0972718
R20710 Vbias Vbias.n346 0.0972718
R20711 Vbias Vbias.n348 0.0972718
R20712 Vbias Vbias.n350 0.0972718
R20713 Vbias Vbias.n290 0.0972718
R20714 Vbias Vbias.n292 0.0972718
R20715 Vbias Vbias.n294 0.0972718
R20716 Vbias Vbias.n296 0.0972718
R20717 Vbias Vbias.n298 0.0972718
R20718 Vbias Vbias.n300 0.0972718
R20719 Vbias Vbias.n302 0.0972718
R20720 Vbias Vbias.n304 0.0972718
R20721 Vbias Vbias.n306 0.0972718
R20722 Vbias Vbias.n308 0.0972718
R20723 Vbias Vbias.n310 0.0972718
R20724 Vbias Vbias.n312 0.0972718
R20725 Vbias Vbias.n314 0.0972718
R20726 Vbias Vbias.n316 0.0972718
R20727 Vbias Vbias.n318 0.0972718
R20728 Vbias Vbias.n258 0.0972718
R20729 Vbias Vbias.n260 0.0972718
R20730 Vbias Vbias.n262 0.0972718
R20731 Vbias Vbias.n264 0.0972718
R20732 Vbias Vbias.n266 0.0972718
R20733 Vbias Vbias.n268 0.0972718
R20734 Vbias Vbias.n270 0.0972718
R20735 Vbias Vbias.n272 0.0972718
R20736 Vbias Vbias.n274 0.0972718
R20737 Vbias Vbias.n276 0.0972718
R20738 Vbias Vbias.n278 0.0972718
R20739 Vbias Vbias.n280 0.0972718
R20740 Vbias Vbias.n282 0.0972718
R20741 Vbias Vbias.n284 0.0972718
R20742 Vbias Vbias.n286 0.0972718
R20743 Vbias Vbias.n226 0.0972718
R20744 Vbias Vbias.n228 0.0972718
R20745 Vbias Vbias.n230 0.0972718
R20746 Vbias Vbias.n232 0.0972718
R20747 Vbias Vbias.n234 0.0972718
R20748 Vbias Vbias.n236 0.0972718
R20749 Vbias Vbias.n238 0.0972718
R20750 Vbias Vbias.n240 0.0972718
R20751 Vbias Vbias.n242 0.0972718
R20752 Vbias Vbias.n244 0.0972718
R20753 Vbias Vbias.n246 0.0972718
R20754 Vbias Vbias.n248 0.0972718
R20755 Vbias Vbias.n250 0.0972718
R20756 Vbias Vbias.n252 0.0972718
R20757 Vbias Vbias.n254 0.0972718
R20758 Vbias Vbias.n194 0.0972718
R20759 Vbias Vbias.n196 0.0972718
R20760 Vbias Vbias.n198 0.0972718
R20761 Vbias Vbias.n200 0.0972718
R20762 Vbias Vbias.n202 0.0972718
R20763 Vbias Vbias.n204 0.0972718
R20764 Vbias Vbias.n206 0.0972718
R20765 Vbias Vbias.n208 0.0972718
R20766 Vbias Vbias.n210 0.0972718
R20767 Vbias Vbias.n212 0.0972718
R20768 Vbias Vbias.n214 0.0972718
R20769 Vbias Vbias.n216 0.0972718
R20770 Vbias Vbias.n218 0.0972718
R20771 Vbias Vbias.n220 0.0972718
R20772 Vbias Vbias.n222 0.0972718
R20773 Vbias Vbias.n162 0.0972718
R20774 Vbias Vbias.n164 0.0972718
R20775 Vbias Vbias.n166 0.0972718
R20776 Vbias Vbias.n168 0.0972718
R20777 Vbias Vbias.n170 0.0972718
R20778 Vbias Vbias.n172 0.0972718
R20779 Vbias Vbias.n174 0.0972718
R20780 Vbias Vbias.n176 0.0972718
R20781 Vbias Vbias.n178 0.0972718
R20782 Vbias Vbias.n180 0.0972718
R20783 Vbias Vbias.n182 0.0972718
R20784 Vbias Vbias.n184 0.0972718
R20785 Vbias Vbias.n186 0.0972718
R20786 Vbias Vbias.n188 0.0972718
R20787 Vbias Vbias.n190 0.0972718
R20788 Vbias Vbias.n130 0.0972718
R20789 Vbias Vbias.n132 0.0972718
R20790 Vbias Vbias.n134 0.0972718
R20791 Vbias Vbias.n136 0.0972718
R20792 Vbias Vbias.n138 0.0972718
R20793 Vbias Vbias.n140 0.0972718
R20794 Vbias Vbias.n142 0.0972718
R20795 Vbias Vbias.n144 0.0972718
R20796 Vbias Vbias.n146 0.0972718
R20797 Vbias Vbias.n148 0.0972718
R20798 Vbias Vbias.n150 0.0972718
R20799 Vbias Vbias.n152 0.0972718
R20800 Vbias Vbias.n154 0.0972718
R20801 Vbias Vbias.n156 0.0972718
R20802 Vbias Vbias.n158 0.0972718
R20803 Vbias Vbias.n98 0.0972718
R20804 Vbias Vbias.n100 0.0972718
R20805 Vbias Vbias.n102 0.0972718
R20806 Vbias Vbias.n104 0.0972718
R20807 Vbias Vbias.n106 0.0972718
R20808 Vbias Vbias.n108 0.0972718
R20809 Vbias Vbias.n110 0.0972718
R20810 Vbias Vbias.n112 0.0972718
R20811 Vbias Vbias.n114 0.0972718
R20812 Vbias Vbias.n116 0.0972718
R20813 Vbias Vbias.n118 0.0972718
R20814 Vbias Vbias.n120 0.0972718
R20815 Vbias Vbias.n122 0.0972718
R20816 Vbias Vbias.n124 0.0972718
R20817 Vbias Vbias.n126 0.0972718
R20818 Vbias Vbias.n66 0.0972718
R20819 Vbias Vbias.n68 0.0972718
R20820 Vbias Vbias.n70 0.0972718
R20821 Vbias Vbias.n72 0.0972718
R20822 Vbias Vbias.n74 0.0972718
R20823 Vbias Vbias.n76 0.0972718
R20824 Vbias Vbias.n78 0.0972718
R20825 Vbias Vbias.n80 0.0972718
R20826 Vbias Vbias.n82 0.0972718
R20827 Vbias Vbias.n84 0.0972718
R20828 Vbias Vbias.n86 0.0972718
R20829 Vbias Vbias.n88 0.0972718
R20830 Vbias Vbias.n90 0.0972718
R20831 Vbias Vbias.n92 0.0972718
R20832 Vbias Vbias.n94 0.0972718
R20833 Vbias Vbias.n34 0.0972718
R20834 Vbias Vbias.n36 0.0972718
R20835 Vbias Vbias.n38 0.0972718
R20836 Vbias Vbias.n40 0.0972718
R20837 Vbias Vbias.n42 0.0972718
R20838 Vbias Vbias.n44 0.0972718
R20839 Vbias Vbias.n46 0.0972718
R20840 Vbias Vbias.n48 0.0972718
R20841 Vbias Vbias.n50 0.0972718
R20842 Vbias Vbias.n52 0.0972718
R20843 Vbias Vbias.n54 0.0972718
R20844 Vbias Vbias.n56 0.0972718
R20845 Vbias Vbias.n58 0.0972718
R20846 Vbias Vbias.n60 0.0972718
R20847 Vbias Vbias.n62 0.0972718
R20848 Vbias Vbias.n2 0.0972718
R20849 Vbias Vbias.n4 0.0972718
R20850 Vbias Vbias.n6 0.0972718
R20851 Vbias Vbias.n8 0.0972718
R20852 Vbias Vbias.n10 0.0972718
R20853 Vbias Vbias.n12 0.0972718
R20854 Vbias Vbias.n14 0.0972718
R20855 Vbias Vbias.n16 0.0972718
R20856 Vbias Vbias.n18 0.0972718
R20857 Vbias Vbias.n20 0.0972718
R20858 Vbias Vbias.n22 0.0972718
R20859 Vbias Vbias.n24 0.0972718
R20860 Vbias Vbias.n26 0.0972718
R20861 Vbias Vbias.n28 0.0972718
R20862 Vbias Vbias.n30 0.0972718
R20863 Vbias.n509 Vbias 0.0489375
R20864 Vbias.n507 Vbias 0.0489375
R20865 Vbias.n505 Vbias 0.0489375
R20866 Vbias.n503 Vbias 0.0489375
R20867 Vbias.n501 Vbias 0.0489375
R20868 Vbias.n499 Vbias 0.0489375
R20869 Vbias.n497 Vbias 0.0489375
R20870 Vbias.n495 Vbias 0.0489375
R20871 Vbias.n493 Vbias 0.0489375
R20872 Vbias.n491 Vbias 0.0489375
R20873 Vbias.n489 Vbias 0.0489375
R20874 Vbias.n487 Vbias 0.0489375
R20875 Vbias.n485 Vbias 0.0489375
R20876 Vbias.n483 Vbias 0.0489375
R20877 Vbias.n481 Vbias 0.0489375
R20878 Vbias.n480 Vbias 0.0489375
R20879 Vbias.n477 Vbias 0.0489375
R20880 Vbias.n475 Vbias 0.0489375
R20881 Vbias.n473 Vbias 0.0489375
R20882 Vbias.n471 Vbias 0.0489375
R20883 Vbias.n469 Vbias 0.0489375
R20884 Vbias.n467 Vbias 0.0489375
R20885 Vbias.n465 Vbias 0.0489375
R20886 Vbias.n463 Vbias 0.0489375
R20887 Vbias.n461 Vbias 0.0489375
R20888 Vbias.n459 Vbias 0.0489375
R20889 Vbias.n457 Vbias 0.0489375
R20890 Vbias.n455 Vbias 0.0489375
R20891 Vbias.n453 Vbias 0.0489375
R20892 Vbias.n451 Vbias 0.0489375
R20893 Vbias.n449 Vbias 0.0489375
R20894 Vbias.n448 Vbias 0.0489375
R20895 Vbias.n445 Vbias 0.0489375
R20896 Vbias.n443 Vbias 0.0489375
R20897 Vbias.n441 Vbias 0.0489375
R20898 Vbias.n439 Vbias 0.0489375
R20899 Vbias.n437 Vbias 0.0489375
R20900 Vbias.n435 Vbias 0.0489375
R20901 Vbias.n433 Vbias 0.0489375
R20902 Vbias.n431 Vbias 0.0489375
R20903 Vbias.n429 Vbias 0.0489375
R20904 Vbias.n427 Vbias 0.0489375
R20905 Vbias.n425 Vbias 0.0489375
R20906 Vbias.n423 Vbias 0.0489375
R20907 Vbias.n421 Vbias 0.0489375
R20908 Vbias.n419 Vbias 0.0489375
R20909 Vbias.n417 Vbias 0.0489375
R20910 Vbias.n416 Vbias 0.0489375
R20911 Vbias.n413 Vbias 0.0489375
R20912 Vbias.n411 Vbias 0.0489375
R20913 Vbias.n409 Vbias 0.0489375
R20914 Vbias.n407 Vbias 0.0489375
R20915 Vbias.n405 Vbias 0.0489375
R20916 Vbias.n403 Vbias 0.0489375
R20917 Vbias.n401 Vbias 0.0489375
R20918 Vbias.n399 Vbias 0.0489375
R20919 Vbias.n397 Vbias 0.0489375
R20920 Vbias.n395 Vbias 0.0489375
R20921 Vbias.n393 Vbias 0.0489375
R20922 Vbias.n391 Vbias 0.0489375
R20923 Vbias.n389 Vbias 0.0489375
R20924 Vbias.n387 Vbias 0.0489375
R20925 Vbias.n385 Vbias 0.0489375
R20926 Vbias.n384 Vbias 0.0489375
R20927 Vbias.n381 Vbias 0.0489375
R20928 Vbias.n379 Vbias 0.0489375
R20929 Vbias.n377 Vbias 0.0489375
R20930 Vbias.n375 Vbias 0.0489375
R20931 Vbias.n373 Vbias 0.0489375
R20932 Vbias.n371 Vbias 0.0489375
R20933 Vbias.n369 Vbias 0.0489375
R20934 Vbias.n367 Vbias 0.0489375
R20935 Vbias.n365 Vbias 0.0489375
R20936 Vbias.n363 Vbias 0.0489375
R20937 Vbias.n361 Vbias 0.0489375
R20938 Vbias.n359 Vbias 0.0489375
R20939 Vbias.n357 Vbias 0.0489375
R20940 Vbias.n355 Vbias 0.0489375
R20941 Vbias.n353 Vbias 0.0489375
R20942 Vbias.n352 Vbias 0.0489375
R20943 Vbias.n349 Vbias 0.0489375
R20944 Vbias.n347 Vbias 0.0489375
R20945 Vbias.n345 Vbias 0.0489375
R20946 Vbias.n343 Vbias 0.0489375
R20947 Vbias.n341 Vbias 0.0489375
R20948 Vbias.n339 Vbias 0.0489375
R20949 Vbias.n337 Vbias 0.0489375
R20950 Vbias.n335 Vbias 0.0489375
R20951 Vbias.n333 Vbias 0.0489375
R20952 Vbias.n331 Vbias 0.0489375
R20953 Vbias.n329 Vbias 0.0489375
R20954 Vbias.n327 Vbias 0.0489375
R20955 Vbias.n325 Vbias 0.0489375
R20956 Vbias.n323 Vbias 0.0489375
R20957 Vbias.n321 Vbias 0.0489375
R20958 Vbias.n320 Vbias 0.0489375
R20959 Vbias.n317 Vbias 0.0489375
R20960 Vbias.n315 Vbias 0.0489375
R20961 Vbias.n313 Vbias 0.0489375
R20962 Vbias.n311 Vbias 0.0489375
R20963 Vbias.n309 Vbias 0.0489375
R20964 Vbias.n307 Vbias 0.0489375
R20965 Vbias.n305 Vbias 0.0489375
R20966 Vbias.n303 Vbias 0.0489375
R20967 Vbias.n301 Vbias 0.0489375
R20968 Vbias.n299 Vbias 0.0489375
R20969 Vbias.n297 Vbias 0.0489375
R20970 Vbias.n295 Vbias 0.0489375
R20971 Vbias.n293 Vbias 0.0489375
R20972 Vbias.n291 Vbias 0.0489375
R20973 Vbias.n289 Vbias 0.0489375
R20974 Vbias.n288 Vbias 0.0489375
R20975 Vbias.n285 Vbias 0.0489375
R20976 Vbias.n283 Vbias 0.0489375
R20977 Vbias.n281 Vbias 0.0489375
R20978 Vbias.n279 Vbias 0.0489375
R20979 Vbias.n277 Vbias 0.0489375
R20980 Vbias.n275 Vbias 0.0489375
R20981 Vbias.n273 Vbias 0.0489375
R20982 Vbias.n271 Vbias 0.0489375
R20983 Vbias.n269 Vbias 0.0489375
R20984 Vbias.n267 Vbias 0.0489375
R20985 Vbias.n265 Vbias 0.0489375
R20986 Vbias.n263 Vbias 0.0489375
R20987 Vbias.n261 Vbias 0.0489375
R20988 Vbias.n259 Vbias 0.0489375
R20989 Vbias.n257 Vbias 0.0489375
R20990 Vbias.n256 Vbias 0.0489375
R20991 Vbias.n253 Vbias 0.0489375
R20992 Vbias.n251 Vbias 0.0489375
R20993 Vbias.n249 Vbias 0.0489375
R20994 Vbias.n247 Vbias 0.0489375
R20995 Vbias.n245 Vbias 0.0489375
R20996 Vbias.n243 Vbias 0.0489375
R20997 Vbias.n241 Vbias 0.0489375
R20998 Vbias.n239 Vbias 0.0489375
R20999 Vbias.n237 Vbias 0.0489375
R21000 Vbias.n235 Vbias 0.0489375
R21001 Vbias.n233 Vbias 0.0489375
R21002 Vbias.n231 Vbias 0.0489375
R21003 Vbias.n229 Vbias 0.0489375
R21004 Vbias.n227 Vbias 0.0489375
R21005 Vbias.n225 Vbias 0.0489375
R21006 Vbias.n224 Vbias 0.0489375
R21007 Vbias.n221 Vbias 0.0489375
R21008 Vbias.n219 Vbias 0.0489375
R21009 Vbias.n217 Vbias 0.0489375
R21010 Vbias.n215 Vbias 0.0489375
R21011 Vbias.n213 Vbias 0.0489375
R21012 Vbias.n211 Vbias 0.0489375
R21013 Vbias.n209 Vbias 0.0489375
R21014 Vbias.n207 Vbias 0.0489375
R21015 Vbias.n205 Vbias 0.0489375
R21016 Vbias.n203 Vbias 0.0489375
R21017 Vbias.n201 Vbias 0.0489375
R21018 Vbias.n199 Vbias 0.0489375
R21019 Vbias.n197 Vbias 0.0489375
R21020 Vbias.n195 Vbias 0.0489375
R21021 Vbias.n193 Vbias 0.0489375
R21022 Vbias.n192 Vbias 0.0489375
R21023 Vbias.n189 Vbias 0.0489375
R21024 Vbias.n187 Vbias 0.0489375
R21025 Vbias.n185 Vbias 0.0489375
R21026 Vbias.n183 Vbias 0.0489375
R21027 Vbias.n181 Vbias 0.0489375
R21028 Vbias.n179 Vbias 0.0489375
R21029 Vbias.n177 Vbias 0.0489375
R21030 Vbias.n175 Vbias 0.0489375
R21031 Vbias.n173 Vbias 0.0489375
R21032 Vbias.n171 Vbias 0.0489375
R21033 Vbias.n169 Vbias 0.0489375
R21034 Vbias.n167 Vbias 0.0489375
R21035 Vbias.n165 Vbias 0.0489375
R21036 Vbias.n163 Vbias 0.0489375
R21037 Vbias.n161 Vbias 0.0489375
R21038 Vbias.n160 Vbias 0.0489375
R21039 Vbias.n157 Vbias 0.0489375
R21040 Vbias.n155 Vbias 0.0489375
R21041 Vbias.n153 Vbias 0.0489375
R21042 Vbias.n151 Vbias 0.0489375
R21043 Vbias.n149 Vbias 0.0489375
R21044 Vbias.n147 Vbias 0.0489375
R21045 Vbias.n145 Vbias 0.0489375
R21046 Vbias.n143 Vbias 0.0489375
R21047 Vbias.n141 Vbias 0.0489375
R21048 Vbias.n139 Vbias 0.0489375
R21049 Vbias.n137 Vbias 0.0489375
R21050 Vbias.n135 Vbias 0.0489375
R21051 Vbias.n133 Vbias 0.0489375
R21052 Vbias.n131 Vbias 0.0489375
R21053 Vbias.n129 Vbias 0.0489375
R21054 Vbias.n128 Vbias 0.0489375
R21055 Vbias.n125 Vbias 0.0489375
R21056 Vbias.n123 Vbias 0.0489375
R21057 Vbias.n121 Vbias 0.0489375
R21058 Vbias.n119 Vbias 0.0489375
R21059 Vbias.n117 Vbias 0.0489375
R21060 Vbias.n115 Vbias 0.0489375
R21061 Vbias.n113 Vbias 0.0489375
R21062 Vbias.n111 Vbias 0.0489375
R21063 Vbias.n109 Vbias 0.0489375
R21064 Vbias.n107 Vbias 0.0489375
R21065 Vbias.n105 Vbias 0.0489375
R21066 Vbias.n103 Vbias 0.0489375
R21067 Vbias.n101 Vbias 0.0489375
R21068 Vbias.n99 Vbias 0.0489375
R21069 Vbias.n97 Vbias 0.0489375
R21070 Vbias.n96 Vbias 0.0489375
R21071 Vbias.n93 Vbias 0.0489375
R21072 Vbias.n91 Vbias 0.0489375
R21073 Vbias.n89 Vbias 0.0489375
R21074 Vbias.n87 Vbias 0.0489375
R21075 Vbias.n85 Vbias 0.0489375
R21076 Vbias.n83 Vbias 0.0489375
R21077 Vbias.n81 Vbias 0.0489375
R21078 Vbias.n79 Vbias 0.0489375
R21079 Vbias.n77 Vbias 0.0489375
R21080 Vbias.n75 Vbias 0.0489375
R21081 Vbias.n73 Vbias 0.0489375
R21082 Vbias.n71 Vbias 0.0489375
R21083 Vbias.n69 Vbias 0.0489375
R21084 Vbias.n67 Vbias 0.0489375
R21085 Vbias.n65 Vbias 0.0489375
R21086 Vbias.n64 Vbias 0.0489375
R21087 Vbias.n61 Vbias 0.0489375
R21088 Vbias.n59 Vbias 0.0489375
R21089 Vbias.n57 Vbias 0.0489375
R21090 Vbias.n55 Vbias 0.0489375
R21091 Vbias.n53 Vbias 0.0489375
R21092 Vbias.n51 Vbias 0.0489375
R21093 Vbias.n49 Vbias 0.0489375
R21094 Vbias.n47 Vbias 0.0489375
R21095 Vbias.n45 Vbias 0.0489375
R21096 Vbias.n43 Vbias 0.0489375
R21097 Vbias.n41 Vbias 0.0489375
R21098 Vbias.n39 Vbias 0.0489375
R21099 Vbias.n37 Vbias 0.0489375
R21100 Vbias.n35 Vbias 0.0489375
R21101 Vbias.n33 Vbias 0.0489375
R21102 Vbias.n32 Vbias 0.0489375
R21103 Vbias.n29 Vbias 0.0489375
R21104 Vbias.n27 Vbias 0.0489375
R21105 Vbias.n25 Vbias 0.0489375
R21106 Vbias.n23 Vbias 0.0489375
R21107 Vbias.n21 Vbias 0.0489375
R21108 Vbias.n19 Vbias 0.0489375
R21109 Vbias.n17 Vbias 0.0489375
R21110 Vbias.n15 Vbias 0.0489375
R21111 Vbias.n13 Vbias 0.0489375
R21112 Vbias.n11 Vbias 0.0489375
R21113 Vbias.n9 Vbias 0.0489375
R21114 Vbias.n7 Vbias 0.0489375
R21115 Vbias.n5 Vbias 0.0489375
R21116 Vbias.n3 Vbias 0.0489375
R21117 Vbias.n1 Vbias 0.0489375
R21118 Vbias.n0 Vbias 0.0489375
R21119 XA.Cn[1].n2 XA.Cn[1].n1 332.332
R21120 XA.Cn[1].n2 XA.Cn[1].n0 296.493
R21121 XA.Cn[1].n12 XA.Cn[1].n10 161.406
R21122 XA.Cn[1].n15 XA.Cn[1].n13 161.406
R21123 XA.Cn[1].n18 XA.Cn[1].n16 161.406
R21124 XA.Cn[1].n21 XA.Cn[1].n19 161.406
R21125 XA.Cn[1].n24 XA.Cn[1].n22 161.406
R21126 XA.Cn[1].n27 XA.Cn[1].n25 161.406
R21127 XA.Cn[1].n30 XA.Cn[1].n28 161.406
R21128 XA.Cn[1].n33 XA.Cn[1].n31 161.406
R21129 XA.Cn[1].n36 XA.Cn[1].n34 161.406
R21130 XA.Cn[1].n39 XA.Cn[1].n37 161.406
R21131 XA.Cn[1].n42 XA.Cn[1].n40 161.406
R21132 XA.Cn[1].n45 XA.Cn[1].n43 161.406
R21133 XA.Cn[1].n48 XA.Cn[1].n46 161.406
R21134 XA.Cn[1].n51 XA.Cn[1].n49 161.406
R21135 XA.Cn[1].n54 XA.Cn[1].n52 161.406
R21136 XA.Cn[1].n57 XA.Cn[1].n55 161.406
R21137 XA.Cn[1].n10 XA.Cn[1].t29 161.202
R21138 XA.Cn[1].n13 XA.Cn[1].t14 161.202
R21139 XA.Cn[1].n16 XA.Cn[1].t16 161.202
R21140 XA.Cn[1].n19 XA.Cn[1].t18 161.202
R21141 XA.Cn[1].n22 XA.Cn[1].t39 161.202
R21142 XA.Cn[1].n25 XA.Cn[1].t40 161.202
R21143 XA.Cn[1].n28 XA.Cn[1].t21 161.202
R21144 XA.Cn[1].n31 XA.Cn[1].t30 161.202
R21145 XA.Cn[1].n34 XA.Cn[1].t32 161.202
R21146 XA.Cn[1].n37 XA.Cn[1].t19 161.202
R21147 XA.Cn[1].n40 XA.Cn[1].t20 161.202
R21148 XA.Cn[1].n43 XA.Cn[1].t33 161.202
R21149 XA.Cn[1].n46 XA.Cn[1].t41 161.202
R21150 XA.Cn[1].n49 XA.Cn[1].t12 161.202
R21151 XA.Cn[1].n52 XA.Cn[1].t25 161.202
R21152 XA.Cn[1].n55 XA.Cn[1].t35 161.202
R21153 XA.Cn[1].n10 XA.Cn[1].t31 145.137
R21154 XA.Cn[1].n13 XA.Cn[1].t17 145.137
R21155 XA.Cn[1].n16 XA.Cn[1].t22 145.137
R21156 XA.Cn[1].n19 XA.Cn[1].t23 145.137
R21157 XA.Cn[1].n22 XA.Cn[1].t42 145.137
R21158 XA.Cn[1].n25 XA.Cn[1].t43 145.137
R21159 XA.Cn[1].n28 XA.Cn[1].t27 145.137
R21160 XA.Cn[1].n31 XA.Cn[1].t34 145.137
R21161 XA.Cn[1].n34 XA.Cn[1].t36 145.137
R21162 XA.Cn[1].n37 XA.Cn[1].t24 145.137
R21163 XA.Cn[1].n40 XA.Cn[1].t26 145.137
R21164 XA.Cn[1].n43 XA.Cn[1].t37 145.137
R21165 XA.Cn[1].n46 XA.Cn[1].t13 145.137
R21166 XA.Cn[1].n49 XA.Cn[1].t15 145.137
R21167 XA.Cn[1].n52 XA.Cn[1].t28 145.137
R21168 XA.Cn[1].n55 XA.Cn[1].t38 145.137
R21169 XA.Cn[1].n5 XA.Cn[1].n3 135.249
R21170 XA.Cn[1].n5 XA.Cn[1].n4 98.981
R21171 XA.Cn[1].n7 XA.Cn[1].n6 98.981
R21172 XA.Cn[1].n9 XA.Cn[1].n8 98.981
R21173 XA.Cn[1].n7 XA.Cn[1].n5 36.2672
R21174 XA.Cn[1].n9 XA.Cn[1].n7 36.2672
R21175 XA.Cn[1].n59 XA.Cn[1].n9 32.6405
R21176 XA.Cn[1].n1 XA.Cn[1].t1 26.5955
R21177 XA.Cn[1].n1 XA.Cn[1].t0 26.5955
R21178 XA.Cn[1].n0 XA.Cn[1].t3 26.5955
R21179 XA.Cn[1].n0 XA.Cn[1].t2 26.5955
R21180 XA.Cn[1].n3 XA.Cn[1].t11 24.9236
R21181 XA.Cn[1].n3 XA.Cn[1].t10 24.9236
R21182 XA.Cn[1].n4 XA.Cn[1].t9 24.9236
R21183 XA.Cn[1].n4 XA.Cn[1].t8 24.9236
R21184 XA.Cn[1].n6 XA.Cn[1].t7 24.9236
R21185 XA.Cn[1].n6 XA.Cn[1].t6 24.9236
R21186 XA.Cn[1].n8 XA.Cn[1].t5 24.9236
R21187 XA.Cn[1].n8 XA.Cn[1].t4 24.9236
R21188 XA.Cn[1] XA.Cn[1].n2 23.3605
R21189 XA.Cn[1].n58 XA.Cn[1] 7.29217
R21190 XA.Cn[1] XA.Cn[1].n59 6.7205
R21191 XA.Cn[1].n59 XA.Cn[1].n58 3.13711
R21192 XA.Cn[1].n15 XA.Cn[1] 0.931056
R21193 XA.Cn[1].n18 XA.Cn[1] 0.931056
R21194 XA.Cn[1].n21 XA.Cn[1] 0.931056
R21195 XA.Cn[1].n24 XA.Cn[1] 0.931056
R21196 XA.Cn[1].n27 XA.Cn[1] 0.931056
R21197 XA.Cn[1].n30 XA.Cn[1] 0.931056
R21198 XA.Cn[1].n33 XA.Cn[1] 0.931056
R21199 XA.Cn[1].n36 XA.Cn[1] 0.931056
R21200 XA.Cn[1].n39 XA.Cn[1] 0.931056
R21201 XA.Cn[1].n42 XA.Cn[1] 0.931056
R21202 XA.Cn[1].n45 XA.Cn[1] 0.931056
R21203 XA.Cn[1].n48 XA.Cn[1] 0.931056
R21204 XA.Cn[1].n51 XA.Cn[1] 0.931056
R21205 XA.Cn[1].n54 XA.Cn[1] 0.931056
R21206 XA.Cn[1].n57 XA.Cn[1] 0.931056
R21207 XA.Cn[1] XA.Cn[1].n12 0.396333
R21208 XA.Cn[1] XA.Cn[1].n15 0.396333
R21209 XA.Cn[1] XA.Cn[1].n18 0.396333
R21210 XA.Cn[1] XA.Cn[1].n21 0.396333
R21211 XA.Cn[1] XA.Cn[1].n24 0.396333
R21212 XA.Cn[1] XA.Cn[1].n27 0.396333
R21213 XA.Cn[1] XA.Cn[1].n30 0.396333
R21214 XA.Cn[1] XA.Cn[1].n33 0.396333
R21215 XA.Cn[1] XA.Cn[1].n36 0.396333
R21216 XA.Cn[1] XA.Cn[1].n39 0.396333
R21217 XA.Cn[1] XA.Cn[1].n42 0.396333
R21218 XA.Cn[1] XA.Cn[1].n45 0.396333
R21219 XA.Cn[1] XA.Cn[1].n48 0.396333
R21220 XA.Cn[1] XA.Cn[1].n51 0.396333
R21221 XA.Cn[1] XA.Cn[1].n54 0.396333
R21222 XA.Cn[1] XA.Cn[1].n57 0.396333
R21223 XA.Cn[1].n11 XA.Cn[1] 0.104667
R21224 XA.Cn[1].n14 XA.Cn[1] 0.104667
R21225 XA.Cn[1].n17 XA.Cn[1] 0.104667
R21226 XA.Cn[1].n20 XA.Cn[1] 0.104667
R21227 XA.Cn[1].n23 XA.Cn[1] 0.104667
R21228 XA.Cn[1].n26 XA.Cn[1] 0.104667
R21229 XA.Cn[1].n29 XA.Cn[1] 0.104667
R21230 XA.Cn[1].n32 XA.Cn[1] 0.104667
R21231 XA.Cn[1].n35 XA.Cn[1] 0.104667
R21232 XA.Cn[1].n38 XA.Cn[1] 0.104667
R21233 XA.Cn[1].n41 XA.Cn[1] 0.104667
R21234 XA.Cn[1].n44 XA.Cn[1] 0.104667
R21235 XA.Cn[1].n47 XA.Cn[1] 0.104667
R21236 XA.Cn[1].n50 XA.Cn[1] 0.104667
R21237 XA.Cn[1].n53 XA.Cn[1] 0.104667
R21238 XA.Cn[1].n56 XA.Cn[1] 0.104667
R21239 XA.Cn[1].n58 XA.Cn[1] 0.0594286
R21240 XA.Cn[1].n11 XA.Cn[1] 0.0309878
R21241 XA.Cn[1].n14 XA.Cn[1] 0.0309878
R21242 XA.Cn[1].n17 XA.Cn[1] 0.0309878
R21243 XA.Cn[1].n20 XA.Cn[1] 0.0309878
R21244 XA.Cn[1].n23 XA.Cn[1] 0.0309878
R21245 XA.Cn[1].n26 XA.Cn[1] 0.0309878
R21246 XA.Cn[1].n29 XA.Cn[1] 0.0309878
R21247 XA.Cn[1].n32 XA.Cn[1] 0.0309878
R21248 XA.Cn[1].n35 XA.Cn[1] 0.0309878
R21249 XA.Cn[1].n38 XA.Cn[1] 0.0309878
R21250 XA.Cn[1].n41 XA.Cn[1] 0.0309878
R21251 XA.Cn[1].n44 XA.Cn[1] 0.0309878
R21252 XA.Cn[1].n47 XA.Cn[1] 0.0309878
R21253 XA.Cn[1].n50 XA.Cn[1] 0.0309878
R21254 XA.Cn[1].n53 XA.Cn[1] 0.0309878
R21255 XA.Cn[1].n56 XA.Cn[1] 0.0309878
R21256 XA.Cn[1].n12 XA.Cn[1].n11 0.027939
R21257 XA.Cn[1].n15 XA.Cn[1].n14 0.027939
R21258 XA.Cn[1].n18 XA.Cn[1].n17 0.027939
R21259 XA.Cn[1].n21 XA.Cn[1].n20 0.027939
R21260 XA.Cn[1].n24 XA.Cn[1].n23 0.027939
R21261 XA.Cn[1].n27 XA.Cn[1].n26 0.027939
R21262 XA.Cn[1].n30 XA.Cn[1].n29 0.027939
R21263 XA.Cn[1].n33 XA.Cn[1].n32 0.027939
R21264 XA.Cn[1].n36 XA.Cn[1].n35 0.027939
R21265 XA.Cn[1].n39 XA.Cn[1].n38 0.027939
R21266 XA.Cn[1].n42 XA.Cn[1].n41 0.027939
R21267 XA.Cn[1].n45 XA.Cn[1].n44 0.027939
R21268 XA.Cn[1].n48 XA.Cn[1].n47 0.027939
R21269 XA.Cn[1].n51 XA.Cn[1].n50 0.027939
R21270 XA.Cn[1].n54 XA.Cn[1].n53 0.027939
R21271 XA.Cn[1].n57 XA.Cn[1].n56 0.027939
R21272 XA.Cn[3].n2 XA.Cn[3].n1 332.332
R21273 XA.Cn[3].n2 XA.Cn[3].n0 296.493
R21274 XA.Cn[3].n12 XA.Cn[3].n10 161.406
R21275 XA.Cn[3].n15 XA.Cn[3].n13 161.406
R21276 XA.Cn[3].n18 XA.Cn[3].n16 161.406
R21277 XA.Cn[3].n21 XA.Cn[3].n19 161.406
R21278 XA.Cn[3].n24 XA.Cn[3].n22 161.406
R21279 XA.Cn[3].n27 XA.Cn[3].n25 161.406
R21280 XA.Cn[3].n30 XA.Cn[3].n28 161.406
R21281 XA.Cn[3].n33 XA.Cn[3].n31 161.406
R21282 XA.Cn[3].n36 XA.Cn[3].n34 161.406
R21283 XA.Cn[3].n39 XA.Cn[3].n37 161.406
R21284 XA.Cn[3].n42 XA.Cn[3].n40 161.406
R21285 XA.Cn[3].n45 XA.Cn[3].n43 161.406
R21286 XA.Cn[3].n48 XA.Cn[3].n46 161.406
R21287 XA.Cn[3].n51 XA.Cn[3].n49 161.406
R21288 XA.Cn[3].n54 XA.Cn[3].n52 161.406
R21289 XA.Cn[3].n57 XA.Cn[3].n55 161.406
R21290 XA.Cn[3].n10 XA.Cn[3].t42 161.202
R21291 XA.Cn[3].n13 XA.Cn[3].t27 161.202
R21292 XA.Cn[3].n16 XA.Cn[3].t29 161.202
R21293 XA.Cn[3].n19 XA.Cn[3].t31 161.202
R21294 XA.Cn[3].n22 XA.Cn[3].t20 161.202
R21295 XA.Cn[3].n25 XA.Cn[3].t21 161.202
R21296 XA.Cn[3].n28 XA.Cn[3].t34 161.202
R21297 XA.Cn[3].n31 XA.Cn[3].t43 161.202
R21298 XA.Cn[3].n34 XA.Cn[3].t13 161.202
R21299 XA.Cn[3].n37 XA.Cn[3].t32 161.202
R21300 XA.Cn[3].n40 XA.Cn[3].t33 161.202
R21301 XA.Cn[3].n43 XA.Cn[3].t14 161.202
R21302 XA.Cn[3].n46 XA.Cn[3].t22 161.202
R21303 XA.Cn[3].n49 XA.Cn[3].t25 161.202
R21304 XA.Cn[3].n52 XA.Cn[3].t38 161.202
R21305 XA.Cn[3].n55 XA.Cn[3].t16 161.202
R21306 XA.Cn[3].n10 XA.Cn[3].t12 145.137
R21307 XA.Cn[3].n13 XA.Cn[3].t30 145.137
R21308 XA.Cn[3].n16 XA.Cn[3].t35 145.137
R21309 XA.Cn[3].n19 XA.Cn[3].t36 145.137
R21310 XA.Cn[3].n22 XA.Cn[3].t23 145.137
R21311 XA.Cn[3].n25 XA.Cn[3].t24 145.137
R21312 XA.Cn[3].n28 XA.Cn[3].t40 145.137
R21313 XA.Cn[3].n31 XA.Cn[3].t15 145.137
R21314 XA.Cn[3].n34 XA.Cn[3].t17 145.137
R21315 XA.Cn[3].n37 XA.Cn[3].t37 145.137
R21316 XA.Cn[3].n40 XA.Cn[3].t39 145.137
R21317 XA.Cn[3].n43 XA.Cn[3].t18 145.137
R21318 XA.Cn[3].n46 XA.Cn[3].t26 145.137
R21319 XA.Cn[3].n49 XA.Cn[3].t28 145.137
R21320 XA.Cn[3].n52 XA.Cn[3].t41 145.137
R21321 XA.Cn[3].n55 XA.Cn[3].t19 145.137
R21322 XA.Cn[3].n7 XA.Cn[3].n6 135.249
R21323 XA.Cn[3].n9 XA.Cn[3].n3 98.981
R21324 XA.Cn[3].n8 XA.Cn[3].n4 98.981
R21325 XA.Cn[3].n7 XA.Cn[3].n5 98.981
R21326 XA.Cn[3].n9 XA.Cn[3].n8 36.2672
R21327 XA.Cn[3].n8 XA.Cn[3].n7 36.2672
R21328 XA.Cn[3].n58 XA.Cn[3].n9 32.6405
R21329 XA.Cn[3].n1 XA.Cn[3].t7 26.5955
R21330 XA.Cn[3].n1 XA.Cn[3].t6 26.5955
R21331 XA.Cn[3].n0 XA.Cn[3].t5 26.5955
R21332 XA.Cn[3].n0 XA.Cn[3].t4 26.5955
R21333 XA.Cn[3].n3 XA.Cn[3].t9 24.9236
R21334 XA.Cn[3].n3 XA.Cn[3].t8 24.9236
R21335 XA.Cn[3].n4 XA.Cn[3].t11 24.9236
R21336 XA.Cn[3].n4 XA.Cn[3].t10 24.9236
R21337 XA.Cn[3].n5 XA.Cn[3].t1 24.9236
R21338 XA.Cn[3].n5 XA.Cn[3].t0 24.9236
R21339 XA.Cn[3].n6 XA.Cn[3].t3 24.9236
R21340 XA.Cn[3].n6 XA.Cn[3].t2 24.9236
R21341 XA.Cn[3] XA.Cn[3].n2 23.3605
R21342 XA.Cn[3] XA.Cn[3].n58 6.7205
R21343 XA.Cn[3].n58 XA.Cn[3] 3.19574
R21344 XA.Cn[3].n15 XA.Cn[3] 0.931056
R21345 XA.Cn[3].n18 XA.Cn[3] 0.931056
R21346 XA.Cn[3].n21 XA.Cn[3] 0.931056
R21347 XA.Cn[3].n24 XA.Cn[3] 0.931056
R21348 XA.Cn[3].n27 XA.Cn[3] 0.931056
R21349 XA.Cn[3].n30 XA.Cn[3] 0.931056
R21350 XA.Cn[3].n33 XA.Cn[3] 0.931056
R21351 XA.Cn[3].n36 XA.Cn[3] 0.931056
R21352 XA.Cn[3].n39 XA.Cn[3] 0.931056
R21353 XA.Cn[3].n42 XA.Cn[3] 0.931056
R21354 XA.Cn[3].n45 XA.Cn[3] 0.931056
R21355 XA.Cn[3].n48 XA.Cn[3] 0.931056
R21356 XA.Cn[3].n51 XA.Cn[3] 0.931056
R21357 XA.Cn[3].n54 XA.Cn[3] 0.931056
R21358 XA.Cn[3].n57 XA.Cn[3] 0.931056
R21359 XA.Cn[3] XA.Cn[3].n12 0.396333
R21360 XA.Cn[3] XA.Cn[3].n15 0.396333
R21361 XA.Cn[3] XA.Cn[3].n18 0.396333
R21362 XA.Cn[3] XA.Cn[3].n21 0.396333
R21363 XA.Cn[3] XA.Cn[3].n24 0.396333
R21364 XA.Cn[3] XA.Cn[3].n27 0.396333
R21365 XA.Cn[3] XA.Cn[3].n30 0.396333
R21366 XA.Cn[3] XA.Cn[3].n33 0.396333
R21367 XA.Cn[3] XA.Cn[3].n36 0.396333
R21368 XA.Cn[3] XA.Cn[3].n39 0.396333
R21369 XA.Cn[3] XA.Cn[3].n42 0.396333
R21370 XA.Cn[3] XA.Cn[3].n45 0.396333
R21371 XA.Cn[3] XA.Cn[3].n48 0.396333
R21372 XA.Cn[3] XA.Cn[3].n51 0.396333
R21373 XA.Cn[3] XA.Cn[3].n54 0.396333
R21374 XA.Cn[3] XA.Cn[3].n57 0.396333
R21375 XA.Cn[3].n11 XA.Cn[3] 0.104667
R21376 XA.Cn[3].n14 XA.Cn[3] 0.104667
R21377 XA.Cn[3].n17 XA.Cn[3] 0.104667
R21378 XA.Cn[3].n20 XA.Cn[3] 0.104667
R21379 XA.Cn[3].n23 XA.Cn[3] 0.104667
R21380 XA.Cn[3].n26 XA.Cn[3] 0.104667
R21381 XA.Cn[3].n29 XA.Cn[3] 0.104667
R21382 XA.Cn[3].n32 XA.Cn[3] 0.104667
R21383 XA.Cn[3].n35 XA.Cn[3] 0.104667
R21384 XA.Cn[3].n38 XA.Cn[3] 0.104667
R21385 XA.Cn[3].n41 XA.Cn[3] 0.104667
R21386 XA.Cn[3].n44 XA.Cn[3] 0.104667
R21387 XA.Cn[3].n47 XA.Cn[3] 0.104667
R21388 XA.Cn[3].n50 XA.Cn[3] 0.104667
R21389 XA.Cn[3].n53 XA.Cn[3] 0.104667
R21390 XA.Cn[3].n56 XA.Cn[3] 0.104667
R21391 XA.Cn[3].n11 XA.Cn[3] 0.0309878
R21392 XA.Cn[3].n14 XA.Cn[3] 0.0309878
R21393 XA.Cn[3].n17 XA.Cn[3] 0.0309878
R21394 XA.Cn[3].n20 XA.Cn[3] 0.0309878
R21395 XA.Cn[3].n23 XA.Cn[3] 0.0309878
R21396 XA.Cn[3].n26 XA.Cn[3] 0.0309878
R21397 XA.Cn[3].n29 XA.Cn[3] 0.0309878
R21398 XA.Cn[3].n32 XA.Cn[3] 0.0309878
R21399 XA.Cn[3].n35 XA.Cn[3] 0.0309878
R21400 XA.Cn[3].n38 XA.Cn[3] 0.0309878
R21401 XA.Cn[3].n41 XA.Cn[3] 0.0309878
R21402 XA.Cn[3].n44 XA.Cn[3] 0.0309878
R21403 XA.Cn[3].n47 XA.Cn[3] 0.0309878
R21404 XA.Cn[3].n50 XA.Cn[3] 0.0309878
R21405 XA.Cn[3].n53 XA.Cn[3] 0.0309878
R21406 XA.Cn[3].n56 XA.Cn[3] 0.0309878
R21407 XA.Cn[3].n12 XA.Cn[3].n11 0.027939
R21408 XA.Cn[3].n15 XA.Cn[3].n14 0.027939
R21409 XA.Cn[3].n18 XA.Cn[3].n17 0.027939
R21410 XA.Cn[3].n21 XA.Cn[3].n20 0.027939
R21411 XA.Cn[3].n24 XA.Cn[3].n23 0.027939
R21412 XA.Cn[3].n27 XA.Cn[3].n26 0.027939
R21413 XA.Cn[3].n30 XA.Cn[3].n29 0.027939
R21414 XA.Cn[3].n33 XA.Cn[3].n32 0.027939
R21415 XA.Cn[3].n36 XA.Cn[3].n35 0.027939
R21416 XA.Cn[3].n39 XA.Cn[3].n38 0.027939
R21417 XA.Cn[3].n42 XA.Cn[3].n41 0.027939
R21418 XA.Cn[3].n45 XA.Cn[3].n44 0.027939
R21419 XA.Cn[3].n48 XA.Cn[3].n47 0.027939
R21420 XA.Cn[3].n51 XA.Cn[3].n50 0.027939
R21421 XA.Cn[3].n54 XA.Cn[3].n53 0.027939
R21422 XA.Cn[3].n57 XA.Cn[3].n56 0.027939
R21423 XThR.Tn[10].n87 XThR.Tn[10].n86 256.103
R21424 XThR.Tn[10].n2 XThR.Tn[10].n0 243.68
R21425 XThR.Tn[10].n5 XThR.Tn[10].n3 241.847
R21426 XThR.Tn[10].n2 XThR.Tn[10].n1 205.28
R21427 XThR.Tn[10].n87 XThR.Tn[10].n85 202.094
R21428 XThR.Tn[10].n5 XThR.Tn[10].n4 185
R21429 XThR.Tn[10] XThR.Tn[10].n78 161.363
R21430 XThR.Tn[10] XThR.Tn[10].n73 161.363
R21431 XThR.Tn[10] XThR.Tn[10].n68 161.363
R21432 XThR.Tn[10] XThR.Tn[10].n63 161.363
R21433 XThR.Tn[10] XThR.Tn[10].n58 161.363
R21434 XThR.Tn[10] XThR.Tn[10].n53 161.363
R21435 XThR.Tn[10] XThR.Tn[10].n48 161.363
R21436 XThR.Tn[10] XThR.Tn[10].n43 161.363
R21437 XThR.Tn[10] XThR.Tn[10].n38 161.363
R21438 XThR.Tn[10] XThR.Tn[10].n33 161.363
R21439 XThR.Tn[10] XThR.Tn[10].n28 161.363
R21440 XThR.Tn[10] XThR.Tn[10].n23 161.363
R21441 XThR.Tn[10] XThR.Tn[10].n18 161.363
R21442 XThR.Tn[10] XThR.Tn[10].n13 161.363
R21443 XThR.Tn[10] XThR.Tn[10].n8 161.363
R21444 XThR.Tn[10] XThR.Tn[10].n6 161.363
R21445 XThR.Tn[10].n80 XThR.Tn[10].n79 161.3
R21446 XThR.Tn[10].n75 XThR.Tn[10].n74 161.3
R21447 XThR.Tn[10].n70 XThR.Tn[10].n69 161.3
R21448 XThR.Tn[10].n65 XThR.Tn[10].n64 161.3
R21449 XThR.Tn[10].n60 XThR.Tn[10].n59 161.3
R21450 XThR.Tn[10].n55 XThR.Tn[10].n54 161.3
R21451 XThR.Tn[10].n50 XThR.Tn[10].n49 161.3
R21452 XThR.Tn[10].n45 XThR.Tn[10].n44 161.3
R21453 XThR.Tn[10].n40 XThR.Tn[10].n39 161.3
R21454 XThR.Tn[10].n35 XThR.Tn[10].n34 161.3
R21455 XThR.Tn[10].n30 XThR.Tn[10].n29 161.3
R21456 XThR.Tn[10].n25 XThR.Tn[10].n24 161.3
R21457 XThR.Tn[10].n20 XThR.Tn[10].n19 161.3
R21458 XThR.Tn[10].n15 XThR.Tn[10].n14 161.3
R21459 XThR.Tn[10].n10 XThR.Tn[10].n9 161.3
R21460 XThR.Tn[10].n78 XThR.Tn[10].t37 161.106
R21461 XThR.Tn[10].n73 XThR.Tn[10].t45 161.106
R21462 XThR.Tn[10].n68 XThR.Tn[10].t27 161.106
R21463 XThR.Tn[10].n63 XThR.Tn[10].t72 161.106
R21464 XThR.Tn[10].n58 XThR.Tn[10].t35 161.106
R21465 XThR.Tn[10].n53 XThR.Tn[10].t61 161.106
R21466 XThR.Tn[10].n48 XThR.Tn[10].t43 161.106
R21467 XThR.Tn[10].n43 XThR.Tn[10].t24 161.106
R21468 XThR.Tn[10].n38 XThR.Tn[10].t69 161.106
R21469 XThR.Tn[10].n33 XThR.Tn[10].t15 161.106
R21470 XThR.Tn[10].n28 XThR.Tn[10].t59 161.106
R21471 XThR.Tn[10].n23 XThR.Tn[10].t26 161.106
R21472 XThR.Tn[10].n18 XThR.Tn[10].t58 161.106
R21473 XThR.Tn[10].n13 XThR.Tn[10].t41 161.106
R21474 XThR.Tn[10].n8 XThR.Tn[10].t63 161.106
R21475 XThR.Tn[10].n6 XThR.Tn[10].t47 161.106
R21476 XThR.Tn[10].n79 XThR.Tn[10].t34 159.978
R21477 XThR.Tn[10].n74 XThR.Tn[10].t39 159.978
R21478 XThR.Tn[10].n69 XThR.Tn[10].t22 159.978
R21479 XThR.Tn[10].n64 XThR.Tn[10].t68 159.978
R21480 XThR.Tn[10].n59 XThR.Tn[10].t32 159.978
R21481 XThR.Tn[10].n54 XThR.Tn[10].t57 159.978
R21482 XThR.Tn[10].n49 XThR.Tn[10].t38 159.978
R21483 XThR.Tn[10].n44 XThR.Tn[10].t20 159.978
R21484 XThR.Tn[10].n39 XThR.Tn[10].t66 159.978
R21485 XThR.Tn[10].n34 XThR.Tn[10].t12 159.978
R21486 XThR.Tn[10].n29 XThR.Tn[10].t56 159.978
R21487 XThR.Tn[10].n24 XThR.Tn[10].t21 159.978
R21488 XThR.Tn[10].n19 XThR.Tn[10].t55 159.978
R21489 XThR.Tn[10].n14 XThR.Tn[10].t36 159.978
R21490 XThR.Tn[10].n9 XThR.Tn[10].t60 159.978
R21491 XThR.Tn[10].n78 XThR.Tn[10].t29 145.038
R21492 XThR.Tn[10].n73 XThR.Tn[10].t49 145.038
R21493 XThR.Tn[10].n68 XThR.Tn[10].t31 145.038
R21494 XThR.Tn[10].n63 XThR.Tn[10].t16 145.038
R21495 XThR.Tn[10].n58 XThR.Tn[10].t46 145.038
R21496 XThR.Tn[10].n53 XThR.Tn[10].t28 145.038
R21497 XThR.Tn[10].n48 XThR.Tn[10].t33 145.038
R21498 XThR.Tn[10].n43 XThR.Tn[10].t17 145.038
R21499 XThR.Tn[10].n38 XThR.Tn[10].t14 145.038
R21500 XThR.Tn[10].n33 XThR.Tn[10].t44 145.038
R21501 XThR.Tn[10].n28 XThR.Tn[10].t67 145.038
R21502 XThR.Tn[10].n23 XThR.Tn[10].t30 145.038
R21503 XThR.Tn[10].n18 XThR.Tn[10].t65 145.038
R21504 XThR.Tn[10].n13 XThR.Tn[10].t48 145.038
R21505 XThR.Tn[10].n8 XThR.Tn[10].t13 145.038
R21506 XThR.Tn[10].n6 XThR.Tn[10].t54 145.038
R21507 XThR.Tn[10].n79 XThR.Tn[10].t64 143.911
R21508 XThR.Tn[10].n74 XThR.Tn[10].t25 143.911
R21509 XThR.Tn[10].n69 XThR.Tn[10].t71 143.911
R21510 XThR.Tn[10].n64 XThR.Tn[10].t52 143.911
R21511 XThR.Tn[10].n59 XThR.Tn[10].t19 143.911
R21512 XThR.Tn[10].n54 XThR.Tn[10].t62 143.911
R21513 XThR.Tn[10].n49 XThR.Tn[10].t73 143.911
R21514 XThR.Tn[10].n44 XThR.Tn[10].t53 143.911
R21515 XThR.Tn[10].n39 XThR.Tn[10].t51 143.911
R21516 XThR.Tn[10].n34 XThR.Tn[10].t18 143.911
R21517 XThR.Tn[10].n29 XThR.Tn[10].t42 143.911
R21518 XThR.Tn[10].n24 XThR.Tn[10].t70 143.911
R21519 XThR.Tn[10].n19 XThR.Tn[10].t40 143.911
R21520 XThR.Tn[10].n14 XThR.Tn[10].t23 143.911
R21521 XThR.Tn[10].n9 XThR.Tn[10].t50 143.911
R21522 XThR.Tn[10] XThR.Tn[10].n2 35.7652
R21523 XThR.Tn[10].n86 XThR.Tn[10].t4 26.5955
R21524 XThR.Tn[10].n86 XThR.Tn[10].t3 26.5955
R21525 XThR.Tn[10].n0 XThR.Tn[10].t10 26.5955
R21526 XThR.Tn[10].n0 XThR.Tn[10].t8 26.5955
R21527 XThR.Tn[10].n1 XThR.Tn[10].t11 26.5955
R21528 XThR.Tn[10].n1 XThR.Tn[10].t9 26.5955
R21529 XThR.Tn[10].n85 XThR.Tn[10].t0 26.5955
R21530 XThR.Tn[10].n85 XThR.Tn[10].t5 26.5955
R21531 XThR.Tn[10].n4 XThR.Tn[10].t1 24.9236
R21532 XThR.Tn[10].n4 XThR.Tn[10].t6 24.9236
R21533 XThR.Tn[10].n3 XThR.Tn[10].t2 24.9236
R21534 XThR.Tn[10].n3 XThR.Tn[10].t7 24.9236
R21535 XThR.Tn[10] XThR.Tn[10].n5 18.8943
R21536 XThR.Tn[10].n88 XThR.Tn[10].n87 13.5534
R21537 XThR.Tn[10].n84 XThR.Tn[10] 7.84567
R21538 XThR.Tn[10].n84 XThR.Tn[10] 6.34069
R21539 XThR.Tn[10] XThR.Tn[10].n7 5.34038
R21540 XThR.Tn[10].n12 XThR.Tn[10].n11 4.5005
R21541 XThR.Tn[10].n17 XThR.Tn[10].n16 4.5005
R21542 XThR.Tn[10].n22 XThR.Tn[10].n21 4.5005
R21543 XThR.Tn[10].n27 XThR.Tn[10].n26 4.5005
R21544 XThR.Tn[10].n32 XThR.Tn[10].n31 4.5005
R21545 XThR.Tn[10].n37 XThR.Tn[10].n36 4.5005
R21546 XThR.Tn[10].n42 XThR.Tn[10].n41 4.5005
R21547 XThR.Tn[10].n47 XThR.Tn[10].n46 4.5005
R21548 XThR.Tn[10].n52 XThR.Tn[10].n51 4.5005
R21549 XThR.Tn[10].n57 XThR.Tn[10].n56 4.5005
R21550 XThR.Tn[10].n62 XThR.Tn[10].n61 4.5005
R21551 XThR.Tn[10].n67 XThR.Tn[10].n66 4.5005
R21552 XThR.Tn[10].n72 XThR.Tn[10].n71 4.5005
R21553 XThR.Tn[10].n77 XThR.Tn[10].n76 4.5005
R21554 XThR.Tn[10].n82 XThR.Tn[10].n81 4.5005
R21555 XThR.Tn[10].n83 XThR.Tn[10] 3.70586
R21556 XThR.Tn[10].n12 XThR.Tn[10] 2.52282
R21557 XThR.Tn[10].n17 XThR.Tn[10] 2.52282
R21558 XThR.Tn[10].n22 XThR.Tn[10] 2.52282
R21559 XThR.Tn[10].n27 XThR.Tn[10] 2.52282
R21560 XThR.Tn[10].n32 XThR.Tn[10] 2.52282
R21561 XThR.Tn[10].n37 XThR.Tn[10] 2.52282
R21562 XThR.Tn[10].n42 XThR.Tn[10] 2.52282
R21563 XThR.Tn[10].n47 XThR.Tn[10] 2.52282
R21564 XThR.Tn[10].n52 XThR.Tn[10] 2.52282
R21565 XThR.Tn[10].n57 XThR.Tn[10] 2.52282
R21566 XThR.Tn[10].n62 XThR.Tn[10] 2.52282
R21567 XThR.Tn[10].n67 XThR.Tn[10] 2.52282
R21568 XThR.Tn[10].n72 XThR.Tn[10] 2.52282
R21569 XThR.Tn[10].n77 XThR.Tn[10] 2.52282
R21570 XThR.Tn[10].n82 XThR.Tn[10] 2.52282
R21571 XThR.Tn[10] XThR.Tn[10].n84 1.79489
R21572 XThR.Tn[10] XThR.Tn[10].n88 1.50638
R21573 XThR.Tn[10].n88 XThR.Tn[10] 1.19676
R21574 XThR.Tn[10].n80 XThR.Tn[10] 1.08677
R21575 XThR.Tn[10].n75 XThR.Tn[10] 1.08677
R21576 XThR.Tn[10].n70 XThR.Tn[10] 1.08677
R21577 XThR.Tn[10].n65 XThR.Tn[10] 1.08677
R21578 XThR.Tn[10].n60 XThR.Tn[10] 1.08677
R21579 XThR.Tn[10].n55 XThR.Tn[10] 1.08677
R21580 XThR.Tn[10].n50 XThR.Tn[10] 1.08677
R21581 XThR.Tn[10].n45 XThR.Tn[10] 1.08677
R21582 XThR.Tn[10].n40 XThR.Tn[10] 1.08677
R21583 XThR.Tn[10].n35 XThR.Tn[10] 1.08677
R21584 XThR.Tn[10].n30 XThR.Tn[10] 1.08677
R21585 XThR.Tn[10].n25 XThR.Tn[10] 1.08677
R21586 XThR.Tn[10].n20 XThR.Tn[10] 1.08677
R21587 XThR.Tn[10].n15 XThR.Tn[10] 1.08677
R21588 XThR.Tn[10].n10 XThR.Tn[10] 1.08677
R21589 XThR.Tn[10] XThR.Tn[10].n12 0.839786
R21590 XThR.Tn[10] XThR.Tn[10].n17 0.839786
R21591 XThR.Tn[10] XThR.Tn[10].n22 0.839786
R21592 XThR.Tn[10] XThR.Tn[10].n27 0.839786
R21593 XThR.Tn[10] XThR.Tn[10].n32 0.839786
R21594 XThR.Tn[10] XThR.Tn[10].n37 0.839786
R21595 XThR.Tn[10] XThR.Tn[10].n42 0.839786
R21596 XThR.Tn[10] XThR.Tn[10].n47 0.839786
R21597 XThR.Tn[10] XThR.Tn[10].n52 0.839786
R21598 XThR.Tn[10] XThR.Tn[10].n57 0.839786
R21599 XThR.Tn[10] XThR.Tn[10].n62 0.839786
R21600 XThR.Tn[10] XThR.Tn[10].n67 0.839786
R21601 XThR.Tn[10] XThR.Tn[10].n72 0.839786
R21602 XThR.Tn[10] XThR.Tn[10].n77 0.839786
R21603 XThR.Tn[10] XThR.Tn[10].n82 0.839786
R21604 XThR.Tn[10].n7 XThR.Tn[10] 0.499542
R21605 XThR.Tn[10].n81 XThR.Tn[10] 0.063
R21606 XThR.Tn[10].n76 XThR.Tn[10] 0.063
R21607 XThR.Tn[10].n71 XThR.Tn[10] 0.063
R21608 XThR.Tn[10].n66 XThR.Tn[10] 0.063
R21609 XThR.Tn[10].n61 XThR.Tn[10] 0.063
R21610 XThR.Tn[10].n56 XThR.Tn[10] 0.063
R21611 XThR.Tn[10].n51 XThR.Tn[10] 0.063
R21612 XThR.Tn[10].n46 XThR.Tn[10] 0.063
R21613 XThR.Tn[10].n41 XThR.Tn[10] 0.063
R21614 XThR.Tn[10].n36 XThR.Tn[10] 0.063
R21615 XThR.Tn[10].n31 XThR.Tn[10] 0.063
R21616 XThR.Tn[10].n26 XThR.Tn[10] 0.063
R21617 XThR.Tn[10].n21 XThR.Tn[10] 0.063
R21618 XThR.Tn[10].n16 XThR.Tn[10] 0.063
R21619 XThR.Tn[10].n11 XThR.Tn[10] 0.063
R21620 XThR.Tn[10].n83 XThR.Tn[10] 0.0540714
R21621 XThR.Tn[10] XThR.Tn[10].n83 0.038
R21622 XThR.Tn[10].n7 XThR.Tn[10] 0.0143889
R21623 XThR.Tn[10].n81 XThR.Tn[10].n80 0.00771154
R21624 XThR.Tn[10].n76 XThR.Tn[10].n75 0.00771154
R21625 XThR.Tn[10].n71 XThR.Tn[10].n70 0.00771154
R21626 XThR.Tn[10].n66 XThR.Tn[10].n65 0.00771154
R21627 XThR.Tn[10].n61 XThR.Tn[10].n60 0.00771154
R21628 XThR.Tn[10].n56 XThR.Tn[10].n55 0.00771154
R21629 XThR.Tn[10].n51 XThR.Tn[10].n50 0.00771154
R21630 XThR.Tn[10].n46 XThR.Tn[10].n45 0.00771154
R21631 XThR.Tn[10].n41 XThR.Tn[10].n40 0.00771154
R21632 XThR.Tn[10].n36 XThR.Tn[10].n35 0.00771154
R21633 XThR.Tn[10].n31 XThR.Tn[10].n30 0.00771154
R21634 XThR.Tn[10].n26 XThR.Tn[10].n25 0.00771154
R21635 XThR.Tn[10].n21 XThR.Tn[10].n20 0.00771154
R21636 XThR.Tn[10].n16 XThR.Tn[10].n15 0.00771154
R21637 XThR.Tn[10].n11 XThR.Tn[10].n10 0.00771154
R21638 XA.Cn[14].n55 XA.Cn[14].n54 256.104
R21639 XA.Cn[14].n59 XA.Cn[14].n58 243.679
R21640 XA.Cn[14].n2 XA.Cn[14].n0 241.847
R21641 XA.Cn[14].n59 XA.Cn[14].n57 205.28
R21642 XA.Cn[14].n55 XA.Cn[14].n53 202.095
R21643 XA.Cn[14].n2 XA.Cn[14].n1 185
R21644 XA.Cn[14].n5 XA.Cn[14].n3 161.406
R21645 XA.Cn[14].n8 XA.Cn[14].n6 161.406
R21646 XA.Cn[14].n11 XA.Cn[14].n9 161.406
R21647 XA.Cn[14].n14 XA.Cn[14].n12 161.406
R21648 XA.Cn[14].n17 XA.Cn[14].n15 161.406
R21649 XA.Cn[14].n20 XA.Cn[14].n18 161.406
R21650 XA.Cn[14].n23 XA.Cn[14].n21 161.406
R21651 XA.Cn[14].n26 XA.Cn[14].n24 161.406
R21652 XA.Cn[14].n29 XA.Cn[14].n27 161.406
R21653 XA.Cn[14].n32 XA.Cn[14].n30 161.406
R21654 XA.Cn[14].n35 XA.Cn[14].n33 161.406
R21655 XA.Cn[14].n38 XA.Cn[14].n36 161.406
R21656 XA.Cn[14].n41 XA.Cn[14].n39 161.406
R21657 XA.Cn[14].n44 XA.Cn[14].n42 161.406
R21658 XA.Cn[14].n47 XA.Cn[14].n45 161.406
R21659 XA.Cn[14].n50 XA.Cn[14].n48 161.406
R21660 XA.Cn[14].n3 XA.Cn[14].t38 161.202
R21661 XA.Cn[14].n6 XA.Cn[14].t22 161.202
R21662 XA.Cn[14].n9 XA.Cn[14].t25 161.202
R21663 XA.Cn[14].n12 XA.Cn[14].t26 161.202
R21664 XA.Cn[14].n15 XA.Cn[14].t14 161.202
R21665 XA.Cn[14].n18 XA.Cn[14].t17 161.202
R21666 XA.Cn[14].n21 XA.Cn[14].t31 161.202
R21667 XA.Cn[14].n24 XA.Cn[14].t39 161.202
R21668 XA.Cn[14].n27 XA.Cn[14].t41 161.202
R21669 XA.Cn[14].n30 XA.Cn[14].t27 161.202
R21670 XA.Cn[14].n33 XA.Cn[14].t30 161.202
R21671 XA.Cn[14].n36 XA.Cn[14].t42 161.202
R21672 XA.Cn[14].n39 XA.Cn[14].t19 161.202
R21673 XA.Cn[14].n42 XA.Cn[14].t21 161.202
R21674 XA.Cn[14].n45 XA.Cn[14].t33 161.202
R21675 XA.Cn[14].n48 XA.Cn[14].t12 161.202
R21676 XA.Cn[14].n3 XA.Cn[14].t43 145.137
R21677 XA.Cn[14].n6 XA.Cn[14].t29 145.137
R21678 XA.Cn[14].n9 XA.Cn[14].t32 145.137
R21679 XA.Cn[14].n12 XA.Cn[14].t34 145.137
R21680 XA.Cn[14].n15 XA.Cn[14].t20 145.137
R21681 XA.Cn[14].n18 XA.Cn[14].t23 145.137
R21682 XA.Cn[14].n21 XA.Cn[14].t37 145.137
R21683 XA.Cn[14].n24 XA.Cn[14].t13 145.137
R21684 XA.Cn[14].n27 XA.Cn[14].t15 145.137
R21685 XA.Cn[14].n30 XA.Cn[14].t35 145.137
R21686 XA.Cn[14].n33 XA.Cn[14].t36 145.137
R21687 XA.Cn[14].n36 XA.Cn[14].t16 145.137
R21688 XA.Cn[14].n39 XA.Cn[14].t24 145.137
R21689 XA.Cn[14].n42 XA.Cn[14].t28 145.137
R21690 XA.Cn[14].n45 XA.Cn[14].t40 145.137
R21691 XA.Cn[14].n48 XA.Cn[14].t18 145.137
R21692 XA.Cn[14].n53 XA.Cn[14].t4 26.5955
R21693 XA.Cn[14].n53 XA.Cn[14].t5 26.5955
R21694 XA.Cn[14].n54 XA.Cn[14].t7 26.5955
R21695 XA.Cn[14].n54 XA.Cn[14].t6 26.5955
R21696 XA.Cn[14].n57 XA.Cn[14].t1 26.5955
R21697 XA.Cn[14].n57 XA.Cn[14].t0 26.5955
R21698 XA.Cn[14].n58 XA.Cn[14].t3 26.5955
R21699 XA.Cn[14].n58 XA.Cn[14].t2 26.5955
R21700 XA.Cn[14].n1 XA.Cn[14].t9 24.9236
R21701 XA.Cn[14].n1 XA.Cn[14].t11 24.9236
R21702 XA.Cn[14].n0 XA.Cn[14].t8 24.9236
R21703 XA.Cn[14].n0 XA.Cn[14].t10 24.9236
R21704 XA.Cn[14] XA.Cn[14].n59 22.9652
R21705 XA.Cn[14] XA.Cn[14].n2 22.9615
R21706 XA.Cn[14].n56 XA.Cn[14].n55 13.9299
R21707 XA.Cn[14] XA.Cn[14].n56 13.9299
R21708 XA.Cn[14].n51 XA.Cn[14] 5.65386
R21709 XA.Cn[14].n52 XA.Cn[14].n51 5.13312
R21710 XA.Cn[14].n56 XA.Cn[14].n52 2.99115
R21711 XA.Cn[14].n56 XA.Cn[14] 2.87153
R21712 XA.Cn[14].n52 XA.Cn[14] 2.2734
R21713 XA.Cn[14].n8 XA.Cn[14] 0.931056
R21714 XA.Cn[14].n11 XA.Cn[14] 0.931056
R21715 XA.Cn[14].n14 XA.Cn[14] 0.931056
R21716 XA.Cn[14].n17 XA.Cn[14] 0.931056
R21717 XA.Cn[14].n20 XA.Cn[14] 0.931056
R21718 XA.Cn[14].n23 XA.Cn[14] 0.931056
R21719 XA.Cn[14].n26 XA.Cn[14] 0.931056
R21720 XA.Cn[14].n29 XA.Cn[14] 0.931056
R21721 XA.Cn[14].n32 XA.Cn[14] 0.931056
R21722 XA.Cn[14].n35 XA.Cn[14] 0.931056
R21723 XA.Cn[14].n38 XA.Cn[14] 0.931056
R21724 XA.Cn[14].n41 XA.Cn[14] 0.931056
R21725 XA.Cn[14].n44 XA.Cn[14] 0.931056
R21726 XA.Cn[14].n47 XA.Cn[14] 0.931056
R21727 XA.Cn[14].n50 XA.Cn[14] 0.931056
R21728 XA.Cn[14] XA.Cn[14].n5 0.396333
R21729 XA.Cn[14] XA.Cn[14].n8 0.396333
R21730 XA.Cn[14] XA.Cn[14].n11 0.396333
R21731 XA.Cn[14] XA.Cn[14].n14 0.396333
R21732 XA.Cn[14] XA.Cn[14].n17 0.396333
R21733 XA.Cn[14] XA.Cn[14].n20 0.396333
R21734 XA.Cn[14] XA.Cn[14].n23 0.396333
R21735 XA.Cn[14] XA.Cn[14].n26 0.396333
R21736 XA.Cn[14] XA.Cn[14].n29 0.396333
R21737 XA.Cn[14] XA.Cn[14].n32 0.396333
R21738 XA.Cn[14] XA.Cn[14].n35 0.396333
R21739 XA.Cn[14] XA.Cn[14].n38 0.396333
R21740 XA.Cn[14] XA.Cn[14].n41 0.396333
R21741 XA.Cn[14] XA.Cn[14].n44 0.396333
R21742 XA.Cn[14] XA.Cn[14].n47 0.396333
R21743 XA.Cn[14] XA.Cn[14].n50 0.396333
R21744 XA.Cn[14].n4 XA.Cn[14] 0.104667
R21745 XA.Cn[14].n7 XA.Cn[14] 0.104667
R21746 XA.Cn[14].n10 XA.Cn[14] 0.104667
R21747 XA.Cn[14].n13 XA.Cn[14] 0.104667
R21748 XA.Cn[14].n16 XA.Cn[14] 0.104667
R21749 XA.Cn[14].n19 XA.Cn[14] 0.104667
R21750 XA.Cn[14].n22 XA.Cn[14] 0.104667
R21751 XA.Cn[14].n25 XA.Cn[14] 0.104667
R21752 XA.Cn[14].n28 XA.Cn[14] 0.104667
R21753 XA.Cn[14].n31 XA.Cn[14] 0.104667
R21754 XA.Cn[14].n34 XA.Cn[14] 0.104667
R21755 XA.Cn[14].n37 XA.Cn[14] 0.104667
R21756 XA.Cn[14].n40 XA.Cn[14] 0.104667
R21757 XA.Cn[14].n43 XA.Cn[14] 0.104667
R21758 XA.Cn[14].n46 XA.Cn[14] 0.104667
R21759 XA.Cn[14].n49 XA.Cn[14] 0.104667
R21760 XA.Cn[14].n4 XA.Cn[14] 0.0309878
R21761 XA.Cn[14].n7 XA.Cn[14] 0.0309878
R21762 XA.Cn[14].n10 XA.Cn[14] 0.0309878
R21763 XA.Cn[14].n13 XA.Cn[14] 0.0309878
R21764 XA.Cn[14].n16 XA.Cn[14] 0.0309878
R21765 XA.Cn[14].n19 XA.Cn[14] 0.0309878
R21766 XA.Cn[14].n22 XA.Cn[14] 0.0309878
R21767 XA.Cn[14].n25 XA.Cn[14] 0.0309878
R21768 XA.Cn[14].n28 XA.Cn[14] 0.0309878
R21769 XA.Cn[14].n31 XA.Cn[14] 0.0309878
R21770 XA.Cn[14].n34 XA.Cn[14] 0.0309878
R21771 XA.Cn[14].n37 XA.Cn[14] 0.0309878
R21772 XA.Cn[14].n40 XA.Cn[14] 0.0309878
R21773 XA.Cn[14].n43 XA.Cn[14] 0.0309878
R21774 XA.Cn[14].n46 XA.Cn[14] 0.0309878
R21775 XA.Cn[14].n49 XA.Cn[14] 0.0309878
R21776 XA.Cn[14].n5 XA.Cn[14].n4 0.027939
R21777 XA.Cn[14].n8 XA.Cn[14].n7 0.027939
R21778 XA.Cn[14].n11 XA.Cn[14].n10 0.027939
R21779 XA.Cn[14].n14 XA.Cn[14].n13 0.027939
R21780 XA.Cn[14].n17 XA.Cn[14].n16 0.027939
R21781 XA.Cn[14].n20 XA.Cn[14].n19 0.027939
R21782 XA.Cn[14].n23 XA.Cn[14].n22 0.027939
R21783 XA.Cn[14].n26 XA.Cn[14].n25 0.027939
R21784 XA.Cn[14].n29 XA.Cn[14].n28 0.027939
R21785 XA.Cn[14].n32 XA.Cn[14].n31 0.027939
R21786 XA.Cn[14].n35 XA.Cn[14].n34 0.027939
R21787 XA.Cn[14].n38 XA.Cn[14].n37 0.027939
R21788 XA.Cn[14].n41 XA.Cn[14].n40 0.027939
R21789 XA.Cn[14].n44 XA.Cn[14].n43 0.027939
R21790 XA.Cn[14].n47 XA.Cn[14].n46 0.027939
R21791 XA.Cn[14].n50 XA.Cn[14].n49 0.027939
R21792 XA.Cn[14].n51 XA.Cn[14] 0.00250754
R21793 thermo15c_0.XTB1.Y.n6 thermo15c_0.XTB1.Y.t11 212.081
R21794 thermo15c_0.XTB1.Y.n5 thermo15c_0.XTB1.Y.t8 212.081
R21795 thermo15c_0.XTB1.Y.n11 thermo15c_0.XTB1.Y.t6 212.081
R21796 thermo15c_0.XTB1.Y.n3 thermo15c_0.XTB1.Y.t17 212.081
R21797 thermo15c_0.XTB1.Y.n15 thermo15c_0.XTB1.Y.t10 212.081
R21798 thermo15c_0.XTB1.Y.n16 thermo15c_0.XTB1.Y.t14 212.081
R21799 thermo15c_0.XTB1.Y.n18 thermo15c_0.XTB1.Y.t7 212.081
R21800 thermo15c_0.XTB1.Y.n14 thermo15c_0.XTB1.Y.t18 212.081
R21801 thermo15c_0.XTB1.Y.n22 thermo15c_0.XTB1.Y.n2 201.288
R21802 thermo15c_0.XTB1.Y.n8 thermo15c_0.XTB1.Y.n7 173.761
R21803 thermo15c_0.XTB1.Y.n17 thermo15c_0.XTB1.Y 158.656
R21804 thermo15c_0.XTB1.Y.n10 thermo15c_0.XTB1.Y.n9 152
R21805 thermo15c_0.XTB1.Y.n8 thermo15c_0.XTB1.Y.n4 152
R21806 thermo15c_0.XTB1.Y.n13 thermo15c_0.XTB1.Y.n12 152
R21807 thermo15c_0.XTB1.Y.n20 thermo15c_0.XTB1.Y.n19 152
R21808 thermo15c_0.XTB1.Y.n6 thermo15c_0.XTB1.Y.t16 139.78
R21809 thermo15c_0.XTB1.Y.n5 thermo15c_0.XTB1.Y.t13 139.78
R21810 thermo15c_0.XTB1.Y.n11 thermo15c_0.XTB1.Y.t12 139.78
R21811 thermo15c_0.XTB1.Y.n3 thermo15c_0.XTB1.Y.t5 139.78
R21812 thermo15c_0.XTB1.Y.n15 thermo15c_0.XTB1.Y.t4 139.78
R21813 thermo15c_0.XTB1.Y.n16 thermo15c_0.XTB1.Y.t3 139.78
R21814 thermo15c_0.XTB1.Y.n18 thermo15c_0.XTB1.Y.t15 139.78
R21815 thermo15c_0.XTB1.Y.n14 thermo15c_0.XTB1.Y.t9 139.78
R21816 thermo15c_0.XTB1.Y.n0 thermo15c_0.XTB1.Y.t1 132.067
R21817 thermo15c_0.XTB1.Y.n21 thermo15c_0.XTB1.Y 83.4676
R21818 thermo15c_0.XTB1.Y.n21 thermo15c_0.XTB1.Y.n13 61.4091
R21819 thermo15c_0.XTB1.Y.n16 thermo15c_0.XTB1.Y.n15 61.346
R21820 thermo15c_0.XTB1.Y.n10 thermo15c_0.XTB1.Y.n4 49.6611
R21821 thermo15c_0.XTB1.Y.n12 thermo15c_0.XTB1.Y.n11 45.2793
R21822 thermo15c_0.XTB1.Y.n7 thermo15c_0.XTB1.Y.n5 42.3581
R21823 thermo15c_0.XTB1.Y.n19 thermo15c_0.XTB1.Y.n14 30.6732
R21824 thermo15c_0.XTB1.Y.n19 thermo15c_0.XTB1.Y.n18 30.6732
R21825 thermo15c_0.XTB1.Y.n18 thermo15c_0.XTB1.Y.n17 30.6732
R21826 thermo15c_0.XTB1.Y.n17 thermo15c_0.XTB1.Y.n16 30.6732
R21827 thermo15c_0.XTB1.Y.n2 thermo15c_0.XTB1.Y.t2 26.5955
R21828 thermo15c_0.XTB1.Y.n2 thermo15c_0.XTB1.Y.t0 26.5955
R21829 thermo15c_0.XTB1.Y thermo15c_0.XTB1.Y.n22 23.489
R21830 thermo15c_0.XTB1.Y.n9 thermo15c_0.XTB1.Y.n8 21.7605
R21831 thermo15c_0.XTB1.Y.n7 thermo15c_0.XTB1.Y.n6 18.9884
R21832 thermo15c_0.XTB1.Y.n12 thermo15c_0.XTB1.Y.n3 16.0672
R21833 thermo15c_0.XTB1.Y.n20 thermo15c_0.XTB1.Y 14.8485
R21834 thermo15c_0.XTB1.Y.n13 thermo15c_0.XTB1.Y 11.5205
R21835 thermo15c_0.XTB1.Y.n22 thermo15c_0.XTB1.Y.n21 10.7939
R21836 thermo15c_0.XTB1.Y.n9 thermo15c_0.XTB1.Y 10.2405
R21837 thermo15c_0.XTB1.Y thermo15c_0.XTB1.Y.n20 8.7045
R21838 thermo15c_0.XTB1.Y.n5 thermo15c_0.XTB1.Y.n4 7.30353
R21839 thermo15c_0.XTB1.Y.n11 thermo15c_0.XTB1.Y.n10 4.38232
R21840 thermo15c_0.XTB1.Y.n1 thermo15c_0.XTB1.Y.n0 4.15748
R21841 thermo15c_0.XTB1.Y thermo15c_0.XTB1.Y.n1 3.76521
R21842 thermo15c_0.XTB1.Y.n0 thermo15c_0.XTB1.Y 1.17559
R21843 thermo15c_0.XTB1.Y.n1 thermo15c_0.XTB1.Y 0.921363
R21844 XA.Cn[8].n56 XA.Cn[8].n55 256.103
R21845 XA.Cn[8].n60 XA.Cn[8].n58 243.68
R21846 XA.Cn[8].n2 XA.Cn[8].n0 241.847
R21847 XA.Cn[8].n60 XA.Cn[8].n59 205.28
R21848 XA.Cn[8].n56 XA.Cn[8].n54 202.095
R21849 XA.Cn[8].n2 XA.Cn[8].n1 185
R21850 XA.Cn[8].n5 XA.Cn[8].n3 161.406
R21851 XA.Cn[8].n8 XA.Cn[8].n6 161.406
R21852 XA.Cn[8].n11 XA.Cn[8].n9 161.406
R21853 XA.Cn[8].n14 XA.Cn[8].n12 161.406
R21854 XA.Cn[8].n17 XA.Cn[8].n15 161.406
R21855 XA.Cn[8].n20 XA.Cn[8].n18 161.406
R21856 XA.Cn[8].n23 XA.Cn[8].n21 161.406
R21857 XA.Cn[8].n26 XA.Cn[8].n24 161.406
R21858 XA.Cn[8].n29 XA.Cn[8].n27 161.406
R21859 XA.Cn[8].n32 XA.Cn[8].n30 161.406
R21860 XA.Cn[8].n35 XA.Cn[8].n33 161.406
R21861 XA.Cn[8].n38 XA.Cn[8].n36 161.406
R21862 XA.Cn[8].n41 XA.Cn[8].n39 161.406
R21863 XA.Cn[8].n44 XA.Cn[8].n42 161.406
R21864 XA.Cn[8].n47 XA.Cn[8].n45 161.406
R21865 XA.Cn[8].n50 XA.Cn[8].n48 161.406
R21866 XA.Cn[8].n3 XA.Cn[8].t41 161.202
R21867 XA.Cn[8].n6 XA.Cn[8].t26 161.202
R21868 XA.Cn[8].n9 XA.Cn[8].t28 161.202
R21869 XA.Cn[8].n12 XA.Cn[8].t30 161.202
R21870 XA.Cn[8].n15 XA.Cn[8].t19 161.202
R21871 XA.Cn[8].n18 XA.Cn[8].t20 161.202
R21872 XA.Cn[8].n21 XA.Cn[8].t33 161.202
R21873 XA.Cn[8].n24 XA.Cn[8].t42 161.202
R21874 XA.Cn[8].n27 XA.Cn[8].t12 161.202
R21875 XA.Cn[8].n30 XA.Cn[8].t31 161.202
R21876 XA.Cn[8].n33 XA.Cn[8].t32 161.202
R21877 XA.Cn[8].n36 XA.Cn[8].t13 161.202
R21878 XA.Cn[8].n39 XA.Cn[8].t21 161.202
R21879 XA.Cn[8].n42 XA.Cn[8].t24 161.202
R21880 XA.Cn[8].n45 XA.Cn[8].t37 161.202
R21881 XA.Cn[8].n48 XA.Cn[8].t15 161.202
R21882 XA.Cn[8].n3 XA.Cn[8].t43 145.137
R21883 XA.Cn[8].n6 XA.Cn[8].t29 145.137
R21884 XA.Cn[8].n9 XA.Cn[8].t34 145.137
R21885 XA.Cn[8].n12 XA.Cn[8].t35 145.137
R21886 XA.Cn[8].n15 XA.Cn[8].t22 145.137
R21887 XA.Cn[8].n18 XA.Cn[8].t23 145.137
R21888 XA.Cn[8].n21 XA.Cn[8].t39 145.137
R21889 XA.Cn[8].n24 XA.Cn[8].t14 145.137
R21890 XA.Cn[8].n27 XA.Cn[8].t16 145.137
R21891 XA.Cn[8].n30 XA.Cn[8].t36 145.137
R21892 XA.Cn[8].n33 XA.Cn[8].t38 145.137
R21893 XA.Cn[8].n36 XA.Cn[8].t17 145.137
R21894 XA.Cn[8].n39 XA.Cn[8].t25 145.137
R21895 XA.Cn[8].n42 XA.Cn[8].t27 145.137
R21896 XA.Cn[8].n45 XA.Cn[8].t40 145.137
R21897 XA.Cn[8].n48 XA.Cn[8].t18 145.137
R21898 XA.Cn[8].n54 XA.Cn[8].t1 26.5955
R21899 XA.Cn[8].n54 XA.Cn[8].t2 26.5955
R21900 XA.Cn[8].n58 XA.Cn[8].t8 26.5955
R21901 XA.Cn[8].n58 XA.Cn[8].t11 26.5955
R21902 XA.Cn[8].n59 XA.Cn[8].t10 26.5955
R21903 XA.Cn[8].n59 XA.Cn[8].t9 26.5955
R21904 XA.Cn[8].n55 XA.Cn[8].t0 26.5955
R21905 XA.Cn[8].n55 XA.Cn[8].t3 26.5955
R21906 XA.Cn[8].n1 XA.Cn[8].t7 24.9236
R21907 XA.Cn[8].n1 XA.Cn[8].t6 24.9236
R21908 XA.Cn[8].n0 XA.Cn[8].t5 24.9236
R21909 XA.Cn[8].n0 XA.Cn[8].t4 24.9236
R21910 XA.Cn[8] XA.Cn[8].n60 22.9652
R21911 XA.Cn[8] XA.Cn[8].n2 22.9615
R21912 XA.Cn[8].n57 XA.Cn[8].n56 13.9299
R21913 XA.Cn[8] XA.Cn[8].n57 13.9299
R21914 XA.Cn[8].n53 XA.Cn[8].n52 5.09639
R21915 XA.Cn[8].n57 XA.Cn[8].n53 2.99115
R21916 XA.Cn[8].n57 XA.Cn[8] 2.87153
R21917 XA.Cn[8].n53 XA.Cn[8] 2.2734
R21918 XA.Cn[8].n51 XA.Cn[8] 1.14336
R21919 XA.Cn[8].n8 XA.Cn[8] 0.931056
R21920 XA.Cn[8].n11 XA.Cn[8] 0.931056
R21921 XA.Cn[8].n14 XA.Cn[8] 0.931056
R21922 XA.Cn[8].n17 XA.Cn[8] 0.931056
R21923 XA.Cn[8].n20 XA.Cn[8] 0.931056
R21924 XA.Cn[8].n23 XA.Cn[8] 0.931056
R21925 XA.Cn[8].n26 XA.Cn[8] 0.931056
R21926 XA.Cn[8].n29 XA.Cn[8] 0.931056
R21927 XA.Cn[8].n32 XA.Cn[8] 0.931056
R21928 XA.Cn[8].n35 XA.Cn[8] 0.931056
R21929 XA.Cn[8].n38 XA.Cn[8] 0.931056
R21930 XA.Cn[8].n41 XA.Cn[8] 0.931056
R21931 XA.Cn[8].n44 XA.Cn[8] 0.931056
R21932 XA.Cn[8].n47 XA.Cn[8] 0.931056
R21933 XA.Cn[8].n50 XA.Cn[8] 0.931056
R21934 XA.Cn[8] XA.Cn[8].n5 0.396333
R21935 XA.Cn[8] XA.Cn[8].n8 0.396333
R21936 XA.Cn[8] XA.Cn[8].n11 0.396333
R21937 XA.Cn[8] XA.Cn[8].n14 0.396333
R21938 XA.Cn[8] XA.Cn[8].n17 0.396333
R21939 XA.Cn[8] XA.Cn[8].n20 0.396333
R21940 XA.Cn[8] XA.Cn[8].n23 0.396333
R21941 XA.Cn[8] XA.Cn[8].n26 0.396333
R21942 XA.Cn[8] XA.Cn[8].n29 0.396333
R21943 XA.Cn[8] XA.Cn[8].n32 0.396333
R21944 XA.Cn[8] XA.Cn[8].n35 0.396333
R21945 XA.Cn[8] XA.Cn[8].n38 0.396333
R21946 XA.Cn[8] XA.Cn[8].n41 0.396333
R21947 XA.Cn[8] XA.Cn[8].n44 0.396333
R21948 XA.Cn[8] XA.Cn[8].n47 0.396333
R21949 XA.Cn[8] XA.Cn[8].n50 0.396333
R21950 XA.Cn[8].n52 XA.Cn[8].n51 0.166125
R21951 XA.Cn[8].n4 XA.Cn[8] 0.104667
R21952 XA.Cn[8].n7 XA.Cn[8] 0.104667
R21953 XA.Cn[8].n10 XA.Cn[8] 0.104667
R21954 XA.Cn[8].n13 XA.Cn[8] 0.104667
R21955 XA.Cn[8].n16 XA.Cn[8] 0.104667
R21956 XA.Cn[8].n19 XA.Cn[8] 0.104667
R21957 XA.Cn[8].n22 XA.Cn[8] 0.104667
R21958 XA.Cn[8].n25 XA.Cn[8] 0.104667
R21959 XA.Cn[8].n28 XA.Cn[8] 0.104667
R21960 XA.Cn[8].n31 XA.Cn[8] 0.104667
R21961 XA.Cn[8].n34 XA.Cn[8] 0.104667
R21962 XA.Cn[8].n37 XA.Cn[8] 0.104667
R21963 XA.Cn[8].n40 XA.Cn[8] 0.104667
R21964 XA.Cn[8].n43 XA.Cn[8] 0.104667
R21965 XA.Cn[8].n46 XA.Cn[8] 0.104667
R21966 XA.Cn[8].n49 XA.Cn[8] 0.104667
R21967 XA.Cn[8].n52 XA.Cn[8] 0.0389615
R21968 XA.Cn[8].n51 XA.Cn[8] 0.038
R21969 XA.Cn[8].n4 XA.Cn[8] 0.0309878
R21970 XA.Cn[8].n7 XA.Cn[8] 0.0309878
R21971 XA.Cn[8].n10 XA.Cn[8] 0.0309878
R21972 XA.Cn[8].n13 XA.Cn[8] 0.0309878
R21973 XA.Cn[8].n16 XA.Cn[8] 0.0309878
R21974 XA.Cn[8].n19 XA.Cn[8] 0.0309878
R21975 XA.Cn[8].n22 XA.Cn[8] 0.0309878
R21976 XA.Cn[8].n25 XA.Cn[8] 0.0309878
R21977 XA.Cn[8].n28 XA.Cn[8] 0.0309878
R21978 XA.Cn[8].n31 XA.Cn[8] 0.0309878
R21979 XA.Cn[8].n34 XA.Cn[8] 0.0309878
R21980 XA.Cn[8].n37 XA.Cn[8] 0.0309878
R21981 XA.Cn[8].n40 XA.Cn[8] 0.0309878
R21982 XA.Cn[8].n43 XA.Cn[8] 0.0309878
R21983 XA.Cn[8].n46 XA.Cn[8] 0.0309878
R21984 XA.Cn[8].n49 XA.Cn[8] 0.0309878
R21985 XA.Cn[8].n5 XA.Cn[8].n4 0.027939
R21986 XA.Cn[8].n8 XA.Cn[8].n7 0.027939
R21987 XA.Cn[8].n11 XA.Cn[8].n10 0.027939
R21988 XA.Cn[8].n14 XA.Cn[8].n13 0.027939
R21989 XA.Cn[8].n17 XA.Cn[8].n16 0.027939
R21990 XA.Cn[8].n20 XA.Cn[8].n19 0.027939
R21991 XA.Cn[8].n23 XA.Cn[8].n22 0.027939
R21992 XA.Cn[8].n26 XA.Cn[8].n25 0.027939
R21993 XA.Cn[8].n29 XA.Cn[8].n28 0.027939
R21994 XA.Cn[8].n32 XA.Cn[8].n31 0.027939
R21995 XA.Cn[8].n35 XA.Cn[8].n34 0.027939
R21996 XA.Cn[8].n38 XA.Cn[8].n37 0.027939
R21997 XA.Cn[8].n41 XA.Cn[8].n40 0.027939
R21998 XA.Cn[8].n44 XA.Cn[8].n43 0.027939
R21999 XA.Cn[8].n47 XA.Cn[8].n46 0.027939
R22000 XA.Cn[8].n50 XA.Cn[8].n49 0.027939
R22001 XThR.Tn[1].n2 XThR.Tn[1].n1 332.332
R22002 XThR.Tn[1].n2 XThR.Tn[1].n0 296.493
R22003 XThR.Tn[1] XThR.Tn[1].n82 161.363
R22004 XThR.Tn[1] XThR.Tn[1].n77 161.363
R22005 XThR.Tn[1] XThR.Tn[1].n72 161.363
R22006 XThR.Tn[1] XThR.Tn[1].n67 161.363
R22007 XThR.Tn[1] XThR.Tn[1].n62 161.363
R22008 XThR.Tn[1] XThR.Tn[1].n57 161.363
R22009 XThR.Tn[1] XThR.Tn[1].n52 161.363
R22010 XThR.Tn[1] XThR.Tn[1].n47 161.363
R22011 XThR.Tn[1] XThR.Tn[1].n42 161.363
R22012 XThR.Tn[1] XThR.Tn[1].n37 161.363
R22013 XThR.Tn[1] XThR.Tn[1].n32 161.363
R22014 XThR.Tn[1] XThR.Tn[1].n27 161.363
R22015 XThR.Tn[1] XThR.Tn[1].n22 161.363
R22016 XThR.Tn[1] XThR.Tn[1].n17 161.363
R22017 XThR.Tn[1] XThR.Tn[1].n12 161.363
R22018 XThR.Tn[1] XThR.Tn[1].n10 161.363
R22019 XThR.Tn[1].n84 XThR.Tn[1].n83 161.3
R22020 XThR.Tn[1].n79 XThR.Tn[1].n78 161.3
R22021 XThR.Tn[1].n74 XThR.Tn[1].n73 161.3
R22022 XThR.Tn[1].n69 XThR.Tn[1].n68 161.3
R22023 XThR.Tn[1].n64 XThR.Tn[1].n63 161.3
R22024 XThR.Tn[1].n59 XThR.Tn[1].n58 161.3
R22025 XThR.Tn[1].n54 XThR.Tn[1].n53 161.3
R22026 XThR.Tn[1].n49 XThR.Tn[1].n48 161.3
R22027 XThR.Tn[1].n44 XThR.Tn[1].n43 161.3
R22028 XThR.Tn[1].n39 XThR.Tn[1].n38 161.3
R22029 XThR.Tn[1].n34 XThR.Tn[1].n33 161.3
R22030 XThR.Tn[1].n29 XThR.Tn[1].n28 161.3
R22031 XThR.Tn[1].n24 XThR.Tn[1].n23 161.3
R22032 XThR.Tn[1].n19 XThR.Tn[1].n18 161.3
R22033 XThR.Tn[1].n14 XThR.Tn[1].n13 161.3
R22034 XThR.Tn[1].n82 XThR.Tn[1].t70 161.106
R22035 XThR.Tn[1].n77 XThR.Tn[1].t14 161.106
R22036 XThR.Tn[1].n72 XThR.Tn[1].t56 161.106
R22037 XThR.Tn[1].n67 XThR.Tn[1].t42 161.106
R22038 XThR.Tn[1].n62 XThR.Tn[1].t68 161.106
R22039 XThR.Tn[1].n57 XThR.Tn[1].t31 161.106
R22040 XThR.Tn[1].n52 XThR.Tn[1].t12 161.106
R22041 XThR.Tn[1].n47 XThR.Tn[1].t54 161.106
R22042 XThR.Tn[1].n42 XThR.Tn[1].t41 161.106
R22043 XThR.Tn[1].n37 XThR.Tn[1].t46 161.106
R22044 XThR.Tn[1].n32 XThR.Tn[1].t29 161.106
R22045 XThR.Tn[1].n27 XThR.Tn[1].t55 161.106
R22046 XThR.Tn[1].n22 XThR.Tn[1].t28 161.106
R22047 XThR.Tn[1].n17 XThR.Tn[1].t73 161.106
R22048 XThR.Tn[1].n12 XThR.Tn[1].t34 161.106
R22049 XThR.Tn[1].n10 XThR.Tn[1].t18 161.106
R22050 XThR.Tn[1].n83 XThR.Tn[1].t66 159.978
R22051 XThR.Tn[1].n78 XThR.Tn[1].t72 159.978
R22052 XThR.Tn[1].n73 XThR.Tn[1].t52 159.978
R22053 XThR.Tn[1].n68 XThR.Tn[1].t39 159.978
R22054 XThR.Tn[1].n63 XThR.Tn[1].t63 159.978
R22055 XThR.Tn[1].n58 XThR.Tn[1].t27 159.978
R22056 XThR.Tn[1].n53 XThR.Tn[1].t71 159.978
R22057 XThR.Tn[1].n48 XThR.Tn[1].t49 159.978
R22058 XThR.Tn[1].n43 XThR.Tn[1].t36 159.978
R22059 XThR.Tn[1].n38 XThR.Tn[1].t43 159.978
R22060 XThR.Tn[1].n33 XThR.Tn[1].t26 159.978
R22061 XThR.Tn[1].n28 XThR.Tn[1].t51 159.978
R22062 XThR.Tn[1].n23 XThR.Tn[1].t25 159.978
R22063 XThR.Tn[1].n18 XThR.Tn[1].t69 159.978
R22064 XThR.Tn[1].n13 XThR.Tn[1].t30 159.978
R22065 XThR.Tn[1].n82 XThR.Tn[1].t58 145.038
R22066 XThR.Tn[1].n77 XThR.Tn[1].t20 145.038
R22067 XThR.Tn[1].n72 XThR.Tn[1].t62 145.038
R22068 XThR.Tn[1].n67 XThR.Tn[1].t47 145.038
R22069 XThR.Tn[1].n62 XThR.Tn[1].t15 145.038
R22070 XThR.Tn[1].n57 XThR.Tn[1].t57 145.038
R22071 XThR.Tn[1].n52 XThR.Tn[1].t64 145.038
R22072 XThR.Tn[1].n47 XThR.Tn[1].t48 145.038
R22073 XThR.Tn[1].n42 XThR.Tn[1].t45 145.038
R22074 XThR.Tn[1].n37 XThR.Tn[1].t13 145.038
R22075 XThR.Tn[1].n32 XThR.Tn[1].t37 145.038
R22076 XThR.Tn[1].n27 XThR.Tn[1].t59 145.038
R22077 XThR.Tn[1].n22 XThR.Tn[1].t35 145.038
R22078 XThR.Tn[1].n17 XThR.Tn[1].t19 145.038
R22079 XThR.Tn[1].n12 XThR.Tn[1].t44 145.038
R22080 XThR.Tn[1].n10 XThR.Tn[1].t24 145.038
R22081 XThR.Tn[1].n83 XThR.Tn[1].t17 143.911
R22082 XThR.Tn[1].n78 XThR.Tn[1].t40 143.911
R22083 XThR.Tn[1].n73 XThR.Tn[1].t22 143.911
R22084 XThR.Tn[1].n68 XThR.Tn[1].t65 143.911
R22085 XThR.Tn[1].n63 XThR.Tn[1].t33 143.911
R22086 XThR.Tn[1].n58 XThR.Tn[1].t16 143.911
R22087 XThR.Tn[1].n53 XThR.Tn[1].t23 143.911
R22088 XThR.Tn[1].n48 XThR.Tn[1].t67 143.911
R22089 XThR.Tn[1].n43 XThR.Tn[1].t60 143.911
R22090 XThR.Tn[1].n38 XThR.Tn[1].t32 143.911
R22091 XThR.Tn[1].n33 XThR.Tn[1].t53 143.911
R22092 XThR.Tn[1].n28 XThR.Tn[1].t21 143.911
R22093 XThR.Tn[1].n23 XThR.Tn[1].t50 143.911
R22094 XThR.Tn[1].n18 XThR.Tn[1].t38 143.911
R22095 XThR.Tn[1].n13 XThR.Tn[1].t61 143.911
R22096 XThR.Tn[1].n7 XThR.Tn[1].n6 135.249
R22097 XThR.Tn[1].n9 XThR.Tn[1].n3 98.981
R22098 XThR.Tn[1].n8 XThR.Tn[1].n4 98.981
R22099 XThR.Tn[1].n7 XThR.Tn[1].n5 98.981
R22100 XThR.Tn[1].n9 XThR.Tn[1].n8 36.2672
R22101 XThR.Tn[1].n8 XThR.Tn[1].n7 36.2672
R22102 XThR.Tn[1].n88 XThR.Tn[1].n9 32.6405
R22103 XThR.Tn[1].n1 XThR.Tn[1].t7 26.5955
R22104 XThR.Tn[1].n1 XThR.Tn[1].t6 26.5955
R22105 XThR.Tn[1].n0 XThR.Tn[1].t4 26.5955
R22106 XThR.Tn[1].n0 XThR.Tn[1].t5 26.5955
R22107 XThR.Tn[1].n3 XThR.Tn[1].t11 24.9236
R22108 XThR.Tn[1].n3 XThR.Tn[1].t8 24.9236
R22109 XThR.Tn[1].n4 XThR.Tn[1].t10 24.9236
R22110 XThR.Tn[1].n4 XThR.Tn[1].t9 24.9236
R22111 XThR.Tn[1].n5 XThR.Tn[1].t2 24.9236
R22112 XThR.Tn[1].n5 XThR.Tn[1].t1 24.9236
R22113 XThR.Tn[1].n6 XThR.Tn[1].t3 24.9236
R22114 XThR.Tn[1].n6 XThR.Tn[1].t0 24.9236
R22115 XThR.Tn[1].n89 XThR.Tn[1].n2 18.5605
R22116 XThR.Tn[1].n89 XThR.Tn[1].n88 11.5205
R22117 XThR.Tn[1].n88 XThR.Tn[1] 6.42118
R22118 XThR.Tn[1] XThR.Tn[1].n11 5.34038
R22119 XThR.Tn[1].n16 XThR.Tn[1].n15 4.5005
R22120 XThR.Tn[1].n21 XThR.Tn[1].n20 4.5005
R22121 XThR.Tn[1].n26 XThR.Tn[1].n25 4.5005
R22122 XThR.Tn[1].n31 XThR.Tn[1].n30 4.5005
R22123 XThR.Tn[1].n36 XThR.Tn[1].n35 4.5005
R22124 XThR.Tn[1].n41 XThR.Tn[1].n40 4.5005
R22125 XThR.Tn[1].n46 XThR.Tn[1].n45 4.5005
R22126 XThR.Tn[1].n51 XThR.Tn[1].n50 4.5005
R22127 XThR.Tn[1].n56 XThR.Tn[1].n55 4.5005
R22128 XThR.Tn[1].n61 XThR.Tn[1].n60 4.5005
R22129 XThR.Tn[1].n66 XThR.Tn[1].n65 4.5005
R22130 XThR.Tn[1].n71 XThR.Tn[1].n70 4.5005
R22131 XThR.Tn[1].n76 XThR.Tn[1].n75 4.5005
R22132 XThR.Tn[1].n81 XThR.Tn[1].n80 4.5005
R22133 XThR.Tn[1].n86 XThR.Tn[1].n85 4.5005
R22134 XThR.Tn[1].n87 XThR.Tn[1] 3.70586
R22135 XThR.Tn[1].n16 XThR.Tn[1] 2.52282
R22136 XThR.Tn[1].n21 XThR.Tn[1] 2.52282
R22137 XThR.Tn[1].n26 XThR.Tn[1] 2.52282
R22138 XThR.Tn[1].n31 XThR.Tn[1] 2.52282
R22139 XThR.Tn[1].n36 XThR.Tn[1] 2.52282
R22140 XThR.Tn[1].n41 XThR.Tn[1] 2.52282
R22141 XThR.Tn[1].n46 XThR.Tn[1] 2.52282
R22142 XThR.Tn[1].n51 XThR.Tn[1] 2.52282
R22143 XThR.Tn[1].n56 XThR.Tn[1] 2.52282
R22144 XThR.Tn[1].n61 XThR.Tn[1] 2.52282
R22145 XThR.Tn[1].n66 XThR.Tn[1] 2.52282
R22146 XThR.Tn[1].n71 XThR.Tn[1] 2.52282
R22147 XThR.Tn[1].n76 XThR.Tn[1] 2.52282
R22148 XThR.Tn[1].n81 XThR.Tn[1] 2.52282
R22149 XThR.Tn[1].n86 XThR.Tn[1] 2.52282
R22150 XThR.Tn[1].n84 XThR.Tn[1] 1.08677
R22151 XThR.Tn[1].n79 XThR.Tn[1] 1.08677
R22152 XThR.Tn[1].n74 XThR.Tn[1] 1.08677
R22153 XThR.Tn[1].n69 XThR.Tn[1] 1.08677
R22154 XThR.Tn[1].n64 XThR.Tn[1] 1.08677
R22155 XThR.Tn[1].n59 XThR.Tn[1] 1.08677
R22156 XThR.Tn[1].n54 XThR.Tn[1] 1.08677
R22157 XThR.Tn[1].n49 XThR.Tn[1] 1.08677
R22158 XThR.Tn[1].n44 XThR.Tn[1] 1.08677
R22159 XThR.Tn[1].n39 XThR.Tn[1] 1.08677
R22160 XThR.Tn[1].n34 XThR.Tn[1] 1.08677
R22161 XThR.Tn[1].n29 XThR.Tn[1] 1.08677
R22162 XThR.Tn[1].n24 XThR.Tn[1] 1.08677
R22163 XThR.Tn[1].n19 XThR.Tn[1] 1.08677
R22164 XThR.Tn[1].n14 XThR.Tn[1] 1.08677
R22165 XThR.Tn[1] XThR.Tn[1].n16 0.839786
R22166 XThR.Tn[1] XThR.Tn[1].n21 0.839786
R22167 XThR.Tn[1] XThR.Tn[1].n26 0.839786
R22168 XThR.Tn[1] XThR.Tn[1].n31 0.839786
R22169 XThR.Tn[1] XThR.Tn[1].n36 0.839786
R22170 XThR.Tn[1] XThR.Tn[1].n41 0.839786
R22171 XThR.Tn[1] XThR.Tn[1].n46 0.839786
R22172 XThR.Tn[1] XThR.Tn[1].n51 0.839786
R22173 XThR.Tn[1] XThR.Tn[1].n56 0.839786
R22174 XThR.Tn[1] XThR.Tn[1].n61 0.839786
R22175 XThR.Tn[1] XThR.Tn[1].n66 0.839786
R22176 XThR.Tn[1] XThR.Tn[1].n71 0.839786
R22177 XThR.Tn[1] XThR.Tn[1].n76 0.839786
R22178 XThR.Tn[1] XThR.Tn[1].n81 0.839786
R22179 XThR.Tn[1] XThR.Tn[1].n86 0.839786
R22180 XThR.Tn[1] XThR.Tn[1].n89 0.6405
R22181 XThR.Tn[1].n11 XThR.Tn[1] 0.499542
R22182 XThR.Tn[1].n85 XThR.Tn[1] 0.063
R22183 XThR.Tn[1].n80 XThR.Tn[1] 0.063
R22184 XThR.Tn[1].n75 XThR.Tn[1] 0.063
R22185 XThR.Tn[1].n70 XThR.Tn[1] 0.063
R22186 XThR.Tn[1].n65 XThR.Tn[1] 0.063
R22187 XThR.Tn[1].n60 XThR.Tn[1] 0.063
R22188 XThR.Tn[1].n55 XThR.Tn[1] 0.063
R22189 XThR.Tn[1].n50 XThR.Tn[1] 0.063
R22190 XThR.Tn[1].n45 XThR.Tn[1] 0.063
R22191 XThR.Tn[1].n40 XThR.Tn[1] 0.063
R22192 XThR.Tn[1].n35 XThR.Tn[1] 0.063
R22193 XThR.Tn[1].n30 XThR.Tn[1] 0.063
R22194 XThR.Tn[1].n25 XThR.Tn[1] 0.063
R22195 XThR.Tn[1].n20 XThR.Tn[1] 0.063
R22196 XThR.Tn[1].n15 XThR.Tn[1] 0.063
R22197 XThR.Tn[1].n87 XThR.Tn[1] 0.0540714
R22198 XThR.Tn[1] XThR.Tn[1].n87 0.038
R22199 XThR.Tn[1].n11 XThR.Tn[1] 0.0143889
R22200 XThR.Tn[1].n85 XThR.Tn[1].n84 0.00771154
R22201 XThR.Tn[1].n80 XThR.Tn[1].n79 0.00771154
R22202 XThR.Tn[1].n75 XThR.Tn[1].n74 0.00771154
R22203 XThR.Tn[1].n70 XThR.Tn[1].n69 0.00771154
R22204 XThR.Tn[1].n65 XThR.Tn[1].n64 0.00771154
R22205 XThR.Tn[1].n60 XThR.Tn[1].n59 0.00771154
R22206 XThR.Tn[1].n55 XThR.Tn[1].n54 0.00771154
R22207 XThR.Tn[1].n50 XThR.Tn[1].n49 0.00771154
R22208 XThR.Tn[1].n45 XThR.Tn[1].n44 0.00771154
R22209 XThR.Tn[1].n40 XThR.Tn[1].n39 0.00771154
R22210 XThR.Tn[1].n35 XThR.Tn[1].n34 0.00771154
R22211 XThR.Tn[1].n30 XThR.Tn[1].n29 0.00771154
R22212 XThR.Tn[1].n25 XThR.Tn[1].n24 0.00771154
R22213 XThR.Tn[1].n20 XThR.Tn[1].n19 0.00771154
R22214 XThR.Tn[1].n15 XThR.Tn[1].n14 0.00771154
R22215 XA.Cn[7].n5 XA.Cn[7].n4 255.096
R22216 XA.Cn[7].n2 XA.Cn[7].n0 236.589
R22217 XA.Cn[7].n5 XA.Cn[7].n3 201.845
R22218 XA.Cn[7].n2 XA.Cn[7].n1 200.321
R22219 XA.Cn[7].n8 XA.Cn[7].n6 161.406
R22220 XA.Cn[7].n11 XA.Cn[7].n9 161.406
R22221 XA.Cn[7].n14 XA.Cn[7].n12 161.406
R22222 XA.Cn[7].n17 XA.Cn[7].n15 161.406
R22223 XA.Cn[7].n20 XA.Cn[7].n18 161.406
R22224 XA.Cn[7].n23 XA.Cn[7].n21 161.406
R22225 XA.Cn[7].n26 XA.Cn[7].n24 161.406
R22226 XA.Cn[7].n29 XA.Cn[7].n27 161.406
R22227 XA.Cn[7].n32 XA.Cn[7].n30 161.406
R22228 XA.Cn[7].n35 XA.Cn[7].n33 161.406
R22229 XA.Cn[7].n38 XA.Cn[7].n36 161.406
R22230 XA.Cn[7].n41 XA.Cn[7].n39 161.406
R22231 XA.Cn[7].n44 XA.Cn[7].n42 161.406
R22232 XA.Cn[7].n47 XA.Cn[7].n45 161.406
R22233 XA.Cn[7].n50 XA.Cn[7].n48 161.406
R22234 XA.Cn[7].n53 XA.Cn[7].n51 161.406
R22235 XA.Cn[7].n6 XA.Cn[7].t11 161.202
R22236 XA.Cn[7].n9 XA.Cn[7].t30 161.202
R22237 XA.Cn[7].n12 XA.Cn[7].t34 161.202
R22238 XA.Cn[7].n15 XA.Cn[7].t35 161.202
R22239 XA.Cn[7].n18 XA.Cn[7].t22 161.202
R22240 XA.Cn[7].n21 XA.Cn[7].t23 161.202
R22241 XA.Cn[7].n24 XA.Cn[7].t39 161.202
R22242 XA.Cn[7].n27 XA.Cn[7].t14 161.202
R22243 XA.Cn[7].n30 XA.Cn[7].t16 161.202
R22244 XA.Cn[7].n33 XA.Cn[7].t36 161.202
R22245 XA.Cn[7].n36 XA.Cn[7].t38 161.202
R22246 XA.Cn[7].n39 XA.Cn[7].t17 161.202
R22247 XA.Cn[7].n42 XA.Cn[7].t26 161.202
R22248 XA.Cn[7].n45 XA.Cn[7].t28 161.202
R22249 XA.Cn[7].n48 XA.Cn[7].t9 161.202
R22250 XA.Cn[7].n51 XA.Cn[7].t19 161.202
R22251 XA.Cn[7].n6 XA.Cn[7].t8 145.137
R22252 XA.Cn[7].n9 XA.Cn[7].t25 145.137
R22253 XA.Cn[7].n12 XA.Cn[7].t27 145.137
R22254 XA.Cn[7].n15 XA.Cn[7].t29 145.137
R22255 XA.Cn[7].n18 XA.Cn[7].t18 145.137
R22256 XA.Cn[7].n21 XA.Cn[7].t20 145.137
R22257 XA.Cn[7].n24 XA.Cn[7].t33 145.137
R22258 XA.Cn[7].n27 XA.Cn[7].t10 145.137
R22259 XA.Cn[7].n30 XA.Cn[7].t12 145.137
R22260 XA.Cn[7].n33 XA.Cn[7].t31 145.137
R22261 XA.Cn[7].n36 XA.Cn[7].t32 145.137
R22262 XA.Cn[7].n39 XA.Cn[7].t13 145.137
R22263 XA.Cn[7].n42 XA.Cn[7].t21 145.137
R22264 XA.Cn[7].n45 XA.Cn[7].t24 145.137
R22265 XA.Cn[7].n48 XA.Cn[7].t37 145.137
R22266 XA.Cn[7].n51 XA.Cn[7].t15 145.137
R22267 XA.Cn[7].n4 XA.Cn[7].t2 26.5955
R22268 XA.Cn[7].n4 XA.Cn[7].t1 26.5955
R22269 XA.Cn[7].n3 XA.Cn[7].t0 26.5955
R22270 XA.Cn[7].n3 XA.Cn[7].t3 26.5955
R22271 XA.Cn[7] XA.Cn[7].n5 26.4992
R22272 XA.Cn[7].n0 XA.Cn[7].t6 24.9236
R22273 XA.Cn[7].n0 XA.Cn[7].t5 24.9236
R22274 XA.Cn[7].n1 XA.Cn[7].t4 24.9236
R22275 XA.Cn[7].n1 XA.Cn[7].t7 24.9236
R22276 XA.Cn[7].n56 XA.Cn[7].n2 12.0894
R22277 XA.Cn[7].n56 XA.Cn[7] 9.64206
R22278 XA.Cn[7].n55 XA.Cn[7] 8.14595
R22279 XA.Cn[7].n55 XA.Cn[7].n54 3.36239
R22280 XA.Cn[7] XA.Cn[7].n55 3.15894
R22281 XA.Cn[7].n54 XA.Cn[7] 2.07622
R22282 XA.Cn[7] XA.Cn[7].n56 1.66284
R22283 XA.Cn[7].n11 XA.Cn[7] 0.931056
R22284 XA.Cn[7].n14 XA.Cn[7] 0.931056
R22285 XA.Cn[7].n17 XA.Cn[7] 0.931056
R22286 XA.Cn[7].n20 XA.Cn[7] 0.931056
R22287 XA.Cn[7].n23 XA.Cn[7] 0.931056
R22288 XA.Cn[7].n26 XA.Cn[7] 0.931056
R22289 XA.Cn[7].n29 XA.Cn[7] 0.931056
R22290 XA.Cn[7].n32 XA.Cn[7] 0.931056
R22291 XA.Cn[7].n35 XA.Cn[7] 0.931056
R22292 XA.Cn[7].n38 XA.Cn[7] 0.931056
R22293 XA.Cn[7].n41 XA.Cn[7] 0.931056
R22294 XA.Cn[7].n44 XA.Cn[7] 0.931056
R22295 XA.Cn[7].n47 XA.Cn[7] 0.931056
R22296 XA.Cn[7].n50 XA.Cn[7] 0.931056
R22297 XA.Cn[7].n53 XA.Cn[7] 0.931056
R22298 XA.Cn[7] XA.Cn[7].n8 0.396333
R22299 XA.Cn[7] XA.Cn[7].n11 0.396333
R22300 XA.Cn[7] XA.Cn[7].n14 0.396333
R22301 XA.Cn[7] XA.Cn[7].n17 0.396333
R22302 XA.Cn[7] XA.Cn[7].n20 0.396333
R22303 XA.Cn[7] XA.Cn[7].n23 0.396333
R22304 XA.Cn[7] XA.Cn[7].n26 0.396333
R22305 XA.Cn[7] XA.Cn[7].n29 0.396333
R22306 XA.Cn[7] XA.Cn[7].n32 0.396333
R22307 XA.Cn[7] XA.Cn[7].n35 0.396333
R22308 XA.Cn[7] XA.Cn[7].n38 0.396333
R22309 XA.Cn[7] XA.Cn[7].n41 0.396333
R22310 XA.Cn[7] XA.Cn[7].n44 0.396333
R22311 XA.Cn[7] XA.Cn[7].n47 0.396333
R22312 XA.Cn[7] XA.Cn[7].n50 0.396333
R22313 XA.Cn[7] XA.Cn[7].n53 0.396333
R22314 XA.Cn[7].n7 XA.Cn[7] 0.104667
R22315 XA.Cn[7].n10 XA.Cn[7] 0.104667
R22316 XA.Cn[7].n13 XA.Cn[7] 0.104667
R22317 XA.Cn[7].n16 XA.Cn[7] 0.104667
R22318 XA.Cn[7].n19 XA.Cn[7] 0.104667
R22319 XA.Cn[7].n22 XA.Cn[7] 0.104667
R22320 XA.Cn[7].n25 XA.Cn[7] 0.104667
R22321 XA.Cn[7].n28 XA.Cn[7] 0.104667
R22322 XA.Cn[7].n31 XA.Cn[7] 0.104667
R22323 XA.Cn[7].n34 XA.Cn[7] 0.104667
R22324 XA.Cn[7].n37 XA.Cn[7] 0.104667
R22325 XA.Cn[7].n40 XA.Cn[7] 0.104667
R22326 XA.Cn[7].n43 XA.Cn[7] 0.104667
R22327 XA.Cn[7].n46 XA.Cn[7] 0.104667
R22328 XA.Cn[7].n49 XA.Cn[7] 0.104667
R22329 XA.Cn[7].n52 XA.Cn[7] 0.104667
R22330 XA.Cn[7].n7 XA.Cn[7] 0.0309878
R22331 XA.Cn[7].n10 XA.Cn[7] 0.0309878
R22332 XA.Cn[7].n13 XA.Cn[7] 0.0309878
R22333 XA.Cn[7].n16 XA.Cn[7] 0.0309878
R22334 XA.Cn[7].n19 XA.Cn[7] 0.0309878
R22335 XA.Cn[7].n22 XA.Cn[7] 0.0309878
R22336 XA.Cn[7].n25 XA.Cn[7] 0.0309878
R22337 XA.Cn[7].n28 XA.Cn[7] 0.0309878
R22338 XA.Cn[7].n31 XA.Cn[7] 0.0309878
R22339 XA.Cn[7].n34 XA.Cn[7] 0.0309878
R22340 XA.Cn[7].n37 XA.Cn[7] 0.0309878
R22341 XA.Cn[7].n40 XA.Cn[7] 0.0309878
R22342 XA.Cn[7].n43 XA.Cn[7] 0.0309878
R22343 XA.Cn[7].n46 XA.Cn[7] 0.0309878
R22344 XA.Cn[7].n49 XA.Cn[7] 0.0309878
R22345 XA.Cn[7].n52 XA.Cn[7] 0.0309878
R22346 XA.Cn[7].n8 XA.Cn[7].n7 0.027939
R22347 XA.Cn[7].n11 XA.Cn[7].n10 0.027939
R22348 XA.Cn[7].n14 XA.Cn[7].n13 0.027939
R22349 XA.Cn[7].n17 XA.Cn[7].n16 0.027939
R22350 XA.Cn[7].n20 XA.Cn[7].n19 0.027939
R22351 XA.Cn[7].n23 XA.Cn[7].n22 0.027939
R22352 XA.Cn[7].n26 XA.Cn[7].n25 0.027939
R22353 XA.Cn[7].n29 XA.Cn[7].n28 0.027939
R22354 XA.Cn[7].n32 XA.Cn[7].n31 0.027939
R22355 XA.Cn[7].n35 XA.Cn[7].n34 0.027939
R22356 XA.Cn[7].n38 XA.Cn[7].n37 0.027939
R22357 XA.Cn[7].n41 XA.Cn[7].n40 0.027939
R22358 XA.Cn[7].n44 XA.Cn[7].n43 0.027939
R22359 XA.Cn[7].n47 XA.Cn[7].n46 0.027939
R22360 XA.Cn[7].n50 XA.Cn[7].n49 0.027939
R22361 XA.Cn[7].n53 XA.Cn[7].n52 0.027939
R22362 XA.Cn[7].n54 XA.Cn[7] 0.00240908
R22363 XThR.Tn[4].n2 XThR.Tn[4].n1 332.332
R22364 XThR.Tn[4].n2 XThR.Tn[4].n0 296.493
R22365 XThR.Tn[4] XThR.Tn[4].n82 161.363
R22366 XThR.Tn[4] XThR.Tn[4].n77 161.363
R22367 XThR.Tn[4] XThR.Tn[4].n72 161.363
R22368 XThR.Tn[4] XThR.Tn[4].n67 161.363
R22369 XThR.Tn[4] XThR.Tn[4].n62 161.363
R22370 XThR.Tn[4] XThR.Tn[4].n57 161.363
R22371 XThR.Tn[4] XThR.Tn[4].n52 161.363
R22372 XThR.Tn[4] XThR.Tn[4].n47 161.363
R22373 XThR.Tn[4] XThR.Tn[4].n42 161.363
R22374 XThR.Tn[4] XThR.Tn[4].n37 161.363
R22375 XThR.Tn[4] XThR.Tn[4].n32 161.363
R22376 XThR.Tn[4] XThR.Tn[4].n27 161.363
R22377 XThR.Tn[4] XThR.Tn[4].n22 161.363
R22378 XThR.Tn[4] XThR.Tn[4].n17 161.363
R22379 XThR.Tn[4] XThR.Tn[4].n12 161.363
R22380 XThR.Tn[4] XThR.Tn[4].n10 161.363
R22381 XThR.Tn[4].n84 XThR.Tn[4].n83 161.3
R22382 XThR.Tn[4].n79 XThR.Tn[4].n78 161.3
R22383 XThR.Tn[4].n74 XThR.Tn[4].n73 161.3
R22384 XThR.Tn[4].n69 XThR.Tn[4].n68 161.3
R22385 XThR.Tn[4].n64 XThR.Tn[4].n63 161.3
R22386 XThR.Tn[4].n59 XThR.Tn[4].n58 161.3
R22387 XThR.Tn[4].n54 XThR.Tn[4].n53 161.3
R22388 XThR.Tn[4].n49 XThR.Tn[4].n48 161.3
R22389 XThR.Tn[4].n44 XThR.Tn[4].n43 161.3
R22390 XThR.Tn[4].n39 XThR.Tn[4].n38 161.3
R22391 XThR.Tn[4].n34 XThR.Tn[4].n33 161.3
R22392 XThR.Tn[4].n29 XThR.Tn[4].n28 161.3
R22393 XThR.Tn[4].n24 XThR.Tn[4].n23 161.3
R22394 XThR.Tn[4].n19 XThR.Tn[4].n18 161.3
R22395 XThR.Tn[4].n14 XThR.Tn[4].n13 161.3
R22396 XThR.Tn[4].n82 XThR.Tn[4].t28 161.106
R22397 XThR.Tn[4].n77 XThR.Tn[4].t34 161.106
R22398 XThR.Tn[4].n72 XThR.Tn[4].t14 161.106
R22399 XThR.Tn[4].n67 XThR.Tn[4].t62 161.106
R22400 XThR.Tn[4].n62 XThR.Tn[4].t26 161.106
R22401 XThR.Tn[4].n57 XThR.Tn[4].t51 161.106
R22402 XThR.Tn[4].n52 XThR.Tn[4].t32 161.106
R22403 XThR.Tn[4].n47 XThR.Tn[4].t12 161.106
R22404 XThR.Tn[4].n42 XThR.Tn[4].t61 161.106
R22405 XThR.Tn[4].n37 XThR.Tn[4].t66 161.106
R22406 XThR.Tn[4].n32 XThR.Tn[4].t49 161.106
R22407 XThR.Tn[4].n27 XThR.Tn[4].t13 161.106
R22408 XThR.Tn[4].n22 XThR.Tn[4].t48 161.106
R22409 XThR.Tn[4].n17 XThR.Tn[4].t31 161.106
R22410 XThR.Tn[4].n12 XThR.Tn[4].t54 161.106
R22411 XThR.Tn[4].n10 XThR.Tn[4].t38 161.106
R22412 XThR.Tn[4].n83 XThR.Tn[4].t24 159.978
R22413 XThR.Tn[4].n78 XThR.Tn[4].t30 159.978
R22414 XThR.Tn[4].n73 XThR.Tn[4].t72 159.978
R22415 XThR.Tn[4].n68 XThR.Tn[4].t59 159.978
R22416 XThR.Tn[4].n63 XThR.Tn[4].t21 159.978
R22417 XThR.Tn[4].n58 XThR.Tn[4].t47 159.978
R22418 XThR.Tn[4].n53 XThR.Tn[4].t29 159.978
R22419 XThR.Tn[4].n48 XThR.Tn[4].t69 159.978
R22420 XThR.Tn[4].n43 XThR.Tn[4].t56 159.978
R22421 XThR.Tn[4].n38 XThR.Tn[4].t63 159.978
R22422 XThR.Tn[4].n33 XThR.Tn[4].t46 159.978
R22423 XThR.Tn[4].n28 XThR.Tn[4].t71 159.978
R22424 XThR.Tn[4].n23 XThR.Tn[4].t45 159.978
R22425 XThR.Tn[4].n18 XThR.Tn[4].t27 159.978
R22426 XThR.Tn[4].n13 XThR.Tn[4].t50 159.978
R22427 XThR.Tn[4].n82 XThR.Tn[4].t16 145.038
R22428 XThR.Tn[4].n77 XThR.Tn[4].t40 145.038
R22429 XThR.Tn[4].n72 XThR.Tn[4].t20 145.038
R22430 XThR.Tn[4].n67 XThR.Tn[4].t67 145.038
R22431 XThR.Tn[4].n62 XThR.Tn[4].t35 145.038
R22432 XThR.Tn[4].n57 XThR.Tn[4].t15 145.038
R22433 XThR.Tn[4].n52 XThR.Tn[4].t22 145.038
R22434 XThR.Tn[4].n47 XThR.Tn[4].t68 145.038
R22435 XThR.Tn[4].n42 XThR.Tn[4].t64 145.038
R22436 XThR.Tn[4].n37 XThR.Tn[4].t33 145.038
R22437 XThR.Tn[4].n32 XThR.Tn[4].t57 145.038
R22438 XThR.Tn[4].n27 XThR.Tn[4].t17 145.038
R22439 XThR.Tn[4].n22 XThR.Tn[4].t55 145.038
R22440 XThR.Tn[4].n17 XThR.Tn[4].t39 145.038
R22441 XThR.Tn[4].n12 XThR.Tn[4].t65 145.038
R22442 XThR.Tn[4].n10 XThR.Tn[4].t44 145.038
R22443 XThR.Tn[4].n83 XThR.Tn[4].t37 143.911
R22444 XThR.Tn[4].n78 XThR.Tn[4].t60 143.911
R22445 XThR.Tn[4].n73 XThR.Tn[4].t42 143.911
R22446 XThR.Tn[4].n68 XThR.Tn[4].t23 143.911
R22447 XThR.Tn[4].n63 XThR.Tn[4].t53 143.911
R22448 XThR.Tn[4].n58 XThR.Tn[4].t36 143.911
R22449 XThR.Tn[4].n53 XThR.Tn[4].t43 143.911
R22450 XThR.Tn[4].n48 XThR.Tn[4].t25 143.911
R22451 XThR.Tn[4].n43 XThR.Tn[4].t18 143.911
R22452 XThR.Tn[4].n38 XThR.Tn[4].t52 143.911
R22453 XThR.Tn[4].n33 XThR.Tn[4].t73 143.911
R22454 XThR.Tn[4].n28 XThR.Tn[4].t41 143.911
R22455 XThR.Tn[4].n23 XThR.Tn[4].t70 143.911
R22456 XThR.Tn[4].n18 XThR.Tn[4].t58 143.911
R22457 XThR.Tn[4].n13 XThR.Tn[4].t19 143.911
R22458 XThR.Tn[4].n7 XThR.Tn[4].n5 135.249
R22459 XThR.Tn[4].n9 XThR.Tn[4].n3 98.982
R22460 XThR.Tn[4].n8 XThR.Tn[4].n4 98.982
R22461 XThR.Tn[4].n7 XThR.Tn[4].n6 98.982
R22462 XThR.Tn[4].n9 XThR.Tn[4].n8 36.2672
R22463 XThR.Tn[4].n8 XThR.Tn[4].n7 36.2672
R22464 XThR.Tn[4].n88 XThR.Tn[4].n9 32.6405
R22465 XThR.Tn[4].n1 XThR.Tn[4].t8 26.5955
R22466 XThR.Tn[4].n1 XThR.Tn[4].t11 26.5955
R22467 XThR.Tn[4].n0 XThR.Tn[4].t9 26.5955
R22468 XThR.Tn[4].n0 XThR.Tn[4].t10 26.5955
R22469 XThR.Tn[4].n3 XThR.Tn[4].t7 24.9236
R22470 XThR.Tn[4].n3 XThR.Tn[4].t4 24.9236
R22471 XThR.Tn[4].n4 XThR.Tn[4].t6 24.9236
R22472 XThR.Tn[4].n4 XThR.Tn[4].t5 24.9236
R22473 XThR.Tn[4].n5 XThR.Tn[4].t0 24.9236
R22474 XThR.Tn[4].n5 XThR.Tn[4].t1 24.9236
R22475 XThR.Tn[4].n6 XThR.Tn[4].t3 24.9236
R22476 XThR.Tn[4].n6 XThR.Tn[4].t2 24.9236
R22477 XThR.Tn[4] XThR.Tn[4].n2 23.3605
R22478 XThR.Tn[4] XThR.Tn[4].n88 6.7205
R22479 XThR.Tn[4].n88 XThR.Tn[4] 5.80883
R22480 XThR.Tn[4] XThR.Tn[4].n11 5.34038
R22481 XThR.Tn[4].n16 XThR.Tn[4].n15 4.5005
R22482 XThR.Tn[4].n21 XThR.Tn[4].n20 4.5005
R22483 XThR.Tn[4].n26 XThR.Tn[4].n25 4.5005
R22484 XThR.Tn[4].n31 XThR.Tn[4].n30 4.5005
R22485 XThR.Tn[4].n36 XThR.Tn[4].n35 4.5005
R22486 XThR.Tn[4].n41 XThR.Tn[4].n40 4.5005
R22487 XThR.Tn[4].n46 XThR.Tn[4].n45 4.5005
R22488 XThR.Tn[4].n51 XThR.Tn[4].n50 4.5005
R22489 XThR.Tn[4].n56 XThR.Tn[4].n55 4.5005
R22490 XThR.Tn[4].n61 XThR.Tn[4].n60 4.5005
R22491 XThR.Tn[4].n66 XThR.Tn[4].n65 4.5005
R22492 XThR.Tn[4].n71 XThR.Tn[4].n70 4.5005
R22493 XThR.Tn[4].n76 XThR.Tn[4].n75 4.5005
R22494 XThR.Tn[4].n81 XThR.Tn[4].n80 4.5005
R22495 XThR.Tn[4].n86 XThR.Tn[4].n85 4.5005
R22496 XThR.Tn[4].n87 XThR.Tn[4] 3.70586
R22497 XThR.Tn[4].n16 XThR.Tn[4] 2.52282
R22498 XThR.Tn[4].n21 XThR.Tn[4] 2.52282
R22499 XThR.Tn[4].n26 XThR.Tn[4] 2.52282
R22500 XThR.Tn[4].n31 XThR.Tn[4] 2.52282
R22501 XThR.Tn[4].n36 XThR.Tn[4] 2.52282
R22502 XThR.Tn[4].n41 XThR.Tn[4] 2.52282
R22503 XThR.Tn[4].n46 XThR.Tn[4] 2.52282
R22504 XThR.Tn[4].n51 XThR.Tn[4] 2.52282
R22505 XThR.Tn[4].n56 XThR.Tn[4] 2.52282
R22506 XThR.Tn[4].n61 XThR.Tn[4] 2.52282
R22507 XThR.Tn[4].n66 XThR.Tn[4] 2.52282
R22508 XThR.Tn[4].n71 XThR.Tn[4] 2.52282
R22509 XThR.Tn[4].n76 XThR.Tn[4] 2.52282
R22510 XThR.Tn[4].n81 XThR.Tn[4] 2.52282
R22511 XThR.Tn[4].n86 XThR.Tn[4] 2.52282
R22512 XThR.Tn[4].n84 XThR.Tn[4] 1.08677
R22513 XThR.Tn[4].n79 XThR.Tn[4] 1.08677
R22514 XThR.Tn[4].n74 XThR.Tn[4] 1.08677
R22515 XThR.Tn[4].n69 XThR.Tn[4] 1.08677
R22516 XThR.Tn[4].n64 XThR.Tn[4] 1.08677
R22517 XThR.Tn[4].n59 XThR.Tn[4] 1.08677
R22518 XThR.Tn[4].n54 XThR.Tn[4] 1.08677
R22519 XThR.Tn[4].n49 XThR.Tn[4] 1.08677
R22520 XThR.Tn[4].n44 XThR.Tn[4] 1.08677
R22521 XThR.Tn[4].n39 XThR.Tn[4] 1.08677
R22522 XThR.Tn[4].n34 XThR.Tn[4] 1.08677
R22523 XThR.Tn[4].n29 XThR.Tn[4] 1.08677
R22524 XThR.Tn[4].n24 XThR.Tn[4] 1.08677
R22525 XThR.Tn[4].n19 XThR.Tn[4] 1.08677
R22526 XThR.Tn[4].n14 XThR.Tn[4] 1.08677
R22527 XThR.Tn[4] XThR.Tn[4].n16 0.839786
R22528 XThR.Tn[4] XThR.Tn[4].n21 0.839786
R22529 XThR.Tn[4] XThR.Tn[4].n26 0.839786
R22530 XThR.Tn[4] XThR.Tn[4].n31 0.839786
R22531 XThR.Tn[4] XThR.Tn[4].n36 0.839786
R22532 XThR.Tn[4] XThR.Tn[4].n41 0.839786
R22533 XThR.Tn[4] XThR.Tn[4].n46 0.839786
R22534 XThR.Tn[4] XThR.Tn[4].n51 0.839786
R22535 XThR.Tn[4] XThR.Tn[4].n56 0.839786
R22536 XThR.Tn[4] XThR.Tn[4].n61 0.839786
R22537 XThR.Tn[4] XThR.Tn[4].n66 0.839786
R22538 XThR.Tn[4] XThR.Tn[4].n71 0.839786
R22539 XThR.Tn[4] XThR.Tn[4].n76 0.839786
R22540 XThR.Tn[4] XThR.Tn[4].n81 0.839786
R22541 XThR.Tn[4] XThR.Tn[4].n86 0.839786
R22542 XThR.Tn[4].n11 XThR.Tn[4] 0.499542
R22543 XThR.Tn[4].n85 XThR.Tn[4] 0.063
R22544 XThR.Tn[4].n80 XThR.Tn[4] 0.063
R22545 XThR.Tn[4].n75 XThR.Tn[4] 0.063
R22546 XThR.Tn[4].n70 XThR.Tn[4] 0.063
R22547 XThR.Tn[4].n65 XThR.Tn[4] 0.063
R22548 XThR.Tn[4].n60 XThR.Tn[4] 0.063
R22549 XThR.Tn[4].n55 XThR.Tn[4] 0.063
R22550 XThR.Tn[4].n50 XThR.Tn[4] 0.063
R22551 XThR.Tn[4].n45 XThR.Tn[4] 0.063
R22552 XThR.Tn[4].n40 XThR.Tn[4] 0.063
R22553 XThR.Tn[4].n35 XThR.Tn[4] 0.063
R22554 XThR.Tn[4].n30 XThR.Tn[4] 0.063
R22555 XThR.Tn[4].n25 XThR.Tn[4] 0.063
R22556 XThR.Tn[4].n20 XThR.Tn[4] 0.063
R22557 XThR.Tn[4].n15 XThR.Tn[4] 0.063
R22558 XThR.Tn[4].n87 XThR.Tn[4] 0.0540714
R22559 XThR.Tn[4] XThR.Tn[4].n87 0.038
R22560 XThR.Tn[4].n11 XThR.Tn[4] 0.0143889
R22561 XThR.Tn[4].n85 XThR.Tn[4].n84 0.00771154
R22562 XThR.Tn[4].n80 XThR.Tn[4].n79 0.00771154
R22563 XThR.Tn[4].n75 XThR.Tn[4].n74 0.00771154
R22564 XThR.Tn[4].n70 XThR.Tn[4].n69 0.00771154
R22565 XThR.Tn[4].n65 XThR.Tn[4].n64 0.00771154
R22566 XThR.Tn[4].n60 XThR.Tn[4].n59 0.00771154
R22567 XThR.Tn[4].n55 XThR.Tn[4].n54 0.00771154
R22568 XThR.Tn[4].n50 XThR.Tn[4].n49 0.00771154
R22569 XThR.Tn[4].n45 XThR.Tn[4].n44 0.00771154
R22570 XThR.Tn[4].n40 XThR.Tn[4].n39 0.00771154
R22571 XThR.Tn[4].n35 XThR.Tn[4].n34 0.00771154
R22572 XThR.Tn[4].n30 XThR.Tn[4].n29 0.00771154
R22573 XThR.Tn[4].n25 XThR.Tn[4].n24 0.00771154
R22574 XThR.Tn[4].n20 XThR.Tn[4].n19 0.00771154
R22575 XThR.Tn[4].n15 XThR.Tn[4].n14 0.00771154
R22576 XThR.Tn[11].n8 XThR.Tn[11].n7 256.104
R22577 XThR.Tn[11].n5 XThR.Tn[11].n3 243.68
R22578 XThR.Tn[11].n2 XThR.Tn[11].n1 241.847
R22579 XThR.Tn[11].n5 XThR.Tn[11].n4 205.28
R22580 XThR.Tn[11].n8 XThR.Tn[11].n6 202.094
R22581 XThR.Tn[11].n2 XThR.Tn[11].n0 185
R22582 XThR.Tn[11] XThR.Tn[11].n82 161.363
R22583 XThR.Tn[11] XThR.Tn[11].n77 161.363
R22584 XThR.Tn[11] XThR.Tn[11].n72 161.363
R22585 XThR.Tn[11] XThR.Tn[11].n67 161.363
R22586 XThR.Tn[11] XThR.Tn[11].n62 161.363
R22587 XThR.Tn[11] XThR.Tn[11].n57 161.363
R22588 XThR.Tn[11] XThR.Tn[11].n52 161.363
R22589 XThR.Tn[11] XThR.Tn[11].n47 161.363
R22590 XThR.Tn[11] XThR.Tn[11].n42 161.363
R22591 XThR.Tn[11] XThR.Tn[11].n37 161.363
R22592 XThR.Tn[11] XThR.Tn[11].n32 161.363
R22593 XThR.Tn[11] XThR.Tn[11].n27 161.363
R22594 XThR.Tn[11] XThR.Tn[11].n22 161.363
R22595 XThR.Tn[11] XThR.Tn[11].n17 161.363
R22596 XThR.Tn[11] XThR.Tn[11].n12 161.363
R22597 XThR.Tn[11] XThR.Tn[11].n10 161.363
R22598 XThR.Tn[11].n84 XThR.Tn[11].n83 161.3
R22599 XThR.Tn[11].n79 XThR.Tn[11].n78 161.3
R22600 XThR.Tn[11].n74 XThR.Tn[11].n73 161.3
R22601 XThR.Tn[11].n69 XThR.Tn[11].n68 161.3
R22602 XThR.Tn[11].n64 XThR.Tn[11].n63 161.3
R22603 XThR.Tn[11].n59 XThR.Tn[11].n58 161.3
R22604 XThR.Tn[11].n54 XThR.Tn[11].n53 161.3
R22605 XThR.Tn[11].n49 XThR.Tn[11].n48 161.3
R22606 XThR.Tn[11].n44 XThR.Tn[11].n43 161.3
R22607 XThR.Tn[11].n39 XThR.Tn[11].n38 161.3
R22608 XThR.Tn[11].n34 XThR.Tn[11].n33 161.3
R22609 XThR.Tn[11].n29 XThR.Tn[11].n28 161.3
R22610 XThR.Tn[11].n24 XThR.Tn[11].n23 161.3
R22611 XThR.Tn[11].n19 XThR.Tn[11].n18 161.3
R22612 XThR.Tn[11].n14 XThR.Tn[11].n13 161.3
R22613 XThR.Tn[11].n82 XThR.Tn[11].t40 161.106
R22614 XThR.Tn[11].n77 XThR.Tn[11].t46 161.106
R22615 XThR.Tn[11].n72 XThR.Tn[11].t24 161.106
R22616 XThR.Tn[11].n67 XThR.Tn[11].t73 161.106
R22617 XThR.Tn[11].n62 XThR.Tn[11].t39 161.106
R22618 XThR.Tn[11].n57 XThR.Tn[11].t63 161.106
R22619 XThR.Tn[11].n52 XThR.Tn[11].t43 161.106
R22620 XThR.Tn[11].n47 XThR.Tn[11].t22 161.106
R22621 XThR.Tn[11].n42 XThR.Tn[11].t71 161.106
R22622 XThR.Tn[11].n37 XThR.Tn[11].t14 161.106
R22623 XThR.Tn[11].n32 XThR.Tn[11].t62 161.106
R22624 XThR.Tn[11].n27 XThR.Tn[11].t23 161.106
R22625 XThR.Tn[11].n22 XThR.Tn[11].t60 161.106
R22626 XThR.Tn[11].n17 XThR.Tn[11].t41 161.106
R22627 XThR.Tn[11].n12 XThR.Tn[11].t67 161.106
R22628 XThR.Tn[11].n10 XThR.Tn[11].t48 161.106
R22629 XThR.Tn[11].n83 XThR.Tn[11].t31 159.978
R22630 XThR.Tn[11].n78 XThR.Tn[11].t38 159.978
R22631 XThR.Tn[11].n73 XThR.Tn[11].t20 159.978
R22632 XThR.Tn[11].n68 XThR.Tn[11].t66 159.978
R22633 XThR.Tn[11].n63 XThR.Tn[11].t29 159.978
R22634 XThR.Tn[11].n58 XThR.Tn[11].t57 159.978
R22635 XThR.Tn[11].n53 XThR.Tn[11].t37 159.978
R22636 XThR.Tn[11].n48 XThR.Tn[11].t17 159.978
R22637 XThR.Tn[11].n43 XThR.Tn[11].t64 159.978
R22638 XThR.Tn[11].n38 XThR.Tn[11].t72 159.978
R22639 XThR.Tn[11].n33 XThR.Tn[11].t55 159.978
R22640 XThR.Tn[11].n28 XThR.Tn[11].t19 159.978
R22641 XThR.Tn[11].n23 XThR.Tn[11].t54 159.978
R22642 XThR.Tn[11].n18 XThR.Tn[11].t36 159.978
R22643 XThR.Tn[11].n13 XThR.Tn[11].t58 159.978
R22644 XThR.Tn[11].n82 XThR.Tn[11].t26 145.038
R22645 XThR.Tn[11].n77 XThR.Tn[11].t53 145.038
R22646 XThR.Tn[11].n72 XThR.Tn[11].t34 145.038
R22647 XThR.Tn[11].n67 XThR.Tn[11].t15 145.038
R22648 XThR.Tn[11].n62 XThR.Tn[11].t47 145.038
R22649 XThR.Tn[11].n57 XThR.Tn[11].t25 145.038
R22650 XThR.Tn[11].n52 XThR.Tn[11].t35 145.038
R22651 XThR.Tn[11].n47 XThR.Tn[11].t16 145.038
R22652 XThR.Tn[11].n42 XThR.Tn[11].t13 145.038
R22653 XThR.Tn[11].n37 XThR.Tn[11].t44 145.038
R22654 XThR.Tn[11].n32 XThR.Tn[11].t70 145.038
R22655 XThR.Tn[11].n27 XThR.Tn[11].t33 145.038
R22656 XThR.Tn[11].n22 XThR.Tn[11].t68 145.038
R22657 XThR.Tn[11].n17 XThR.Tn[11].t49 145.038
R22658 XThR.Tn[11].n12 XThR.Tn[11].t12 145.038
R22659 XThR.Tn[11].n10 XThR.Tn[11].t56 145.038
R22660 XThR.Tn[11].n83 XThR.Tn[11].t45 143.911
R22661 XThR.Tn[11].n78 XThR.Tn[11].t69 143.911
R22662 XThR.Tn[11].n73 XThR.Tn[11].t51 143.911
R22663 XThR.Tn[11].n68 XThR.Tn[11].t30 143.911
R22664 XThR.Tn[11].n63 XThR.Tn[11].t61 143.911
R22665 XThR.Tn[11].n58 XThR.Tn[11].t42 143.911
R22666 XThR.Tn[11].n53 XThR.Tn[11].t52 143.911
R22667 XThR.Tn[11].n48 XThR.Tn[11].t32 143.911
R22668 XThR.Tn[11].n43 XThR.Tn[11].t28 143.911
R22669 XThR.Tn[11].n38 XThR.Tn[11].t59 143.911
R22670 XThR.Tn[11].n33 XThR.Tn[11].t21 143.911
R22671 XThR.Tn[11].n28 XThR.Tn[11].t50 143.911
R22672 XThR.Tn[11].n23 XThR.Tn[11].t18 143.911
R22673 XThR.Tn[11].n18 XThR.Tn[11].t65 143.911
R22674 XThR.Tn[11].n13 XThR.Tn[11].t27 143.911
R22675 XThR.Tn[11] XThR.Tn[11].n5 35.7652
R22676 XThR.Tn[11].n6 XThR.Tn[11].t3 26.5955
R22677 XThR.Tn[11].n6 XThR.Tn[11].t7 26.5955
R22678 XThR.Tn[11].n7 XThR.Tn[11].t1 26.5955
R22679 XThR.Tn[11].n7 XThR.Tn[11].t6 26.5955
R22680 XThR.Tn[11].n3 XThR.Tn[11].t8 26.5955
R22681 XThR.Tn[11].n3 XThR.Tn[11].t10 26.5955
R22682 XThR.Tn[11].n4 XThR.Tn[11].t9 26.5955
R22683 XThR.Tn[11].n4 XThR.Tn[11].t11 26.5955
R22684 XThR.Tn[11].n0 XThR.Tn[11].t5 24.9236
R22685 XThR.Tn[11].n0 XThR.Tn[11].t2 24.9236
R22686 XThR.Tn[11].n1 XThR.Tn[11].t4 24.9236
R22687 XThR.Tn[11].n1 XThR.Tn[11].t0 24.9236
R22688 XThR.Tn[11] XThR.Tn[11].n2 22.9615
R22689 XThR.Tn[11].n9 XThR.Tn[11].n8 13.5534
R22690 XThR.Tn[11].n88 XThR.Tn[11] 8.41462
R22691 XThR.Tn[11] XThR.Tn[11].n11 5.34038
R22692 XThR.Tn[11].n16 XThR.Tn[11].n15 4.5005
R22693 XThR.Tn[11].n21 XThR.Tn[11].n20 4.5005
R22694 XThR.Tn[11].n26 XThR.Tn[11].n25 4.5005
R22695 XThR.Tn[11].n31 XThR.Tn[11].n30 4.5005
R22696 XThR.Tn[11].n36 XThR.Tn[11].n35 4.5005
R22697 XThR.Tn[11].n41 XThR.Tn[11].n40 4.5005
R22698 XThR.Tn[11].n46 XThR.Tn[11].n45 4.5005
R22699 XThR.Tn[11].n51 XThR.Tn[11].n50 4.5005
R22700 XThR.Tn[11].n56 XThR.Tn[11].n55 4.5005
R22701 XThR.Tn[11].n61 XThR.Tn[11].n60 4.5005
R22702 XThR.Tn[11].n66 XThR.Tn[11].n65 4.5005
R22703 XThR.Tn[11].n71 XThR.Tn[11].n70 4.5005
R22704 XThR.Tn[11].n76 XThR.Tn[11].n75 4.5005
R22705 XThR.Tn[11].n81 XThR.Tn[11].n80 4.5005
R22706 XThR.Tn[11].n86 XThR.Tn[11].n85 4.5005
R22707 XThR.Tn[11].n87 XThR.Tn[11] 3.70586
R22708 XThR.Tn[11].n88 XThR.Tn[11].n9 2.99115
R22709 XThR.Tn[11].n9 XThR.Tn[11] 2.87153
R22710 XThR.Tn[11].n16 XThR.Tn[11] 2.52282
R22711 XThR.Tn[11].n21 XThR.Tn[11] 2.52282
R22712 XThR.Tn[11].n26 XThR.Tn[11] 2.52282
R22713 XThR.Tn[11].n31 XThR.Tn[11] 2.52282
R22714 XThR.Tn[11].n36 XThR.Tn[11] 2.52282
R22715 XThR.Tn[11].n41 XThR.Tn[11] 2.52282
R22716 XThR.Tn[11].n46 XThR.Tn[11] 2.52282
R22717 XThR.Tn[11].n51 XThR.Tn[11] 2.52282
R22718 XThR.Tn[11].n56 XThR.Tn[11] 2.52282
R22719 XThR.Tn[11].n61 XThR.Tn[11] 2.52282
R22720 XThR.Tn[11].n66 XThR.Tn[11] 2.52282
R22721 XThR.Tn[11].n71 XThR.Tn[11] 2.52282
R22722 XThR.Tn[11].n76 XThR.Tn[11] 2.52282
R22723 XThR.Tn[11].n81 XThR.Tn[11] 2.52282
R22724 XThR.Tn[11].n86 XThR.Tn[11] 2.52282
R22725 XThR.Tn[11] XThR.Tn[11].n88 2.2734
R22726 XThR.Tn[11].n9 XThR.Tn[11] 1.50638
R22727 XThR.Tn[11].n84 XThR.Tn[11] 1.08677
R22728 XThR.Tn[11].n79 XThR.Tn[11] 1.08677
R22729 XThR.Tn[11].n74 XThR.Tn[11] 1.08677
R22730 XThR.Tn[11].n69 XThR.Tn[11] 1.08677
R22731 XThR.Tn[11].n64 XThR.Tn[11] 1.08677
R22732 XThR.Tn[11].n59 XThR.Tn[11] 1.08677
R22733 XThR.Tn[11].n54 XThR.Tn[11] 1.08677
R22734 XThR.Tn[11].n49 XThR.Tn[11] 1.08677
R22735 XThR.Tn[11].n44 XThR.Tn[11] 1.08677
R22736 XThR.Tn[11].n39 XThR.Tn[11] 1.08677
R22737 XThR.Tn[11].n34 XThR.Tn[11] 1.08677
R22738 XThR.Tn[11].n29 XThR.Tn[11] 1.08677
R22739 XThR.Tn[11].n24 XThR.Tn[11] 1.08677
R22740 XThR.Tn[11].n19 XThR.Tn[11] 1.08677
R22741 XThR.Tn[11].n14 XThR.Tn[11] 1.08677
R22742 XThR.Tn[11] XThR.Tn[11].n16 0.839786
R22743 XThR.Tn[11] XThR.Tn[11].n21 0.839786
R22744 XThR.Tn[11] XThR.Tn[11].n26 0.839786
R22745 XThR.Tn[11] XThR.Tn[11].n31 0.839786
R22746 XThR.Tn[11] XThR.Tn[11].n36 0.839786
R22747 XThR.Tn[11] XThR.Tn[11].n41 0.839786
R22748 XThR.Tn[11] XThR.Tn[11].n46 0.839786
R22749 XThR.Tn[11] XThR.Tn[11].n51 0.839786
R22750 XThR.Tn[11] XThR.Tn[11].n56 0.839786
R22751 XThR.Tn[11] XThR.Tn[11].n61 0.839786
R22752 XThR.Tn[11] XThR.Tn[11].n66 0.839786
R22753 XThR.Tn[11] XThR.Tn[11].n71 0.839786
R22754 XThR.Tn[11] XThR.Tn[11].n76 0.839786
R22755 XThR.Tn[11] XThR.Tn[11].n81 0.839786
R22756 XThR.Tn[11] XThR.Tn[11].n86 0.839786
R22757 XThR.Tn[11].n11 XThR.Tn[11] 0.499542
R22758 XThR.Tn[11].n85 XThR.Tn[11] 0.063
R22759 XThR.Tn[11].n80 XThR.Tn[11] 0.063
R22760 XThR.Tn[11].n75 XThR.Tn[11] 0.063
R22761 XThR.Tn[11].n70 XThR.Tn[11] 0.063
R22762 XThR.Tn[11].n65 XThR.Tn[11] 0.063
R22763 XThR.Tn[11].n60 XThR.Tn[11] 0.063
R22764 XThR.Tn[11].n55 XThR.Tn[11] 0.063
R22765 XThR.Tn[11].n50 XThR.Tn[11] 0.063
R22766 XThR.Tn[11].n45 XThR.Tn[11] 0.063
R22767 XThR.Tn[11].n40 XThR.Tn[11] 0.063
R22768 XThR.Tn[11].n35 XThR.Tn[11] 0.063
R22769 XThR.Tn[11].n30 XThR.Tn[11] 0.063
R22770 XThR.Tn[11].n25 XThR.Tn[11] 0.063
R22771 XThR.Tn[11].n20 XThR.Tn[11] 0.063
R22772 XThR.Tn[11].n15 XThR.Tn[11] 0.063
R22773 XThR.Tn[11].n87 XThR.Tn[11] 0.0540714
R22774 XThR.Tn[11] XThR.Tn[11].n87 0.038
R22775 XThR.Tn[11].n11 XThR.Tn[11] 0.0143889
R22776 XThR.Tn[11].n85 XThR.Tn[11].n84 0.00771154
R22777 XThR.Tn[11].n80 XThR.Tn[11].n79 0.00771154
R22778 XThR.Tn[11].n75 XThR.Tn[11].n74 0.00771154
R22779 XThR.Tn[11].n70 XThR.Tn[11].n69 0.00771154
R22780 XThR.Tn[11].n65 XThR.Tn[11].n64 0.00771154
R22781 XThR.Tn[11].n60 XThR.Tn[11].n59 0.00771154
R22782 XThR.Tn[11].n55 XThR.Tn[11].n54 0.00771154
R22783 XThR.Tn[11].n50 XThR.Tn[11].n49 0.00771154
R22784 XThR.Tn[11].n45 XThR.Tn[11].n44 0.00771154
R22785 XThR.Tn[11].n40 XThR.Tn[11].n39 0.00771154
R22786 XThR.Tn[11].n35 XThR.Tn[11].n34 0.00771154
R22787 XThR.Tn[11].n30 XThR.Tn[11].n29 0.00771154
R22788 XThR.Tn[11].n25 XThR.Tn[11].n24 0.00771154
R22789 XThR.Tn[11].n20 XThR.Tn[11].n19 0.00771154
R22790 XThR.Tn[11].n15 XThR.Tn[11].n14 0.00771154
R22791 XThR.Tn[7].n5 XThR.Tn[7].n3 244.067
R22792 XThR.Tn[7].n2 XThR.Tn[7].n0 236.589
R22793 XThR.Tn[7].n5 XThR.Tn[7].n4 204.893
R22794 XThR.Tn[7].n2 XThR.Tn[7].n1 200.321
R22795 XThR.Tn[7] XThR.Tn[7].n79 161.363
R22796 XThR.Tn[7] XThR.Tn[7].n74 161.363
R22797 XThR.Tn[7] XThR.Tn[7].n69 161.363
R22798 XThR.Tn[7] XThR.Tn[7].n64 161.363
R22799 XThR.Tn[7] XThR.Tn[7].n59 161.363
R22800 XThR.Tn[7] XThR.Tn[7].n54 161.363
R22801 XThR.Tn[7] XThR.Tn[7].n49 161.363
R22802 XThR.Tn[7] XThR.Tn[7].n44 161.363
R22803 XThR.Tn[7] XThR.Tn[7].n39 161.363
R22804 XThR.Tn[7] XThR.Tn[7].n34 161.363
R22805 XThR.Tn[7] XThR.Tn[7].n29 161.363
R22806 XThR.Tn[7] XThR.Tn[7].n24 161.363
R22807 XThR.Tn[7] XThR.Tn[7].n19 161.363
R22808 XThR.Tn[7] XThR.Tn[7].n14 161.363
R22809 XThR.Tn[7] XThR.Tn[7].n9 161.363
R22810 XThR.Tn[7] XThR.Tn[7].n7 161.363
R22811 XThR.Tn[7].n81 XThR.Tn[7].n80 161.3
R22812 XThR.Tn[7].n76 XThR.Tn[7].n75 161.3
R22813 XThR.Tn[7].n71 XThR.Tn[7].n70 161.3
R22814 XThR.Tn[7].n66 XThR.Tn[7].n65 161.3
R22815 XThR.Tn[7].n61 XThR.Tn[7].n60 161.3
R22816 XThR.Tn[7].n56 XThR.Tn[7].n55 161.3
R22817 XThR.Tn[7].n51 XThR.Tn[7].n50 161.3
R22818 XThR.Tn[7].n46 XThR.Tn[7].n45 161.3
R22819 XThR.Tn[7].n41 XThR.Tn[7].n40 161.3
R22820 XThR.Tn[7].n36 XThR.Tn[7].n35 161.3
R22821 XThR.Tn[7].n31 XThR.Tn[7].n30 161.3
R22822 XThR.Tn[7].n26 XThR.Tn[7].n25 161.3
R22823 XThR.Tn[7].n21 XThR.Tn[7].n20 161.3
R22824 XThR.Tn[7].n16 XThR.Tn[7].n15 161.3
R22825 XThR.Tn[7].n11 XThR.Tn[7].n10 161.3
R22826 XThR.Tn[7].n79 XThR.Tn[7].t35 161.106
R22827 XThR.Tn[7].n74 XThR.Tn[7].t41 161.106
R22828 XThR.Tn[7].n69 XThR.Tn[7].t22 161.106
R22829 XThR.Tn[7].n64 XThR.Tn[7].t69 161.106
R22830 XThR.Tn[7].n59 XThR.Tn[7].t33 161.106
R22831 XThR.Tn[7].n54 XThR.Tn[7].t57 161.106
R22832 XThR.Tn[7].n49 XThR.Tn[7].t39 161.106
R22833 XThR.Tn[7].n44 XThR.Tn[7].t20 161.106
R22834 XThR.Tn[7].n39 XThR.Tn[7].t68 161.106
R22835 XThR.Tn[7].n34 XThR.Tn[7].t11 161.106
R22836 XThR.Tn[7].n29 XThR.Tn[7].t56 161.106
R22837 XThR.Tn[7].n24 XThR.Tn[7].t21 161.106
R22838 XThR.Tn[7].n19 XThR.Tn[7].t55 161.106
R22839 XThR.Tn[7].n14 XThR.Tn[7].t37 161.106
R22840 XThR.Tn[7].n9 XThR.Tn[7].t60 161.106
R22841 XThR.Tn[7].n7 XThR.Tn[7].t45 161.106
R22842 XThR.Tn[7].n80 XThR.Tn[7].t13 159.978
R22843 XThR.Tn[7].n75 XThR.Tn[7].t17 159.978
R22844 XThR.Tn[7].n70 XThR.Tn[7].t64 159.978
R22845 XThR.Tn[7].n65 XThR.Tn[7].t48 159.978
R22846 XThR.Tn[7].n60 XThR.Tn[7].t10 159.978
R22847 XThR.Tn[7].n55 XThR.Tn[7].t36 159.978
R22848 XThR.Tn[7].n50 XThR.Tn[7].t16 159.978
R22849 XThR.Tn[7].n45 XThR.Tn[7].t61 159.978
R22850 XThR.Tn[7].n40 XThR.Tn[7].t46 159.978
R22851 XThR.Tn[7].n35 XThR.Tn[7].t54 159.978
R22852 XThR.Tn[7].n30 XThR.Tn[7].t34 159.978
R22853 XThR.Tn[7].n25 XThR.Tn[7].t63 159.978
R22854 XThR.Tn[7].n20 XThR.Tn[7].t32 159.978
R22855 XThR.Tn[7].n15 XThR.Tn[7].t15 159.978
R22856 XThR.Tn[7].n10 XThR.Tn[7].t38 159.978
R22857 XThR.Tn[7].n79 XThR.Tn[7].t24 145.038
R22858 XThR.Tn[7].n74 XThR.Tn[7].t49 145.038
R22859 XThR.Tn[7].n69 XThR.Tn[7].t28 145.038
R22860 XThR.Tn[7].n64 XThR.Tn[7].t12 145.038
R22861 XThR.Tn[7].n59 XThR.Tn[7].t42 145.038
R22862 XThR.Tn[7].n54 XThR.Tn[7].t23 145.038
R22863 XThR.Tn[7].n49 XThR.Tn[7].t29 145.038
R22864 XThR.Tn[7].n44 XThR.Tn[7].t14 145.038
R22865 XThR.Tn[7].n39 XThR.Tn[7].t9 145.038
R22866 XThR.Tn[7].n34 XThR.Tn[7].t40 145.038
R22867 XThR.Tn[7].n29 XThR.Tn[7].t65 145.038
R22868 XThR.Tn[7].n24 XThR.Tn[7].t25 145.038
R22869 XThR.Tn[7].n19 XThR.Tn[7].t62 145.038
R22870 XThR.Tn[7].n14 XThR.Tn[7].t47 145.038
R22871 XThR.Tn[7].n9 XThR.Tn[7].t8 145.038
R22872 XThR.Tn[7].n7 XThR.Tn[7].t53 145.038
R22873 XThR.Tn[7].n80 XThR.Tn[7].t44 143.911
R22874 XThR.Tn[7].n75 XThR.Tn[7].t67 143.911
R22875 XThR.Tn[7].n70 XThR.Tn[7].t51 143.911
R22876 XThR.Tn[7].n65 XThR.Tn[7].t30 143.911
R22877 XThR.Tn[7].n60 XThR.Tn[7].t59 143.911
R22878 XThR.Tn[7].n55 XThR.Tn[7].t43 143.911
R22879 XThR.Tn[7].n50 XThR.Tn[7].t52 143.911
R22880 XThR.Tn[7].n45 XThR.Tn[7].t31 143.911
R22881 XThR.Tn[7].n40 XThR.Tn[7].t27 143.911
R22882 XThR.Tn[7].n35 XThR.Tn[7].t58 143.911
R22883 XThR.Tn[7].n30 XThR.Tn[7].t19 143.911
R22884 XThR.Tn[7].n25 XThR.Tn[7].t50 143.911
R22885 XThR.Tn[7].n20 XThR.Tn[7].t18 143.911
R22886 XThR.Tn[7].n15 XThR.Tn[7].t66 143.911
R22887 XThR.Tn[7].n10 XThR.Tn[7].t26 143.911
R22888 XThR.Tn[7].n4 XThR.Tn[7].t1 26.5955
R22889 XThR.Tn[7].n4 XThR.Tn[7].t0 26.5955
R22890 XThR.Tn[7].n3 XThR.Tn[7].t2 26.5955
R22891 XThR.Tn[7].n3 XThR.Tn[7].t3 26.5955
R22892 XThR.Tn[7].n0 XThR.Tn[7].t7 24.9236
R22893 XThR.Tn[7].n0 XThR.Tn[7].t4 24.9236
R22894 XThR.Tn[7].n1 XThR.Tn[7].t6 24.9236
R22895 XThR.Tn[7].n1 XThR.Tn[7].t5 24.9236
R22896 XThR.Tn[7] XThR.Tn[7].n2 16.079
R22897 XThR.Tn[7].n6 XThR.Tn[7].n5 11.4531
R22898 XThR.Tn[7] XThR.Tn[7].n6 10.4732
R22899 XThR.Tn[7] XThR.Tn[7].n85 8.81089
R22900 XThR.Tn[7] XThR.Tn[7].n8 5.34038
R22901 XThR.Tn[7].n85 XThR.Tn[7] 5.25732
R22902 XThR.Tn[7].n13 XThR.Tn[7].n12 4.5005
R22903 XThR.Tn[7].n18 XThR.Tn[7].n17 4.5005
R22904 XThR.Tn[7].n23 XThR.Tn[7].n22 4.5005
R22905 XThR.Tn[7].n28 XThR.Tn[7].n27 4.5005
R22906 XThR.Tn[7].n33 XThR.Tn[7].n32 4.5005
R22907 XThR.Tn[7].n38 XThR.Tn[7].n37 4.5005
R22908 XThR.Tn[7].n43 XThR.Tn[7].n42 4.5005
R22909 XThR.Tn[7].n48 XThR.Tn[7].n47 4.5005
R22910 XThR.Tn[7].n53 XThR.Tn[7].n52 4.5005
R22911 XThR.Tn[7].n58 XThR.Tn[7].n57 4.5005
R22912 XThR.Tn[7].n63 XThR.Tn[7].n62 4.5005
R22913 XThR.Tn[7].n68 XThR.Tn[7].n67 4.5005
R22914 XThR.Tn[7].n73 XThR.Tn[7].n72 4.5005
R22915 XThR.Tn[7].n78 XThR.Tn[7].n77 4.5005
R22916 XThR.Tn[7].n83 XThR.Tn[7].n82 4.5005
R22917 XThR.Tn[7].n84 XThR.Tn[7] 3.70586
R22918 XThR.Tn[7].n13 XThR.Tn[7] 2.52282
R22919 XThR.Tn[7].n18 XThR.Tn[7] 2.52282
R22920 XThR.Tn[7].n23 XThR.Tn[7] 2.52282
R22921 XThR.Tn[7].n28 XThR.Tn[7] 2.52282
R22922 XThR.Tn[7].n33 XThR.Tn[7] 2.52282
R22923 XThR.Tn[7].n38 XThR.Tn[7] 2.52282
R22924 XThR.Tn[7].n43 XThR.Tn[7] 2.52282
R22925 XThR.Tn[7].n48 XThR.Tn[7] 2.52282
R22926 XThR.Tn[7].n53 XThR.Tn[7] 2.52282
R22927 XThR.Tn[7].n58 XThR.Tn[7] 2.52282
R22928 XThR.Tn[7].n63 XThR.Tn[7] 2.52282
R22929 XThR.Tn[7].n68 XThR.Tn[7] 2.52282
R22930 XThR.Tn[7].n73 XThR.Tn[7] 2.52282
R22931 XThR.Tn[7].n78 XThR.Tn[7] 2.52282
R22932 XThR.Tn[7].n83 XThR.Tn[7] 2.52282
R22933 XThR.Tn[7].n85 XThR.Tn[7] 2.49401
R22934 XThR.Tn[7].n81 XThR.Tn[7] 1.08677
R22935 XThR.Tn[7].n76 XThR.Tn[7] 1.08677
R22936 XThR.Tn[7].n71 XThR.Tn[7] 1.08677
R22937 XThR.Tn[7].n66 XThR.Tn[7] 1.08677
R22938 XThR.Tn[7].n61 XThR.Tn[7] 1.08677
R22939 XThR.Tn[7].n56 XThR.Tn[7] 1.08677
R22940 XThR.Tn[7].n51 XThR.Tn[7] 1.08677
R22941 XThR.Tn[7].n46 XThR.Tn[7] 1.08677
R22942 XThR.Tn[7].n41 XThR.Tn[7] 1.08677
R22943 XThR.Tn[7].n36 XThR.Tn[7] 1.08677
R22944 XThR.Tn[7].n31 XThR.Tn[7] 1.08677
R22945 XThR.Tn[7].n26 XThR.Tn[7] 1.08677
R22946 XThR.Tn[7].n21 XThR.Tn[7] 1.08677
R22947 XThR.Tn[7].n16 XThR.Tn[7] 1.08677
R22948 XThR.Tn[7].n11 XThR.Tn[7] 1.08677
R22949 XThR.Tn[7] XThR.Tn[7].n13 0.839786
R22950 XThR.Tn[7] XThR.Tn[7].n18 0.839786
R22951 XThR.Tn[7] XThR.Tn[7].n23 0.839786
R22952 XThR.Tn[7] XThR.Tn[7].n28 0.839786
R22953 XThR.Tn[7] XThR.Tn[7].n33 0.839786
R22954 XThR.Tn[7] XThR.Tn[7].n38 0.839786
R22955 XThR.Tn[7] XThR.Tn[7].n43 0.839786
R22956 XThR.Tn[7] XThR.Tn[7].n48 0.839786
R22957 XThR.Tn[7] XThR.Tn[7].n53 0.839786
R22958 XThR.Tn[7] XThR.Tn[7].n58 0.839786
R22959 XThR.Tn[7] XThR.Tn[7].n63 0.839786
R22960 XThR.Tn[7] XThR.Tn[7].n68 0.839786
R22961 XThR.Tn[7] XThR.Tn[7].n73 0.839786
R22962 XThR.Tn[7] XThR.Tn[7].n78 0.839786
R22963 XThR.Tn[7] XThR.Tn[7].n83 0.839786
R22964 XThR.Tn[7].n6 XThR.Tn[7] 0.830612
R22965 XThR.Tn[7].n8 XThR.Tn[7] 0.499542
R22966 XThR.Tn[7].n82 XThR.Tn[7] 0.063
R22967 XThR.Tn[7].n77 XThR.Tn[7] 0.063
R22968 XThR.Tn[7].n72 XThR.Tn[7] 0.063
R22969 XThR.Tn[7].n67 XThR.Tn[7] 0.063
R22970 XThR.Tn[7].n62 XThR.Tn[7] 0.063
R22971 XThR.Tn[7].n57 XThR.Tn[7] 0.063
R22972 XThR.Tn[7].n52 XThR.Tn[7] 0.063
R22973 XThR.Tn[7].n47 XThR.Tn[7] 0.063
R22974 XThR.Tn[7].n42 XThR.Tn[7] 0.063
R22975 XThR.Tn[7].n37 XThR.Tn[7] 0.063
R22976 XThR.Tn[7].n32 XThR.Tn[7] 0.063
R22977 XThR.Tn[7].n27 XThR.Tn[7] 0.063
R22978 XThR.Tn[7].n22 XThR.Tn[7] 0.063
R22979 XThR.Tn[7].n17 XThR.Tn[7] 0.063
R22980 XThR.Tn[7].n12 XThR.Tn[7] 0.063
R22981 XThR.Tn[7].n84 XThR.Tn[7] 0.0540714
R22982 XThR.Tn[7] XThR.Tn[7].n84 0.038
R22983 XThR.Tn[7].n8 XThR.Tn[7] 0.0143889
R22984 XThR.Tn[7].n82 XThR.Tn[7].n81 0.00771154
R22985 XThR.Tn[7].n77 XThR.Tn[7].n76 0.00771154
R22986 XThR.Tn[7].n72 XThR.Tn[7].n71 0.00771154
R22987 XThR.Tn[7].n67 XThR.Tn[7].n66 0.00771154
R22988 XThR.Tn[7].n62 XThR.Tn[7].n61 0.00771154
R22989 XThR.Tn[7].n57 XThR.Tn[7].n56 0.00771154
R22990 XThR.Tn[7].n52 XThR.Tn[7].n51 0.00771154
R22991 XThR.Tn[7].n47 XThR.Tn[7].n46 0.00771154
R22992 XThR.Tn[7].n42 XThR.Tn[7].n41 0.00771154
R22993 XThR.Tn[7].n37 XThR.Tn[7].n36 0.00771154
R22994 XThR.Tn[7].n32 XThR.Tn[7].n31 0.00771154
R22995 XThR.Tn[7].n27 XThR.Tn[7].n26 0.00771154
R22996 XThR.Tn[7].n22 XThR.Tn[7].n21 0.00771154
R22997 XThR.Tn[7].n17 XThR.Tn[7].n16 0.00771154
R22998 XThR.Tn[7].n12 XThR.Tn[7].n11 0.00771154
R22999 XThR.Tn[0].n2 XThR.Tn[0].n1 332.332
R23000 XThR.Tn[0].n2 XThR.Tn[0].n0 296.493
R23001 XThR.Tn[0] XThR.Tn[0].n82 161.363
R23002 XThR.Tn[0] XThR.Tn[0].n77 161.363
R23003 XThR.Tn[0] XThR.Tn[0].n72 161.363
R23004 XThR.Tn[0] XThR.Tn[0].n67 161.363
R23005 XThR.Tn[0] XThR.Tn[0].n62 161.363
R23006 XThR.Tn[0] XThR.Tn[0].n57 161.363
R23007 XThR.Tn[0] XThR.Tn[0].n52 161.363
R23008 XThR.Tn[0] XThR.Tn[0].n47 161.363
R23009 XThR.Tn[0] XThR.Tn[0].n42 161.363
R23010 XThR.Tn[0] XThR.Tn[0].n37 161.363
R23011 XThR.Tn[0] XThR.Tn[0].n32 161.363
R23012 XThR.Tn[0] XThR.Tn[0].n27 161.363
R23013 XThR.Tn[0] XThR.Tn[0].n22 161.363
R23014 XThR.Tn[0] XThR.Tn[0].n17 161.363
R23015 XThR.Tn[0] XThR.Tn[0].n12 161.363
R23016 XThR.Tn[0] XThR.Tn[0].n10 161.363
R23017 XThR.Tn[0].n84 XThR.Tn[0].n83 161.3
R23018 XThR.Tn[0].n79 XThR.Tn[0].n78 161.3
R23019 XThR.Tn[0].n74 XThR.Tn[0].n73 161.3
R23020 XThR.Tn[0].n69 XThR.Tn[0].n68 161.3
R23021 XThR.Tn[0].n64 XThR.Tn[0].n63 161.3
R23022 XThR.Tn[0].n59 XThR.Tn[0].n58 161.3
R23023 XThR.Tn[0].n54 XThR.Tn[0].n53 161.3
R23024 XThR.Tn[0].n49 XThR.Tn[0].n48 161.3
R23025 XThR.Tn[0].n44 XThR.Tn[0].n43 161.3
R23026 XThR.Tn[0].n39 XThR.Tn[0].n38 161.3
R23027 XThR.Tn[0].n34 XThR.Tn[0].n33 161.3
R23028 XThR.Tn[0].n29 XThR.Tn[0].n28 161.3
R23029 XThR.Tn[0].n24 XThR.Tn[0].n23 161.3
R23030 XThR.Tn[0].n19 XThR.Tn[0].n18 161.3
R23031 XThR.Tn[0].n14 XThR.Tn[0].n13 161.3
R23032 XThR.Tn[0].n82 XThR.Tn[0].t32 161.106
R23033 XThR.Tn[0].n77 XThR.Tn[0].t36 161.106
R23034 XThR.Tn[0].n72 XThR.Tn[0].t16 161.106
R23035 XThR.Tn[0].n67 XThR.Tn[0].t65 161.106
R23036 XThR.Tn[0].n62 XThR.Tn[0].t31 161.106
R23037 XThR.Tn[0].n57 XThR.Tn[0].t53 161.106
R23038 XThR.Tn[0].n52 XThR.Tn[0].t34 161.106
R23039 XThR.Tn[0].n47 XThR.Tn[0].t14 161.106
R23040 XThR.Tn[0].n42 XThR.Tn[0].t63 161.106
R23041 XThR.Tn[0].n37 XThR.Tn[0].t68 161.106
R23042 XThR.Tn[0].n32 XThR.Tn[0].t52 161.106
R23043 XThR.Tn[0].n27 XThR.Tn[0].t15 161.106
R23044 XThR.Tn[0].n22 XThR.Tn[0].t51 161.106
R23045 XThR.Tn[0].n17 XThR.Tn[0].t33 161.106
R23046 XThR.Tn[0].n12 XThR.Tn[0].t58 161.106
R23047 XThR.Tn[0].n10 XThR.Tn[0].t40 161.106
R23048 XThR.Tn[0].n83 XThR.Tn[0].t20 159.978
R23049 XThR.Tn[0].n78 XThR.Tn[0].t30 159.978
R23050 XThR.Tn[0].n73 XThR.Tn[0].t73 159.978
R23051 XThR.Tn[0].n68 XThR.Tn[0].t57 159.978
R23052 XThR.Tn[0].n63 XThR.Tn[0].t19 159.978
R23053 XThR.Tn[0].n58 XThR.Tn[0].t49 159.978
R23054 XThR.Tn[0].n53 XThR.Tn[0].t29 159.978
R23055 XThR.Tn[0].n48 XThR.Tn[0].t71 159.978
R23056 XThR.Tn[0].n43 XThR.Tn[0].t55 159.978
R23057 XThR.Tn[0].n38 XThR.Tn[0].t64 159.978
R23058 XThR.Tn[0].n33 XThR.Tn[0].t46 159.978
R23059 XThR.Tn[0].n28 XThR.Tn[0].t72 159.978
R23060 XThR.Tn[0].n23 XThR.Tn[0].t44 159.978
R23061 XThR.Tn[0].n18 XThR.Tn[0].t26 159.978
R23062 XThR.Tn[0].n13 XThR.Tn[0].t50 159.978
R23063 XThR.Tn[0].n82 XThR.Tn[0].t18 145.038
R23064 XThR.Tn[0].n77 XThR.Tn[0].t42 145.038
R23065 XThR.Tn[0].n72 XThR.Tn[0].t22 145.038
R23066 XThR.Tn[0].n67 XThR.Tn[0].t69 145.038
R23067 XThR.Tn[0].n62 XThR.Tn[0].t37 145.038
R23068 XThR.Tn[0].n57 XThR.Tn[0].t17 145.038
R23069 XThR.Tn[0].n52 XThR.Tn[0].t25 145.038
R23070 XThR.Tn[0].n47 XThR.Tn[0].t70 145.038
R23071 XThR.Tn[0].n42 XThR.Tn[0].t66 145.038
R23072 XThR.Tn[0].n37 XThR.Tn[0].t35 145.038
R23073 XThR.Tn[0].n32 XThR.Tn[0].t60 145.038
R23074 XThR.Tn[0].n27 XThR.Tn[0].t21 145.038
R23075 XThR.Tn[0].n22 XThR.Tn[0].t59 145.038
R23076 XThR.Tn[0].n17 XThR.Tn[0].t41 145.038
R23077 XThR.Tn[0].n12 XThR.Tn[0].t67 145.038
R23078 XThR.Tn[0].n10 XThR.Tn[0].t48 145.038
R23079 XThR.Tn[0].n83 XThR.Tn[0].t39 143.911
R23080 XThR.Tn[0].n78 XThR.Tn[0].t62 143.911
R23081 XThR.Tn[0].n73 XThR.Tn[0].t45 143.911
R23082 XThR.Tn[0].n68 XThR.Tn[0].t27 143.911
R23083 XThR.Tn[0].n63 XThR.Tn[0].t56 143.911
R23084 XThR.Tn[0].n58 XThR.Tn[0].t38 143.911
R23085 XThR.Tn[0].n53 XThR.Tn[0].t47 143.911
R23086 XThR.Tn[0].n48 XThR.Tn[0].t28 143.911
R23087 XThR.Tn[0].n43 XThR.Tn[0].t23 143.911
R23088 XThR.Tn[0].n38 XThR.Tn[0].t54 143.911
R23089 XThR.Tn[0].n33 XThR.Tn[0].t13 143.911
R23090 XThR.Tn[0].n28 XThR.Tn[0].t43 143.911
R23091 XThR.Tn[0].n23 XThR.Tn[0].t12 143.911
R23092 XThR.Tn[0].n18 XThR.Tn[0].t61 143.911
R23093 XThR.Tn[0].n13 XThR.Tn[0].t24 143.911
R23094 XThR.Tn[0].n7 XThR.Tn[0].n5 135.249
R23095 XThR.Tn[0].n9 XThR.Tn[0].n3 98.982
R23096 XThR.Tn[0].n8 XThR.Tn[0].n4 98.982
R23097 XThR.Tn[0].n7 XThR.Tn[0].n6 98.982
R23098 XThR.Tn[0].n9 XThR.Tn[0].n8 36.2672
R23099 XThR.Tn[0].n8 XThR.Tn[0].n7 36.2672
R23100 XThR.Tn[0].n88 XThR.Tn[0].n9 32.6405
R23101 XThR.Tn[0].n1 XThR.Tn[0].t5 26.5955
R23102 XThR.Tn[0].n1 XThR.Tn[0].t4 26.5955
R23103 XThR.Tn[0].n0 XThR.Tn[0].t6 26.5955
R23104 XThR.Tn[0].n0 XThR.Tn[0].t7 26.5955
R23105 XThR.Tn[0].n3 XThR.Tn[0].t9 24.9236
R23106 XThR.Tn[0].n3 XThR.Tn[0].t10 24.9236
R23107 XThR.Tn[0].n4 XThR.Tn[0].t8 24.9236
R23108 XThR.Tn[0].n4 XThR.Tn[0].t11 24.9236
R23109 XThR.Tn[0].n5 XThR.Tn[0].t1 24.9236
R23110 XThR.Tn[0].n5 XThR.Tn[0].t2 24.9236
R23111 XThR.Tn[0].n6 XThR.Tn[0].t0 24.9236
R23112 XThR.Tn[0].n6 XThR.Tn[0].t3 24.9236
R23113 XThR.Tn[0] XThR.Tn[0].n2 23.3605
R23114 XThR.Tn[0] XThR.Tn[0].n88 6.7205
R23115 XThR.Tn[0].n88 XThR.Tn[0] 6.36522
R23116 XThR.Tn[0] XThR.Tn[0].n11 5.34038
R23117 XThR.Tn[0].n16 XThR.Tn[0].n15 4.5005
R23118 XThR.Tn[0].n21 XThR.Tn[0].n20 4.5005
R23119 XThR.Tn[0].n26 XThR.Tn[0].n25 4.5005
R23120 XThR.Tn[0].n31 XThR.Tn[0].n30 4.5005
R23121 XThR.Tn[0].n36 XThR.Tn[0].n35 4.5005
R23122 XThR.Tn[0].n41 XThR.Tn[0].n40 4.5005
R23123 XThR.Tn[0].n46 XThR.Tn[0].n45 4.5005
R23124 XThR.Tn[0].n51 XThR.Tn[0].n50 4.5005
R23125 XThR.Tn[0].n56 XThR.Tn[0].n55 4.5005
R23126 XThR.Tn[0].n61 XThR.Tn[0].n60 4.5005
R23127 XThR.Tn[0].n66 XThR.Tn[0].n65 4.5005
R23128 XThR.Tn[0].n71 XThR.Tn[0].n70 4.5005
R23129 XThR.Tn[0].n76 XThR.Tn[0].n75 4.5005
R23130 XThR.Tn[0].n81 XThR.Tn[0].n80 4.5005
R23131 XThR.Tn[0].n86 XThR.Tn[0].n85 4.5005
R23132 XThR.Tn[0].n87 XThR.Tn[0] 3.70586
R23133 XThR.Tn[0].n16 XThR.Tn[0] 2.52282
R23134 XThR.Tn[0].n21 XThR.Tn[0] 2.52282
R23135 XThR.Tn[0].n26 XThR.Tn[0] 2.52282
R23136 XThR.Tn[0].n31 XThR.Tn[0] 2.52282
R23137 XThR.Tn[0].n36 XThR.Tn[0] 2.52282
R23138 XThR.Tn[0].n41 XThR.Tn[0] 2.52282
R23139 XThR.Tn[0].n46 XThR.Tn[0] 2.52282
R23140 XThR.Tn[0].n51 XThR.Tn[0] 2.52282
R23141 XThR.Tn[0].n56 XThR.Tn[0] 2.52282
R23142 XThR.Tn[0].n61 XThR.Tn[0] 2.52282
R23143 XThR.Tn[0].n66 XThR.Tn[0] 2.52282
R23144 XThR.Tn[0].n71 XThR.Tn[0] 2.52282
R23145 XThR.Tn[0].n76 XThR.Tn[0] 2.52282
R23146 XThR.Tn[0].n81 XThR.Tn[0] 2.52282
R23147 XThR.Tn[0].n86 XThR.Tn[0] 2.52282
R23148 XThR.Tn[0].n84 XThR.Tn[0] 1.08677
R23149 XThR.Tn[0].n79 XThR.Tn[0] 1.08677
R23150 XThR.Tn[0].n74 XThR.Tn[0] 1.08677
R23151 XThR.Tn[0].n69 XThR.Tn[0] 1.08677
R23152 XThR.Tn[0].n64 XThR.Tn[0] 1.08677
R23153 XThR.Tn[0].n59 XThR.Tn[0] 1.08677
R23154 XThR.Tn[0].n54 XThR.Tn[0] 1.08677
R23155 XThR.Tn[0].n49 XThR.Tn[0] 1.08677
R23156 XThR.Tn[0].n44 XThR.Tn[0] 1.08677
R23157 XThR.Tn[0].n39 XThR.Tn[0] 1.08677
R23158 XThR.Tn[0].n34 XThR.Tn[0] 1.08677
R23159 XThR.Tn[0].n29 XThR.Tn[0] 1.08677
R23160 XThR.Tn[0].n24 XThR.Tn[0] 1.08677
R23161 XThR.Tn[0].n19 XThR.Tn[0] 1.08677
R23162 XThR.Tn[0].n14 XThR.Tn[0] 1.08677
R23163 XThR.Tn[0] XThR.Tn[0].n16 0.839786
R23164 XThR.Tn[0] XThR.Tn[0].n21 0.839786
R23165 XThR.Tn[0] XThR.Tn[0].n26 0.839786
R23166 XThR.Tn[0] XThR.Tn[0].n31 0.839786
R23167 XThR.Tn[0] XThR.Tn[0].n36 0.839786
R23168 XThR.Tn[0] XThR.Tn[0].n41 0.839786
R23169 XThR.Tn[0] XThR.Tn[0].n46 0.839786
R23170 XThR.Tn[0] XThR.Tn[0].n51 0.839786
R23171 XThR.Tn[0] XThR.Tn[0].n56 0.839786
R23172 XThR.Tn[0] XThR.Tn[0].n61 0.839786
R23173 XThR.Tn[0] XThR.Tn[0].n66 0.839786
R23174 XThR.Tn[0] XThR.Tn[0].n71 0.839786
R23175 XThR.Tn[0] XThR.Tn[0].n76 0.839786
R23176 XThR.Tn[0] XThR.Tn[0].n81 0.839786
R23177 XThR.Tn[0] XThR.Tn[0].n86 0.839786
R23178 XThR.Tn[0].n11 XThR.Tn[0] 0.499542
R23179 XThR.Tn[0].n85 XThR.Tn[0] 0.063
R23180 XThR.Tn[0].n80 XThR.Tn[0] 0.063
R23181 XThR.Tn[0].n75 XThR.Tn[0] 0.063
R23182 XThR.Tn[0].n70 XThR.Tn[0] 0.063
R23183 XThR.Tn[0].n65 XThR.Tn[0] 0.063
R23184 XThR.Tn[0].n60 XThR.Tn[0] 0.063
R23185 XThR.Tn[0].n55 XThR.Tn[0] 0.063
R23186 XThR.Tn[0].n50 XThR.Tn[0] 0.063
R23187 XThR.Tn[0].n45 XThR.Tn[0] 0.063
R23188 XThR.Tn[0].n40 XThR.Tn[0] 0.063
R23189 XThR.Tn[0].n35 XThR.Tn[0] 0.063
R23190 XThR.Tn[0].n30 XThR.Tn[0] 0.063
R23191 XThR.Tn[0].n25 XThR.Tn[0] 0.063
R23192 XThR.Tn[0].n20 XThR.Tn[0] 0.063
R23193 XThR.Tn[0].n15 XThR.Tn[0] 0.063
R23194 XThR.Tn[0].n87 XThR.Tn[0] 0.0540714
R23195 XThR.Tn[0] XThR.Tn[0].n87 0.038
R23196 XThR.Tn[0].n11 XThR.Tn[0] 0.0143889
R23197 XThR.Tn[0].n85 XThR.Tn[0].n84 0.00771154
R23198 XThR.Tn[0].n80 XThR.Tn[0].n79 0.00771154
R23199 XThR.Tn[0].n75 XThR.Tn[0].n74 0.00771154
R23200 XThR.Tn[0].n70 XThR.Tn[0].n69 0.00771154
R23201 XThR.Tn[0].n65 XThR.Tn[0].n64 0.00771154
R23202 XThR.Tn[0].n60 XThR.Tn[0].n59 0.00771154
R23203 XThR.Tn[0].n55 XThR.Tn[0].n54 0.00771154
R23204 XThR.Tn[0].n50 XThR.Tn[0].n49 0.00771154
R23205 XThR.Tn[0].n45 XThR.Tn[0].n44 0.00771154
R23206 XThR.Tn[0].n40 XThR.Tn[0].n39 0.00771154
R23207 XThR.Tn[0].n35 XThR.Tn[0].n34 0.00771154
R23208 XThR.Tn[0].n30 XThR.Tn[0].n29 0.00771154
R23209 XThR.Tn[0].n25 XThR.Tn[0].n24 0.00771154
R23210 XThR.Tn[0].n20 XThR.Tn[0].n19 0.00771154
R23211 XThR.Tn[0].n15 XThR.Tn[0].n14 0.00771154
R23212 XThR.Tn[8].n87 XThR.Tn[8].n86 256.103
R23213 XThR.Tn[8].n2 XThR.Tn[8].n0 243.68
R23214 XThR.Tn[8].n5 XThR.Tn[8].n3 241.847
R23215 XThR.Tn[8].n2 XThR.Tn[8].n1 205.28
R23216 XThR.Tn[8].n87 XThR.Tn[8].n85 202.095
R23217 XThR.Tn[8].n5 XThR.Tn[8].n4 185
R23218 XThR.Tn[8] XThR.Tn[8].n78 161.363
R23219 XThR.Tn[8] XThR.Tn[8].n73 161.363
R23220 XThR.Tn[8] XThR.Tn[8].n68 161.363
R23221 XThR.Tn[8] XThR.Tn[8].n63 161.363
R23222 XThR.Tn[8] XThR.Tn[8].n58 161.363
R23223 XThR.Tn[8] XThR.Tn[8].n53 161.363
R23224 XThR.Tn[8] XThR.Tn[8].n48 161.363
R23225 XThR.Tn[8] XThR.Tn[8].n43 161.363
R23226 XThR.Tn[8] XThR.Tn[8].n38 161.363
R23227 XThR.Tn[8] XThR.Tn[8].n33 161.363
R23228 XThR.Tn[8] XThR.Tn[8].n28 161.363
R23229 XThR.Tn[8] XThR.Tn[8].n23 161.363
R23230 XThR.Tn[8] XThR.Tn[8].n18 161.363
R23231 XThR.Tn[8] XThR.Tn[8].n13 161.363
R23232 XThR.Tn[8] XThR.Tn[8].n8 161.363
R23233 XThR.Tn[8] XThR.Tn[8].n6 161.363
R23234 XThR.Tn[8].n80 XThR.Tn[8].n79 161.3
R23235 XThR.Tn[8].n75 XThR.Tn[8].n74 161.3
R23236 XThR.Tn[8].n70 XThR.Tn[8].n69 161.3
R23237 XThR.Tn[8].n65 XThR.Tn[8].n64 161.3
R23238 XThR.Tn[8].n60 XThR.Tn[8].n59 161.3
R23239 XThR.Tn[8].n55 XThR.Tn[8].n54 161.3
R23240 XThR.Tn[8].n50 XThR.Tn[8].n49 161.3
R23241 XThR.Tn[8].n45 XThR.Tn[8].n44 161.3
R23242 XThR.Tn[8].n40 XThR.Tn[8].n39 161.3
R23243 XThR.Tn[8].n35 XThR.Tn[8].n34 161.3
R23244 XThR.Tn[8].n30 XThR.Tn[8].n29 161.3
R23245 XThR.Tn[8].n25 XThR.Tn[8].n24 161.3
R23246 XThR.Tn[8].n20 XThR.Tn[8].n19 161.3
R23247 XThR.Tn[8].n15 XThR.Tn[8].n14 161.3
R23248 XThR.Tn[8].n10 XThR.Tn[8].n9 161.3
R23249 XThR.Tn[8].n78 XThR.Tn[8].t23 161.106
R23250 XThR.Tn[8].n73 XThR.Tn[8].t29 161.106
R23251 XThR.Tn[8].n68 XThR.Tn[8].t71 161.106
R23252 XThR.Tn[8].n63 XThR.Tn[8].t57 161.106
R23253 XThR.Tn[8].n58 XThR.Tn[8].t21 161.106
R23254 XThR.Tn[8].n53 XThR.Tn[8].t46 161.106
R23255 XThR.Tn[8].n48 XThR.Tn[8].t27 161.106
R23256 XThR.Tn[8].n43 XThR.Tn[8].t69 161.106
R23257 XThR.Tn[8].n38 XThR.Tn[8].t56 161.106
R23258 XThR.Tn[8].n33 XThR.Tn[8].t61 161.106
R23259 XThR.Tn[8].n28 XThR.Tn[8].t44 161.106
R23260 XThR.Tn[8].n23 XThR.Tn[8].t70 161.106
R23261 XThR.Tn[8].n18 XThR.Tn[8].t43 161.106
R23262 XThR.Tn[8].n13 XThR.Tn[8].t26 161.106
R23263 XThR.Tn[8].n8 XThR.Tn[8].t49 161.106
R23264 XThR.Tn[8].n6 XThR.Tn[8].t33 161.106
R23265 XThR.Tn[8].n79 XThR.Tn[8].t19 159.978
R23266 XThR.Tn[8].n74 XThR.Tn[8].t25 159.978
R23267 XThR.Tn[8].n69 XThR.Tn[8].t67 159.978
R23268 XThR.Tn[8].n64 XThR.Tn[8].t54 159.978
R23269 XThR.Tn[8].n59 XThR.Tn[8].t16 159.978
R23270 XThR.Tn[8].n54 XThR.Tn[8].t42 159.978
R23271 XThR.Tn[8].n49 XThR.Tn[8].t24 159.978
R23272 XThR.Tn[8].n44 XThR.Tn[8].t64 159.978
R23273 XThR.Tn[8].n39 XThR.Tn[8].t51 159.978
R23274 XThR.Tn[8].n34 XThR.Tn[8].t58 159.978
R23275 XThR.Tn[8].n29 XThR.Tn[8].t41 159.978
R23276 XThR.Tn[8].n24 XThR.Tn[8].t66 159.978
R23277 XThR.Tn[8].n19 XThR.Tn[8].t40 159.978
R23278 XThR.Tn[8].n14 XThR.Tn[8].t22 159.978
R23279 XThR.Tn[8].n9 XThR.Tn[8].t45 159.978
R23280 XThR.Tn[8].n78 XThR.Tn[8].t73 145.038
R23281 XThR.Tn[8].n73 XThR.Tn[8].t35 145.038
R23282 XThR.Tn[8].n68 XThR.Tn[8].t15 145.038
R23283 XThR.Tn[8].n63 XThR.Tn[8].t62 145.038
R23284 XThR.Tn[8].n58 XThR.Tn[8].t30 145.038
R23285 XThR.Tn[8].n53 XThR.Tn[8].t72 145.038
R23286 XThR.Tn[8].n48 XThR.Tn[8].t17 145.038
R23287 XThR.Tn[8].n43 XThR.Tn[8].t63 145.038
R23288 XThR.Tn[8].n38 XThR.Tn[8].t60 145.038
R23289 XThR.Tn[8].n33 XThR.Tn[8].t28 145.038
R23290 XThR.Tn[8].n28 XThR.Tn[8].t52 145.038
R23291 XThR.Tn[8].n23 XThR.Tn[8].t12 145.038
R23292 XThR.Tn[8].n18 XThR.Tn[8].t50 145.038
R23293 XThR.Tn[8].n13 XThR.Tn[8].t34 145.038
R23294 XThR.Tn[8].n8 XThR.Tn[8].t59 145.038
R23295 XThR.Tn[8].n6 XThR.Tn[8].t39 145.038
R23296 XThR.Tn[8].n79 XThR.Tn[8].t32 143.911
R23297 XThR.Tn[8].n74 XThR.Tn[8].t55 143.911
R23298 XThR.Tn[8].n69 XThR.Tn[8].t37 143.911
R23299 XThR.Tn[8].n64 XThR.Tn[8].t18 143.911
R23300 XThR.Tn[8].n59 XThR.Tn[8].t48 143.911
R23301 XThR.Tn[8].n54 XThR.Tn[8].t31 143.911
R23302 XThR.Tn[8].n49 XThR.Tn[8].t38 143.911
R23303 XThR.Tn[8].n44 XThR.Tn[8].t20 143.911
R23304 XThR.Tn[8].n39 XThR.Tn[8].t14 143.911
R23305 XThR.Tn[8].n34 XThR.Tn[8].t47 143.911
R23306 XThR.Tn[8].n29 XThR.Tn[8].t68 143.911
R23307 XThR.Tn[8].n24 XThR.Tn[8].t36 143.911
R23308 XThR.Tn[8].n19 XThR.Tn[8].t65 143.911
R23309 XThR.Tn[8].n14 XThR.Tn[8].t53 143.911
R23310 XThR.Tn[8].n9 XThR.Tn[8].t13 143.911
R23311 XThR.Tn[8] XThR.Tn[8].n2 35.7652
R23312 XThR.Tn[8].n85 XThR.Tn[8].t2 26.5955
R23313 XThR.Tn[8].n85 XThR.Tn[8].t0 26.5955
R23314 XThR.Tn[8].n0 XThR.Tn[8].t10 26.5955
R23315 XThR.Tn[8].n0 XThR.Tn[8].t8 26.5955
R23316 XThR.Tn[8].n1 XThR.Tn[8].t11 26.5955
R23317 XThR.Tn[8].n1 XThR.Tn[8].t9 26.5955
R23318 XThR.Tn[8].n86 XThR.Tn[8].t3 26.5955
R23319 XThR.Tn[8].n86 XThR.Tn[8].t1 26.5955
R23320 XThR.Tn[8].n4 XThR.Tn[8].t4 24.9236
R23321 XThR.Tn[8].n4 XThR.Tn[8].t6 24.9236
R23322 XThR.Tn[8].n3 XThR.Tn[8].t5 24.9236
R23323 XThR.Tn[8].n3 XThR.Tn[8].t7 24.9236
R23324 XThR.Tn[8] XThR.Tn[8].n5 18.8943
R23325 XThR.Tn[8].n88 XThR.Tn[8].n87 13.5534
R23326 XThR.Tn[8].n84 XThR.Tn[8] 7.82692
R23327 XThR.Tn[8].n84 XThR.Tn[8] 6.34069
R23328 XThR.Tn[8] XThR.Tn[8].n7 5.34038
R23329 XThR.Tn[8].n12 XThR.Tn[8].n11 4.5005
R23330 XThR.Tn[8].n17 XThR.Tn[8].n16 4.5005
R23331 XThR.Tn[8].n22 XThR.Tn[8].n21 4.5005
R23332 XThR.Tn[8].n27 XThR.Tn[8].n26 4.5005
R23333 XThR.Tn[8].n32 XThR.Tn[8].n31 4.5005
R23334 XThR.Tn[8].n37 XThR.Tn[8].n36 4.5005
R23335 XThR.Tn[8].n42 XThR.Tn[8].n41 4.5005
R23336 XThR.Tn[8].n47 XThR.Tn[8].n46 4.5005
R23337 XThR.Tn[8].n52 XThR.Tn[8].n51 4.5005
R23338 XThR.Tn[8].n57 XThR.Tn[8].n56 4.5005
R23339 XThR.Tn[8].n62 XThR.Tn[8].n61 4.5005
R23340 XThR.Tn[8].n67 XThR.Tn[8].n66 4.5005
R23341 XThR.Tn[8].n72 XThR.Tn[8].n71 4.5005
R23342 XThR.Tn[8].n77 XThR.Tn[8].n76 4.5005
R23343 XThR.Tn[8].n82 XThR.Tn[8].n81 4.5005
R23344 XThR.Tn[8].n83 XThR.Tn[8] 3.70586
R23345 XThR.Tn[8].n12 XThR.Tn[8] 2.52282
R23346 XThR.Tn[8].n17 XThR.Tn[8] 2.52282
R23347 XThR.Tn[8].n22 XThR.Tn[8] 2.52282
R23348 XThR.Tn[8].n27 XThR.Tn[8] 2.52282
R23349 XThR.Tn[8].n32 XThR.Tn[8] 2.52282
R23350 XThR.Tn[8].n37 XThR.Tn[8] 2.52282
R23351 XThR.Tn[8].n42 XThR.Tn[8] 2.52282
R23352 XThR.Tn[8].n47 XThR.Tn[8] 2.52282
R23353 XThR.Tn[8].n52 XThR.Tn[8] 2.52282
R23354 XThR.Tn[8].n57 XThR.Tn[8] 2.52282
R23355 XThR.Tn[8].n62 XThR.Tn[8] 2.52282
R23356 XThR.Tn[8].n67 XThR.Tn[8] 2.52282
R23357 XThR.Tn[8].n72 XThR.Tn[8] 2.52282
R23358 XThR.Tn[8].n77 XThR.Tn[8] 2.52282
R23359 XThR.Tn[8].n82 XThR.Tn[8] 2.52282
R23360 XThR.Tn[8] XThR.Tn[8].n84 1.79489
R23361 XThR.Tn[8] XThR.Tn[8].n88 1.50638
R23362 XThR.Tn[8].n88 XThR.Tn[8] 1.19676
R23363 XThR.Tn[8].n80 XThR.Tn[8] 1.08677
R23364 XThR.Tn[8].n75 XThR.Tn[8] 1.08677
R23365 XThR.Tn[8].n70 XThR.Tn[8] 1.08677
R23366 XThR.Tn[8].n65 XThR.Tn[8] 1.08677
R23367 XThR.Tn[8].n60 XThR.Tn[8] 1.08677
R23368 XThR.Tn[8].n55 XThR.Tn[8] 1.08677
R23369 XThR.Tn[8].n50 XThR.Tn[8] 1.08677
R23370 XThR.Tn[8].n45 XThR.Tn[8] 1.08677
R23371 XThR.Tn[8].n40 XThR.Tn[8] 1.08677
R23372 XThR.Tn[8].n35 XThR.Tn[8] 1.08677
R23373 XThR.Tn[8].n30 XThR.Tn[8] 1.08677
R23374 XThR.Tn[8].n25 XThR.Tn[8] 1.08677
R23375 XThR.Tn[8].n20 XThR.Tn[8] 1.08677
R23376 XThR.Tn[8].n15 XThR.Tn[8] 1.08677
R23377 XThR.Tn[8].n10 XThR.Tn[8] 1.08677
R23378 XThR.Tn[8] XThR.Tn[8].n12 0.839786
R23379 XThR.Tn[8] XThR.Tn[8].n17 0.839786
R23380 XThR.Tn[8] XThR.Tn[8].n22 0.839786
R23381 XThR.Tn[8] XThR.Tn[8].n27 0.839786
R23382 XThR.Tn[8] XThR.Tn[8].n32 0.839786
R23383 XThR.Tn[8] XThR.Tn[8].n37 0.839786
R23384 XThR.Tn[8] XThR.Tn[8].n42 0.839786
R23385 XThR.Tn[8] XThR.Tn[8].n47 0.839786
R23386 XThR.Tn[8] XThR.Tn[8].n52 0.839786
R23387 XThR.Tn[8] XThR.Tn[8].n57 0.839786
R23388 XThR.Tn[8] XThR.Tn[8].n62 0.839786
R23389 XThR.Tn[8] XThR.Tn[8].n67 0.839786
R23390 XThR.Tn[8] XThR.Tn[8].n72 0.839786
R23391 XThR.Tn[8] XThR.Tn[8].n77 0.839786
R23392 XThR.Tn[8] XThR.Tn[8].n82 0.839786
R23393 XThR.Tn[8].n7 XThR.Tn[8] 0.499542
R23394 XThR.Tn[8].n81 XThR.Tn[8] 0.063
R23395 XThR.Tn[8].n76 XThR.Tn[8] 0.063
R23396 XThR.Tn[8].n71 XThR.Tn[8] 0.063
R23397 XThR.Tn[8].n66 XThR.Tn[8] 0.063
R23398 XThR.Tn[8].n61 XThR.Tn[8] 0.063
R23399 XThR.Tn[8].n56 XThR.Tn[8] 0.063
R23400 XThR.Tn[8].n51 XThR.Tn[8] 0.063
R23401 XThR.Tn[8].n46 XThR.Tn[8] 0.063
R23402 XThR.Tn[8].n41 XThR.Tn[8] 0.063
R23403 XThR.Tn[8].n36 XThR.Tn[8] 0.063
R23404 XThR.Tn[8].n31 XThR.Tn[8] 0.063
R23405 XThR.Tn[8].n26 XThR.Tn[8] 0.063
R23406 XThR.Tn[8].n21 XThR.Tn[8] 0.063
R23407 XThR.Tn[8].n16 XThR.Tn[8] 0.063
R23408 XThR.Tn[8].n11 XThR.Tn[8] 0.063
R23409 XThR.Tn[8].n83 XThR.Tn[8] 0.0540714
R23410 XThR.Tn[8] XThR.Tn[8].n83 0.038
R23411 XThR.Tn[8].n7 XThR.Tn[8] 0.0143889
R23412 XThR.Tn[8].n81 XThR.Tn[8].n80 0.00771154
R23413 XThR.Tn[8].n76 XThR.Tn[8].n75 0.00771154
R23414 XThR.Tn[8].n71 XThR.Tn[8].n70 0.00771154
R23415 XThR.Tn[8].n66 XThR.Tn[8].n65 0.00771154
R23416 XThR.Tn[8].n61 XThR.Tn[8].n60 0.00771154
R23417 XThR.Tn[8].n56 XThR.Tn[8].n55 0.00771154
R23418 XThR.Tn[8].n51 XThR.Tn[8].n50 0.00771154
R23419 XThR.Tn[8].n46 XThR.Tn[8].n45 0.00771154
R23420 XThR.Tn[8].n41 XThR.Tn[8].n40 0.00771154
R23421 XThR.Tn[8].n36 XThR.Tn[8].n35 0.00771154
R23422 XThR.Tn[8].n31 XThR.Tn[8].n30 0.00771154
R23423 XThR.Tn[8].n26 XThR.Tn[8].n25 0.00771154
R23424 XThR.Tn[8].n21 XThR.Tn[8].n20 0.00771154
R23425 XThR.Tn[8].n16 XThR.Tn[8].n15 0.00771154
R23426 XThR.Tn[8].n11 XThR.Tn[8].n10 0.00771154
R23427 thermo15c_0.XTB3.Y.n6 thermo15c_0.XTB3.Y.t3 212.081
R23428 thermo15c_0.XTB3.Y.n5 thermo15c_0.XTB3.Y.t15 212.081
R23429 thermo15c_0.XTB3.Y.n11 thermo15c_0.XTB3.Y.t14 212.081
R23430 thermo15c_0.XTB3.Y.n3 thermo15c_0.XTB3.Y.t10 212.081
R23431 thermo15c_0.XTB3.Y.n15 thermo15c_0.XTB3.Y.t11 212.081
R23432 thermo15c_0.XTB3.Y.n16 thermo15c_0.XTB3.Y.t12 212.081
R23433 thermo15c_0.XTB3.Y.n18 thermo15c_0.XTB3.Y.t4 212.081
R23434 thermo15c_0.XTB3.Y.n14 thermo15c_0.XTB3.Y.t16 212.081
R23435 thermo15c_0.XTB3.Y.n22 thermo15c_0.XTB3.Y.n2 201.288
R23436 thermo15c_0.XTB3.Y.n8 thermo15c_0.XTB3.Y.n7 173.761
R23437 thermo15c_0.XTB3.Y.n17 thermo15c_0.XTB3.Y 158.656
R23438 thermo15c_0.XTB3.Y.n10 thermo15c_0.XTB3.Y.n9 152
R23439 thermo15c_0.XTB3.Y.n8 thermo15c_0.XTB3.Y.n4 152
R23440 thermo15c_0.XTB3.Y.n13 thermo15c_0.XTB3.Y.n12 152
R23441 thermo15c_0.XTB3.Y.n20 thermo15c_0.XTB3.Y.n19 152
R23442 thermo15c_0.XTB3.Y.n6 thermo15c_0.XTB3.Y.t9 139.78
R23443 thermo15c_0.XTB3.Y.n5 thermo15c_0.XTB3.Y.t6 139.78
R23444 thermo15c_0.XTB3.Y.n11 thermo15c_0.XTB3.Y.t5 139.78
R23445 thermo15c_0.XTB3.Y.n3 thermo15c_0.XTB3.Y.t17 139.78
R23446 thermo15c_0.XTB3.Y.n15 thermo15c_0.XTB3.Y.t8 139.78
R23447 thermo15c_0.XTB3.Y.n16 thermo15c_0.XTB3.Y.t18 139.78
R23448 thermo15c_0.XTB3.Y.n18 thermo15c_0.XTB3.Y.t13 139.78
R23449 thermo15c_0.XTB3.Y.n14 thermo15c_0.XTB3.Y.t7 139.78
R23450 thermo15c_0.XTB3.Y.n0 thermo15c_0.XTB3.Y.t1 132.067
R23451 thermo15c_0.XTB3.Y.n21 thermo15c_0.XTB3.Y.n13 61.4096
R23452 thermo15c_0.XTB3.Y.n16 thermo15c_0.XTB3.Y.n15 61.346
R23453 thermo15c_0.XTB3.Y.n21 thermo15c_0.XTB3.Y 54.2785
R23454 thermo15c_0.XTB3.Y.n10 thermo15c_0.XTB3.Y.n4 49.6611
R23455 thermo15c_0.XTB3.Y.n12 thermo15c_0.XTB3.Y.n11 45.2793
R23456 thermo15c_0.XTB3.Y.n7 thermo15c_0.XTB3.Y.n5 42.3581
R23457 thermo15c_0.XTB3.Y.n19 thermo15c_0.XTB3.Y.n14 30.6732
R23458 thermo15c_0.XTB3.Y.n19 thermo15c_0.XTB3.Y.n18 30.6732
R23459 thermo15c_0.XTB3.Y.n18 thermo15c_0.XTB3.Y.n17 30.6732
R23460 thermo15c_0.XTB3.Y.n17 thermo15c_0.XTB3.Y.n16 30.6732
R23461 thermo15c_0.XTB3.Y.n2 thermo15c_0.XTB3.Y.t2 26.5955
R23462 thermo15c_0.XTB3.Y.n2 thermo15c_0.XTB3.Y.t0 26.5955
R23463 thermo15c_0.XTB3.Y thermo15c_0.XTB3.Y.n22 23.489
R23464 thermo15c_0.XTB3.Y.n9 thermo15c_0.XTB3.Y.n8 21.7605
R23465 thermo15c_0.XTB3.Y.n7 thermo15c_0.XTB3.Y.n6 18.9884
R23466 thermo15c_0.XTB3.Y.n12 thermo15c_0.XTB3.Y.n3 16.0672
R23467 thermo15c_0.XTB3.Y.n20 thermo15c_0.XTB3.Y 14.8485
R23468 thermo15c_0.XTB3.Y.n13 thermo15c_0.XTB3.Y 11.5205
R23469 thermo15c_0.XTB3.Y.n22 thermo15c_0.XTB3.Y.n21 10.8207
R23470 thermo15c_0.XTB3.Y.n9 thermo15c_0.XTB3.Y 10.2405
R23471 thermo15c_0.XTB3.Y thermo15c_0.XTB3.Y.n20 8.7045
R23472 thermo15c_0.XTB3.Y.n5 thermo15c_0.XTB3.Y.n4 7.30353
R23473 thermo15c_0.XTB3.Y.n11 thermo15c_0.XTB3.Y.n10 4.38232
R23474 thermo15c_0.XTB3.Y.n1 thermo15c_0.XTB3.Y.n0 4.15748
R23475 thermo15c_0.XTB3.Y thermo15c_0.XTB3.Y.n1 3.76521
R23476 thermo15c_0.XTB3.Y.n0 thermo15c_0.XTB3.Y 1.17559
R23477 thermo15c_0.XTB3.Y.n1 thermo15c_0.XTB3.Y 0.921363
R23478 data[4].n3 data[4].t0 231.835
R23479 data[4].n0 data[4].t3 230.155
R23480 data[4].n0 data[4].t1 157.856
R23481 data[4].n3 data[4].t2 157.07
R23482 data[4].n1 data[4].n0 152
R23483 data[4].n4 data[4].n3 152
R23484 data[4].n2 data[4].n1 25.6681
R23485 data[4].n4 data[4].n2 10.7642
R23486 data[4].n2 data[4] 2.763
R23487 data[4].n1 data[4] 2.10199
R23488 data[4] data[4].n4 2.01193
R23489 XThR.Tn[13].n87 XThR.Tn[13].n86 256.103
R23490 XThR.Tn[13].n2 XThR.Tn[13].n0 243.68
R23491 XThR.Tn[13].n5 XThR.Tn[13].n3 241.847
R23492 XThR.Tn[13].n2 XThR.Tn[13].n1 205.28
R23493 XThR.Tn[13].n87 XThR.Tn[13].n85 202.094
R23494 XThR.Tn[13].n5 XThR.Tn[13].n4 185
R23495 XThR.Tn[13] XThR.Tn[13].n78 161.363
R23496 XThR.Tn[13] XThR.Tn[13].n73 161.363
R23497 XThR.Tn[13] XThR.Tn[13].n68 161.363
R23498 XThR.Tn[13] XThR.Tn[13].n63 161.363
R23499 XThR.Tn[13] XThR.Tn[13].n58 161.363
R23500 XThR.Tn[13] XThR.Tn[13].n53 161.363
R23501 XThR.Tn[13] XThR.Tn[13].n48 161.363
R23502 XThR.Tn[13] XThR.Tn[13].n43 161.363
R23503 XThR.Tn[13] XThR.Tn[13].n38 161.363
R23504 XThR.Tn[13] XThR.Tn[13].n33 161.363
R23505 XThR.Tn[13] XThR.Tn[13].n28 161.363
R23506 XThR.Tn[13] XThR.Tn[13].n23 161.363
R23507 XThR.Tn[13] XThR.Tn[13].n18 161.363
R23508 XThR.Tn[13] XThR.Tn[13].n13 161.363
R23509 XThR.Tn[13] XThR.Tn[13].n8 161.363
R23510 XThR.Tn[13] XThR.Tn[13].n6 161.363
R23511 XThR.Tn[13].n80 XThR.Tn[13].n79 161.3
R23512 XThR.Tn[13].n75 XThR.Tn[13].n74 161.3
R23513 XThR.Tn[13].n70 XThR.Tn[13].n69 161.3
R23514 XThR.Tn[13].n65 XThR.Tn[13].n64 161.3
R23515 XThR.Tn[13].n60 XThR.Tn[13].n59 161.3
R23516 XThR.Tn[13].n55 XThR.Tn[13].n54 161.3
R23517 XThR.Tn[13].n50 XThR.Tn[13].n49 161.3
R23518 XThR.Tn[13].n45 XThR.Tn[13].n44 161.3
R23519 XThR.Tn[13].n40 XThR.Tn[13].n39 161.3
R23520 XThR.Tn[13].n35 XThR.Tn[13].n34 161.3
R23521 XThR.Tn[13].n30 XThR.Tn[13].n29 161.3
R23522 XThR.Tn[13].n25 XThR.Tn[13].n24 161.3
R23523 XThR.Tn[13].n20 XThR.Tn[13].n19 161.3
R23524 XThR.Tn[13].n15 XThR.Tn[13].n14 161.3
R23525 XThR.Tn[13].n10 XThR.Tn[13].n9 161.3
R23526 XThR.Tn[13].n78 XThR.Tn[13].t56 161.106
R23527 XThR.Tn[13].n73 XThR.Tn[13].t62 161.106
R23528 XThR.Tn[13].n68 XThR.Tn[13].t40 161.106
R23529 XThR.Tn[13].n63 XThR.Tn[13].t27 161.106
R23530 XThR.Tn[13].n58 XThR.Tn[13].t55 161.106
R23531 XThR.Tn[13].n53 XThR.Tn[13].t17 161.106
R23532 XThR.Tn[13].n48 XThR.Tn[13].t59 161.106
R23533 XThR.Tn[13].n43 XThR.Tn[13].t38 161.106
R23534 XThR.Tn[13].n38 XThR.Tn[13].t25 161.106
R23535 XThR.Tn[13].n33 XThR.Tn[13].t30 161.106
R23536 XThR.Tn[13].n28 XThR.Tn[13].t16 161.106
R23537 XThR.Tn[13].n23 XThR.Tn[13].t39 161.106
R23538 XThR.Tn[13].n18 XThR.Tn[13].t14 161.106
R23539 XThR.Tn[13].n13 XThR.Tn[13].t57 161.106
R23540 XThR.Tn[13].n8 XThR.Tn[13].t21 161.106
R23541 XThR.Tn[13].n6 XThR.Tn[13].t64 161.106
R23542 XThR.Tn[13].n79 XThR.Tn[13].t47 159.978
R23543 XThR.Tn[13].n74 XThR.Tn[13].t54 159.978
R23544 XThR.Tn[13].n69 XThR.Tn[13].t36 159.978
R23545 XThR.Tn[13].n64 XThR.Tn[13].t20 159.978
R23546 XThR.Tn[13].n59 XThR.Tn[13].t45 159.978
R23547 XThR.Tn[13].n54 XThR.Tn[13].t73 159.978
R23548 XThR.Tn[13].n49 XThR.Tn[13].t53 159.978
R23549 XThR.Tn[13].n44 XThR.Tn[13].t33 159.978
R23550 XThR.Tn[13].n39 XThR.Tn[13].t18 159.978
R23551 XThR.Tn[13].n34 XThR.Tn[13].t26 159.978
R23552 XThR.Tn[13].n29 XThR.Tn[13].t71 159.978
R23553 XThR.Tn[13].n24 XThR.Tn[13].t35 159.978
R23554 XThR.Tn[13].n19 XThR.Tn[13].t70 159.978
R23555 XThR.Tn[13].n14 XThR.Tn[13].t52 159.978
R23556 XThR.Tn[13].n9 XThR.Tn[13].t12 159.978
R23557 XThR.Tn[13].n78 XThR.Tn[13].t42 145.038
R23558 XThR.Tn[13].n73 XThR.Tn[13].t69 145.038
R23559 XThR.Tn[13].n68 XThR.Tn[13].t50 145.038
R23560 XThR.Tn[13].n63 XThR.Tn[13].t31 145.038
R23561 XThR.Tn[13].n58 XThR.Tn[13].t63 145.038
R23562 XThR.Tn[13].n53 XThR.Tn[13].t41 145.038
R23563 XThR.Tn[13].n48 XThR.Tn[13].t51 145.038
R23564 XThR.Tn[13].n43 XThR.Tn[13].t32 145.038
R23565 XThR.Tn[13].n38 XThR.Tn[13].t29 145.038
R23566 XThR.Tn[13].n33 XThR.Tn[13].t60 145.038
R23567 XThR.Tn[13].n28 XThR.Tn[13].t24 145.038
R23568 XThR.Tn[13].n23 XThR.Tn[13].t49 145.038
R23569 XThR.Tn[13].n18 XThR.Tn[13].t22 145.038
R23570 XThR.Tn[13].n13 XThR.Tn[13].t65 145.038
R23571 XThR.Tn[13].n8 XThR.Tn[13].t28 145.038
R23572 XThR.Tn[13].n6 XThR.Tn[13].t72 145.038
R23573 XThR.Tn[13].n79 XThR.Tn[13].t61 143.911
R23574 XThR.Tn[13].n74 XThR.Tn[13].t23 143.911
R23575 XThR.Tn[13].n69 XThR.Tn[13].t67 143.911
R23576 XThR.Tn[13].n64 XThR.Tn[13].t46 143.911
R23577 XThR.Tn[13].n59 XThR.Tn[13].t15 143.911
R23578 XThR.Tn[13].n54 XThR.Tn[13].t58 143.911
R23579 XThR.Tn[13].n49 XThR.Tn[13].t68 143.911
R23580 XThR.Tn[13].n44 XThR.Tn[13].t48 143.911
R23581 XThR.Tn[13].n39 XThR.Tn[13].t43 143.911
R23582 XThR.Tn[13].n34 XThR.Tn[13].t13 143.911
R23583 XThR.Tn[13].n29 XThR.Tn[13].t37 143.911
R23584 XThR.Tn[13].n24 XThR.Tn[13].t66 143.911
R23585 XThR.Tn[13].n19 XThR.Tn[13].t34 143.911
R23586 XThR.Tn[13].n14 XThR.Tn[13].t19 143.911
R23587 XThR.Tn[13].n9 XThR.Tn[13].t44 143.911
R23588 XThR.Tn[13] XThR.Tn[13].n2 35.7652
R23589 XThR.Tn[13].n85 XThR.Tn[13].t2 26.5955
R23590 XThR.Tn[13].n85 XThR.Tn[13].t0 26.5955
R23591 XThR.Tn[13].n0 XThR.Tn[13].t9 26.5955
R23592 XThR.Tn[13].n0 XThR.Tn[13].t11 26.5955
R23593 XThR.Tn[13].n1 XThR.Tn[13].t10 26.5955
R23594 XThR.Tn[13].n1 XThR.Tn[13].t8 26.5955
R23595 XThR.Tn[13].n86 XThR.Tn[13].t3 26.5955
R23596 XThR.Tn[13].n86 XThR.Tn[13].t1 26.5955
R23597 XThR.Tn[13].n4 XThR.Tn[13].t6 24.9236
R23598 XThR.Tn[13].n4 XThR.Tn[13].t4 24.9236
R23599 XThR.Tn[13].n3 XThR.Tn[13].t7 24.9236
R23600 XThR.Tn[13].n3 XThR.Tn[13].t5 24.9236
R23601 XThR.Tn[13] XThR.Tn[13].n5 22.9615
R23602 XThR.Tn[13].n88 XThR.Tn[13].n87 13.5534
R23603 XThR.Tn[13].n84 XThR.Tn[13] 8.8494
R23604 XThR.Tn[13] XThR.Tn[13].n7 5.34038
R23605 XThR.Tn[13].n12 XThR.Tn[13].n11 4.5005
R23606 XThR.Tn[13].n17 XThR.Tn[13].n16 4.5005
R23607 XThR.Tn[13].n22 XThR.Tn[13].n21 4.5005
R23608 XThR.Tn[13].n27 XThR.Tn[13].n26 4.5005
R23609 XThR.Tn[13].n32 XThR.Tn[13].n31 4.5005
R23610 XThR.Tn[13].n37 XThR.Tn[13].n36 4.5005
R23611 XThR.Tn[13].n42 XThR.Tn[13].n41 4.5005
R23612 XThR.Tn[13].n47 XThR.Tn[13].n46 4.5005
R23613 XThR.Tn[13].n52 XThR.Tn[13].n51 4.5005
R23614 XThR.Tn[13].n57 XThR.Tn[13].n56 4.5005
R23615 XThR.Tn[13].n62 XThR.Tn[13].n61 4.5005
R23616 XThR.Tn[13].n67 XThR.Tn[13].n66 4.5005
R23617 XThR.Tn[13].n72 XThR.Tn[13].n71 4.5005
R23618 XThR.Tn[13].n77 XThR.Tn[13].n76 4.5005
R23619 XThR.Tn[13].n82 XThR.Tn[13].n81 4.5005
R23620 XThR.Tn[13].n83 XThR.Tn[13] 3.70586
R23621 XThR.Tn[13].n88 XThR.Tn[13].n84 2.99115
R23622 XThR.Tn[13].n88 XThR.Tn[13] 2.87153
R23623 XThR.Tn[13].n12 XThR.Tn[13] 2.52282
R23624 XThR.Tn[13].n17 XThR.Tn[13] 2.52282
R23625 XThR.Tn[13].n22 XThR.Tn[13] 2.52282
R23626 XThR.Tn[13].n27 XThR.Tn[13] 2.52282
R23627 XThR.Tn[13].n32 XThR.Tn[13] 2.52282
R23628 XThR.Tn[13].n37 XThR.Tn[13] 2.52282
R23629 XThR.Tn[13].n42 XThR.Tn[13] 2.52282
R23630 XThR.Tn[13].n47 XThR.Tn[13] 2.52282
R23631 XThR.Tn[13].n52 XThR.Tn[13] 2.52282
R23632 XThR.Tn[13].n57 XThR.Tn[13] 2.52282
R23633 XThR.Tn[13].n62 XThR.Tn[13] 2.52282
R23634 XThR.Tn[13].n67 XThR.Tn[13] 2.52282
R23635 XThR.Tn[13].n72 XThR.Tn[13] 2.52282
R23636 XThR.Tn[13].n77 XThR.Tn[13] 2.52282
R23637 XThR.Tn[13].n82 XThR.Tn[13] 2.52282
R23638 XThR.Tn[13].n84 XThR.Tn[13] 2.2734
R23639 XThR.Tn[13] XThR.Tn[13].n88 1.50638
R23640 XThR.Tn[13].n80 XThR.Tn[13] 1.08677
R23641 XThR.Tn[13].n75 XThR.Tn[13] 1.08677
R23642 XThR.Tn[13].n70 XThR.Tn[13] 1.08677
R23643 XThR.Tn[13].n65 XThR.Tn[13] 1.08677
R23644 XThR.Tn[13].n60 XThR.Tn[13] 1.08677
R23645 XThR.Tn[13].n55 XThR.Tn[13] 1.08677
R23646 XThR.Tn[13].n50 XThR.Tn[13] 1.08677
R23647 XThR.Tn[13].n45 XThR.Tn[13] 1.08677
R23648 XThR.Tn[13].n40 XThR.Tn[13] 1.08677
R23649 XThR.Tn[13].n35 XThR.Tn[13] 1.08677
R23650 XThR.Tn[13].n30 XThR.Tn[13] 1.08677
R23651 XThR.Tn[13].n25 XThR.Tn[13] 1.08677
R23652 XThR.Tn[13].n20 XThR.Tn[13] 1.08677
R23653 XThR.Tn[13].n15 XThR.Tn[13] 1.08677
R23654 XThR.Tn[13].n10 XThR.Tn[13] 1.08677
R23655 XThR.Tn[13] XThR.Tn[13].n12 0.839786
R23656 XThR.Tn[13] XThR.Tn[13].n17 0.839786
R23657 XThR.Tn[13] XThR.Tn[13].n22 0.839786
R23658 XThR.Tn[13] XThR.Tn[13].n27 0.839786
R23659 XThR.Tn[13] XThR.Tn[13].n32 0.839786
R23660 XThR.Tn[13] XThR.Tn[13].n37 0.839786
R23661 XThR.Tn[13] XThR.Tn[13].n42 0.839786
R23662 XThR.Tn[13] XThR.Tn[13].n47 0.839786
R23663 XThR.Tn[13] XThR.Tn[13].n52 0.839786
R23664 XThR.Tn[13] XThR.Tn[13].n57 0.839786
R23665 XThR.Tn[13] XThR.Tn[13].n62 0.839786
R23666 XThR.Tn[13] XThR.Tn[13].n67 0.839786
R23667 XThR.Tn[13] XThR.Tn[13].n72 0.839786
R23668 XThR.Tn[13] XThR.Tn[13].n77 0.839786
R23669 XThR.Tn[13] XThR.Tn[13].n82 0.839786
R23670 XThR.Tn[13].n7 XThR.Tn[13] 0.499542
R23671 XThR.Tn[13].n81 XThR.Tn[13] 0.063
R23672 XThR.Tn[13].n76 XThR.Tn[13] 0.063
R23673 XThR.Tn[13].n71 XThR.Tn[13] 0.063
R23674 XThR.Tn[13].n66 XThR.Tn[13] 0.063
R23675 XThR.Tn[13].n61 XThR.Tn[13] 0.063
R23676 XThR.Tn[13].n56 XThR.Tn[13] 0.063
R23677 XThR.Tn[13].n51 XThR.Tn[13] 0.063
R23678 XThR.Tn[13].n46 XThR.Tn[13] 0.063
R23679 XThR.Tn[13].n41 XThR.Tn[13] 0.063
R23680 XThR.Tn[13].n36 XThR.Tn[13] 0.063
R23681 XThR.Tn[13].n31 XThR.Tn[13] 0.063
R23682 XThR.Tn[13].n26 XThR.Tn[13] 0.063
R23683 XThR.Tn[13].n21 XThR.Tn[13] 0.063
R23684 XThR.Tn[13].n16 XThR.Tn[13] 0.063
R23685 XThR.Tn[13].n11 XThR.Tn[13] 0.063
R23686 XThR.Tn[13].n83 XThR.Tn[13] 0.0540714
R23687 XThR.Tn[13] XThR.Tn[13].n83 0.038
R23688 XThR.Tn[13].n7 XThR.Tn[13] 0.0143889
R23689 XThR.Tn[13].n81 XThR.Tn[13].n80 0.00771154
R23690 XThR.Tn[13].n76 XThR.Tn[13].n75 0.00771154
R23691 XThR.Tn[13].n71 XThR.Tn[13].n70 0.00771154
R23692 XThR.Tn[13].n66 XThR.Tn[13].n65 0.00771154
R23693 XThR.Tn[13].n61 XThR.Tn[13].n60 0.00771154
R23694 XThR.Tn[13].n56 XThR.Tn[13].n55 0.00771154
R23695 XThR.Tn[13].n51 XThR.Tn[13].n50 0.00771154
R23696 XThR.Tn[13].n46 XThR.Tn[13].n45 0.00771154
R23697 XThR.Tn[13].n41 XThR.Tn[13].n40 0.00771154
R23698 XThR.Tn[13].n36 XThR.Tn[13].n35 0.00771154
R23699 XThR.Tn[13].n31 XThR.Tn[13].n30 0.00771154
R23700 XThR.Tn[13].n26 XThR.Tn[13].n25 0.00771154
R23701 XThR.Tn[13].n21 XThR.Tn[13].n20 0.00771154
R23702 XThR.Tn[13].n16 XThR.Tn[13].n15 0.00771154
R23703 XThR.Tn[13].n11 XThR.Tn[13].n10 0.00771154
R23704 data[0].n1 data[0].t0 230.155
R23705 data[0].n0 data[0].t2 228.463
R23706 data[0].n1 data[0].t1 157.856
R23707 data[0].n0 data[0].t3 157.07
R23708 data[0].n2 data[0].n1 152.768
R23709 data[0].n4 data[0].n0 152.256
R23710 data[0].n3 data[0].n2 24.1398
R23711 data[0].n4 data[0].n3 9.48418
R23712 data[0] data[0].n4 6.1445
R23713 data[0].n2 data[0] 5.6325
R23714 data[0].n3 data[0] 2.638
R23715 XThR.XTB4.Y XThR.XTB4.Y.t0 230.518
R23716 XThR.XTB4.Y.n10 XThR.XTB4.Y.t12 212.081
R23717 XThR.XTB4.Y.n11 XThR.XTB4.Y.t2 212.081
R23718 XThR.XTB4.Y.n16 XThR.XTB4.Y.t7 212.081
R23719 XThR.XTB4.Y.n17 XThR.XTB4.Y.t6 212.081
R23720 XThR.XTB4.Y.n0 XThR.XTB4.Y.t17 212.081
R23721 XThR.XTB4.Y.n1 XThR.XTB4.Y.t5 212.081
R23722 XThR.XTB4.Y.n3 XThR.XTB4.Y.t15 212.081
R23723 XThR.XTB4.Y.n4 XThR.XTB4.Y.t4 212.081
R23724 XThR.XTB4.Y.n13 XThR.XTB4.Y.n12 173.761
R23725 XThR.XTB4.Y.n2 XThR.XTB4.Y 167.361
R23726 XThR.XTB4.Y.n19 XThR.XTB4.Y.n18 152
R23727 XThR.XTB4.Y.n15 XThR.XTB4.Y.n14 152
R23728 XThR.XTB4.Y.n13 XThR.XTB4.Y.n9 152
R23729 XThR.XTB4.Y.n6 XThR.XTB4.Y.n5 152
R23730 XThR.XTB4.Y.n10 XThR.XTB4.Y.t3 139.78
R23731 XThR.XTB4.Y.n11 XThR.XTB4.Y.t9 139.78
R23732 XThR.XTB4.Y.n16 XThR.XTB4.Y.t14 139.78
R23733 XThR.XTB4.Y.n17 XThR.XTB4.Y.t11 139.78
R23734 XThR.XTB4.Y.n0 XThR.XTB4.Y.t10 139.78
R23735 XThR.XTB4.Y.n1 XThR.XTB4.Y.t16 139.78
R23736 XThR.XTB4.Y.n3 XThR.XTB4.Y.t8 139.78
R23737 XThR.XTB4.Y.n4 XThR.XTB4.Y.t13 139.78
R23738 XThR.XTB4.Y.n21 XThR.XTB4.Y.t1 133.386
R23739 XThR.XTB4.Y.n20 XThR.XTB4.Y.n19 72.9296
R23740 XThR.XTB4.Y.n1 XThR.XTB4.Y.n0 61.346
R23741 XThR.XTB4.Y.n15 XThR.XTB4.Y.n9 49.6611
R23742 XThR.XTB4.Y.n18 XThR.XTB4.Y.n16 45.2793
R23743 XThR.XTB4.Y.n12 XThR.XTB4.Y.n11 42.3581
R23744 XThR.XTB4.Y.n20 XThR.XTB4.Y.n8 38.1854
R23745 XThR.XTB4.Y.n2 XThR.XTB4.Y.n1 30.6732
R23746 XThR.XTB4.Y.n3 XThR.XTB4.Y.n2 30.6732
R23747 XThR.XTB4.Y.n5 XThR.XTB4.Y.n3 30.6732
R23748 XThR.XTB4.Y.n5 XThR.XTB4.Y.n4 30.6732
R23749 XThR.XTB4.Y XThR.XTB4.Y.n21 28.966
R23750 XThR.XTB4.Y.n14 XThR.XTB4.Y.n13 21.7605
R23751 XThR.XTB4.Y.n14 XThR.XTB4.Y 21.1205
R23752 XThR.XTB4.Y.n12 XThR.XTB4.Y.n10 18.9884
R23753 XThR.XTB4.Y.n18 XThR.XTB4.Y.n17 16.0672
R23754 XThR.XTB4.Y.n21 XThR.XTB4.Y.n20 11.994
R23755 XThR.XTB4.Y.n22 XThR.XTB4.Y 11.6875
R23756 XThR.XTB4.Y.n8 XThR.XTB4.Y.n7 8.21182
R23757 XThR.XTB4.Y.n11 XThR.XTB4.Y.n9 7.30353
R23758 XThR.XTB4.Y.n8 XThR.XTB4.Y.n6 7.24578
R23759 XThR.XTB4.Y.n22 XThR.XTB4.Y 7.23528
R23760 XThR.XTB4.Y.n6 XThR.XTB4.Y 6.08654
R23761 XThR.XTB4.Y XThR.XTB4.Y.n22 5.04292
R23762 XThR.XTB4.Y.n16 XThR.XTB4.Y.n15 4.38232
R23763 XThR.XTB4.Y.n7 XThR.XTB4.Y 1.79489
R23764 XThR.XTB4.Y.n7 XThR.XTB4.Y 0.966538
R23765 XThR.XTB4.Y.n19 XThR.XTB4.Y 0.6405
R23766 XThR.XTB3.Y.n9 XThR.XTB3.Y.t7 212.081
R23767 XThR.XTB3.Y.n10 XThR.XTB3.Y.t11 212.081
R23768 XThR.XTB3.Y.n15 XThR.XTB3.Y.t18 212.081
R23769 XThR.XTB3.Y.n16 XThR.XTB3.Y.t14 212.081
R23770 XThR.XTB3.Y.n1 XThR.XTB3.Y.t9 212.081
R23771 XThR.XTB3.Y.n2 XThR.XTB3.Y.t13 212.081
R23772 XThR.XTB3.Y.n4 XThR.XTB3.Y.t8 212.081
R23773 XThR.XTB3.Y.n5 XThR.XTB3.Y.t12 212.081
R23774 XThR.XTB3.Y.n21 XThR.XTB3.Y.n20 201.288
R23775 XThR.XTB3.Y.n12 XThR.XTB3.Y.n11 173.761
R23776 XThR.XTB3.Y.n3 XThR.XTB3.Y 167.361
R23777 XThR.XTB3.Y.n18 XThR.XTB3.Y.n17 152
R23778 XThR.XTB3.Y.n14 XThR.XTB3.Y.n13 152
R23779 XThR.XTB3.Y.n12 XThR.XTB3.Y.n8 152
R23780 XThR.XTB3.Y.n7 XThR.XTB3.Y.n6 152
R23781 XThR.XTB3.Y.n9 XThR.XTB3.Y.t10 139.78
R23782 XThR.XTB3.Y.n10 XThR.XTB3.Y.t16 139.78
R23783 XThR.XTB3.Y.n15 XThR.XTB3.Y.t5 139.78
R23784 XThR.XTB3.Y.n16 XThR.XTB3.Y.t3 139.78
R23785 XThR.XTB3.Y.n1 XThR.XTB3.Y.t17 139.78
R23786 XThR.XTB3.Y.n2 XThR.XTB3.Y.t6 139.78
R23787 XThR.XTB3.Y.n4 XThR.XTB3.Y.t15 139.78
R23788 XThR.XTB3.Y.n5 XThR.XTB3.Y.t4 139.78
R23789 XThR.XTB3.Y.n0 XThR.XTB3.Y.t1 130.548
R23790 XThR.XTB3.Y.n19 XThR.XTB3.Y.n18 61.4096
R23791 XThR.XTB3.Y.n2 XThR.XTB3.Y.n1 61.346
R23792 XThR.XTB3.Y.n14 XThR.XTB3.Y.n8 49.6611
R23793 XThR.XTB3.Y.n19 XThR.XTB3.Y 45.5863
R23794 XThR.XTB3.Y.n17 XThR.XTB3.Y.n15 45.2793
R23795 XThR.XTB3.Y.n11 XThR.XTB3.Y.n10 42.3581
R23796 XThR.XTB3.Y XThR.XTB3.Y.n21 36.289
R23797 XThR.XTB3.Y.n3 XThR.XTB3.Y.n2 30.6732
R23798 XThR.XTB3.Y.n4 XThR.XTB3.Y.n3 30.6732
R23799 XThR.XTB3.Y.n6 XThR.XTB3.Y.n4 30.6732
R23800 XThR.XTB3.Y.n6 XThR.XTB3.Y.n5 30.6732
R23801 XThR.XTB3.Y.n20 XThR.XTB3.Y.t0 26.5955
R23802 XThR.XTB3.Y.n20 XThR.XTB3.Y.t2 26.5955
R23803 XThR.XTB3.Y.n13 XThR.XTB3.Y.n12 21.7605
R23804 XThR.XTB3.Y.n13 XThR.XTB3.Y 21.1205
R23805 XThR.XTB3.Y.n11 XThR.XTB3.Y.n9 18.9884
R23806 XThR.XTB3.Y XThR.XTB3.Y.n7 17.4085
R23807 XThR.XTB3.Y.n22 XThR.XTB3.Y 16.5652
R23808 XThR.XTB3.Y.n17 XThR.XTB3.Y.n16 16.0672
R23809 XThR.XTB3.Y.n21 XThR.XTB3.Y.n19 10.8207
R23810 XThR.XTB3.Y XThR.XTB3.Y.n22 9.03579
R23811 XThR.XTB3.Y.n10 XThR.XTB3.Y.n8 7.30353
R23812 XThR.XTB3.Y.n7 XThR.XTB3.Y 6.1445
R23813 XThR.XTB3.Y.n15 XThR.XTB3.Y.n14 4.38232
R23814 XThR.XTB3.Y XThR.XTB3.Y.n0 3.46739
R23815 XThR.XTB3.Y.n0 XThR.XTB3.Y 2.74112
R23816 XThR.XTB3.Y.n22 XThR.XTB3.Y 2.21057
R23817 XThR.XTB3.Y.n18 XThR.XTB3.Y 0.6405
R23818 data[6].n0 data[6].t0 230.576
R23819 data[6].n0 data[6].t1 158.275
R23820 data[6].n1 data[6].n0 152
R23821 data[6].n1 data[6] 11.9995
R23822 data[6] data[6].n1 6.66717
R23823 data[1].n4 data[1].t2 230.576
R23824 data[1].n1 data[1].t0 230.363
R23825 data[1].n0 data[1].t4 229.369
R23826 data[1].n4 data[1].t5 158.275
R23827 data[1].n1 data[1].t3 158.064
R23828 data[1].n0 data[1].t1 157.07
R23829 data[1].n2 data[1].n1 153.28
R23830 data[1].n7 data[1].n0 153.147
R23831 data[1].n5 data[1].n4 152
R23832 data[1].n7 data[1].n6 16.3874
R23833 data[1].n6 data[1].n5 14.9641
R23834 data[1].n3 data[1].n2 9.3005
R23835 data[1].n6 data[1].n3 6.49639
R23836 data[1] data[1].n7 3.24826
R23837 data[1].n2 data[1] 2.92621
R23838 data[1].n3 data[1] 2.15819
R23839 data[1].n5 data[1] 2.13383
R23840 data[2].n0 data[2].t0 230.576
R23841 data[2].n0 data[2].t1 158.275
R23842 data[2].n1 data[2].n0 152
R23843 data[2].n1 data[2] 12.7714
R23844 data[2] data[2].n1 2.13383
R23845 data[5].n4 data[5].t2 230.576
R23846 data[5].n1 data[5].t0 230.363
R23847 data[5].n0 data[5].t1 229.369
R23848 data[5].n4 data[5].t5 158.275
R23849 data[5].n1 data[5].t3 158.064
R23850 data[5].n0 data[5].t4 157.07
R23851 data[5].n2 data[5].n1 152.256
R23852 data[5].n7 data[5].n0 152.238
R23853 data[5].n5 data[5].n4 152
R23854 data[5].n7 data[5].n6 16.3874
R23855 data[5].n6 data[5].n5 14.6005
R23856 data[5].n3 data[5].n2 9.3005
R23857 data[5].n5 data[5] 6.66717
R23858 data[5].n6 data[5].n3 6.49639
R23859 data[5].n2 data[5] 6.1445
R23860 data[5] data[5].n7 5.68939
R23861 data[5].n3 data[5] 2.28319
R23862 bias[0] bias[0].t0 12.1467
R23863 bias[2].n0 bias[2].t0 56.8043
R23864 bias[2].n0 bias[2] 6.35112
R23865 bias[2] bias[2].n0 0.828709
R23866 data[3].n0 data[3].t1 230.576
R23867 data[3].n0 data[3].t0 158.275
R23868 data[3].n1 data[3].n0 153.553
R23869 data[3].n1 data[3] 11.6078
R23870 data[3] data[3].n1 2.90959
R23871 data[7].n0 data[7].t0 230.576
R23872 data[7].n0 data[7].t1 158.275
R23873 data[7].n1 data[7].n0 152
R23874 data[7].n1 data[7] 11.9995
R23875 data[7] data[7].n1 6.66717
R23876 bias[1] bias[1].t0 23.8076
C0 XA.XIR[10].XIC[9].icell.PDM VPWR 0.01171f
C1 XA.XIR[7].XIC[13].icell.Ien Vbias 0.19161f
C2 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.Ien 0.04854f
C3 XThR.XTBN.Y XThR.Tn[3] 0.62501f
C4 XA.XIR[11].XIC_dummy_left.icell.Ien XThR.Tn[11] 0.01244f
C5 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.PDM 0.02104f
C6 a_n1049_8581# XThR.Tn[0] 0.2685f
C7 XThR.XTB7.B XThR.Tn[11] 0.03888f
C8 XA.XIR[13].XIC[0].icell.Ien Vbias 0.19149f
C9 XA.XIR[15].XIC[7].icell.Ien VPWR 0.31713f
C10 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.Ien 0.04854f
C11 XThR.Tn[2] XA.XIR[2].XIC[11].icell.Ien 0.14211f
C12 XA.Cn[14] XThR.Tn[7] 0.40742f
C13 XA.Cn[8] XA.XIR[13].XIC[8].icell.PDM 0.02601f
C14 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR 0.38902f
C15 XThR.XTBN.Y XThR.XTB7.Y 0.50018f
C16 XA.XIR[4].XIC[10].icell.Ien VPWR 0.18829f
C17 a_9827_9569# XA.Cn[12] 0.20217f
C18 XA.XIR[0].XIC[1].icell.Ien VPWR 0.18776f
C19 XA.XIR[2].XIC[1].icell.PDM VPWR 0.01171f
C20 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.PDM 0.02104f
C21 XA.XIR[8].XIC[4].icell.Ien VPWR 0.18829f
C22 XA.XIR[7].XIC[13].icell.PDM Vbias 0.03928f
C23 XThR.XTB4.Y XThR.Tn[3] 0.1895f
C24 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.Ien 0.04854f
C25 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PDM 0.04035f
C26 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.PDM 0.02104f
C27 XA.XIR[9].XIC[13].icell.Ien VPWR 0.18829f
C28 XThR.XTB4.Y XThR.XTB7.Y 0.03475f
C29 thermo15c_0.XTBN.Y a_9827_9569# 0.22873f
C30 XThR.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.14211f
C31 thermo15c_0.XTB2.Y a_4067_9615# 0.02133f
C32 XA.XIR[9].XIC[9].icell.PDM Vbias 0.03928f
C33 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.Ien 0.04854f
C34 XA.XIR[0].XIC[6].icell.Ien VPWR 0.1878f
C35 XA.Cn[0] XA.XIR[3].XIC[0].icell.PDM 0.02601f
C36 XThR.Tn[7] Iout 1.1276f
C37 XA.XIR[0].XIC[1].icell.PDM Vbias 0.03945f
C38 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR 0.01604f
C39 XThR.XTB7.Y XThR.Tn[10] 0.07406f
C40 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR 0.01691f
C41 XA.Cn[11] XA.XIR[10].XIC[11].icell.Ien 0.04604f
C42 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.Ien 0.04854f
C43 XA.Cn[12] XThR.Tn[3] 0.40738f
C44 XThR.Tn[5] XA.XIR[5].XIC[0].icell.Ien 0.1423f
C45 XA.XIR[7].XIC[9].icell.Ien VPWR 0.18829f
C46 XA.XIR[4].XIC[2].icell.Ien Iout 0.06801f
C47 XThR.Tn[14] XA.XIR[14].XIC[13].icell.Ien 0.14211f
C48 XA.Cn[4] XA.XIR[11].XIC[4].icell.PDM 0.02601f
C49 VPWR bias[2] 1.20331f
C50 a_4067_9615# VPWR 0.70663f
C51 XA.XIR[3].XIC[10].icell.Ien Vbias 0.19161f
C52 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PDM 0.04035f
C53 XA.Cn[4] XA.Cn[5] 0.31867f
C54 XA.XIR[1].XIC[14].icell.PDM Vbias 0.03928f
C55 XThR.XTBN.Y a_n997_2667# 0.22784f
C56 XA.XIR[10].XIC[14].icell.PDM Vbias 0.03928f
C57 XA.Cn[14] XA.XIR[5].XIC[14].icell.Ien 0.04604f
C58 XA.XIR[9].XIC_dummy_left.icell.Iout XA.XIR[10].XIC_dummy_left.icell.Iout 0.03665f
C59 XA.Cn[13] XThR.Tn[5] 0.40739f
C60 XA.XIR[2].XIC[3].icell.Ien Vbias 0.19161f
C61 XA.XIR[4].XIC[14].icell.PDM Vbias 0.03928f
C62 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.PDM 0.02104f
C63 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR 0.08221f
C64 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.PDM 0.02104f
C65 XA.Cn[14] XA.XIR[3].XIC[14].icell.PDM 0.02601f
C66 XThR.Tn[8] a_n997_3979# 0.1927f
C67 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.Ien 0.04854f
C68 XA.XIR[13].XIC_15.icell.PDM Vbias 0.03927f
C69 XA.XIR[1].XIC[5].icell.Ien Vbias 0.19173f
C70 XA.XIR[2].XIC[0].icell.Ien VPWR 0.18829f
C71 XA.Cn[7] XA.XIR[7].XIC[7].icell.Ien 0.04604f
C72 XA.Cn[6] XA.XIR[12].XIC[6].icell.Ien 0.04604f
C73 XA.XIR[9].XIC[5].icell.Ien Iout 0.06801f
C74 XA.Cn[9] XThR.Tn[0] 0.40759f
C75 XThR.Tn[11] XA.XIR[11].XIC[5].icell.Ien 0.14211f
C76 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PDM 0.04035f
C77 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Ien 0.01557f
C78 XA.Cn[6] VPWR 3.63495f
C79 XA.XIR[8].XIC[13].icell.Ien Vbias 0.19161f
C80 XA.XIR[7].XIC[1].icell.PDM VPWR 0.01171f
C81 XA.XIR[10].XIC[1].icell.Ien VPWR 0.18829f
C82 XThR.XTB4.Y a_n997_2667# 0.07199f
C83 XA.XIR[6].XIC[8].icell.PDM VPWR 0.01171f
C84 XThR.Tn[0] XA.XIR[0].XIC[10].icell.Ien 0.14211f
C85 XThR.Tn[10] XA.XIR[10].XIC[9].icell.Ien 0.14211f
C86 thermo15c_0.XTB7.Y XA.Cn[10] 0.07427f
C87 XThR.Tn[6] XA.XIR[6].XIC[4].icell.Ien 0.14211f
C88 XA.XIR[5].XIC_15.icell.PDM VPWR 0.07527f
C89 XA.XIR[14].XIC[5].icell.PDM VPWR 0.01171f
C90 XA.XIR[5].XIC[14].icell.Ien Iout 0.06801f
C91 thermo15c_0.XTB6.Y a_5949_9615# 0.26831f
C92 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.Ien 0.04854f
C93 XThR.XTBN.Y XThR.Tn[11] 0.52268f
C94 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.Ien 0.04854f
C95 XA.Cn[4] XA.XIR[11].XIC[4].icell.Ien 0.04604f
C96 XA.XIR[13].XIC[9].icell.PDM VPWR 0.01171f
C97 XThR.Tn[7] XA.XIR[7].XIC[11].icell.Ien 0.14211f
C98 XA.XIR[0].XIC_15.icell.Ien Vbias 0.19241f
C99 XThR.XTB7.A XThR.XTB3.Y 0.57441f
C100 XA.Cn[11] XA.XIR[1].XIC[11].icell.PDM 0.02602f
C101 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR 0.01604f
C102 thermo15c_0.XTB7.A thermo15c_0.XTB6.Y 0.19112f
C103 thermo15c_0.XTB6.A thermo15c_0.XTB7.Y 0.01596f
C104 thermo15c_0.XTB3.Y thermo15c_0.XTBN.A 0.03907f
C105 XA.XIR[6].XIC[0].icell.Ien Vbias 0.19149f
C106 XA.XIR[12].XIC[9].icell.Ien Iout 0.06801f
C107 XA.Cn[11] XA.XIR[4].XIC[11].icell.PDM 0.02601f
C108 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout 0.06446f
C109 XThR.Tn[7] XThR.Tn[8] 0.12208f
C110 XA.XIR[11].XIC[13].icell.Ien VPWR 0.18829f
C111 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.PDM 0.02104f
C112 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.Ien 0.04854f
C113 thermo15c_0.XTB7.B XA.Cn[11] 0.03651f
C114 XThR.XTB4.Y XThR.Tn[11] 0.3042f
C115 XA.XIR[3].XIC[6].icell.Ien VPWR 0.18829f
C116 XThR.Tn[14] XA.XIR[14].XIC[11].icell.Ien 0.14211f
C117 XA.XIR[1].XIC[2].icell.PDM VPWR 0.01171f
C118 XA.XIR[11].XIC[4].icell.PDM Vbias 0.03928f
C119 XA.XIR[9].XIC[0].icell.Ien Iout 0.06795f
C120 XA.Cn[5] Vbias 0.82298f
C121 XA.Cn[2] XA.XIR[0].XIC[2].icell.Ien 0.04658f
C122 XA.XIR[4].XIC[2].icell.PDM VPWR 0.01171f
C123 XA.XIR[10].XIC[8].icell.PDM Vbias 0.03928f
C124 XA.Cn[1] XA.XIR[8].XIC[1].icell.PDM 0.02601f
C125 XThR.Tn[10] XThR.Tn[11] 0.10691f
C126 XA.Cn[13] XA.XIR[15].XIC[13].icell.Ien 0.04292f
C127 XA.XIR[3].XIC[10].icell.PDM VPWR 0.01171f
C128 XA.XIR[8].XIC[12].icell.PDM VPWR 0.01171f
C129 XA.XIR[4].XIC_15.icell.Ien VPWR 0.26829f
C130 XA.XIR[6].XIC[5].icell.Ien Vbias 0.19161f
C131 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout 0.06446f
C132 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR 0.08209f
C133 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PDM 0.04035f
C134 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PDM 0.04035f
C135 XA.XIR[8].XIC[9].icell.Ien VPWR 0.18829f
C136 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.Ien 0.04854f
C137 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.Ien 0.04854f
C138 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.PDM 0.02104f
C139 XThR.XTB7.Y XThR.Tn[13] 0.10781f
C140 XA.Cn[12] XThR.Tn[11] 0.40738f
C141 XA.Cn[8] XThR.Tn[6] 0.40738f
C142 XA.XIR[2].XIC[0].icell.PDM Vbias 0.03915f
C143 XA.Cn[11] XA.XIR[13].XIC[11].icell.Ien 0.04604f
C144 XA.XIR[10].XIC[13].icell.PDM Vbias 0.03928f
C145 XA.Cn[4] XA.XIR[14].XIC[4].icell.PDM 0.02601f
C146 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.Ien 0.04854f
C147 XThR.Tn[9] XA.XIR[9].XIC[14].icell.Ien 0.144f
C148 XA.Cn[7] XA.XIR[8].XIC[7].icell.Ien 0.04604f
C149 XA.XIR[0].XIC[11].icell.Ien VPWR 0.18882f
C150 XThR.Tn[12] XA.XIR[12].XIC_dummy_left.icell.Iout 0.03385f
C151 XA.XIR[4].XIC_dummy_right.icell.Iout VPWR 0.11567f
C152 XA.XIR[11].XIC[4].icell.Ien Vbias 0.19161f
C153 XA.XIR[13].XIC[14].icell.PDM Vbias 0.03928f
C154 XA.XIR[15].XIC[4].icell.Ien Iout 0.07192f
C155 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PDM 0.04056f
C156 XA.Cn[14] XA.XIR[12].XIC[14].icell.Ien 0.04604f
C157 XA.XIR[10].XIC[6].icell.Ien Vbias 0.19161f
C158 thermo15c_0.XTBN.A a_9827_9569# 0.09118f
C159 XA.XIR[6].XIC_dummy_left.icell.Iout XA.XIR[7].XIC_dummy_left.icell.Iout 0.03665f
C160 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PDM 0.0404f
C161 XA.XIR[4].XIC[7].icell.Ien Iout 0.06801f
C162 XA.XIR[7].XIC[14].icell.Ien VPWR 0.18835f
C163 XThR.XTB5.Y XThR.XTBN.A 0.10854f
C164 XThR.Tn[13] XA.XIR[13].XIC[4].icell.Ien 0.14211f
C165 XThR.XTB7.A VPWR 0.88595f
C166 XThR.Tn[10] XA.XIR[10].XIC[14].icell.Ien 0.144f
C167 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Iout 0.03842f
C168 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR 0.01691f
C169 XA.XIR[3].XIC_15.icell.Ien Vbias 0.19195f
C170 XA.XIR[11].XIC[11].icell.Ien VPWR 0.18829f
C171 XA.Cn[9] XThR.Tn[1] 0.40744f
C172 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.PDM 0.02104f
C173 XA.XIR[2].XIC[8].icell.Ien Vbias 0.19161f
C174 XA.XIR[13].XIC[1].icell.Ien VPWR 0.18829f
C175 XA.Cn[11] XA.XIR[12].XIC[11].icell.PDM 0.02601f
C176 XA.Cn[2] XA.XIR[12].XIC[2].icell.PDM 0.02601f
C177 XA.XIR[7].XIC[1].icell.Ien Iout 0.06801f
C178 a_3773_9615# Vbias 0.01444f
C179 XA.Cn[1] XThR.Tn[7] 0.40738f
C180 XA.XIR[1].XIC[10].icell.Ien Vbias 0.19173f
C181 XA.Cn[9] XThR.Tn[12] 0.40738f
C182 XA.XIR[9].XIC[10].icell.Ien Iout 0.06801f
C183 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.Ien 0.04854f
C184 XThR.XTB7.B XThR.XTB3.Y 0.23315f
C185 XThR.XTBN.Y XThR.Tn[14] 0.47807f
C186 XA.XIR[12].XIC[14].icell.Ien Iout 0.06801f
C187 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.Ien 0.04854f
C188 XA.Cn[4] XA.XIR[14].XIC[4].icell.Ien 0.04604f
C189 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR 0.08209f
C190 XA.XIR[0].XIC[3].icell.Ien Iout 0.0675f
C191 XA.Cn[2] XA.XIR[3].XIC[2].icell.Ien 0.04604f
C192 XThR.Tn[0] XA.XIR[0].XIC_15.icell.Ien 0.13564f
C193 XA.Cn[8] XThR.Tn[4] 0.40738f
C194 thermo15c_0.XTB5.A data[1] 0.11102f
C195 XThR.Tn[6] XA.XIR[6].XIC[9].icell.Ien 0.14211f
C196 XA.XIR[7].XIC[6].icell.Ien Iout 0.06801f
C197 XA.XIR[7].XIC[0].icell.PDM Vbias 0.03915f
C198 XA.Cn[1] XA.XIR[9].XIC[1].icell.PDM 0.02601f
C199 XA.XIR[14].XIC[13].icell.Ien VPWR 0.18883f
C200 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.PDM 0.02104f
C201 XA.XIR[9].XIC[12].icell.PDM VPWR 0.01171f
C202 XA.XIR[6].XIC[7].icell.PDM Vbias 0.03928f
C203 XA.XIR[0].XIC[4].icell.PDM VPWR 0.01136f
C204 XThR.XTB1.Y XThR.XTBN.A 0.12307f
C205 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout 0.06446f
C206 XA.XIR[14].XIC[4].icell.PDM Vbias 0.03928f
C207 XA.XIR[5].XIC[14].icell.PDM Vbias 0.03928f
C208 XA.XIR[1].XIC[1].icell.Ien VPWR 0.18829f
C209 thermo15c_0.XTB1.Y XA.Cn[0] 0.1842f
C210 thermo15c_0.XTB6.Y XA.Cn[13] 0.32317f
C211 XThR.XTB3.Y XThR.Tn[2] 0.18254f
C212 XA.XIR[10].XIC[2].icell.Ien VPWR 0.18829f
C213 XA.XIR[13].XIC[8].icell.PDM Vbias 0.03928f
C214 XA.Cn[5] XThR.Tn[0] 0.40765f
C215 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.Ien 0.04854f
C216 XA.Cn[8] XA.XIR[5].XIC[8].icell.Ien 0.04604f
C217 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PDM 0.04035f
C218 XThR.XTB5.Y XThR.Tn[4] 0.19957f
C219 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PDM 0.04035f
C220 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PDM 0.04035f
C221 XA.Cn[6] XA.XIR[10].XIC[6].icell.PDM 0.02601f
C222 thermo15c_0.XTB2.Y a_3523_10575# 0.01006f
C223 XA.XIR[3].XIC[11].icell.Ien VPWR 0.18829f
C224 XA.Cn[9] XA.Cn[10] 0.0671f
C225 XThR.Tn[10] XA.XIR[10].XIC[12].icell.Ien 0.14211f
C226 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR 0.01691f
C227 thermo15c_0.XTB7.Y XA.Cn[6] 0.2182f
C228 XA.Cn[14] Iout 0.22441f
C229 XA.XIR[2].XIC[4].icell.Ien VPWR 0.18829f
C230 XA.Cn[0] XThR.Tn[5] 0.40739f
C231 XThR.Tn[1] a_n1049_7787# 0.26879f
C232 XA.Cn[6] XA.XIR[15].XIC[6].icell.Ien 0.04292f
C233 XA.Cn[10] XA.XIR[0].XIC[10].icell.Ien 0.04662f
C234 XA.XIR[1].XIC[6].icell.Ien VPWR 0.18829f
C235 XA.XIR[10].XIC[12].icell.PDM Vbias 0.03928f
C236 XA.Cn[12] XThR.Tn[14] 0.40738f
C237 XA.XIR[1].XIC[1].icell.PDM Vbias 0.03928f
C238 XThR.XTB5.Y XThR.XTB6.Y 2.12831f
C239 XA.XIR[6].XIC[10].icell.Ien Vbias 0.19161f
C240 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.PDM 0.02104f
C241 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.Ien 0.04854f
C242 XA.XIR[13].XIC[13].icell.PDM Vbias 0.03928f
C243 XA.XIR[4].XIC[1].icell.PDM Vbias 0.03928f
C244 XA.XIR[8].XIC[14].icell.Ien VPWR 0.18835f
C245 XA.Cn[12] XA.XIR[10].XIC[12].icell.Ien 0.04604f
C246 XA.XIR[12].XIC[12].icell.Ien Iout 0.06801f
C247 XA.XIR[3].XIC[9].icell.PDM Vbias 0.03928f
C248 XA.XIR[8].XIC[11].icell.PDM Vbias 0.03928f
C249 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR 0.38914f
C250 XA.XIR[14].XIC[4].icell.Ien Vbias 0.19161f
C251 XThR.Tn[7] XA.XIR[7].XIC_dummy_left.icell.Iout 0.0402f
C252 XThR.XTB7.B VPWR 1.67447f
C253 XA.Cn[11] XA.XIR[5].XIC[11].icell.PDM 0.02601f
C254 thermo15c_0.XTB7.B XA.Cn[7] 0.07854f
C255 XA.XIR[2].XIC_15.icell.PDM Vbias 0.03927f
C256 XA.XIR[13].XIC[6].icell.Ien Vbias 0.19161f
C257 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.PDM 0.02104f
C258 thermo15c_0.XTB7.A XA.Cn[2] 0.1255f
C259 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.PDM 0.02104f
C260 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PDM 0.0404f
C261 XA.XIR[8].XIC[1].icell.Ien Iout 0.06801f
C262 XA.Cn[3] XThR.Tn[2] 0.40741f
C263 XA.XIR[3].XIC[3].icell.Ien Iout 0.06801f
C264 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PDM 0.04035f
C265 XA.XIR[14].XIC[11].icell.Ien VPWR 0.18883f
C266 XA.XIR[11].XIC[9].icell.Ien Vbias 0.19161f
C267 XThR.Tn[1] XA.XIR[1].XIC[5].icell.Ien 0.14211f
C268 XThR.Tn[14] XA.XIR[14].XIC[5].icell.Ien 0.14211f
C269 XA.XIR[15].XIC[9].icell.Ien Iout 0.07192f
C270 XA.XIR[5].XIC[2].icell.PDM VPWR 0.01171f
C271 XA.Cn[11] XA.XIR[15].XIC[11].icell.PDM 0.02601f
C272 XA.XIR[6].XIC[1].icell.Ien VPWR 0.18829f
C273 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PDM 0.04035f
C274 XThR.XTBN.Y XThR.XTB3.Y 0.17246f
C275 XA.Cn[2] XA.XIR[15].XIC[2].icell.PDM 0.02601f
C276 XA.XIR[4].XIC[12].icell.Ien Iout 0.06801f
C277 XA.Cn[12] XA.XIR[0].XIC[12].icell.PDM 0.0279f
C278 XThR.Tn[13] XA.XIR[13].XIC[9].icell.Ien 0.14211f
C279 XA.XIR[12].XIC[1].icell.PDM VPWR 0.01171f
C280 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.PDM 0.02104f
C281 XThR.Tn[2] VPWR 8.04926f
C282 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.PDM 0.02104f
C283 XA.XIR[8].XIC[6].icell.Ien Iout 0.06801f
C284 XA.XIR[11].XIC[7].icell.PDM VPWR 0.01171f
C285 XThR.XTB1.Y XThR.XTB6.Y 0.05751f
C286 XA.Cn[4] XThR.Tn[6] 0.40738f
C287 XA.XIR[2].XIC[13].icell.Ien Vbias 0.19161f
C288 thermo15c_0.XTB4.Y XA.Cn[11] 0.30457f
C289 XThR.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.14211f
C290 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.PDM 0.02104f
C291 XA.Cn[0] XA.XIR[6].XIC[0].icell.PDM 0.02601f
C292 XA.Cn[9] XA.XIR[10].XIC[9].icell.PDM 0.02601f
C293 XA.XIR[1].XIC_15.icell.Ien Vbias 0.19206f
C294 XA.Cn[3] XA.XIR[2].XIC[3].icell.PDM 0.02602f
C295 XA.XIR[9].XIC_15.icell.Ien Iout 0.0694f
C296 XThR.XTB3.Y XThR.XTB4.Y 2.13136f
C297 XA.XIR[6].XIC[6].icell.Ien VPWR 0.18829f
C298 XA.Cn[13] XThR.Tn[9] 0.40739f
C299 XA.Cn[14] XThR.Tn[8] 0.40742f
C300 XA.XIR[0].XIC[8].icell.Ien Iout 0.0675f
C301 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.PDM 0.02104f
C302 XThR.XTB3.Y XThR.Tn[10] 0.29462f
C303 XA.Cn[10] XA.XIR[3].XIC[10].icell.Ien 0.04604f
C304 XA.XIR[0].XIC_dummy_left.icell.Iout VPWR 0.1175f
C305 XA.XIR[12].XIC[10].icell.Ien Iout 0.06801f
C306 XA.XIR[2].XIC[3].icell.PDM VPWR 0.01171f
C307 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14] 0.14211f
C308 XThR.Tn[6] XA.XIR[6].XIC[14].icell.Ien 0.144f
C309 XA.XIR[13].XIC[2].icell.Ien VPWR 0.18829f
C310 XA.XIR[7].XIC[11].icell.Ien Iout 0.06801f
C311 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.Ien 0.04854f
C312 XA.XIR[7].XIC_15.icell.PDM Vbias 0.03927f
C313 XA.XIR[5].XIC[3].icell.Ien Vbias 0.19161f
C314 XA.Cn[14] XA.XIR[6].XIC[14].icell.PDM 0.02601f
C315 XThR.Tn[13] XThR.Tn[14] 0.20347f
C316 XA.Cn[2] XA.XIR[1].XIC[2].icell.Ien 0.04606f
C317 XA.Cn[5] XThR.Tn[1] 0.40744f
C318 XA.Cn[1] XA.XIR[7].XIC[1].icell.Ien 0.04604f
C319 XA.Cn[6] XA.XIR[13].XIC[6].icell.PDM 0.02601f
C320 XA.Cn[14] XA.XIR[15].XIC[14].icell.Ien 0.04292f
C321 XA.XIR[11].XIC[5].icell.Ien VPWR 0.18829f
C322 XA.XIR[9].XIC_dummy_right.icell.Iout Iout 0.01732f
C323 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PDM 0.04035f
C324 XA.XIR[10].XIC[11].icell.PDM Vbias 0.03928f
C325 XThR.Tn[8] Iout 1.12761f
C326 XA.XIR[3].XIC[0].icell.Ien Iout 0.06795f
C327 XA.Cn[5] XThR.Tn[12] 0.40738f
C328 XThR.Tn[8] XA.XIR[8].XIC[1].icell.Ien 0.14211f
C329 XA.XIR[10].XIC[7].icell.Ien VPWR 0.18829f
C330 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.PDM 0.02104f
C331 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.PDM 0.02104f
C332 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR 0.35722f
C333 thermo15c_0.XTB4.Y a_4861_9615# 0.23756f
C334 thermo15c_0.XTBN.Y a_10915_9569# 0.21503f
C335 XThR.XTB7.Y XThR.Tn[7] 0.0835f
C336 XA.XIR[9].XIC[11].icell.PDM Vbias 0.03928f
C337 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Iout 0.01728f
C338 XA.XIR[13].XIC[12].icell.PDM Vbias 0.03928f
C339 XA.XIR[0].XIC[3].icell.PDM Vbias 0.03945f
C340 thermo15c_0.XTB5.Y a_5155_10571# 0.01188f
C341 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.PDM 0.02104f
C342 XA.XIR[11].XIC[1].icell.Ien Iout 0.06801f
C343 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR 0.01604f
C344 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PDM 0.04035f
C345 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.PDM 0.02104f
C346 XThR.XTBN.Y VPWR 4.54335f
C347 XA.Cn[4] XThR.Tn[4] 0.40738f
C348 XA.Cn[5] XA.XIR[4].XIC[5].icell.Ien 0.04604f
C349 XA.Cn[12] XA.XIR[13].XIC[12].icell.Ien 0.04604f
C350 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PDM 0.0404f
C351 XA.XIR[2].XIC[9].icell.Ien VPWR 0.18829f
C352 XA.Cn[9] XA.XIR[7].XIC[9].icell.Ien 0.04604f
C353 XThR.XTB2.Y data[5] 0.017f
C354 thermo15c_0.XTB5.A thermo15c_0.XTB2.Y 0.02203f
C355 XA.Cn[8] XA.XIR[12].XIC[8].icell.Ien 0.04604f
C356 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.PDM 0.02104f
C357 XA.XIR[1].XIC[11].icell.Ien VPWR 0.18829f
C358 XThR.Tn[6] Vbias 1.39526f
C359 a_5155_9615# VPWR 0.7051f
C360 XA.XIR[11].XIC[14].icell.Ien Vbias 0.19161f
C361 XThR.Tn[8] XA.XIR[8].XIC[6].icell.Ien 0.14211f
C362 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PDM 0.04035f
C363 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.Ien 0.04854f
C364 XA.XIR[15].XIC[14].icell.Ien Iout 0.07192f
C365 XA.Cn[3] XThR.Tn[10] 0.40738f
C366 XA.XIR[6].XIC_15.icell.Ien Vbias 0.19195f
C367 XA.Cn[3] XA.XIR[7].XIC[3].icell.PDM 0.02601f
C368 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.Ien 0.04854f
C369 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.PDM 0.02104f
C370 XThR.Tn[13] XA.XIR[13].XIC[14].icell.Ien 0.144f
C371 XThR.XTB4.Y VPWR 0.92827f
C372 XA.Cn[7] XA.XIR[2].XIC[7].icell.Ien 0.04605f
C373 thermo15c_0.XTB5.A VPWR 0.82807f
C374 XA.XIR[14].XIC[9].icell.Ien Vbias 0.19161f
C375 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.PDM 0.02104f
C376 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PDM 0.04056f
C377 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.Ien 0.04854f
C378 thermo15c_0.XTBN.A data[1] 0.01444f
C379 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PDM 0.04035f
C380 XThR.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.14211f
C381 XA.Cn[7] XA.Cn[8] 0.06603f
C382 XThR.Tn[10] XA.XIR[10].XIC_15.icell.Ien 0.13564f
C383 XA.XIR[7].XIC[3].icell.PDM VPWR 0.01171f
C384 XThR.Tn[10] VPWR 8.95184f
C385 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Ien 0.01557f
C386 XA.XIR[3].XIC[8].icell.Ien Iout 0.06801f
C387 XA.XIR[6].XIC[10].icell.PDM VPWR 0.01171f
C388 XA.XIR[15].XIC[1].icell.PDM VPWR 0.01512f
C389 XA.Cn[2] XA.XIR[6].XIC[2].icell.Ien 0.04604f
C390 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.Ien 0.04854f
C391 XThR.XTB5.A a_n1335_4229# 0.01243f
C392 XA.XIR[14].XIC[7].icell.PDM VPWR 0.01171f
C393 XThR.Tn[1] XA.XIR[1].XIC[10].icell.Ien 0.14211f
C394 XA.XIR[1].XIC[3].icell.Ien Iout 0.06801f
C395 XA.Cn[9] XA.XIR[13].XIC[9].icell.PDM 0.02601f
C396 XA.Cn[12] VPWR 4.5561f
C397 a_10051_9569# XA.Cn[13] 0.1927f
C398 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.Ien 0.04854f
C399 thermo15c_0.XTBN.Y XA.Cn[3] 0.49586f
C400 XA.XIR[12].XIC_15.icell.Ien Iout 0.0694f
C401 XA.XIR[5].XIC[1].icell.PDM Vbias 0.03928f
C402 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.Ien 0.04854f
C403 XA.XIR[1].XIC_dummy_left.icell.Iout XA.XIR[2].XIC_dummy_left.icell.Iout 0.03665f
C404 thermo15c_0.XTB7.B data[0] 0.0138f
C405 XA.XIR[8].XIC[11].icell.Ien Iout 0.06801f
C406 thermo15c_0.XTB2.Y thermo15c_0.XTBN.Y 0.2075f
C407 thermo15c_0.XTB3.Y a_8739_9569# 0.07285f
C408 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.Ien 0.04854f
C409 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.PDM 0.02104f
C410 XA.Cn[1] XA.XIR[8].XIC[1].icell.Ien 0.04604f
C411 XA.Cn[1] Iout 0.22482f
C412 XThR.Tn[4] Vbias 1.39526f
C413 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.Ien 0.04854f
C414 XA.XIR[12].XIC[0].icell.PDM Vbias 0.03915f
C415 XA.XIR[1].XIC[4].icell.PDM VPWR 0.01171f
C416 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.PDM 0.02104f
C417 XA.XIR[11].XIC[6].icell.PDM Vbias 0.03928f
C418 XA.XIR[6].XIC[11].icell.Ien VPWR 0.18829f
C419 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.Ien 0.04854f
C420 XA.XIR[11].XIC[12].icell.Ien Vbias 0.19161f
C421 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.Ien 0.04854f
C422 thermo15c_0.XTBN.Y VPWR 4.12335f
C423 XA.XIR[10].XIC[10].icell.PDM Vbias 0.03928f
C424 XA.XIR[15].XIC[12].icell.Ien Iout 0.07192f
C425 XA.XIR[0].XIC[13].icell.Ien Iout 0.0675f
C426 XA.XIR[4].XIC[4].icell.PDM VPWR 0.01171f
C427 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PDM 0.04042f
C428 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.Ien 0.04854f
C429 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.Ien 0.04854f
C430 XA.Cn[1] XA.XIR[3].XIC[1].icell.PDM 0.02601f
C431 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.PDM 0.02104f
C432 XA.XIR[3].XIC[12].icell.PDM VPWR 0.01171f
C433 XA.XIR[8].XIC[14].icell.PDM VPWR 0.0118f
C434 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout 0.06446f
C435 XA.XIR[12].XIC_dummy_right.icell.Iout Iout 0.01732f
C436 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.Ien 0.04854f
C437 XA.XIR[14].XIC[5].icell.Ien VPWR 0.18883f
C438 XThR.Tn[13] XA.XIR[13].XIC[12].icell.Ien 0.14211f
C439 XA.XIR[13].XIC[11].icell.PDM Vbias 0.03928f
C440 XA.XIR[13].XIC[7].icell.Ien VPWR 0.18829f
C441 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PDM 0.04035f
C442 XThR.XTB6.A XThR.XTBN.A 0.0512f
C443 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PDM 0.04035f
C444 XA.XIR[5].XIC[8].icell.Ien Vbias 0.19161f
C445 XA.Cn[9] XA.XIR[8].XIC[9].icell.Ien 0.04604f
C446 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR 0.08209f
C447 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR 0.01691f
C448 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.PDM 0.02104f
C449 XA.Cn[5] XA.XIR[11].XIC[5].icell.PDM 0.02601f
C450 XThR.XTB7.Y a_n997_1579# 0.013f
C451 XA.Cn[11] Vbias 0.82596f
C452 XA.XIR[14].XIC[1].icell.Ien Iout 0.06801f
C453 XA.Cn[10] XA.XIR[1].XIC[10].icell.Ien 0.04606f
C454 thermo15c_0.XTB4.Y XA.Cn[7] 0.01805f
C455 a_n997_1803# VPWR 0.01991f
C456 XA.XIR[2].XIC[2].icell.PDM Vbias 0.03928f
C457 XA.XIR[9].XIC_dummy_left.icell.Ien XThR.Tn[9] 0.01244f
C458 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PDM 0.0404f
C459 XA.XIR[12].XIC[3].icell.Ien Vbias 0.19161f
C460 XA.Cn[13] XA.XIR[10].XIC[13].icell.Ien 0.04604f
C461 XA.XIR[14].XIC[14].icell.Ien Vbias 0.19161f
C462 XA.XIR[6].XIC[3].icell.Ien Iout 0.06801f
C463 XA.Cn[3] XThR.Tn[13] 0.40738f
C464 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PDM 0.0404f
C465 XThR.XTB5.A data[4] 0.14415f
C466 XA.XIR[2].XIC[14].icell.Ien VPWR 0.18835f
C467 XA.Cn[13] XA.XIR[12].XIC[13].icell.PDM 0.02601f
C468 thermo15c_0.XTB7.A thermo15c_0.XTB7.B 0.35844f
C469 XA.Cn[13] XA.XIR[4].XIC[13].icell.Ien 0.04604f
C470 thermo15c_0.XTB3.Y thermo15c_0.XTB5.Y 0.04438f
C471 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.PDM 0.02104f
C472 XA.Cn[4] XA.XIR[9].XIC[4].icell.Ien 0.04604f
C473 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.Ien 0.04854f
C474 XThR.Tn[8] XA.XIR[8].XIC[11].icell.Ien 0.14211f
C475 XA.XIR[14].XIC[0].icell.Ien VPWR 0.18883f
C476 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.Ien 0.04854f
C477 XA.Cn[0] XThR.Tn[9] 0.40738f
C478 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.Ien 0.04854f
C479 XA.Cn[1] XThR.Tn[8] 0.40738f
C480 XThR.Tn[13] VPWR 9.0331f
C481 XA.XIR[11].XIC[10].icell.Ien Vbias 0.19161f
C482 XA.XIR[7].XIC_dummy_left.icell.Iout Iout 0.03553f
C483 XA.XIR[2].XIC[1].icell.Ien Iout 0.06801f
C484 XA.XIR[11].XIC[2].icell.Ien Iout 0.06801f
C485 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.PDM 0.02104f
C486 XA.XIR[15].XIC[10].icell.Ien Iout 0.07192f
C487 XA.Cn[1] XA.XIR[11].XIC[1].icell.Ien 0.04604f
C488 XA.Cn[12] XA.XIR[1].XIC[12].icell.PDM 0.02602f
C489 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.PDM 0.02104f
C490 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.PDM 0.02104f
C491 XA.XIR[10].XIC[4].icell.Ien Iout 0.06801f
C492 XThR.Tn[5] XA.XIR[5].XIC[10].icell.Ien 0.14211f
C493 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.Ien 0.04854f
C494 XA.Cn[12] XA.XIR[4].XIC[12].icell.PDM 0.02601f
C495 XThR.Tn[13] XA.XIR[13].XIC[10].icell.Ien 0.14211f
C496 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.PDM 0.02104f
C497 XA.XIR[5].XIC[4].icell.Ien VPWR 0.18829f
C498 XA.Cn[0] XA.XIR[15].XIC[0].icell.Ien 0.04292f
C499 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.PDM 0.02104f
C500 XA.XIR[3].XIC[13].icell.Ien Iout 0.06801f
C501 XThR.Tn[3] a_n1049_6699# 0.27008f
C502 VPWR data[6] 0.21221f
C503 XA.XIR[11].XIC[0].icell.Ien Vbias 0.19149f
C504 XA.Cn[10] XA.XIR[6].XIC[10].icell.Ien 0.04604f
C505 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.PDM 0.02104f
C506 XThR.Tn[1] XA.XIR[1].XIC_15.icell.Ien 0.13564f
C507 XA.XIR[2].XIC[6].icell.Ien Iout 0.06801f
C508 XA.XIR[7].XIC[2].icell.PDM Vbias 0.03928f
C509 XA.Cn[8] XA.XIR[11].XIC[8].icell.PDM 0.02601f
C510 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.PDM 0.02104f
C511 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.PDM 0.02104f
C512 XA.Cn[2] XA.XIR[8].XIC[2].icell.PDM 0.02601f
C513 XA.XIR[1].XIC[8].icell.Ien Iout 0.06801f
C514 XThR.XTB6.A XThR.XTB6.Y 0.10153f
C515 XA.XIR[15].XIC[0].icell.PDM Vbias 0.03915f
C516 XA.XIR[9].XIC[14].icell.PDM VPWR 0.0118f
C517 XA.XIR[6].XIC[9].icell.PDM Vbias 0.03928f
C518 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.PDM 0.02104f
C519 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.Ien 0.04854f
C520 XA.XIR[0].XIC[6].icell.PDM VPWR 0.01138f
C521 XA.XIR[14].XIC[6].icell.PDM Vbias 0.03928f
C522 XA.XIR[1].XIC_dummy_left.icell.Iout VPWR 0.11048f
C523 XA.XIR[14].XIC[12].icell.Ien Vbias 0.19161f
C524 XA.Cn[14] XThR.Tn[3] 0.40742f
C525 XA.XIR[13].XIC[10].icell.PDM Vbias 0.03928f
C526 XA.Cn[8] data[0] 0.01744f
C527 thermo15c_0.XTB5.Y a_9827_9569# 0.06458f
C528 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.Ien 0.04854f
C529 XA.Cn[8] XA.XIR[15].XIC[8].icell.Ien 0.04292f
C530 XA.Cn[5] XA.Cn[6] 0.14629f
C531 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PDM 0.04035f
C532 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PDM 0.0404f
C533 thermo15c_0.XTB1.Y thermo15c_0.XTB6.Y 0.05752f
C534 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PDM 0.04035f
C535 thermo15c_0.XTB2.Y thermo15c_0.XTBN.A 0.04716f
C536 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.PDM 0.02104f
C537 XA.XIR[9].XIC[4].icell.Ien Vbias 0.19161f
C538 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.PDM 0.02104f
C539 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR 0.08209f
C540 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR 0.01691f
C541 XA.Cn[5] XA.XIR[14].XIC[5].icell.PDM 0.02601f
C542 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.PDM 0.02104f
C543 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout 0.06446f
C544 XA.XIR[1].XIC[3].icell.PDM Vbias 0.03928f
C545 XA.Cn[11] XThR.Tn[0] 0.40763f
C546 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.Ien 0.04854f
C547 thermo15c_0.XTBN.A VPWR 0.88815f
C548 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Ien 0.01263f
C549 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR 0.38999f
C550 XA.XIR[4].XIC[3].icell.PDM Vbias 0.03928f
C551 XA.XIR[5].XIC[13].icell.Ien Vbias 0.19161f
C552 XThR.Tn[3] Iout 1.12764f
C553 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.04035f
C554 XThR.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.14211f
C555 XA.Cn[13] XA.XIR[13].XIC[13].icell.Ien 0.04604f
C556 thermo15c_0.XTB7.Y XA.Cn[12] 0.07091f
C557 XA.XIR[3].XIC[11].icell.PDM Vbias 0.03928f
C558 XA.XIR[8].XIC[13].icell.PDM Vbias 0.03928f
C559 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.PDM 0.02104f
C560 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.Ien 0.04854f
C561 XThR.XTBN.A XThR.Tn[12] 0.22096f
C562 XA.XIR[11].XIC_15.icell.PDM Vbias 0.03927f
C563 XA.Cn[3] XA.XIR[12].XIC[3].icell.PDM 0.02601f
C564 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.PDM 0.02104f
C565 XA.XIR[11].XIC_15.icell.Ien Vbias 0.19195f
C566 XA.XIR[8].XIC_dummy_left.icell.Iout Iout 0.03553f
C567 XA.XIR[12].XIC[8].icell.Ien Vbias 0.19161f
C568 XA.Cn[13] XA.XIR[15].XIC[13].icell.PDM 0.02601f
C569 XA.Cn[6] XA.XIR[10].XIC[6].icell.Ien 0.04604f
C570 XThR.XTB2.Y a_n997_3755# 0.06476f
C571 XA.XIR[15].XIC_15.icell.Ien Iout 0.0733f
C572 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.Ien 0.04854f
C573 XA.XIR[6].XIC[8].icell.Ien Iout 0.06801f
C574 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PDM 0.04035f
C575 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.PDM 0.02104f
C576 XA.XIR[5].XIC[4].icell.PDM VPWR 0.01171f
C577 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout 0.06446f
C578 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.PDM 0.02104f
C579 XThR.XTBN.Y a_n1049_8581# 0.0607f
C580 XThR.Tn[13] XA.XIR[13].XIC_15.icell.Ien 0.13564f
C581 thermo15c_0.XTB7.Y thermo15c_0.XTBN.Y 0.50018f
C582 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.PDM 0.02104f
C583 XA.XIR[6].XIC_dummy_left.icell.Iout VPWR 0.11008f
C584 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PDM 0.04056f
C585 XA.XIR[14].XIC[10].icell.Ien Vbias 0.19161f
C586 XA.XIR[14].XIC[2].icell.Ien Iout 0.06801f
C587 XA.XIR[12].XIC[3].icell.PDM VPWR 0.01171f
C588 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.Ien 0.04854f
C589 XA.Cn[1] XA.XIR[14].XIC[1].icell.Ien 0.04604f
C590 XA.XIR[13].XIC[4].icell.Ien Iout 0.06801f
C591 XA.Cn[12] XA.XIR[9].XIC[12].icell.Ien 0.04604f
C592 XA.Cn[7] Vbias 0.82088f
C593 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.PDM 0.02104f
C594 XA.Cn[9] XThR.Tn[2] 0.40741f
C595 XA.XIR[11].XIC[9].icell.PDM VPWR 0.01171f
C596 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.Ien 0.04854f
C597 XA.Cn[2] XA.XIR[9].XIC[2].icell.PDM 0.02601f
C598 XA.XIR[15].XIC_dummy_right.icell.Iout Iout 0.01732f
C599 XA.XIR[11].XIC[7].icell.Ien Iout 0.06801f
C600 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PDM 0.04035f
C601 XA.XIR[4].XIC[1].icell.Ien Vbias 0.19161f
C602 XA.XIR[10].XIC[9].icell.Ien Iout 0.06801f
C603 XThR.Tn[5] XA.XIR[5].XIC_15.icell.Ien 0.13564f
C604 XA.Cn[8] XA.XIR[14].XIC[8].icell.PDM 0.02601f
C605 XThR.XTB3.Y a_n997_2891# 0.07285f
C606 XA.XIR[5].XIC[9].icell.Ien VPWR 0.18829f
C607 XA.Cn[14] XThR.Tn[11] 0.40742f
C608 XThR.Tn[4] XA.XIR[4].XIC[0].icell.Ien 0.1423f
C609 XA.Cn[7] XA.XIR[10].XIC[7].icell.PDM 0.02601f
C610 XA.XIR[8].XIC[1].icell.PDM VPWR 0.01171f
C611 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10] 0.14211f
C612 XA.Cn[10] XThR.Tn[6] 0.40738f
C613 a_n1049_5317# XThR.Tn[6] 0.26047f
C614 XA.XIR[2].XIC[5].icell.PDM VPWR 0.01171f
C615 XThR.Tn[3] XA.XIR[3].XIC[0].icell.Ien 0.14251f
C616 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout 0.06446f
C617 XA.XIR[15].XIC[3].icell.Ien Vbias 0.15966f
C618 XA.XIR[2].XIC[11].icell.Ien Iout 0.06801f
C619 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.PDM 0.02104f
C620 XA.XIR[12].XIC[4].icell.Ien VPWR 0.18829f
C621 XA.Cn[1] XA.XIR[2].XIC[1].icell.Ien 0.04605f
C622 XA.XIR[1].XIC[13].icell.Ien Iout 0.06801f
C623 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout 0.06446f
C624 XA.Cn[7] XA.XIR[5].XIC[7].icell.Ien 0.04604f
C625 XA.XIR[4].XIC[6].icell.Ien Vbias 0.19161f
C626 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.PDM 0.02104f
C627 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.Ien 0.04854f
C628 a_n997_3979# VPWR 0.01662f
C629 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PDM 0.04035f
C630 XThR.XTB7.Y XThR.Tn[8] 0.07806f
C631 XThR.Tn[8] XA.XIR[8].XIC_dummy_left.icell.Iout 0.03962f
C632 XA.XIR[9].XIC_15.icell.PUM VPWR 0.01655f
C633 XThR.Tn[4] XA.XIR[4].XIC[5].icell.Ien 0.14211f
C634 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR 0.01604f
C635 XA.XIR[12].XIC[0].icell.Ien Iout 0.06795f
C636 XThR.XTB6.Y XThR.Tn[12] 0.02431f
C637 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.Ien 0.04854f
C638 XA.XIR[9].XIC[13].icell.PDM Vbias 0.03928f
C639 XA.XIR[0].XIC[5].icell.PDM Vbias 0.03945f
C640 XA.XIR[7].XIC[0].icell.Ien Vbias 0.19149f
C641 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.Ien 0.04854f
C642 XThR.Tn[11] Iout 1.12764f
C643 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PDM 0.04035f
C644 XA.Cn[12] XA.XIR[5].XIC[12].icell.PDM 0.02601f
C645 thermo15c_0.XTB7.B a_7875_9569# 0.01174f
C646 XA.Cn[11] XThR.Tn[1] 0.40744f
C647 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PDM 0.04035f
C648 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.PDM 0.02104f
C649 XA.XIR[9].XIC[9].icell.Ien Vbias 0.19161f
C650 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PDM 0.04035f
C651 thermo15c_0.XTB7.A thermo15c_0.XTB4.Y 0.14536f
C652 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR 0.38939f
C653 XA.XIR[0].XIC[2].icell.Ien Vbias 0.19213f
C654 XA.Cn[9] XA.XIR[2].XIC[9].icell.Ien 0.04605f
C655 XA.Cn[3] XThR.Tn[7] 0.40738f
C656 XA.Cn[11] XThR.Tn[12] 0.40738f
C657 XA.XIR[11].XIC[14].icell.PDM Vbias 0.03928f
C658 XA.Cn[14] XA.XIR[10].XIC[14].icell.Ien 0.04604f
C659 a_6243_9615# VPWR 0.7055f
C660 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.04035f
C661 XA.XIR[14].XIC_15.icell.PDM Vbias 0.03927f
C662 XA.Cn[3] XA.XIR[15].XIC[3].icell.PDM 0.02601f
C663 XA.XIR[14].XIC_15.icell.Ien Vbias 0.19195f
C664 XThR.Tn[12] XA.XIR[12].XIC[3].icell.Ien 0.14211f
C665 XA.XIR[7].XIC[5].icell.Ien Vbias 0.19161f
C666 XA.Cn[13] XA.XIR[0].XIC[13].icell.PDM 0.0279f
C667 XA.Cn[6] XA.XIR[13].XIC[6].icell.Ien 0.04604f
C668 XA.Cn[10] XThR.Tn[4] 0.40738f
C669 XThR.Tn[3] XA.XIR[3].XIC[8].icell.Ien 0.14211f
C670 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.Ien 0.04854f
C671 XThR.Tn[7] VPWR 8.3986f
C672 a_n997_2891# VPWR 0.01347f
C673 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PDM 0.04035f
C674 XA.XIR[7].XIC[5].icell.PDM VPWR 0.01171f
C675 XA.Cn[9] XThR.Tn[10] 0.40738f
C676 XThR.Tn[2] XA.XIR[2].XIC[3].icell.Ien 0.14211f
C677 XA.Cn[10] XA.XIR[10].XIC[10].icell.PDM 0.02601f
C678 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout 0.06446f
C679 XA.Cn[1] XA.XIR[6].XIC[1].icell.PDM 0.02601f
C680 XA.Cn[4] XA.XIR[2].XIC[4].icell.PDM 0.02602f
C681 XThR.XTB6.Y a_n1049_5317# 0.01199f
C682 XA.XIR[4].XIC[2].icell.Ien VPWR 0.18829f
C683 XA.XIR[15].XIC[3].icell.PDM VPWR 0.01512f
C684 XA.XIR[6].XIC[12].icell.PDM VPWR 0.01171f
C685 XA.XIR[3].XIC_dummy_right.icell.Iout XA.XIR[4].XIC_dummy_right.icell.Iout 0.04047f
C686 XA.XIR[6].XIC[13].icell.Ien Iout 0.06801f
C687 XA.XIR[10].XIC[14].icell.Ien Iout 0.06801f
C688 XA.XIR[14].XIC[9].icell.PDM VPWR 0.01171f
C689 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.Ien 0.04854f
C690 XA.Cn[7] XThR.Tn[0] 0.40759f
C691 XA.Cn[1] XThR.Tn[3] 0.40738f
C692 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.Ien 0.04854f
C693 XA.XIR[9].XIC[1].icell.PDM VPWR 0.01171f
C694 XA.XIR[14].XIC[7].icell.Ien Iout 0.06801f
C695 XA.Cn[10] XA.Cn[11] 0.07237f
C696 XA.XIR[5].XIC[3].icell.PDM Vbias 0.03928f
C697 thermo15c_0.XTBN.A thermo15c_0.XTB7.Y 1.11562f
C698 XA.XIR[13].XIC[9].icell.Ien Iout 0.06801f
C699 XA.XIR[9].XIC[5].icell.Ien VPWR 0.18829f
C700 XA.Cn[2] XThR.Tn[5] 0.40738f
C701 XThR.XTBN.Y a_n1049_7787# 0.08456f
C702 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.Ien 0.04854f
C703 XA.Cn[7] XA.XIR[13].XIC[7].icell.PDM 0.02601f
C704 XA.Cn[14] XThR.Tn[14] 0.40742f
C705 XA.XIR[12].XIC[2].icell.PDM Vbias 0.03928f
C706 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PDM 0.0404f
C707 XThR.XTB2.Y XThR.XTB7.Y 0.0437f
C708 XA.XIR[1].XIC[6].icell.PDM VPWR 0.01171f
C709 XA.XIR[11].XIC[8].icell.PDM Vbias 0.03928f
C710 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11] 0.14211f
C711 XA.XIR[5].XIC_dummy_left.icell.Iout XA.XIR[6].XIC_dummy_left.icell.Iout 0.03665f
C712 a_n1049_6405# XThR.Tn[4] 0.26564f
C713 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR 0.01604f
C714 XA.XIR[4].XIC[6].icell.PDM VPWR 0.01171f
C715 thermo15c_0.XTBN.Y XA.Cn[9] 0.39932f
C716 XA.XIR[5].XIC[14].icell.Ien VPWR 0.18835f
C717 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PDM 0.04035f
C718 XA.XIR[3].XIC[2].icell.Ien Vbias 0.19161f
C719 XA.XIR[3].XIC[14].icell.PDM VPWR 0.0118f
C720 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR 0.08209f
C721 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.PDM 0.02104f
C722 XA.XIR[12].XIC_15.icell.PUM VPWR 0.01655f
C723 thermo15c_0.XTB7.A XA.Cn[4] 0.02779f
C724 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PDM 0.04035f
C725 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PDM 0.04035f
C726 XA.XIR[15].XIC[8].icell.Ien Vbias 0.15966f
C727 XA.Cn[5] XThR.Tn[2] 0.40741f
C728 XA.XIR[5].XIC[1].icell.Ien Iout 0.06801f
C729 XA.Cn[10] XA.XIR[11].XIC[10].icell.Ien 0.04604f
C730 XA.XIR[12].XIC[9].icell.Ien VPWR 0.18829f
C731 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.Ien 0.04854f
C732 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR 0.01604f
C733 XA.XIR[4].XIC[11].icell.Ien Vbias 0.19161f
C734 XA.XIR[8].XIC[0].icell.PDM Vbias 0.03915f
C735 XThR.Tn[14] Iout 1.12763f
C736 XA.Cn[4] XA.XIR[7].XIC[4].icell.PDM 0.02601f
C737 XA.XIR[11].XIC[13].icell.PDM Vbias 0.03928f
C738 XA.XIR[2].XIC[4].icell.PDM Vbias 0.03928f
C739 XA.XIR[8].XIC[5].icell.Ien Vbias 0.19161f
C740 XA.XIR[10].XIC[12].icell.Ien Iout 0.06801f
C741 XA.XIR[9].XIC[0].icell.Ien VPWR 0.18829f
C742 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PDM 0.04035f
C743 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Iout 0.01828f
C744 XThR.Tn[4] XA.XIR[4].XIC[10].icell.Ien 0.14211f
C745 XA.XIR[14].XIC[14].icell.PDM Vbias 0.03928f
C746 XThR.Tn[0] XA.XIR[0].XIC[2].icell.Ien 0.14211f
C747 XA.Cn[14] XA.XIR[13].XIC[14].icell.Ien 0.04604f
C748 XA.Cn[7] XA.XIR[12].XIC[7].icell.Ien 0.04604f
C749 XA.XIR[9].XIC[14].icell.Ien Vbias 0.19161f
C750 XA.XIR[5].XIC[6].icell.Ien Iout 0.06801f
C751 XA.Cn[6] XThR.Tn[6] 0.40738f
C752 data[6] data[7] 0.04128f
C753 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PDM 0.04035f
C754 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.Ien 0.04854f
C755 XThR.Tn[7] XA.XIR[7].XIC[3].icell.Ien 0.14211f
C756 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR 0.01691f
C757 XA.XIR[0].XIC[7].icell.Ien Vbias 0.19213f
C758 a_n997_1579# VPWR 0.02417f
C759 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout 0.06446f
C760 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.PDM 0.02104f
C761 XA.Cn[5] XA.XIR[11].XIC[5].icell.Ien 0.04604f
C762 XA.XIR[7].XIC[10].icell.Ien Vbias 0.19161f
C763 XA.Cn[10] XA.XIR[13].XIC[10].icell.PDM 0.02601f
C764 XThR.Tn[12] XA.XIR[12].XIC[8].icell.Ien 0.14211f
C765 XA.Cn[9] XThR.Tn[13] 0.40738f
C766 XA.XIR[10].XIC[0].icell.PDM VPWR 0.01171f
C767 XA.XIR[2].XIC_dummy_left.icell.Iout Iout 0.03553f
C768 XA.XIR[7].XIC_dummy_left.icell.Iout XA.XIR[8].XIC_dummy_left.icell.Iout 0.03665f
C769 XThR.Tn[3] XA.XIR[3].XIC[13].icell.Ien 0.14211f
C770 a_10915_9569# XA.Cn[14] 0.20879f
C771 bias[1] bias[0] 0.56718f
C772 XA.Cn[1] XThR.Tn[11] 0.40738f
C773 XA.XIR[13].XIC[14].icell.Ien Iout 0.06801f
C774 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.Ien 0.04854f
C775 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout 0.06446f
C776 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.Ien 0.04854f
C777 XA.XIR[15].XIC[4].icell.Ien VPWR 0.31713f
C778 XA.Cn[7] XThR.Tn[1] 0.40744f
C779 XA.XIR[8].XIC[0].icell.Ien Vbias 0.19149f
C780 XThR.Tn[2] XA.XIR[2].XIC[8].icell.Ien 0.14211f
C781 thermo15c_0.XTB7.A Vbias 0.0148f
C782 XA.XIR[4].XIC[7].icell.Ien VPWR 0.18829f
C783 XThR.Tn[9] XA.XIR[9].XIC[1].icell.Ien 0.14211f
C784 XA.Cn[7] XThR.Tn[12] 0.40738f
C785 XThR.XTB7.Y a_n997_715# 0.06874f
C786 XA.Cn[3] XA.XIR[0].XIC[3].icell.Ien 0.04658f
C787 XA.XIR[7].XIC[4].icell.PDM Vbias 0.03928f
C788 XA.Cn[2] XA.XIR[3].XIC[2].icell.PDM 0.02601f
C789 XA.XIR[3].XIC_dummy_left.icell.Iout XA.XIR[4].XIC_dummy_left.icell.Iout 0.03665f
C790 XA.XIR[15].XIC[2].icell.PDM Vbias 0.03928f
C791 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR 0.08209f
C792 XA.XIR[6].XIC[11].icell.PDM Vbias 0.03928f
C793 XA.XIR[10].XIC[10].icell.Ien Iout 0.06801f
C794 XA.XIR[7].XIC[1].icell.Ien VPWR 0.18829f
C795 thermo15c_0.XTB7.Y a_6243_9615# 0.27822f
C796 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13] 0.14211f
C797 XA.XIR[0].XIC[8].icell.PDM VPWR 0.01451f
C798 XA.Cn[6] XThR.Tn[4] 0.40738f
C799 XA.XIR[14].XIC[8].icell.PDM Vbias 0.03928f
C800 XA.XIR[9].XIC[10].icell.Ien VPWR 0.18829f
C801 XA.XIR[12].XIC[14].icell.Ien VPWR 0.18835f
C802 XA.Cn[6] XA.XIR[11].XIC[6].icell.PDM 0.02601f
C803 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.Ien 0.04854f
C804 XThR.Tn[9] XA.XIR[9].XIC[6].icell.Ien 0.14211f
C805 XA.XIR[9].XIC[0].icell.PDM Vbias 0.03915f
C806 XA.XIR[0].XIC[3].icell.Ien VPWR 0.18776f
C807 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PDM 0.04035f
C808 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PDM 0.04035f
C809 XA.Cn[5] XThR.Tn[10] 0.40738f
C810 VPWR data[5] 0.4402f
C811 XA.XIR[11].XIC[12].icell.PDM Vbias 0.03928f
C812 XA.XIR[7].XIC[6].icell.Ien VPWR 0.18829f
C813 XA.Cn[10] XA.XIR[14].XIC[10].icell.Ien 0.04604f
C814 XA.XIR[3].XIC[7].icell.Ien Vbias 0.19161f
C815 XA.XIR[1].XIC[5].icell.PDM Vbias 0.03928f
C816 XA.XIR[14].XIC[13].icell.PDM Vbias 0.03928f
C817 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.PDM 0.02104f
C818 XThR.XTB7.A XThR.XTBN.A 0.19736f
C819 a_n1049_6699# VPWR 0.72162f
C820 thermo15c_0.XTBN.A XA.Cn[9] 0.12399f
C821 XA.XIR[13].XIC[12].icell.Ien Iout 0.06801f
C822 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.PDM 0.02104f
C823 XA.XIR[4].XIC[5].icell.PDM Vbias 0.03928f
C824 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR 0.01691f
C825 XA.Cn[8] XA.XIR[10].XIC[8].icell.Ien 0.04604f
C826 XThR.XTB7.A XThR.Tn[6] 0.1056f
C827 XA.XIR[3].XIC[13].icell.PDM Vbias 0.03928f
C828 XA.XIR[1].XIC[2].icell.Ien Vbias 0.19173f
C829 XA.XIR[8].XIC_15.icell.PDM Vbias 0.03927f
C830 XA.XIR[9].XIC[2].icell.Ien Iout 0.06801f
C831 XThR.Tn[11] XA.XIR[11].XIC[2].icell.Ien 0.14211f
C832 XA.XIR[8].XIC[10].icell.Ien Vbias 0.19161f
C833 XThR.Tn[4] XA.XIR[4].XIC_15.icell.Ien 0.13564f
C834 XA.Cn[14] VPWR 4.55561f
C835 XA.Cn[13] XA.XIR[1].XIC[13].icell.PDM 0.02602f
C836 XThR.Tn[0] XA.XIR[0].XIC[7].icell.Ien 0.14211f
C837 XThR.Tn[10] XA.XIR[10].XIC[6].icell.Ien 0.14211f
C838 thermo15c_0.XTBN.Y XA.Cn[5] 0.49425f
C839 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR 0.08221f
C840 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PDM 0.04035f
C841 XA.XIR[5].XIC[6].icell.PDM VPWR 0.01171f
C842 XA.XIR[5].XIC[11].icell.Ien Iout 0.06801f
C843 XA.Cn[13] XA.XIR[4].XIC[13].icell.PDM 0.02601f
C844 XA.Cn[3] Iout 0.22443f
C845 XA.Cn[5] XA.XIR[14].XIC[5].icell.Ien 0.04604f
C846 XA.XIR[13].XIC[0].icell.PDM VPWR 0.01171f
C847 XA.Cn[3] XA.XIR[3].XIC[3].icell.Ien 0.04604f
C848 XA.Cn[1] XA.XIR[5].XIC[1].icell.Ien 0.04604f
C849 XA.XIR[0].XIC[12].icell.Ien Vbias 0.19213f
C850 thermo15c_0.XTB6.Y a_10051_9569# 0.07626f
C851 XThR.Tn[7] XA.XIR[7].XIC[8].icell.Ien 0.14211f
C852 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.PDM 0.02104f
C853 XA.XIR[12].XIC[5].icell.PDM VPWR 0.01171f
C854 XA.Cn[1] XThR.Tn[14] 0.40738f
C855 XA.XIR[12].XIC[12].icell.Ien VPWR 0.18829f
C856 thermo15c_0.XTB1.Y thermo15c_0.XTB7.B 1.61695f
C857 thermo15c_0.XTB2.Y thermo15c_0.XTB5.Y 0.0451f
C858 XA.Cn[9] XA.XIR[11].XIC[9].icell.PDM 0.02601f
C859 XA.XIR[12].XIC[6].icell.Ien Iout 0.06801f
C860 XA.XIR[7].XIC_15.icell.Ien Vbias 0.19195f
C861 XA.Cn[3] XA.XIR[8].XIC[3].icell.PDM 0.02601f
C862 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.Ien 0.04854f
C863 XA.XIR[8].XIC[1].icell.Ien VPWR 0.18829f
C864 XA.XIR[10].XIC_15.icell.Ien Iout 0.0694f
C865 XA.XIR[5].XIC[0].icell.Ien Vbias 0.19149f
C866 VPWR Iout 57.8523f
C867 XA.XIR[3].XIC[3].icell.Ien VPWR 0.18829f
C868 XA.XIR[15].XIC_15.icell.PUM VPWR 0.01655f
C869 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PDM 0.04035f
C870 thermo15c_0.XTB5.Y VPWR 1.01219f
C871 XThR.XTB7.A XThR.Tn[4] 0.02736f
C872 XA.XIR[15].XIC[9].icell.Ien VPWR 0.31713f
C873 XThR.Tn[2] XA.XIR[2].XIC[13].icell.Ien 0.14211f
C874 XA.Cn[13] Vbias 0.82511f
C875 XA.Cn[9] XA.XIR[5].XIC[9].icell.Ien 0.04604f
C876 XA.XIR[13].XIC[10].icell.Ien Iout 0.06801f
C877 XThR.XTB7.A a_n1049_7493# 0.0127f
C878 XA.XIR[3].XIC[1].icell.PDM VPWR 0.01171f
C879 XA.XIR[4].XIC[12].icell.Ien VPWR 0.18829f
C880 XA.XIR[8].XIC[3].icell.PDM VPWR 0.01171f
C881 XA.XIR[6].XIC[2].icell.Ien Vbias 0.19161f
C882 XA.XIR[2].XIC[7].icell.PDM VPWR 0.01171f
C883 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14] 0.14211f
C884 XA.Cn[2] XA.XIR[7].XIC[2].icell.Ien 0.04604f
C885 XA.XIR[8].XIC[6].icell.Ien VPWR 0.18829f
C886 XA.Cn[6] XA.XIR[14].XIC[6].icell.PDM 0.02601f
C887 XThR.XTB7.A XThR.XTB6.Y 0.19112f
C888 XA.Cn[11] XA.XIR[0].XIC[11].icell.Ien 0.04662f
C889 XA.Cn[7] XA.XIR[15].XIC[7].icell.Ien 0.04292f
C890 XA.XIR[10].XIC_dummy_right.icell.Iout Iout 0.01732f
C891 XA.XIR[11].XIC[11].icell.PDM Vbias 0.03928f
C892 XA.Cn[5] XThR.Tn[13] 0.40738f
C893 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PDM 0.04035f
C894 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.Ien 0.04854f
C895 XA.XIR[9].XIC_15.icell.Ien VPWR 0.26829f
C896 thermo15c_0.XTBN.Y a_3773_9615# 0.08456f
C897 XA.XIR[14].XIC[12].icell.PDM Vbias 0.03928f
C898 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.PDM 0.02104f
C899 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.PDM 0.02104f
C900 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR 0.01604f
C901 XThR.XTB7.B XThR.XTBN.A 0.35142f
C902 XA.XIR[9].XIC_15.icell.PDM Vbias 0.03927f
C903 XThR.Tn[9] XA.XIR[9].XIC[11].icell.Ien 0.14211f
C904 XThR.XTB7.Y XThR.Tn[11] 0.07412f
C905 XA.XIR[0].XIC[8].icell.Ien VPWR 0.18959f
C906 XA.XIR[0].XIC[7].icell.PDM Vbias 0.03945f
C907 XA.Cn[11] XA.XIR[11].XIC[11].icell.Ien 0.04604f
C908 thermo15c_0.XTB7.B a_8963_9569# 0.02071f
C909 XThR.XTB7.B XThR.Tn[6] 0.04822f
C910 XA.Cn[2] XThR.Tn[9] 0.40738f
C911 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PDM 0.04035f
C912 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.PDM 0.02104f
C913 XA.Cn[3] XThR.Tn[8] 0.40738f
C914 XA.XIR[10].XIC[3].icell.Ien Vbias 0.19161f
C915 XA.XIR[12].XIC[10].icell.Ien VPWR 0.18829f
C916 XA.Cn[4] XA.XIR[12].XIC[4].icell.PDM 0.02601f
C917 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PDM 0.04035f
C918 XA.Cn[8] XA.XIR[13].XIC[8].icell.Ien 0.04604f
C919 XA.XIR[7].XIC[11].icell.Ien VPWR 0.18829f
C920 XA.XIR[4].XIC[4].icell.Ien Iout 0.06801f
C921 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.Ien 0.04854f
C922 XA.XIR[3].XIC[12].icell.Ien Vbias 0.19161f
C923 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.Ien 0.04854f
C924 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PDM 0.04035f
C925 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.Ien 0.04854f
C926 XA.XIR[9].XIC_dummy_right.icell.Iout VPWR 0.11567f
C927 XThR.Tn[6] XA.XIR[6].XIC[1].icell.Ien 0.14211f
C928 XA.XIR[2].XIC[5].icell.Ien Vbias 0.19161f
C929 XA.XIR[3].XIC[0].icell.Ien VPWR 0.18829f
C930 XThR.Tn[8] VPWR 8.93422f
C931 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.PDM 0.02104f
C932 XA.Cn[12] XA.XIR[10].XIC[12].icell.PDM 0.02601f
C933 XA.XIR[1].XIC[7].icell.Ien Vbias 0.19173f
C934 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR 0.08221f
C935 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.PDM 0.02104f
C936 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.PDM 0.02104f
C937 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.Ien 0.04854f
C938 XA.XIR[9].XIC[7].icell.Ien Iout 0.06801f
C939 XA.Cn[9] XThR.Tn[7] 0.40738f
C940 XThR.Tn[11] XA.XIR[11].XIC[7].icell.Ien 0.14211f
C941 XA.XIR[11].XIC[1].icell.Ien VPWR 0.18829f
C942 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PDM 0.04035f
C943 XA.XIR[8].XIC_15.icell.Ien Vbias 0.19195f
C944 XA.Cn[3] XA.XIR[9].XIC[3].icell.PDM 0.02601f
C945 XA.XIR[7].XIC[7].icell.PDM VPWR 0.01171f
C946 XThR.XTB2.Y XThR.XTB3.Y 2.04808f
C947 XThR.Tn[14] a_n997_715# 0.1927f
C948 XA.XIR[6].XIC[14].icell.PDM VPWR 0.0118f
C949 XA.XIR[15].XIC[5].icell.PDM VPWR 0.01512f
C950 XThR.Tn[0] XA.XIR[0].XIC[12].icell.Ien 0.14211f
C951 XThR.Tn[11] a_n997_2667# 0.19413f
C952 XThR.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.14211f
C953 XA.XIR[9].XIC_dummy_right.icell.Iout XA.XIR[10].XIC_dummy_right.icell.Iout 0.04047f
C954 XA.Cn[9] XA.XIR[14].XIC[9].icell.PDM 0.02601f
C955 XA.XIR[7].XIC[3].icell.Ien Iout 0.06801f
C956 XA.XIR[15].XIC[14].icell.Ien VPWR 0.31908f
C957 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Ien 0.01569f
C958 XA.Cn[6] XA.Cn[7] 0.0974f
C959 XA.XIR[13].XIC_15.icell.Ien Iout 0.0694f
C960 XThR.Tn[7] XA.XIR[7].XIC[13].icell.Ien 0.14211f
C961 XA.XIR[9].XIC[3].icell.PDM VPWR 0.01171f
C962 XA.Cn[11] XA.XIR[3].XIC[11].icell.Ien 0.04604f
C963 XA.XIR[5].XIC[5].icell.PDM Vbias 0.03928f
C964 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.Ien 0.04854f
C965 XA.Cn[2] XA.XIR[8].XIC[2].icell.Ien 0.04604f
C966 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.Ien 0.04854f
C967 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.Ien 0.04854f
C968 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.PDM 0.02104f
C969 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.PDM 0.02104f
C970 XA.Cn[3] XA.XIR[1].XIC[3].icell.Ien 0.04607f
C971 thermo15c_0.XTB1.Y XA.Cn[8] 0.29214f
C972 thermo15c_0.XTB6.A data[0] 0.48493f
C973 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.PDM 0.02104f
C974 XA.XIR[12].XIC[4].icell.PDM Vbias 0.03928f
C975 XA.Cn[13] XThR.Tn[0] 0.40764f
C976 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PDM 0.04035f
C977 XThR.XTB7.B XThR.XTB6.Y 0.30244f
C978 XA.XIR[3].XIC[8].icell.Ien VPWR 0.18829f
C979 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.Ien 0.04854f
C980 XA.XIR[1].XIC[8].icell.PDM VPWR 0.01171f
C981 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.PDM 0.02104f
C982 XA.XIR[11].XIC[10].icell.PDM Vbias 0.03928f
C983 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.Ien 0.04854f
C984 XA.XIR[4].XIC[8].icell.PDM VPWR 0.01171f
C985 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout 0.06446f
C986 XA.XIR[13].XIC_dummy_right.icell.Iout Iout 0.01732f
C987 thermo15c_0.XTB7.Y XA.Cn[14] 0.4237f
C988 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PDM 0.04035f
C989 thermo15c_0.XTB2.Y XA.Cn[1] 0.18085f
C990 XA.XIR[14].XIC[11].icell.PDM Vbias 0.03928f
C991 XThR.XTBN.Y XThR.XTBN.A 0.77119f
C992 XA.Cn[8] XThR.Tn[5] 0.40738f
C993 XA.Cn[0] XA.XIR[0].XIC[0].icell.PDM 0.02804f
C994 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.PDM 0.02104f
C995 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR 0.08209f
C996 XA.XIR[1].XIC[3].icell.Ien VPWR 0.18829f
C997 XA.Cn[13] XA.XIR[5].XIC[13].icell.PDM 0.02601f
C998 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.Ien 0.04854f
C999 XA.XIR[6].XIC[7].icell.Ien Vbias 0.19161f
C1000 a_n1049_7493# XThR.Tn[2] 0.26564f
C1001 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.Ien 0.04854f
C1002 XA.Cn[6] XA.XIR[4].XIC[6].icell.Ien 0.04604f
C1003 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.Ien 0.04854f
C1004 XA.XIR[12].XIC_15.icell.Ien VPWR 0.26829f
C1005 XThR.XTBN.Y XThR.Tn[6] 0.59897f
C1006 XThR.XTB1.Y data[4] 0.06453f
C1007 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PDM 0.04035f
C1008 XA.XIR[8].XIC[11].icell.Ien VPWR 0.18829f
C1009 XA.XIR[15].XIC[1].icell.Ien Iout 0.07192f
C1010 XA.Cn[10] XA.XIR[7].XIC[10].icell.Ien 0.04604f
C1011 XThR.XTB7.Y XThR.Tn[14] 0.4222f
C1012 XA.XIR[5].XIC_dummy_left.icell.Iout Iout 0.03553f
C1013 XA.XIR[3].XIC[0].icell.PDM Vbias 0.03915f
C1014 XA.Cn[9] XA.XIR[12].XIC[9].icell.Ien 0.04604f
C1015 XA.Cn[1] VPWR 3.60376f
C1016 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.PDM 0.02104f
C1017 XA.XIR[8].XIC[2].icell.PDM Vbias 0.03928f
C1018 XA.Cn[11] XA.XIR[14].XIC[11].icell.Ien 0.04604f
C1019 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.Ien 0.04854f
C1020 XA.XIR[2].XIC[6].icell.PDM Vbias 0.03928f
C1021 XA.XIR[13].XIC[3].icell.Ien Vbias 0.19161f
C1022 XThR.XTB4.Y XThR.XTBN.A 0.03415f
C1023 XA.Cn[4] XA.XIR[15].XIC[4].icell.PDM 0.02601f
C1024 a_n997_3755# VPWR 0.0133f
C1025 XThR.XTB2.Y VPWR 0.98845f
C1026 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PDM 0.04035f
C1027 XA.Cn[14] XA.XIR[0].XIC[14].icell.PDM 0.02792f
C1028 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout 0.06446f
C1029 XA.XIR[15].XIC[12].icell.Ien VPWR 0.31713f
C1030 XA.XIR[0].XIC[13].icell.Ien VPWR 0.18776f
C1031 XThR.XTB5.Y XThR.Tn[5] 0.01094f
C1032 XA.XIR[11].XIC[6].icell.Ien Vbias 0.19161f
C1033 XA.Cn[11] XThR.Tn[2] 0.40741f
C1034 XThR.XTBN.A XThR.Tn[10] 0.12147f
C1035 XThR.Tn[1] XA.XIR[1].XIC[2].icell.Ien 0.14211f
C1036 XThR.Tn[14] XA.XIR[14].XIC[2].icell.Ien 0.14211f
C1037 XA.XIR[15].XIC[6].icell.Ien Iout 0.07192f
C1038 XA.XIR[12].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1039 thermo15c_0.XTB7.B thermo15c_0.XTB6.Y 0.30244f
C1040 XA.XIR[10].XIC[8].icell.Ien Vbias 0.19161f
C1041 thermo15c_0.XTB5.Y thermo15c_0.XTB7.Y 0.036f
C1042 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PDM 0.04035f
C1043 XA.Cn[2] XA.XIR[6].XIC[2].icell.PDM 0.02601f
C1044 XA.XIR[4].XIC[9].icell.Ien Iout 0.06801f
C1045 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1046 XA.Cn[12] XA.XIR[13].XIC[12].icell.PDM 0.02601f
C1047 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.PDM 0.02104f
C1048 XA.Cn[5] XA.XIR[2].XIC[5].icell.PDM 0.02602f
C1049 XA.Cn[3] XA.XIR[6].XIC[3].icell.Ien 0.04604f
C1050 XThR.Tn[13] XA.XIR[13].XIC[6].icell.Ien 0.14211f
C1051 XA.XIR[0].XIC[0].icell.Ien Iout 0.06743f
C1052 a_n1049_5611# VPWR 0.71817f
C1053 thermo15c_0.XTB3.Y XA.Cn[3] 0.01335f
C1054 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.Ien 0.04854f
C1055 thermo15c_0.XTB2.Y thermo15c_0.XTB3.Y 2.04808f
C1056 thermo15c_0.XTB6.A thermo15c_0.XTB7.A 0.44014f
C1057 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.Ien 0.04854f
C1058 thermo15c_0.XTB1.Y thermo15c_0.XTB4.Y 0.05121f
C1059 XA.XIR[14].XIC[1].icell.Ien VPWR 0.18883f
C1060 XA.XIR[8].XIC[3].icell.Ien Iout 0.06801f
C1061 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.Ien 0.04854f
C1062 XA.XIR[2].XIC[10].icell.Ien Vbias 0.19161f
C1063 XA.XIR[10].XIC[2].icell.PDM VPWR 0.01171f
C1064 XA.Cn[0] Vbias 0.27573f
C1065 XA.XIR[1].XIC[12].icell.Ien Vbias 0.19173f
C1066 XA.Cn[12] XThR.Tn[6] 0.40738f
C1067 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.PDM 0.02104f
C1068 XThR.XTBN.Y XThR.Tn[4] 0.6035f
C1069 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.PDM 0.02104f
C1070 XA.XIR[9].XIC[12].icell.Ien Iout 0.06801f
C1071 XA.XIR[6].XIC[3].icell.Ien VPWR 0.18829f
C1072 thermo15c_0.XTB3.Y VPWR 1.07064f
C1073 XThR.XTBN.Y a_n1049_7493# 0.08456f
C1074 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.Ien 0.04854f
C1075 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.PDM 0.02104f
C1076 XA.XIR[0].XIC[5].icell.Ien Iout 0.0675f
C1077 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.PDM 0.02104f
C1078 XThR.Tn[9] XA.XIR[9].XIC_dummy_left.icell.Iout 0.03386f
C1079 XThR.XTBN.Y XThR.XTB6.Y 0.1894f
C1080 XThR.Tn[6] XA.XIR[6].XIC[11].icell.Ien 0.14211f
C1081 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.PDM 0.02104f
C1082 XA.XIR[7].XIC[6].icell.PDM Vbias 0.03928f
C1083 XA.XIR[7].XIC[8].icell.Ien Iout 0.06801f
C1084 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.PDM 0.02104f
C1085 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout 0.06446f
C1086 XA.XIR[15].XIC[4].icell.PDM Vbias 0.03928f
C1087 XA.XIR[6].XIC[13].icell.PDM Vbias 0.03928f
C1088 XA.XIR[7].XIC_dummy_left.icell.Iout VPWR 0.10954f
C1089 XA.XIR[2].XIC[1].icell.Ien VPWR 0.18829f
C1090 XThR.XTB3.Y XThR.Tn[3] 0.01287f
C1091 XA.Cn[13] XThR.Tn[1] 0.40745f
C1092 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.Ien 0.04854f
C1093 XA.XIR[0].XIC[10].icell.PDM VPWR 0.01132f
C1094 XA.XIR[11].XIC[2].icell.Ien VPWR 0.18829f
C1095 XA.XIR[15].XIC[10].icell.Ien VPWR 0.31713f
C1096 XA.XIR[14].XIC[10].icell.PDM Vbias 0.03928f
C1097 XA.XIR[10].XIC[4].icell.Ien VPWR 0.18829f
C1098 XA.Cn[5] XThR.Tn[7] 0.40738f
C1099 XA.Cn[10] XA.XIR[8].XIC[10].icell.Ien 0.04604f
C1100 XA.Cn[13] XThR.Tn[12] 0.40739f
C1101 XThR.XTBN.A a_n997_1803# 0.09118f
C1102 XA.XIR[9].XIC[2].icell.PDM Vbias 0.03928f
C1103 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PDM 0.04035f
C1104 XThR.XTB4.Y XThR.XTB6.Y 0.04273f
C1105 XThR.XTB3.Y XThR.XTB7.Y 0.03772f
C1106 XA.Cn[11] XA.XIR[1].XIC[11].icell.Ien 0.04606f
C1107 XA.Cn[5] XA.XIR[7].XIC[5].icell.PDM 0.02601f
C1108 thermo15c_0.XTB4.Y a_8963_9569# 0.07199f
C1109 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PDM 0.04035f
C1110 XA.XIR[3].XIC[13].icell.Ien VPWR 0.18829f
C1111 XA.XIR[12].XIC[13].icell.Ien Vbias 0.19161f
C1112 XA.XIR[10].XIC[0].icell.Ien Iout 0.06795f
C1113 XThR.XTB6.Y XThR.Tn[10] 0.02461f
C1114 XA.Cn[8] XA.XIR[2].XIC[8].icell.PDM 0.02602f
C1115 XA.Cn[12] XThR.Tn[4] 0.40738f
C1116 XA.XIR[2].XIC[6].icell.Ien VPWR 0.18829f
C1117 a_n997_715# VPWR 0.02818f
C1118 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.PDM 0.02104f
C1119 XA.XIR[1].XIC[8].icell.Ien VPWR 0.18829f
C1120 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1121 XA.XIR[1].XIC[7].icell.PDM Vbias 0.03928f
C1122 XThR.Tn[8] XA.XIR[8].XIC[3].icell.Ien 0.14211f
C1123 XA.XIR[6].XIC[12].icell.Ien Vbias 0.19161f
C1124 XA.Cn[12] XA.XIR[11].XIC[12].icell.Ien 0.04604f
C1125 XThR.Tn[10] XA.XIR[10].XIC_dummy_left.icell.Iout 0.03385f
C1126 XA.Cn[11] XThR.Tn[10] 0.40738f
C1127 XA.XIR[4].XIC[7].icell.PDM Vbias 0.03928f
C1128 XA.Cn[14] XA.XIR[4].XIC[14].icell.Ien 0.04604f
C1129 XA.Cn[5] XA.XIR[9].XIC[5].icell.Ien 0.04604f
C1130 XA.XIR[3].XIC_15.icell.PDM Vbias 0.03927f
C1131 XA.XIR[14].XIC[6].icell.Ien Vbias 0.19161f
C1132 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.PDM 0.02104f
C1133 XThR.Tn[5] XA.XIR[5].XIC[2].icell.Ien 0.14211f
C1134 XA.XIR[13].XIC[8].icell.Ien Vbias 0.19161f
C1135 XA.Cn[3] XThR.Tn[3] 0.40738f
C1136 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.PDM 0.02104f
C1137 XA.Cn[11] XA.Cn[12] 0.12311f
C1138 a_2979_9615# XA.Cn[0] 0.27729f
C1139 XA.XIR[12].XIC_dummy_left.icell.Iout Iout 0.03553f
C1140 XA.XIR[3].XIC[5].icell.Ien Iout 0.06801f
C1141 XA.XIR[6].XIC[1].icell.PDM VPWR 0.01171f
C1142 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.Ien 0.04854f
C1143 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PDM 0.04035f
C1144 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.PDM 0.02104f
C1145 XThR.Tn[1] XA.XIR[1].XIC[7].icell.Ien 0.14211f
C1146 XThR.Tn[14] XA.XIR[14].XIC[7].icell.Ien 0.14211f
C1147 XA.Cn[4] XThR.Tn[5] 0.40738f
C1148 XA.XIR[5].XIC[8].icell.PDM VPWR 0.01171f
C1149 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.PDM 0.02104f
C1150 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.PDM 0.02104f
C1151 XA.Cn[1] XA.XIR[15].XIC[1].icell.Ien 0.04292f
C1152 XA.XIR[13].XIC[2].icell.PDM VPWR 0.01171f
C1153 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.PDM 0.02104f
C1154 thermo15c_0.XTB7.A a_4067_9615# 0.0127f
C1155 XA.XIR[4].XIC[14].icell.Ien Iout 0.06801f
C1156 XThR.Tn[3] VPWR 8.06517f
C1157 thermo15c_0.XTB6.Y XA.Cn[8] 0.02463f
C1158 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.PDM 0.02104f
C1159 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout 0.06446f
C1160 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.Ien 0.04854f
C1161 XA.XIR[12].XIC[7].icell.PDM VPWR 0.01171f
C1162 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.Ien 0.04854f
C1163 XA.Cn[0] XThR.Tn[0] 0.41303f
C1164 XA.XIR[12].XIC_dummy_right.icell.Iout XA.XIR[13].XIC_dummy_right.icell.Iout 0.04047f
C1165 XA.Cn[11] XA.XIR[6].XIC[11].icell.Ien 0.04604f
C1166 XA.XIR[8].XIC[8].icell.Ien Iout 0.06801f
C1167 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.Ien 0.04854f
C1168 thermo15c_0.XTBN.Y XA.Cn[11] 0.40412f
C1169 XThR.XTB7.Y VPWR 1.14768f
C1170 XA.Cn[3] XA.XIR[3].XIC[3].icell.PDM 0.02601f
C1171 XA.XIR[2].XIC_15.icell.Ien Vbias 0.19195f
C1172 XA.XIR[12].XIC[11].icell.Ien Vbias 0.19161f
C1173 XA.Cn[8] XA.XIR[7].XIC[8].icell.PDM 0.02601f
C1174 XThR.XTB5.A XThR.XTB5.Y 0.0538f
C1175 XA.XIR[8].XIC_dummy_left.icell.Iout VPWR 0.11f
C1176 XA.Cn[9] Iout 0.22393f
C1177 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.Ien 0.04854f
C1178 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.Ien 0.04854f
C1179 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PDM 0.04035f
C1180 XA.XIR[15].XIC_15.icell.Ien VPWR 0.37868f
C1181 thermo15c_0.XTB7.A XA.Cn[6] 0.10502f
C1182 XA.XIR[6].XIC[8].icell.Ien VPWR 0.18829f
C1183 XA.Cn[7] XThR.Tn[2] 0.40741f
C1184 XA.XIR[10].XIC[1].icell.PDM Vbias 0.03928f
C1185 XA.Cn[7] XA.XIR[11].XIC[7].icell.PDM 0.02601f
C1186 XA.XIR[0].XIC[10].icell.Ien Iout 0.0675f
C1187 thermo15c_0.XTB5.Y XA.Cn[9] 0.01732f
C1188 XA.Cn[9] XA.XIR[15].XIC[9].icell.Ien 0.04292f
C1189 XA.XIR[3].XIC[3].icell.PDM VPWR 0.01171f
C1190 XA.XIR[8].XIC[5].icell.PDM VPWR 0.01171f
C1191 XA.XIR[14].XIC[2].icell.Ien VPWR 0.18883f
C1192 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.Ien 0.04854f
C1193 thermo15c_0.XTB1.Y Vbias 0.01576f
C1194 XA.XIR[2].XIC[9].icell.PDM VPWR 0.01171f
C1195 XA.Cn[2] XA.XIR[2].XIC[2].icell.Ien 0.04605f
C1196 XA.XIR[13].XIC[4].icell.Ien VPWR 0.18829f
C1197 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.PDM 0.02104f
C1198 XA.XIR[7].XIC[13].icell.Ien Iout 0.06801f
C1199 XA.XIR[5].XIC[5].icell.Ien Vbias 0.19161f
C1200 XA.XIR[10].XIC_15.icell.PUM VPWR 0.01655f
C1201 XA.XIR[15].XIC_dummy_right.icell.Iout VPWR 0.21463f
C1202 XA.XIR[11].XIC[7].icell.Ien VPWR 0.18829f
C1203 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.Ien 0.04854f
C1204 XA.Cn[0] XA.XIR[1].XIC[0].icell.PDM 0.02602f
C1205 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PDM 0.04035f
C1206 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.PDM 0.02104f
C1207 XA.XIR[13].XIC[0].icell.Ien Iout 0.06795f
C1208 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.PDM 0.02104f
C1209 thermo15c_0.XTBN.Y a_4861_9615# 0.07601f
C1210 XA.XIR[10].XIC[9].icell.Ien VPWR 0.18829f
C1211 XThR.XTB6.Y XThR.Tn[13] 0.32265f
C1212 XA.Cn[0] XA.XIR[4].XIC[0].icell.PDM 0.02601f
C1213 XThR.Tn[5] Vbias 1.39526f
C1214 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.Ien 0.04854f
C1215 XA.XIR[0].XIC[9].icell.PDM Vbias 0.03945f
C1216 a_n997_2667# VPWR 0.01642f
C1217 bias[1] Vbias 0.05009f
C1218 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1219 XThR.XTB5.A XThR.XTB1.Y 0.1098f
C1220 XA.Cn[12] XA.XIR[14].XIC[12].icell.Ien 0.04604f
C1221 thermo15c_0.XTB3.Y thermo15c_0.XTB7.Y 0.03772f
C1222 thermo15c_0.XTB4.Y thermo15c_0.XTB6.Y 0.04273f
C1223 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PDM 0.04035f
C1224 XA.Cn[11] XThR.Tn[13] 0.40738f
C1225 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR 0.38522f
C1226 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PDM 0.04035f
C1227 XA.XIR[2].XIC[11].icell.Ien VPWR 0.18829f
C1228 XA.Cn[7] XA.XIR[10].XIC[7].icell.Ien 0.04604f
C1229 XA.Cn[14] XA.XIR[1].XIC[14].icell.PDM 0.02602f
C1230 XA.Cn[3] XThR.Tn[11] 0.40738f
C1231 XThR.XTB6.A data[4] 0.48493f
C1232 XA.Cn[14] XA.XIR[10].XIC[14].icell.PDM 0.02601f
C1233 XA.XIR[1].XIC[13].icell.Ien VPWR 0.18829f
C1234 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PDM 0.04035f
C1235 XThR.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.14211f
C1236 XA.Cn[14] XA.XIR[4].XIC[14].icell.PDM 0.02601f
C1237 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.Ien 0.04854f
C1238 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Iout 0.03777f
C1239 XA.Cn[8] XThR.Tn[9] 0.40738f
C1240 XA.Cn[9] XThR.Tn[8] 0.40738f
C1241 XA.XIR[12].XIC[0].icell.Ien VPWR 0.18829f
C1242 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.Ien 0.04854f
C1243 XA.Cn[13] XA.XIR[9].XIC[13].icell.Ien 0.04604f
C1244 XThR.Tn[11] VPWR 9.00382f
C1245 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PDM 0.04035f
C1246 XThR.Tn[5] XA.XIR[5].XIC[7].icell.Ien 0.14211f
C1247 XA.Cn[10] XA.XIR[11].XIC[10].icell.PDM 0.02601f
C1248 XA.Cn[4] XA.XIR[8].XIC[4].icell.PDM 0.02601f
C1249 XA.XIR[7].XIC[9].icell.PDM VPWR 0.01171f
C1250 XA.Cn[0] XA.XIR[1].XIC[0].icell.Ien 0.04606f
C1251 XA.XIR[3].XIC[10].icell.Ien Iout 0.06801f
C1252 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1253 XA.XIR[15].XIC[7].icell.PDM VPWR 0.01512f
C1254 XA.Cn[0] XA.XIR[4].XIC[0].icell.Ien 0.04604f
C1255 XA.Cn[0] XThR.Tn[1] 0.40748f
C1256 XThR.Tn[1] XA.XIR[1].XIC[12].icell.Ien 0.14211f
C1257 XA.XIR[2].XIC[3].icell.Ien Iout 0.06801f
C1258 XThR.XTB5.Y XThR.Tn[9] 0.01732f
C1259 XA.XIR[1].XIC[5].icell.Ien Iout 0.06801f
C1260 XA.Cn[0] XThR.Tn[12] 0.40738f
C1261 XA.XIR[6].XIC[0].icell.PDM Vbias 0.03915f
C1262 XA.XIR[9].XIC[5].icell.PDM VPWR 0.01171f
C1263 XA.Cn[7] XThR.Tn[10] 0.40738f
C1264 XA.XIR[15].XIC[13].icell.Ien Vbias 0.15966f
C1265 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.Ien 0.04854f
C1266 XA.XIR[5].XIC[7].icell.PDM Vbias 0.03928f
C1267 XA.XIR[8].XIC[13].icell.Ien Iout 0.06801f
C1268 thermo15c_0.XTB1.Y a_2979_9615# 0.21263f
C1269 thermo15c_0.XTBN.A data[3] 0.07741f
C1270 data[1] data[2] 0.01393f
C1271 XA.Cn[7] XA.XIR[14].XIC[7].icell.PDM 0.02601f
C1272 XA.XIR[13].XIC[1].icell.PDM Vbias 0.03928f
C1273 XThR.XTBN.A a_n997_3979# 0.02087f
C1274 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.PDM 0.02104f
C1275 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.Ien 0.04854f
C1276 XA.XIR[12].XIC[6].icell.PDM Vbias 0.03928f
C1277 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.Ien 0.04854f
C1278 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.04035f
C1279 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.PDM 0.02104f
C1280 XA.Cn[8] XA.XIR[4].XIC[8].icell.Ien 0.04604f
C1281 XA.XIR[1].XIC[10].icell.PDM VPWR 0.01171f
C1282 thermo15c_0.XTBN.A XA.Cn[11] 0.11997f
C1283 XA.XIR[6].XIC[13].icell.Ien VPWR 0.18829f
C1284 XA.XIR[10].XIC[14].icell.Ien VPWR 0.18835f
C1285 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1286 XA.XIR[0].XIC_15.icell.Ien Iout 0.06774f
C1287 XA.XIR[4].XIC[10].icell.PDM VPWR 0.01171f
C1288 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PDM 0.04035f
C1289 XA.XIR[13].XIC_15.icell.PUM VPWR 0.01655f
C1290 XA.XIR[14].XIC[7].icell.Ien VPWR 0.18883f
C1291 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1292 XA.XIR[6].XIC[0].icell.Ien Iout 0.06795f
C1293 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PDM 0.04035f
C1294 XA.Cn[5] XA.XIR[12].XIC[5].icell.PDM 0.02601f
C1295 XA.XIR[13].XIC[9].icell.Ien VPWR 0.18829f
C1296 XA.XIR[5].XIC[10].icell.Ien Vbias 0.19161f
C1297 XA.XIR[15].XIC_dummy_left.icell.Iout Iout 0.03553f
C1298 XA.Cn[10] XA.XIR[2].XIC[10].icell.Ien 0.04605f
C1299 thermo15c_0.XTBN.Y XA.Cn[7] 0.85979f
C1300 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.Ien 0.04854f
C1301 XA.XIR[3].XIC[2].icell.PDM Vbias 0.03928f
C1302 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1303 XA.XIR[8].XIC[4].icell.PDM Vbias 0.03928f
C1304 thermo15c_0.XTB2.Y data[1] 0.017f
C1305 XThR.Tn[13] XA.XIR[13].XIC_dummy_left.icell.Iout 0.03385f
C1306 XThR.Tn[12] XA.XIR[12].XIC[13].icell.Ien 0.14211f
C1307 XA.XIR[2].XIC[8].icell.PDM Vbias 0.03928f
C1308 XA.Cn[5] Iout 0.22432f
C1309 XA.Cn[13] XA.XIR[11].XIC[13].icell.Ien 0.04604f
C1310 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PDM 0.04035f
C1311 XThR.XTBN.A XThR.Tn[7] 0.01439f
C1312 XA.XIR[0].XIC_dummy_right.icell.Iout Iout 0.01732f
C1313 XA.XIR[12].XIC[5].icell.Ien Vbias 0.19161f
C1314 XA.Cn[7] XA.XIR[13].XIC[7].icell.Ien 0.04604f
C1315 XThR.XTBN.A a_n997_2891# 0.01719f
C1316 XA.Cn[3] XThR.Tn[14] 0.40738f
C1317 thermo15c_0.XTB5.Y XA.Cn[5] 0.01168f
C1318 XA.Cn[14] XA.XIR[13].XIC[14].icell.PDM 0.02601f
C1319 XA.XIR[6].XIC[5].icell.Ien Iout 0.06801f
C1320 VPWR data[1] 0.44103f
C1321 XThR.Tn[6] XThR.Tn[7] 0.11401f
C1322 XA.Cn[4] XA.XIR[9].XIC[4].icell.PDM 0.02601f
C1323 XA.XIR[15].XIC[11].icell.Ien Vbias 0.15966f
C1324 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PDM 0.04056f
C1325 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PDM 0.04035f
C1326 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.Ien 0.04854f
C1327 XA.XIR[5].XIC[1].icell.Ien VPWR 0.18829f
C1328 XThR.Tn[8] XA.XIR[8].XIC[13].icell.Ien 0.14211f
C1329 XThR.Tn[14] VPWR 9.25423f
C1330 XA.Cn[10] XA.XIR[14].XIC[10].icell.PDM 0.02601f
C1331 XA.XIR[11].XIC[0].icell.PDM VPWR 0.01171f
C1332 XA.XIR[10].XIC[4].icell.PDM VPWR 0.01171f
C1333 XA.XIR[10].XIC[12].icell.Ien VPWR 0.18829f
C1334 XThR.XTB2.Y a_n1335_8107# 0.01006f
C1335 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.Ien 0.04854f
C1336 XA.XIR[11].XIC[4].icell.Ien Iout 0.06801f
C1337 XA.Cn[0] XA.XIR[5].XIC[0].icell.PDM 0.02601f
C1338 XA.XIR[10].XIC[6].icell.Ien Iout 0.06801f
C1339 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.Ien 0.04854f
C1340 XThR.Tn[5] XA.XIR[5].XIC[12].icell.Ien 0.14211f
C1341 thermo15c_0.XTB6.Y Vbias 0.01779f
C1342 XA.XIR[5].XIC[6].icell.Ien VPWR 0.18829f
C1343 XA.Cn[7] XThR.Tn[13] 0.40738f
C1344 XA.XIR[3].XIC_15.icell.Ien Iout 0.0694f
C1345 XA.Cn[8] XA.XIR[12].XIC[8].icell.PDM 0.02601f
C1346 XA.XIR[2].XIC[8].icell.Ien Iout 0.06801f
C1347 XA.XIR[7].XIC[8].icell.PDM Vbias 0.03928f
C1348 XA.XIR[9].XIC[1].icell.Ien Vbias 0.19161f
C1349 XThR.Tn[12] XA.XIR[12].XIC[11].icell.Ien 0.14211f
C1350 XA.Cn[1] XA.XIR[0].XIC[1].icell.PDM 0.02803f
C1351 XA.XIR[1].XIC[10].icell.Ien Iout 0.06801f
C1352 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR 0.3367f
C1353 XA.XIR[6].XIC_15.icell.PDM Vbias 0.03927f
C1354 XA.XIR[4].XIC[3].icell.Ien Vbias 0.19161f
C1355 XA.XIR[15].XIC[6].icell.PDM Vbias 0.03928f
C1356 XThR.XTB2.Y a_n1049_7787# 0.2342f
C1357 XA.Cn[14] XA.XIR[5].XIC[14].icell.PDM 0.02601f
C1358 XA.XIR[2].XIC_dummy_left.icell.Iout VPWR 0.10954f
C1359 XA.Cn[4] XThR.Tn[9] 0.40738f
C1360 XA.XIR[0].XIC[12].icell.PDM VPWR 0.01451f
C1361 XA.Cn[5] XThR.Tn[8] 0.40738f
C1362 XA.XIR[13].XIC[14].icell.Ien VPWR 0.18835f
C1363 XThR.Tn[4] XA.XIR[4].XIC[2].icell.Ien 0.14211f
C1364 XA.XIR[9].XIC[4].icell.PDM Vbias 0.03928f
C1365 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.Ien 0.04854f
C1366 XA.XIR[3].XIC_dummy_right.icell.Iout Iout 0.01732f
C1367 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PDM 0.04035f
C1368 XThR.XTB6.Y XThR.Tn[7] 0.01462f
C1369 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PDM 0.04035f
C1370 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.Ien 0.04854f
C1371 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.PDM 0.02104f
C1372 XA.XIR[9].XIC[6].icell.Ien Vbias 0.19161f
C1373 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR 0.0824f
C1374 thermo15c_0.XTB5.A data[0] 0.14415f
C1375 XA.Cn[5] XA.XIR[15].XIC[5].icell.PDM 0.02601f
C1376 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.PDM 0.02104f
C1377 XA.Cn[11] XThR.Tn[7] 0.40738f
C1378 XA.XIR[10].XIC[10].icell.Ien VPWR 0.18829f
C1379 XA.XIR[1].XIC[9].icell.PDM Vbias 0.03928f
C1380 XA.Cn[13] XA.XIR[14].XIC[13].icell.Ien 0.04604f
C1381 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.PDM 0.02104f
C1382 XA.XIR[7].XIC[2].icell.Ien Vbias 0.19161f
C1383 XA.XIR[4].XIC[9].icell.PDM Vbias 0.03928f
C1384 XA.XIR[5].XIC_15.icell.Ien Vbias 0.19195f
C1385 XA.Cn[3] XA.XIR[6].XIC[3].icell.PDM 0.02601f
C1386 XA.Cn[6] XA.XIR[2].XIC[6].icell.PDM 0.02602f
C1387 XThR.Tn[3] XA.XIR[3].XIC[5].icell.Ien 0.14211f
C1388 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PDM 0.0404f
C1389 XA.XIR[12].XIC_15.icell.PDM Vbias 0.03927f
C1390 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.Ien 0.04854f
C1391 XThR.XTB3.Y VPWR 1.07975f
C1392 XA.Cn[6] XA.XIR[11].XIC[6].icell.Ien 0.04604f
C1393 thermo15c_0.XTBN.A XA.Cn[7] 0.01451f
C1394 XThR.XTB5.A XThR.XTB6.A 1.80461f
C1395 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1396 XA.XIR[6].XIC[3].icell.PDM VPWR 0.01171f
C1397 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PDM 0.0404f
C1398 XA.XIR[6].XIC[10].icell.Ien Iout 0.06801f
C1399 XA.XIR[14].XIC[0].icell.PDM VPWR 0.01171f
C1400 XA.Cn[2] XA.XIR[5].XIC[2].icell.Ien 0.04604f
C1401 XA.XIR[5].XIC[10].icell.PDM VPWR 0.01171f
C1402 XThR.Tn[9] Vbias 1.39532f
C1403 VPWR data[2] 0.21031f
C1404 XA.XIR[13].XIC[4].icell.PDM VPWR 0.01171f
C1405 XA.XIR[13].XIC[12].icell.Ien VPWR 0.18829f
C1406 thermo15c_0.XTB7.A a_5155_9615# 0.02287f
C1407 XA.XIR[14].XIC[4].icell.Ien Iout 0.06801f
C1408 XA.Cn[0] XA.XIR[2].XIC[0].icell.Ien 0.04605f
C1409 XA.Cn[9] XThR.Tn[3] 0.40738f
C1410 XA.XIR[12].XIC[9].icell.PDM VPWR 0.01171f
C1411 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.PDM 0.02104f
C1412 XA.XIR[13].XIC[6].icell.Ien Iout 0.06801f
C1413 XA.XIR[9].XIC[2].icell.Ien VPWR 0.18829f
C1414 XA.Cn[4] XA.XIR[0].XIC[4].icell.Ien 0.04658f
C1415 thermo15c_0.XTB1.Y thermo15c_0.XTB6.A 0.01609f
C1416 XA.Cn[10] XThR.Tn[5] 0.40738f
C1417 XA.XIR[15].XIC[0].icell.Ien Vbias 0.15953f
C1418 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.Ien 0.04854f
C1419 thermo15c_0.XTB5.A thermo15c_0.XTB7.A 0.07824f
C1420 XA.XIR[11].XIC[9].icell.Ien Iout 0.06801f
C1421 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PDM 0.04035f
C1422 XA.Cn[8] XA.XIR[15].XIC[8].icell.PDM 0.02601f
C1423 XA.XIR[10].XIC[3].icell.PDM Vbias 0.03928f
C1424 XA.XIR[5].XIC[11].icell.Ien VPWR 0.18829f
C1425 XA.Cn[3] VPWR 3.60513f
C1426 XThR.XTBN.A data[5] 0.0148f
C1427 thermo15c_0.XTB2.Y VPWR 0.97668f
C1428 XA.XIR[3].XIC[5].icell.PDM VPWR 0.01171f
C1429 XA.Cn[6] XA.XIR[7].XIC[6].icell.PDM 0.02601f
C1430 XA.XIR[8].XIC[7].icell.PDM VPWR 0.01171f
C1431 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.PDM 0.02104f
C1432 XA.XIR[2].XIC[11].icell.PDM VPWR 0.01171f
C1433 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PDM 0.04035f
C1434 XA.XIR[2].XIC[13].icell.Ien Iout 0.06801f
C1435 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.PDM 0.02104f
C1436 XA.XIR[15].XIC[5].icell.Ien Vbias 0.15966f
C1437 XA.Cn[9] XA.XIR[2].XIC[9].icell.PDM 0.02602f
C1438 XA.XIR[12].XIC[6].icell.Ien VPWR 0.18829f
C1439 XA.XIR[1].XIC_15.icell.Ien Iout 0.0694f
C1440 XA.XIR[4].XIC[8].icell.Ien Vbias 0.19161f
C1441 XA.Cn[13] XThR.Tn[2] 0.40742f
C1442 XA.XIR[10].XIC_15.icell.Ien VPWR 0.26829f
C1443 XThR.XTB6.Y a_n997_1579# 0.07626f
C1444 XA.XIR[8].XIC[2].icell.Ien Vbias 0.19161f
C1445 thermo15c_0.XTBN.Y a_5949_9615# 0.07703f
C1446 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.PDM 0.02104f
C1447 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.PDM 0.02104f
C1448 XThR.Tn[4] XA.XIR[4].XIC[7].icell.Ien 0.14211f
C1449 XA.Cn[9] XA.XIR[10].XIC[9].icell.Ien 0.04604f
C1450 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.Ien 0.04854f
C1451 XA.XIR[0].XIC[11].icell.PDM Vbias 0.03945f
C1452 XA.XIR[13].XIC[10].icell.Ien VPWR 0.18829f
C1453 thermo15c_0.XTB7.B XA.Cn[8] 0.05151f
C1454 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PDM 0.04035f
C1455 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PDM 0.04035f
C1456 XA.XIR[9].XIC[11].icell.Ien Vbias 0.19161f
C1457 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Iout 0.02485f
C1458 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.PDM 0.02104f
C1459 thermo15c_0.XTB7.A thermo15c_0.XTBN.Y 0.59539f
C1460 XA.XIR[5].XIC[3].icell.Ien Iout 0.06801f
C1461 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PDM 0.04035f
C1462 XA.XIR[12].XIC[14].icell.PDM Vbias 0.03928f
C1463 XA.Cn[2] Vbias 0.83223f
C1464 XA.Cn[14] XThR.Tn[6] 0.40742f
C1465 XA.Cn[14] XA.XIR[11].XIC[14].icell.Ien 0.04604f
C1466 XA.XIR[0].XIC[4].icell.Ien Vbias 0.19213f
C1467 XA.XIR[1].XIC_dummy_right.icell.Iout Iout 0.01732f
C1468 a_3773_9615# XA.Cn[1] 0.26251f
C1469 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.PDM 0.02104f
C1470 XA.XIR[10].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1471 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PDM 0.0404f
C1472 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.Ien 0.04854f
C1473 XA.XIR[15].XIC_15.icell.PDM Vbias 0.03927f
C1474 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PDM 0.04056f
C1475 XA.Cn[6] XA.XIR[14].XIC[6].icell.Ien 0.04604f
C1476 XA.Cn[12] XA.XIR[11].XIC[12].icell.PDM 0.02601f
C1477 XThR.Tn[12] XA.XIR[12].XIC[5].icell.Ien 0.14211f
C1478 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1479 XA.XIR[7].XIC[7].icell.Ien Vbias 0.19161f
C1480 XA.Cn[4] XA.XIR[3].XIC[4].icell.Ien 0.04604f
C1481 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.PDM 0.02104f
C1482 XThR.Tn[3] XA.XIR[3].XIC[10].icell.Ien 0.14211f
C1483 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.PDM 0.02104f
C1484 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.Ien 0.04854f
C1485 a_10051_9569# Vbias 0.0105f
C1486 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PDM 0.04056f
C1487 XA.Cn[9] XThR.Tn[11] 0.40738f
C1488 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.Ien 0.04854f
C1489 XA.Cn[4] XA.XIR[3].XIC[4].icell.PDM 0.02601f
C1490 XThR.XTB7.Y a_n1319_5317# 0.01283f
C1491 XA.XIR[7].XIC[11].icell.PDM VPWR 0.01171f
C1492 XThR.Tn[2] XA.XIR[2].XIC[5].icell.Ien 0.14211f
C1493 XA.Cn[9] XA.XIR[7].XIC[9].icell.PDM 0.02601f
C1494 XThR.Tn[6] Iout 1.12758f
C1495 XA.XIR[11].XIC[14].icell.Ien Iout 0.06801f
C1496 XA.XIR[15].XIC[9].icell.PDM VPWR 0.01512f
C1497 XA.XIR[4].XIC[4].icell.Ien VPWR 0.18829f
C1498 XA.XIR[6].XIC_15.icell.Ien Iout 0.0694f
C1499 XA.Cn[7] XThR.Tn[7] 0.40738f
C1500 XA.Cn[10] XA.XIR[5].XIC[10].icell.Ien 0.04604f
C1501 XA.XIR[6].XIC[2].icell.PDM Vbias 0.03928f
C1502 XA.XIR[14].XIC[9].icell.Ien Iout 0.06801f
C1503 XA.XIR[9].XIC[7].icell.PDM VPWR 0.01171f
C1504 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.Ien 0.04854f
C1505 XA.XIR[5].XIC[9].icell.PDM Vbias 0.03928f
C1506 thermo15c_0.XTB7.Y a_10915_9569# 0.06874f
C1507 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.Ien 0.04854f
C1508 XA.Cn[3] XA.XIR[7].XIC[3].icell.Ien 0.04604f
C1509 XA.XIR[9].XIC[7].icell.Ien VPWR 0.18829f
C1510 XA.Cn[2] XA.XIR[12].XIC[2].icell.Ien 0.04604f
C1511 XA.Cn[14] XThR.Tn[4] 0.40742f
C1512 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.Ien 0.04854f
C1513 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.PDM 0.02104f
C1514 thermo15c_0.XTBN.A data[0] 0.02545f
C1515 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.PDM 0.02104f
C1516 XA.XIR[13].XIC[3].icell.PDM Vbias 0.03928f
C1517 thermo15c_0.XTB4.Y thermo15c_0.XTB7.B 0.33064f
C1518 XThR.Tn[9] XA.XIR[9].XIC[3].icell.Ien 0.14211f
C1519 XA.Cn[12] XA.XIR[0].XIC[12].icell.Ien 0.04662f
C1520 XA.XIR[12].XIC[8].icell.PDM Vbias 0.03928f
C1521 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.PDM 0.02104f
C1522 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PDM 0.04035f
C1523 XA.Cn[1] XA.XIR[1].XIC[1].icell.PDM 0.02602f
C1524 XA.XIR[6].XIC_dummy_right.icell.Iout Iout 0.01732f
C1525 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.Ien 0.04854f
C1526 XA.XIR[1].XIC[12].icell.PDM VPWR 0.01171f
C1527 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.PDM 0.02104f
C1528 XA.Cn[13] XThR.Tn[10] 0.40739f
C1529 XA.Cn[1] XA.XIR[4].XIC[1].icell.PDM 0.02601f
C1530 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.Ien 0.04854f
C1531 XA.XIR[4].XIC[12].icell.PDM VPWR 0.01171f
C1532 XA.XIR[7].XIC[3].icell.Ien VPWR 0.18829f
C1533 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PDM 0.04035f
C1534 Vbias bias[0] 0.21039f
C1535 bias[1] bias[2] 0.16429f
C1536 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.Ien 0.04854f
C1537 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.Ien 0.04854f
C1538 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.PDM 0.02104f
C1539 XA.XIR[10].XIC[13].icell.Ien Vbias 0.19161f
C1540 XA.XIR[13].XIC_15.icell.Ien VPWR 0.26829f
C1541 XA.XIR[3].XIC[4].icell.Ien Vbias 0.19161f
C1542 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.Ien 0.04854f
C1543 XA.Cn[5] XThR.Tn[3] 0.40738f
C1544 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.Ien 0.04854f
C1545 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PDM 0.04035f
C1546 XA.Cn[9] XA.XIR[13].XIC[9].icell.Ien 0.04604f
C1547 XThR.Tn[4] Iout 1.12761f
C1548 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PDM 0.04035f
C1549 XA.Cn[12] XA.Cn[13] 0.17915f
C1550 XA.XIR[12].XIC[13].icell.PDM Vbias 0.03928f
C1551 XA.XIR[4].XIC[13].icell.Ien Vbias 0.19161f
C1552 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.PDM 0.02104f
C1553 XA.XIR[8].XIC[6].icell.PDM Vbias 0.03928f
C1554 XA.XIR[3].XIC[4].icell.PDM Vbias 0.03928f
C1555 XThR.Tn[7] XA.XIR[7].XIC[0].icell.Ien 0.14211f
C1556 XThR.XTBN.A XThR.Tn[8] 0.1369f
C1557 XA.Cn[6] XThR.Tn[5] 0.40738f
C1558 XA.XIR[2].XIC[10].icell.PDM Vbias 0.03928f
C1559 XA.XIR[11].XIC[12].icell.Ien Iout 0.06801f
C1560 XA.XIR[8].XIC[7].icell.Ien Vbias 0.19161f
C1561 XA.XIR[15].XIC[14].icell.PDM Vbias 0.03928f
C1562 thermo15c_0.XTB6.Y XA.Cn[10] 0.02478f
C1563 XA.Cn[14] XA.XIR[14].XIC[14].icell.Ien 0.04604f
C1564 XThR.Tn[4] XA.XIR[4].XIC[12].icell.Ien 0.14211f
C1565 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PDM 0.04035f
C1566 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.0404f
C1567 XA.Cn[2] XThR.Tn[0] 0.40765f
C1568 XA.XIR[0].XIC_15.icell.PUM VPWR 0.01577f
C1569 XThR.Tn[0] XA.XIR[0].XIC[4].icell.Ien 0.14211f
C1570 XA.XIR[13].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1571 XThR.Tn[10] XA.XIR[10].XIC[3].icell.Ien 0.14211f
C1572 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PDM 0.0404f
C1573 thermo15c_0.XTBN.Y XA.Cn[13] 0.41509f
C1574 XA.XIR[5].XIC[8].icell.Ien Iout 0.06801f
C1575 XA.Cn[5] XA.XIR[8].XIC[5].icell.PDM 0.02601f
C1576 XA.Cn[12] XA.XIR[14].XIC[12].icell.PDM 0.02601f
C1577 XA.XIR[10].XIC_dummy_left.icell.Iout Iout 0.03553f
C1578 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PDM 0.04035f
C1579 XA.Cn[11] Iout 0.22485f
C1580 XThR.XTB7.A data[4] 0.8689f
C1581 XA.XIR[0].XIC[9].icell.Ien Vbias 0.19213f
C1582 XThR.Tn[7] XA.XIR[7].XIC[5].icell.Ien 0.14211f
C1583 XA.XIR[15].XIC[1].icell.Ien VPWR 0.31713f
C1584 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.PDM 0.02104f
C1585 thermo15c_0.XTB2.Y thermo15c_0.XTB7.Y 0.0437f
C1586 thermo15c_0.XTB6.A thermo15c_0.XTB6.Y 0.10153f
C1587 XA.XIR[5].XIC_dummy_left.icell.Iout VPWR 0.11011f
C1588 thermo15c_0.XTB7.A thermo15c_0.XTBN.A 0.197f
C1589 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.Ien 0.04854f
C1590 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.Ien 0.04854f
C1591 XA.XIR[11].XIC[2].icell.PDM VPWR 0.01171f
C1592 XA.Cn[9] XThR.Tn[14] 0.40738f
C1593 thermo15c_0.XTB5.Y XA.Cn[11] 0.02112f
C1594 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.Ien 0.04854f
C1595 XA.XIR[12].XIC[3].icell.Ien Iout 0.06801f
C1596 XA.XIR[7].XIC[12].icell.Ien Vbias 0.19161f
C1597 XA.XIR[10].XIC[6].icell.PDM VPWR 0.01171f
C1598 XA.XIR[14].XIC[14].icell.Ien Iout 0.06801f
C1599 XThR.Tn[3] XA.XIR[3].XIC_15.icell.Ien 0.13564f
C1600 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.PDM 0.02104f
C1601 XA.Cn[12] XA.XIR[3].XIC[12].icell.Ien 0.04604f
C1602 thermo15c_0.XTB7.Y VPWR 1.07721f
C1603 XA.Cn[3] XA.XIR[8].XIC[3].icell.Ien 0.04604f
C1604 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout 0.06446f
C1605 XA.XIR[10].XIC[11].icell.Ien Vbias 0.19161f
C1606 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.Ien 0.04854f
C1607 XA.XIR[15].XIC[6].icell.Ien VPWR 0.31713f
C1608 XA.Cn[4] XA.XIR[1].XIC[4].icell.Ien 0.04607f
C1609 XA.XIR[3].XIC[1].icell.Ien Vbias 0.19161f
C1610 XThR.Tn[2] XA.XIR[2].XIC[10].icell.Ien 0.14211f
C1611 XA.XIR[4].XIC[9].icell.Ien VPWR 0.18829f
C1612 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.PDM 0.02104f
C1613 XA.Cn[0] XThR.Tn[2] 0.40744f
C1614 XA.XIR[0].XIC[0].icell.Ien VPWR 0.18776f
C1615 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.PDM 0.02104f
C1616 XA.XIR[7].XIC[10].icell.PDM Vbias 0.03928f
C1617 XA.XIR[8].XIC[3].icell.Ien VPWR 0.18829f
C1618 XA.XIR[11].XIC[10].icell.Ien Iout 0.06801f
C1619 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.Ien 0.04854f
C1620 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.Ien 0.04854f
C1621 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.PDM 0.02104f
C1622 XA.XIR[15].XIC[8].icell.PDM Vbias 0.03928f
C1623 XA.XIR[0].XIC[14].icell.PDM VPWR 0.01141f
C1624 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.Ien 0.04854f
C1625 XA.Cn[7] XA.XIR[4].XIC[7].icell.Ien 0.04604f
C1626 XA.Cn[6] XA.XIR[12].XIC[6].icell.PDM 0.02601f
C1627 XA.Cn[13] XThR.Tn[13] 0.40739f
C1628 XA.XIR[9].XIC[12].icell.Ien VPWR 0.18829f
C1629 XThR.XTB6.Y XThR.Tn[8] 0.02461f
C1630 XA.Cn[11] XA.XIR[7].XIC[11].icell.Ien 0.04604f
C1631 XA.Cn[5] XThR.Tn[11] 0.40738f
C1632 thermo15c_0.XTBN.Y a_7875_9569# 0.229f
C1633 XThR.Tn[9] XA.XIR[9].XIC[8].icell.Ien 0.14211f
C1634 XA.XIR[9].XIC[6].icell.PDM Vbias 0.03928f
C1635 XA.XIR[0].XIC[5].icell.Ien VPWR 0.18797f
C1636 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.04035f
C1637 XA.Cn[1] XThR.Tn[6] 0.40738f
C1638 XA.XIR[13].XIC[13].icell.Ien Vbias 0.19161f
C1639 XThR.XTBN.A a_n997_3755# 0.01939f
C1640 XA.XIR[11].XIC[0].icell.Ien Iout 0.06795f
C1641 thermo15c_0.XTB4.Y XA.Cn[8] 0.01307f
C1642 XThR.XTB2.Y XThR.XTBN.A 0.04716f
C1643 XA.XIR[3].XIC_15.icell.PUM VPWR 0.01655f
C1644 XA.XIR[12].XIC[12].icell.PDM Vbias 0.03928f
C1645 XA.Cn[8] XA.XIR[8].XIC[8].icell.PDM 0.02601f
C1646 XA.Cn[10] XThR.Tn[9] 0.40738f
C1647 XThR.XTB7.A XThR.Tn[5] 0.02751f
C1648 XA.Cn[11] XThR.Tn[8] 0.40738f
C1649 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.Ien 0.04854f
C1650 XA.XIR[7].XIC[8].icell.Ien VPWR 0.18829f
C1651 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1652 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.Ien 0.04854f
C1653 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.PDM 0.02104f
C1654 XA.XIR[15].XIC[13].icell.PDM Vbias 0.03928f
C1655 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PDM 0.04035f
C1656 XA.XIR[3].XIC[9].icell.Ien Vbias 0.19161f
C1657 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PDM 0.0404f
C1658 XA.XIR[1].XIC[11].icell.PDM Vbias 0.03928f
C1659 XA.XIR[14].XIC[12].icell.Ien Iout 0.06801f
C1660 XA.Cn[5] XA.XIR[9].XIC[5].icell.PDM 0.02601f
C1661 XA.Cn[8] XA.XIR[11].XIC[8].icell.Ien 0.04604f
C1662 XA.XIR[2].XIC[2].icell.Ien Vbias 0.19161f
C1663 XA.XIR[4].XIC[11].icell.PDM Vbias 0.03928f
C1664 XA.Cn[4] XA.XIR[6].XIC[4].icell.Ien 0.04604f
C1665 thermo15c_0.XTB7.B Vbias 0.12116f
C1666 XA.XIR[1].XIC[4].icell.Ien Vbias 0.19173f
C1667 XA.Cn[2] XThR.Tn[1] 0.40744f
C1668 XThR.XTB7.B data[4] 0.01382f
C1669 XA.XIR[9].XIC[4].icell.Ien Iout 0.06801f
C1670 a_n1049_8581# VPWR 0.71708f
C1671 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.PDM 0.02104f
C1672 XThR.Tn[11] XA.XIR[11].XIC[4].icell.Ien 0.14211f
C1673 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PDM 0.04035f
C1674 XA.XIR[8].XIC[12].icell.Ien Vbias 0.19161f
C1675 XA.XIR[13].XIC_dummy_left.icell.Iout Iout 0.03553f
C1676 XA.XIR[10].XIC[0].icell.Ien VPWR 0.18829f
C1677 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout 0.06446f
C1678 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.PDM 0.02104f
C1679 XA.Cn[2] XThR.Tn[12] 0.40738f
C1680 XThR.XTB1.Y XThR.XTB5.Y 0.05054f
C1681 XThR.Tn[0] XA.XIR[0].XIC[9].icell.Ien 0.14211f
C1682 XA.XIR[6].XIC[5].icell.PDM VPWR 0.01171f
C1683 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.Ien 0.04854f
C1684 XThR.Tn[10] XA.XIR[10].XIC[8].icell.Ien 0.14211f
C1685 XA.Cn[1] XA.XIR[5].XIC[1].icell.PDM 0.02601f
C1686 XA.XIR[14].XIC[2].icell.PDM VPWR 0.01171f
C1687 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.PDM 0.02104f
C1688 XA.Cn[2] XA.XIR[15].XIC[2].icell.Ien 0.04292f
C1689 XThR.Tn[6] XA.XIR[6].XIC[3].icell.Ien 0.14211f
C1690 XA.XIR[5].XIC[12].icell.PDM VPWR 0.01171f
C1691 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.PDM 0.02104f
C1692 XA.XIR[5].XIC[13].icell.Ien Iout 0.06801f
C1693 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.PDM 0.02104f
C1694 XA.Cn[1] XThR.Tn[4] 0.40738f
C1695 XA.XIR[13].XIC[6].icell.PDM VPWR 0.01171f
C1696 thermo15c_0.XTB7.A a_6243_9615# 0.02018f
C1697 XThR.Tn[7] XA.XIR[7].XIC[10].icell.Ien 0.14211f
C1698 XA.XIR[0].XIC[14].icell.Ien Vbias 0.19213f
C1699 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.Ien 0.04854f
C1700 XA.Cn[9] XA.XIR[12].XIC[9].icell.PDM 0.02601f
C1701 XA.XIR[13].XIC[11].icell.Ien Vbias 0.19161f
C1702 XA.XIR[12].XIC_dummy_left.icell.Ien XThR.Tn[12] 0.01244f
C1703 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.PDM 0.02104f
C1704 XA.XIR[11].XIC_15.icell.Ien Iout 0.0694f
C1705 XA.Cn[0] XThR.Tn[10] 0.40734f
C1706 XThR.XTB2.Y a_n1049_7493# 0.02133f
C1707 XA.XIR[12].XIC[8].icell.Ien Iout 0.06801f
C1708 VPWR data[7] 0.212f
C1709 XA.Cn[2] XA.XIR[0].XIC[2].icell.PDM 0.02803f
C1710 thermo15c_0.XTB6.Y XA.Cn[6] 0.01038f
C1711 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Iout 0.01728f
C1712 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.PDM 0.02104f
C1713 XA.XIR[12].XIC_dummy_left.icell.Iout VPWR 0.10997f
C1714 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.04035f
C1715 XA.XIR[3].XIC[5].icell.Ien VPWR 0.18829f
C1716 XA.XIR[11].XIC[1].icell.PDM Vbias 0.03928f
C1717 XThR.XTB2.Y XThR.XTB6.Y 0.04959f
C1718 XA.Cn[11] XA.XIR[8].XIC[11].icell.Ien 0.04604f
C1719 XA.XIR[14].XIC[10].icell.Ien Iout 0.06801f
C1720 XA.XIR[10].XIC[5].icell.PDM Vbias 0.03928f
C1721 XThR.Tn[2] XA.XIR[2].XIC_15.icell.Ien 0.13564f
C1722 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.PDM 0.02104f
C1723 XA.Cn[12] XA.XIR[1].XIC[12].icell.Ien 0.04606f
C1724 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Iout 0.0203f
C1725 XA.XIR[4].XIC[14].icell.Ien VPWR 0.18835f
C1726 XA.XIR[3].XIC[7].icell.PDM VPWR 0.01171f
C1727 thermo15c_0.XTB2.Y XA.Cn[9] 0.292f
C1728 XA.XIR[8].XIC[9].icell.PDM VPWR 0.01171f
C1729 XA.Cn[8] XA.XIR[9].XIC[8].icell.PDM 0.02601f
C1730 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.Ien 0.04854f
C1731 XA.Cn[7] Iout 0.22453f
C1732 XA.XIR[6].XIC[4].icell.Ien Vbias 0.19161f
C1733 XA.Cn[6] XA.XIR[15].XIC[6].icell.PDM 0.02601f
C1734 XA.XIR[2].XIC[13].icell.PDM VPWR 0.01171f
C1735 XA.XIR[11].XIC_dummy_right.icell.Iout Iout 0.01732f
C1736 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PDM 0.04035f
C1737 XA.XIR[8].XIC[8].icell.Ien VPWR 0.18829f
C1738 XA.XIR[12].XIC[11].icell.PDM Vbias 0.03928f
C1739 XA.Cn[5] XThR.Tn[14] 0.40738f
C1740 XThR.XTB6.Y a_n1049_5611# 0.26831f
C1741 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.Ien 0.04854f
C1742 XA.XIR[10].XIC_15.icell.PDM VPWR 0.07527f
C1743 XA.XIR[4].XIC[1].icell.Ien Iout 0.06801f
C1744 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.Ien 0.04854f
C1745 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.PDM 0.02104f
C1746 XA.XIR[15].XIC[12].icell.PDM Vbias 0.03928f
C1747 XA.Cn[9] VPWR 4.54443f
C1748 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR 0.39107f
C1749 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PDM 0.04035f
C1750 thermo15c_0.XTBN.Y XA.Cn[0] 0.45269f
C1751 XA.Cn[4] XA.XIR[6].XIC[4].icell.PDM 0.02601f
C1752 XA.Cn[7] XA.XIR[2].XIC[7].icell.PDM 0.02602f
C1753 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1754 XA.Cn[6] XA.XIR[9].XIC[6].icell.Ien 0.04604f
C1755 XThR.Tn[9] XA.XIR[9].XIC[13].icell.Ien 0.14211f
C1756 XA.XIR[0].XIC[10].icell.Ien VPWR 0.18776f
C1757 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.Ien 0.04854f
C1758 XA.XIR[0].XIC[13].icell.PDM Vbias 0.03945f
C1759 XA.XIR[11].XIC[3].icell.Ien Vbias 0.19161f
C1760 thermo15c_0.XTB6.Y a_5949_10571# 0.01283f
C1761 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PDM 0.04035f
C1762 XA.XIR[15].XIC[3].icell.Ien Iout 0.07192f
C1763 XA.Cn[8] XA.XIR[14].XIC[8].icell.Ien 0.04604f
C1764 XA.XIR[10].XIC[5].icell.Ien Vbias 0.19161f
C1765 thermo15c_0.XTBN.A a_7875_9569# 0.01939f
C1766 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PDM 0.04035f
C1767 XA.Cn[14] XA.XIR[11].XIC[14].icell.PDM 0.02601f
C1768 XA.XIR[4].XIC[6].icell.Ien Iout 0.06801f
C1769 XA.XIR[7].XIC[13].icell.Ien VPWR 0.18829f
C1770 XThR.Tn[13] XA.XIR[13].XIC[3].icell.Ien 0.14211f
C1771 XA.XIR[3].XIC[14].icell.Ien Vbias 0.19161f
C1772 XA.XIR[1].XIC_15.icell.PUM VPWR 0.01655f
C1773 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.Ien 0.04854f
C1774 XA.XIR[2].XIC[7].icell.Ien Vbias 0.19161f
C1775 XA.XIR[13].XIC[0].icell.Ien VPWR 0.18829f
C1776 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.Ien 0.04854f
C1777 XA.XIR[7].XIC[0].icell.Ien Iout 0.06795f
C1778 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.Ien 0.04854f
C1779 XA.XIR[1].XIC[9].icell.Ien Vbias 0.19173f
C1780 XA.Cn[12] XA.XIR[6].XIC[12].icell.Ien 0.04604f
C1781 XA.XIR[9].XIC[9].icell.Ien Iout 0.06801f
C1782 XThR.XTB7.Y XThR.XTBN.A 1.11559f
C1783 XA.Cn[8] Vbias 0.79784f
C1784 XThR.Tn[11] XA.XIR[11].XIC[9].icell.Ien 0.14211f
C1785 XThR.XTB5.A XThR.XTB7.A 0.07862f
C1786 XThR.XTB7.Y XThR.Tn[6] 0.21438f
C1787 XA.XIR[0].XIC[2].icell.Ien Iout 0.0675f
C1788 XA.XIR[7].XIC[13].icell.PDM VPWR 0.01171f
C1789 XA.Cn[6] XThR.Tn[9] 0.40738f
C1790 XA.Cn[7] XThR.Tn[8] 0.40738f
C1791 XThR.Tn[0] XA.XIR[0].XIC[14].icell.Ien 0.144f
C1792 XA.Cn[9] XA.XIR[15].XIC[9].icell.PDM 0.02601f
C1793 XA.Cn[0] XA.XIR[14].XIC[0].icell.Ien 0.04604f
C1794 XThR.Tn[6] XA.XIR[6].XIC[8].icell.Ien 0.14211f
C1795 XA.XIR[14].XIC_15.icell.Ien Iout 0.0694f
C1796 XA.XIR[7].XIC[5].icell.Ien Iout 0.06801f
C1797 XA.Cn[0] XThR.Tn[13] 0.40741f
C1798 a_n1049_7787# VPWR 0.72173f
C1799 XThR.Tn[7] XA.XIR[7].XIC_15.icell.Ien 0.13564f
C1800 XA.XIR[9].XIC[9].icell.PDM VPWR 0.01171f
C1801 XA.Cn[7] XA.XIR[7].XIC[7].icell.PDM 0.02601f
C1802 XA.XIR[6].XIC[4].icell.PDM Vbias 0.03928f
C1803 XA.XIR[0].XIC[1].icell.PDM VPWR 0.01132f
C1804 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.Ien 0.04854f
C1805 XA.XIR[14].XIC[1].icell.PDM Vbias 0.03928f
C1806 XA.XIR[5].XIC[11].icell.PDM Vbias 0.03928f
C1807 XA.Cn[3] XA.XIR[2].XIC[3].icell.Ien 0.04605f
C1808 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.Ien 0.04854f
C1809 XA.Cn[10] XA.XIR[2].XIC[10].icell.PDM 0.02602f
C1810 XA.XIR[13].XIC[5].icell.PDM Vbias 0.03928f
C1811 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.Ien 0.04854f
C1812 XA.Cn[13] XThR.Tn[7] 0.40739f
C1813 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.Ien 0.04854f
C1814 XA.XIR[12].XIC[10].icell.PDM Vbias 0.03928f
C1815 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PDM 0.04035f
C1816 XThR.XTBN.Y XThR.Tn[5] 0.59911f
C1817 XA.XIR[3].XIC[10].icell.Ien VPWR 0.18829f
C1818 XA.XIR[1].XIC[14].icell.PDM VPWR 0.0118f
C1819 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout 0.06446f
C1820 XA.XIR[6].XIC_15.icell.PUM VPWR 0.01655f
C1821 XA.XIR[10].XIC[14].icell.PDM VPWR 0.0118f
C1822 thermo15c_0.XTB5.A thermo15c_0.XTB1.Y 0.1098f
C1823 XA.XIR[14].XIC_dummy_right.icell.Iout Iout 0.01732f
C1824 XThR.XTBN.A a_n997_2667# 0.01679f
C1825 XThR.Tn[3] XThR.Tn[4] 0.1175f
C1826 XA.XIR[15].XIC[11].icell.PDM Vbias 0.03928f
C1827 XA.XIR[2].XIC[3].icell.Ien VPWR 0.18829f
C1828 XA.XIR[4].XIC[14].icell.PDM VPWR 0.0118f
C1829 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR 0.01493f
C1830 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PDM 0.04035f
C1831 XA.XIR[13].XIC_15.icell.PDM VPWR 0.07527f
C1832 XA.XIR[1].XIC[5].icell.Ien VPWR 0.18829f
C1833 XA.XIR[6].XIC[9].icell.Ien Vbias 0.19161f
C1834 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PDM 0.0404f
C1835 XA.XIR[8].XIC[13].icell.Ien VPWR 0.18829f
C1836 a_4067_9615# XA.Cn[2] 0.27296f
C1837 thermo15c_0.XTB4.Y Vbias 0.01644f
C1838 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.Ien 0.04854f
C1839 XA.XIR[3].XIC[6].icell.PDM Vbias 0.03928f
C1840 XA.XIR[14].XIC[3].icell.Ien Vbias 0.19161f
C1841 XA.XIR[8].XIC[8].icell.PDM Vbias 0.03928f
C1842 XA.XIR[2].XIC[12].icell.PDM Vbias 0.03928f
C1843 XA.XIR[13].XIC[5].icell.Ien Vbias 0.19161f
C1844 XThR.XTB6.Y XThR.XTB7.Y 2.05133f
C1845 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PDM 0.04035f
C1846 XA.Cn[14] XA.XIR[14].XIC[14].icell.PDM 0.02601f
C1847 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.Ien 0.04854f
C1848 XA.Cn[11] XThR.Tn[3] 0.40738f
C1849 XThR.XTBN.A XThR.Tn[11] 0.11968f
C1850 XA.XIR[3].XIC[2].icell.Ien Iout 0.06801f
C1851 XA.XIR[0].XIC_15.icell.Ien VPWR 0.26622f
C1852 XA.XIR[11].XIC[8].icell.Ien Vbias 0.19161f
C1853 XA.Cn[14] XA.XIR[9].XIC[14].icell.Ien 0.04604f
C1854 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.04035f
C1855 XThR.Tn[14] XA.XIR[14].XIC[4].icell.Ien 0.14211f
C1856 XThR.Tn[11] XA.XIR[11].XIC[14].icell.Ien 0.144f
C1857 XThR.Tn[1] XA.XIR[1].XIC[4].icell.Ien 0.14211f
C1858 XA.XIR[15].XIC[8].icell.Ien Iout 0.07192f
C1859 XA.Cn[5] XA.XIR[3].XIC[5].icell.PDM 0.02601f
C1860 XA.XIR[4].XIC_dummy_right.icell.Iout XA.XIR[5].XIC_dummy_right.icell.Iout 0.04047f
C1861 XA.XIR[6].XIC[0].icell.Ien VPWR 0.18829f
C1862 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PDM 0.04035f
C1863 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout 0.06446f
C1864 XA.Cn[12] XThR.Tn[5] 0.40738f
C1865 XA.Cn[10] XA.XIR[7].XIC[10].icell.PDM 0.02601f
C1866 XThR.XTB5.A XThR.XTB7.B 0.30355f
C1867 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.Ien 0.04854f
C1868 XA.XIR[4].XIC[11].icell.Ien Iout 0.06801f
C1869 XA.XIR[15].XIC_dummy_left.icell.Iout VPWR 0.24997f
C1870 thermo15c_0.XTB1.Y thermo15c_0.XTBN.Y 0.1979f
C1871 XThR.Tn[13] XA.XIR[13].XIC[8].icell.Ien 0.14211f
C1872 XA.Cn[1] XA.XIR[4].XIC[1].icell.Ien 0.04604f
C1873 XA.XIR[8].XIC[5].icell.Ien Iout 0.06801f
C1874 XA.Cn[8] XThR.Tn[0] 0.40759f
C1875 XA.XIR[11].XIC[4].icell.PDM VPWR 0.01171f
C1876 XA.Cn[5] VPWR 3.59867f
C1877 XA.XIR[2].XIC[12].icell.Ien Vbias 0.19161f
C1878 XA.XIR[10].XIC[8].icell.PDM VPWR 0.01171f
C1879 XA.XIR[0].XIC_dummy_right.icell.Iout VPWR 0.12361f
C1880 XA.XIR[11].XIC_dummy_right.icell.Iout XA.XIR[12].XIC_dummy_right.icell.Iout 0.04047f
C1881 XA.XIR[1].XIC[14].icell.Ien Vbias 0.19173f
C1882 XA.XIR[9].XIC[14].icell.Ien Iout 0.06801f
C1883 thermo15c_0.XTB7.Y XA.Cn[9] 0.07413f
C1884 XA.XIR[6].XIC[5].icell.Ien VPWR 0.18829f
C1885 XThR.XTB6.A XThR.XTB5.Y 0.01866f
C1886 XA.XIR[0].XIC[7].icell.Ien Iout 0.0675f
C1887 XA.XIR[12].XIC[1].icell.Ien Vbias 0.19161f
C1888 XA.Cn[2] XA.XIR[1].XIC[2].icell.PDM 0.02602f
C1889 XA.Cn[9] XA.XIR[4].XIC[9].icell.Ien 0.04604f
C1890 XThR.Tn[6] XA.XIR[6].XIC[13].icell.Ien 0.14211f
C1891 XA.Cn[2] XA.XIR[4].XIC[2].icell.PDM 0.02601f
C1892 XA.XIR[2].XIC[0].icell.PDM VPWR 0.01171f
C1893 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR 0.01669f
C1894 XA.XIR[7].XIC[10].icell.Ien Iout 0.06801f
C1895 XA.XIR[5].XIC[2].icell.Ien Vbias 0.19161f
C1896 XA.XIR[7].XIC[12].icell.PDM Vbias 0.03928f
C1897 XA.XIR[10].XIC[13].icell.PDM VPWR 0.01171f
C1898 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.Ien 0.04854f
C1899 XA.XIR[15].XIC[10].icell.PDM Vbias 0.03928f
C1900 thermo15c_0.XTB7.B XA.Cn[10] 0.0672f
C1901 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR 0.08055f
C1902 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PDM 0.04042f
C1903 XA.XIR[11].XIC[4].icell.Ien VPWR 0.18829f
C1904 XA.XIR[13].XIC[14].icell.PDM VPWR 0.0118f
C1905 XA.XIR[8].XIC[0].icell.Ien Iout 0.06795f
C1906 XA.XIR[10].XIC[6].icell.Ien VPWR 0.18829f
C1907 XA.Cn[4] Vbias 0.84011f
C1908 XThR.Tn[11] XA.XIR[11].XIC[12].icell.Ien 0.14211f
C1909 XA.Cn[11] XA.XIR[2].XIC[11].icell.Ien 0.04605f
C1910 thermo15c_0.XTBN.Y a_8963_9569# 0.22784f
C1911 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.Ien 0.04854f
C1912 XA.XIR[9].XIC[8].icell.PDM Vbias 0.03928f
C1913 thermo15c_0.XTB2.Y a_3773_9615# 0.2342f
C1914 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.Ien 0.04854f
C1915 XA.XIR[0].XIC[0].icell.PDM Vbias 0.03932f
C1916 XA.XIR[3].XIC_15.icell.Ien VPWR 0.26829f
C1917 XA.Cn[8] XA.XIR[3].XIC[8].icell.PDM 0.02601f
C1918 XThR.XTB6.Y XThR.Tn[11] 0.02465f
C1919 thermo15c_0.XTB7.A thermo15c_0.XTB5.Y 0.11935f
C1920 thermo15c_0.XTB6.A thermo15c_0.XTB7.B 1.47641f
C1921 XThR.XTB1.Y XThR.XTB6.A 0.01609f
C1922 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR 0.39039f
C1923 XA.XIR[2].XIC[8].icell.Ien VPWR 0.18829f
C1924 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Iout 0.01758f
C1925 a_3773_9615# VPWR 0.70508f
C1926 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR 0.38912f
C1927 XA.XIR[1].XIC[10].icell.Ien VPWR 0.18829f
C1928 XThR.Tn[8] XA.XIR[8].XIC[5].icell.Ien 0.14211f
C1929 XA.XIR[1].XIC[13].icell.PDM Vbias 0.03928f
C1930 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PDM 0.04035f
C1931 XA.Cn[11] XThR.Tn[11] 0.40738f
C1932 XA.XIR[6].XIC[14].icell.Ien Vbias 0.19161f
C1933 XA.Cn[6] XA.XIR[8].XIC[6].icell.PDM 0.02601f
C1934 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.PDM 0.02104f
C1935 XA.XIR[4].XIC[13].icell.PDM Vbias 0.03928f
C1936 XThR.XTB1.Y XThR.Tn[0] 0.1837f
C1937 XA.XIR[14].XIC[8].icell.Ien Vbias 0.19161f
C1938 XA.XIR[3].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1939 XThR.Tn[5] XA.XIR[5].XIC[4].icell.Ien 0.14211f
C1940 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.Ien 0.04854f
C1941 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.04035f
C1942 XA.XIR[7].XIC[0].icell.PDM VPWR 0.01171f
C1943 XThR.XTB7.B XThR.Tn[9] 0.0565f
C1944 XA.XIR[3].XIC[7].icell.Ien Iout 0.06801f
C1945 XA.XIR[6].XIC[7].icell.PDM VPWR 0.01171f
C1946 XThR.Tn[1] XA.XIR[1].XIC[9].icell.Ien 0.14211f
C1947 XThR.Tn[14] XA.XIR[14].XIC[9].icell.Ien 0.14211f
C1948 XA.XIR[5].XIC[14].icell.PDM VPWR 0.0118f
C1949 XA.XIR[14].XIC[4].icell.PDM VPWR 0.01171f
C1950 XThR.XTB5.A XThR.XTB4.Y 0.02767f
C1951 XA.Cn[8] XThR.Tn[1] 0.40744f
C1952 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.PDM 0.02104f
C1953 XA.XIR[13].XIC[8].icell.PDM VPWR 0.01171f
C1954 XA.XIR[1].XIC[2].icell.Ien Iout 0.06801f
C1955 XThR.Tn[11] XA.XIR[11].XIC[10].icell.Ien 0.14211f
C1956 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.PDM 0.02104f
C1957 XA.Cn[0] XThR.Tn[7] 0.40736f
C1958 XA.Cn[8] XThR.Tn[12] 0.40738f
C1959 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8] 0.14211f
C1960 XA.XIR[8].XIC[10].icell.Ien Iout 0.06801f
C1961 thermo15c_0.XTB1.Y thermo15c_0.XTBN.A 0.12307f
C1962 thermo15c_0.XTB1.Y a_7651_9569# 0.06353f
C1963 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1964 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.Ien 0.04854f
C1965 XA.XIR[10].XIC[12].icell.PDM VPWR 0.01171f
C1966 XA.Cn[7] XThR.Tn[3] 0.40738f
C1967 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.Ien 0.04854f
C1968 XA.XIR[1].XIC[1].icell.PDM VPWR 0.01171f
C1969 XA.Cn[2] XA.XIR[10].XIC[2].icell.Ien 0.04604f
C1970 XA.XIR[11].XIC[3].icell.PDM Vbias 0.03928f
C1971 XA.XIR[6].XIC[10].icell.Ien VPWR 0.18829f
C1972 XA.Cn[7] XA.XIR[12].XIC[7].icell.PDM 0.02601f
C1973 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11] 0.14211f
C1974 XA.Cn[13] XA.Cn[14] 0.3543f
C1975 XA.XIR[4].XIC[1].icell.PDM VPWR 0.01171f
C1976 XA.XIR[0].XIC[12].icell.Ien Iout 0.0675f
C1977 XA.XIR[10].XIC[7].icell.PDM Vbias 0.03928f
C1978 XA.XIR[13].XIC[13].icell.PDM VPWR 0.01171f
C1979 XA.XIR[8].XIC[11].icell.PDM VPWR 0.01171f
C1980 XA.XIR[3].XIC[9].icell.PDM VPWR 0.01171f
C1981 XA.XIR[14].XIC[4].icell.Ien VPWR 0.18883f
C1982 XThR.XTB5.Y XThR.Tn[12] 0.32095f
C1983 XA.Cn[9] XA.XIR[8].XIC[9].icell.PDM 0.02601f
C1984 XA.XIR[2].XIC_15.icell.PDM VPWR 0.07527f
C1985 thermo15c_0.XTB6.Y XA.Cn[12] 0.0253f
C1986 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.PDM 0.02104f
C1987 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PDM 0.0404f
C1988 XA.XIR[13].XIC[6].icell.Ien VPWR 0.18829f
C1989 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PDM 0.04035f
C1990 XA.XIR[7].XIC_15.icell.Ien Iout 0.0694f
C1991 XA.XIR[5].XIC[7].icell.Ien Vbias 0.19161f
C1992 XA.Cn[8] XA.XIR[9].XIC[8].icell.Ien 0.04604f
C1993 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout 0.06446f
C1994 XA.XIR[11].XIC_15.icell.PUM VPWR 0.01655f
C1995 XA.XIR[5].XIC[0].icell.Ien Iout 0.06795f
C1996 XA.Cn[4] XThR.Tn[0] 0.40763f
C1997 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1998 XA.XIR[4].XIC_dummy_left.icell.Iout Iout 0.03553f
C1999 XA.XIR[11].XIC[9].icell.Ien VPWR 0.18829f
C2000 XA.Cn[6] XA.XIR[9].XIC[6].icell.PDM 0.02601f
C2001 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2002 XA.Cn[13] Iout 0.22423f
C2003 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.PDM 0.02104f
C2004 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.PDM 0.02104f
C2005 XA.XIR[12].XIC[2].icell.Ien Vbias 0.19161f
C2006 XThR.XTB3.Y XThR.XTBN.A 0.03907f
C2007 XA.XIR[0].XIC_15.icell.PDM Vbias 0.03947f
C2008 thermo15c_0.XTB6.Y thermo15c_0.XTBN.Y 0.18947f
C2009 XA.XIR[6].XIC[2].icell.Ien Iout 0.06801f
C2010 XA.Cn[11] XThR.Tn[14] 0.40738f
C2011 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.PDM 0.02104f
C2012 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Iout 0.01728f
C2013 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PDM 0.0404f
C2014 XA.Cn[7] XA.XIR[11].XIC[7].icell.Ien 0.04604f
C2015 thermo15c_0.XTBN.A a_8963_9569# 0.01679f
C2016 XA.XIR[7].XIC_dummy_right.icell.Iout Iout 0.01732f
C2017 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PDM 0.04035f
C2018 thermo15c_0.XTB3.Y data[0] 0.03253f
C2019 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.Ien 0.04854f
C2020 XA.XIR[2].XIC[13].icell.Ien VPWR 0.18829f
C2021 XThR.XTBN.Y XThR.Tn[9] 0.48067f
C2022 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2023 XA.Cn[2] XA.XIR[5].XIC[2].icell.PDM 0.02601f
C2024 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.PDM 0.02104f
C2025 XA.XIR[1].XIC_15.icell.Ien VPWR 0.26829f
C2026 XThR.Tn[8] XA.XIR[8].XIC[10].icell.Ien 0.14211f
C2027 XThR.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.144f
C2028 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.Ien 0.04854f
C2029 XA.Cn[3] XA.XIR[5].XIC[3].icell.Ien 0.04604f
C2030 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.PDM 0.02104f
C2031 thermo15c_0.XTB7.B XA.Cn[6] 0.04318f
C2032 XA.Cn[0] XA.XIR[9].XIC[0].icell.Ien 0.04604f
C2033 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR 0.35555f
C2034 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.PDM 0.02104f
C2035 XThR.Tn[11] XA.XIR[11].XIC_15.icell.Ien 0.13564f
C2036 XA.Cn[2] XThR.Tn[2] 0.40741f
C2037 a_2979_9615# Vbias 0.01381f
C2038 XA.Cn[10] XA.XIR[12].XIC[10].icell.PDM 0.02601f
C2039 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.Ien 0.04854f
C2040 XA.XIR[10].XIC[3].icell.Ien Iout 0.06801f
C2041 XThR.Tn[5] XA.XIR[5].XIC[9].icell.Ien 0.14211f
C2042 XA.Cn[5] XA.XIR[0].XIC[5].icell.Ien 0.04659f
C2043 XThR.XTB4.Y XThR.Tn[9] 0.01318f
C2044 XA.XIR[5].XIC[3].icell.Ien VPWR 0.18829f
C2045 XA.XIR[7].XIC_15.icell.PDM VPWR 0.07527f
C2046 XA.Cn[3] XA.XIR[0].XIC[3].icell.PDM 0.02804f
C2047 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.Ien 0.04854f
C2048 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.Ien 0.04854f
C2049 XA.XIR[3].XIC[12].icell.Ien Iout 0.06801f
C2050 XThR.Tn[9] XThR.Tn[10] 0.12586f
C2051 XA.XIR[1].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2052 XThR.Tn[0] Vbias 1.40808f
C2053 XThR.Tn[1] XA.XIR[1].XIC[14].icell.Ien 0.144f
C2054 XA.XIR[10].XIC[11].icell.PDM VPWR 0.01171f
C2055 XA.XIR[2].XIC[5].icell.Ien Iout 0.06801f
C2056 XA.Cn[7] XThR.Tn[11] 0.40738f
C2057 XA.Cn[0] XA.XIR[10].XIC[0].icell.PDM 0.02601f
C2058 XA.Cn[3] XThR.Tn[6] 0.40738f
C2059 XA.XIR[1].XIC[7].icell.Ien Iout 0.06801f
C2060 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.Ien 0.04854f
C2061 thermo15c_0.XTB4.Y XA.Cn[10] 0.01405f
C2062 XA.XIR[6].XIC[6].icell.PDM Vbias 0.03928f
C2063 XA.XIR[9].XIC[11].icell.PDM VPWR 0.01171f
C2064 XA.XIR[13].XIC[12].icell.PDM VPWR 0.01171f
C2065 XA.Cn[9] XA.XIR[9].XIC[9].icell.PDM 0.02601f
C2066 XA.XIR[0].XIC[3].icell.PDM VPWR 0.01132f
C2067 XA.Cn[2] XA.XIR[13].XIC[2].icell.Ien 0.04604f
C2068 XA.Cn[7] XA.XIR[15].XIC[7].icell.PDM 0.02601f
C2069 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.Ien 0.04854f
C2070 XA.XIR[14].XIC[3].icell.PDM Vbias 0.03928f
C2071 XA.XIR[5].XIC[13].icell.PDM Vbias 0.03928f
C2072 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.Ien 0.04854f
C2073 XThR.XTB3.Y a_n1049_7493# 0.23056f
C2074 XA.Cn[12] XThR.Tn[9] 0.40738f
C2075 XA.XIR[8].XIC_15.icell.Ien Iout 0.0694f
C2076 XA.Cn[13] XThR.Tn[8] 0.40739f
C2077 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.Ien 0.04854f
C2078 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.Ien 0.04854f
C2079 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.PDM 0.02104f
C2080 XThR.XTBN.A VPWR 0.90694f
C2081 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.PDM 0.02104f
C2082 XA.XIR[13].XIC[7].icell.PDM Vbias 0.03928f
C2083 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12] 0.14211f
C2084 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.PDM 0.02104f
C2085 XThR.XTB5.Y a_n1049_6405# 0.24821f
C2086 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PDM 0.04035f
C2087 XThR.Tn[6] VPWR 7.9997f
C2088 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PDM 0.04042f
C2089 XA.XIR[11].XIC[14].icell.Ien VPWR 0.18835f
C2090 thermo15c_0.XTB6.A thermo15c_0.XTB4.Y 0.04137f
C2091 thermo15c_0.XTB7.A thermo15c_0.XTB3.Y 0.57441f
C2092 XThR.XTB3.Y XThR.XTB6.Y 0.04428f
C2093 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2094 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.PDM 0.02104f
C2095 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Ien 0.01532f
C2096 XA.XIR[6].XIC_15.icell.Ien VPWR 0.26829f
C2097 XA.XIR[9].XIC[3].icell.Ien Vbias 0.19161f
C2098 XA.Cn[5] XA.XIR[6].XIC[5].icell.PDM 0.02601f
C2099 XThR.Tn[14] XA.XIR[14].XIC[12].icell.Ien 0.14211f
C2100 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.Ien 0.04854f
C2101 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2102 XA.XIR[14].XIC_15.icell.PUM VPWR 0.01655f
C2103 XA.Cn[4] XThR.Tn[1] 0.40744f
C2104 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.PDM 0.02104f
C2105 XA.XIR[1].XIC[0].icell.PDM Vbias 0.03915f
C2106 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.Ien 0.04854f
C2107 XA.XIR[14].XIC[9].icell.Ien VPWR 0.18883f
C2108 XA.XIR[8].XIC_dummy_right.icell.Iout Iout 0.01732f
C2109 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.Ien 0.04854f
C2110 XA.Cn[4] XThR.Tn[12] 0.40738f
C2111 XA.XIR[5].XIC[12].icell.Ien Vbias 0.19161f
C2112 XA.XIR[4].XIC[0].icell.PDM Vbias 0.03915f
C2113 data[2] data[3] 0.04128f
C2114 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR 0.38902f
C2115 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2116 XThR.Tn[3] XA.XIR[3].XIC[2].icell.Ien 0.14211f
C2117 XA.XIR[8].XIC[10].icell.PDM Vbias 0.03928f
C2118 XA.XIR[3].XIC[8].icell.PDM Vbias 0.03928f
C2119 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0222f
C2120 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.PDM 0.02104f
C2121 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.Ien 0.04854f
C2122 XA.XIR[2].XIC[14].icell.PDM Vbias 0.03928f
C2123 XA.XIR[6].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2124 XA.Cn[7] XA.XIR[14].XIC[7].icell.Ien 0.04604f
C2125 XA.Cn[3] XThR.Tn[4] 0.40738f
C2126 XA.Cn[5] XA.XIR[3].XIC[5].icell.Ien 0.04604f
C2127 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PDM 0.04035f
C2128 XA.XIR[14].XIC_dummy_right.icell.Iout XA.XIR[15].XIC_dummy_right.icell.Iout 0.04047f
C2129 XA.XIR[12].XIC[7].icell.Ien Vbias 0.19161f
C2130 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PDM 0.04035f
C2131 XA.XIR[6].XIC[7].icell.Ien Iout 0.06801f
C2132 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.PDM 0.02104f
C2133 XA.XIR[5].XIC[1].icell.PDM VPWR 0.01171f
C2134 XA.Cn[2] XThR.Tn[10] 0.40738f
C2135 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PDM 0.04035f
C2136 thermo15c_0.XTBN.A thermo15c_0.XTB6.Y 0.06405f
C2137 XThR.Tn[4] VPWR 8.03623f
C2138 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.PDM 0.02104f
C2139 XA.Cn[10] XA.XIR[15].XIC[10].icell.PDM 0.02601f
C2140 XA.XIR[12].XIC[0].icell.PDM VPWR 0.01171f
C2141 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.Ien 0.04854f
C2142 XA.XIR[13].XIC[3].icell.Ien Iout 0.06801f
C2143 a_n1049_7493# VPWR 0.72084f
C2144 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.Ien 0.04854f
C2145 XThR.Tn[8] XA.XIR[8].XIC_15.icell.Ien 0.13564f
C2146 XA.XIR[11].XIC[6].icell.PDM VPWR 0.01171f
C2147 XA.XIR[11].XIC[12].icell.Ien VPWR 0.18829f
C2148 XA.Cn[11] XA.XIR[5].XIC[11].icell.Ien 0.04604f
C2149 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.Ien 0.04854f
C2150 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.PDM 0.02104f
C2151 XA.XIR[10].XIC[10].icell.PDM VPWR 0.01171f
C2152 XA.XIR[1].XIC[0].icell.Ien Vbias 0.1916f
C2153 XThR.Tn[14] XA.XIR[14].XIC[10].icell.Ien 0.14211f
C2154 XA.XIR[11].XIC[6].icell.Ien Iout 0.06801f
C2155 XThR.XTB6.Y VPWR 1.05512f
C2156 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.PDM 0.02104f
C2157 XA.Cn[8] XA.XIR[6].XIC[8].icell.PDM 0.02601f
C2158 XA.Cn[4] XA.XIR[7].XIC[4].icell.Ien 0.04604f
C2159 XA.XIR[4].XIC[0].icell.Ien Vbias 0.19149f
C2160 XA.Cn[11] XA.XIR[2].XIC[11].icell.PDM 0.02602f
C2161 XThR.Tn[1] Vbias 1.39552f
C2162 XA.XIR[10].XIC[8].icell.Ien Iout 0.06801f
C2163 VPWR data[3] 0.20846f
C2164 XA.XIR[13].XIC[11].icell.PDM VPWR 0.01171f
C2165 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.PDM 0.02104f
C2166 XThR.Tn[5] XA.XIR[5].XIC[14].icell.Ien 0.144f
C2167 XA.Cn[3] XA.XIR[12].XIC[3].icell.Ien 0.04604f
C2168 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.Ien 0.04854f
C2169 XA.Cn[7] XThR.Tn[14] 0.40738f
C2170 XA.Cn[0] XA.XIR[13].XIC[0].icell.PDM 0.02601f
C2171 XA.Cn[13] XA.XIR[0].XIC[13].icell.Ien 0.04662f
C2172 XA.XIR[5].XIC[8].icell.Ien VPWR 0.18829f
C2173 XA.XIR[10].XIC_dummy_left.icell.Iout VPWR 0.11161f
C2174 XA.XIR[8].XIC_dummy_right.icell.Iout XA.XIR[9].XIC_dummy_right.icell.Iout 0.04047f
C2175 XThR.Tn[12] Vbias 1.39531f
C2176 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.PDM 0.02104f
C2177 XA.Cn[11] VPWR 4.57828f
C2178 thermo15c_0.XTBN.Y XA.Cn[2] 0.49723f
C2179 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.PDM 0.02104f
C2180 XA.XIR[2].XIC[2].icell.PDM VPWR 0.01171f
C2181 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.PDM 0.02104f
C2182 XA.XIR[15].XIC[2].icell.Ien Vbias 0.15966f
C2183 XA.XIR[2].XIC[10].icell.Ien Iout 0.06801f
C2184 XA.XIR[7].XIC[14].icell.PDM Vbias 0.03928f
C2185 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.PDM 0.02104f
C2186 XA.XIR[1].XIC[12].icell.Ien Iout 0.06801f
C2187 XA.XIR[12].XIC[3].icell.Ien VPWR 0.18829f
C2188 XA.Cn[0] Iout 0.07042f
C2189 XA.XIR[4].XIC[5].icell.Ien Vbias 0.19161f
C2190 XA.XIR[14].XIC[14].icell.Ien VPWR 0.1889f
C2191 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.Ien 0.04854f
C2192 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PDM 0.04035f
C2193 a_4861_9615# XA.Cn[3] 0.26251f
C2194 thermo15c_0.XTBN.Y a_10051_9569# 0.23006f
C2195 XThR.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.14211f
C2196 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.PDM 0.02104f
C2197 XA.XIR[9].XIC[10].icell.PDM Vbias 0.03928f
C2198 XA.XIR[0].XIC[2].icell.PDM Vbias 0.03945f
C2199 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.PDM 0.02104f
C2200 data[5] data[4] 0.64735f
C2201 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.0404f
C2202 XA.XIR[9].XIC[8].icell.Ien Vbias 0.19161f
C2203 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.Ien 0.04854f
C2204 XThR.Tn[10] XA.XIR[10].XIC[13].icell.Ien 0.14211f
C2205 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.PDM 0.02104f
C2206 XA.XIR[11].XIC[10].icell.Ien VPWR 0.18829f
C2207 a_4861_9615# VPWR 0.70519f
C2208 XA.Cn[10] Vbias 0.81591f
C2209 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PDM 0.04035f
C2210 XA.XIR[1].XIC_15.icell.PDM Vbias 0.03927f
C2211 XA.Cn[6] XA.XIR[3].XIC[6].icell.PDM 0.02601f
C2212 XA.Cn[11] XA.XIR[7].XIC[11].icell.PDM 0.02601f
C2213 XA.XIR[7].XIC[4].icell.Ien Vbias 0.19161f
C2214 XA.XIR[4].XIC_15.icell.PDM Vbias 0.03927f
C2215 XThR.Tn[12] XA.XIR[12].XIC[2].icell.Ien 0.14211f
C2216 XThR.Tn[3] XA.XIR[3].XIC[7].icell.Ien 0.14211f
C2217 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.PDM 0.02104f
C2218 XA.XIR[12].XIC[13].icell.Ien Iout 0.06801f
C2219 XA.XIR[11].XIC[0].icell.Ien VPWR 0.18829f
C2220 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.PDM 0.02104f
C2221 XA.Cn[2] XThR.Tn[13] 0.40738f
C2222 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PDM 0.04035f
C2223 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2224 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.PDM 0.02104f
C2225 XA.XIR[7].XIC[2].icell.PDM VPWR 0.01171f
C2226 XThR.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.14211f
C2227 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2228 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.PDM 0.02104f
C2229 XThR.Tn[14] XA.XIR[14].XIC_15.icell.Ien 0.13564f
C2230 XA.Cn[13] XA.XIR[3].XIC[13].icell.Ien 0.04604f
C2231 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.Ien 0.04854f
C2232 XA.XIR[6].XIC[9].icell.PDM VPWR 0.01171f
C2233 XA.XIR[15].XIC[0].icell.PDM VPWR 0.01512f
C2234 XA.XIR[6].XIC[12].icell.Ien Iout 0.06801f
C2235 XA.Cn[4] XA.XIR[8].XIC[4].icell.Ien 0.04604f
C2236 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.PDM 0.02104f
C2237 XA.XIR[14].XIC[6].icell.PDM VPWR 0.01171f
C2238 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.PDM 0.02104f
C2239 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2240 XA.XIR[14].XIC[12].icell.Ien VPWR 0.18883f
C2241 XA.Cn[5] XA.XIR[1].XIC[5].icell.Ien 0.04606f
C2242 thermo15c_0.XTB6.Y a_6243_9615# 0.01199f
C2243 XA.Cn[0] XA.XIR[3].XIC[0].icell.Ien 0.04604f
C2244 XA.Cn[0] XThR.Tn[8] 0.40736f
C2245 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.PDM 0.02104f
C2246 XA.XIR[13].XIC[10].icell.PDM VPWR 0.01171f
C2247 XA.XIR[14].XIC[6].icell.Ien Iout 0.06801f
C2248 XA.Cn[3] XA.XIR[1].XIC[3].icell.PDM 0.02602f
C2249 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.Ien 0.04854f
C2250 XA.XIR[5].XIC[0].icell.PDM Vbias 0.03915f
C2251 XA.XIR[13].XIC[8].icell.Ien Iout 0.06801f
C2252 XA.Cn[3] XA.XIR[4].XIC[3].icell.PDM 0.02601f
C2253 XA.XIR[9].XIC[4].icell.Ien VPWR 0.18829f
C2254 XThR.Tn[0] XThR.Tn[1] 0.27134f
C2255 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.Ien 0.04854f
C2256 XA.XIR[13].XIC_dummy_left.icell.Iout VPWR 0.11047f
C2257 XThR.XTB7.A XThR.XTB5.Y 0.11935f
C2258 XThR.Tn[10] XA.XIR[10].XIC[11].icell.Ien 0.14211f
C2259 XA.XIR[1].XIC[3].icell.PDM VPWR 0.01171f
C2260 XA.XIR[11].XIC[5].icell.PDM Vbias 0.03928f
C2261 XA.Cn[12] XA.XIR[7].XIC[12].icell.Ien 0.04604f
C2262 XA.XIR[10].XIC[9].icell.PDM Vbias 0.03928f
C2263 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Iout 0.01728f
C2264 XA.XIR[4].XIC[3].icell.PDM VPWR 0.01171f
C2265 XA.XIR[5].XIC[13].icell.Ien VPWR 0.18829f
C2266 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.PDM 0.02104f
C2267 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Iout 0.01728f
C2268 XA.XIR[8].XIC[13].icell.PDM VPWR 0.01171f
C2269 XA.XIR[3].XIC[11].icell.PDM VPWR 0.01171f
C2270 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2271 XA.Cn[9] XA.XIR[3].XIC[9].icell.PDM 0.02601f
C2272 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PDM 0.04035f
C2273 data[1] data[0] 0.64735f
C2274 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PDM 0.04035f
C2275 XA.XIR[2].XIC_15.icell.Ien Iout 0.0694f
C2276 XA.XIR[15].XIC[7].icell.Ien Vbias 0.15966f
C2277 XA.XIR[12].XIC[11].icell.Ien Iout 0.06801f
C2278 XA.Cn[13] XThR.Tn[3] 0.40739f
C2279 XA.XIR[11].XIC_15.icell.PDM VPWR 0.07527f
C2280 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.PDM 0.02104f
C2281 XA.XIR[11].XIC_15.icell.Ien VPWR 0.26829f
C2282 XA.XIR[12].XIC[8].icell.Ien VPWR 0.18829f
C2283 XA.XIR[4].XIC[10].icell.Ien Vbias 0.19161f
C2284 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.Ien 0.04854f
C2285 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2286 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.Ien 0.04854f
C2287 XA.XIR[0].XIC[1].icell.Ien Vbias 0.19213f
C2288 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.PDM 0.02104f
C2289 XA.Cn[9] XA.XIR[11].XIC[9].icell.Ien 0.04604f
C2290 XA.XIR[2].XIC[1].icell.PDM Vbias 0.03928f
C2291 XA.Cn[7] XA.XIR[8].XIC[7].icell.PDM 0.02601f
C2292 XA.Cn[14] XThR.Tn[5] 0.40742f
C2293 XA.XIR[8].XIC[4].icell.Ien Vbias 0.19161f
C2294 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.Ien 0.04854f
C2295 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.PDM 0.02104f
C2296 XThR.Tn[4] XA.XIR[4].XIC[9].icell.Ien 0.14211f
C2297 XA.Cn[5] XA.XIR[6].XIC[5].icell.Ien 0.04604f
C2298 XA.XIR[14].XIC[10].icell.Ien VPWR 0.18883f
C2299 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.Ien 0.04854f
C2300 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.Ien 0.04854f
C2301 XA.Cn[10] XThR.Tn[0] 0.40762f
C2302 XThR.XTB1.Y XThR.XTB7.A 0.48957f
C2303 XA.XIR[9].XIC[13].icell.Ien Vbias 0.19161f
C2304 XA.XIR[5].XIC[5].icell.Ien Iout 0.06801f
C2305 XA.Cn[7] VPWR 3.9785f
C2306 XA.XIR[2].XIC_dummy_right.icell.Iout Iout 0.01732f
C2307 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PDM 0.04056f
C2308 XA.XIR[11].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2309 XThR.Tn[7] XA.XIR[7].XIC[2].icell.Ien 0.14211f
C2310 XA.XIR[7].XIC_15.icell.PUM VPWR 0.01655f
C2311 XA.XIR[0].XIC[6].icell.Ien Vbias 0.19213f
C2312 XA.Cn[0] XA.Cn[1] 0.88262f
C2313 thermo15c_0.XTB1.Y thermo15c_0.XTB5.Y 0.05054f
C2314 thermo15c_0.XTB5.A thermo15c_0.XTB7.B 0.30355f
C2315 thermo15c_0.XTB7.Y XA.Cn[11] 0.07422f
C2316 XA.Cn[3] XA.XIR[15].XIC[3].icell.Ien 0.04292f
C2317 XA.Cn[12] XA.XIR[12].XIC[12].icell.PDM 0.02601f
C2318 XA.XIR[4].XIC[1].icell.Ien VPWR 0.18829f
C2319 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR 0.08252f
C2320 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.Ien 0.04854f
C2321 XThR.Tn[5] Iout 1.12761f
C2322 XThR.Tn[12] XA.XIR[12].XIC[7].icell.Ien 0.14211f
C2323 XA.XIR[7].XIC[9].icell.Ien Vbias 0.19161f
C2324 XThR.Tn[8] data[4] 0.01643f
C2325 Vbias bias[2] 0.06133f
C2326 XThR.Tn[3] XA.XIR[3].XIC[12].icell.Ien 0.14211f
C2327 XThR.XTBN.A data[7] 0.07741f
C2328 XA.XIR[15].XIC[3].icell.Ien VPWR 0.31713f
C2329 XA.XIR[10].XIC_dummy_right.icell.Iout XA.XIR[11].XIC_dummy_right.icell.Iout 0.04047f
C2330 XThR.Tn[2] XA.XIR[2].XIC[7].icell.Ien 0.14211f
C2331 XA.XIR[2].XIC[0].icell.Ien Vbias 0.19149f
C2332 thermo15c_0.XTB7.A data[1] 0.06544f
C2333 XA.XIR[14].XIC_dummy_left.icell.Ien XThR.Tn[14] 0.01244f
C2334 XA.XIR[4].XIC[6].icell.Ien VPWR 0.18829f
C2335 XThR.Tn[1] XA.XIR[1].XIC[0].icell.Ien 0.14251f
C2336 XA.Cn[6] Vbias 0.81928f
C2337 XA.Cn[12] XA.XIR[8].XIC[12].icell.Ien 0.04604f
C2338 XThR.XTB7.B XThR.XTB5.Y 0.30227f
C2339 XA.Cn[8] XThR.Tn[2] 0.40741f
C2340 XA.XIR[10].XIC[1].icell.Ien Vbias 0.19161f
C2341 XA.XIR[7].XIC[1].icell.PDM Vbias 0.03928f
C2342 XA.Cn[13] XA.XIR[1].XIC[13].icell.Ien 0.04606f
C2343 XA.XIR[9].XIC[13].icell.PDM VPWR 0.01171f
C2344 XA.XIR[6].XIC[8].icell.PDM Vbias 0.03928f
C2345 XA.Cn[10] XA.XIR[8].XIC[10].icell.PDM 0.02601f
C2346 XA.XIR[0].XIC[5].icell.PDM VPWR 0.01261f
C2347 XA.XIR[7].XIC[0].icell.Ien VPWR 0.18829f
C2348 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.PDM 0.02104f
C2349 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.Ien 0.04854f
C2350 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.PDM 0.02104f
C2351 XA.XIR[14].XIC[5].icell.PDM Vbias 0.03928f
C2352 XA.XIR[5].XIC_15.icell.PDM Vbias 0.03927f
C2353 XA.XIR[9].XIC[9].icell.Ien VPWR 0.18829f
C2354 thermo15c_0.XTB7.B thermo15c_0.XTBN.Y 0.38751f
C2355 XA.XIR[13].XIC[9].icell.PDM Vbias 0.03928f
C2356 XThR.Tn[9] XA.XIR[9].XIC[5].icell.Ien 0.14211f
C2357 XA.XIR[0].XIC[2].icell.Ien VPWR 0.18776f
C2358 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.Ien 0.04854f
C2359 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PDM 0.04035f
C2360 XA.XIR[11].XIC[14].icell.PDM VPWR 0.0118f
C2361 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PDM 0.04035f
C2362 XA.Cn[13] XThR.Tn[11] 0.40739f
C2363 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PDM 0.04035f
C2364 XA.Cn[7] XA.XIR[9].XIC[7].icell.PDM 0.02601f
C2365 XA.Cn[9] XThR.Tn[6] 0.40738f
C2366 XA.XIR[14].XIC_15.icell.PDM VPWR 0.07527f
C2367 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.PDM 0.02104f
C2368 XA.Cn[7] XA.XIR[9].XIC[7].icell.Ien 0.04604f
C2369 XA.XIR[7].XIC[5].icell.Ien VPWR 0.18829f
C2370 XA.XIR[11].XIC[13].icell.Ien Vbias 0.19161f
C2371 XA.XIR[14].XIC_15.icell.Ien VPWR 0.26861f
C2372 XA.XIR[15].XIC[13].icell.Ien Iout 0.07192f
C2373 XA.XIR[3].XIC[6].icell.Ien Vbias 0.19161f
C2374 XA.XIR[1].XIC[2].icell.PDM Vbias 0.03928f
C2375 XA.Cn[9] XA.XIR[14].XIC[9].icell.Ien 0.04604f
C2376 XThR.Tn[0] XA.XIR[0].XIC[1].icell.Ien 0.14211f
C2377 XThR.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.14211f
C2378 XA.XIR[4].XIC[2].icell.PDM Vbias 0.03928f
C2379 XA.XIR[8].XIC_15.icell.PUM VPWR 0.01655f
C2380 XThR.XTB7.B XThR.XTB1.Y 1.61695f
C2381 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.Ien 0.04854f
C2382 XA.Cn[3] XA.XIR[5].XIC[3].icell.PDM 0.02601f
C2383 XA.XIR[4].XIC_15.icell.Ien Vbias 0.19195f
C2384 XThR.XTB5.A data[5] 0.11096f
C2385 XA.XIR[3].XIC[10].icell.PDM Vbias 0.03928f
C2386 XA.XIR[8].XIC[12].icell.PDM Vbias 0.03928f
C2387 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.PDM 0.02104f
C2388 XA.Cn[10] XThR.Tn[1] 0.40744f
C2389 XA.XIR[8].XIC[9].icell.Ien Vbias 0.19161f
C2390 XA.XIR[14].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2391 XThR.Tn[4] XA.XIR[4].XIC[14].icell.Ien 0.144f
C2392 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PDM 0.04056f
C2393 XA.Cn[2] XThR.Tn[7] 0.40738f
C2394 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9] 0.14211f
C2395 XThR.Tn[0] XA.XIR[0].XIC[6].icell.Ien 0.14211f
C2396 XA.Cn[10] XThR.Tn[12] 0.40738f
C2397 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PDM 0.04035f
C2398 XA.Cn[13] XA.XIR[6].XIC[13].icell.Ien 0.04604f
C2399 XThR.Tn[10] XA.XIR[10].XIC[5].icell.Ien 0.14211f
C2400 XA.Cn[12] XA.XIR[15].XIC[12].icell.PDM 0.02601f
C2401 XA.XIR[11].XIC_dummy_left.icell.Iout Iout 0.03553f
C2402 XA.XIR[5].XIC[3].icell.PDM VPWR 0.01171f
C2403 XA.XIR[5].XIC[10].icell.Ien Iout 0.06801f
C2404 thermo15c_0.XTB7.Y a_6243_10571# 0.01283f
C2405 XA.Cn[4] XA.XIR[0].XIC[4].icell.PDM 0.02803f
C2406 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PDM 0.0404f
C2407 XA.Cn[2] XA.XIR[4].XIC[2].icell.Ien 0.04604f
C2408 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.Ien 0.04854f
C2409 XThR.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.14211f
C2410 XA.XIR[0].XIC[11].icell.Ien Vbias 0.19213f
C2411 XA.Cn[9] XThR.Tn[4] 0.40738f
C2412 thermo15c_0.XTB5.A a_7331_10587# 0.01243f
C2413 XA.XIR[12].XIC[2].icell.PDM VPWR 0.01171f
C2414 XA.XIR[11].XIC[8].icell.PDM VPWR 0.01171f
C2415 XA.Cn[1] XA.XIR[10].XIC[1].icell.PDM 0.02601f
C2416 XThR.XTBN.Y XThR.XTB5.Y 0.16186f
C2417 XA.XIR[12].XIC[5].icell.Ien Iout 0.06801f
C2418 XA.XIR[7].XIC[14].icell.Ien Vbias 0.19161f
C2419 XA.Cn[8] XThR.Tn[10] 0.40738f
C2420 XA.Cn[10] XA.XIR[9].XIC[10].icell.PDM 0.02601f
C2421 XA.XIR[11].XIC[11].icell.Ien Vbias 0.19161f
C2422 XA.XIR[3].XIC[2].icell.Ien VPWR 0.18829f
C2423 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PDM 0.04042f
C2424 XA.Cn[4] XA.XIR[2].XIC[4].icell.Ien 0.04605f
C2425 XA.XIR[15].XIC[11].icell.Ien Iout 0.07192f
C2426 thermo15c_0.XTB1.Y XA.Cn[1] 0.01068f
C2427 VPWR data[0] 0.52929f
C2428 XA.XIR[13].XIC[1].icell.Ien Vbias 0.19161f
C2429 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.PDM 0.02104f
C2430 XA.Cn[6] XThR.Tn[0] 0.40767f
C2431 XA.XIR[15].XIC[8].icell.Ien VPWR 0.31713f
C2432 XA.Cn[0] XThR.Tn[3] 0.40742f
C2433 XThR.Tn[2] XA.XIR[2].XIC[12].icell.Ien 0.14211f
C2434 XThR.Tn[13] XA.XIR[13].XIC[11].icell.Ien 0.14211f
C2435 XA.XIR[4].XIC[11].icell.Ien VPWR 0.18829f
C2436 XA.XIR[8].XIC[0].icell.PDM VPWR 0.01171f
C2437 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.PDM 0.02104f
C2438 XThR.XTB4.Y XThR.XTB5.Y 2.06459f
C2439 XA.XIR[2].XIC[4].icell.PDM VPWR 0.01171f
C2440 thermo15c_0.XTB7.Y XA.Cn[7] 0.08399f
C2441 XA.Cn[6] XA.XIR[6].XIC[6].icell.PDM 0.02601f
C2442 XA.XIR[11].XIC[13].icell.PDM VPWR 0.01171f
C2443 XA.XIR[8].XIC[5].icell.Ien VPWR 0.18829f
C2444 XA.Cn[1] XThR.Tn[5] 0.40738f
C2445 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Iout 0.01728f
C2446 XThR.XTB5.Y XThR.Tn[10] 0.01742f
C2447 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.Ien 0.04854f
C2448 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.Ien 0.04854f
C2449 XA.XIR[14].XIC[14].icell.PDM VPWR 0.0118f
C2450 XA.Cn[13] XThR.Tn[14] 0.40739f
C2451 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PDM 0.04035f
C2452 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout 0.06446f
C2453 XA.XIR[9].XIC[14].icell.Ien VPWR 0.18835f
C2454 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.PDM 0.02104f
C2455 XA.XIR[14].XIC[13].icell.Ien Vbias 0.19161f
C2456 thermo15c_0.XTB4.Y a_5155_9615# 0.01546f
C2457 thermo15c_0.XTBN.Y XA.Cn[8] 0.41222f
C2458 XThR.Tn[9] XA.XIR[9].XIC[10].icell.Ien 0.14211f
C2459 XA.XIR[9].XIC[12].icell.PDM Vbias 0.03928f
C2460 XThR.XTB1.Y XThR.XTBN.Y 0.20262f
C2461 XA.XIR[0].XIC[7].icell.Ien VPWR 0.18776f
C2462 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.Ien 0.04854f
C2463 XA.XIR[0].XIC[4].icell.PDM Vbias 0.03945f
C2464 thermo15c_0.XTB5.Y thermo15c_0.XTB6.Y 2.12831f
C2465 thermo15c_0.XTBN.A thermo15c_0.XTB7.B 0.35142f
C2466 thermo15c_0.XTB7.B a_7651_9569# 0.01152f
C2467 XA.XIR[1].XIC[1].icell.Ien Vbias 0.19173f
C2468 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PDM 0.04035f
C2469 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2470 XA.XIR[10].XIC[2].icell.Ien Vbias 0.19161f
C2471 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.PDM 0.02104f
C2472 XA.XIR[9].XIC[1].icell.Ien Iout 0.06801f
C2473 thermo15c_0.XTB7.A XA.Cn[3] 0.0337f
C2474 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.04035f
C2475 XThR.Tn[5] a_n1049_5611# 0.27042f
C2476 thermo15c_0.XTB1.Y thermo15c_0.XTB3.Y 0.04033f
C2477 thermo15c_0.XTB5.A thermo15c_0.XTB4.Y 0.02767f
C2478 XA.Cn[4] XThR.Tn[2] 0.40741f
C2479 thermo15c_0.XTB2.Y thermo15c_0.XTB7.A 0.2319f
C2480 XA.XIR[4].XIC[3].icell.Ien Iout 0.06801f
C2481 XA.XIR[7].XIC[10].icell.Ien VPWR 0.18829f
C2482 XA.XIR[0].XIC_dummy_right.icell.Iout XA.XIR[1].XIC_dummy_right.icell.Iout 0.04047f
C2483 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR 0.38902f
C2484 a_5949_9615# VPWR 0.7053f
C2485 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PDM 0.04035f
C2486 XA.XIR[3].XIC[11].icell.Ien Vbias 0.19161f
C2487 XThR.XTB1.Y XThR.XTB4.Y 0.05121f
C2488 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.PDM 0.02104f
C2489 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.Ien 0.04854f
C2490 XA.XIR[2].XIC[4].icell.Ien Vbias 0.19161f
C2491 XThR.Tn[6] XA.XIR[6].XIC[0].icell.Ien 0.14211f
C2492 XA.XIR[8].XIC[0].icell.Ien VPWR 0.18829f
C2493 thermo15c_0.XTB7.A VPWR 0.87269f
C2494 XA.XIR[1].XIC[6].icell.Ien Vbias 0.19173f
C2495 XA.XIR[9].XIC[6].icell.Ien Iout 0.06801f
C2496 XA.XIR[14].XIC_dummy_left.icell.Iout Iout 0.03553f
C2497 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.Ien 0.04854f
C2498 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PDM 0.04035f
C2499 XThR.Tn[11] XA.XIR[11].XIC[6].icell.Ien 0.14211f
C2500 XA.XIR[8].XIC[14].icell.Ien Vbias 0.19161f
C2501 XA.Cn[5] XThR.Tn[6] 0.40738f
C2502 XA.XIR[7].XIC[4].icell.PDM VPWR 0.01171f
C2503 XThR.XTB6.A XThR.XTB7.A 0.44014f
C2504 XA.XIR[12].XIC_dummy_left.icell.Iout XA.XIR[13].XIC_dummy_left.icell.Iout 0.03665f
C2505 XA.XIR[15].XIC[2].icell.PDM VPWR 0.01512f
C2506 XThR.Tn[0] XA.XIR[0].XIC[11].icell.Ien 0.14211f
C2507 XA.XIR[6].XIC[11].icell.PDM VPWR 0.01171f
C2508 XA.Cn[9] XA.XIR[6].XIC[9].icell.PDM 0.02601f
C2509 XA.Cn[14] XThR.Tn[9] 0.40742f
C2510 XA.Cn[12] XA.XIR[2].XIC[12].icell.PDM 0.02602f
C2511 XA.XIR[14].XIC[8].icell.PDM VPWR 0.01171f
C2512 XThR.Tn[6] XA.XIR[6].XIC[5].icell.Ien 0.14211f
C2513 XThR.XTB5.Y a_n997_1803# 0.06458f
C2514 XA.XIR[7].XIC[2].icell.Ien Iout 0.06801f
C2515 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.Ien 0.04854f
C2516 XA.XIR[5].XIC_15.icell.Ien Iout 0.0694f
C2517 XA.XIR[13].XIC_dummy_right.icell.Iout XA.XIR[14].XIC_dummy_right.icell.Iout 0.04047f
C2518 XA.Cn[1] XA.XIR[13].XIC[1].icell.PDM 0.02601f
C2519 XThR.Tn[7] XA.XIR[7].XIC[12].icell.Ien 0.14211f
C2520 XA.Cn[8] XThR.Tn[13] 0.40738f
C2521 XA.Cn[0] XA.XIR[12].XIC[0].icell.Ien 0.04604f
C2522 XA.XIR[9].XIC[0].icell.PDM VPWR 0.01171f
C2523 XA.Cn[10] XA.XIR[4].XIC[10].icell.Ien 0.04604f
C2524 XA.XIR[14].XIC[11].icell.Ien Vbias 0.19161f
C2525 XA.Cn[0] XThR.Tn[11] 0.4074f
C2526 thermo15c_0.XTB4.Y thermo15c_0.XTBN.Y 0.15636f
C2527 XA.XIR[5].XIC[2].icell.PDM Vbias 0.03928f
C2528 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2529 XA.XIR[6].XIC[1].icell.Ien Vbias 0.19161f
C2530 XA.Cn[6] XThR.Tn[1] 0.40744f
C2531 XA.XIR[11].XIC[12].icell.PDM VPWR 0.01171f
C2532 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.Ien 0.04854f
C2533 XA.XIR[12].XIC[1].icell.PDM Vbias 0.03928f
C2534 XThR.Tn[2] Vbias 1.39527f
C2535 XA.XIR[3].XIC[7].icell.Ien VPWR 0.18829f
C2536 XA.XIR[1].XIC[5].icell.PDM VPWR 0.01171f
C2537 XA.XIR[14].XIC[13].icell.PDM VPWR 0.01171f
C2538 XA.XIR[11].XIC[7].icell.PDM Vbias 0.03928f
C2539 XA.Cn[6] XThR.Tn[12] 0.40738f
C2540 XThR.Tn[9] Iout 1.12762f
C2541 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.Ien 0.04854f
C2542 XA.XIR[5].XIC_dummy_right.icell.Iout Iout 0.01732f
C2543 a_5155_9615# XA.Cn[4] 0.27224f
C2544 XA.Cn[12] XA.XIR[2].XIC[12].icell.Ien 0.04605f
C2545 XA.XIR[4].XIC[5].icell.PDM VPWR 0.01171f
C2546 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PDM 0.04035f
C2547 XA.XIR[1].XIC[2].icell.Ien VPWR 0.18829f
C2548 XA.XIR[3].XIC[13].icell.PDM VPWR 0.01171f
C2549 XA.XIR[8].XIC_15.icell.PDM VPWR 0.07527f
C2550 XA.XIR[6].XIC[6].icell.Ien Vbias 0.19161f
C2551 XA.Cn[5] XThR.Tn[4] 0.40738f
C2552 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PDM 0.04035f
C2553 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PDM 0.04035f
C2554 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.PDM 0.02104f
C2555 XA.XIR[8].XIC[10].icell.Ien VPWR 0.18829f
C2556 XA.XIR[15].XIC[0].icell.Ien Iout 0.07185f
C2557 XA.Cn[4] XThR.Tn[10] 0.40738f
C2558 XA.XIR[2].XIC[3].icell.PDM Vbias 0.03928f
C2559 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2560 XA.Cn[7] XA.XIR[3].XIC[7].icell.PDM 0.02601f
C2561 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2562 XA.XIR[13].XIC[2].icell.Ien Vbias 0.19161f
C2563 XA.Cn[12] XA.XIR[7].XIC[12].icell.PDM 0.02601f
C2564 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.PDM 0.02104f
C2565 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.PDM 0.02104f
C2566 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PDM 0.04035f
C2567 XThR.Tn[9] XA.XIR[9].XIC_15.icell.Ien 0.13564f
C2568 XA.XIR[0].XIC[12].icell.Ien VPWR 0.1902f
C2569 thermo15c_0.XTB7.B a_6243_9615# 0.01743f
C2570 XA.XIR[11].XIC[5].icell.Ien Vbias 0.19161f
C2571 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.PDM 0.02104f
C2572 XA.Cn[14] XA.XIR[12].XIC[14].icell.PDM 0.02601f
C2573 XA.XIR[15].XIC[5].icell.Ien Iout 0.07192f
C2574 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.PDM 0.02104f
C2575 XA.XIR[10].XIC[7].icell.Ien Vbias 0.19161f
C2576 a_7651_9569# XA.Cn[8] 0.1927f
C2577 thermo15c_0.XTBN.A XA.Cn[8] 0.13691f
C2578 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PDM 0.04039f
C2579 XA.XIR[2].XIC_15.icell.PUM VPWR 0.01655f
C2580 XA.XIR[7].XIC_15.icell.Ien VPWR 0.26829f
C2581 XA.XIR[4].XIC[8].icell.Ien Iout 0.06801f
C2582 XThR.Tn[13] XA.XIR[13].XIC[5].icell.Ien 0.14211f
C2583 XA.XIR[5].XIC[0].icell.Ien VPWR 0.18829f
C2584 XThR.XTB5.A XThR.XTB2.Y 0.02203f
C2585 XThR.XTB7.B XThR.XTB6.A 1.47641f
C2586 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.PDM 0.02104f
C2587 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.Ien 0.04854f
C2588 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.PDM 0.02104f
C2589 XA.XIR[4].XIC_dummy_left.icell.Iout VPWR 0.10954f
C2590 XA.XIR[8].XIC[2].icell.Ien Iout 0.06801f
C2591 XA.XIR[2].XIC[9].icell.Ien Vbias 0.19161f
C2592 XA.Cn[4] XA.XIR[1].XIC[4].icell.PDM 0.02602f
C2593 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.PDM 0.02104f
C2594 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout 0.06446f
C2595 XA.Cn[13] VPWR 4.60106f
C2596 XA.XIR[1].XIC[11].icell.Ien Vbias 0.19173f
C2597 thermo15c_0.XTBN.Y XA.Cn[4] 0.49752f
C2598 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.Ien 0.04854f
C2599 XThR.Tn[8] XThR.Tn[9] 0.10569f
C2600 XA.XIR[9].XIC[11].icell.Ien Iout 0.06801f
C2601 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2602 XA.Cn[4] XA.XIR[4].XIC[4].icell.PDM 0.02601f
C2603 XA.XIR[6].XIC[2].icell.Ien VPWR 0.18829f
C2604 XA.Cn[1] XA.XIR[9].XIC[1].icell.Ien 0.04604f
C2605 XA.Cn[2] Iout 0.22439f
C2606 XA.XIR[0].XIC[4].icell.Ien Iout 0.0675f
C2607 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Ien 0.01546f
C2608 XA.XIR[7].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2609 XA.XIR[10].XIC_dummy_left.icell.Ien XThR.Tn[10] 0.01244f
C2610 XA.XIR[11].XIC[11].icell.PDM VPWR 0.01171f
C2611 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Ien 0.01597f
C2612 XA.Cn[3] XA.XIR[10].XIC[3].icell.Ien 0.04604f
C2613 XA.Cn[0] XThR.Tn[14] 0.40739f
C2614 XA.Cn[0] XA.XIR[11].XIC[0].icell.PDM 0.02601f
C2615 XThR.Tn[6] XA.XIR[6].XIC[10].icell.Ien 0.14211f
C2616 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.PDM 0.02104f
C2617 XA.XIR[7].XIC[7].icell.Ien Iout 0.06801f
C2618 XA.XIR[7].XIC[3].icell.PDM Vbias 0.03928f
C2619 XThR.Tn[10] Vbias 1.39532f
C2620 XA.XIR[14].XIC[12].icell.PDM VPWR 0.01171f
C2621 XA.XIR[9].XIC_15.icell.PDM VPWR 0.07527f
C2622 XA.XIR[15].XIC[1].icell.PDM Vbias 0.03928f
C2623 XA.XIR[6].XIC[10].icell.PDM Vbias 0.03928f
C2624 XA.XIR[0].XIC[7].icell.PDM VPWR 0.01132f
C2625 XA.Cn[10] XA.XIR[3].XIC[10].icell.PDM 0.02601f
C2626 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.Ien 0.04854f
C2627 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.Ien 0.04854f
C2628 XA.XIR[14].XIC[7].icell.PDM Vbias 0.03928f
C2629 XA.XIR[10].XIC[3].icell.Ien VPWR 0.18829f
C2630 XA.Cn[9] XA.XIR[9].XIC[9].icell.Ien 0.04604f
C2631 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.PDM 0.02104f
C2632 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.Ien 0.04854f
C2633 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.PDM 0.02104f
C2634 thermo15c_0.XTB3.Y thermo15c_0.XTB6.Y 0.04428f
C2635 XA.Cn[12] Vbias 0.8219f
C2636 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PDM 0.04035f
C2637 thermo15c_0.XTB7.A thermo15c_0.XTB7.Y 0.37429f
C2638 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PDM 0.04056f
C2639 thermo15c_0.XTB4.Y thermo15c_0.XTBN.A 0.03415f
C2640 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PDM 0.04035f
C2641 thermo15c_0.XTB2.Y a_7875_9569# 0.06476f
C2642 XA.XIR[3].XIC[12].icell.Ien VPWR 0.18829f
C2643 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.PDM 0.02104f
C2644 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.Ien 0.04854f
C2645 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.Ien 0.04854f
C2646 XA.XIR[2].XIC[5].icell.Ien VPWR 0.18829f
C2647 XA.XIR[1].XIC[7].icell.Ien VPWR 0.18829f
C2648 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.PDM 0.02104f
C2649 XThR.Tn[8] XA.XIR[8].XIC[2].icell.Ien 0.14211f
C2650 XA.XIR[1].XIC[4].icell.PDM Vbias 0.03928f
C2651 XA.Cn[4] XThR.Tn[13] 0.40738f
C2652 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.Ien 0.04854f
C2653 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.03838f
C2654 XA.XIR[6].XIC[11].icell.Ien Vbias 0.19161f
C2655 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.Ien 0.04854f
C2656 thermo15c_0.XTBN.Y Vbias 0.22975f
C2657 XA.XIR[4].XIC[4].icell.PDM Vbias 0.03928f
C2658 XA.XIR[8].XIC_15.icell.Ien VPWR 0.26829f
C2659 XThR.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.14211f
C2660 XThR.XTB7.A a_n1049_5317# 0.02018f
C2661 XA.XIR[3].XIC[12].icell.PDM Vbias 0.03928f
C2662 XA.XIR[8].XIC[14].icell.PDM Vbias 0.03928f
C2663 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.PDM 0.02104f
C2664 XA.XIR[14].XIC[5].icell.Ien Vbias 0.19161f
C2665 XA.Cn[4] XA.XIR[5].XIC[4].icell.Ien 0.04604f
C2666 XA.Cn[14] XA.XIR[15].XIC[14].icell.PDM 0.02601f
C2667 XThR.XTBN.Y XThR.XTB6.A 0.03867f
C2668 XA.Cn[1] XThR.Tn[9] 0.40738f
C2669 XA.XIR[13].XIC[7].icell.Ien Vbias 0.19161f
C2670 XA.Cn[2] XThR.Tn[8] 0.40738f
C2671 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.PDM 0.02104f
C2672 XA.XIR[10].XIC[13].icell.Ien Iout 0.06801f
C2673 XA.XIR[3].XIC[4].icell.Ien Iout 0.06801f
C2674 XThR.XTB2.Y XThR.Tn[9] 0.292f
C2675 a_n997_3755# XThR.Tn[9] 0.19352f
C2676 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PDM 0.04035f
C2677 XThR.Tn[14] XA.XIR[14].XIC[6].icell.Ien 0.14211f
C2678 XA.Cn[6] XA.XIR[0].XIC[6].icell.Ien 0.04659f
C2679 XThR.Tn[1] XA.XIR[1].XIC[6].icell.Ien 0.14211f
C2680 XA.XIR[5].XIC[5].icell.PDM VPWR 0.01171f
C2681 XThR.XTBN.Y XThR.Tn[0] 0.55717f
C2682 XA.XIR[8].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2683 XA.XIR[4].XIC[13].icell.Ien Iout 0.06801f
C2684 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.PDM 0.02104f
C2685 XThR.XTB6.A XThR.XTB4.Y 0.04137f
C2686 XA.XIR[12].XIC[4].icell.PDM VPWR 0.01171f
C2687 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.Ien 0.04854f
C2688 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.Ien 0.04854f
C2689 XA.XIR[8].XIC[7].icell.Ien Iout 0.06801f
C2690 XA.XIR[11].XIC[10].icell.PDM VPWR 0.01171f
C2691 XA.Cn[8] XThR.Tn[7] 0.40738f
C2692 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.Ien 0.04854f
C2693 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.PDM 0.02104f
C2694 XA.XIR[2].XIC[14].icell.Ien Vbias 0.19161f
C2695 XA.Cn[11] XA.XIR[8].XIC[11].icell.PDM 0.02601f
C2696 XA.XIR[14].XIC[11].icell.PDM VPWR 0.01171f
C2697 XA.Cn[3] XA.XIR[13].XIC[3].icell.Ien 0.04604f
C2698 XA.XIR[14].XIC[0].icell.Ien Vbias 0.19149f
C2699 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PDM 0.04035f
C2700 XA.Cn[0] XA.XIR[14].XIC[0].icell.PDM 0.02601f
C2701 XA.XIR[6].XIC[7].icell.Ien VPWR 0.18829f
C2702 XThR.Tn[13] Vbias 1.39532f
C2703 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.Ien 0.04854f
C2704 XThR.XTB7.A a_n1049_6405# 0.02287f
C2705 XA.XIR[0].XIC[9].icell.Ien Iout 0.0675f
C2706 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.PDM 0.02104f
C2707 XA.XIR[3].XIC[0].icell.PDM VPWR 0.01171f
C2708 XA.XIR[8].XIC[2].icell.PDM VPWR 0.01171f
C2709 XA.XIR[4].XIC_dummy_left.icell.Iout XA.XIR[5].XIC_dummy_left.icell.Iout 0.03665f
C2710 XThR.Tn[6] XA.XIR[6].XIC_15.icell.Ien 0.13564f
C2711 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.PDM 0.02104f
C2712 XA.XIR[2].XIC[6].icell.PDM VPWR 0.01171f
C2713 XThR.Tn[1] XThR.Tn[2] 0.15279f
C2714 XA.XIR[13].XIC[3].icell.Ien VPWR 0.18829f
C2715 XA.XIR[7].XIC[12].icell.Ien Iout 0.06801f
C2716 XA.XIR[5].XIC[4].icell.Ien Vbias 0.19161f
C2717 XThR.XTB1.Y a_n997_3979# 0.06353f
C2718 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.PDM 0.02104f
C2719 XA.Cn[12] XThR.Tn[0] 0.40763f
C2720 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.Ien 0.04854f
C2721 XA.XIR[11].XIC[6].icell.Ien VPWR 0.18829f
C2722 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR 0.38914f
C2723 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PDM 0.04035f
C2724 XA.XIR[10].XIC[11].icell.Ien Iout 0.06801f
C2725 XA.XIR[3].XIC[1].icell.Ien Iout 0.06801f
C2726 thermo15c_0.XTBN.Y a_2979_9615# 0.0607f
C2727 XA.XIR[10].XIC[8].icell.Ien VPWR 0.18829f
C2728 XA.Cn[1] XA.Cn[2] 0.71417f
C2729 XA.XIR[9].XIC[14].icell.PDM Vbias 0.03928f
C2730 thermo15c_0.XTB7.Y XA.Cn[13] 0.10846f
C2731 XA.Cn[4] XA.XIR[5].XIC[4].icell.PDM 0.02601f
C2732 XA.XIR[0].XIC[6].icell.PDM Vbias 0.03945f
C2733 thermo15c_0.XTB7.B a_8739_9569# 0.0168f
C2734 XThR.XTB7.B a_n1049_5317# 0.01743f
C2735 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PDM 0.04035f
C2736 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.PDM 0.02104f
C2737 XA.XIR[9].XIC_dummy_left.icell.Iout Iout 0.03553f
C2738 XA.Cn[6] XA.XIR[3].XIC[6].icell.Ien 0.04604f
C2739 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.Ien 0.04854f
C2740 XThR.Tn[11] XA.XIR[11].XIC_dummy_left.icell.Iout 0.03385f
C2741 XThR.Tn[5] XA.XIR[5].XIC[1].icell.Ien 0.14211f
C2742 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PDM 0.04035f
C2743 XA.XIR[2].XIC[10].icell.Ien VPWR 0.18829f
C2744 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.PDM 0.02104f
C2745 XA.Cn[0] VPWR 3.67891f
C2746 XA.XIR[1].XIC[12].icell.Ien VPWR 0.18829f
C2747 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.Ien 0.04854f
C2748 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PDM 0.04035f
C2749 XThR.Tn[8] XA.XIR[8].XIC[7].icell.Ien 0.14211f
C2750 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.Ien 0.04854f
C2751 XA.Cn[5] XA.XIR[0].XIC[5].icell.PDM 0.02803f
C2752 XA.XIR[13].XIC[13].icell.Ien Iout 0.06801f
C2753 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.PDM 0.02104f
C2754 XA.Cn[10] XThR.Tn[2] 0.40741f
C2755 thermo15c_0.XTBN.A Vbias 0.01693f
C2756 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.PDM 0.02104f
C2757 XA.Cn[11] XA.XIR[10].XIC[11].icell.PDM 0.02601f
C2758 XThR.XTB3.Y data[4] 0.03253f
C2759 XThR.Tn[5] XA.XIR[5].XIC[6].icell.Ien 0.14211f
C2760 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PDM 0.04035f
C2761 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2762 XA.Cn[2] XA.XIR[10].XIC[2].icell.PDM 0.02601f
C2763 XThR.XTB6.Y XThR.XTBN.A 0.06405f
C2764 XA.Cn[12] XA.XIR[5].XIC[12].icell.Ien 0.04604f
C2765 XA.XIR[7].XIC[6].icell.PDM VPWR 0.01171f
C2766 XThR.XTBN.Y XThR.Tn[1] 0.61094f
C2767 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.PDM 0.02104f
C2768 XA.Cn[11] XA.XIR[9].XIC[11].icell.PDM 0.02601f
C2769 XA.XIR[6].XIC[13].icell.PDM VPWR 0.01171f
C2770 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.Ien 0.04854f
C2771 XA.XIR[15].XIC[4].icell.PDM VPWR 0.01512f
C2772 XA.XIR[3].XIC[9].icell.Ien Iout 0.06801f
C2773 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.Ien 0.04854f
C2774 thermo15c_0.XTB3.Y XA.Cn[2] 0.18399f
C2775 XA.Cn[5] XA.XIR[7].XIC[5].icell.Ien 0.04604f
C2776 XThR.XTBN.Y XThR.Tn[12] 0.50762f
C2777 XThR.Tn[1] XA.XIR[1].XIC[11].icell.Ien 0.14211f
C2778 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.PDM 0.02104f
C2779 XA.XIR[14].XIC[10].icell.PDM VPWR 0.01171f
C2780 XA.Cn[4] XA.XIR[12].XIC[4].icell.Ien 0.04604f
C2781 XA.XIR[2].XIC[2].icell.Ien Iout 0.06801f
C2782 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.PDM 0.02104f
C2783 XA.Cn[14] XA.XIR[0].XIC[14].icell.Ien 0.04662f
C2784 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.PDM 0.02104f
C2785 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.PDM 0.02104f
C2786 XA.XIR[1].XIC[4].icell.Ien Iout 0.06801f
C2787 XA.XIR[13].XIC_dummy_left.icell.Ien XThR.Tn[13] 0.01244f
C2788 XA.XIR[9].XIC[2].icell.PDM VPWR 0.01171f
C2789 XA.Cn[11] XThR.Tn[6] 0.40738f
C2790 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.Ien 0.04854f
C2791 XA.XIR[5].XIC[4].icell.PDM Vbias 0.03928f
C2792 XA.Cn[7] XA.XIR[6].XIC[7].icell.PDM 0.02601f
C2793 XA.XIR[8].XIC[12].icell.Ien Iout 0.06801f
C2794 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2795 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.PDM 0.02104f
C2796 XA.XIR[12].XIC[13].icell.Ien VPWR 0.18829f
C2797 thermo15c_0.XTB5.Y thermo15c_0.XTB7.B 0.30234f
C2798 XA.Cn[2] XA.XIR[11].XIC[2].icell.Ien 0.04604f
C2799 XA.XIR[12].XIC[3].icell.PDM Vbias 0.03928f
C2800 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PDM 0.04035f
C2801 XThR.XTB7.Y XThR.Tn[9] 0.07413f
C2802 XA.XIR[1].XIC[7].icell.PDM VPWR 0.01171f
C2803 XA.XIR[6].XIC[12].icell.Ien VPWR 0.18829f
C2804 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Iout 0.01728f
C2805 XA.XIR[11].XIC[9].icell.PDM Vbias 0.03928f
C2806 XA.XIR[4].XIC[7].icell.PDM VPWR 0.01171f
C2807 XA.XIR[0].XIC[14].icell.Ien Iout 0.0675f
C2808 XA.XIR[5].XIC_15.icell.PUM VPWR 0.01655f
C2809 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.PDM 0.02104f
C2810 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PDM 0.04035f
C2811 XA.XIR[3].XIC_15.icell.PDM VPWR 0.07527f
C2812 XA.XIR[14].XIC[6].icell.Ien VPWR 0.18883f
C2813 XA.Cn[12] XThR.Tn[1] 0.40744f
C2814 XA.XIR[13].XIC[11].icell.Ien Iout 0.06801f
C2815 XA.Cn[8] XA.XIR[0].XIC[8].icell.PDM 0.02805f
C2816 XThR.XTBN.Y a_n1049_5317# 0.07731f
C2817 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PDM 0.04035f
C2818 XA.XIR[13].XIC[8].icell.Ien VPWR 0.18829f
C2819 XA.XIR[5].XIC[9].icell.Ien Vbias 0.19161f
C2820 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout 0.06446f
C2821 XA.Cn[4] XThR.Tn[7] 0.40738f
C2822 XA.Cn[12] XThR.Tn[12] 0.40738f
C2823 XA.XIR[8].XIC[1].icell.PDM Vbias 0.03928f
C2824 VPWR data[4] 0.5303f
C2825 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.Ien 0.04854f
C2826 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.PDM 0.02104f
C2827 XA.XIR[2].XIC[5].icell.PDM Vbias 0.03928f
C2828 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.01728f
C2829 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.Ien 0.04854f
C2830 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PDM 0.04035f
C2831 XA.XIR[12].XIC[4].icell.Ien Vbias 0.19161f
C2832 XA.Cn[11] XThR.Tn[4] 0.40738f
C2833 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.Ien 0.04854f
C2834 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.Ien 0.04854f
C2835 XA.XIR[6].XIC[4].icell.Ien Iout 0.06801f
C2836 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2837 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PDM 0.04035f
C2838 XA.Cn[10] XThR.Tn[10] 0.40738f
C2839 XA.XIR[2].XIC_15.icell.Ien VPWR 0.26829f
C2840 XA.XIR[12].XIC[11].icell.Ien VPWR 0.18829f
C2841 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.Ien 0.04854f
C2842 XA.Cn[14] XA.XIR[3].XIC[14].icell.Ien 0.04604f
C2843 XA.Cn[5] XA.XIR[8].XIC[5].icell.Ien 0.04604f
C2844 XA.Cn[10] XA.XIR[6].XIC[10].icell.PDM 0.02601f
C2845 XA.Cn[13] XA.XIR[2].XIC[13].icell.PDM 0.02602f
C2846 XThR.Tn[8] XA.XIR[8].XIC[12].icell.Ien 0.14211f
C2847 XA.Cn[11] XA.XIR[13].XIC[11].icell.PDM 0.02601f
C2848 XA.Cn[2] XA.XIR[13].XIC[2].icell.PDM 0.02601f
C2849 XA.Cn[6] XA.XIR[1].XIC[6].icell.Ien 0.04606f
C2850 thermo15c_0.XTB1.Y thermo15c_0.XTB2.Y 2.14864f
C2851 thermo15c_0.XTB5.A thermo15c_0.XTB6.A 1.80461f
C2852 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.Ien 0.04854f
C2853 XA.Cn[1] XA.XIR[3].XIC[1].icell.Ien 0.04604f
C2854 XA.Cn[2] XThR.Tn[3] 0.40738f
C2855 XA.XIR[10].XIC[1].icell.PDM VPWR 0.01171f
C2856 XA.XIR[11].XIC[3].icell.Ien Iout 0.06801f
C2857 a_6243_9615# Vbias 0.01011f
C2858 XThR.XTBN.Y a_n1049_6405# 0.07602f
C2859 XThR.Tn[12] a_n997_1803# 0.18719f
C2860 XA.XIR[10].XIC[5].icell.Ien Iout 0.06801f
C2861 XThR.Tn[5] XA.XIR[5].XIC[11].icell.Ien 0.14211f
C2862 XA.Cn[3] XThR.Tn[5] 0.40738f
C2863 thermo15c_0.XTB1.Y VPWR 1.11809f
C2864 XA.XIR[5].XIC[5].icell.Ien VPWR 0.18829f
C2865 XA.XIR[2].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2866 XA.XIR[3].XIC[14].icell.Ien Iout 0.06801f
C2867 XThR.Tn[7] Vbias 1.39526f
C2868 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.Ien 0.04854f
C2869 XA.XIR[2].XIC[7].icell.Ien Iout 0.06801f
C2870 XA.Cn[13] XA.XIR[7].XIC[13].icell.Ien 0.04604f
C2871 a_5949_9615# XA.Cn[5] 0.26251f
C2872 thermo15c_0.XTBN.Y XA.Cn[10] 0.4511f
C2873 XA.XIR[7].XIC[5].icell.PDM Vbias 0.03928f
C2874 XThR.XTB4.Y a_n1049_6405# 0.01546f
C2875 XA.Cn[2] XA.XIR[14].XIC[2].icell.Ien 0.04604f
C2876 XA.XIR[1].XIC[9].icell.Ien Iout 0.06801f
C2877 XThR.Tn[5] VPWR 8.03417f
C2878 XA.XIR[15].XIC[3].icell.PDM Vbias 0.03928f
C2879 XA.XIR[6].XIC[12].icell.PDM Vbias 0.03928f
C2880 XA.XIR[4].XIC[2].icell.Ien Vbias 0.19161f
C2881 XThR.Tn[2] XA.XIR[2].XIC[0].icell.Ien 0.14251f
C2882 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.Ien 0.04854f
C2883 VPWR bias[1] 1.33312f
C2884 XA.Cn[8] Iout 0.22393f
C2885 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.PDM 0.02104f
C2886 XA.XIR[0].XIC[9].icell.PDM VPWR 0.01451f
C2887 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.PDM 0.02104f
C2888 XA.XIR[14].XIC[9].icell.PDM Vbias 0.03928f
C2889 thermo15c_0.XTB7.A XA.Cn[5] 0.02777f
C2890 XThR.Tn[12] XThR.Tn[13] 0.11103f
C2891 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.Ien 0.04854f
C2892 XA.Cn[6] XThR.Tn[2] 0.40741f
C2893 thermo15c_0.XTB5.Y XA.Cn[8] 0.0173f
C2894 XA.XIR[9].XIC[1].icell.PDM Vbias 0.03928f
C2895 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PDM 0.04035f
C2896 thermo15c_0.XTB6.A thermo15c_0.XTBN.Y 0.03867f
C2897 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.Ien 0.04854f
C2898 XA.Cn[0] XA.XIR[0].XIC[0].icell.Ien 0.04657f
C2899 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PDM 0.04035f
C2900 XA.XIR[9].XIC[5].icell.Ien Vbias 0.19161f
C2901 XA.Cn[13] XA.XIR[7].XIC[13].icell.PDM 0.02601f
C2902 XA.Cn[6] XA.XIR[6].XIC[6].icell.Ien 0.04604f
C2903 XA.XIR[1].XIC[6].icell.PDM Vbias 0.03928f
C2904 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR 0.38998f
C2905 XA.Cn[7] XThR.Tn[6] 0.40738f
C2906 a_7875_9569# XA.Cn[9] 0.19271f
C2907 XA.XIR[5].XIC[14].icell.Ien Vbias 0.19161f
C2908 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Iout 0.03842f
C2909 XThR.Tn[14] XA.XIR[14].XIC_dummy_left.icell.Iout 0.03385f
C2910 XA.XIR[4].XIC[6].icell.PDM Vbias 0.03928f
C2911 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.Ien 0.04854f
C2912 XThR.Tn[3] XA.XIR[3].XIC[4].icell.Ien 0.14211f
C2913 XA.XIR[3].XIC[14].icell.PDM Vbias 0.03928f
C2914 XA.Cn[4] XA.XIR[15].XIC[4].icell.Ien 0.04292f
C2915 XA.Cn[8] XA.XIR[0].XIC[8].icell.Ien 0.04654f
C2916 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout 0.06446f
C2917 XA.Cn[10] XThR.Tn[13] 0.40738f
C2918 XA.Cn[5] XA.XIR[1].XIC[5].icell.PDM 0.02602f
C2919 XA.XIR[12].XIC[9].icell.Ien Vbias 0.19161f
C2920 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PDM 0.04056f
C2921 XA.XIR[6].XIC[0].icell.PDM VPWR 0.01171f
C2922 XA.Cn[2] XThR.Tn[11] 0.40738f
C2923 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PDM 0.04035f
C2924 XA.XIR[6].XIC[9].icell.Ien Iout 0.06801f
C2925 XA.Cn[5] XA.XIR[4].XIC[5].icell.PDM 0.02601f
C2926 XA.XIR[15].XIC[13].icell.Ien VPWR 0.31713f
C2927 XA.XIR[5].XIC[7].icell.PDM VPWR 0.01171f
C2928 XA.XIR[9].XIC[0].icell.Ien Vbias 0.19149f
C2929 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.Ien 0.04854f
C2930 XA.XIR[13].XIC[1].icell.PDM VPWR 0.01171f
C2931 XA.XIR[14].XIC[3].icell.Ien Iout 0.06801f
C2932 XThR.XTB7.B XThR.XTB7.A 0.35833f
C2933 XA.Cn[8] XThR.Tn[8] 0.40738f
C2934 XThR.XTB5.A XThR.XTB3.Y 0.01152f
C2935 XA.XIR[12].XIC[6].icell.PDM VPWR 0.01171f
C2936 XA.XIR[13].XIC[5].icell.Ien Iout 0.06801f
C2937 XA.Cn[1] XA.XIR[11].XIC[1].icell.PDM 0.02601f
C2938 thermo15c_0.XTB4.Y thermo15c_0.XTB5.Y 2.06459f
C2939 thermo15c_0.XTB3.Y thermo15c_0.XTB7.B 0.23315f
C2940 XA.Cn[13] XA.XIR[8].XIC[13].icell.Ien 0.04604f
C2941 XA.Cn[0] XA.XIR[10].XIC[0].icell.Ien 0.04604f
C2942 XA.Cn[14] XA.XIR[1].XIC[14].icell.Ien 0.04606f
C2943 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout 0.06446f
C2944 XA.XIR[11].XIC[8].icell.Ien Iout 0.06801f
C2945 XA.Cn[11] XA.XIR[3].XIC[11].icell.PDM 0.02601f
C2946 XA.Cn[7] XThR.Tn[4] 0.40738f
C2947 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PDM 0.04035f
C2948 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.Ien 0.04854f
C2949 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.PDM 0.02104f
C2950 XA.XIR[11].XIC_dummy_left.icell.Iout VPWR 0.10954f
C2951 XA.XIR[10].XIC[0].icell.PDM Vbias 0.03915f
C2952 XA.XIR[5].XIC[10].icell.Ien VPWR 0.18829f
C2953 XThR.XTB5.Y XThR.Tn[8] 0.01728f
C2954 XThR.XTB7.A XThR.Tn[2] 0.12549f
C2955 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.Ien 0.04854f
C2956 XA.XIR[8].XIC[4].icell.PDM VPWR 0.01171f
C2957 XThR.Tn[4] XA.XIR[4].XIC[1].icell.Ien 0.14211f
C2958 XA.Cn[6] XThR.Tn[10] 0.40738f
C2959 XA.XIR[3].XIC[2].icell.PDM VPWR 0.01171f
C2960 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10] 0.14211f
C2961 XThR.Tn[3] XA.XIR[3].XIC[1].icell.Ien 0.14211f
C2962 XA.XIR[2].XIC[8].icell.PDM VPWR 0.01171f
C2963 XA.XIR[15].XIC[4].icell.Ien Vbias 0.15966f
C2964 XA.XIR[2].XIC[12].icell.Ien Iout 0.06801f
C2965 XA.XIR[12].XIC[5].icell.Ien VPWR 0.18829f
C2966 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.Ien 0.04854f
C2967 XA.XIR[1].XIC[14].icell.Ien Iout 0.06801f
C2968 XA.XIR[4].XIC[7].icell.Ien Vbias 0.19161f
C2969 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.Ien 0.04854f
C2970 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PDM 0.04035f
C2971 XA.Cn[8] XA.XIR[3].XIC[8].icell.Ien 0.04604f
C2972 thermo15c_0.XTBN.A XA.Cn[10] 0.12208f
C2973 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2974 XA.Cn[8] XA.XIR[1].XIC[8].icell.PDM 0.02602f
C2975 thermo15c_0.XTBN.Y a_4067_9615# 0.08456f
C2976 XA.XIR[3].XIC_dummy_left.icell.Iout Iout 0.03553f
C2977 XA.XIR[15].XIC[11].icell.Ien VPWR 0.31713f
C2978 XThR.Tn[4] XA.XIR[4].XIC[6].icell.Ien 0.14211f
C2979 XA.XIR[12].XIC[1].icell.Ien Iout 0.06801f
C2980 XA.Cn[8] XA.XIR[4].XIC[8].icell.PDM 0.02601f
C2981 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.Ien 0.04854f
C2982 XA.XIR[7].XIC[1].icell.Ien Vbias 0.19161f
C2983 XA.XIR[0].XIC[8].icell.PDM Vbias 0.03945f
C2984 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PDM 0.04035f
C2985 XA.XIR[5].XIC[2].icell.Ien Iout 0.06801f
C2986 XA.XIR[9].XIC[10].icell.Ien Vbias 0.19161f
C2987 thermo15c_0.XTB1.Y thermo15c_0.XTB7.Y 0.05222f
C2988 thermo15c_0.XTB2.Y thermo15c_0.XTB6.Y 0.04959f
C2989 XA.XIR[8].XIC_dummy_left.icell.Iout XA.XIR[9].XIC_dummy_left.icell.Iout 0.03665f
C2990 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout 0.06446f
C2991 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PDM 0.04035f
C2992 thermo15c_0.XTB6.A thermo15c_0.XTBN.A 0.0513f
C2993 XThR.XTB5.A VPWR 0.83125f
C2994 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Iout 0.03935f
C2995 XA.XIR[12].XIC[14].icell.Ien Vbias 0.19161f
C2996 XA.XIR[0].XIC[3].icell.Ien Vbias 0.19213f
C2997 thermo15c_0.XTBN.Y XA.Cn[6] 0.49549f
C2998 XA.Cn[14] XA.XIR[6].XIC[14].icell.Ien 0.04604f
C2999 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PDM 0.04035f
C3000 XThR.XTB1.Y XThR.Tn[8] 0.29191f
C3001 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PDM 0.0404f
C3002 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3003 XA.Cn[13] XA.XIR[10].XIC[13].icell.PDM 0.02601f
C3004 XA.Cn[4] Iout 0.22518f
C3005 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.PDM 0.02104f
C3006 thermo15c_0.XTB6.Y VPWR 1.03165f
C3007 XA.XIR[7].XIC[6].icell.Ien Vbias 0.19161f
C3008 XThR.Tn[12] XA.XIR[12].XIC[4].icell.Ien 0.14211f
C3009 XA.Cn[3] XA.XIR[4].XIC[3].icell.Ien 0.04604f
C3010 XThR.Tn[3] XA.XIR[3].XIC[9].icell.Ien 0.14211f
C3011 XA.Cn[2] XThR.Tn[14] 0.40738f
C3012 thermo15c_0.XTB5.Y XA.Cn[4] 0.20108f
C3013 XThR.XTBN.Y XThR.XTB7.A 0.59539f
C3014 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.Ien 0.04854f
C3015 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3016 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PDM 0.04035f
C3017 XA.XIR[7].XIC[8].icell.PDM VPWR 0.01171f
C3018 XA.XIR[9].XIC[1].icell.Ien VPWR 0.18829f
C3019 XThR.Tn[2] XA.XIR[2].XIC[4].icell.Ien 0.14211f
C3020 XA.Cn[12] XA.XIR[8].XIC[12].icell.PDM 0.02601f
C3021 XA.XIR[6].XIC_15.icell.PDM VPWR 0.07527f
C3022 XA.XIR[15].XIC[6].icell.PDM VPWR 0.01512f
C3023 XA.XIR[4].XIC[3].icell.Ien VPWR 0.18829f
C3024 XA.Cn[5] XA.XIR[2].XIC[5].icell.Ien 0.04605f
C3025 XA.Cn[1] XA.XIR[14].XIC[1].icell.PDM 0.02601f
C3026 XA.XIR[6].XIC[14].icell.Ien Iout 0.06801f
C3027 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout 0.06446f
C3028 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.PDM 0.02104f
C3029 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.Ien 0.04854f
C3030 XA.Cn[0] XA.XIR[13].XIC[0].icell.Ien 0.04604f
C3031 XA.Cn[14] Vbias 0.8291f
C3032 XThR.XTB2.Y XThR.XTB5.Y 0.0451f
C3033 XThR.XTB7.A XThR.XTB4.Y 0.14536f
C3034 XA.XIR[14].XIC[8].icell.Ien Iout 0.06801f
C3035 XA.XIR[9].XIC[4].icell.PDM VPWR 0.01171f
C3036 XA.XIR[5].XIC[6].icell.PDM Vbias 0.03928f
C3037 XA.XIR[9].XIC[6].icell.Ien VPWR 0.18829f
C3038 XA.XIR[14].XIC_dummy_left.icell.Iout VPWR 0.10954f
C3039 XA.XIR[13].XIC[0].icell.PDM Vbias 0.03915f
C3040 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.Ien 0.04854f
C3041 XThR.Tn[9] XA.XIR[9].XIC[2].icell.Ien 0.14211f
C3042 XA.XIR[12].XIC[5].icell.PDM Vbias 0.03928f
C3043 XA.Cn[6] XThR.Tn[13] 0.40738f
C3044 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PDM 0.04035f
C3045 XA.XIR[12].XIC[12].icell.Ien Vbias 0.19161f
C3046 XA.XIR[1].XIC[9].icell.PDM VPWR 0.01171f
C3047 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.Ien 0.04854f
C3048 XA.XIR[5].XIC_15.icell.Ien VPWR 0.26829f
C3049 XA.XIR[4].XIC[9].icell.PDM VPWR 0.01171f
C3050 XA.XIR[7].XIC[2].icell.Ien VPWR 0.18829f
C3051 XA.Cn[5] XA.XIR[5].XIC[5].icell.PDM 0.02601f
C3052 Vbias Iout 74.00211f
C3053 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PDM 0.04035f
C3054 XA.XIR[8].XIC[1].icell.Ien Vbias 0.19161f
C3055 XA.XIR[3].XIC[3].icell.Ien Vbias 0.19161f
C3056 XA.Cn[3] XThR.Tn[9] 0.40738f
C3057 XA.Cn[4] XThR.Tn[8] 0.40738f
C3058 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.Ien 0.04854f
C3059 XA.XIR[12].XIC_15.icell.PDM VPWR 0.07527f
C3060 thermo15c_0.XTB5.Y Vbias 0.01606f
C3061 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3062 XA.XIR[15].XIC[9].icell.Ien Vbias 0.15966f
C3063 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.04035f
C3064 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.PDM 0.02104f
C3065 XA.XIR[4].XIC[12].icell.Ien Vbias 0.19161f
C3066 XA.XIR[8].XIC[3].icell.PDM Vbias 0.03928f
C3067 XA.XIR[3].XIC[1].icell.PDM Vbias 0.03928f
C3068 XThR.XTB1.Y XThR.XTB2.Y 2.14864f
C3069 XThR.XTB6.A data[5] 0.37233f
C3070 XA.XIR[2].XIC[7].icell.PDM Vbias 0.03928f
C3071 XA.Cn[6] XA.XIR[0].XIC[6].icell.PDM 0.02803f
C3072 XA.XIR[8].XIC[6].icell.Ien Vbias 0.19161f
C3073 XThR.Tn[9] VPWR 8.97014f
C3074 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PDM 0.04035f
C3075 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.PDM 0.02104f
C3076 XA.XIR[5].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3077 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.PDM 0.02104f
C3078 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.04035f
C3079 XThR.Tn[4] XA.XIR[4].XIC[11].icell.Ien 0.14211f
C3080 XThR.Tn[0] XA.XIR[0].XIC[3].icell.Ien 0.14211f
C3081 XThR.Tn[10] XA.XIR[10].XIC[2].icell.Ien 0.14211f
C3082 XA.Cn[10] XThR.Tn[7] 0.40738f
C3083 XA.Cn[8] XA.XIR[1].XIC[8].icell.Ien 0.04606f
C3084 XA.Cn[13] XA.XIR[13].XIC[13].icell.PDM 0.02601f
C3085 XA.XIR[5].XIC[7].icell.Ien Iout 0.06801f
C3086 XA.Cn[3] XA.XIR[10].XIC[3].icell.PDM 0.02601f
C3087 XA.XIR[9].XIC_15.icell.Ien Vbias 0.19195f
C3088 XThR.XTB7.B XThR.XTBN.Y 0.3875f
C3089 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PDM 0.04035f
C3090 XThR.Tn[7] XA.XIR[7].XIC[4].icell.Ien 0.14211f
C3091 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.04056f
C3092 XA.Cn[12] XA.XIR[9].XIC[12].icell.PDM 0.02601f
C3093 XA.XIR[0].XIC[8].icell.Ien Vbias 0.19213f
C3094 XA.XIR[15].XIC[0].icell.Ien VPWR 0.31713f
C3095 thermo15c_0.XTB3.Y thermo15c_0.XTB4.Y 2.13136f
C3096 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.PDM 0.02104f
C3097 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.Ien 0.04854f
C3098 XA.XIR[12].XIC[10].icell.Ien Vbias 0.19161f
C3099 XA.XIR[12].XIC[2].icell.Ien Iout 0.06801f
C3100 XA.XIR[7].XIC[11].icell.Ien Vbias 0.19161f
C3101 XThR.Tn[12] XA.XIR[12].XIC[9].icell.Ien 0.14211f
C3102 XA.XIR[10].XIC[3].icell.PDM VPWR 0.01171f
C3103 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.PDM 0.02104f
C3104 XA.Cn[1] XA.XIR[12].XIC[1].icell.Ien 0.04604f
C3105 XThR.Tn[3] XA.XIR[3].XIC[14].icell.Ien 0.144f
C3106 XA.Cn[11] XA.XIR[4].XIC[11].icell.Ien 0.04604f
C3107 XThR.XTB7.B XThR.XTB4.Y 0.33064f
C3108 XA.Cn[2] XA.XIR[9].XIC[2].icell.Ien 0.04604f
C3109 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.Ien 0.04854f
C3110 XThR.XTBN.Y XThR.Tn[2] 0.6189f
C3111 XA.Cn[0] XA.XIR[6].XIC[0].icell.Ien 0.04604f
C3112 XA.Cn[8] XA.XIR[5].XIC[8].icell.PDM 0.02601f
C3113 XThR.Tn[8] Vbias 1.39526f
C3114 XA.XIR[15].XIC[5].icell.Ien VPWR 0.31713f
C3115 XA.XIR[3].XIC[0].icell.Ien Vbias 0.19149f
C3116 XThR.XTB7.B XThR.Tn[10] 0.06102f
C3117 XThR.Tn[2] XA.XIR[2].XIC[9].icell.Ien 0.14211f
C3118 XA.Cn[14] XThR.Tn[0] 0.40766f
C3119 XA.XIR[4].XIC[8].icell.Ien VPWR 0.18829f
C3120 XA.Cn[8] XThR.Tn[3] 0.40738f
C3121 XA.XIR[11].XIC[1].icell.Ien Vbias 0.19161f
C3122 XA.Cn[2] XA.Cn[3] 0.59596f
C3123 XA.Cn[13] XA.XIR[2].XIC[13].icell.Ien 0.04605f
C3124 XA.XIR[7].XIC[7].icell.PDM Vbias 0.03928f
C3125 XA.XIR[8].XIC[2].icell.Ien VPWR 0.18829f
C3126 XA.XIR[6].XIC[14].icell.PDM Vbias 0.03928f
C3127 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.Ien 0.04854f
C3128 XA.Cn[9] XThR.Tn[5] 0.40738f
C3129 XA.XIR[15].XIC[5].icell.PDM Vbias 0.03928f
C3130 XA.XIR[0].XIC[11].icell.PDM VPWR 0.01132f
C3131 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13] 0.14211f
C3132 XA.Cn[9] XA.XIR[0].XIC[9].icell.PDM 0.02801f
C3133 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.Ien 0.04854f
C3134 XA.XIR[15].XIC[14].icell.Ien Vbias 0.15966f
C3135 XA.XIR[9].XIC[11].icell.Ien VPWR 0.18829f
C3136 XA.Cn[8] XA.XIR[6].XIC[8].icell.Ien 0.04604f
C3137 thermo15c_0.XTB6.Y thermo15c_0.XTB7.Y 2.05133f
C3138 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.PDM 0.02104f
C3139 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.PDM 0.02104f
C3140 XA.XIR[12].XIC[14].icell.PDM VPWR 0.0118f
C3141 XA.XIR[9].XIC[3].icell.PDM Vbias 0.03928f
C3142 XThR.Tn[9] XA.XIR[9].XIC[7].icell.Ien 0.14211f
C3143 XA.XIR[0].XIC[4].icell.Ien VPWR 0.18788f
C3144 XA.Cn[2] VPWR 3.64821f
C3145 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PDM 0.04035f
C3146 XThR.Tn[0] Iout 1.12768f
C3147 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PDM 0.04035f
C3148 XA.XIR[15].XIC_15.icell.PDM VPWR 0.07867f
C3149 XA.Cn[0] XA.XIR[2].XIC[0].icell.PDM 0.02602f
C3150 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.PDM 0.02104f
C3151 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.Ien 0.04854f
C3152 XA.XIR[7].XIC[7].icell.Ien VPWR 0.18829f
C3153 XThR.XTB5.Y XThR.XTB7.Y 0.036f
C3154 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.04035f
C3155 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.PDM 0.02104f
C3156 XA.Cn[12] XThR.Tn[2] 0.40741f
C3157 XA.XIR[7].XIC_dummy_left.icell.Ien XThR.Tn[7] 0.01256f
C3158 XA.XIR[3].XIC[8].icell.Ien Vbias 0.19161f
C3159 XA.XIR[1].XIC[8].icell.PDM Vbias 0.03928f
C3160 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.Ien 0.04854f
C3161 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.Ien 0.04854f
C3162 XA.XIR[4].XIC[8].icell.PDM Vbias 0.03928f
C3163 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR 0.38922f
C3164 XA.Cn[11] XA.XIR[6].XIC[11].icell.PDM 0.02601f
C3165 XA.XIR[1].XIC[3].icell.Ien Vbias 0.19173f
C3166 XA.Cn[14] XA.XIR[2].XIC[14].icell.PDM 0.02602f
C3167 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.Ien 0.04854f
C3168 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.PDM 0.02104f
C3169 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PDM 0.0404f
C3170 XA.XIR[9].XIC[3].icell.Ien Iout 0.06801f
C3171 XThR.Tn[11] XA.XIR[11].XIC[3].icell.Ien 0.14211f
C3172 XA.Cn[3] XA.XIR[13].XIC[3].icell.PDM 0.02601f
C3173 XA.XIR[12].XIC_15.icell.Ien Vbias 0.19195f
C3174 XA.XIR[8].XIC[11].icell.Ien Vbias 0.19161f
C3175 XThR.Tn[12] XA.XIR[12].XIC[14].icell.Ien 0.144f
C3176 XA.Cn[1] Vbias 0.83728f
C3177 XA.Cn[13] XThR.Tn[6] 0.40739f
C3178 XThR.Tn[0] XA.XIR[0].XIC[8].icell.Ien 0.14211f
C3179 XA.XIR[6].XIC[2].icell.PDM VPWR 0.01171f
C3180 XThR.Tn[10] XA.XIR[10].XIC[7].icell.Ien 0.14211f
C3181 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PDM 0.04035f
C3182 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.Ien 0.04854f
C3183 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.Ien 0.04854f
C3184 XThR.XTBN.Y XThR.XTB4.Y 0.15627f
C3185 XThR.Tn[6] XA.XIR[6].XIC[2].icell.Ien 0.14211f
C3186 XA.XIR[5].XIC[9].icell.PDM VPWR 0.01171f
C3187 XA.XIR[5].XIC[12].icell.Ien Iout 0.06801f
C3188 XA.XIR[11].XIC_dummy_left.icell.Iout XA.XIR[12].XIC_dummy_left.icell.Iout 0.03665f
C3189 XA.XIR[13].XIC[3].icell.PDM VPWR 0.01171f
C3190 XThR.Tn[7] XA.XIR[7].XIC[9].icell.Ien 0.14211f
C3191 XA.XIR[15].XIC[12].icell.Ien Vbias 0.15966f
C3192 thermo15c_0.XTB7.A a_4861_9615# 0.02294f
C3193 XA.XIR[0].XIC[13].icell.Ien Vbias 0.19213f
C3194 XThR.XTBN.Y XThR.Tn[10] 0.46535f
C3195 XA.XIR[12].XIC[8].icell.PDM VPWR 0.01171f
C3196 XA.Cn[4] XA.XIR[10].XIC[4].icell.Ien 0.04604f
C3197 XThR.XTB1.Y XThR.XTB7.Y 0.05211f
C3198 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.Ien 0.04854f
C3199 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.Ien 0.04854f
C3200 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.Ien 0.04854f
C3201 a_6243_9615# XA.Cn[6] 0.26385f
C3202 XA.Cn[8] XThR.Tn[11] 0.40738f
C3203 XA.Cn[0] XA.XIR[7].XIC[0].icell.PDM 0.02601f
C3204 XA.XIR[12].XIC[7].icell.Ien Iout 0.06801f
C3205 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.Ien 0.04854f
C3206 XA.Cn[14] XThR.Tn[1] 0.40747f
C3207 VPWR bias[0] 2.10172f
C3208 XA.XIR[10].XIC[13].icell.Ien VPWR 0.18829f
C3209 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3210 XA.XIR[14].XIC[1].icell.Ien Vbias 0.19161f
C3211 XA.XIR[3].XIC[4].icell.Ien VPWR 0.18829f
C3212 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PDM 0.04035f
C3213 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.PDM 0.02104f
C3214 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.Ien 0.04854f
C3215 XA.Cn[10] XA.XIR[9].XIC[10].icell.Ien 0.04604f
C3216 XA.Cn[6] XThR.Tn[7] 0.40738f
C3217 XThR.XTB4.Y XThR.Tn[10] 0.01391f
C3218 XA.XIR[10].XIC[2].icell.PDM Vbias 0.03928f
C3219 XA.Cn[14] XThR.Tn[12] 0.40742f
C3220 XThR.Tn[2] XA.XIR[2].XIC[14].icell.Ien 0.144f
C3221 XA.XIR[6].XIC_dummy_right.icell.Iout XA.XIR[7].XIC_dummy_right.icell.Iout 0.04047f
C3222 XA.XIR[12].XIC[13].icell.PDM VPWR 0.01171f
C3223 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.PDM 0.02104f
C3224 XA.XIR[8].XIC[6].icell.PDM VPWR 0.01171f
C3225 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Iout 0.03908f
C3226 XA.XIR[3].XIC[4].icell.PDM VPWR 0.01171f
C3227 XA.XIR[4].XIC[13].icell.Ien VPWR 0.18829f
C3228 XA.XIR[6].XIC[3].icell.Ien Vbias 0.19161f
C3229 XThR.XTB7.B data[6] 0.07481f
C3230 XA.Cn[14] XA.XIR[7].XIC[14].icell.PDM 0.02601f
C3231 thermo15c_0.XTB3.Y Vbias 0.01224f
C3232 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.PDM 0.02104f
C3233 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Iout 0.03843f
C3234 XA.XIR[2].XIC[10].icell.PDM VPWR 0.01171f
C3235 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PDM 0.04041f
C3236 XThR.XTB5.Y XThR.Tn[11] 0.02067f
C3237 XA.XIR[8].XIC[7].icell.Ien VPWR 0.18829f
C3238 XA.Cn[13] XThR.Tn[4] 0.40739f
C3239 XA.XIR[1].XIC[0].icell.Ien Iout 0.06795f
C3240 XA.XIR[15].XIC[14].icell.PDM VPWR 0.01521f
C3241 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.PDM 0.02104f
C3242 XThR.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.14211f
C3243 XA.XIR[4].XIC[0].icell.Ien Iout 0.06795f
C3244 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.Ien 0.04854f
C3245 XThR.Tn[1] Iout 1.12765f
C3246 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.Ien 0.04854f
C3247 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PDM 0.04035f
C3248 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3249 a_8739_9569# XA.Cn[10] 0.21014f
C3250 thermo15c_0.XTBN.Y a_5155_9615# 0.07602f
C3251 XA.Cn[12] XThR.Tn[10] 0.40738f
C3252 XThR.Tn[12] Iout 1.12762f
C3253 XA.XIR[0].XIC[9].icell.Ien VPWR 0.18925f
C3254 XThR.Tn[9] XA.XIR[9].XIC[12].icell.Ien 0.14211f
C3255 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR 0.01604f
C3256 XA.XIR[2].XIC[1].icell.Ien Vbias 0.19161f
C3257 XA.XIR[0].XIC[10].icell.PDM Vbias 0.03945f
C3258 XA.XIR[11].XIC[2].icell.Ien Vbias 0.19161f
C3259 XA.Cn[5] XA.XIR[5].XIC[5].icell.Ien 0.04604f
C3260 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.PDM 0.02104f
C3261 XA.XIR[15].XIC[10].icell.Ien Vbias 0.15966f
C3262 XA.XIR[15].XIC[2].icell.Ien Iout 0.07192f
C3263 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PDM 0.04035f
C3264 XA.Cn[4] XThR.Tn[3] 0.40738f
C3265 XA.XIR[10].XIC[4].icell.Ien Vbias 0.19161f
C3266 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PDM 0.04035f
C3267 XThR.XTBN.Y a_n997_1803# 0.22873f
C3268 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PDM 0.04035f
C3269 XA.Cn[6] XA.XIR[1].XIC[6].icell.PDM 0.02602f
C3270 XA.XIR[7].XIC[12].icell.Ien VPWR 0.18829f
C3271 XA.XIR[4].XIC[5].icell.Ien Iout 0.06801f
C3272 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.PDM 0.02104f
C3273 XThR.Tn[13] XA.XIR[13].XIC[2].icell.Ien 0.14211f
C3274 XA.Cn[6] XA.XIR[4].XIC[6].icell.PDM 0.02601f
C3275 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.Ien 0.04854f
C3276 XA.XIR[3].XIC[13].icell.Ien Vbias 0.19161f
C3277 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PDM 0.04035f
C3278 XA.Cn[7] XA.XIR[0].XIC[7].icell.Ien 0.04658f
C3279 XA.Cn[5] XThR.Tn[5] 0.40738f
C3280 XA.XIR[10].XIC[11].icell.Ien VPWR 0.18829f
C3281 XThR.XTB6.A XThR.XTB2.Y 0.18237f
C3282 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.Ien 0.04854f
C3283 XA.XIR[2].XIC[6].icell.Ien Vbias 0.19161f
C3284 XA.XIR[3].XIC[1].icell.Ien VPWR 0.18829f
C3285 thermo15c_0.XTB6.Y XA.Cn[9] 0.0246f
C3286 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.PDM 0.02104f
C3287 XA.Cn[11] XA.XIR[11].XIC[11].icell.PDM 0.02601f
C3288 XA.Cn[1] XThR.Tn[0] 0.40762f
C3289 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout 0.06446f
C3290 XA.XIR[1].XIC[8].icell.Ien Vbias 0.19173f
C3291 XA.Cn[2] XA.XIR[11].XIC[2].icell.PDM 0.02601f
C3292 XA.XIR[9].XIC[8].icell.Ien Iout 0.06801f
C3293 thermo15c_0.XTB7.B data[2] 0.07481f
C3294 XThR.Tn[11] XA.XIR[11].XIC[8].icell.Ien 0.14211f
C3295 thermo15c_0.XTBN.Y XA.Cn[12] 0.46758f
C3296 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PDM 0.0404f
C3297 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.PDM 0.02104f
C3298 XA.XIR[7].XIC[10].icell.PDM VPWR 0.01171f
C3299 XA.XIR[9].XIC_dummy_left.icell.Iout VPWR 0.10954f
C3300 XA.Cn[12] XA.XIR[3].XIC[12].icell.PDM 0.02601f
C3301 XThR.XTBN.Y XThR.Tn[13] 0.56841f
C3302 XA.Cn[10] Iout 0.22426f
C3303 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.PDM 0.02104f
C3304 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.PDM 0.02104f
C3305 XA.Cn[4] XA.XIR[13].XIC[4].icell.Ien 0.04604f
C3306 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.Ien 0.04854f
C3307 XA.XIR[15].XIC[8].icell.PDM VPWR 0.01512f
C3308 XThR.Tn[0] XA.XIR[0].XIC[13].icell.Ien 0.14211f
C3309 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.PDM 0.02104f
C3310 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.PDM 0.02104f
C3311 XThR.Tn[6] XA.XIR[6].XIC[7].icell.Ien 0.14211f
C3312 XThR.Tn[12] XA.XIR[12].XIC[10].icell.Ien 0.14211f
C3313 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.PDM 0.02104f
C3314 XA.XIR[7].XIC[4].icell.Ien Iout 0.06801f
C3315 XA.XIR[0].XIC_dummy_left.icell.Iout XA.XIR[1].XIC_dummy_left.icell.Iout 0.03665f
C3316 XA.Cn[8] XThR.Tn[14] 0.40738f
C3317 thermo15c_0.XTB5.Y XA.Cn[10] 0.01755f
C3318 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.PDM 0.02104f
C3319 XThR.Tn[7] XA.XIR[7].XIC[14].icell.Ien 0.144f
C3320 XA.XIR[6].XIC[1].icell.PDM Vbias 0.03928f
C3321 XA.XIR[9].XIC[6].icell.PDM VPWR 0.01171f
C3322 XA.XIR[13].XIC[13].icell.Ien VPWR 0.18829f
C3323 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.Ien 0.04854f
C3324 thermo15c_0.XTB7.Y a_10051_9569# 0.013f
C3325 XA.XIR[5].XIC[8].icell.PDM Vbias 0.03928f
C3326 XA.XIR[12].XIC[12].icell.PDM VPWR 0.01171f
C3327 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.Ien 0.04854f
C3328 XA.XIR[13].XIC[2].icell.PDM Vbias 0.03928f
C3329 XThR.Tn[3] Vbias 1.39527f
C3330 thermo15c_0.XTB6.A thermo15c_0.XTB5.Y 0.01866f
C3331 thermo15c_0.XTB2.Y thermo15c_0.XTB7.B 0.22599f
C3332 XA.XIR[15].XIC[13].icell.PDM VPWR 0.01512f
C3333 XA.XIR[12].XIC[7].icell.PDM Vbias 0.03928f
C3334 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PDM 0.04035f
C3335 XA.XIR[1].XIC[11].icell.PDM VPWR 0.01171f
C3336 XA.XIR[3].XIC[9].icell.Ien VPWR 0.18829f
C3337 XA.Cn[9] XA.XIR[1].XIC[9].icell.PDM 0.02602f
C3338 XA.XIR[2].XIC[2].icell.Ien VPWR 0.18829f
C3339 XA.XIR[2].XIC_dummy_right.icell.Iout XA.XIR[3].XIC_dummy_right.icell.Iout 0.04047f
C3340 XA.XIR[4].XIC[11].icell.PDM VPWR 0.01171f
C3341 XA.Cn[9] XA.XIR[4].XIC[9].icell.PDM 0.02601f
C3342 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PDM 0.04035f
C3343 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.PDM 0.02104f
C3344 XA.XIR[1].XIC[4].icell.Ien VPWR 0.18829f
C3345 thermo15c_0.XTB7.B VPWR 1.33508f
C3346 XA.XIR[15].XIC_15.icell.Ien Vbias 0.15966f
C3347 XA.XIR[6].XIC[8].icell.Ien Vbias 0.19161f
C3348 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PDM 0.04035f
C3349 XA.Cn[7] XA.XIR[3].XIC[7].icell.Ien 0.04604f
C3350 XA.Cn[12] XThR.Tn[13] 0.40738f
C3351 XA.Cn[10] XA.XIR[12].XIC[10].icell.Ien 0.04604f
C3352 XA.XIR[8].XIC[12].icell.Ien VPWR 0.18829f
C3353 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PDM 0.04035f
C3354 XA.Cn[4] XThR.Tn[11] 0.40738f
C3355 XA.XIR[8].XIC[5].icell.PDM Vbias 0.03928f
C3356 XA.XIR[3].XIC[3].icell.PDM Vbias 0.03928f
C3357 XA.Cn[0] XThR.Tn[6] 0.40736f
C3358 XA.XIR[14].XIC[2].icell.Ien Vbias 0.19161f
C3359 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.Ien 0.04854f
C3360 XThR.XTB7.B a_n997_3979# 0.01152f
C3361 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.PDM 0.02104f
C3362 XA.XIR[2].XIC[9].icell.PDM Vbias 0.03928f
C3363 XA.XIR[13].XIC[4].icell.Ien Vbias 0.19161f
C3364 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.Ien 0.04854f
C3365 XA.Cn[9] XThR.Tn[9] 0.40738f
C3366 XA.Cn[10] XThR.Tn[8] 0.40738f
C3367 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PDM 0.04035f
C3368 XA.XIR[0].XIC[14].icell.Ien VPWR 0.18783f
C3369 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.Ien 0.04854f
C3370 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.Ien 0.04854f
C3371 XA.XIR[11].XIC[7].icell.Ien Vbias 0.19161f
C3372 XThR.Tn[14] XA.XIR[14].XIC[3].icell.Ien 0.14211f
C3373 XThR.Tn[1] XA.XIR[1].XIC[3].icell.Ien 0.14211f
C3374 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.PDM 0.02104f
C3375 XA.XIR[15].XIC[7].icell.Ien Iout 0.07192f
C3376 XA.XIR[10].XIC[9].icell.Ien Vbias 0.19161f
C3377 XA.Cn[13] XA.XIR[5].XIC[13].icell.Ien 0.04604f
C3378 XA.XIR[13].XIC[11].icell.Ien VPWR 0.18829f
C3379 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.04035f
C3380 XA.XIR[4].XIC[10].icell.Ien Iout 0.06801f
C3381 XA.Cn[13] XA.XIR[8].XIC[13].icell.PDM 0.02601f
C3382 XA.Cn[11] XA.XIR[14].XIC[11].icell.PDM 0.02601f
C3383 XThR.Tn[13] XA.XIR[13].XIC[7].icell.Ien 0.14211f
C3384 XA.XIR[0].XIC[1].icell.Ien Iout 0.0675f
C3385 XA.Cn[6] XA.XIR[7].XIC[6].icell.Ien 0.04604f
C3386 XA.Cn[2] XA.XIR[14].XIC[2].icell.PDM 0.02601f
C3387 XA.Cn[1] XThR.Tn[1] 0.40744f
C3388 XThR.Tn[12] XA.XIR[12].XIC_15.icell.Ien 0.13564f
C3389 thermo15c_0.XTB5.A thermo15c_0.XTBN.A 0.06305f
C3390 XA.Cn[5] XA.XIR[12].XIC[5].icell.Ien 0.04604f
C3391 XA.XIR[8].XIC[4].icell.Ien Iout 0.06801f
C3392 XA.XIR[11].XIC[1].icell.PDM VPWR 0.01171f
C3393 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.Ien 0.04854f
C3394 XA.XIR[2].XIC[11].icell.Ien Vbias 0.19161f
C3395 XA.XIR[10].XIC[5].icell.PDM VPWR 0.01171f
C3396 XThR.XTB2.Y XThR.Tn[1] 0.17876f
C3397 XA.Cn[1] XThR.Tn[12] 0.40738f
C3398 XA.XIR[1].XIC[13].icell.Ien Vbias 0.19173f
C3399 XA.XIR[9].XIC[13].icell.Ien Iout 0.06801f
C3400 XThR.XTB7.B XThR.Tn[7] 0.07415f
C3401 XA.XIR[6].XIC[4].icell.Ien VPWR 0.18829f
C3402 XThR.XTB7.B a_n997_2891# 0.0168f
C3403 XA.XIR[12].XIC[11].icell.PDM VPWR 0.01171f
C3404 XA.XIR[0].XIC[6].icell.Ien Iout 0.0675f
C3405 XA.Cn[3] XA.XIR[11].XIC[3].icell.Ien 0.04604f
C3406 XA.Cn[0] XThR.Tn[4] 0.40739f
C3407 XA.XIR[12].XIC[0].icell.Ien Vbias 0.19149f
C3408 XA.Cn[0] XA.XIR[12].XIC[0].icell.PDM 0.02601f
C3409 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.Ien 0.04854f
C3410 thermo15c_0.XTBN.A XA.Cn[12] 0.22871f
C3411 XThR.Tn[11] Vbias 1.39532f
C3412 XA.XIR[15].XIC[12].icell.PDM VPWR 0.01512f
C3413 XThR.Tn[6] XA.XIR[6].XIC[12].icell.Ien 0.14211f
C3414 XA.XIR[7].XIC[9].icell.Ien Iout 0.06801f
C3415 XA.XIR[7].XIC[9].icell.PDM Vbias 0.03928f
C3416 XThR.XTB6.A XThR.XTB7.Y 0.01596f
C3417 XThR.XTB3.Y XThR.XTB5.Y 0.04438f
C3418 XA.Cn[6] XA.XIR[5].XIC[6].icell.PDM 0.02601f
C3419 XA.XIR[15].XIC[7].icell.PDM Vbias 0.03928f
C3420 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.PDM 0.02104f
C3421 XA.XIR[0].XIC[13].icell.PDM VPWR 0.01132f
C3422 thermo15c_0.XTB6.Y XA.Cn[5] 0.20249f
C3423 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.Ien 0.04854f
C3424 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.PDM 0.02104f
C3425 XA.XIR[11].XIC[3].icell.Ien VPWR 0.18829f
C3426 XThR.XTBN.A data[4] 0.02581f
C3427 XA.XIR[10].XIC[5].icell.Ien VPWR 0.18829f
C3428 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout 0.06446f
C3429 thermo15c_0.XTBN.A thermo15c_0.XTBN.Y 0.77125f
C3430 thermo15c_0.XTBN.Y a_7651_9569# 0.23021f
C3431 XA.XIR[9].XIC[5].icell.PDM Vbias 0.03928f
C3432 XA.XIR[2].XIC[0].icell.Ien Iout 0.06795f
C3433 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.Ien 0.04854f
C3434 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PDM 0.04035f
C3435 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PDM 0.04035f
C3436 XA.XIR[3].XIC[14].icell.Ien VPWR 0.18835f
C3437 XA.Cn[6] Iout 0.22423f
C3438 thermo15c_0.XTB7.A data[0] 0.86893f
C3439 XA.Cn[7] XA.XIR[0].XIC[7].icell.PDM 0.02803f
C3440 XA.XIR[10].XIC[1].icell.Ien Iout 0.06801f
C3441 XThR.XTBN.Y a_n997_3979# 0.23021f
C3442 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.Ien 0.04854f
C3443 XA.XIR[2].XIC[7].icell.Ien VPWR 0.18829f
C3444 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PDM 0.04056f
C3445 XA.Cn[4] XThR.Tn[14] 0.40738f
C3446 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.PDM 0.02104f
C3447 XA.XIR[1].XIC[9].icell.Ien VPWR 0.18829f
C3448 XA.XIR[1].XIC[10].icell.PDM Vbias 0.03928f
C3449 XThR.Tn[8] XA.XIR[8].XIC[4].icell.Ien 0.14211f
C3450 XA.XIR[14].XIC_dummy_left.icell.Iout XA.XIR[15].XIC_dummy_left.icell.Iout 0.03665f
C3451 XA.Cn[4] XA.XIR[10].XIC[4].icell.PDM 0.02601f
C3452 XA.XIR[6].XIC[13].icell.Ien Vbias 0.19161f
C3453 XA.XIR[10].XIC[14].icell.Ien Vbias 0.19161f
C3454 XA.Cn[8] VPWR 4.5473f
C3455 XA.XIR[2].XIC_dummy_left.icell.Iout XA.XIR[3].XIC_dummy_left.icell.Iout 0.03665f
C3456 XA.XIR[4].XIC[10].icell.PDM Vbias 0.03928f
C3457 XA.XIR[1].XIC_dummy_right.icell.Iout XA.XIR[2].XIC_dummy_right.icell.Iout 0.04047f
C3458 XA.Cn[13] XA.XIR[9].XIC[13].icell.PDM 0.02601f
C3459 XThR.XTB1.Y XThR.XTB3.Y 0.04033f
C3460 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.Ien 0.04854f
C3461 XA.Cn[6] XA.XIR[8].XIC[6].icell.Ien 0.04604f
C3462 XA.XIR[14].XIC[7].icell.Ien Vbias 0.19161f
C3463 XThR.XTB7.A data[5] 0.06538f
C3464 XA.Cn[7] XA.XIR[1].XIC[7].icell.Ien 0.04606f
C3465 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PDM 0.0404f
C3466 XThR.Tn[5] XA.XIR[5].XIC[3].icell.Ien 0.14211f
C3467 XA.XIR[13].XIC[9].icell.Ien Vbias 0.19161f
C3468 XA.XIR[11].XIC[13].icell.Ien Iout 0.06801f
C3469 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout 0.06446f
C3470 XA.XIR[3].XIC[6].icell.Ien Iout 0.06801f
C3471 XA.XIR[6].XIC[4].icell.PDM VPWR 0.01171f
C3472 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PDM 0.04056f
C3473 XThR.XTB7.A a_n1049_6699# 0.02294f
C3474 XThR.Tn[14] XA.XIR[14].XIC[8].icell.Ien 0.14211f
C3475 XA.XIR[14].XIC[1].icell.PDM VPWR 0.01171f
C3476 XThR.XTB5.Y VPWR 1.0269f
C3477 XA.XIR[5].XIC[11].icell.PDM VPWR 0.01171f
C3478 XThR.Tn[1] XA.XIR[1].XIC[8].icell.Ien 0.14211f
C3479 thermo15c_0.XTB3.Y XA.Cn[10] 0.29566f
C3480 XA.Cn[9] XA.XIR[5].XIC[9].icell.PDM 0.02601f
C3481 XThR.XTBN.Y XThR.Tn[7] 0.89994f
C3482 XThR.XTBN.Y a_n997_2891# 0.22804f
C3483 XA.XIR[13].XIC[5].icell.PDM VPWR 0.01171f
C3484 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.Ien 0.04854f
C3485 XA.XIR[4].XIC_15.icell.Ien Iout 0.0694f
C3486 thermo15c_0.XTB7.A a_5949_9615# 0.01824f
C3487 thermo15c_0.XTB7.B thermo15c_0.XTB7.Y 0.33493f
C3488 XA.XIR[12].XIC[10].icell.PDM VPWR 0.01171f
C3489 XA.Cn[0] XA.XIR[11].XIC[0].icell.Ien 0.04604f
C3490 XA.XIR[8].XIC[9].icell.Ien Iout 0.06801f
C3491 XA.Cn[14] XA.XIR[7].XIC[14].icell.Ien 0.04604f
C3492 thermo15c_0.XTB4.Y XA.Cn[3] 0.1917f
C3493 XA.XIR[15].XIC[11].icell.PDM VPWR 0.01512f
C3494 thermo15c_0.XTB2.Y thermo15c_0.XTB4.Y 0.04006f
C3495 thermo15c_0.XTB6.A thermo15c_0.XTB3.Y 0.03869f
C3496 XA.Cn[3] XA.XIR[14].XIC[3].icell.Ien 0.04604f
C3497 XThR.Tn[5] XThR.Tn[6] 0.11432f
C3498 XA.Cn[0] XA.XIR[15].XIC[0].icell.PDM 0.02601f
C3499 XA.XIR[5].XIC[1].icell.Ien Vbias 0.19161f
C3500 XA.Cn[5] XThR.Tn[9] 0.40738f
C3501 XA.Cn[6] XThR.Tn[8] 0.40738f
C3502 XA.Cn[10] XA.XIR[0].XIC[10].icell.PDM 0.02792f
C3503 XThR.XTB4.Y XThR.Tn[7] 0.01797f
C3504 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PDM 0.04035f
C3505 XThR.Tn[14] Vbias 1.39537f
C3506 XA.Cn[10] XA.XIR[15].XIC[10].icell.Ien 0.04292f
C3507 XA.XIR[11].XIC[0].icell.PDM Vbias 0.03915f
C3508 XA.XIR[6].XIC[9].icell.Ien VPWR 0.18829f
C3509 XA.XIR[10].XIC[4].icell.PDM Vbias 0.03928f
C3510 XA.XIR[0].XIC[11].icell.Ien Iout 0.0675f
C3511 XA.XIR[10].XIC[12].icell.Ien Vbias 0.19161f
C3512 XA.XIR[4].XIC_dummy_right.icell.Iout Iout 0.01732f
C3513 XThR.Tn[10] a_n997_2891# 0.1927f
C3514 thermo15c_0.XTB4.Y VPWR 0.91479f
C3515 XA.Cn[1] XA.XIR[0].XIC[1].icell.Ien 0.04659f
C3516 XA.XIR[3].XIC[6].icell.PDM VPWR 0.01171f
C3517 XA.XIR[8].XIC[8].icell.PDM VPWR 0.01171f
C3518 XA.XIR[14].XIC[3].icell.Ien VPWR 0.18883f
C3519 XA.Cn[1] XA.XIR[2].XIC[1].icell.PDM 0.02602f
C3520 XA.XIR[2].XIC[12].icell.PDM VPWR 0.01171f
C3521 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.PDM 0.02104f
C3522 XA.XIR[13].XIC[5].icell.Ien VPWR 0.18829f
C3523 XA.XIR[7].XIC[14].icell.Ien Iout 0.06801f
C3524 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PDM 0.04035f
C3525 XA.Cn[7] XA.XIR[6].XIC[7].icell.Ien 0.04604f
C3526 XA.XIR[5].XIC[6].icell.Ien Vbias 0.19161f
C3527 XThR.XTB1.Y VPWR 1.13148f
C3528 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.Ien 0.04854f
C3529 XThR.XTB6.Y a_n1319_5611# 0.01283f
C3530 XA.XIR[11].XIC[11].icell.Ien Iout 0.06801f
C3531 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.PDM 0.02104f
C3532 XA.Cn[12] XThR.Tn[7] 0.40738f
C3533 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3534 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PDM 0.0404f
C3535 XA.XIR[11].XIC[8].icell.Ien VPWR 0.18829f
C3536 XA.XIR[13].XIC[1].icell.Ien Iout 0.06801f
C3537 XThR.XTB7.Y XThR.Tn[12] 0.07066f
C3538 thermo15c_0.XTBN.Y a_6243_9615# 0.07767f
C3539 XA.Cn[11] XA.XIR[12].XIC[11].icell.Ien 0.04604f
C3540 XA.Cn[12] XA.XIR[6].XIC[12].icell.PDM 0.02601f
C3541 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.Ien 0.04854f
C3542 XA.XIR[0].XIC[12].icell.PDM Vbias 0.03945f
C3543 XA.Cn[9] XA.XIR[0].XIC[9].icell.Ien 0.04656f
C3544 XA.Cn[5] XA.XIR[15].XIC[5].icell.Ien 0.04292f
C3545 XA.Cn[4] XA.XIR[13].XIC[4].icell.PDM 0.02601f
C3546 XA.XIR[13].XIC[14].icell.Ien Vbias 0.19161f
C3547 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PDM 0.04035f
C3548 XThR.Tn[4] XThR.Tn[5] 0.12171f
C3549 thermo15c_0.XTBN.A a_7651_9569# 0.02087f
C3550 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PDM 0.04035f
C3551 XA.XIR[2].XIC[12].icell.Ien VPWR 0.18829f
C3552 XA.Cn[13] XA.XIR[11].XIC[13].icell.PDM 0.02601f
C3553 XA.XIR[1].XIC[14].icell.Ien VPWR 0.18835f
C3554 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PDM 0.04056f
C3555 XThR.Tn[8] XA.XIR[8].XIC[9].icell.Ien 0.14211f
C3556 XA.XIR[14].XIC[13].icell.Ien Iout 0.06801f
C3557 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.PDM 0.02104f
C3558 XThR.XTB6.Y XThR.Tn[5] 0.20186f
C3559 XA.XIR[3].XIC_dummy_left.icell.Iout VPWR 0.11229f
C3560 XA.Cn[10] XThR.Tn[3] 0.40738f
C3561 XA.XIR[12].XIC[1].icell.Ien VPWR 0.18829f
C3562 XA.XIR[10].XIC[10].icell.Ien Vbias 0.19161f
C3563 XA.XIR[1].XIC[1].icell.Ien Iout 0.06801f
C3564 a_10915_9569# Vbias 0.01451f
C3565 XA.Cn[14] XA.XIR[8].XIC[14].icell.Ien 0.04604f
C3566 XA.XIR[10].XIC[2].icell.Ien Iout 0.06801f
C3567 XA.Cn[3] XA.Cn[4] 0.45992f
C3568 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.Ien 0.04854f
C3569 XThR.Tn[5] XA.XIR[5].XIC[8].icell.Ien 0.14211f
C3570 XA.Cn[1] XA.XIR[7].XIC[1].icell.PDM 0.02601f
C3571 XA.Cn[1] XA.XIR[10].XIC[1].icell.Ien 0.04604f
C3572 XThR.XTBN.Y a_n997_1579# 0.23006f
C3573 XA.XIR[5].XIC[2].icell.Ien VPWR 0.18829f
C3574 XThR.XTB7.Y a_n1049_5317# 0.27822f
C3575 XA.XIR[7].XIC[12].icell.PDM VPWR 0.01171f
C3576 XA.Cn[11] XThR.Tn[5] 0.40738f
C3577 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout 0.06446f
C3578 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.PDM 0.02104f
C3579 XA.XIR[15].XIC[10].icell.PDM VPWR 0.01512f
C3580 XA.XIR[3].XIC[11].icell.Ien Iout 0.06801f
C3581 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.Ien 0.04854f
C3582 XThR.Tn[1] XA.XIR[1].XIC[13].icell.Ien 0.14211f
C3583 XA.XIR[2].XIC[4].icell.Ien Iout 0.06801f
C3584 XA.Cn[4] VPWR 3.6464f
C3585 XA.XIR[1].XIC[6].icell.Ien Iout 0.06801f
C3586 XA.XIR[9].XIC[8].icell.PDM VPWR 0.01171f
C3587 XA.XIR[6].XIC[3].icell.PDM Vbias 0.03928f
C3588 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.Ien 0.04854f
C3589 XA.XIR[0].XIC[0].icell.PDM VPWR 0.01132f
C3590 XA.XIR[14].XIC[0].icell.PDM Vbias 0.03915f
C3591 XA.XIR[5].XIC[10].icell.PDM Vbias 0.03928f
C3592 thermo15c_0.XTB7.Y XA.Cn[8] 0.07809f
C3593 thermo15c_0.XTB3.Y a_4067_9615# 0.23056f
C3594 XA.XIR[8].XIC[14].icell.Ien Iout 0.06801f
C3595 XA.XIR[13].XIC[4].icell.PDM Vbias 0.03928f
C3596 XA.XIR[13].XIC[12].icell.Ien Vbias 0.19161f
C3597 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12] 0.14211f
C3598 XA.Cn[14] XThR.Tn[2] 0.40744f
C3599 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.Ien 0.04854f
C3600 XA.XIR[12].XIC[9].icell.PDM Vbias 0.03928f
C3601 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PDM 0.04035f
C3602 XThR.Tn[11] XThR.Tn[12] 0.1626f
C3603 a_8963_9569# XA.Cn[11] 0.1927f
C3604 XA.XIR[1].XIC[13].icell.PDM VPWR 0.01171f
C3605 XA.XIR[9].XIC[2].icell.Ien Vbias 0.19161f
C3606 XA.Cn[9] XA.XIR[3].XIC[9].icell.Ien 0.04604f
C3607 XA.XIR[6].XIC[14].icell.Ien VPWR 0.18835f
C3608 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PDM 0.04035f
C3609 XA.XIR[4].XIC[13].icell.PDM VPWR 0.01171f
C3610 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PDM 0.04035f
C3611 XA.XIR[14].XIC[11].icell.Ien Iout 0.06801f
C3612 XA.Cn[0] XA.XIR[7].XIC[0].icell.Ien 0.04604f
C3613 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3614 XA.XIR[14].XIC[8].icell.Ien VPWR 0.18883f
C3615 thermo15c_0.XTB7.B XA.Cn[9] 0.05542f
C3616 XThR.XTB5.A XThR.XTBN.A 0.06303f
C3617 XA.XIR[6].XIC[1].icell.Ien Iout 0.06801f
C3618 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.PDM 0.02104f
C3619 XA.Cn[7] XA.XIR[1].XIC[7].icell.PDM 0.02602f
C3620 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PDM 0.04035f
C3621 XA.XIR[5].XIC[11].icell.Ien Vbias 0.19161f
C3622 XA.Cn[3] Vbias 0.84088f
C3623 a_3773_9615# XA.Cn[2] 0.01043f
C3624 XA.XIR[3].XIC[5].icell.PDM Vbias 0.03928f
C3625 thermo15c_0.XTB2.Y Vbias 0.01484f
C3626 XThR.Tn[2] Iout 1.12764f
C3627 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.PDM 0.02104f
C3628 XA.XIR[8].XIC[7].icell.PDM Vbias 0.03928f
C3629 XA.Cn[7] XA.XIR[4].XIC[7].icell.PDM 0.02601f
C3630 XA.XIR[2].XIC[11].icell.PDM Vbias 0.03928f
C3631 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR 0.39005f
C3632 XA.Cn[4] XA.XIR[4].XIC[4].icell.Ien 0.04604f
C3633 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.PDM 0.02104f
C3634 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PDM 0.04035f
C3635 XThR.XTBN.Y a_n1049_6699# 0.07601f
C3636 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.PDM 0.02104f
C3637 XA.XIR[12].XIC[6].icell.Ien Vbias 0.19161f
C3638 XA.Cn[8] XA.XIR[7].XIC[8].icell.Ien 0.04604f
C3639 XA.XIR[10].XIC_15.icell.Ien Vbias 0.19195f
C3640 XA.Cn[3] XA.XIR[11].XIC[3].icell.PDM 0.02601f
C3641 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PDM 0.04035f
C3642 XA.XIR[6].XIC[6].icell.Ien Iout 0.06801f
C3643 XA.Cn[13] XA.XIR[14].XIC[13].icell.PDM 0.02601f
C3644 VPWR Vbias 98.23621f
C3645 XA.Cn[10] XThR.Tn[11] 0.40738f
C3646 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PDM 0.04035f
C3647 XA.Cn[13] XA.XIR[3].XIC[13].icell.PDM 0.02601f
C3648 thermo15c_0.XTB4.Y thermo15c_0.XTB7.Y 0.03475f
C3649 XA.XIR[0].XIC_dummy_left.icell.Iout Iout 0.03553f
C3650 XA.Cn[6] XA.XIR[2].XIC[6].icell.Ien 0.04605f
C3651 XA.XIR[13].XIC[10].icell.Ien Vbias 0.19161f
C3652 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.PDM 0.02104f
C3653 XA.XIR[10].XIC_dummy_left.icell.Iout XA.XIR[11].XIC_dummy_left.icell.Iout 0.03665f
C3654 XThR.Tn[8] XA.XIR[8].XIC[14].icell.Ien 0.144f
C3655 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.Ien 0.04854f
C3656 XA.XIR[13].XIC[2].icell.Ien Iout 0.06801f
C3657 XThR.XTB4.Y a_n1049_6699# 0.23756f
C3658 XThR.XTB6.A XThR.XTB3.Y 0.03869f
C3659 XThR.XTB2.Y XThR.XTB7.A 0.2319f
C3660 XA.XIR[11].XIC[3].icell.PDM VPWR 0.01171f
C3661 XA.Cn[1] XA.XIR[13].XIC[1].icell.Ien 0.04604f
C3662 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.Ien 0.04854f
C3663 XA.XIR[10].XIC[7].icell.PDM VPWR 0.01171f
C3664 XThR.XTB7.B XThR.Tn[8] 0.05091f
C3665 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.PDM 0.02104f
C3666 XA.XIR[11].XIC[5].icell.Ien Iout 0.06801f
C3667 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.Ien 0.04854f
C3668 XA.XIR[10].XIC[7].icell.Ien Iout 0.06801f
C3669 XThR.Tn[5] XA.XIR[5].XIC[13].icell.Ien 0.14211f
C3670 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR 0.08547f
C3671 XA.XIR[5].XIC[7].icell.Ien VPWR 0.18829f
C3672 XThR.XTB7.A a_n1049_5611# 0.01824f
C3673 XA.Cn[10] XA.XIR[1].XIC[10].icell.PDM 0.02602f
C3674 XA.Cn[14] XThR.Tn[10] 0.40742f
C3675 XA.XIR[2].XIC[9].icell.Ien Iout 0.06801f
C3676 XA.Cn[11] XA.XIR[15].XIC[11].icell.Ien 0.04292f
C3677 XA.XIR[7].XIC[11].icell.PDM Vbias 0.03928f
C3678 XThR.Tn[13] a_n997_1579# 0.19413f
C3679 XA.Cn[10] XA.XIR[4].XIC[10].icell.PDM 0.02601f
C3680 XA.XIR[12].XIC[2].icell.Ien VPWR 0.18829f
C3681 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PDM 0.04035f
C3682 XA.XIR[1].XIC[11].icell.Ien Iout 0.06801f
C3683 XA.XIR[15].XIC[9].icell.PDM Vbias 0.03928f
C3684 XA.XIR[4].XIC[4].icell.Ien Vbias 0.19161f
C3685 XA.XIR[0].XIC_15.icell.PDM VPWR 0.07389f
C3686 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.PDM 0.02104f
C3687 XA.Cn[1] XA.XIR[1].XIC[1].icell.Ien 0.04606f
C3688 XA.Cn[6] XThR.Tn[3] 0.40738f
C3689 thermo15c_0.XTB5.Y a_5155_9615# 0.24821f
C3690 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.PDM 0.02104f
C3691 XThR.Tn[4] XA.XIR[4].XIC[3].icell.Ien 0.14211f
C3692 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.PDM 0.02104f
C3693 thermo15c_0.XTBN.Y a_8739_9569# 0.22804f
C3694 XA.XIR[9].XIC[7].icell.PDM Vbias 0.03928f
C3695 XA.Cn[0] XA.XIR[8].XIC[0].icell.PDM 0.02601f
C3696 XThR.XTBN.A XThR.Tn[9] 0.12398f
C3697 XA.Cn[7] XThR.Tn[5] 0.40738f
C3698 XA.XIR[9].XIC[7].icell.Ien Vbias 0.19161f
C3699 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.PDM 0.02104f
C3700 XThR.Tn[10] Iout 1.12758f
C3701 thermo15c_0.XTB5.A thermo15c_0.XTB5.Y 0.0538f
C3702 thermo15c_0.XTB6.Y XA.Cn[11] 0.02473f
C3703 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.Ien 0.04854f
C3704 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR 0.01604f
C3705 XA.Cn[8] XA.XIR[8].XIC[8].icell.Ien 0.04604f
C3706 XA.Cn[3] XThR.Tn[0] 0.40763f
C3707 XA.Cn[12] XA.XIR[12].XIC[12].icell.Ien 0.04604f
C3708 a_2979_9615# VPWR 0.70527f
C3709 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.PDM 0.02104f
C3710 XThR.XTB6.A VPWR 0.68638f
C3711 XA.XIR[1].XIC[12].icell.PDM Vbias 0.03928f
C3712 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PDM 0.04035f
C3713 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.Ien 0.04854f
C3714 XA.Cn[9] XA.XIR[1].XIC[9].icell.Ien 0.04606f
C3715 thermo15c_0.XTBN.Y XA.Cn[14] 0.42645f
C3716 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Iout 0.01728f
C3717 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR 0.39002f
C3718 XA.Cn[8] XA.Cn[9] 0.0619f
C3719 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.Ien 0.04854f
C3720 XA.XIR[4].XIC[12].icell.PDM Vbias 0.03928f
C3721 XA.XIR[7].XIC[3].icell.Ien Vbias 0.19161f
C3722 XThR.XTB1.Y a_n1049_8581# 0.21263f
C3723 XA.Cn[14] XA.XIR[8].XIC[14].icell.PDM 0.02601f
C3724 XA.Cn[12] Iout 0.2243f
C3725 XThR.Tn[3] XA.XIR[3].XIC[6].icell.Ien 0.14211f
C3726 XA.Cn[3] XA.XIR[14].XIC[3].icell.PDM 0.02601f
C3727 XA.XIR[13].XIC_15.icell.Ien Vbias 0.19195f
C3728 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.PDM 0.02104f
C3729 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.Ien 0.04854f
C3730 XA.Cn[10] XThR.Tn[14] 0.40738f
C3731 XThR.Tn[0] VPWR 8.08835f
C3732 thermo15c_0.XTB5.Y XA.Cn[12] 0.32158f
C3733 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PDM 0.04035f
C3734 thermo15c_0.XTB6.A data[1] 0.37233f
C3735 XThR.XTB7.B a_n997_3755# 0.01174f
C3736 XThR.XTB7.B XThR.XTB2.Y 0.22599f
C3737 XA.XIR[5].XIC_dummy_right.icell.Iout XA.XIR[6].XIC_dummy_right.icell.Iout 0.04047f
C3738 XA.Cn[12] XA.XIR[4].XIC[12].icell.Ien 0.04604f
C3739 XThR.XTBN.Y XThR.Tn[8] 0.4783f
C3740 XA.XIR[6].XIC[6].icell.PDM VPWR 0.01171f
C3741 XA.Cn[3] XA.XIR[9].XIC[3].icell.Ien 0.04604f
C3742 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.Ien 0.04854f
C3743 XA.XIR[6].XIC[11].icell.Ien Iout 0.06801f
C3744 XA.XIR[5].XIC[13].icell.PDM VPWR 0.01171f
C3745 XA.XIR[14].XIC[3].icell.PDM VPWR 0.01171f
C3746 XA.Cn[1] XA.XIR[6].XIC[1].icell.Ien 0.04604f
C3747 XA.Cn[0] XA.XIR[8].XIC[0].icell.Ien 0.04604f
C3748 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.PDM 0.02104f
C3749 XA.XIR[13].XIC[7].icell.PDM VPWR 0.01171f
C3750 XA.Cn[1] XA.XIR[12].XIC[1].icell.PDM 0.02601f
C3751 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.PDM 0.02104f
C3752 XA.XIR[14].XIC[5].icell.Ien Iout 0.06801f
C3753 XA.Cn[1] XThR.Tn[2] 0.40741f
C3754 thermo15c_0.XTB5.Y thermo15c_0.XTBN.Y 0.162f
C3755 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.Ien 0.04854f
C3756 XA.XIR[13].XIC[7].icell.Ien Iout 0.06801f
C3757 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.Ien 0.04854f
C3758 XA.Cn[14] XA.XIR[2].XIC[14].icell.Ien 0.04605f
C3759 data[5] data[6] 0.01513f
C3760 XA.XIR[9].XIC[3].icell.Ien VPWR 0.18829f
C3761 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.Ien 0.04854f
C3762 XThR.XTB4.Y XThR.Tn[8] 0.01306f
C3763 XA.Cn[7] XA.XIR[5].XIC[7].icell.PDM 0.02601f
C3764 XA.XIR[15].XIC[1].icell.Ien Vbias 0.15966f
C3765 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PDM 0.04035f
C3766 XA.Cn[14] XThR.Tn[13] 0.40742f
C3767 XA.XIR[1].XIC[0].icell.PDM VPWR 0.01171f
C3768 XA.XIR[11].XIC[2].icell.PDM Vbias 0.03928f
C3769 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.PDM 0.02104f
C3770 XA.Cn[9] XA.XIR[6].XIC[9].icell.Ien 0.04604f
C3771 XThR.XTB6.Y XThR.Tn[9] 0.0246f
C3772 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.Ien 0.04854f
C3773 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.PDM 0.02104f
C3774 XThR.XTB7.A XThR.Tn[3] 0.0306f
C3775 XA.Cn[6] XThR.Tn[11] 0.40738f
C3776 XA.XIR[10].XIC[6].icell.PDM Vbias 0.03928f
C3777 XA.XIR[4].XIC[0].icell.PDM VPWR 0.01171f
C3778 XA.XIR[5].XIC[12].icell.Ien VPWR 0.18829f
C3779 XA.Cn[0] XA.XIR[9].XIC[0].icell.PDM 0.02601f
C3780 XA.Cn[2] XThR.Tn[6] 0.40738f
C3781 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.PDM 0.02104f
C3782 thermo15c_0.XTB4.Y XA.Cn[9] 0.01318f
C3783 XA.XIR[3].XIC[8].icell.PDM VPWR 0.01171f
C3784 XA.XIR[4].XIC_15.icell.PUM VPWR 0.01655f
C3785 thermo15c_0.XTB7.Y Vbias 0.01962f
C3786 XA.XIR[8].XIC[10].icell.PDM VPWR 0.01171f
C3787 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Iout 0.01779f
C3788 XThR.XTB7.A XThR.XTB7.Y 0.37429f
C3789 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.PDM 0.02104f
C3790 XA.XIR[2].XIC[14].icell.PDM VPWR 0.0118f
C3791 XA.XIR[2].XIC[14].icell.Ien Iout 0.06801f
C3792 XA.XIR[15].XIC[6].icell.Ien Vbias 0.15966f
C3793 XA.Cn[11] XThR.Tn[9] 0.40738f
C3794 XA.Cn[12] XThR.Tn[8] 0.40738f
C3795 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PDM 0.04035f
C3796 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.PDM 0.02104f
C3797 XA.XIR[12].XIC[7].icell.Ien VPWR 0.18829f
C3798 XA.XIR[4].XIC[9].icell.Ien Vbias 0.19161f
C3799 XA.XIR[14].XIC[0].icell.Ien Iout 0.06795f
C3800 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3801 XA.XIR[0].XIC[0].icell.Ien Vbias 0.19209f
C3802 XA.Cn[10] XA.XIR[10].XIC[10].icell.Ien 0.04604f
C3803 XA.Cn[5] XA.XIR[10].XIC[5].icell.PDM 0.02601f
C3804 XA.XIR[7].XIC_dummy_right.icell.Iout XA.XIR[8].XIC_dummy_right.icell.Iout 0.04047f
C3805 XThR.Tn[13] Iout 1.12765f
C3806 XA.XIR[8].XIC[3].icell.Ien Vbias 0.19161f
C3807 XA.Cn[14] XA.XIR[9].XIC[14].icell.PDM 0.02601f
C3808 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR 0.01669f
C3809 XThR.Tn[4] XA.XIR[4].XIC[8].icell.Ien 0.14211f
C3810 XThR.Tn[11] XA.XIR[11].XIC[13].icell.Ien 0.14211f
C3811 XA.Cn[3] XThR.Tn[1] 0.40744f
C3812 XA.XIR[0].XIC[14].icell.PDM Vbias 0.03945f
C3813 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.PDM 0.02104f
C3814 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR 0.38995f
C3815 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PDM 0.04035f
C3816 XA.XIR[9].XIC[12].icell.Ien Vbias 0.19161f
C3817 XA.XIR[5].XIC[4].icell.Ien Iout 0.06801f
C3818 thermo15c_0.XTBN.A a_8739_9569# 0.01719f
C3819 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PDM 0.04035f
C3820 XA.Cn[3] XThR.Tn[12] 0.40738f
C3821 XThR.XTBN.Y XThR.XTB2.Y 0.2075f
C3822 XA.XIR[0].XIC[5].icell.Ien Vbias 0.19213f
C3823 XThR.XTBN.Y a_n997_3755# 0.229f
C3824 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.PDM 0.02104f
C3825 XA.XIR[1].XIC[0].icell.Ien VPWR 0.18829f
C3826 thermo15c_0.XTB1.Y data[0] 0.06453f
C3827 XThR.Tn[2] XA.XIR[2].XIC[1].icell.Ien 0.14211f
C3828 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.Ien 0.04854f
C3829 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.Ien 0.04854f
C3830 XA.XIR[4].XIC[0].icell.Ien VPWR 0.18829f
C3831 XA.Cn[10] XA.XIR[5].XIC[10].icell.PDM 0.02601f
C3832 XThR.Tn[1] VPWR 8.09331f
C3833 XA.Cn[2] XThR.Tn[4] 0.40738f
C3834 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.Ien 0.04854f
C3835 XThR.Tn[12] XA.XIR[12].XIC[6].icell.Ien 0.14211f
C3836 XA.XIR[7].XIC[8].icell.Ien Vbias 0.19161f
C3837 XThR.Tn[3] XA.XIR[3].XIC[11].icell.Ien 0.14211f
C3838 XThR.Tn[12] VPWR 8.99609f
C3839 XA.Cn[5] XA.XIR[10].XIC[5].icell.Ien 0.04604f
C3840 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.PDM 0.02104f
C3841 XA.XIR[1].XIC_dummy_left.icell.Iout Iout 0.03553f
C3842 XA.XIR[13].XIC_dummy_left.icell.Iout XA.XIR[14].XIC_dummy_left.icell.Iout 0.03665f
C3843 XThR.XTBN.Y a_n1049_5611# 0.0768f
C3844 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.Ien 0.04854f
C3845 XThR.XTB2.Y XThR.XTB4.Y 0.04006f
C3846 XA.Cn[1] XThR.Tn[10] 0.40738f
C3847 XA.XIR[15].XIC[2].icell.Ien VPWR 0.31713f
C3848 XA.XIR[7].XIC[14].icell.PDM VPWR 0.0118f
C3849 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.Ien 0.04854f
C3850 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.PDM 0.02104f
C3851 XA.Cn[1] XA.XIR[15].XIC[1].icell.PDM 0.02601f
C3852 XThR.Tn[2] XA.XIR[2].XIC[6].icell.Ien 0.14211f
C3853 XA.Cn[0] XA.XIR[5].XIC[0].icell.Ien 0.04604f
C3854 thermo15c_0.XTB6.Y XA.Cn[7] 0.01474f
C3855 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.PDM 0.02104f
C3856 XA.XIR[4].XIC[5].icell.Ien VPWR 0.18829f
C3857 XA.Cn[11] XA.XIR[0].XIC[11].icell.PDM 0.0279f
C3858 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.Ien 0.04854f
C3859 XA.Cn[11] XA.XIR[9].XIC[11].icell.Ien 0.04604f
C3860 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.PDM 0.02104f
C3861 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3862 XA.XIR[10].XIC[0].icell.Ien Vbias 0.19149f
C3863 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.PDM 0.02104f
C3864 XA.XIR[9].XIC[10].icell.PDM VPWR 0.01171f
C3865 XA.XIR[6].XIC[5].icell.PDM Vbias 0.03928f
C3866 XA.Cn[8] XA.XIR[10].XIC[8].icell.PDM 0.02601f
C3867 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3868 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.Ien 0.04854f
C3869 XA.Cn[2] XA.XIR[2].XIC[2].icell.PDM 0.02602f
C3870 XA.XIR[0].XIC[2].icell.PDM VPWR 0.01132f
C3871 XA.XIR[5].XIC[12].icell.PDM Vbias 0.03928f
C3872 XA.XIR[14].XIC[2].icell.PDM Vbias 0.03928f
C3873 XThR.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.14211f
C3874 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.Ien 0.04854f
C3875 XA.XIR[9].XIC[8].icell.Ien VPWR 0.18829f
C3876 XA.XIR[13].XIC[6].icell.PDM Vbias 0.03928f
C3877 XA.Cn[6] XThR.Tn[14] 0.40738f
C3878 XThR.XTB7.B XThR.XTB7.Y 0.33493f
C3879 thermo15c_0.XTBN.A thermo15c_0.XTB5.Y 0.10854f
C3880 XA.Cn[12] XA.XIR[15].XIC[12].icell.Ien 0.04292f
C3881 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.Ien 0.04854f
C3882 XThR.Tn[9] XA.XIR[9].XIC[4].icell.Ien 0.14211f
C3883 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PDM 0.04035f
C3884 XThR.XTB5.Y a_n1319_6405# 0.01188f
C3885 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.PDM 0.02104f
C3886 a_n1049_5317# VPWR 0.72036f
C3887 XA.Cn[10] VPWR 4.54895f
C3888 XA.XIR[1].XIC_15.icell.PDM VPWR 0.07527f
C3889 thermo15c_0.XTB2.Y thermo15c_0.XTB6.A 0.18237f
C3890 thermo15c_0.XTB5.A thermo15c_0.XTB3.Y 0.01156f
C3891 thermo15c_0.XTB1.Y thermo15c_0.XTB7.A 0.48957f
C3892 thermo15c_0.XTBN.Y XA.Cn[1] 0.49539f
C3893 XA.XIR[4].XIC_15.icell.PDM VPWR 0.07527f
C3894 XA.XIR[7].XIC[4].icell.Ien VPWR 0.18829f
C3895 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.PDM 0.02104f
C3896 XA.Cn[13] XA.XIR[6].XIC[13].icell.PDM 0.02601f
C3897 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.Ien 0.04854f
C3898 XThR.Tn[2] XThR.Tn[3] 0.15335f
C3899 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.PDM 0.02104f
C3900 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3901 XA.Cn[6] XA.XIR[5].XIC[6].icell.Ien 0.04604f
C3902 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout 0.06446f
C3903 XA.XIR[3].XIC[5].icell.Ien Vbias 0.19161f
C3904 XA.Cn[5] XA.XIR[13].XIC[5].icell.PDM 0.02601f
C3905 XA.Cn[10] XA.XIR[13].XIC[10].icell.Ien 0.04604f
C3906 XThR.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.14251f
C3907 XA.XIR[6].XIC_dummy_left.icell.Iout Iout 0.03553f
C3908 thermo15c_0.XTB6.A VPWR 0.68179f
C3909 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PDM 0.04056f
C3910 XA.XIR[3].XIC[7].icell.PDM Vbias 0.03928f
C3911 XA.XIR[4].XIC[14].icell.Ien Vbias 0.19161f
C3912 XA.XIR[8].XIC[9].icell.PDM Vbias 0.03928f
C3913 XThR.XTBN.Y a_n997_715# 0.21503f
C3914 XThR.Tn[7] XA.XIR[7].XIC[1].icell.Ien 0.14211f
C3915 XA.Cn[13] XA.XIR[12].XIC[13].icell.Ien 0.04604f
C3916 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.Ien 0.04854f
C3917 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.PDM 0.02104f
C3918 XA.XIR[2].XIC[13].icell.PDM Vbias 0.03928f
C3919 XA.XIR[8].XIC[8].icell.Ien Vbias 0.19161f
C3920 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PDM 0.04035f
C3921 XThR.Tn[4] XA.XIR[4].XIC[13].icell.Ien 0.14211f
C3922 XA.Cn[8] XA.XIR[2].XIC[8].icell.Ien 0.04605f
C3923 XThR.Tn[0] XA.XIR[0].XIC[5].icell.Ien 0.14211f
C3924 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR 0.01499f
C3925 XA.XIR[10].XIC_15.icell.PDM Vbias 0.03927f
C3926 XThR.Tn[10] XA.XIR[10].XIC[4].icell.Ien 0.14211f
C3927 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.Ien 0.04854f
C3928 XThR.XTB7.B a_n997_2667# 0.02071f
C3929 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PDM 0.04035f
C3930 XA.Cn[9] Vbias 0.79809f
C3931 XA.Cn[2] XA.XIR[7].XIC[2].icell.PDM 0.02601f
C3932 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.PDM 0.02104f
C3933 XA.XIR[5].XIC[0].icell.PDM VPWR 0.01171f
C3934 XA.XIR[5].XIC[9].icell.Ien Iout 0.06801f
C3935 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PDM 0.04035f
C3936 XThR.Tn[7] XA.XIR[7].XIC[6].icell.Ien 0.14211f
C3937 thermo15c_0.XTB3.Y thermo15c_0.XTBN.Y 0.17246f
C3938 XA.XIR[0].XIC[10].icell.Ien Vbias 0.19213f
C3939 a_n1049_6405# VPWR 0.72095f
C3940 XA.Cn[7] XThR.Tn[9] 0.40738f
C3941 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.Ien 0.04854f
C3942 XA.Cn[5] XA.XIR[13].XIC[5].icell.Ien 0.04604f
C3943 XA.XIR[8].XIC_dummy_left.icell.Ien XThR.Tn[8] 0.0125f
C3944 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.Ien 0.04854f
C3945 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.PDM 0.02104f
C3946 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.Ien 0.04854f
C3947 XA.XIR[11].XIC[5].icell.PDM VPWR 0.01171f
C3948 XA.Cn[1] XThR.Tn[13] 0.40738f
C3949 XA.XIR[12].XIC[4].icell.Ien Iout 0.06801f
C3950 data[7] VGND 0.49949f
C3951 data[6] VGND 0.47974f
C3952 data[4] VGND 0.59317f
C3953 data[5] VGND 1.17814f
C3954 Iout VGND 0.32108p
C3955 bias[2] VGND 0.8011f
C3956 bias[0] VGND 2.64942f
C3957 Vbias VGND 0.17035p
C3958 bias[1] VGND 0.72457f
C3959 data[3] VGND 0.49926f
C3960 data[2] VGND 0.48064f
C3961 data[0] VGND 0.59269f
C3962 data[1] VGND 1.17844f
C3963 VPWR VGND 0.37297p
C3964 a_n997_715# VGND 0.5638f
C3965 XA.XIR[15].XIC_dummy_right.icell.Iout VGND 0.7524f
C3966 XA.XIR[15].XIC_dummy_right.icell.SM VGND 0.01013f
C3967 XA.XIR[15].XIC_dummy_right.icell.Ien VGND 0.64532f
C3968 XA.XIR[15].XIC_15.icell.Ien VGND 0.44493f
C3969 XA.XIR[15].XIC[14].icell.Ien VGND 0.4451f
C3970 XA.XIR[15].XIC[13].icell.Ien VGND 0.44506f
C3971 XA.XIR[15].XIC[12].icell.Ien VGND 0.44506f
C3972 XA.XIR[15].XIC[11].icell.Ien VGND 0.44506f
C3973 XA.XIR[15].XIC[10].icell.Ien VGND 0.44506f
C3974 XA.XIR[15].XIC[9].icell.Ien VGND 0.44506f
C3975 XA.XIR[15].XIC[8].icell.Ien VGND 0.44506f
C3976 XA.XIR[15].XIC[7].icell.Ien VGND 0.44506f
C3977 XA.XIR[15].XIC[6].icell.Ien VGND 0.44506f
C3978 XA.XIR[15].XIC[5].icell.Ien VGND 0.44506f
C3979 XA.XIR[15].XIC[4].icell.Ien VGND 0.44506f
C3980 XA.XIR[15].XIC[3].icell.Ien VGND 0.44506f
C3981 XA.XIR[15].XIC[2].icell.Ien VGND 0.44506f
C3982 XA.XIR[15].XIC_dummy_left.icell.Iout VGND 0.70682f
C3983 XA.XIR[15].XIC[1].icell.Ien VGND 0.44506f
C3984 XA.XIR[15].XIC[0].icell.Ien VGND 0.44521f
C3985 XA.XIR[15].XIC_dummy_left.icell.SM VGND 0.01033f
C3986 XA.XIR[15].XIC_dummy_left.icell.Ien VGND 0.6116f
C3987 XA.XIR[15].XIC_dummy_right.icell.PDM VGND 0.23278f
C3988 XA.XIR[15].XIC_15.icell.PDM VGND 0.18786f
C3989 XA.XIR[15].XIC[14].icell.PDM VGND 0.18744f
C3990 XA.XIR[15].XIC[13].icell.PDM VGND 0.18744f
C3991 XA.XIR[15].XIC[12].icell.PDM VGND 0.18744f
C3992 XA.XIR[15].XIC[11].icell.PDM VGND 0.18744f
C3993 XA.XIR[15].XIC[10].icell.PDM VGND 0.18744f
C3994 XA.XIR[15].XIC[9].icell.PDM VGND 0.18744f
C3995 XA.XIR[15].XIC[8].icell.PDM VGND 0.18744f
C3996 XA.XIR[15].XIC[7].icell.PDM VGND 0.18744f
C3997 XA.XIR[15].XIC[6].icell.PDM VGND 0.18744f
C3998 XA.XIR[15].XIC[5].icell.PDM VGND 0.18744f
C3999 XA.XIR[15].XIC[4].icell.PDM VGND 0.18744f
C4000 XA.XIR[15].XIC[3].icell.PDM VGND 0.18744f
C4001 XA.XIR[15].XIC[2].icell.PDM VGND 0.18744f
C4002 XA.XIR[15].XIC[1].icell.PDM VGND 0.18744f
C4003 XA.XIR[15].XIC[0].icell.PDM VGND 0.1876f
C4004 XA.XIR[15].XIC_dummy_left.icell.PDM VGND 0.22703f
C4005 XA.XIR[14].XIC_dummy_right.icell.Iout VGND 0.85788f
C4006 XA.XIR[14].XIC_dummy_right.icell.SM VGND 0.01013f
C4007 XA.XIR[14].XIC_dummy_right.icell.Ien VGND 0.60818f
C4008 XA.XIR[14].XIC_15.icell.Ien VGND 0.37264f
C4009 XA.XIR[14].XIC[14].icell.Ien VGND 0.37333f
C4010 XA.XIR[14].XIC[13].icell.Ien VGND 0.3733f
C4011 XA.XIR[14].XIC[12].icell.Ien VGND 0.3733f
C4012 XA.XIR[14].XIC[11].icell.Ien VGND 0.3733f
C4013 XA.XIR[14].XIC[10].icell.Ien VGND 0.3733f
C4014 XA.XIR[14].XIC[9].icell.Ien VGND 0.3733f
C4015 XA.XIR[14].XIC[8].icell.Ien VGND 0.3733f
C4016 XA.XIR[14].XIC[7].icell.Ien VGND 0.3733f
C4017 XA.XIR[14].XIC[6].icell.Ien VGND 0.3733f
C4018 XA.XIR[14].XIC[5].icell.Ien VGND 0.3733f
C4019 XA.XIR[14].XIC[4].icell.Ien VGND 0.3733f
C4020 XA.XIR[14].XIC[3].icell.Ien VGND 0.3733f
C4021 XA.XIR[14].XIC[2].icell.Ien VGND 0.3733f
C4022 XA.XIR[14].XIC_dummy_left.icell.Iout VGND 0.8066f
C4023 XThR.Tn[14] VGND 13.06755f
C4024 XA.XIR[14].XIC[1].icell.Ien VGND 0.3733f
C4025 a_n997_1579# VGND 0.54776f
C4026 XA.XIR[14].XIC[0].icell.Ien VGND 0.37345f
C4027 XA.XIR[14].XIC_dummy_left.icell.SM VGND 0.01033f
C4028 XA.XIR[14].XIC_dummy_left.icell.Ien VGND 0.57576f
C4029 a_n997_1803# VGND 0.53619f
C4030 XA.XIR[14].XIC_dummy_right.icell.PDM VGND 0.23384f
C4031 XA.XIR[14].XIC_15.icell.PDM VGND 0.18862f
C4032 XA.XIR[14].XIC[14].icell.PDM VGND 0.1882f
C4033 XA.XIR[14].XIC[13].icell.PDM VGND 0.1882f
C4034 XA.XIR[14].XIC[12].icell.PDM VGND 0.1882f
C4035 XA.XIR[14].XIC[11].icell.PDM VGND 0.1882f
C4036 XA.XIR[14].XIC[10].icell.PDM VGND 0.1882f
C4037 XA.XIR[14].XIC[9].icell.PDM VGND 0.1882f
C4038 XA.XIR[14].XIC[8].icell.PDM VGND 0.1882f
C4039 XA.XIR[14].XIC[7].icell.PDM VGND 0.1882f
C4040 XA.XIR[14].XIC[6].icell.PDM VGND 0.1882f
C4041 XA.XIR[14].XIC[5].icell.PDM VGND 0.1882f
C4042 XA.XIR[14].XIC[4].icell.PDM VGND 0.1882f
C4043 XA.XIR[14].XIC[3].icell.PDM VGND 0.1882f
C4044 XA.XIR[14].XIC[2].icell.PDM VGND 0.1882f
C4045 XA.XIR[14].XIC[1].icell.PDM VGND 0.1882f
C4046 XA.XIR[14].XIC[0].icell.PDM VGND 0.18836f
C4047 XA.XIR[14].XIC_dummy_left.icell.PDM VGND 0.22809f
C4048 XA.XIR[13].XIC_dummy_right.icell.Iout VGND 0.85788f
C4049 XA.XIR[13].XIC_dummy_right.icell.SM VGND 0.01013f
C4050 XA.XIR[13].XIC_dummy_right.icell.Ien VGND 0.60818f
C4051 XA.XIR[13].XIC_15.icell.Ien VGND 0.37264f
C4052 XA.XIR[13].XIC[14].icell.Ien VGND 0.37333f
C4053 XA.XIR[13].XIC[13].icell.Ien VGND 0.3733f
C4054 XA.XIR[13].XIC[12].icell.Ien VGND 0.3733f
C4055 XA.XIR[13].XIC[11].icell.Ien VGND 0.3733f
C4056 XA.XIR[13].XIC[10].icell.Ien VGND 0.3733f
C4057 XA.XIR[13].XIC[9].icell.Ien VGND 0.3733f
C4058 XA.XIR[13].XIC[8].icell.Ien VGND 0.3733f
C4059 XA.XIR[13].XIC[7].icell.Ien VGND 0.3733f
C4060 XA.XIR[13].XIC[6].icell.Ien VGND 0.3733f
C4061 XA.XIR[13].XIC[5].icell.Ien VGND 0.3733f
C4062 XA.XIR[13].XIC[4].icell.Ien VGND 0.3733f
C4063 XA.XIR[13].XIC[3].icell.Ien VGND 0.3733f
C4064 XA.XIR[13].XIC[2].icell.Ien VGND 0.3733f
C4065 XA.XIR[13].XIC_dummy_left.icell.Iout VGND 0.80664f
C4066 XThR.Tn[13] VGND 12.91167f
C4067 XA.XIR[13].XIC[1].icell.Ien VGND 0.3733f
C4068 XA.XIR[13].XIC[0].icell.Ien VGND 0.37345f
C4069 XA.XIR[13].XIC_dummy_left.icell.SM VGND 0.01033f
C4070 XA.XIR[13].XIC_dummy_left.icell.Ien VGND 0.57422f
C4071 XA.XIR[13].XIC_dummy_right.icell.PDM VGND 0.23384f
C4072 XA.XIR[13].XIC_15.icell.PDM VGND 0.18862f
C4073 XA.XIR[13].XIC[14].icell.PDM VGND 0.1882f
C4074 XA.XIR[13].XIC[13].icell.PDM VGND 0.1882f
C4075 XA.XIR[13].XIC[12].icell.PDM VGND 0.1882f
C4076 XA.XIR[13].XIC[11].icell.PDM VGND 0.1882f
C4077 XA.XIR[13].XIC[10].icell.PDM VGND 0.1882f
C4078 XA.XIR[13].XIC[9].icell.PDM VGND 0.1882f
C4079 XA.XIR[13].XIC[8].icell.PDM VGND 0.1882f
C4080 XA.XIR[13].XIC[7].icell.PDM VGND 0.1882f
C4081 XA.XIR[13].XIC[6].icell.PDM VGND 0.1882f
C4082 XA.XIR[13].XIC[5].icell.PDM VGND 0.1882f
C4083 XA.XIR[13].XIC[4].icell.PDM VGND 0.1882f
C4084 XA.XIR[13].XIC[3].icell.PDM VGND 0.1882f
C4085 XA.XIR[13].XIC[2].icell.PDM VGND 0.1882f
C4086 XA.XIR[13].XIC[1].icell.PDM VGND 0.1882f
C4087 XA.XIR[13].XIC[0].icell.PDM VGND 0.18836f
C4088 XA.XIR[13].XIC_dummy_left.icell.PDM VGND 0.22809f
C4089 XA.XIR[12].XIC_dummy_right.icell.Iout VGND 0.85788f
C4090 XA.XIR[12].XIC_dummy_right.icell.SM VGND 0.01013f
C4091 XA.XIR[12].XIC_dummy_right.icell.Ien VGND 0.60818f
C4092 XA.XIR[12].XIC_15.icell.Ien VGND 0.37264f
C4093 XA.XIR[12].XIC[14].icell.Ien VGND 0.37333f
C4094 XA.XIR[12].XIC[13].icell.Ien VGND 0.3733f
C4095 XA.XIR[12].XIC[12].icell.Ien VGND 0.3733f
C4096 XA.XIR[12].XIC[11].icell.Ien VGND 0.3733f
C4097 XA.XIR[12].XIC[10].icell.Ien VGND 0.3733f
C4098 XA.XIR[12].XIC[9].icell.Ien VGND 0.3733f
C4099 XA.XIR[12].XIC[8].icell.Ien VGND 0.3733f
C4100 XA.XIR[12].XIC[7].icell.Ien VGND 0.3733f
C4101 XA.XIR[12].XIC[6].icell.Ien VGND 0.3733f
C4102 XA.XIR[12].XIC[5].icell.Ien VGND 0.3733f
C4103 XA.XIR[12].XIC[4].icell.Ien VGND 0.3733f
C4104 XA.XIR[12].XIC[3].icell.Ien VGND 0.3733f
C4105 XA.XIR[12].XIC[2].icell.Ien VGND 0.3733f
C4106 XA.XIR[12].XIC_dummy_left.icell.Iout VGND 0.80529f
C4107 XThR.Tn[12] VGND 12.80173f
C4108 XA.XIR[12].XIC[1].icell.Ien VGND 0.3733f
C4109 XA.XIR[12].XIC[0].icell.Ien VGND 0.37345f
C4110 XA.XIR[12].XIC_dummy_left.icell.SM VGND 0.01033f
C4111 XA.XIR[12].XIC_dummy_left.icell.Ien VGND 0.5728f
C4112 a_n997_2667# VGND 0.5457f
C4113 XA.XIR[12].XIC_dummy_right.icell.PDM VGND 0.23384f
C4114 XA.XIR[12].XIC_15.icell.PDM VGND 0.18862f
C4115 XA.XIR[12].XIC[14].icell.PDM VGND 0.1882f
C4116 XA.XIR[12].XIC[13].icell.PDM VGND 0.1882f
C4117 XA.XIR[12].XIC[12].icell.PDM VGND 0.1882f
C4118 XA.XIR[12].XIC[11].icell.PDM VGND 0.1882f
C4119 XA.XIR[12].XIC[10].icell.PDM VGND 0.1882f
C4120 XA.XIR[12].XIC[9].icell.PDM VGND 0.1882f
C4121 XA.XIR[12].XIC[8].icell.PDM VGND 0.1882f
C4122 XA.XIR[12].XIC[7].icell.PDM VGND 0.1882f
C4123 XA.XIR[12].XIC[6].icell.PDM VGND 0.1882f
C4124 XA.XIR[12].XIC[5].icell.PDM VGND 0.1882f
C4125 XA.XIR[12].XIC[4].icell.PDM VGND 0.1882f
C4126 XA.XIR[12].XIC[3].icell.PDM VGND 0.1882f
C4127 XA.XIR[12].XIC[2].icell.PDM VGND 0.1882f
C4128 XA.XIR[12].XIC[1].icell.PDM VGND 0.1882f
C4129 XA.XIR[12].XIC[0].icell.PDM VGND 0.18836f
C4130 XA.XIR[12].XIC_dummy_left.icell.PDM VGND 0.22809f
C4131 XA.XIR[11].XIC_dummy_right.icell.Iout VGND 0.85788f
C4132 XA.XIR[11].XIC_dummy_right.icell.SM VGND 0.01013f
C4133 XA.XIR[11].XIC_dummy_right.icell.Ien VGND 0.60818f
C4134 XA.XIR[11].XIC_15.icell.Ien VGND 0.37264f
C4135 XA.XIR[11].XIC[14].icell.Ien VGND 0.37333f
C4136 XA.XIR[11].XIC[13].icell.Ien VGND 0.3733f
C4137 XA.XIR[11].XIC[12].icell.Ien VGND 0.3733f
C4138 XA.XIR[11].XIC[11].icell.Ien VGND 0.3733f
C4139 XA.XIR[11].XIC[10].icell.Ien VGND 0.3733f
C4140 XA.XIR[11].XIC[9].icell.Ien VGND 0.3733f
C4141 XA.XIR[11].XIC[8].icell.Ien VGND 0.3733f
C4142 XA.XIR[11].XIC[7].icell.Ien VGND 0.3733f
C4143 XA.XIR[11].XIC[6].icell.Ien VGND 0.3733f
C4144 XA.XIR[11].XIC[5].icell.Ien VGND 0.3733f
C4145 XA.XIR[11].XIC[4].icell.Ien VGND 0.3733f
C4146 XA.XIR[11].XIC[3].icell.Ien VGND 0.3733f
C4147 XA.XIR[11].XIC[2].icell.Ien VGND 0.3733f
C4148 XA.XIR[11].XIC_dummy_left.icell.Iout VGND 0.80765f
C4149 XThR.Tn[11] VGND 12.86402f
C4150 XA.XIR[11].XIC[1].icell.Ien VGND 0.3733f
C4151 a_n997_2891# VGND 0.54795f
C4152 XA.XIR[11].XIC[0].icell.Ien VGND 0.37345f
C4153 XA.XIR[11].XIC_dummy_left.icell.SM VGND 0.01033f
C4154 XA.XIR[11].XIC_dummy_left.icell.Ien VGND 0.57294f
C4155 XA.XIR[11].XIC_dummy_right.icell.PDM VGND 0.23384f
C4156 XA.XIR[11].XIC_15.icell.PDM VGND 0.18862f
C4157 XA.XIR[11].XIC[14].icell.PDM VGND 0.1882f
C4158 XA.XIR[11].XIC[13].icell.PDM VGND 0.1882f
C4159 XA.XIR[11].XIC[12].icell.PDM VGND 0.1882f
C4160 XA.XIR[11].XIC[11].icell.PDM VGND 0.1882f
C4161 XA.XIR[11].XIC[10].icell.PDM VGND 0.1882f
C4162 XA.XIR[11].XIC[9].icell.PDM VGND 0.1882f
C4163 XA.XIR[11].XIC[8].icell.PDM VGND 0.1882f
C4164 XA.XIR[11].XIC[7].icell.PDM VGND 0.1882f
C4165 XA.XIR[11].XIC[6].icell.PDM VGND 0.1882f
C4166 XA.XIR[11].XIC[5].icell.PDM VGND 0.1882f
C4167 XA.XIR[11].XIC[4].icell.PDM VGND 0.1882f
C4168 XA.XIR[11].XIC[3].icell.PDM VGND 0.1882f
C4169 XA.XIR[11].XIC[2].icell.PDM VGND 0.1882f
C4170 XA.XIR[11].XIC[1].icell.PDM VGND 0.1882f
C4171 XA.XIR[11].XIC[0].icell.PDM VGND 0.18836f
C4172 XA.XIR[11].XIC_dummy_left.icell.PDM VGND 0.22809f
C4173 XA.XIR[10].XIC_dummy_right.icell.Iout VGND 0.85788f
C4174 XA.XIR[10].XIC_dummy_right.icell.SM VGND 0.01013f
C4175 XA.XIR[10].XIC_dummy_right.icell.Ien VGND 0.60818f
C4176 XA.XIR[10].XIC_15.icell.Ien VGND 0.37264f
C4177 XA.XIR[10].XIC[14].icell.Ien VGND 0.37333f
C4178 XA.XIR[10].XIC[13].icell.Ien VGND 0.3733f
C4179 XA.XIR[10].XIC[12].icell.Ien VGND 0.3733f
C4180 XA.XIR[10].XIC[11].icell.Ien VGND 0.3733f
C4181 XA.XIR[10].XIC[10].icell.Ien VGND 0.3733f
C4182 XA.XIR[10].XIC[9].icell.Ien VGND 0.3733f
C4183 XA.XIR[10].XIC[8].icell.Ien VGND 0.3733f
C4184 XA.XIR[10].XIC[7].icell.Ien VGND 0.3733f
C4185 XA.XIR[10].XIC[6].icell.Ien VGND 0.3733f
C4186 XA.XIR[10].XIC[5].icell.Ien VGND 0.3733f
C4187 XA.XIR[10].XIC[4].icell.Ien VGND 0.3733f
C4188 XA.XIR[10].XIC[3].icell.Ien VGND 0.3733f
C4189 XA.XIR[10].XIC[2].icell.Ien VGND 0.3733f
C4190 XA.XIR[10].XIC_dummy_left.icell.Iout VGND 0.80648f
C4191 XThR.Tn[10] VGND 12.83941f
C4192 XA.XIR[10].XIC[1].icell.Ien VGND 0.3733f
C4193 XA.XIR[10].XIC[0].icell.Ien VGND 0.37345f
C4194 XA.XIR[10].XIC_dummy_left.icell.SM VGND 0.01033f
C4195 XA.XIR[10].XIC_dummy_left.icell.Ien VGND 0.57422f
C4196 XA.XIR[10].XIC_dummy_right.icell.PDM VGND 0.23384f
C4197 XA.XIR[10].XIC_15.icell.PDM VGND 0.18862f
C4198 XA.XIR[10].XIC[14].icell.PDM VGND 0.1882f
C4199 XA.XIR[10].XIC[13].icell.PDM VGND 0.1882f
C4200 XA.XIR[10].XIC[12].icell.PDM VGND 0.1882f
C4201 XA.XIR[10].XIC[11].icell.PDM VGND 0.1882f
C4202 XA.XIR[10].XIC[10].icell.PDM VGND 0.1882f
C4203 XA.XIR[10].XIC[9].icell.PDM VGND 0.1882f
C4204 XA.XIR[10].XIC[8].icell.PDM VGND 0.1882f
C4205 XA.XIR[10].XIC[7].icell.PDM VGND 0.1882f
C4206 XA.XIR[10].XIC[6].icell.PDM VGND 0.1882f
C4207 XA.XIR[10].XIC[5].icell.PDM VGND 0.1882f
C4208 XA.XIR[10].XIC[4].icell.PDM VGND 0.1882f
C4209 XA.XIR[10].XIC[3].icell.PDM VGND 0.1882f
C4210 XA.XIR[10].XIC[2].icell.PDM VGND 0.1882f
C4211 XA.XIR[10].XIC[1].icell.PDM VGND 0.1882f
C4212 XA.XIR[10].XIC[0].icell.PDM VGND 0.18836f
C4213 XA.XIR[10].XIC_dummy_left.icell.PDM VGND 0.22809f
C4214 XA.XIR[9].XIC_dummy_right.icell.Iout VGND 0.85788f
C4215 XA.XIR[9].XIC_dummy_right.icell.SM VGND 0.01013f
C4216 XA.XIR[9].XIC_dummy_right.icell.Ien VGND 0.60818f
C4217 XA.XIR[9].XIC_15.icell.Ien VGND 0.37264f
C4218 XA.XIR[9].XIC[14].icell.Ien VGND 0.37333f
C4219 XA.XIR[9].XIC[13].icell.Ien VGND 0.3733f
C4220 XA.XIR[9].XIC[12].icell.Ien VGND 0.3733f
C4221 XA.XIR[9].XIC[11].icell.Ien VGND 0.3733f
C4222 XA.XIR[9].XIC[10].icell.Ien VGND 0.3733f
C4223 XA.XIR[9].XIC[9].icell.Ien VGND 0.3733f
C4224 XA.XIR[9].XIC[8].icell.Ien VGND 0.3733f
C4225 XA.XIR[9].XIC[7].icell.Ien VGND 0.3733f
C4226 XA.XIR[9].XIC[6].icell.Ien VGND 0.3733f
C4227 XA.XIR[9].XIC[5].icell.Ien VGND 0.3733f
C4228 XA.XIR[9].XIC[4].icell.Ien VGND 0.3733f
C4229 XA.XIR[9].XIC[3].icell.Ien VGND 0.3733f
C4230 XA.XIR[9].XIC[2].icell.Ien VGND 0.3733f
C4231 XA.XIR[9].XIC_dummy_left.icell.Iout VGND 0.80834f
C4232 XA.XIR[9].XIC[1].icell.Ien VGND 0.3733f
C4233 XThR.Tn[9] VGND 12.8472f
C4234 a_n997_3755# VGND 0.54861f
C4235 XA.XIR[9].XIC[0].icell.Ien VGND 0.37345f
C4236 XA.XIR[9].XIC_dummy_left.icell.SM VGND 0.01033f
C4237 XA.XIR[9].XIC_dummy_left.icell.Ien VGND 0.5732f
C4238 a_n997_3979# VGND 0.54721f
C4239 XA.XIR[9].XIC_dummy_right.icell.PDM VGND 0.23384f
C4240 XA.XIR[9].XIC_15.icell.PDM VGND 0.18862f
C4241 XA.XIR[9].XIC[14].icell.PDM VGND 0.1882f
C4242 XA.XIR[9].XIC[13].icell.PDM VGND 0.1882f
C4243 XA.XIR[9].XIC[12].icell.PDM VGND 0.1882f
C4244 XA.XIR[9].XIC[11].icell.PDM VGND 0.1882f
C4245 XA.XIR[9].XIC[10].icell.PDM VGND 0.1882f
C4246 XA.XIR[9].XIC[9].icell.PDM VGND 0.1882f
C4247 XA.XIR[9].XIC[8].icell.PDM VGND 0.1882f
C4248 XA.XIR[9].XIC[7].icell.PDM VGND 0.1882f
C4249 XA.XIR[9].XIC[6].icell.PDM VGND 0.1882f
C4250 XA.XIR[9].XIC[5].icell.PDM VGND 0.1882f
C4251 XA.XIR[9].XIC[4].icell.PDM VGND 0.1882f
C4252 XA.XIR[9].XIC[3].icell.PDM VGND 0.1882f
C4253 XA.XIR[9].XIC[2].icell.PDM VGND 0.1882f
C4254 XA.XIR[9].XIC[1].icell.PDM VGND 0.1882f
C4255 XA.XIR[9].XIC[0].icell.PDM VGND 0.18836f
C4256 XA.XIR[9].XIC_dummy_left.icell.PDM VGND 0.22809f
C4257 XA.XIR[8].XIC_dummy_right.icell.Iout VGND 0.85788f
C4258 XA.XIR[8].XIC_dummy_right.icell.SM VGND 0.01013f
C4259 XA.XIR[8].XIC_dummy_right.icell.Ien VGND 0.60818f
C4260 XA.XIR[8].XIC_15.icell.Ien VGND 0.37264f
C4261 XA.XIR[8].XIC[14].icell.Ien VGND 0.37333f
C4262 XA.XIR[8].XIC[13].icell.Ien VGND 0.3733f
C4263 XA.XIR[8].XIC[12].icell.Ien VGND 0.3733f
C4264 XA.XIR[8].XIC[11].icell.Ien VGND 0.3733f
C4265 XA.XIR[8].XIC[10].icell.Ien VGND 0.3733f
C4266 XA.XIR[8].XIC[9].icell.Ien VGND 0.3733f
C4267 XA.XIR[8].XIC[8].icell.Ien VGND 0.3733f
C4268 XA.XIR[8].XIC[7].icell.Ien VGND 0.3733f
C4269 XA.XIR[8].XIC[6].icell.Ien VGND 0.3733f
C4270 XA.XIR[8].XIC[5].icell.Ien VGND 0.3733f
C4271 XA.XIR[8].XIC[4].icell.Ien VGND 0.3733f
C4272 XA.XIR[8].XIC[3].icell.Ien VGND 0.3733f
C4273 XA.XIR[8].XIC[2].icell.Ien VGND 0.3733f
C4274 XA.XIR[8].XIC_dummy_left.icell.Iout VGND 0.80566f
C4275 XA.XIR[8].XIC[1].icell.Ien VGND 0.3733f
C4276 XThR.Tn[8] VGND 12.78722f
C4277 XA.XIR[8].XIC[0].icell.Ien VGND 0.37345f
C4278 XA.XIR[8].XIC_dummy_left.icell.SM VGND 0.01033f
C4279 XA.XIR[8].XIC_dummy_left.icell.Ien VGND 0.57308f
C4280 XA.XIR[8].XIC_dummy_right.icell.PDM VGND 0.23384f
C4281 XA.XIR[8].XIC_15.icell.PDM VGND 0.18862f
C4282 XA.XIR[8].XIC[14].icell.PDM VGND 0.1882f
C4283 XA.XIR[8].XIC[13].icell.PDM VGND 0.1882f
C4284 XA.XIR[8].XIC[12].icell.PDM VGND 0.1882f
C4285 XA.XIR[8].XIC[11].icell.PDM VGND 0.1882f
C4286 XA.XIR[8].XIC[10].icell.PDM VGND 0.1882f
C4287 XA.XIR[8].XIC[9].icell.PDM VGND 0.1882f
C4288 XA.XIR[8].XIC[8].icell.PDM VGND 0.1882f
C4289 XA.XIR[8].XIC[7].icell.PDM VGND 0.1882f
C4290 XA.XIR[8].XIC[6].icell.PDM VGND 0.1882f
C4291 XA.XIR[8].XIC[5].icell.PDM VGND 0.1882f
C4292 XA.XIR[8].XIC[4].icell.PDM VGND 0.1882f
C4293 XA.XIR[8].XIC[3].icell.PDM VGND 0.1882f
C4294 XA.XIR[8].XIC[2].icell.PDM VGND 0.1882f
C4295 XA.XIR[8].XIC[1].icell.PDM VGND 0.1882f
C4296 XA.XIR[8].XIC[0].icell.PDM VGND 0.18836f
C4297 XA.XIR[8].XIC_dummy_left.icell.PDM VGND 0.22809f
C4298 XA.XIR[7].XIC_dummy_right.icell.Iout VGND 0.85788f
C4299 XA.XIR[7].XIC_dummy_right.icell.SM VGND 0.01013f
C4300 XA.XIR[7].XIC_dummy_right.icell.Ien VGND 0.60818f
C4301 XA.XIR[7].XIC_15.icell.Ien VGND 0.37264f
C4302 XA.XIR[7].XIC[14].icell.Ien VGND 0.37333f
C4303 XA.XIR[7].XIC[13].icell.Ien VGND 0.3733f
C4304 XA.XIR[7].XIC[12].icell.Ien VGND 0.3733f
C4305 XA.XIR[7].XIC[11].icell.Ien VGND 0.3733f
C4306 XA.XIR[7].XIC[10].icell.Ien VGND 0.3733f
C4307 XA.XIR[7].XIC[9].icell.Ien VGND 0.3733f
C4308 XA.XIR[7].XIC[8].icell.Ien VGND 0.3733f
C4309 XA.XIR[7].XIC[7].icell.Ien VGND 0.3733f
C4310 XA.XIR[7].XIC[6].icell.Ien VGND 0.3733f
C4311 XA.XIR[7].XIC[5].icell.Ien VGND 0.3733f
C4312 XA.XIR[7].XIC[4].icell.Ien VGND 0.3733f
C4313 XA.XIR[7].XIC[3].icell.Ien VGND 0.3733f
C4314 XA.XIR[7].XIC[2].icell.Ien VGND 0.3733f
C4315 XA.XIR[7].XIC_dummy_left.icell.Iout VGND 0.80598f
C4316 XA.XIR[7].XIC[1].icell.Ien VGND 0.3733f
C4317 XA.XIR[7].XIC[0].icell.Ien VGND 0.37345f
C4318 XA.XIR[7].XIC_dummy_left.icell.SM VGND 0.01033f
C4319 XThR.Tn[7] VGND 13.23029f
C4320 XThR.XTBN.A VGND 1.22814f
C4321 XA.XIR[7].XIC_dummy_left.icell.Ien VGND 0.57576f
C4322 XA.XIR[7].XIC_dummy_right.icell.PDM VGND 0.23384f
C4323 XA.XIR[7].XIC_15.icell.PDM VGND 0.18862f
C4324 XA.XIR[7].XIC[14].icell.PDM VGND 0.1882f
C4325 XA.XIR[7].XIC[13].icell.PDM VGND 0.1882f
C4326 XA.XIR[7].XIC[12].icell.PDM VGND 0.1882f
C4327 XA.XIR[7].XIC[11].icell.PDM VGND 0.1882f
C4328 XA.XIR[7].XIC[10].icell.PDM VGND 0.1882f
C4329 XA.XIR[7].XIC[9].icell.PDM VGND 0.1882f
C4330 XA.XIR[7].XIC[8].icell.PDM VGND 0.1882f
C4331 XA.XIR[7].XIC[7].icell.PDM VGND 0.1882f
C4332 XA.XIR[7].XIC[6].icell.PDM VGND 0.1882f
C4333 XA.XIR[7].XIC[5].icell.PDM VGND 0.1882f
C4334 XA.XIR[7].XIC[4].icell.PDM VGND 0.1882f
C4335 XA.XIR[7].XIC[3].icell.PDM VGND 0.1882f
C4336 XA.XIR[7].XIC[2].icell.PDM VGND 0.1882f
C4337 XA.XIR[7].XIC[1].icell.PDM VGND 0.1882f
C4338 XA.XIR[7].XIC[0].icell.PDM VGND 0.18836f
C4339 XA.XIR[7].XIC_dummy_left.icell.PDM VGND 0.22809f
C4340 XA.XIR[6].XIC_dummy_right.icell.Iout VGND 0.85788f
C4341 XA.XIR[6].XIC_dummy_right.icell.SM VGND 0.01013f
C4342 XA.XIR[6].XIC_dummy_right.icell.Ien VGND 0.60818f
C4343 XA.XIR[6].XIC_15.icell.Ien VGND 0.37264f
C4344 XA.XIR[6].XIC[14].icell.Ien VGND 0.37333f
C4345 XA.XIR[6].XIC[13].icell.Ien VGND 0.3733f
C4346 XA.XIR[6].XIC[12].icell.Ien VGND 0.3733f
C4347 XA.XIR[6].XIC[11].icell.Ien VGND 0.3733f
C4348 XA.XIR[6].XIC[10].icell.Ien VGND 0.3733f
C4349 XA.XIR[6].XIC[9].icell.Ien VGND 0.3733f
C4350 XA.XIR[6].XIC[8].icell.Ien VGND 0.3733f
C4351 XA.XIR[6].XIC[7].icell.Ien VGND 0.3733f
C4352 XA.XIR[6].XIC[6].icell.Ien VGND 0.3733f
C4353 XA.XIR[6].XIC[5].icell.Ien VGND 0.3733f
C4354 XA.XIR[6].XIC[4].icell.Ien VGND 0.3733f
C4355 XA.XIR[6].XIC[3].icell.Ien VGND 0.3733f
C4356 XA.XIR[6].XIC[2].icell.Ien VGND 0.3733f
C4357 XA.XIR[6].XIC_dummy_left.icell.Iout VGND 0.80693f
C4358 XA.XIR[6].XIC[1].icell.Ien VGND 0.3733f
C4359 XA.XIR[6].XIC[0].icell.Ien VGND 0.37345f
C4360 XA.XIR[6].XIC_dummy_left.icell.SM VGND 0.01033f
C4361 XA.XIR[6].XIC_dummy_left.icell.Ien VGND 0.57422f
C4362 XThR.Tn[6] VGND 12.9018f
C4363 a_n1049_5317# VGND 0.02283f
C4364 XThR.XTB7.Y VGND 1.36132f
C4365 XA.XIR[6].XIC_dummy_right.icell.PDM VGND 0.23384f
C4366 XA.XIR[6].XIC_15.icell.PDM VGND 0.18862f
C4367 XA.XIR[6].XIC[14].icell.PDM VGND 0.1882f
C4368 XA.XIR[6].XIC[13].icell.PDM VGND 0.1882f
C4369 XA.XIR[6].XIC[12].icell.PDM VGND 0.1882f
C4370 XA.XIR[6].XIC[11].icell.PDM VGND 0.1882f
C4371 XA.XIR[6].XIC[10].icell.PDM VGND 0.1882f
C4372 XA.XIR[6].XIC[9].icell.PDM VGND 0.1882f
C4373 XA.XIR[6].XIC[8].icell.PDM VGND 0.1882f
C4374 XA.XIR[6].XIC[7].icell.PDM VGND 0.1882f
C4375 XA.XIR[6].XIC[6].icell.PDM VGND 0.1882f
C4376 XA.XIR[6].XIC[5].icell.PDM VGND 0.1882f
C4377 XA.XIR[6].XIC[4].icell.PDM VGND 0.1882f
C4378 XA.XIR[6].XIC[3].icell.PDM VGND 0.1882f
C4379 XA.XIR[6].XIC[2].icell.PDM VGND 0.1882f
C4380 XA.XIR[6].XIC[1].icell.PDM VGND 0.1882f
C4381 XA.XIR[6].XIC[0].icell.PDM VGND 0.18836f
C4382 XA.XIR[6].XIC_dummy_left.icell.PDM VGND 0.22809f
C4383 XA.XIR[5].XIC_dummy_right.icell.Iout VGND 0.85788f
C4384 XA.XIR[5].XIC_dummy_right.icell.SM VGND 0.01013f
C4385 XA.XIR[5].XIC_dummy_right.icell.Ien VGND 0.60818f
C4386 XA.XIR[5].XIC_15.icell.Ien VGND 0.37264f
C4387 XA.XIR[5].XIC[14].icell.Ien VGND 0.37333f
C4388 XA.XIR[5].XIC[13].icell.Ien VGND 0.3733f
C4389 XA.XIR[5].XIC[12].icell.Ien VGND 0.3733f
C4390 XA.XIR[5].XIC[11].icell.Ien VGND 0.3733f
C4391 XA.XIR[5].XIC[10].icell.Ien VGND 0.3733f
C4392 XA.XIR[5].XIC[9].icell.Ien VGND 0.3733f
C4393 XA.XIR[5].XIC[8].icell.Ien VGND 0.3733f
C4394 XA.XIR[5].XIC[7].icell.Ien VGND 0.3733f
C4395 XA.XIR[5].XIC[6].icell.Ien VGND 0.3733f
C4396 XA.XIR[5].XIC[5].icell.Ien VGND 0.3733f
C4397 XA.XIR[5].XIC[4].icell.Ien VGND 0.3733f
C4398 XA.XIR[5].XIC[3].icell.Ien VGND 0.3733f
C4399 XA.XIR[5].XIC[2].icell.Ien VGND 0.3733f
C4400 XA.XIR[5].XIC_dummy_left.icell.Iout VGND 0.80562f
C4401 XA.XIR[5].XIC[1].icell.Ien VGND 0.3733f
C4402 a_n1049_5611# VGND 0.02888f
C4403 XA.XIR[5].XIC[0].icell.Ien VGND 0.37345f
C4404 XA.XIR[5].XIC_dummy_left.icell.SM VGND 0.01033f
C4405 XA.XIR[5].XIC_dummy_left.icell.Ien VGND 0.57288f
C4406 XThR.Tn[5] VGND 12.89248f
C4407 XThR.XTB6.Y VGND 1.38212f
C4408 XA.XIR[5].XIC_dummy_right.icell.PDM VGND 0.23384f
C4409 XA.XIR[5].XIC_15.icell.PDM VGND 0.18862f
C4410 XA.XIR[5].XIC[14].icell.PDM VGND 0.1882f
C4411 XA.XIR[5].XIC[13].icell.PDM VGND 0.1882f
C4412 XA.XIR[5].XIC[12].icell.PDM VGND 0.1882f
C4413 XA.XIR[5].XIC[11].icell.PDM VGND 0.1882f
C4414 XA.XIR[5].XIC[10].icell.PDM VGND 0.1882f
C4415 XA.XIR[5].XIC[9].icell.PDM VGND 0.1882f
C4416 XA.XIR[5].XIC[8].icell.PDM VGND 0.1882f
C4417 XA.XIR[5].XIC[7].icell.PDM VGND 0.1882f
C4418 XA.XIR[5].XIC[6].icell.PDM VGND 0.1882f
C4419 XA.XIR[5].XIC[5].icell.PDM VGND 0.1882f
C4420 XA.XIR[5].XIC[4].icell.PDM VGND 0.1882f
C4421 XA.XIR[5].XIC[3].icell.PDM VGND 0.1882f
C4422 XA.XIR[5].XIC[2].icell.PDM VGND 0.1882f
C4423 XA.XIR[5].XIC[1].icell.PDM VGND 0.1882f
C4424 XA.XIR[5].XIC[0].icell.PDM VGND 0.18836f
C4425 XA.XIR[5].XIC_dummy_left.icell.PDM VGND 0.22809f
C4426 XA.XIR[4].XIC_dummy_right.icell.Iout VGND 0.85788f
C4427 XA.XIR[4].XIC_dummy_right.icell.SM VGND 0.01013f
C4428 XA.XIR[4].XIC_dummy_right.icell.Ien VGND 0.60818f
C4429 XA.XIR[4].XIC_15.icell.Ien VGND 0.37264f
C4430 XA.XIR[4].XIC[14].icell.Ien VGND 0.37333f
C4431 XA.XIR[4].XIC[13].icell.Ien VGND 0.3733f
C4432 XA.XIR[4].XIC[12].icell.Ien VGND 0.3733f
C4433 XA.XIR[4].XIC[11].icell.Ien VGND 0.3733f
C4434 XA.XIR[4].XIC[10].icell.Ien VGND 0.3733f
C4435 XA.XIR[4].XIC[9].icell.Ien VGND 0.3733f
C4436 XA.XIR[4].XIC[8].icell.Ien VGND 0.3733f
C4437 XA.XIR[4].XIC[7].icell.Ien VGND 0.3733f
C4438 XA.XIR[4].XIC[6].icell.Ien VGND 0.3733f
C4439 XA.XIR[4].XIC[5].icell.Ien VGND 0.3733f
C4440 XA.XIR[4].XIC[4].icell.Ien VGND 0.3733f
C4441 XA.XIR[4].XIC[3].icell.Ien VGND 0.3733f
C4442 XA.XIR[4].XIC[2].icell.Ien VGND 0.3733f
C4443 XA.XIR[4].XIC_dummy_left.icell.Iout VGND 0.80734f
C4444 XA.XIR[4].XIC[1].icell.Ien VGND 0.3733f
C4445 XA.XIR[4].XIC[0].icell.Ien VGND 0.37345f
C4446 XA.XIR[4].XIC_dummy_left.icell.SM VGND 0.01033f
C4447 XA.XIR[4].XIC_dummy_left.icell.Ien VGND 0.57333f
C4448 XA.XIR[4].XIC_dummy_right.icell.PDM VGND 0.23384f
C4449 XA.XIR[4].XIC_15.icell.PDM VGND 0.18862f
C4450 XA.XIR[4].XIC[14].icell.PDM VGND 0.1882f
C4451 XA.XIR[4].XIC[13].icell.PDM VGND 0.1882f
C4452 XA.XIR[4].XIC[12].icell.PDM VGND 0.1882f
C4453 XA.XIR[4].XIC[11].icell.PDM VGND 0.1882f
C4454 XA.XIR[4].XIC[10].icell.PDM VGND 0.1882f
C4455 XA.XIR[4].XIC[9].icell.PDM VGND 0.1882f
C4456 XA.XIR[4].XIC[8].icell.PDM VGND 0.1882f
C4457 XA.XIR[4].XIC[7].icell.PDM VGND 0.1882f
C4458 XA.XIR[4].XIC[6].icell.PDM VGND 0.1882f
C4459 XA.XIR[4].XIC[5].icell.PDM VGND 0.1882f
C4460 XA.XIR[4].XIC[4].icell.PDM VGND 0.1882f
C4461 XA.XIR[4].XIC[3].icell.PDM VGND 0.1882f
C4462 XA.XIR[4].XIC[2].icell.PDM VGND 0.1882f
C4463 XA.XIR[4].XIC[1].icell.PDM VGND 0.1882f
C4464 XA.XIR[4].XIC[0].icell.PDM VGND 0.18836f
C4465 XA.XIR[4].XIC_dummy_left.icell.PDM VGND 0.22809f
C4466 XThR.Tn[4] VGND 12.95212f
C4467 a_n1049_6405# VGND 0.02935f
C4468 XA.XIR[3].XIC_dummy_right.icell.Iout VGND 0.85788f
C4469 XA.XIR[3].XIC_dummy_right.icell.SM VGND 0.01013f
C4470 XA.XIR[3].XIC_dummy_right.icell.Ien VGND 0.60818f
C4471 XA.XIR[3].XIC_15.icell.Ien VGND 0.37264f
C4472 XA.XIR[3].XIC[14].icell.Ien VGND 0.37333f
C4473 XA.XIR[3].XIC[13].icell.Ien VGND 0.3733f
C4474 XA.XIR[3].XIC[12].icell.Ien VGND 0.3733f
C4475 XA.XIR[3].XIC[11].icell.Ien VGND 0.3733f
C4476 XA.XIR[3].XIC[10].icell.Ien VGND 0.3733f
C4477 XA.XIR[3].XIC[9].icell.Ien VGND 0.3733f
C4478 XA.XIR[3].XIC[8].icell.Ien VGND 0.3733f
C4479 XA.XIR[3].XIC[7].icell.Ien VGND 0.3733f
C4480 XA.XIR[3].XIC[6].icell.Ien VGND 0.3733f
C4481 XA.XIR[3].XIC[5].icell.Ien VGND 0.3733f
C4482 XA.XIR[3].XIC[4].icell.Ien VGND 0.3733f
C4483 XA.XIR[3].XIC[3].icell.Ien VGND 0.3733f
C4484 XA.XIR[3].XIC[2].icell.Ien VGND 0.3733f
C4485 XThR.XTB5.Y VGND 1.32753f
C4486 XA.XIR[3].XIC_dummy_left.icell.Iout VGND 0.80575f
C4487 XA.XIR[3].XIC[1].icell.Ien VGND 0.3733f
C4488 XA.XIR[3].XIC[0].icell.Ien VGND 0.37345f
C4489 XA.XIR[3].XIC_dummy_left.icell.SM VGND 0.01033f
C4490 XA.XIR[3].XIC_dummy_left.icell.Ien VGND 0.57422f
C4491 a_n1049_6699# VGND 0.02979f
C4492 XA.XIR[3].XIC_dummy_right.icell.PDM VGND 0.23384f
C4493 XA.XIR[3].XIC_15.icell.PDM VGND 0.18862f
C4494 XA.XIR[3].XIC[14].icell.PDM VGND 0.1882f
C4495 XA.XIR[3].XIC[13].icell.PDM VGND 0.1882f
C4496 XA.XIR[3].XIC[12].icell.PDM VGND 0.1882f
C4497 XA.XIR[3].XIC[11].icell.PDM VGND 0.1882f
C4498 XA.XIR[3].XIC[10].icell.PDM VGND 0.1882f
C4499 XA.XIR[3].XIC[9].icell.PDM VGND 0.1882f
C4500 XA.XIR[3].XIC[8].icell.PDM VGND 0.1882f
C4501 XA.XIR[3].XIC[7].icell.PDM VGND 0.1882f
C4502 XA.XIR[3].XIC[6].icell.PDM VGND 0.1882f
C4503 XA.XIR[3].XIC[5].icell.PDM VGND 0.1882f
C4504 XA.XIR[3].XIC[4].icell.PDM VGND 0.1882f
C4505 XA.XIR[3].XIC[3].icell.PDM VGND 0.1882f
C4506 XA.XIR[3].XIC[2].icell.PDM VGND 0.1882f
C4507 XA.XIR[3].XIC[1].icell.PDM VGND 0.1882f
C4508 XA.XIR[3].XIC[0].icell.PDM VGND 0.18836f
C4509 XA.XIR[3].XIC_dummy_left.icell.PDM VGND 0.22809f
C4510 XA.XIR[2].XIC_dummy_right.icell.Iout VGND 0.85788f
C4511 XA.XIR[2].XIC_dummy_right.icell.SM VGND 0.01013f
C4512 XA.XIR[2].XIC_dummy_right.icell.Ien VGND 0.60818f
C4513 XA.XIR[2].XIC_15.icell.Ien VGND 0.37264f
C4514 XA.XIR[2].XIC[14].icell.Ien VGND 0.37333f
C4515 XA.XIR[2].XIC[13].icell.Ien VGND 0.3733f
C4516 XA.XIR[2].XIC[12].icell.Ien VGND 0.3733f
C4517 XA.XIR[2].XIC[11].icell.Ien VGND 0.3733f
C4518 XA.XIR[2].XIC[10].icell.Ien VGND 0.3733f
C4519 XA.XIR[2].XIC[9].icell.Ien VGND 0.3733f
C4520 XA.XIR[2].XIC[8].icell.Ien VGND 0.3733f
C4521 XA.XIR[2].XIC[7].icell.Ien VGND 0.3733f
C4522 XA.XIR[2].XIC[6].icell.Ien VGND 0.3733f
C4523 XA.XIR[2].XIC[5].icell.Ien VGND 0.3733f
C4524 XA.XIR[2].XIC[4].icell.Ien VGND 0.3733f
C4525 XA.XIR[2].XIC[3].icell.Ien VGND 0.3733f
C4526 XA.XIR[2].XIC[2].icell.Ien VGND 0.3733f
C4527 XA.XIR[2].XIC_dummy_left.icell.Iout VGND 0.80789f
C4528 XA.XIR[2].XIC[1].icell.Ien VGND 0.3733f
C4529 XThR.Tn[3] VGND 12.94485f
C4530 XThR.XTB4.Y VGND 1.76953f
C4531 XA.XIR[2].XIC[0].icell.Ien VGND 0.37345f
C4532 XA.XIR[2].XIC_dummy_left.icell.SM VGND 0.01033f
C4533 XA.XIR[2].XIC_dummy_left.icell.Ien VGND 0.57556f
C4534 XA.XIR[2].XIC_dummy_right.icell.PDM VGND 0.23384f
C4535 XA.XIR[2].XIC_15.icell.PDM VGND 0.18862f
C4536 XA.XIR[2].XIC[14].icell.PDM VGND 0.1882f
C4537 XA.XIR[2].XIC[13].icell.PDM VGND 0.1882f
C4538 XA.XIR[2].XIC[12].icell.PDM VGND 0.1882f
C4539 XA.XIR[2].XIC[11].icell.PDM VGND 0.1882f
C4540 XA.XIR[2].XIC[10].icell.PDM VGND 0.1882f
C4541 XA.XIR[2].XIC[9].icell.PDM VGND 0.1882f
C4542 XA.XIR[2].XIC[8].icell.PDM VGND 0.1882f
C4543 XA.XIR[2].XIC[7].icell.PDM VGND 0.1882f
C4544 XA.XIR[2].XIC[6].icell.PDM VGND 0.1882f
C4545 XA.XIR[2].XIC[5].icell.PDM VGND 0.1882f
C4546 XA.XIR[2].XIC[4].icell.PDM VGND 0.1882f
C4547 XA.XIR[2].XIC[3].icell.PDM VGND 0.1882f
C4548 XA.XIR[2].XIC[2].icell.PDM VGND 0.1882f
C4549 XA.XIR[2].XIC[1].icell.PDM VGND 0.1882f
C4550 XA.XIR[2].XIC[0].icell.PDM VGND 0.18836f
C4551 XA.XIR[2].XIC_dummy_left.icell.PDM VGND 0.22809f
C4552 XA.XIR[1].XIC_dummy_right.icell.Iout VGND 0.85788f
C4553 XA.XIR[1].XIC_dummy_right.icell.SM VGND 0.01013f
C4554 XA.XIR[1].XIC_dummy_right.icell.Ien VGND 0.60818f
C4555 XA.XIR[1].XIC_15.icell.Ien VGND 0.37264f
C4556 XA.XIR[1].XIC[14].icell.Ien VGND 0.37333f
C4557 XA.XIR[1].XIC[13].icell.Ien VGND 0.3733f
C4558 XA.XIR[1].XIC[12].icell.Ien VGND 0.3733f
C4559 XA.XIR[1].XIC[11].icell.Ien VGND 0.3733f
C4560 XA.XIR[1].XIC[10].icell.Ien VGND 0.3733f
C4561 XA.XIR[1].XIC[9].icell.Ien VGND 0.3733f
C4562 XA.XIR[1].XIC[8].icell.Ien VGND 0.3733f
C4563 XA.XIR[1].XIC[7].icell.Ien VGND 0.3733f
C4564 XA.XIR[1].XIC[6].icell.Ien VGND 0.3733f
C4565 XA.XIR[1].XIC[5].icell.Ien VGND 0.3733f
C4566 XA.XIR[1].XIC[4].icell.Ien VGND 0.3733f
C4567 XA.XIR[1].XIC[3].icell.Ien VGND 0.3733f
C4568 XA.XIR[1].XIC[2].icell.Ien VGND 0.3733f
C4569 XA.XIR[1].XIC_dummy_left.icell.Iout VGND 0.80575f
C4570 XA.XIR[1].XIC[1].icell.Ien VGND 0.3733f
C4571 XThR.Tn[2] VGND 12.94933f
C4572 a_n1049_7493# VGND 0.02484f
C4573 XThR.XTB3.Y VGND 2.09162f
C4574 XThR.XTB7.A VGND 1.95537f
C4575 XA.XIR[1].XIC[0].icell.Ien VGND 0.37345f
C4576 XA.XIR[1].XIC_dummy_left.icell.SM VGND 0.01033f
C4577 XA.XIR[1].XIC_dummy_left.icell.Ien VGND 0.57376f
C4578 XA.XIR[1].XIC_dummy_right.icell.PDM VGND 0.23384f
C4579 XA.XIR[1].XIC_15.icell.PDM VGND 0.18862f
C4580 XA.XIR[1].XIC[14].icell.PDM VGND 0.1882f
C4581 XA.XIR[1].XIC[13].icell.PDM VGND 0.1882f
C4582 XA.XIR[1].XIC[12].icell.PDM VGND 0.1882f
C4583 XA.XIR[1].XIC[11].icell.PDM VGND 0.1882f
C4584 XA.XIR[1].XIC[10].icell.PDM VGND 0.1882f
C4585 XA.XIR[1].XIC[9].icell.PDM VGND 0.1882f
C4586 XA.XIR[1].XIC[8].icell.PDM VGND 0.1882f
C4587 XA.XIR[1].XIC[7].icell.PDM VGND 0.1882f
C4588 XA.XIR[1].XIC[6].icell.PDM VGND 0.1882f
C4589 XA.XIR[1].XIC[5].icell.PDM VGND 0.1882f
C4590 XA.XIR[1].XIC[4].icell.PDM VGND 0.1882f
C4591 XA.XIR[1].XIC[3].icell.PDM VGND 0.1882f
C4592 XA.XIR[1].XIC[2].icell.PDM VGND 0.1882f
C4593 XA.XIR[1].XIC[1].icell.PDM VGND 0.1882f
C4594 XA.XIR[1].XIC[0].icell.PDM VGND 0.18836f
C4595 XA.XIR[1].XIC_dummy_left.icell.PDM VGND 0.22809f
C4596 a_n1049_7787# VGND 0.03397f
C4597 XA.XIR[0].XIC_dummy_right.icell.Iout VGND 0.87403f
C4598 XA.XIR[0].XIC_dummy_right.icell.SM VGND 0.01013f
C4599 XA.XIR[0].XIC_dummy_right.icell.Ien VGND 0.61797f
C4600 XA.XIR[0].XIC_15.icell.Ien VGND 0.37874f
C4601 XA.XIR[0].XIC[14].icell.Ien VGND 0.39158f
C4602 XA.XIR[0].XIC[13].icell.Ien VGND 0.39155f
C4603 XA.XIR[0].XIC[12].icell.Ien VGND 0.38822f
C4604 XA.XIR[0].XIC[11].icell.Ien VGND 0.3889f
C4605 XA.XIR[0].XIC[10].icell.Ien VGND 0.39022f
C4606 XA.XIR[0].XIC[9].icell.Ien VGND 0.3885f
C4607 XA.XIR[0].XIC[8].icell.Ien VGND 0.38898f
C4608 XA.XIR[0].XIC[7].icell.Ien VGND 0.38927f
C4609 XA.XIR[0].XIC[6].icell.Ien VGND 0.38927f
C4610 XA.XIR[0].XIC[5].icell.Ien VGND 0.38822f
C4611 XA.XIR[0].XIC[4].icell.Ien VGND 0.38827f
C4612 XA.XIR[0].XIC[3].icell.Ien VGND 0.38951f
C4613 XA.XIR[0].XIC[2].icell.Ien VGND 0.39155f
C4614 XA.XIR[0].XIC_dummy_left.icell.Iout VGND 0.83191f
C4615 XA.XIR[0].XIC[1].icell.Ien VGND 0.39155f
C4616 XA.XIR[0].XIC[0].icell.Ien VGND 0.39086f
C4617 XA.XIR[0].XIC_dummy_left.icell.SM VGND 0.01033f
C4618 XThR.Tn[1] VGND 12.98843f
C4619 XThR.XTB2.Y VGND 1.47619f
C4620 XThR.XTB6.A VGND 0.95635f
C4621 XA.XIR[0].XIC_dummy_left.icell.Ien VGND 0.58431f
C4622 XA.XIR[0].XIC_dummy_right.icell.PDM VGND 0.251f
C4623 XA.XIR[0].XIC_15.icell.PDM VGND 0.20773f
C4624 XA.XIR[0].XIC[14].icell.PDM VGND 0.24601f
C4625 XA.XIR[0].XIC[13].icell.PDM VGND 0.24585f
C4626 XA.XIR[0].XIC[12].icell.PDM VGND 0.24146f
C4627 XA.XIR[0].XIC[11].icell.PDM VGND 0.24184f
C4628 XA.XIR[0].XIC[10].icell.PDM VGND 0.24174f
C4629 XA.XIR[0].XIC[9].icell.PDM VGND 0.24147f
C4630 XA.XIR[0].XIC[8].icell.PDM VGND 0.24147f
C4631 XA.XIR[0].XIC[7].icell.PDM VGND 0.2442f
C4632 XA.XIR[0].XIC[6].icell.PDM VGND 0.24156f
C4633 XA.XIR[0].XIC[5].icell.PDM VGND 0.24321f
C4634 XA.XIR[0].XIC[4].icell.PDM VGND 0.24159f
C4635 XA.XIR[0].XIC[3].icell.PDM VGND 0.24451f
C4636 XA.XIR[0].XIC[2].icell.PDM VGND 0.2458f
C4637 XA.XIR[0].XIC[1].icell.PDM VGND 0.2458f
C4638 XA.XIR[0].XIC[0].icell.PDM VGND 0.2446f
C4639 XA.XIR[0].XIC_dummy_left.icell.PDM VGND 0.24577f
C4640 XThR.Tn[0] VGND 13.29619f
C4641 a_n1049_8581# VGND 0.04333f
C4642 XThR.XTBN.Y VGND 7.54415f
C4643 XThR.XTB1.Y VGND 1.45322f
C4644 XThR.XTB7.B VGND 2.61063f
C4645 XThR.XTB5.A VGND 1.75777f
C4646 XA.Cn[14] VGND 5.52615f
C4647 XA.Cn[13] VGND 5.16689f
C4648 XA.Cn[12] VGND 5.1562f
C4649 XA.Cn[11] VGND 5.52379f
C4650 XA.Cn[10] VGND 5.0515f
C4651 XA.Cn[9] VGND 5.34336f
C4652 XA.Cn[8] VGND 4.89287f
C4653 a_10915_9569# VGND 0.55912f
C4654 a_10051_9569# VGND 0.55747f
C4655 a_9827_9569# VGND 0.54584f
C4656 a_8963_9569# VGND 0.55439f
C4657 a_8739_9569# VGND 0.553f
C4658 a_7875_9569# VGND 0.55432f
C4659 a_7651_9569# VGND 0.55717f
C4660 XA.Cn[7] VGND 5.47379f
C4661 XA.Cn[6] VGND 5.48958f
C4662 XA.Cn[5] VGND 5.60438f
C4663 XA.Cn[4] VGND 5.55465f
C4664 XA.Cn[3] VGND 5.88113f
C4665 XA.Cn[2] VGND 5.58437f
C4666 XA.Cn[1] VGND 5.71923f
C4667 XA.Cn[0] VGND 6.86777f
C4668 a_6243_9615# VGND 0.03028f
C4669 a_5949_9615# VGND 0.03456f
C4670 a_5155_9615# VGND 0.03624f
C4671 a_4861_9615# VGND 0.03647f
C4672 a_4067_9615# VGND 0.03118f
C4673 a_3773_9615# VGND 0.03896f
C4674 a_2979_9615# VGND 0.04122f
C4675 thermo15c_0.XTBN.Y VGND 8.71711f
C4676 thermo15c_0.XTB7.Y VGND 1.35988f
C4677 thermo15c_0.XTB6.Y VGND 1.3794f
C4678 thermo15c_0.XTB7.B VGND 2.83799f
C4679 thermo15c_0.XTB5.Y VGND 1.32558f
C4680 thermo15c_0.XTBN.A VGND 1.2246f
C4681 thermo15c_0.XTB4.Y VGND 1.69704f
C4682 thermo15c_0.XTB3.Y VGND 1.96717f
C4683 thermo15c_0.XTB7.A VGND 1.94951f
C4684 thermo15c_0.XTB6.A VGND 0.95452f
C4685 thermo15c_0.XTB2.Y VGND 1.4752f
C4686 thermo15c_0.XTB1.Y VGND 1.77643f
C4687 thermo15c_0.XTB5.A VGND 1.75974f
C4688 bias[0].t0 VGND 0.94587f
C4689 XThR.XTB3.Y.t1 VGND 0.06176f
C4690 XThR.XTB3.Y.n0 VGND 0.01521f
C4691 XThR.XTB3.Y.t8 VGND 0.04903f
C4692 XThR.XTB3.Y.t15 VGND 0.02889f
C4693 XThR.XTB3.Y.t13 VGND 0.04903f
C4694 XThR.XTB3.Y.t6 VGND 0.02889f
C4695 XThR.XTB3.Y.t9 VGND 0.04903f
C4696 XThR.XTB3.Y.t17 VGND 0.02889f
C4697 XThR.XTB3.Y.n1 VGND 0.08226f
C4698 XThR.XTB3.Y.n2 VGND 0.08688f
C4699 XThR.XTB3.Y.n3 VGND 0.03573f
C4700 XThR.XTB3.Y.n4 VGND 0.0707f
C4701 XThR.XTB3.Y.t12 VGND 0.04903f
C4702 XThR.XTB3.Y.t4 VGND 0.02889f
C4703 XThR.XTB3.Y.n5 VGND 0.06608f
C4704 XThR.XTB3.Y.n6 VGND 0.03236f
C4705 XThR.XTB3.Y.n7 VGND 0.02685f
C4706 XThR.XTB3.Y.t18 VGND 0.04903f
C4707 XThR.XTB3.Y.t5 VGND 0.02889f
C4708 XThR.XTB3.Y.n8 VGND 0.03005f
C4709 XThR.XTB3.Y.t7 VGND 0.04903f
C4710 XThR.XTB3.Y.t10 VGND 0.02889f
C4711 XThR.XTB3.Y.n9 VGND 0.05992f
C4712 XThR.XTB3.Y.t11 VGND 0.04903f
C4713 XThR.XTB3.Y.t16 VGND 0.02889f
C4714 XThR.XTB3.Y.n10 VGND 0.06454f
C4715 XThR.XTB3.Y.n11 VGND 0.03645f
C4716 XThR.XTB3.Y.n12 VGND 0.06034f
C4717 XThR.XTB3.Y.n13 VGND 0.03128f
C4718 XThR.XTB3.Y.n14 VGND 0.02851f
C4719 XThR.XTB3.Y.n15 VGND 0.06454f
C4720 XThR.XTB3.Y.t14 VGND 0.04903f
C4721 XThR.XTB3.Y.t3 VGND 0.02889f
C4722 XThR.XTB3.Y.n16 VGND 0.05838f
C4723 XThR.XTB3.Y.n17 VGND 0.03236f
C4724 XThR.XTB3.Y.n18 VGND 0.04707f
C4725 XThR.XTB3.Y.n19 VGND 1.31347f
C4726 XThR.XTB3.Y.t0 VGND 0.03152f
C4727 XThR.XTB3.Y.t2 VGND 0.03152f
C4728 XThR.XTB3.Y.n20 VGND 0.06766f
C4729 XThR.XTB3.Y.n21 VGND 0.157f
C4730 XThR.XTB3.Y.n22 VGND 0.03296f
C4731 XThR.XTB4.Y.t8 VGND 0.02956f
C4732 XThR.XTB4.Y.t15 VGND 0.05016f
C4733 XThR.XTB4.Y.t16 VGND 0.02956f
C4734 XThR.XTB4.Y.t5 VGND 0.05016f
C4735 XThR.XTB4.Y.t10 VGND 0.02956f
C4736 XThR.XTB4.Y.t17 VGND 0.05016f
C4737 XThR.XTB4.Y.n0 VGND 0.08416f
C4738 XThR.XTB4.Y.n1 VGND 0.08889f
C4739 XThR.XTB4.Y.n2 VGND 0.03656f
C4740 XThR.XTB4.Y.n3 VGND 0.07234f
C4741 XThR.XTB4.Y.t13 VGND 0.02956f
C4742 XThR.XTB4.Y.t4 VGND 0.05016f
C4743 XThR.XTB4.Y.n4 VGND 0.06761f
C4744 XThR.XTB4.Y.n5 VGND 0.0331f
C4745 XThR.XTB4.Y.n6 VGND 0.01685f
C4746 XThR.XTB4.Y.n7 VGND 0.05355f
C4747 XThR.XTB4.Y.n8 VGND 0.64921f
C4748 XThR.XTB4.Y.t14 VGND 0.02956f
C4749 XThR.XTB4.Y.t7 VGND 0.05016f
C4750 XThR.XTB4.Y.n9 VGND 0.03074f
C4751 XThR.XTB4.Y.t3 VGND 0.02956f
C4752 XThR.XTB4.Y.t12 VGND 0.05016f
C4753 XThR.XTB4.Y.n10 VGND 0.0613f
C4754 XThR.XTB4.Y.t9 VGND 0.02956f
C4755 XThR.XTB4.Y.t2 VGND 0.05016f
C4756 XThR.XTB4.Y.n11 VGND 0.06603f
C4757 XThR.XTB4.Y.n12 VGND 0.03729f
C4758 XThR.XTB4.Y.n13 VGND 0.06174f
C4759 XThR.XTB4.Y.n14 VGND 0.03201f
C4760 XThR.XTB4.Y.n15 VGND 0.02916f
C4761 XThR.XTB4.Y.n16 VGND 0.06603f
C4762 XThR.XTB4.Y.t11 VGND 0.02956f
C4763 XThR.XTB4.Y.t6 VGND 0.05016f
C4764 XThR.XTB4.Y.n17 VGND 0.05972f
C4765 XThR.XTB4.Y.n18 VGND 0.0331f
C4766 XThR.XTB4.Y.n19 VGND 0.05647f
C4767 XThR.XTB4.Y.n20 VGND 1.3092f
C4768 XThR.XTB4.Y.t1 VGND 0.06491f
C4769 XThR.XTB4.Y.n21 VGND 0.12281f
C4770 XThR.XTB4.Y.n22 VGND 0.02892f
C4771 XThR.XTB4.Y.t0 VGND 0.11919f
C4772 XThR.Tn[13].t9 VGND 0.01909f
C4773 XThR.Tn[13].t11 VGND 0.01909f
C4774 XThR.Tn[13].n0 VGND 0.05796f
C4775 XThR.Tn[13].t10 VGND 0.01909f
C4776 XThR.Tn[13].t8 VGND 0.01909f
C4777 XThR.Tn[13].n1 VGND 0.04243f
C4778 XThR.Tn[13].n2 VGND 0.19293f
C4779 XThR.Tn[13].t7 VGND 0.01241f
C4780 XThR.Tn[13].t5 VGND 0.01241f
C4781 XThR.Tn[13].n3 VGND 0.03094f
C4782 XThR.Tn[13].t6 VGND 0.01241f
C4783 XThR.Tn[13].t4 VGND 0.01241f
C4784 XThR.Tn[13].n4 VGND 0.02481f
C4785 XThR.Tn[13].n5 VGND 0.06242f
C4786 XThR.Tn[13].t72 VGND 0.01492f
C4787 XThR.Tn[13].t64 VGND 0.01633f
C4788 XThR.Tn[13].n6 VGND 0.03989f
C4789 XThR.Tn[13].n7 VGND 0.07663f
C4790 XThR.Tn[13].t28 VGND 0.01492f
C4791 XThR.Tn[13].t21 VGND 0.01633f
C4792 XThR.Tn[13].n8 VGND 0.03989f
C4793 XThR.Tn[13].t44 VGND 0.01487f
C4794 XThR.Tn[13].t12 VGND 0.01628f
C4795 XThR.Tn[13].n9 VGND 0.0415f
C4796 XThR.Tn[13].n10 VGND 0.02916f
C4797 XThR.Tn[13].n12 VGND 0.09357f
C4798 XThR.Tn[13].t65 VGND 0.01492f
C4799 XThR.Tn[13].t57 VGND 0.01633f
C4800 XThR.Tn[13].n13 VGND 0.03989f
C4801 XThR.Tn[13].t19 VGND 0.01487f
C4802 XThR.Tn[13].t52 VGND 0.01628f
C4803 XThR.Tn[13].n14 VGND 0.0415f
C4804 XThR.Tn[13].n15 VGND 0.02916f
C4805 XThR.Tn[13].n17 VGND 0.09357f
C4806 XThR.Tn[13].t22 VGND 0.01492f
C4807 XThR.Tn[13].t14 VGND 0.01633f
C4808 XThR.Tn[13].n18 VGND 0.03989f
C4809 XThR.Tn[13].t34 VGND 0.01487f
C4810 XThR.Tn[13].t70 VGND 0.01628f
C4811 XThR.Tn[13].n19 VGND 0.0415f
C4812 XThR.Tn[13].n20 VGND 0.02916f
C4813 XThR.Tn[13].n22 VGND 0.09357f
C4814 XThR.Tn[13].t49 VGND 0.01492f
C4815 XThR.Tn[13].t39 VGND 0.01633f
C4816 XThR.Tn[13].n23 VGND 0.03989f
C4817 XThR.Tn[13].t66 VGND 0.01487f
C4818 XThR.Tn[13].t35 VGND 0.01628f
C4819 XThR.Tn[13].n24 VGND 0.0415f
C4820 XThR.Tn[13].n25 VGND 0.02916f
C4821 XThR.Tn[13].n27 VGND 0.09357f
C4822 XThR.Tn[13].t24 VGND 0.01492f
C4823 XThR.Tn[13].t16 VGND 0.01633f
C4824 XThR.Tn[13].n28 VGND 0.03989f
C4825 XThR.Tn[13].t37 VGND 0.01487f
C4826 XThR.Tn[13].t71 VGND 0.01628f
C4827 XThR.Tn[13].n29 VGND 0.0415f
C4828 XThR.Tn[13].n30 VGND 0.02916f
C4829 XThR.Tn[13].n32 VGND 0.09357f
C4830 XThR.Tn[13].t60 VGND 0.01492f
C4831 XThR.Tn[13].t30 VGND 0.01633f
C4832 XThR.Tn[13].n33 VGND 0.03989f
C4833 XThR.Tn[13].t13 VGND 0.01487f
C4834 XThR.Tn[13].t26 VGND 0.01628f
C4835 XThR.Tn[13].n34 VGND 0.0415f
C4836 XThR.Tn[13].n35 VGND 0.02916f
C4837 XThR.Tn[13].n37 VGND 0.09357f
C4838 XThR.Tn[13].t29 VGND 0.01492f
C4839 XThR.Tn[13].t25 VGND 0.01633f
C4840 XThR.Tn[13].n38 VGND 0.03989f
C4841 XThR.Tn[13].t43 VGND 0.01487f
C4842 XThR.Tn[13].t18 VGND 0.01628f
C4843 XThR.Tn[13].n39 VGND 0.0415f
C4844 XThR.Tn[13].n40 VGND 0.02916f
C4845 XThR.Tn[13].n42 VGND 0.09357f
C4846 XThR.Tn[13].t32 VGND 0.01492f
C4847 XThR.Tn[13].t38 VGND 0.01633f
C4848 XThR.Tn[13].n43 VGND 0.03989f
C4849 XThR.Tn[13].t48 VGND 0.01487f
C4850 XThR.Tn[13].t33 VGND 0.01628f
C4851 XThR.Tn[13].n44 VGND 0.0415f
C4852 XThR.Tn[13].n45 VGND 0.02916f
C4853 XThR.Tn[13].n47 VGND 0.09357f
C4854 XThR.Tn[13].t51 VGND 0.01492f
C4855 XThR.Tn[13].t59 VGND 0.01633f
C4856 XThR.Tn[13].n48 VGND 0.03989f
C4857 XThR.Tn[13].t68 VGND 0.01487f
C4858 XThR.Tn[13].t53 VGND 0.01628f
C4859 XThR.Tn[13].n49 VGND 0.0415f
C4860 XThR.Tn[13].n50 VGND 0.02916f
C4861 XThR.Tn[13].n52 VGND 0.09357f
C4862 XThR.Tn[13].t41 VGND 0.01492f
C4863 XThR.Tn[13].t17 VGND 0.01633f
C4864 XThR.Tn[13].n53 VGND 0.03989f
C4865 XThR.Tn[13].t58 VGND 0.01487f
C4866 XThR.Tn[13].t73 VGND 0.01628f
C4867 XThR.Tn[13].n54 VGND 0.0415f
C4868 XThR.Tn[13].n55 VGND 0.02916f
C4869 XThR.Tn[13].n57 VGND 0.09357f
C4870 XThR.Tn[13].t63 VGND 0.01492f
C4871 XThR.Tn[13].t55 VGND 0.01633f
C4872 XThR.Tn[13].n58 VGND 0.03989f
C4873 XThR.Tn[13].t15 VGND 0.01487f
C4874 XThR.Tn[13].t45 VGND 0.01628f
C4875 XThR.Tn[13].n59 VGND 0.0415f
C4876 XThR.Tn[13].n60 VGND 0.02916f
C4877 XThR.Tn[13].n62 VGND 0.09357f
C4878 XThR.Tn[13].t31 VGND 0.01492f
C4879 XThR.Tn[13].t27 VGND 0.01633f
C4880 XThR.Tn[13].n63 VGND 0.03989f
C4881 XThR.Tn[13].t46 VGND 0.01487f
C4882 XThR.Tn[13].t20 VGND 0.01628f
C4883 XThR.Tn[13].n64 VGND 0.0415f
C4884 XThR.Tn[13].n65 VGND 0.02916f
C4885 XThR.Tn[13].n67 VGND 0.09357f
C4886 XThR.Tn[13].t50 VGND 0.01492f
C4887 XThR.Tn[13].t40 VGND 0.01633f
C4888 XThR.Tn[13].n68 VGND 0.03989f
C4889 XThR.Tn[13].t67 VGND 0.01487f
C4890 XThR.Tn[13].t36 VGND 0.01628f
C4891 XThR.Tn[13].n69 VGND 0.0415f
C4892 XThR.Tn[13].n70 VGND 0.02916f
C4893 XThR.Tn[13].n72 VGND 0.09357f
C4894 XThR.Tn[13].t69 VGND 0.01492f
C4895 XThR.Tn[13].t62 VGND 0.01633f
C4896 XThR.Tn[13].n73 VGND 0.03989f
C4897 XThR.Tn[13].t23 VGND 0.01487f
C4898 XThR.Tn[13].t54 VGND 0.01628f
C4899 XThR.Tn[13].n74 VGND 0.0415f
C4900 XThR.Tn[13].n75 VGND 0.02916f
C4901 XThR.Tn[13].n77 VGND 0.09357f
C4902 XThR.Tn[13].t42 VGND 0.01492f
C4903 XThR.Tn[13].t56 VGND 0.01633f
C4904 XThR.Tn[13].n78 VGND 0.03989f
C4905 XThR.Tn[13].t61 VGND 0.01487f
C4906 XThR.Tn[13].t47 VGND 0.01628f
C4907 XThR.Tn[13].n79 VGND 0.0415f
C4908 XThR.Tn[13].n80 VGND 0.02916f
C4909 XThR.Tn[13].n82 VGND 0.09357f
C4910 XThR.Tn[13].n83 VGND 0.08503f
C4911 XThR.Tn[13].n84 VGND 0.33338f
C4912 XThR.Tn[13].t2 VGND 0.01909f
C4913 XThR.Tn[13].t0 VGND 0.01909f
C4914 XThR.Tn[13].n85 VGND 0.04124f
C4915 XThR.Tn[13].t3 VGND 0.01909f
C4916 XThR.Tn[13].t1 VGND 0.01909f
C4917 XThR.Tn[13].n86 VGND 0.06277f
C4918 XThR.Tn[13].n87 VGND 0.17429f
C4919 XThR.Tn[13].n88 VGND 0.02334f
C4920 thermo15c_0.XTB3.Y.t1 VGND 0.06296f
C4921 thermo15c_0.XTB3.Y.n0 VGND 0.04069f
C4922 thermo15c_0.XTB3.Y.n1 VGND 0.05192f
C4923 thermo15c_0.XTB3.Y.t2 VGND 0.03159f
C4924 thermo15c_0.XTB3.Y.t0 VGND 0.03159f
C4925 thermo15c_0.XTB3.Y.n2 VGND 0.06782f
C4926 thermo15c_0.XTB3.Y.t10 VGND 0.04914f
C4927 thermo15c_0.XTB3.Y.t17 VGND 0.02896f
C4928 thermo15c_0.XTB3.Y.n3 VGND 0.05852f
C4929 thermo15c_0.XTB3.Y.t14 VGND 0.04914f
C4930 thermo15c_0.XTB3.Y.t5 VGND 0.02896f
C4931 thermo15c_0.XTB3.Y.n4 VGND 0.03012f
C4932 thermo15c_0.XTB3.Y.t15 VGND 0.04914f
C4933 thermo15c_0.XTB3.Y.t6 VGND 0.02896f
C4934 thermo15c_0.XTB3.Y.n5 VGND 0.06469f
C4935 thermo15c_0.XTB3.Y.t3 VGND 0.04914f
C4936 thermo15c_0.XTB3.Y.t9 VGND 0.02896f
C4937 thermo15c_0.XTB3.Y.n6 VGND 0.06006f
C4938 thermo15c_0.XTB3.Y.n7 VGND 0.03654f
C4939 thermo15c_0.XTB3.Y.n8 VGND 0.06049f
C4940 thermo15c_0.XTB3.Y.n9 VGND 0.0234f
C4941 thermo15c_0.XTB3.Y.n10 VGND 0.02857f
C4942 thermo15c_0.XTB3.Y.n11 VGND 0.06469f
C4943 thermo15c_0.XTB3.Y.n12 VGND 0.03243f
C4944 thermo15c_0.XTB3.Y.n13 VGND 0.05514f
C4945 thermo15c_0.XTB3.Y.t16 VGND 0.04914f
C4946 thermo15c_0.XTB3.Y.t7 VGND 0.02896f
C4947 thermo15c_0.XTB3.Y.n14 VGND 0.06624f
C4948 thermo15c_0.XTB3.Y.t4 VGND 0.04914f
C4949 thermo15c_0.XTB3.Y.t13 VGND 0.02896f
C4950 thermo15c_0.XTB3.Y.t12 VGND 0.04914f
C4951 thermo15c_0.XTB3.Y.t18 VGND 0.02896f
C4952 thermo15c_0.XTB3.Y.t11 VGND 0.04914f
C4953 thermo15c_0.XTB3.Y.t8 VGND 0.02896f
C4954 thermo15c_0.XTB3.Y.n15 VGND 0.08245f
C4955 thermo15c_0.XTB3.Y.n16 VGND 0.08709f
C4956 thermo15c_0.XTB3.Y.n17 VGND 0.03356f
C4957 thermo15c_0.XTB3.Y.n18 VGND 0.07087f
C4958 thermo15c_0.XTB3.Y.n19 VGND 0.03243f
C4959 thermo15c_0.XTB3.Y.n20 VGND 0.02691f
C4960 thermo15c_0.XTB3.Y.n21 VGND 1.39635f
C4961 thermo15c_0.XTB3.Y.n22 VGND 0.14933f
C4962 XThR.Tn[8].t10 VGND 0.01919f
C4963 XThR.Tn[8].t8 VGND 0.01919f
C4964 XThR.Tn[8].n0 VGND 0.05828f
C4965 XThR.Tn[8].t11 VGND 0.01919f
C4966 XThR.Tn[8].t9 VGND 0.01919f
C4967 XThR.Tn[8].n1 VGND 0.04267f
C4968 XThR.Tn[8].n2 VGND 0.19401f
C4969 XThR.Tn[8].t5 VGND 0.01248f
C4970 XThR.Tn[8].t7 VGND 0.01248f
C4971 XThR.Tn[8].n3 VGND 0.03112f
C4972 XThR.Tn[8].t4 VGND 0.01248f
C4973 XThR.Tn[8].t6 VGND 0.01248f
C4974 XThR.Tn[8].n4 VGND 0.02495f
C4975 XThR.Tn[8].n5 VGND 0.05754f
C4976 XThR.Tn[8].t39 VGND 0.015f
C4977 XThR.Tn[8].t33 VGND 0.01643f
C4978 XThR.Tn[8].n6 VGND 0.04011f
C4979 XThR.Tn[8].n7 VGND 0.07706f
C4980 XThR.Tn[8].t59 VGND 0.015f
C4981 XThR.Tn[8].t49 VGND 0.01643f
C4982 XThR.Tn[8].n8 VGND 0.04011f
C4983 XThR.Tn[8].t13 VGND 0.01495f
C4984 XThR.Tn[8].t45 VGND 0.01637f
C4985 XThR.Tn[8].n9 VGND 0.04174f
C4986 XThR.Tn[8].n10 VGND 0.02932f
C4987 XThR.Tn[8].n12 VGND 0.09409f
C4988 XThR.Tn[8].t34 VGND 0.015f
C4989 XThR.Tn[8].t26 VGND 0.01643f
C4990 XThR.Tn[8].n13 VGND 0.04011f
C4991 XThR.Tn[8].t53 VGND 0.01495f
C4992 XThR.Tn[8].t22 VGND 0.01637f
C4993 XThR.Tn[8].n14 VGND 0.04174f
C4994 XThR.Tn[8].n15 VGND 0.02932f
C4995 XThR.Tn[8].n17 VGND 0.09409f
C4996 XThR.Tn[8].t50 VGND 0.015f
C4997 XThR.Tn[8].t43 VGND 0.01643f
C4998 XThR.Tn[8].n18 VGND 0.04011f
C4999 XThR.Tn[8].t65 VGND 0.01495f
C5000 XThR.Tn[8].t40 VGND 0.01637f
C5001 XThR.Tn[8].n19 VGND 0.04174f
C5002 XThR.Tn[8].n20 VGND 0.02932f
C5003 XThR.Tn[8].n22 VGND 0.09409f
C5004 XThR.Tn[8].t12 VGND 0.015f
C5005 XThR.Tn[8].t70 VGND 0.01643f
C5006 XThR.Tn[8].n23 VGND 0.04011f
C5007 XThR.Tn[8].t36 VGND 0.01495f
C5008 XThR.Tn[8].t66 VGND 0.01637f
C5009 XThR.Tn[8].n24 VGND 0.04174f
C5010 XThR.Tn[8].n25 VGND 0.02932f
C5011 XThR.Tn[8].n27 VGND 0.09409f
C5012 XThR.Tn[8].t52 VGND 0.015f
C5013 XThR.Tn[8].t44 VGND 0.01643f
C5014 XThR.Tn[8].n28 VGND 0.04011f
C5015 XThR.Tn[8].t68 VGND 0.01495f
C5016 XThR.Tn[8].t41 VGND 0.01637f
C5017 XThR.Tn[8].n29 VGND 0.04174f
C5018 XThR.Tn[8].n30 VGND 0.02932f
C5019 XThR.Tn[8].n32 VGND 0.09409f
C5020 XThR.Tn[8].t28 VGND 0.015f
C5021 XThR.Tn[8].t61 VGND 0.01643f
C5022 XThR.Tn[8].n33 VGND 0.04011f
C5023 XThR.Tn[8].t47 VGND 0.01495f
C5024 XThR.Tn[8].t58 VGND 0.01637f
C5025 XThR.Tn[8].n34 VGND 0.04174f
C5026 XThR.Tn[8].n35 VGND 0.02932f
C5027 XThR.Tn[8].n37 VGND 0.09409f
C5028 XThR.Tn[8].t60 VGND 0.015f
C5029 XThR.Tn[8].t56 VGND 0.01643f
C5030 XThR.Tn[8].n38 VGND 0.04011f
C5031 XThR.Tn[8].t14 VGND 0.01495f
C5032 XThR.Tn[8].t51 VGND 0.01637f
C5033 XThR.Tn[8].n39 VGND 0.04174f
C5034 XThR.Tn[8].n40 VGND 0.02932f
C5035 XThR.Tn[8].n42 VGND 0.09409f
C5036 XThR.Tn[8].t63 VGND 0.015f
C5037 XThR.Tn[8].t69 VGND 0.01643f
C5038 XThR.Tn[8].n43 VGND 0.04011f
C5039 XThR.Tn[8].t20 VGND 0.01495f
C5040 XThR.Tn[8].t64 VGND 0.01637f
C5041 XThR.Tn[8].n44 VGND 0.04174f
C5042 XThR.Tn[8].n45 VGND 0.02932f
C5043 XThR.Tn[8].n47 VGND 0.09409f
C5044 XThR.Tn[8].t17 VGND 0.015f
C5045 XThR.Tn[8].t27 VGND 0.01643f
C5046 XThR.Tn[8].n48 VGND 0.04011f
C5047 XThR.Tn[8].t38 VGND 0.01495f
C5048 XThR.Tn[8].t24 VGND 0.01637f
C5049 XThR.Tn[8].n49 VGND 0.04174f
C5050 XThR.Tn[8].n50 VGND 0.02932f
C5051 XThR.Tn[8].n52 VGND 0.09409f
C5052 XThR.Tn[8].t72 VGND 0.015f
C5053 XThR.Tn[8].t46 VGND 0.01643f
C5054 XThR.Tn[8].n53 VGND 0.04011f
C5055 XThR.Tn[8].t31 VGND 0.01495f
C5056 XThR.Tn[8].t42 VGND 0.01637f
C5057 XThR.Tn[8].n54 VGND 0.04174f
C5058 XThR.Tn[8].n55 VGND 0.02932f
C5059 XThR.Tn[8].n57 VGND 0.09409f
C5060 XThR.Tn[8].t30 VGND 0.015f
C5061 XThR.Tn[8].t21 VGND 0.01643f
C5062 XThR.Tn[8].n58 VGND 0.04011f
C5063 XThR.Tn[8].t48 VGND 0.01495f
C5064 XThR.Tn[8].t16 VGND 0.01637f
C5065 XThR.Tn[8].n59 VGND 0.04174f
C5066 XThR.Tn[8].n60 VGND 0.02932f
C5067 XThR.Tn[8].n62 VGND 0.09409f
C5068 XThR.Tn[8].t62 VGND 0.015f
C5069 XThR.Tn[8].t57 VGND 0.01643f
C5070 XThR.Tn[8].n63 VGND 0.04011f
C5071 XThR.Tn[8].t18 VGND 0.01495f
C5072 XThR.Tn[8].t54 VGND 0.01637f
C5073 XThR.Tn[8].n64 VGND 0.04174f
C5074 XThR.Tn[8].n65 VGND 0.02932f
C5075 XThR.Tn[8].n67 VGND 0.09409f
C5076 XThR.Tn[8].t15 VGND 0.015f
C5077 XThR.Tn[8].t71 VGND 0.01643f
C5078 XThR.Tn[8].n68 VGND 0.04011f
C5079 XThR.Tn[8].t37 VGND 0.01495f
C5080 XThR.Tn[8].t67 VGND 0.01637f
C5081 XThR.Tn[8].n69 VGND 0.04174f
C5082 XThR.Tn[8].n70 VGND 0.02932f
C5083 XThR.Tn[8].n72 VGND 0.09409f
C5084 XThR.Tn[8].t35 VGND 0.015f
C5085 XThR.Tn[8].t29 VGND 0.01643f
C5086 XThR.Tn[8].n73 VGND 0.04011f
C5087 XThR.Tn[8].t55 VGND 0.01495f
C5088 XThR.Tn[8].t25 VGND 0.01637f
C5089 XThR.Tn[8].n74 VGND 0.04174f
C5090 XThR.Tn[8].n75 VGND 0.02932f
C5091 XThR.Tn[8].n77 VGND 0.09409f
C5092 XThR.Tn[8].t73 VGND 0.015f
C5093 XThR.Tn[8].t23 VGND 0.01643f
C5094 XThR.Tn[8].n78 VGND 0.04011f
C5095 XThR.Tn[8].t32 VGND 0.01495f
C5096 XThR.Tn[8].t19 VGND 0.01637f
C5097 XThR.Tn[8].n79 VGND 0.04174f
C5098 XThR.Tn[8].n80 VGND 0.02932f
C5099 XThR.Tn[8].n82 VGND 0.09409f
C5100 XThR.Tn[8].n83 VGND 0.08551f
C5101 XThR.Tn[8].n84 VGND 0.26201f
C5102 XThR.Tn[8].t2 VGND 0.01919f
C5103 XThR.Tn[8].t0 VGND 0.01919f
C5104 XThR.Tn[8].n85 VGND 0.04147f
C5105 XThR.Tn[8].t3 VGND 0.01919f
C5106 XThR.Tn[8].t1 VGND 0.01919f
C5107 XThR.Tn[8].n86 VGND 0.06312f
C5108 XThR.Tn[8].n87 VGND 0.17526f
C5109 XThR.Tn[0].t6 VGND 0.01769f
C5110 XThR.Tn[0].t7 VGND 0.01769f
C5111 XThR.Tn[0].n0 VGND 0.03571f
C5112 XThR.Tn[0].t5 VGND 0.01769f
C5113 XThR.Tn[0].t4 VGND 0.01769f
C5114 XThR.Tn[0].n1 VGND 0.04178f
C5115 XThR.Tn[0].n2 VGND 0.12532f
C5116 XThR.Tn[0].t9 VGND 0.0115f
C5117 XThR.Tn[0].t10 VGND 0.0115f
C5118 XThR.Tn[0].n3 VGND 0.02618f
C5119 XThR.Tn[0].t8 VGND 0.0115f
C5120 XThR.Tn[0].t11 VGND 0.0115f
C5121 XThR.Tn[0].n4 VGND 0.02618f
C5122 XThR.Tn[0].t1 VGND 0.0115f
C5123 XThR.Tn[0].t2 VGND 0.0115f
C5124 XThR.Tn[0].n5 VGND 0.04363f
C5125 XThR.Tn[0].t0 VGND 0.0115f
C5126 XThR.Tn[0].t3 VGND 0.0115f
C5127 XThR.Tn[0].n6 VGND 0.02618f
C5128 XThR.Tn[0].n7 VGND 0.12469f
C5129 XThR.Tn[0].n8 VGND 0.07708f
C5130 XThR.Tn[0].n9 VGND 0.08699f
C5131 XThR.Tn[0].t48 VGND 0.01383f
C5132 XThR.Tn[0].t40 VGND 0.01514f
C5133 XThR.Tn[0].n10 VGND 0.03697f
C5134 XThR.Tn[0].n11 VGND 0.07101f
C5135 XThR.Tn[0].t67 VGND 0.01383f
C5136 XThR.Tn[0].t58 VGND 0.01514f
C5137 XThR.Tn[0].n12 VGND 0.03697f
C5138 XThR.Tn[0].t24 VGND 0.01378f
C5139 XThR.Tn[0].t50 VGND 0.01509f
C5140 XThR.Tn[0].n13 VGND 0.03846f
C5141 XThR.Tn[0].n14 VGND 0.02702f
C5142 XThR.Tn[0].n16 VGND 0.08671f
C5143 XThR.Tn[0].t41 VGND 0.01383f
C5144 XThR.Tn[0].t33 VGND 0.01514f
C5145 XThR.Tn[0].n17 VGND 0.03697f
C5146 XThR.Tn[0].t61 VGND 0.01378f
C5147 XThR.Tn[0].t26 VGND 0.01509f
C5148 XThR.Tn[0].n18 VGND 0.03846f
C5149 XThR.Tn[0].n19 VGND 0.02702f
C5150 XThR.Tn[0].n21 VGND 0.08671f
C5151 XThR.Tn[0].t59 VGND 0.01383f
C5152 XThR.Tn[0].t51 VGND 0.01514f
C5153 XThR.Tn[0].n22 VGND 0.03697f
C5154 XThR.Tn[0].t12 VGND 0.01378f
C5155 XThR.Tn[0].t44 VGND 0.01509f
C5156 XThR.Tn[0].n23 VGND 0.03846f
C5157 XThR.Tn[0].n24 VGND 0.02702f
C5158 XThR.Tn[0].n26 VGND 0.08671f
C5159 XThR.Tn[0].t21 VGND 0.01383f
C5160 XThR.Tn[0].t15 VGND 0.01514f
C5161 XThR.Tn[0].n27 VGND 0.03697f
C5162 XThR.Tn[0].t43 VGND 0.01378f
C5163 XThR.Tn[0].t72 VGND 0.01509f
C5164 XThR.Tn[0].n28 VGND 0.03846f
C5165 XThR.Tn[0].n29 VGND 0.02702f
C5166 XThR.Tn[0].n31 VGND 0.08671f
C5167 XThR.Tn[0].t60 VGND 0.01383f
C5168 XThR.Tn[0].t52 VGND 0.01514f
C5169 XThR.Tn[0].n32 VGND 0.03697f
C5170 XThR.Tn[0].t13 VGND 0.01378f
C5171 XThR.Tn[0].t46 VGND 0.01509f
C5172 XThR.Tn[0].n33 VGND 0.03846f
C5173 XThR.Tn[0].n34 VGND 0.02702f
C5174 XThR.Tn[0].n36 VGND 0.08671f
C5175 XThR.Tn[0].t35 VGND 0.01383f
C5176 XThR.Tn[0].t68 VGND 0.01514f
C5177 XThR.Tn[0].n37 VGND 0.03697f
C5178 XThR.Tn[0].t54 VGND 0.01378f
C5179 XThR.Tn[0].t64 VGND 0.01509f
C5180 XThR.Tn[0].n38 VGND 0.03846f
C5181 XThR.Tn[0].n39 VGND 0.02702f
C5182 XThR.Tn[0].n41 VGND 0.08671f
C5183 XThR.Tn[0].t66 VGND 0.01383f
C5184 XThR.Tn[0].t63 VGND 0.01514f
C5185 XThR.Tn[0].n42 VGND 0.03697f
C5186 XThR.Tn[0].t23 VGND 0.01378f
C5187 XThR.Tn[0].t55 VGND 0.01509f
C5188 XThR.Tn[0].n43 VGND 0.03846f
C5189 XThR.Tn[0].n44 VGND 0.02702f
C5190 XThR.Tn[0].n46 VGND 0.08671f
C5191 XThR.Tn[0].t70 VGND 0.01383f
C5192 XThR.Tn[0].t14 VGND 0.01514f
C5193 XThR.Tn[0].n47 VGND 0.03697f
C5194 XThR.Tn[0].t28 VGND 0.01378f
C5195 XThR.Tn[0].t71 VGND 0.01509f
C5196 XThR.Tn[0].n48 VGND 0.03846f
C5197 XThR.Tn[0].n49 VGND 0.02702f
C5198 XThR.Tn[0].n51 VGND 0.08671f
C5199 XThR.Tn[0].t25 VGND 0.01383f
C5200 XThR.Tn[0].t34 VGND 0.01514f
C5201 XThR.Tn[0].n52 VGND 0.03697f
C5202 XThR.Tn[0].t47 VGND 0.01378f
C5203 XThR.Tn[0].t29 VGND 0.01509f
C5204 XThR.Tn[0].n53 VGND 0.03846f
C5205 XThR.Tn[0].n54 VGND 0.02702f
C5206 XThR.Tn[0].n56 VGND 0.08671f
C5207 XThR.Tn[0].t17 VGND 0.01383f
C5208 XThR.Tn[0].t53 VGND 0.01514f
C5209 XThR.Tn[0].n57 VGND 0.03697f
C5210 XThR.Tn[0].t38 VGND 0.01378f
C5211 XThR.Tn[0].t49 VGND 0.01509f
C5212 XThR.Tn[0].n58 VGND 0.03846f
C5213 XThR.Tn[0].n59 VGND 0.02702f
C5214 XThR.Tn[0].n61 VGND 0.08671f
C5215 XThR.Tn[0].t37 VGND 0.01383f
C5216 XThR.Tn[0].t31 VGND 0.01514f
C5217 XThR.Tn[0].n62 VGND 0.03697f
C5218 XThR.Tn[0].t56 VGND 0.01378f
C5219 XThR.Tn[0].t19 VGND 0.01509f
C5220 XThR.Tn[0].n63 VGND 0.03846f
C5221 XThR.Tn[0].n64 VGND 0.02702f
C5222 XThR.Tn[0].n66 VGND 0.08671f
C5223 XThR.Tn[0].t69 VGND 0.01383f
C5224 XThR.Tn[0].t65 VGND 0.01514f
C5225 XThR.Tn[0].n67 VGND 0.03697f
C5226 XThR.Tn[0].t27 VGND 0.01378f
C5227 XThR.Tn[0].t57 VGND 0.01509f
C5228 XThR.Tn[0].n68 VGND 0.03846f
C5229 XThR.Tn[0].n69 VGND 0.02702f
C5230 XThR.Tn[0].n71 VGND 0.08671f
C5231 XThR.Tn[0].t22 VGND 0.01383f
C5232 XThR.Tn[0].t16 VGND 0.01514f
C5233 XThR.Tn[0].n72 VGND 0.03697f
C5234 XThR.Tn[0].t45 VGND 0.01378f
C5235 XThR.Tn[0].t73 VGND 0.01509f
C5236 XThR.Tn[0].n73 VGND 0.03846f
C5237 XThR.Tn[0].n74 VGND 0.02702f
C5238 XThR.Tn[0].n76 VGND 0.08671f
C5239 XThR.Tn[0].t42 VGND 0.01383f
C5240 XThR.Tn[0].t36 VGND 0.01514f
C5241 XThR.Tn[0].n77 VGND 0.03697f
C5242 XThR.Tn[0].t62 VGND 0.01378f
C5243 XThR.Tn[0].t30 VGND 0.01509f
C5244 XThR.Tn[0].n78 VGND 0.03846f
C5245 XThR.Tn[0].n79 VGND 0.02702f
C5246 XThR.Tn[0].n81 VGND 0.08671f
C5247 XThR.Tn[0].t18 VGND 0.01383f
C5248 XThR.Tn[0].t32 VGND 0.01514f
C5249 XThR.Tn[0].n82 VGND 0.03697f
C5250 XThR.Tn[0].t39 VGND 0.01378f
C5251 XThR.Tn[0].t20 VGND 0.01509f
C5252 XThR.Tn[0].n83 VGND 0.03846f
C5253 XThR.Tn[0].n84 VGND 0.02702f
C5254 XThR.Tn[0].n86 VGND 0.08671f
C5255 XThR.Tn[0].n87 VGND 0.0788f
C5256 XThR.Tn[0].n88 VGND 0.22563f
C5257 XThR.Tn[7].t7 VGND 0.0118f
C5258 XThR.Tn[7].t4 VGND 0.0118f
C5259 XThR.Tn[7].n0 VGND 0.03641f
C5260 XThR.Tn[7].t6 VGND 0.0118f
C5261 XThR.Tn[7].t5 VGND 0.0118f
C5262 XThR.Tn[7].n1 VGND 0.02606f
C5263 XThR.Tn[7].n2 VGND 0.13363f
C5264 XThR.Tn[7].t2 VGND 0.01815f
C5265 XThR.Tn[7].t3 VGND 0.01815f
C5266 XThR.Tn[7].n3 VGND 0.05527f
C5267 XThR.Tn[7].t1 VGND 0.01815f
C5268 XThR.Tn[7].t0 VGND 0.01815f
C5269 XThR.Tn[7].n4 VGND 0.04021f
C5270 XThR.Tn[7].n5 VGND 0.17693f
C5271 XThR.Tn[7].n6 VGND 0.02205f
C5272 XThR.Tn[7].t53 VGND 0.01419f
C5273 XThR.Tn[7].t45 VGND 0.01553f
C5274 XThR.Tn[7].n7 VGND 0.03793f
C5275 XThR.Tn[7].n8 VGND 0.07287f
C5276 XThR.Tn[7].t8 VGND 0.01419f
C5277 XThR.Tn[7].t60 VGND 0.01553f
C5278 XThR.Tn[7].n9 VGND 0.03793f
C5279 XThR.Tn[7].t26 VGND 0.01414f
C5280 XThR.Tn[7].t38 VGND 0.01548f
C5281 XThR.Tn[7].n10 VGND 0.03947f
C5282 XThR.Tn[7].n11 VGND 0.02773f
C5283 XThR.Tn[7].n13 VGND 0.08897f
C5284 XThR.Tn[7].t47 VGND 0.01419f
C5285 XThR.Tn[7].t37 VGND 0.01553f
C5286 XThR.Tn[7].n14 VGND 0.03793f
C5287 XThR.Tn[7].t66 VGND 0.01414f
C5288 XThR.Tn[7].t15 VGND 0.01548f
C5289 XThR.Tn[7].n15 VGND 0.03947f
C5290 XThR.Tn[7].n16 VGND 0.02773f
C5291 XThR.Tn[7].n18 VGND 0.08897f
C5292 XThR.Tn[7].t62 VGND 0.01419f
C5293 XThR.Tn[7].t55 VGND 0.01553f
C5294 XThR.Tn[7].n19 VGND 0.03793f
C5295 XThR.Tn[7].t18 VGND 0.01414f
C5296 XThR.Tn[7].t32 VGND 0.01548f
C5297 XThR.Tn[7].n20 VGND 0.03947f
C5298 XThR.Tn[7].n21 VGND 0.02773f
C5299 XThR.Tn[7].n23 VGND 0.08897f
C5300 XThR.Tn[7].t25 VGND 0.01419f
C5301 XThR.Tn[7].t21 VGND 0.01553f
C5302 XThR.Tn[7].n24 VGND 0.03793f
C5303 XThR.Tn[7].t50 VGND 0.01414f
C5304 XThR.Tn[7].t63 VGND 0.01548f
C5305 XThR.Tn[7].n25 VGND 0.03947f
C5306 XThR.Tn[7].n26 VGND 0.02773f
C5307 XThR.Tn[7].n28 VGND 0.08897f
C5308 XThR.Tn[7].t65 VGND 0.01419f
C5309 XThR.Tn[7].t56 VGND 0.01553f
C5310 XThR.Tn[7].n29 VGND 0.03793f
C5311 XThR.Tn[7].t19 VGND 0.01414f
C5312 XThR.Tn[7].t34 VGND 0.01548f
C5313 XThR.Tn[7].n30 VGND 0.03947f
C5314 XThR.Tn[7].n31 VGND 0.02773f
C5315 XThR.Tn[7].n33 VGND 0.08897f
C5316 XThR.Tn[7].t40 VGND 0.01419f
C5317 XThR.Tn[7].t11 VGND 0.01553f
C5318 XThR.Tn[7].n34 VGND 0.03793f
C5319 XThR.Tn[7].t58 VGND 0.01414f
C5320 XThR.Tn[7].t54 VGND 0.01548f
C5321 XThR.Tn[7].n35 VGND 0.03947f
C5322 XThR.Tn[7].n36 VGND 0.02773f
C5323 XThR.Tn[7].n38 VGND 0.08897f
C5324 XThR.Tn[7].t9 VGND 0.01419f
C5325 XThR.Tn[7].t68 VGND 0.01553f
C5326 XThR.Tn[7].n39 VGND 0.03793f
C5327 XThR.Tn[7].t27 VGND 0.01414f
C5328 XThR.Tn[7].t46 VGND 0.01548f
C5329 XThR.Tn[7].n40 VGND 0.03947f
C5330 XThR.Tn[7].n41 VGND 0.02773f
C5331 XThR.Tn[7].n43 VGND 0.08897f
C5332 XThR.Tn[7].t14 VGND 0.01419f
C5333 XThR.Tn[7].t20 VGND 0.01553f
C5334 XThR.Tn[7].n44 VGND 0.03793f
C5335 XThR.Tn[7].t31 VGND 0.01414f
C5336 XThR.Tn[7].t61 VGND 0.01548f
C5337 XThR.Tn[7].n45 VGND 0.03947f
C5338 XThR.Tn[7].n46 VGND 0.02773f
C5339 XThR.Tn[7].n48 VGND 0.08897f
C5340 XThR.Tn[7].t29 VGND 0.01419f
C5341 XThR.Tn[7].t39 VGND 0.01553f
C5342 XThR.Tn[7].n49 VGND 0.03793f
C5343 XThR.Tn[7].t52 VGND 0.01414f
C5344 XThR.Tn[7].t16 VGND 0.01548f
C5345 XThR.Tn[7].n50 VGND 0.03947f
C5346 XThR.Tn[7].n51 VGND 0.02773f
C5347 XThR.Tn[7].n53 VGND 0.08897f
C5348 XThR.Tn[7].t23 VGND 0.01419f
C5349 XThR.Tn[7].t57 VGND 0.01553f
C5350 XThR.Tn[7].n54 VGND 0.03793f
C5351 XThR.Tn[7].t43 VGND 0.01414f
C5352 XThR.Tn[7].t36 VGND 0.01548f
C5353 XThR.Tn[7].n55 VGND 0.03947f
C5354 XThR.Tn[7].n56 VGND 0.02773f
C5355 XThR.Tn[7].n58 VGND 0.08897f
C5356 XThR.Tn[7].t42 VGND 0.01419f
C5357 XThR.Tn[7].t33 VGND 0.01553f
C5358 XThR.Tn[7].n59 VGND 0.03793f
C5359 XThR.Tn[7].t59 VGND 0.01414f
C5360 XThR.Tn[7].t10 VGND 0.01548f
C5361 XThR.Tn[7].n60 VGND 0.03947f
C5362 XThR.Tn[7].n61 VGND 0.02773f
C5363 XThR.Tn[7].n63 VGND 0.08897f
C5364 XThR.Tn[7].t12 VGND 0.01419f
C5365 XThR.Tn[7].t69 VGND 0.01553f
C5366 XThR.Tn[7].n64 VGND 0.03793f
C5367 XThR.Tn[7].t30 VGND 0.01414f
C5368 XThR.Tn[7].t48 VGND 0.01548f
C5369 XThR.Tn[7].n65 VGND 0.03947f
C5370 XThR.Tn[7].n66 VGND 0.02773f
C5371 XThR.Tn[7].n68 VGND 0.08897f
C5372 XThR.Tn[7].t28 VGND 0.01419f
C5373 XThR.Tn[7].t22 VGND 0.01553f
C5374 XThR.Tn[7].n69 VGND 0.03793f
C5375 XThR.Tn[7].t51 VGND 0.01414f
C5376 XThR.Tn[7].t64 VGND 0.01548f
C5377 XThR.Tn[7].n70 VGND 0.03947f
C5378 XThR.Tn[7].n71 VGND 0.02773f
C5379 XThR.Tn[7].n73 VGND 0.08897f
C5380 XThR.Tn[7].t49 VGND 0.01419f
C5381 XThR.Tn[7].t41 VGND 0.01553f
C5382 XThR.Tn[7].n74 VGND 0.03793f
C5383 XThR.Tn[7].t67 VGND 0.01414f
C5384 XThR.Tn[7].t17 VGND 0.01548f
C5385 XThR.Tn[7].n75 VGND 0.03947f
C5386 XThR.Tn[7].n76 VGND 0.02773f
C5387 XThR.Tn[7].n78 VGND 0.08897f
C5388 XThR.Tn[7].t24 VGND 0.01419f
C5389 XThR.Tn[7].t35 VGND 0.01553f
C5390 XThR.Tn[7].n79 VGND 0.03793f
C5391 XThR.Tn[7].t44 VGND 0.01414f
C5392 XThR.Tn[7].t13 VGND 0.01548f
C5393 XThR.Tn[7].n80 VGND 0.03947f
C5394 XThR.Tn[7].n81 VGND 0.02773f
C5395 XThR.Tn[7].n83 VGND 0.08897f
C5396 XThR.Tn[7].n84 VGND 0.08086f
C5397 XThR.Tn[7].n85 VGND 0.32824f
C5398 XThR.Tn[11].t5 VGND 0.01248f
C5399 XThR.Tn[11].t2 VGND 0.01248f
C5400 XThR.Tn[11].n0 VGND 0.02496f
C5401 XThR.Tn[11].t4 VGND 0.01248f
C5402 XThR.Tn[11].t0 VGND 0.01248f
C5403 XThR.Tn[11].n1 VGND 0.03112f
C5404 XThR.Tn[11].n2 VGND 0.06279f
C5405 XThR.Tn[11].t8 VGND 0.0192f
C5406 XThR.Tn[11].t10 VGND 0.0192f
C5407 XThR.Tn[11].n3 VGND 0.05829f
C5408 XThR.Tn[11].t9 VGND 0.0192f
C5409 XThR.Tn[11].t11 VGND 0.0192f
C5410 XThR.Tn[11].n4 VGND 0.04268f
C5411 XThR.Tn[11].n5 VGND 0.19406f
C5412 XThR.Tn[11].t3 VGND 0.0192f
C5413 XThR.Tn[11].t7 VGND 0.0192f
C5414 XThR.Tn[11].n6 VGND 0.04148f
C5415 XThR.Tn[11].t1 VGND 0.0192f
C5416 XThR.Tn[11].t6 VGND 0.0192f
C5417 XThR.Tn[11].n7 VGND 0.06313f
C5418 XThR.Tn[11].n8 VGND 0.1753f
C5419 XThR.Tn[11].n9 VGND 0.02347f
C5420 XThR.Tn[11].t56 VGND 0.015f
C5421 XThR.Tn[11].t48 VGND 0.01643f
C5422 XThR.Tn[11].n10 VGND 0.04012f
C5423 XThR.Tn[11].n11 VGND 0.07707f
C5424 XThR.Tn[11].t12 VGND 0.015f
C5425 XThR.Tn[11].t67 VGND 0.01643f
C5426 XThR.Tn[11].n12 VGND 0.04012f
C5427 XThR.Tn[11].t27 VGND 0.01496f
C5428 XThR.Tn[11].t58 VGND 0.01638f
C5429 XThR.Tn[11].n13 VGND 0.04174f
C5430 XThR.Tn[11].n14 VGND 0.02933f
C5431 XThR.Tn[11].n16 VGND 0.09411f
C5432 XThR.Tn[11].t49 VGND 0.015f
C5433 XThR.Tn[11].t41 VGND 0.01643f
C5434 XThR.Tn[11].n17 VGND 0.04012f
C5435 XThR.Tn[11].t65 VGND 0.01496f
C5436 XThR.Tn[11].t36 VGND 0.01638f
C5437 XThR.Tn[11].n18 VGND 0.04174f
C5438 XThR.Tn[11].n19 VGND 0.02933f
C5439 XThR.Tn[11].n21 VGND 0.09411f
C5440 XThR.Tn[11].t68 VGND 0.015f
C5441 XThR.Tn[11].t60 VGND 0.01643f
C5442 XThR.Tn[11].n22 VGND 0.04012f
C5443 XThR.Tn[11].t18 VGND 0.01496f
C5444 XThR.Tn[11].t54 VGND 0.01638f
C5445 XThR.Tn[11].n23 VGND 0.04174f
C5446 XThR.Tn[11].n24 VGND 0.02933f
C5447 XThR.Tn[11].n26 VGND 0.09411f
C5448 XThR.Tn[11].t33 VGND 0.015f
C5449 XThR.Tn[11].t23 VGND 0.01643f
C5450 XThR.Tn[11].n27 VGND 0.04012f
C5451 XThR.Tn[11].t50 VGND 0.01496f
C5452 XThR.Tn[11].t19 VGND 0.01638f
C5453 XThR.Tn[11].n28 VGND 0.04174f
C5454 XThR.Tn[11].n29 VGND 0.02933f
C5455 XThR.Tn[11].n31 VGND 0.09411f
C5456 XThR.Tn[11].t70 VGND 0.015f
C5457 XThR.Tn[11].t62 VGND 0.01643f
C5458 XThR.Tn[11].n32 VGND 0.04012f
C5459 XThR.Tn[11].t21 VGND 0.01496f
C5460 XThR.Tn[11].t55 VGND 0.01638f
C5461 XThR.Tn[11].n33 VGND 0.04174f
C5462 XThR.Tn[11].n34 VGND 0.02933f
C5463 XThR.Tn[11].n36 VGND 0.09411f
C5464 XThR.Tn[11].t44 VGND 0.015f
C5465 XThR.Tn[11].t14 VGND 0.01643f
C5466 XThR.Tn[11].n37 VGND 0.04012f
C5467 XThR.Tn[11].t59 VGND 0.01496f
C5468 XThR.Tn[11].t72 VGND 0.01638f
C5469 XThR.Tn[11].n38 VGND 0.04174f
C5470 XThR.Tn[11].n39 VGND 0.02933f
C5471 XThR.Tn[11].n41 VGND 0.09411f
C5472 XThR.Tn[11].t13 VGND 0.015f
C5473 XThR.Tn[11].t71 VGND 0.01643f
C5474 XThR.Tn[11].n42 VGND 0.04012f
C5475 XThR.Tn[11].t28 VGND 0.01496f
C5476 XThR.Tn[11].t64 VGND 0.01638f
C5477 XThR.Tn[11].n43 VGND 0.04174f
C5478 XThR.Tn[11].n44 VGND 0.02933f
C5479 XThR.Tn[11].n46 VGND 0.09411f
C5480 XThR.Tn[11].t16 VGND 0.015f
C5481 XThR.Tn[11].t22 VGND 0.01643f
C5482 XThR.Tn[11].n47 VGND 0.04012f
C5483 XThR.Tn[11].t32 VGND 0.01496f
C5484 XThR.Tn[11].t17 VGND 0.01638f
C5485 XThR.Tn[11].n48 VGND 0.04174f
C5486 XThR.Tn[11].n49 VGND 0.02933f
C5487 XThR.Tn[11].n51 VGND 0.09411f
C5488 XThR.Tn[11].t35 VGND 0.015f
C5489 XThR.Tn[11].t43 VGND 0.01643f
C5490 XThR.Tn[11].n52 VGND 0.04012f
C5491 XThR.Tn[11].t52 VGND 0.01496f
C5492 XThR.Tn[11].t37 VGND 0.01638f
C5493 XThR.Tn[11].n53 VGND 0.04174f
C5494 XThR.Tn[11].n54 VGND 0.02933f
C5495 XThR.Tn[11].n56 VGND 0.09411f
C5496 XThR.Tn[11].t25 VGND 0.015f
C5497 XThR.Tn[11].t63 VGND 0.01643f
C5498 XThR.Tn[11].n57 VGND 0.04012f
C5499 XThR.Tn[11].t42 VGND 0.01496f
C5500 XThR.Tn[11].t57 VGND 0.01638f
C5501 XThR.Tn[11].n58 VGND 0.04174f
C5502 XThR.Tn[11].n59 VGND 0.02933f
C5503 XThR.Tn[11].n61 VGND 0.09411f
C5504 XThR.Tn[11].t47 VGND 0.015f
C5505 XThR.Tn[11].t39 VGND 0.01643f
C5506 XThR.Tn[11].n62 VGND 0.04012f
C5507 XThR.Tn[11].t61 VGND 0.01496f
C5508 XThR.Tn[11].t29 VGND 0.01638f
C5509 XThR.Tn[11].n63 VGND 0.04174f
C5510 XThR.Tn[11].n64 VGND 0.02933f
C5511 XThR.Tn[11].n66 VGND 0.09411f
C5512 XThR.Tn[11].t15 VGND 0.015f
C5513 XThR.Tn[11].t73 VGND 0.01643f
C5514 XThR.Tn[11].n67 VGND 0.04012f
C5515 XThR.Tn[11].t30 VGND 0.01496f
C5516 XThR.Tn[11].t66 VGND 0.01638f
C5517 XThR.Tn[11].n68 VGND 0.04174f
C5518 XThR.Tn[11].n69 VGND 0.02933f
C5519 XThR.Tn[11].n71 VGND 0.09411f
C5520 XThR.Tn[11].t34 VGND 0.015f
C5521 XThR.Tn[11].t24 VGND 0.01643f
C5522 XThR.Tn[11].n72 VGND 0.04012f
C5523 XThR.Tn[11].t51 VGND 0.01496f
C5524 XThR.Tn[11].t20 VGND 0.01638f
C5525 XThR.Tn[11].n73 VGND 0.04174f
C5526 XThR.Tn[11].n74 VGND 0.02933f
C5527 XThR.Tn[11].n76 VGND 0.09411f
C5528 XThR.Tn[11].t53 VGND 0.015f
C5529 XThR.Tn[11].t46 VGND 0.01643f
C5530 XThR.Tn[11].n77 VGND 0.04012f
C5531 XThR.Tn[11].t69 VGND 0.01496f
C5532 XThR.Tn[11].t38 VGND 0.01638f
C5533 XThR.Tn[11].n78 VGND 0.04174f
C5534 XThR.Tn[11].n79 VGND 0.02933f
C5535 XThR.Tn[11].n81 VGND 0.09411f
C5536 XThR.Tn[11].t26 VGND 0.015f
C5537 XThR.Tn[11].t40 VGND 0.01643f
C5538 XThR.Tn[11].n82 VGND 0.04012f
C5539 XThR.Tn[11].t45 VGND 0.01496f
C5540 XThR.Tn[11].t31 VGND 0.01638f
C5541 XThR.Tn[11].n83 VGND 0.04174f
C5542 XThR.Tn[11].n84 VGND 0.02933f
C5543 XThR.Tn[11].n86 VGND 0.09411f
C5544 XThR.Tn[11].n87 VGND 0.08553f
C5545 XThR.Tn[11].n88 VGND 0.30653f
C5546 XThR.Tn[4].t9 VGND 0.01806f
C5547 XThR.Tn[4].t10 VGND 0.01806f
C5548 XThR.Tn[4].n0 VGND 0.03645f
C5549 XThR.Tn[4].t8 VGND 0.01806f
C5550 XThR.Tn[4].t11 VGND 0.01806f
C5551 XThR.Tn[4].n1 VGND 0.04265f
C5552 XThR.Tn[4].n2 VGND 0.12794f
C5553 XThR.Tn[4].t7 VGND 0.01174f
C5554 XThR.Tn[4].t4 VGND 0.01174f
C5555 XThR.Tn[4].n3 VGND 0.02673f
C5556 XThR.Tn[4].t6 VGND 0.01174f
C5557 XThR.Tn[4].t5 VGND 0.01174f
C5558 XThR.Tn[4].n4 VGND 0.02673f
C5559 XThR.Tn[4].t0 VGND 0.01174f
C5560 XThR.Tn[4].t1 VGND 0.01174f
C5561 XThR.Tn[4].n5 VGND 0.04454f
C5562 XThR.Tn[4].t3 VGND 0.01174f
C5563 XThR.Tn[4].t2 VGND 0.01174f
C5564 XThR.Tn[4].n6 VGND 0.02673f
C5565 XThR.Tn[4].n7 VGND 0.1273f
C5566 XThR.Tn[4].n8 VGND 0.0787f
C5567 XThR.Tn[4].n9 VGND 0.08881f
C5568 XThR.Tn[4].t44 VGND 0.01411f
C5569 XThR.Tn[4].t38 VGND 0.01545f
C5570 XThR.Tn[4].n10 VGND 0.03774f
C5571 XThR.Tn[4].n11 VGND 0.0725f
C5572 XThR.Tn[4].t65 VGND 0.01411f
C5573 XThR.Tn[4].t54 VGND 0.01545f
C5574 XThR.Tn[4].n12 VGND 0.03774f
C5575 XThR.Tn[4].t19 VGND 0.01407f
C5576 XThR.Tn[4].t50 VGND 0.01541f
C5577 XThR.Tn[4].n13 VGND 0.03927f
C5578 XThR.Tn[4].n14 VGND 0.02759f
C5579 XThR.Tn[4].n16 VGND 0.08853f
C5580 XThR.Tn[4].t39 VGND 0.01411f
C5581 XThR.Tn[4].t31 VGND 0.01545f
C5582 XThR.Tn[4].n17 VGND 0.03774f
C5583 XThR.Tn[4].t58 VGND 0.01407f
C5584 XThR.Tn[4].t27 VGND 0.01541f
C5585 XThR.Tn[4].n18 VGND 0.03927f
C5586 XThR.Tn[4].n19 VGND 0.02759f
C5587 XThR.Tn[4].n21 VGND 0.08853f
C5588 XThR.Tn[4].t55 VGND 0.01411f
C5589 XThR.Tn[4].t48 VGND 0.01545f
C5590 XThR.Tn[4].n22 VGND 0.03774f
C5591 XThR.Tn[4].t70 VGND 0.01407f
C5592 XThR.Tn[4].t45 VGND 0.01541f
C5593 XThR.Tn[4].n23 VGND 0.03927f
C5594 XThR.Tn[4].n24 VGND 0.02759f
C5595 XThR.Tn[4].n26 VGND 0.08853f
C5596 XThR.Tn[4].t17 VGND 0.01411f
C5597 XThR.Tn[4].t13 VGND 0.01545f
C5598 XThR.Tn[4].n27 VGND 0.03774f
C5599 XThR.Tn[4].t41 VGND 0.01407f
C5600 XThR.Tn[4].t71 VGND 0.01541f
C5601 XThR.Tn[4].n28 VGND 0.03927f
C5602 XThR.Tn[4].n29 VGND 0.02759f
C5603 XThR.Tn[4].n31 VGND 0.08853f
C5604 XThR.Tn[4].t57 VGND 0.01411f
C5605 XThR.Tn[4].t49 VGND 0.01545f
C5606 XThR.Tn[4].n32 VGND 0.03774f
C5607 XThR.Tn[4].t73 VGND 0.01407f
C5608 XThR.Tn[4].t46 VGND 0.01541f
C5609 XThR.Tn[4].n33 VGND 0.03927f
C5610 XThR.Tn[4].n34 VGND 0.02759f
C5611 XThR.Tn[4].n36 VGND 0.08853f
C5612 XThR.Tn[4].t33 VGND 0.01411f
C5613 XThR.Tn[4].t66 VGND 0.01545f
C5614 XThR.Tn[4].n37 VGND 0.03774f
C5615 XThR.Tn[4].t52 VGND 0.01407f
C5616 XThR.Tn[4].t63 VGND 0.01541f
C5617 XThR.Tn[4].n38 VGND 0.03927f
C5618 XThR.Tn[4].n39 VGND 0.02759f
C5619 XThR.Tn[4].n41 VGND 0.08853f
C5620 XThR.Tn[4].t64 VGND 0.01411f
C5621 XThR.Tn[4].t61 VGND 0.01545f
C5622 XThR.Tn[4].n42 VGND 0.03774f
C5623 XThR.Tn[4].t18 VGND 0.01407f
C5624 XThR.Tn[4].t56 VGND 0.01541f
C5625 XThR.Tn[4].n43 VGND 0.03927f
C5626 XThR.Tn[4].n44 VGND 0.02759f
C5627 XThR.Tn[4].n46 VGND 0.08853f
C5628 XThR.Tn[4].t68 VGND 0.01411f
C5629 XThR.Tn[4].t12 VGND 0.01545f
C5630 XThR.Tn[4].n47 VGND 0.03774f
C5631 XThR.Tn[4].t25 VGND 0.01407f
C5632 XThR.Tn[4].t69 VGND 0.01541f
C5633 XThR.Tn[4].n48 VGND 0.03927f
C5634 XThR.Tn[4].n49 VGND 0.02759f
C5635 XThR.Tn[4].n51 VGND 0.08853f
C5636 XThR.Tn[4].t22 VGND 0.01411f
C5637 XThR.Tn[4].t32 VGND 0.01545f
C5638 XThR.Tn[4].n52 VGND 0.03774f
C5639 XThR.Tn[4].t43 VGND 0.01407f
C5640 XThR.Tn[4].t29 VGND 0.01541f
C5641 XThR.Tn[4].n53 VGND 0.03927f
C5642 XThR.Tn[4].n54 VGND 0.02759f
C5643 XThR.Tn[4].n56 VGND 0.08853f
C5644 XThR.Tn[4].t15 VGND 0.01411f
C5645 XThR.Tn[4].t51 VGND 0.01545f
C5646 XThR.Tn[4].n57 VGND 0.03774f
C5647 XThR.Tn[4].t36 VGND 0.01407f
C5648 XThR.Tn[4].t47 VGND 0.01541f
C5649 XThR.Tn[4].n58 VGND 0.03927f
C5650 XThR.Tn[4].n59 VGND 0.02759f
C5651 XThR.Tn[4].n61 VGND 0.08853f
C5652 XThR.Tn[4].t35 VGND 0.01411f
C5653 XThR.Tn[4].t26 VGND 0.01545f
C5654 XThR.Tn[4].n62 VGND 0.03774f
C5655 XThR.Tn[4].t53 VGND 0.01407f
C5656 XThR.Tn[4].t21 VGND 0.01541f
C5657 XThR.Tn[4].n63 VGND 0.03927f
C5658 XThR.Tn[4].n64 VGND 0.02759f
C5659 XThR.Tn[4].n66 VGND 0.08853f
C5660 XThR.Tn[4].t67 VGND 0.01411f
C5661 XThR.Tn[4].t62 VGND 0.01545f
C5662 XThR.Tn[4].n67 VGND 0.03774f
C5663 XThR.Tn[4].t23 VGND 0.01407f
C5664 XThR.Tn[4].t59 VGND 0.01541f
C5665 XThR.Tn[4].n68 VGND 0.03927f
C5666 XThR.Tn[4].n69 VGND 0.02759f
C5667 XThR.Tn[4].n71 VGND 0.08853f
C5668 XThR.Tn[4].t20 VGND 0.01411f
C5669 XThR.Tn[4].t14 VGND 0.01545f
C5670 XThR.Tn[4].n72 VGND 0.03774f
C5671 XThR.Tn[4].t42 VGND 0.01407f
C5672 XThR.Tn[4].t72 VGND 0.01541f
C5673 XThR.Tn[4].n73 VGND 0.03927f
C5674 XThR.Tn[4].n74 VGND 0.02759f
C5675 XThR.Tn[4].n76 VGND 0.08853f
C5676 XThR.Tn[4].t40 VGND 0.01411f
C5677 XThR.Tn[4].t34 VGND 0.01545f
C5678 XThR.Tn[4].n77 VGND 0.03774f
C5679 XThR.Tn[4].t60 VGND 0.01407f
C5680 XThR.Tn[4].t30 VGND 0.01541f
C5681 XThR.Tn[4].n78 VGND 0.03927f
C5682 XThR.Tn[4].n79 VGND 0.02759f
C5683 XThR.Tn[4].n81 VGND 0.08853f
C5684 XThR.Tn[4].t16 VGND 0.01411f
C5685 XThR.Tn[4].t28 VGND 0.01545f
C5686 XThR.Tn[4].n82 VGND 0.03774f
C5687 XThR.Tn[4].t37 VGND 0.01407f
C5688 XThR.Tn[4].t24 VGND 0.01541f
C5689 XThR.Tn[4].n83 VGND 0.03927f
C5690 XThR.Tn[4].n84 VGND 0.02759f
C5691 XThR.Tn[4].n86 VGND 0.08853f
C5692 XThR.Tn[4].n87 VGND 0.08045f
C5693 XThR.Tn[4].n88 VGND 0.15199f
C5694 XA.Cn[7].n0 VGND 0.02617f
C5695 XA.Cn[7].n1 VGND 0.01873f
C5696 XA.Cn[7].n2 VGND 0.09263f
C5697 XA.Cn[7].t0 VGND 0.01305f
C5698 XA.Cn[7].t3 VGND 0.01305f
C5699 XA.Cn[7].n3 VGND 0.0281f
C5700 XA.Cn[7].t2 VGND 0.01305f
C5701 XA.Cn[7].t1 VGND 0.01305f
C5702 XA.Cn[7].n4 VGND 0.04266f
C5703 XA.Cn[7].n5 VGND 0.12542f
C5704 XA.Cn[7].t8 VGND 0.01034f
C5705 XA.Cn[7].t11 VGND 0.01129f
C5706 XA.Cn[7].n6 VGND 0.02522f
C5707 XA.Cn[7].n7 VGND 0.01441f
C5708 XA.Cn[7].n8 VGND 0.01753f
C5709 XA.Cn[7].t25 VGND 0.01034f
C5710 XA.Cn[7].t30 VGND 0.01129f
C5711 XA.Cn[7].n9 VGND 0.02522f
C5712 XA.Cn[7].n10 VGND 0.01441f
C5713 XA.Cn[7].n11 VGND 0.08328f
C5714 XA.Cn[7].t27 VGND 0.01034f
C5715 XA.Cn[7].t34 VGND 0.01129f
C5716 XA.Cn[7].n12 VGND 0.02522f
C5717 XA.Cn[7].n13 VGND 0.01441f
C5718 XA.Cn[7].n14 VGND 0.08328f
C5719 XA.Cn[7].t29 VGND 0.01034f
C5720 XA.Cn[7].t35 VGND 0.01129f
C5721 XA.Cn[7].n15 VGND 0.02522f
C5722 XA.Cn[7].n16 VGND 0.01441f
C5723 XA.Cn[7].n17 VGND 0.08328f
C5724 XA.Cn[7].t18 VGND 0.01034f
C5725 XA.Cn[7].t22 VGND 0.01129f
C5726 XA.Cn[7].n18 VGND 0.02522f
C5727 XA.Cn[7].n19 VGND 0.01441f
C5728 XA.Cn[7].n20 VGND 0.08328f
C5729 XA.Cn[7].t20 VGND 0.01034f
C5730 XA.Cn[7].t23 VGND 0.01129f
C5731 XA.Cn[7].n21 VGND 0.02522f
C5732 XA.Cn[7].n22 VGND 0.01441f
C5733 XA.Cn[7].n23 VGND 0.08328f
C5734 XA.Cn[7].t33 VGND 0.01034f
C5735 XA.Cn[7].t39 VGND 0.01129f
C5736 XA.Cn[7].n24 VGND 0.02522f
C5737 XA.Cn[7].n25 VGND 0.01441f
C5738 XA.Cn[7].n26 VGND 0.08328f
C5739 XA.Cn[7].t10 VGND 0.01034f
C5740 XA.Cn[7].t14 VGND 0.01129f
C5741 XA.Cn[7].n27 VGND 0.02522f
C5742 XA.Cn[7].n28 VGND 0.01441f
C5743 XA.Cn[7].n29 VGND 0.08328f
C5744 XA.Cn[7].t12 VGND 0.01034f
C5745 XA.Cn[7].t16 VGND 0.01129f
C5746 XA.Cn[7].n30 VGND 0.02522f
C5747 XA.Cn[7].n31 VGND 0.01441f
C5748 XA.Cn[7].n32 VGND 0.08328f
C5749 XA.Cn[7].t31 VGND 0.01034f
C5750 XA.Cn[7].t36 VGND 0.01129f
C5751 XA.Cn[7].n33 VGND 0.02522f
C5752 XA.Cn[7].n34 VGND 0.01441f
C5753 XA.Cn[7].n35 VGND 0.08328f
C5754 XA.Cn[7].t32 VGND 0.01034f
C5755 XA.Cn[7].t38 VGND 0.01129f
C5756 XA.Cn[7].n36 VGND 0.02522f
C5757 XA.Cn[7].n37 VGND 0.01441f
C5758 XA.Cn[7].n38 VGND 0.08328f
C5759 XA.Cn[7].t13 VGND 0.01034f
C5760 XA.Cn[7].t17 VGND 0.01129f
C5761 XA.Cn[7].n39 VGND 0.02522f
C5762 XA.Cn[7].n40 VGND 0.01441f
C5763 XA.Cn[7].n41 VGND 0.08328f
C5764 XA.Cn[7].t21 VGND 0.01034f
C5765 XA.Cn[7].t26 VGND 0.01129f
C5766 XA.Cn[7].n42 VGND 0.02522f
C5767 XA.Cn[7].n43 VGND 0.01441f
C5768 XA.Cn[7].n44 VGND 0.08328f
C5769 XA.Cn[7].t24 VGND 0.01034f
C5770 XA.Cn[7].t28 VGND 0.01129f
C5771 XA.Cn[7].n45 VGND 0.02522f
C5772 XA.Cn[7].n46 VGND 0.01441f
C5773 XA.Cn[7].n47 VGND 0.08328f
C5774 XA.Cn[7].t37 VGND 0.01034f
C5775 XA.Cn[7].t9 VGND 0.01129f
C5776 XA.Cn[7].n48 VGND 0.02522f
C5777 XA.Cn[7].n49 VGND 0.01441f
C5778 XA.Cn[7].n50 VGND 0.08328f
C5779 XA.Cn[7].t15 VGND 0.01034f
C5780 XA.Cn[7].t19 VGND 0.01129f
C5781 XA.Cn[7].n51 VGND 0.02522f
C5782 XA.Cn[7].n52 VGND 0.01441f
C5783 XA.Cn[7].n53 VGND 0.08328f
C5784 XA.Cn[7].n54 VGND 0.52699f
C5785 XA.Cn[7].n55 VGND 0.03388f
C5786 XA.Cn[7].n56 VGND 0.01561f
C5787 XThR.Tn[1].t4 VGND 0.01794f
C5788 XThR.Tn[1].t5 VGND 0.01794f
C5789 XThR.Tn[1].n0 VGND 0.03622f
C5790 XThR.Tn[1].t7 VGND 0.01794f
C5791 XThR.Tn[1].t6 VGND 0.01794f
C5792 XThR.Tn[1].n1 VGND 0.04238f
C5793 XThR.Tn[1].n2 VGND 0.11863f
C5794 XThR.Tn[1].t11 VGND 0.01166f
C5795 XThR.Tn[1].t8 VGND 0.01166f
C5796 XThR.Tn[1].n3 VGND 0.02656f
C5797 XThR.Tn[1].t10 VGND 0.01166f
C5798 XThR.Tn[1].t9 VGND 0.01166f
C5799 XThR.Tn[1].n4 VGND 0.02656f
C5800 XThR.Tn[1].t2 VGND 0.01166f
C5801 XThR.Tn[1].t1 VGND 0.01166f
C5802 XThR.Tn[1].n5 VGND 0.02656f
C5803 XThR.Tn[1].t3 VGND 0.01166f
C5804 XThR.Tn[1].t0 VGND 0.01166f
C5805 XThR.Tn[1].n6 VGND 0.04425f
C5806 XThR.Tn[1].n7 VGND 0.12648f
C5807 XThR.Tn[1].n8 VGND 0.07819f
C5808 XThR.Tn[1].n9 VGND 0.08824f
C5809 XThR.Tn[1].t24 VGND 0.01402f
C5810 XThR.Tn[1].t18 VGND 0.01536f
C5811 XThR.Tn[1].n10 VGND 0.0375f
C5812 XThR.Tn[1].n11 VGND 0.07203f
C5813 XThR.Tn[1].t44 VGND 0.01402f
C5814 XThR.Tn[1].t34 VGND 0.01536f
C5815 XThR.Tn[1].n12 VGND 0.0375f
C5816 XThR.Tn[1].t61 VGND 0.01398f
C5817 XThR.Tn[1].t30 VGND 0.01531f
C5818 XThR.Tn[1].n13 VGND 0.03901f
C5819 XThR.Tn[1].n14 VGND 0.02741f
C5820 XThR.Tn[1].n16 VGND 0.08795f
C5821 XThR.Tn[1].t19 VGND 0.01402f
C5822 XThR.Tn[1].t73 VGND 0.01536f
C5823 XThR.Tn[1].n17 VGND 0.0375f
C5824 XThR.Tn[1].t38 VGND 0.01398f
C5825 XThR.Tn[1].t69 VGND 0.01531f
C5826 XThR.Tn[1].n18 VGND 0.03901f
C5827 XThR.Tn[1].n19 VGND 0.02741f
C5828 XThR.Tn[1].n21 VGND 0.08795f
C5829 XThR.Tn[1].t35 VGND 0.01402f
C5830 XThR.Tn[1].t28 VGND 0.01536f
C5831 XThR.Tn[1].n22 VGND 0.0375f
C5832 XThR.Tn[1].t50 VGND 0.01398f
C5833 XThR.Tn[1].t25 VGND 0.01531f
C5834 XThR.Tn[1].n23 VGND 0.03901f
C5835 XThR.Tn[1].n24 VGND 0.02741f
C5836 XThR.Tn[1].n26 VGND 0.08795f
C5837 XThR.Tn[1].t59 VGND 0.01402f
C5838 XThR.Tn[1].t55 VGND 0.01536f
C5839 XThR.Tn[1].n27 VGND 0.0375f
C5840 XThR.Tn[1].t21 VGND 0.01398f
C5841 XThR.Tn[1].t51 VGND 0.01531f
C5842 XThR.Tn[1].n28 VGND 0.03901f
C5843 XThR.Tn[1].n29 VGND 0.02741f
C5844 XThR.Tn[1].n31 VGND 0.08795f
C5845 XThR.Tn[1].t37 VGND 0.01402f
C5846 XThR.Tn[1].t29 VGND 0.01536f
C5847 XThR.Tn[1].n32 VGND 0.0375f
C5848 XThR.Tn[1].t53 VGND 0.01398f
C5849 XThR.Tn[1].t26 VGND 0.01531f
C5850 XThR.Tn[1].n33 VGND 0.03901f
C5851 XThR.Tn[1].n34 VGND 0.02741f
C5852 XThR.Tn[1].n36 VGND 0.08795f
C5853 XThR.Tn[1].t13 VGND 0.01402f
C5854 XThR.Tn[1].t46 VGND 0.01536f
C5855 XThR.Tn[1].n37 VGND 0.0375f
C5856 XThR.Tn[1].t32 VGND 0.01398f
C5857 XThR.Tn[1].t43 VGND 0.01531f
C5858 XThR.Tn[1].n38 VGND 0.03901f
C5859 XThR.Tn[1].n39 VGND 0.02741f
C5860 XThR.Tn[1].n41 VGND 0.08795f
C5861 XThR.Tn[1].t45 VGND 0.01402f
C5862 XThR.Tn[1].t41 VGND 0.01536f
C5863 XThR.Tn[1].n42 VGND 0.0375f
C5864 XThR.Tn[1].t60 VGND 0.01398f
C5865 XThR.Tn[1].t36 VGND 0.01531f
C5866 XThR.Tn[1].n43 VGND 0.03901f
C5867 XThR.Tn[1].n44 VGND 0.02741f
C5868 XThR.Tn[1].n46 VGND 0.08795f
C5869 XThR.Tn[1].t48 VGND 0.01402f
C5870 XThR.Tn[1].t54 VGND 0.01536f
C5871 XThR.Tn[1].n47 VGND 0.0375f
C5872 XThR.Tn[1].t67 VGND 0.01398f
C5873 XThR.Tn[1].t49 VGND 0.01531f
C5874 XThR.Tn[1].n48 VGND 0.03901f
C5875 XThR.Tn[1].n49 VGND 0.02741f
C5876 XThR.Tn[1].n51 VGND 0.08795f
C5877 XThR.Tn[1].t64 VGND 0.01402f
C5878 XThR.Tn[1].t12 VGND 0.01536f
C5879 XThR.Tn[1].n52 VGND 0.0375f
C5880 XThR.Tn[1].t23 VGND 0.01398f
C5881 XThR.Tn[1].t71 VGND 0.01531f
C5882 XThR.Tn[1].n53 VGND 0.03901f
C5883 XThR.Tn[1].n54 VGND 0.02741f
C5884 XThR.Tn[1].n56 VGND 0.08795f
C5885 XThR.Tn[1].t57 VGND 0.01402f
C5886 XThR.Tn[1].t31 VGND 0.01536f
C5887 XThR.Tn[1].n57 VGND 0.0375f
C5888 XThR.Tn[1].t16 VGND 0.01398f
C5889 XThR.Tn[1].t27 VGND 0.01531f
C5890 XThR.Tn[1].n58 VGND 0.03901f
C5891 XThR.Tn[1].n59 VGND 0.02741f
C5892 XThR.Tn[1].n61 VGND 0.08795f
C5893 XThR.Tn[1].t15 VGND 0.01402f
C5894 XThR.Tn[1].t68 VGND 0.01536f
C5895 XThR.Tn[1].n62 VGND 0.0375f
C5896 XThR.Tn[1].t33 VGND 0.01398f
C5897 XThR.Tn[1].t63 VGND 0.01531f
C5898 XThR.Tn[1].n63 VGND 0.03901f
C5899 XThR.Tn[1].n64 VGND 0.02741f
C5900 XThR.Tn[1].n66 VGND 0.08795f
C5901 XThR.Tn[1].t47 VGND 0.01402f
C5902 XThR.Tn[1].t42 VGND 0.01536f
C5903 XThR.Tn[1].n67 VGND 0.0375f
C5904 XThR.Tn[1].t65 VGND 0.01398f
C5905 XThR.Tn[1].t39 VGND 0.01531f
C5906 XThR.Tn[1].n68 VGND 0.03901f
C5907 XThR.Tn[1].n69 VGND 0.02741f
C5908 XThR.Tn[1].n71 VGND 0.08795f
C5909 XThR.Tn[1].t62 VGND 0.01402f
C5910 XThR.Tn[1].t56 VGND 0.01536f
C5911 XThR.Tn[1].n72 VGND 0.0375f
C5912 XThR.Tn[1].t22 VGND 0.01398f
C5913 XThR.Tn[1].t52 VGND 0.01531f
C5914 XThR.Tn[1].n73 VGND 0.03901f
C5915 XThR.Tn[1].n74 VGND 0.02741f
C5916 XThR.Tn[1].n76 VGND 0.08795f
C5917 XThR.Tn[1].t20 VGND 0.01402f
C5918 XThR.Tn[1].t14 VGND 0.01536f
C5919 XThR.Tn[1].n77 VGND 0.0375f
C5920 XThR.Tn[1].t40 VGND 0.01398f
C5921 XThR.Tn[1].t72 VGND 0.01531f
C5922 XThR.Tn[1].n78 VGND 0.03901f
C5923 XThR.Tn[1].n79 VGND 0.02741f
C5924 XThR.Tn[1].n81 VGND 0.08795f
C5925 XThR.Tn[1].t58 VGND 0.01402f
C5926 XThR.Tn[1].t70 VGND 0.01536f
C5927 XThR.Tn[1].n82 VGND 0.0375f
C5928 XThR.Tn[1].t17 VGND 0.01398f
C5929 XThR.Tn[1].t66 VGND 0.01531f
C5930 XThR.Tn[1].n83 VGND 0.03901f
C5931 XThR.Tn[1].n84 VGND 0.02741f
C5932 XThR.Tn[1].n86 VGND 0.08795f
C5933 XThR.Tn[1].n87 VGND 0.07993f
C5934 XThR.Tn[1].n88 VGND 0.23008f
C5935 XThR.Tn[1].n89 VGND 0.03755f
C5936 XA.Cn[8].n0 VGND 0.02379f
C5937 XA.Cn[8].n1 VGND 0.01907f
C5938 XA.Cn[8].n2 VGND 0.04799f
C5939 XA.Cn[8].t43 VGND 0.01163f
C5940 XA.Cn[8].t41 VGND 0.0127f
C5941 XA.Cn[8].n3 VGND 0.02837f
C5942 XA.Cn[8].n4 VGND 0.01621f
C5943 XA.Cn[8].n5 VGND 0.01972f
C5944 XA.Cn[8].t29 VGND 0.01163f
C5945 XA.Cn[8].t26 VGND 0.0127f
C5946 XA.Cn[8].n6 VGND 0.02837f
C5947 XA.Cn[8].n7 VGND 0.01621f
C5948 XA.Cn[8].n8 VGND 0.09367f
C5949 XA.Cn[8].t34 VGND 0.01163f
C5950 XA.Cn[8].t28 VGND 0.0127f
C5951 XA.Cn[8].n9 VGND 0.02837f
C5952 XA.Cn[8].n10 VGND 0.01621f
C5953 XA.Cn[8].n11 VGND 0.09367f
C5954 XA.Cn[8].t35 VGND 0.01163f
C5955 XA.Cn[8].t30 VGND 0.0127f
C5956 XA.Cn[8].n12 VGND 0.02837f
C5957 XA.Cn[8].n13 VGND 0.01621f
C5958 XA.Cn[8].n14 VGND 0.09367f
C5959 XA.Cn[8].t22 VGND 0.01163f
C5960 XA.Cn[8].t19 VGND 0.0127f
C5961 XA.Cn[8].n15 VGND 0.02837f
C5962 XA.Cn[8].n16 VGND 0.01621f
C5963 XA.Cn[8].n17 VGND 0.09367f
C5964 XA.Cn[8].t23 VGND 0.01163f
C5965 XA.Cn[8].t20 VGND 0.0127f
C5966 XA.Cn[8].n18 VGND 0.02837f
C5967 XA.Cn[8].n19 VGND 0.01621f
C5968 XA.Cn[8].n20 VGND 0.09367f
C5969 XA.Cn[8].t39 VGND 0.01163f
C5970 XA.Cn[8].t33 VGND 0.0127f
C5971 XA.Cn[8].n21 VGND 0.02837f
C5972 XA.Cn[8].n22 VGND 0.01621f
C5973 XA.Cn[8].n23 VGND 0.09367f
C5974 XA.Cn[8].t14 VGND 0.01163f
C5975 XA.Cn[8].t42 VGND 0.0127f
C5976 XA.Cn[8].n24 VGND 0.02837f
C5977 XA.Cn[8].n25 VGND 0.01621f
C5978 XA.Cn[8].n26 VGND 0.09367f
C5979 XA.Cn[8].t16 VGND 0.01163f
C5980 XA.Cn[8].t12 VGND 0.0127f
C5981 XA.Cn[8].n27 VGND 0.02837f
C5982 XA.Cn[8].n28 VGND 0.01621f
C5983 XA.Cn[8].n29 VGND 0.09367f
C5984 XA.Cn[8].t36 VGND 0.01163f
C5985 XA.Cn[8].t31 VGND 0.0127f
C5986 XA.Cn[8].n30 VGND 0.02837f
C5987 XA.Cn[8].n31 VGND 0.01621f
C5988 XA.Cn[8].n32 VGND 0.09367f
C5989 XA.Cn[8].t38 VGND 0.01163f
C5990 XA.Cn[8].t32 VGND 0.0127f
C5991 XA.Cn[8].n33 VGND 0.02837f
C5992 XA.Cn[8].n34 VGND 0.01621f
C5993 XA.Cn[8].n35 VGND 0.09367f
C5994 XA.Cn[8].t17 VGND 0.01163f
C5995 XA.Cn[8].t13 VGND 0.0127f
C5996 XA.Cn[8].n36 VGND 0.02837f
C5997 XA.Cn[8].n37 VGND 0.01621f
C5998 XA.Cn[8].n38 VGND 0.09367f
C5999 XA.Cn[8].t25 VGND 0.01163f
C6000 XA.Cn[8].t21 VGND 0.0127f
C6001 XA.Cn[8].n39 VGND 0.02837f
C6002 XA.Cn[8].n40 VGND 0.01621f
C6003 XA.Cn[8].n41 VGND 0.09367f
C6004 XA.Cn[8].t27 VGND 0.01163f
C6005 XA.Cn[8].t24 VGND 0.0127f
C6006 XA.Cn[8].n42 VGND 0.02837f
C6007 XA.Cn[8].n43 VGND 0.01621f
C6008 XA.Cn[8].n44 VGND 0.09367f
C6009 XA.Cn[8].t40 VGND 0.01163f
C6010 XA.Cn[8].t37 VGND 0.0127f
C6011 XA.Cn[8].n45 VGND 0.02837f
C6012 XA.Cn[8].n46 VGND 0.01621f
C6013 XA.Cn[8].n47 VGND 0.09367f
C6014 XA.Cn[8].t18 VGND 0.01163f
C6015 XA.Cn[8].t15 VGND 0.0127f
C6016 XA.Cn[8].n48 VGND 0.02837f
C6017 XA.Cn[8].n49 VGND 0.01621f
C6018 XA.Cn[8].n50 VGND 0.09367f
C6019 XA.Cn[8].n51 VGND 0.04332f
C6020 XA.Cn[8].n52 VGND 0.41007f
C6021 XA.Cn[8].n53 VGND 0.03291f
C6022 XA.Cn[8].t1 VGND 0.01467f
C6023 XA.Cn[8].t2 VGND 0.01467f
C6024 XA.Cn[8].n54 VGND 0.0317f
C6025 XA.Cn[8].t0 VGND 0.01467f
C6026 XA.Cn[8].t3 VGND 0.01467f
C6027 XA.Cn[8].n55 VGND 0.04825f
C6028 XA.Cn[8].n56 VGND 0.13407f
C6029 XA.Cn[8].n57 VGND 0.02108f
C6030 XA.Cn[8].t8 VGND 0.01467f
C6031 XA.Cn[8].t11 VGND 0.01467f
C6032 XA.Cn[8].n58 VGND 0.04455f
C6033 XA.Cn[8].t10 VGND 0.01467f
C6034 XA.Cn[8].t9 VGND 0.01467f
C6035 XA.Cn[8].n59 VGND 0.03262f
C6036 XA.Cn[8].n60 VGND 0.14517f
C6037 thermo15c_0.XTB1.Y.t1 VGND 0.03224f
C6038 thermo15c_0.XTB1.Y.n0 VGND 0.02084f
C6039 thermo15c_0.XTB1.Y.n1 VGND 0.02659f
C6040 thermo15c_0.XTB1.Y.t2 VGND 0.01618f
C6041 thermo15c_0.XTB1.Y.t0 VGND 0.01618f
C6042 thermo15c_0.XTB1.Y.n2 VGND 0.03473f
C6043 thermo15c_0.XTB1.Y.t17 VGND 0.02517f
C6044 thermo15c_0.XTB1.Y.t5 VGND 0.01483f
C6045 thermo15c_0.XTB1.Y.n3 VGND 0.02997f
C6046 thermo15c_0.XTB1.Y.t6 VGND 0.02517f
C6047 thermo15c_0.XTB1.Y.t12 VGND 0.01483f
C6048 thermo15c_0.XTB1.Y.n4 VGND 0.01542f
C6049 thermo15c_0.XTB1.Y.t8 VGND 0.02517f
C6050 thermo15c_0.XTB1.Y.t13 VGND 0.01483f
C6051 thermo15c_0.XTB1.Y.n5 VGND 0.03313f
C6052 thermo15c_0.XTB1.Y.t11 VGND 0.02517f
C6053 thermo15c_0.XTB1.Y.t16 VGND 0.01483f
C6054 thermo15c_0.XTB1.Y.n6 VGND 0.03076f
C6055 thermo15c_0.XTB1.Y.n7 VGND 0.01871f
C6056 thermo15c_0.XTB1.Y.n8 VGND 0.03098f
C6057 thermo15c_0.XTB1.Y.n9 VGND 0.01198f
C6058 thermo15c_0.XTB1.Y.n10 VGND 0.01463f
C6059 thermo15c_0.XTB1.Y.n11 VGND 0.03313f
C6060 thermo15c_0.XTB1.Y.n12 VGND 0.01661f
C6061 thermo15c_0.XTB1.Y.n13 VGND 0.02824f
C6062 thermo15c_0.XTB1.Y.t18 VGND 0.02517f
C6063 thermo15c_0.XTB1.Y.t9 VGND 0.01483f
C6064 thermo15c_0.XTB1.Y.n14 VGND 0.03392f
C6065 thermo15c_0.XTB1.Y.t7 VGND 0.02517f
C6066 thermo15c_0.XTB1.Y.t15 VGND 0.01483f
C6067 thermo15c_0.XTB1.Y.t14 VGND 0.02517f
C6068 thermo15c_0.XTB1.Y.t3 VGND 0.01483f
C6069 thermo15c_0.XTB1.Y.t10 VGND 0.02517f
C6070 thermo15c_0.XTB1.Y.t4 VGND 0.01483f
C6071 thermo15c_0.XTB1.Y.n15 VGND 0.04223f
C6072 thermo15c_0.XTB1.Y.n16 VGND 0.0446f
C6073 thermo15c_0.XTB1.Y.n17 VGND 0.01719f
C6074 thermo15c_0.XTB1.Y.n18 VGND 0.0363f
C6075 thermo15c_0.XTB1.Y.n19 VGND 0.01661f
C6076 thermo15c_0.XTB1.Y.n20 VGND 0.01378f
C6077 thermo15c_0.XTB1.Y.n21 VGND 0.77148f
C6078 thermo15c_0.XTB1.Y.n22 VGND 0.07634f
C6079 XA.Cn[14].n0 VGND 0.02301f
C6080 XA.Cn[14].n1 VGND 0.01845f
C6081 XA.Cn[14].n2 VGND 0.04642f
C6082 XA.Cn[14].t43 VGND 0.01125f
C6083 XA.Cn[14].t38 VGND 0.01229f
C6084 XA.Cn[14].n3 VGND 0.02744f
C6085 XA.Cn[14].n4 VGND 0.01568f
C6086 XA.Cn[14].n5 VGND 0.01907f
C6087 XA.Cn[14].t29 VGND 0.01125f
C6088 XA.Cn[14].t22 VGND 0.01229f
C6089 XA.Cn[14].n6 VGND 0.02744f
C6090 XA.Cn[14].n7 VGND 0.01568f
C6091 XA.Cn[14].n8 VGND 0.09061f
C6092 XA.Cn[14].t32 VGND 0.01125f
C6093 XA.Cn[14].t25 VGND 0.01229f
C6094 XA.Cn[14].n9 VGND 0.02744f
C6095 XA.Cn[14].n10 VGND 0.01568f
C6096 XA.Cn[14].n11 VGND 0.09061f
C6097 XA.Cn[14].t34 VGND 0.01125f
C6098 XA.Cn[14].t26 VGND 0.01229f
C6099 XA.Cn[14].n12 VGND 0.02744f
C6100 XA.Cn[14].n13 VGND 0.01568f
C6101 XA.Cn[14].n14 VGND 0.09061f
C6102 XA.Cn[14].t20 VGND 0.01125f
C6103 XA.Cn[14].t14 VGND 0.01229f
C6104 XA.Cn[14].n15 VGND 0.02744f
C6105 XA.Cn[14].n16 VGND 0.01568f
C6106 XA.Cn[14].n17 VGND 0.09061f
C6107 XA.Cn[14].t23 VGND 0.01125f
C6108 XA.Cn[14].t17 VGND 0.01229f
C6109 XA.Cn[14].n18 VGND 0.02744f
C6110 XA.Cn[14].n19 VGND 0.01568f
C6111 XA.Cn[14].n20 VGND 0.09061f
C6112 XA.Cn[14].t37 VGND 0.01125f
C6113 XA.Cn[14].t31 VGND 0.01229f
C6114 XA.Cn[14].n21 VGND 0.02744f
C6115 XA.Cn[14].n22 VGND 0.01568f
C6116 XA.Cn[14].n23 VGND 0.09061f
C6117 XA.Cn[14].t13 VGND 0.01125f
C6118 XA.Cn[14].t39 VGND 0.01229f
C6119 XA.Cn[14].n24 VGND 0.02744f
C6120 XA.Cn[14].n25 VGND 0.01568f
C6121 XA.Cn[14].n26 VGND 0.09061f
C6122 XA.Cn[14].t15 VGND 0.01125f
C6123 XA.Cn[14].t41 VGND 0.01229f
C6124 XA.Cn[14].n27 VGND 0.02744f
C6125 XA.Cn[14].n28 VGND 0.01568f
C6126 XA.Cn[14].n29 VGND 0.09061f
C6127 XA.Cn[14].t35 VGND 0.01125f
C6128 XA.Cn[14].t27 VGND 0.01229f
C6129 XA.Cn[14].n30 VGND 0.02744f
C6130 XA.Cn[14].n31 VGND 0.01568f
C6131 XA.Cn[14].n32 VGND 0.09061f
C6132 XA.Cn[14].t36 VGND 0.01125f
C6133 XA.Cn[14].t30 VGND 0.01229f
C6134 XA.Cn[14].n33 VGND 0.02744f
C6135 XA.Cn[14].n34 VGND 0.01568f
C6136 XA.Cn[14].n35 VGND 0.09061f
C6137 XA.Cn[14].t16 VGND 0.01125f
C6138 XA.Cn[14].t42 VGND 0.01229f
C6139 XA.Cn[14].n36 VGND 0.02744f
C6140 XA.Cn[14].n37 VGND 0.01568f
C6141 XA.Cn[14].n38 VGND 0.09061f
C6142 XA.Cn[14].t24 VGND 0.01125f
C6143 XA.Cn[14].t19 VGND 0.01229f
C6144 XA.Cn[14].n39 VGND 0.02744f
C6145 XA.Cn[14].n40 VGND 0.01568f
C6146 XA.Cn[14].n41 VGND 0.09061f
C6147 XA.Cn[14].t28 VGND 0.01125f
C6148 XA.Cn[14].t21 VGND 0.01229f
C6149 XA.Cn[14].n42 VGND 0.02744f
C6150 XA.Cn[14].n43 VGND 0.01568f
C6151 XA.Cn[14].n44 VGND 0.09061f
C6152 XA.Cn[14].t40 VGND 0.01125f
C6153 XA.Cn[14].t33 VGND 0.01229f
C6154 XA.Cn[14].n45 VGND 0.02744f
C6155 XA.Cn[14].n46 VGND 0.01568f
C6156 XA.Cn[14].n47 VGND 0.09061f
C6157 XA.Cn[14].t18 VGND 0.01125f
C6158 XA.Cn[14].t12 VGND 0.01229f
C6159 XA.Cn[14].n48 VGND 0.02744f
C6160 XA.Cn[14].n49 VGND 0.01568f
C6161 XA.Cn[14].n50 VGND 0.09061f
C6162 XA.Cn[14].n51 VGND 0.54091f
C6163 XA.Cn[14].n52 VGND 0.03454f
C6164 XA.Cn[14].t4 VGND 0.01419f
C6165 XA.Cn[14].t5 VGND 0.01419f
C6166 XA.Cn[14].n53 VGND 0.03067f
C6167 XA.Cn[14].t7 VGND 0.01419f
C6168 XA.Cn[14].t6 VGND 0.01419f
C6169 XA.Cn[14].n54 VGND 0.04667f
C6170 XA.Cn[14].n55 VGND 0.12968f
C6171 XA.Cn[14].n56 VGND 0.02039f
C6172 XA.Cn[14].t1 VGND 0.01419f
C6173 XA.Cn[14].t0 VGND 0.01419f
C6174 XA.Cn[14].n57 VGND 0.03155f
C6175 XA.Cn[14].t3 VGND 0.01419f
C6176 XA.Cn[14].t2 VGND 0.01419f
C6177 XA.Cn[14].n58 VGND 0.04309f
C6178 XA.Cn[14].n59 VGND 0.14042f
C6179 XThR.Tn[10].t10 VGND 0.01941f
C6180 XThR.Tn[10].t8 VGND 0.01941f
C6181 XThR.Tn[10].n0 VGND 0.05892f
C6182 XThR.Tn[10].t11 VGND 0.01941f
C6183 XThR.Tn[10].t9 VGND 0.01941f
C6184 XThR.Tn[10].n1 VGND 0.04314f
C6185 XThR.Tn[10].n2 VGND 0.19615f
C6186 XThR.Tn[10].t2 VGND 0.01261f
C6187 XThR.Tn[10].t7 VGND 0.01261f
C6188 XThR.Tn[10].n3 VGND 0.03146f
C6189 XThR.Tn[10].t1 VGND 0.01261f
C6190 XThR.Tn[10].t6 VGND 0.01261f
C6191 XThR.Tn[10].n4 VGND 0.02523f
C6192 XThR.Tn[10].n5 VGND 0.05817f
C6193 XThR.Tn[10].t54 VGND 0.01517f
C6194 XThR.Tn[10].t47 VGND 0.01661f
C6195 XThR.Tn[10].n6 VGND 0.04056f
C6196 XThR.Tn[10].n7 VGND 0.07791f
C6197 XThR.Tn[10].t13 VGND 0.01517f
C6198 XThR.Tn[10].t63 VGND 0.01661f
C6199 XThR.Tn[10].n8 VGND 0.04056f
C6200 XThR.Tn[10].t50 VGND 0.01512f
C6201 XThR.Tn[10].t60 VGND 0.01655f
C6202 XThR.Tn[10].n9 VGND 0.0422f
C6203 XThR.Tn[10].n10 VGND 0.02964f
C6204 XThR.Tn[10].n12 VGND 0.09513f
C6205 XThR.Tn[10].t48 VGND 0.01517f
C6206 XThR.Tn[10].t41 VGND 0.01661f
C6207 XThR.Tn[10].n13 VGND 0.04056f
C6208 XThR.Tn[10].t23 VGND 0.01512f
C6209 XThR.Tn[10].t36 VGND 0.01655f
C6210 XThR.Tn[10].n14 VGND 0.0422f
C6211 XThR.Tn[10].n15 VGND 0.02964f
C6212 XThR.Tn[10].n17 VGND 0.09513f
C6213 XThR.Tn[10].t65 VGND 0.01517f
C6214 XThR.Tn[10].t58 VGND 0.01661f
C6215 XThR.Tn[10].n18 VGND 0.04056f
C6216 XThR.Tn[10].t40 VGND 0.01512f
C6217 XThR.Tn[10].t55 VGND 0.01655f
C6218 XThR.Tn[10].n19 VGND 0.0422f
C6219 XThR.Tn[10].n20 VGND 0.02964f
C6220 XThR.Tn[10].n22 VGND 0.09513f
C6221 XThR.Tn[10].t30 VGND 0.01517f
C6222 XThR.Tn[10].t26 VGND 0.01661f
C6223 XThR.Tn[10].n23 VGND 0.04056f
C6224 XThR.Tn[10].t70 VGND 0.01512f
C6225 XThR.Tn[10].t21 VGND 0.01655f
C6226 XThR.Tn[10].n24 VGND 0.0422f
C6227 XThR.Tn[10].n25 VGND 0.02964f
C6228 XThR.Tn[10].n27 VGND 0.09513f
C6229 XThR.Tn[10].t67 VGND 0.01517f
C6230 XThR.Tn[10].t59 VGND 0.01661f
C6231 XThR.Tn[10].n28 VGND 0.04056f
C6232 XThR.Tn[10].t42 VGND 0.01512f
C6233 XThR.Tn[10].t56 VGND 0.01655f
C6234 XThR.Tn[10].n29 VGND 0.0422f
C6235 XThR.Tn[10].n30 VGND 0.02964f
C6236 XThR.Tn[10].n32 VGND 0.09513f
C6237 XThR.Tn[10].t44 VGND 0.01517f
C6238 XThR.Tn[10].t15 VGND 0.01661f
C6239 XThR.Tn[10].n33 VGND 0.04056f
C6240 XThR.Tn[10].t18 VGND 0.01512f
C6241 XThR.Tn[10].t12 VGND 0.01655f
C6242 XThR.Tn[10].n34 VGND 0.0422f
C6243 XThR.Tn[10].n35 VGND 0.02964f
C6244 XThR.Tn[10].n37 VGND 0.09513f
C6245 XThR.Tn[10].t14 VGND 0.01517f
C6246 XThR.Tn[10].t69 VGND 0.01661f
C6247 XThR.Tn[10].n38 VGND 0.04056f
C6248 XThR.Tn[10].t51 VGND 0.01512f
C6249 XThR.Tn[10].t66 VGND 0.01655f
C6250 XThR.Tn[10].n39 VGND 0.0422f
C6251 XThR.Tn[10].n40 VGND 0.02964f
C6252 XThR.Tn[10].n42 VGND 0.09513f
C6253 XThR.Tn[10].t17 VGND 0.01517f
C6254 XThR.Tn[10].t24 VGND 0.01661f
C6255 XThR.Tn[10].n43 VGND 0.04056f
C6256 XThR.Tn[10].t53 VGND 0.01512f
C6257 XThR.Tn[10].t20 VGND 0.01655f
C6258 XThR.Tn[10].n44 VGND 0.0422f
C6259 XThR.Tn[10].n45 VGND 0.02964f
C6260 XThR.Tn[10].n47 VGND 0.09513f
C6261 XThR.Tn[10].t33 VGND 0.01517f
C6262 XThR.Tn[10].t43 VGND 0.01661f
C6263 XThR.Tn[10].n48 VGND 0.04056f
C6264 XThR.Tn[10].t73 VGND 0.01512f
C6265 XThR.Tn[10].t38 VGND 0.01655f
C6266 XThR.Tn[10].n49 VGND 0.0422f
C6267 XThR.Tn[10].n50 VGND 0.02964f
C6268 XThR.Tn[10].n52 VGND 0.09513f
C6269 XThR.Tn[10].t28 VGND 0.01517f
C6270 XThR.Tn[10].t61 VGND 0.01661f
C6271 XThR.Tn[10].n53 VGND 0.04056f
C6272 XThR.Tn[10].t62 VGND 0.01512f
C6273 XThR.Tn[10].t57 VGND 0.01655f
C6274 XThR.Tn[10].n54 VGND 0.0422f
C6275 XThR.Tn[10].n55 VGND 0.02964f
C6276 XThR.Tn[10].n57 VGND 0.09513f
C6277 XThR.Tn[10].t46 VGND 0.01517f
C6278 XThR.Tn[10].t35 VGND 0.01661f
C6279 XThR.Tn[10].n58 VGND 0.04056f
C6280 XThR.Tn[10].t19 VGND 0.01512f
C6281 XThR.Tn[10].t32 VGND 0.01655f
C6282 XThR.Tn[10].n59 VGND 0.0422f
C6283 XThR.Tn[10].n60 VGND 0.02964f
C6284 XThR.Tn[10].n62 VGND 0.09513f
C6285 XThR.Tn[10].t16 VGND 0.01517f
C6286 XThR.Tn[10].t72 VGND 0.01661f
C6287 XThR.Tn[10].n63 VGND 0.04056f
C6288 XThR.Tn[10].t52 VGND 0.01512f
C6289 XThR.Tn[10].t68 VGND 0.01655f
C6290 XThR.Tn[10].n64 VGND 0.0422f
C6291 XThR.Tn[10].n65 VGND 0.02964f
C6292 XThR.Tn[10].n67 VGND 0.09513f
C6293 XThR.Tn[10].t31 VGND 0.01517f
C6294 XThR.Tn[10].t27 VGND 0.01661f
C6295 XThR.Tn[10].n68 VGND 0.04056f
C6296 XThR.Tn[10].t71 VGND 0.01512f
C6297 XThR.Tn[10].t22 VGND 0.01655f
C6298 XThR.Tn[10].n69 VGND 0.0422f
C6299 XThR.Tn[10].n70 VGND 0.02964f
C6300 XThR.Tn[10].n72 VGND 0.09513f
C6301 XThR.Tn[10].t49 VGND 0.01517f
C6302 XThR.Tn[10].t45 VGND 0.01661f
C6303 XThR.Tn[10].n73 VGND 0.04056f
C6304 XThR.Tn[10].t25 VGND 0.01512f
C6305 XThR.Tn[10].t39 VGND 0.01655f
C6306 XThR.Tn[10].n74 VGND 0.0422f
C6307 XThR.Tn[10].n75 VGND 0.02964f
C6308 XThR.Tn[10].n77 VGND 0.09513f
C6309 XThR.Tn[10].t29 VGND 0.01517f
C6310 XThR.Tn[10].t37 VGND 0.01661f
C6311 XThR.Tn[10].n78 VGND 0.04056f
C6312 XThR.Tn[10].t64 VGND 0.01512f
C6313 XThR.Tn[10].t34 VGND 0.01655f
C6314 XThR.Tn[10].n79 VGND 0.0422f
C6315 XThR.Tn[10].n80 VGND 0.02964f
C6316 XThR.Tn[10].n82 VGND 0.09513f
C6317 XThR.Tn[10].n83 VGND 0.08645f
C6318 XThR.Tn[10].n84 VGND 0.26614f
C6319 XThR.Tn[10].t0 VGND 0.01941f
C6320 XThR.Tn[10].t5 VGND 0.01941f
C6321 XThR.Tn[10].n85 VGND 0.04193f
C6322 XThR.Tn[10].t4 VGND 0.01941f
C6323 XThR.Tn[10].t3 VGND 0.01941f
C6324 XThR.Tn[10].n86 VGND 0.06382f
C6325 XThR.Tn[10].n87 VGND 0.1772f
C6326 XA.Cn[3].t5 VGND 0.01185f
C6327 XA.Cn[3].t4 VGND 0.01185f
C6328 XA.Cn[3].n0 VGND 0.02391f
C6329 XA.Cn[3].t7 VGND 0.01185f
C6330 XA.Cn[3].t6 VGND 0.01185f
C6331 XA.Cn[3].n1 VGND 0.02797f
C6332 XA.Cn[3].n2 VGND 0.08391f
C6333 XA.Cn[3].n3 VGND 0.01753f
C6334 XA.Cn[3].n4 VGND 0.01753f
C6335 XA.Cn[3].n5 VGND 0.01753f
C6336 XA.Cn[3].n6 VGND 0.02921f
C6337 XA.Cn[3].n7 VGND 0.0835f
C6338 XA.Cn[3].n8 VGND 0.05162f
C6339 XA.Cn[3].n9 VGND 0.05825f
C6340 XA.Cn[3].t42 VGND 0.01025f
C6341 XA.Cn[3].n10 VGND 0.0229f
C6342 XA.Cn[3].n11 VGND 0.01309f
C6343 XA.Cn[3].n12 VGND 0.01592f
C6344 XA.Cn[3].t27 VGND 0.01025f
C6345 XA.Cn[3].n13 VGND 0.0229f
C6346 XA.Cn[3].n14 VGND 0.01309f
C6347 XA.Cn[3].n15 VGND 0.07562f
C6348 XA.Cn[3].t29 VGND 0.01025f
C6349 XA.Cn[3].n16 VGND 0.0229f
C6350 XA.Cn[3].n17 VGND 0.01309f
C6351 XA.Cn[3].n18 VGND 0.07562f
C6352 XA.Cn[3].t31 VGND 0.01025f
C6353 XA.Cn[3].n19 VGND 0.0229f
C6354 XA.Cn[3].n20 VGND 0.01309f
C6355 XA.Cn[3].n21 VGND 0.07562f
C6356 XA.Cn[3].t20 VGND 0.01025f
C6357 XA.Cn[3].n22 VGND 0.0229f
C6358 XA.Cn[3].n23 VGND 0.01309f
C6359 XA.Cn[3].n24 VGND 0.07562f
C6360 XA.Cn[3].t21 VGND 0.01025f
C6361 XA.Cn[3].n25 VGND 0.0229f
C6362 XA.Cn[3].n26 VGND 0.01309f
C6363 XA.Cn[3].n27 VGND 0.07562f
C6364 XA.Cn[3].t34 VGND 0.01025f
C6365 XA.Cn[3].n28 VGND 0.0229f
C6366 XA.Cn[3].n29 VGND 0.01309f
C6367 XA.Cn[3].n30 VGND 0.07562f
C6368 XA.Cn[3].t43 VGND 0.01025f
C6369 XA.Cn[3].n31 VGND 0.0229f
C6370 XA.Cn[3].n32 VGND 0.01309f
C6371 XA.Cn[3].n33 VGND 0.07562f
C6372 XA.Cn[3].t13 VGND 0.01025f
C6373 XA.Cn[3].n34 VGND 0.0229f
C6374 XA.Cn[3].n35 VGND 0.01309f
C6375 XA.Cn[3].n36 VGND 0.07562f
C6376 XA.Cn[3].t32 VGND 0.01025f
C6377 XA.Cn[3].n37 VGND 0.0229f
C6378 XA.Cn[3].n38 VGND 0.01309f
C6379 XA.Cn[3].n39 VGND 0.07562f
C6380 XA.Cn[3].t33 VGND 0.01025f
C6381 XA.Cn[3].n40 VGND 0.0229f
C6382 XA.Cn[3].n41 VGND 0.01309f
C6383 XA.Cn[3].n42 VGND 0.07562f
C6384 XA.Cn[3].t14 VGND 0.01025f
C6385 XA.Cn[3].n43 VGND 0.0229f
C6386 XA.Cn[3].n44 VGND 0.01309f
C6387 XA.Cn[3].n45 VGND 0.07562f
C6388 XA.Cn[3].t22 VGND 0.01025f
C6389 XA.Cn[3].n46 VGND 0.0229f
C6390 XA.Cn[3].n47 VGND 0.01309f
C6391 XA.Cn[3].n48 VGND 0.07562f
C6392 XA.Cn[3].t25 VGND 0.01025f
C6393 XA.Cn[3].n49 VGND 0.0229f
C6394 XA.Cn[3].n50 VGND 0.01309f
C6395 XA.Cn[3].n51 VGND 0.07562f
C6396 XA.Cn[3].t38 VGND 0.01025f
C6397 XA.Cn[3].n52 VGND 0.0229f
C6398 XA.Cn[3].n53 VGND 0.01309f
C6399 XA.Cn[3].n54 VGND 0.07562f
C6400 XA.Cn[3].t16 VGND 0.01025f
C6401 XA.Cn[3].n55 VGND 0.0229f
C6402 XA.Cn[3].n56 VGND 0.01309f
C6403 XA.Cn[3].n57 VGND 0.07562f
C6404 XA.Cn[3].n58 VGND 0.03994f
C6405 XA.Cn[1].t3 VGND 0.0116f
C6406 XA.Cn[1].t2 VGND 0.0116f
C6407 XA.Cn[1].n0 VGND 0.02342f
C6408 XA.Cn[1].t1 VGND 0.0116f
C6409 XA.Cn[1].t0 VGND 0.0116f
C6410 XA.Cn[1].n1 VGND 0.02741f
C6411 XA.Cn[1].n2 VGND 0.08221f
C6412 XA.Cn[1].n3 VGND 0.02862f
C6413 XA.Cn[1].n4 VGND 0.01718f
C6414 XA.Cn[1].n5 VGND 0.0818f
C6415 XA.Cn[1].n6 VGND 0.01718f
C6416 XA.Cn[1].n7 VGND 0.05057f
C6417 XA.Cn[1].n8 VGND 0.01718f
C6418 XA.Cn[1].n9 VGND 0.05707f
C6419 XA.Cn[1].t29 VGND 0.01005f
C6420 XA.Cn[1].n10 VGND 0.02244f
C6421 XA.Cn[1].n11 VGND 0.01282f
C6422 XA.Cn[1].n12 VGND 0.01559f
C6423 XA.Cn[1].t14 VGND 0.01005f
C6424 XA.Cn[1].n13 VGND 0.02244f
C6425 XA.Cn[1].n14 VGND 0.01282f
C6426 XA.Cn[1].n15 VGND 0.07408f
C6427 XA.Cn[1].t16 VGND 0.01005f
C6428 XA.Cn[1].n16 VGND 0.02244f
C6429 XA.Cn[1].n17 VGND 0.01282f
C6430 XA.Cn[1].n18 VGND 0.07408f
C6431 XA.Cn[1].t18 VGND 0.01005f
C6432 XA.Cn[1].n19 VGND 0.02244f
C6433 XA.Cn[1].n20 VGND 0.01282f
C6434 XA.Cn[1].n21 VGND 0.07408f
C6435 XA.Cn[1].t39 VGND 0.01005f
C6436 XA.Cn[1].n22 VGND 0.02244f
C6437 XA.Cn[1].n23 VGND 0.01282f
C6438 XA.Cn[1].n24 VGND 0.07408f
C6439 XA.Cn[1].t40 VGND 0.01005f
C6440 XA.Cn[1].n25 VGND 0.02244f
C6441 XA.Cn[1].n26 VGND 0.01282f
C6442 XA.Cn[1].n27 VGND 0.07408f
C6443 XA.Cn[1].t21 VGND 0.01005f
C6444 XA.Cn[1].n28 VGND 0.02244f
C6445 XA.Cn[1].n29 VGND 0.01282f
C6446 XA.Cn[1].n30 VGND 0.07408f
C6447 XA.Cn[1].t30 VGND 0.01005f
C6448 XA.Cn[1].n31 VGND 0.02244f
C6449 XA.Cn[1].n32 VGND 0.01282f
C6450 XA.Cn[1].n33 VGND 0.07408f
C6451 XA.Cn[1].t32 VGND 0.01005f
C6452 XA.Cn[1].n34 VGND 0.02244f
C6453 XA.Cn[1].n35 VGND 0.01282f
C6454 XA.Cn[1].n36 VGND 0.07408f
C6455 XA.Cn[1].t19 VGND 0.01005f
C6456 XA.Cn[1].n37 VGND 0.02244f
C6457 XA.Cn[1].n38 VGND 0.01282f
C6458 XA.Cn[1].n39 VGND 0.07408f
C6459 XA.Cn[1].t20 VGND 0.01005f
C6460 XA.Cn[1].n40 VGND 0.02244f
C6461 XA.Cn[1].n41 VGND 0.01282f
C6462 XA.Cn[1].n42 VGND 0.07408f
C6463 XA.Cn[1].t33 VGND 0.01005f
C6464 XA.Cn[1].n43 VGND 0.02244f
C6465 XA.Cn[1].n44 VGND 0.01282f
C6466 XA.Cn[1].n45 VGND 0.07408f
C6467 XA.Cn[1].t41 VGND 0.01005f
C6468 XA.Cn[1].n46 VGND 0.02244f
C6469 XA.Cn[1].n47 VGND 0.01282f
C6470 XA.Cn[1].n48 VGND 0.07408f
C6471 XA.Cn[1].t12 VGND 0.01005f
C6472 XA.Cn[1].n49 VGND 0.02244f
C6473 XA.Cn[1].n50 VGND 0.01282f
C6474 XA.Cn[1].n51 VGND 0.07408f
C6475 XA.Cn[1].t25 VGND 0.01005f
C6476 XA.Cn[1].n52 VGND 0.02244f
C6477 XA.Cn[1].n53 VGND 0.01282f
C6478 XA.Cn[1].n54 VGND 0.07408f
C6479 XA.Cn[1].t35 VGND 0.01005f
C6480 XA.Cn[1].n55 VGND 0.02244f
C6481 XA.Cn[1].n56 VGND 0.01282f
C6482 XA.Cn[1].n57 VGND 0.07408f
C6483 XA.Cn[1].n58 VGND 0.27353f
C6484 XA.Cn[1].n59 VGND 0.0276f
C6485 Vbias.t260 VGND 0.17882f
C6486 Vbias.n0 VGND 0.19466f
C6487 Vbias.t79 VGND 0.17882f
C6488 Vbias.n1 VGND 0.19501f
C6489 Vbias.n2 VGND 0.12932f
C6490 Vbias.t174 VGND 0.17882f
C6491 Vbias.n3 VGND 0.19501f
C6492 Vbias.n4 VGND 0.12932f
C6493 Vbias.t182 VGND 0.17882f
C6494 Vbias.n5 VGND 0.19501f
C6495 Vbias.n6 VGND 0.12932f
C6496 Vbias.t15 VGND 0.17882f
C6497 Vbias.n7 VGND 0.19501f
C6498 Vbias.n8 VGND 0.12932f
C6499 Vbias.t101 VGND 0.17882f
C6500 Vbias.n9 VGND 0.19501f
C6501 Vbias.n10 VGND 0.12932f
C6502 Vbias.t184 VGND 0.17882f
C6503 Vbias.n11 VGND 0.19501f
C6504 Vbias.n12 VGND 0.12932f
C6505 Vbias.t19 VGND 0.17882f
C6506 Vbias.n13 VGND 0.19501f
C6507 Vbias.n14 VGND 0.12932f
C6508 Vbias.t39 VGND 0.17882f
C6509 Vbias.n15 VGND 0.19501f
C6510 Vbias.n16 VGND 0.12932f
C6511 Vbias.t111 VGND 0.17882f
C6512 Vbias.n17 VGND 0.19501f
C6513 Vbias.n18 VGND 0.12932f
C6514 Vbias.t202 VGND 0.17882f
C6515 Vbias.n19 VGND 0.19501f
C6516 Vbias.n20 VGND 0.12932f
C6517 Vbias.t223 VGND 0.17882f
C6518 Vbias.n21 VGND 0.19501f
C6519 Vbias.n22 VGND 0.12932f
C6520 Vbias.t114 VGND 0.17882f
C6521 Vbias.n23 VGND 0.19501f
C6522 Vbias.n24 VGND 0.12932f
C6523 Vbias.t142 VGND 0.17882f
C6524 Vbias.n25 VGND 0.19501f
C6525 Vbias.n26 VGND 0.12932f
C6526 Vbias.t151 VGND 0.17882f
C6527 Vbias.n27 VGND 0.19501f
C6528 Vbias.n28 VGND 0.12932f
C6529 Vbias.t61 VGND 0.17882f
C6530 Vbias.n29 VGND 0.19501f
C6531 Vbias.n30 VGND 0.12932f
C6532 Vbias.n31 VGND 0.54269f
C6533 Vbias.t140 VGND 0.17882f
C6534 Vbias.n32 VGND 0.19466f
C6535 Vbias.t216 VGND 0.17882f
C6536 Vbias.n33 VGND 0.19501f
C6537 Vbias.n34 VGND 0.12932f
C6538 Vbias.t59 VGND 0.17882f
C6539 Vbias.n35 VGND 0.19501f
C6540 Vbias.n36 VGND 0.12932f
C6541 Vbias.t67 VGND 0.17882f
C6542 Vbias.n37 VGND 0.19501f
C6543 Vbias.n38 VGND 0.12932f
C6544 Vbias.t152 VGND 0.17882f
C6545 Vbias.n39 VGND 0.19501f
C6546 Vbias.n40 VGND 0.12932f
C6547 Vbias.t245 VGND 0.17882f
C6548 Vbias.n41 VGND 0.19501f
C6549 Vbias.n42 VGND 0.12932f
C6550 Vbias.t72 VGND 0.17882f
C6551 Vbias.n43 VGND 0.19501f
C6552 Vbias.n44 VGND 0.12932f
C6553 Vbias.t158 VGND 0.17882f
C6554 Vbias.n45 VGND 0.19501f
C6555 Vbias.n46 VGND 0.12932f
C6556 Vbias.t178 VGND 0.17882f
C6557 Vbias.n47 VGND 0.19501f
C6558 Vbias.n48 VGND 0.12932f
C6559 Vbias.t254 VGND 0.17882f
C6560 Vbias.n49 VGND 0.19501f
C6561 Vbias.n50 VGND 0.12932f
C6562 Vbias.t84 VGND 0.17882f
C6563 Vbias.n51 VGND 0.19501f
C6564 Vbias.n52 VGND 0.12932f
C6565 Vbias.t106 VGND 0.17882f
C6566 Vbias.n53 VGND 0.19501f
C6567 Vbias.n54 VGND 0.12932f
C6568 Vbias.t259 VGND 0.17882f
C6569 Vbias.n55 VGND 0.19501f
C6570 Vbias.n56 VGND 0.12932f
C6571 Vbias.t26 VGND 0.17882f
C6572 Vbias.n57 VGND 0.19501f
C6573 Vbias.n58 VGND 0.12932f
C6574 Vbias.t35 VGND 0.17882f
C6575 Vbias.n59 VGND 0.19501f
C6576 Vbias.n60 VGND 0.12932f
C6577 Vbias.t194 VGND 0.17882f
C6578 Vbias.n61 VGND 0.19501f
C6579 Vbias.n62 VGND 0.12932f
C6580 Vbias.n63 VGND 0.55831f
C6581 Vbias.t215 VGND 0.17882f
C6582 Vbias.n64 VGND 0.19466f
C6583 Vbias.t31 VGND 0.17882f
C6584 Vbias.n65 VGND 0.19501f
C6585 Vbias.n66 VGND 0.12932f
C6586 Vbias.t132 VGND 0.17882f
C6587 Vbias.n67 VGND 0.19501f
C6588 Vbias.n68 VGND 0.12932f
C6589 Vbias.t139 VGND 0.17882f
C6590 Vbias.n69 VGND 0.19501f
C6591 Vbias.n70 VGND 0.12932f
C6592 Vbias.t224 VGND 0.17882f
C6593 Vbias.n71 VGND 0.19501f
C6594 Vbias.n72 VGND 0.12932f
C6595 Vbias.t58 VGND 0.17882f
C6596 Vbias.n73 VGND 0.19501f
C6597 Vbias.n74 VGND 0.12932f
C6598 Vbias.t145 VGND 0.17882f
C6599 Vbias.n75 VGND 0.19501f
C6600 Vbias.n76 VGND 0.12932f
C6601 Vbias.t230 VGND 0.17882f
C6602 Vbias.n77 VGND 0.19501f
C6603 Vbias.n78 VGND 0.12932f
C6604 Vbias.t253 VGND 0.17882f
C6605 Vbias.n79 VGND 0.19501f
C6606 Vbias.n80 VGND 0.12932f
C6607 Vbias.t71 VGND 0.17882f
C6608 Vbias.n81 VGND 0.19501f
C6609 Vbias.n82 VGND 0.12932f
C6610 Vbias.t157 VGND 0.17882f
C6611 Vbias.n83 VGND 0.19501f
C6612 Vbias.n84 VGND 0.12932f
C6613 Vbias.t177 VGND 0.17882f
C6614 Vbias.n85 VGND 0.19501f
C6615 Vbias.n86 VGND 0.12932f
C6616 Vbias.t77 VGND 0.17882f
C6617 Vbias.n87 VGND 0.19501f
C6618 Vbias.n88 VGND 0.12932f
C6619 Vbias.t97 VGND 0.17882f
C6620 Vbias.n89 VGND 0.19501f
C6621 Vbias.n90 VGND 0.12932f
C6622 Vbias.t104 VGND 0.17882f
C6623 Vbias.n91 VGND 0.19501f
C6624 Vbias.n92 VGND 0.12932f
C6625 Vbias.t13 VGND 0.17882f
C6626 Vbias.n93 VGND 0.19501f
C6627 Vbias.n94 VGND 0.12932f
C6628 Vbias.n95 VGND 0.55831f
C6629 Vbias.t30 VGND 0.17882f
C6630 Vbias.n96 VGND 0.19466f
C6631 Vbias.t100 VGND 0.17882f
C6632 Vbias.n97 VGND 0.19501f
C6633 Vbias.n98 VGND 0.12932f
C6634 Vbias.t203 VGND 0.17882f
C6635 Vbias.n99 VGND 0.19501f
C6636 Vbias.n100 VGND 0.12932f
C6637 Vbias.t214 VGND 0.17882f
C6638 Vbias.n101 VGND 0.19501f
C6639 Vbias.n102 VGND 0.12932f
C6640 Vbias.t38 VGND 0.17882f
C6641 Vbias.n103 VGND 0.19501f
C6642 Vbias.n104 VGND 0.12932f
C6643 Vbias.t131 VGND 0.17882f
C6644 Vbias.n105 VGND 0.19501f
C6645 Vbias.n106 VGND 0.12932f
C6646 Vbias.t218 VGND 0.17882f
C6647 Vbias.n107 VGND 0.19501f
C6648 Vbias.n108 VGND 0.12932f
C6649 Vbias.t42 VGND 0.17882f
C6650 Vbias.n109 VGND 0.19501f
C6651 Vbias.n110 VGND 0.12932f
C6652 Vbias.t70 VGND 0.17882f
C6653 Vbias.n111 VGND 0.19501f
C6654 Vbias.n112 VGND 0.12932f
C6655 Vbias.t143 VGND 0.17882f
C6656 Vbias.n113 VGND 0.19501f
C6657 Vbias.n114 VGND 0.12932f
C6658 Vbias.t228 VGND 0.17882f
C6659 Vbias.n115 VGND 0.19501f
C6660 Vbias.n116 VGND 0.12932f
C6661 Vbias.t252 VGND 0.17882f
C6662 Vbias.n117 VGND 0.19501f
C6663 Vbias.n118 VGND 0.12932f
C6664 Vbias.t148 VGND 0.17882f
C6665 Vbias.n119 VGND 0.19501f
C6666 Vbias.n120 VGND 0.12932f
C6667 Vbias.t170 VGND 0.17882f
C6668 Vbias.n121 VGND 0.19501f
C6669 Vbias.n122 VGND 0.12932f
C6670 Vbias.t175 VGND 0.17882f
C6671 Vbias.n123 VGND 0.19501f
C6672 Vbias.n124 VGND 0.12932f
C6673 Vbias.t86 VGND 0.17882f
C6674 Vbias.n125 VGND 0.19501f
C6675 Vbias.n126 VGND 0.12932f
C6676 Vbias.n127 VGND 0.55831f
C6677 Vbias.t186 VGND 0.17882f
C6678 Vbias.n128 VGND 0.19466f
C6679 Vbias.t6 VGND 0.17882f
C6680 Vbias.n129 VGND 0.19501f
C6681 Vbias.n130 VGND 0.12932f
C6682 Vbias.t103 VGND 0.17882f
C6683 Vbias.n131 VGND 0.19501f
C6684 Vbias.n132 VGND 0.12932f
C6685 Vbias.t115 VGND 0.17882f
C6686 Vbias.n133 VGND 0.19501f
C6687 Vbias.n134 VGND 0.12932f
C6688 Vbias.t206 VGND 0.17882f
C6689 Vbias.n135 VGND 0.19501f
C6690 Vbias.n136 VGND 0.12932f
C6691 Vbias.t34 VGND 0.17882f
C6692 Vbias.n137 VGND 0.19501f
C6693 Vbias.n138 VGND 0.12932f
C6694 Vbias.t116 VGND 0.17882f
C6695 Vbias.n139 VGND 0.19501f
C6696 Vbias.n140 VGND 0.12932f
C6697 Vbias.t209 VGND 0.17882f
C6698 Vbias.n141 VGND 0.19501f
C6699 Vbias.n142 VGND 0.12932f
C6700 Vbias.t231 VGND 0.17882f
C6701 Vbias.n143 VGND 0.19501f
C6702 Vbias.n144 VGND 0.12932f
C6703 Vbias.t43 VGND 0.17882f
C6704 Vbias.n145 VGND 0.19501f
C6705 Vbias.n146 VGND 0.12932f
C6706 Vbias.t134 VGND 0.17882f
C6707 Vbias.n147 VGND 0.19501f
C6708 Vbias.n148 VGND 0.12932f
C6709 Vbias.t159 VGND 0.17882f
C6710 Vbias.n149 VGND 0.19501f
C6711 Vbias.n150 VGND 0.12932f
C6712 Vbias.t47 VGND 0.17882f
C6713 Vbias.n151 VGND 0.19501f
C6714 Vbias.n152 VGND 0.12932f
C6715 Vbias.t78 VGND 0.17882f
C6716 Vbias.n153 VGND 0.19501f
C6717 Vbias.n154 VGND 0.12932f
C6718 Vbias.t85 VGND 0.17882f
C6719 Vbias.n155 VGND 0.19501f
C6720 Vbias.n156 VGND 0.12932f
C6721 Vbias.t249 VGND 0.17882f
C6722 Vbias.n157 VGND 0.19501f
C6723 Vbias.n158 VGND 0.12932f
C6724 Vbias.n159 VGND 0.55831f
C6725 Vbias.t55 VGND 0.17882f
C6726 Vbias.n160 VGND 0.19466f
C6727 Vbias.t128 VGND 0.17882f
C6728 Vbias.n161 VGND 0.19501f
C6729 Vbias.n162 VGND 0.12932f
C6730 Vbias.t226 VGND 0.17882f
C6731 Vbias.n163 VGND 0.19501f
C6732 Vbias.n164 VGND 0.12932f
C6733 Vbias.t241 VGND 0.17882f
C6734 Vbias.n165 VGND 0.19501f
C6735 Vbias.n166 VGND 0.12932f
C6736 Vbias.t66 VGND 0.17882f
C6737 Vbias.n167 VGND 0.19501f
C6738 Vbias.n168 VGND 0.12932f
C6739 Vbias.t155 VGND 0.17882f
C6740 Vbias.n169 VGND 0.19501f
C6741 Vbias.n170 VGND 0.12932f
C6742 Vbias.t244 VGND 0.17882f
C6743 Vbias.n171 VGND 0.19501f
C6744 Vbias.n172 VGND 0.12932f
C6745 Vbias.t74 VGND 0.17882f
C6746 Vbias.n173 VGND 0.19501f
C6747 Vbias.n174 VGND 0.12932f
C6748 Vbias.t94 VGND 0.17882f
C6749 Vbias.n175 VGND 0.19501f
C6750 Vbias.n176 VGND 0.12932f
C6751 Vbias.t167 VGND 0.17882f
C6752 Vbias.n177 VGND 0.19501f
C6753 Vbias.n178 VGND 0.12932f
C6754 Vbias.t256 VGND 0.17882f
C6755 Vbias.n179 VGND 0.19501f
C6756 Vbias.n180 VGND 0.12932f
C6757 Vbias.t22 VGND 0.17882f
C6758 Vbias.n181 VGND 0.19501f
C6759 Vbias.n182 VGND 0.12932f
C6760 Vbias.t172 VGND 0.17882f
C6761 Vbias.n183 VGND 0.19501f
C6762 Vbias.n184 VGND 0.12932f
C6763 Vbias.t191 VGND 0.17882f
C6764 Vbias.n185 VGND 0.19501f
C6765 Vbias.n186 VGND 0.12932f
C6766 Vbias.t207 VGND 0.17882f
C6767 Vbias.n187 VGND 0.19501f
C6768 Vbias.n188 VGND 0.12932f
C6769 Vbias.t109 VGND 0.17882f
C6770 Vbias.n189 VGND 0.19501f
C6771 Vbias.n190 VGND 0.12932f
C6772 Vbias.n191 VGND 0.55831f
C6773 Vbias.t189 VGND 0.17882f
C6774 Vbias.n192 VGND 0.19466f
C6775 Vbias.t10 VGND 0.17882f
C6776 Vbias.n193 VGND 0.19501f
C6777 Vbias.n194 VGND 0.12932f
C6778 Vbias.t108 VGND 0.17882f
C6779 Vbias.n195 VGND 0.19501f
C6780 Vbias.n196 VGND 0.12932f
C6781 Vbias.t117 VGND 0.17882f
C6782 Vbias.n197 VGND 0.19501f
C6783 Vbias.n198 VGND 0.12932f
C6784 Vbias.t208 VGND 0.17882f
C6785 Vbias.n199 VGND 0.19501f
C6786 Vbias.n200 VGND 0.12932f
C6787 Vbias.t36 VGND 0.17882f
C6788 Vbias.n201 VGND 0.19501f
C6789 Vbias.n202 VGND 0.12932f
C6790 Vbias.t120 VGND 0.17882f
C6791 Vbias.n203 VGND 0.19501f
C6792 Vbias.n204 VGND 0.12932f
C6793 Vbias.t212 VGND 0.17882f
C6794 Vbias.n205 VGND 0.19501f
C6795 Vbias.n206 VGND 0.12932f
C6796 Vbias.t234 VGND 0.17882f
C6797 Vbias.n207 VGND 0.19501f
C6798 Vbias.n208 VGND 0.12932f
C6799 Vbias.t46 VGND 0.17882f
C6800 Vbias.n209 VGND 0.19501f
C6801 Vbias.n210 VGND 0.12932f
C6802 Vbias.t136 VGND 0.17882f
C6803 Vbias.n211 VGND 0.19501f
C6804 Vbias.n212 VGND 0.12932f
C6805 Vbias.t162 VGND 0.17882f
C6806 Vbias.n213 VGND 0.19501f
C6807 Vbias.n214 VGND 0.12932f
C6808 Vbias.t51 VGND 0.17882f
C6809 Vbias.n215 VGND 0.19501f
C6810 Vbias.n216 VGND 0.12932f
C6811 Vbias.t80 VGND 0.17882f
C6812 Vbias.n217 VGND 0.19501f
C6813 Vbias.n218 VGND 0.12932f
C6814 Vbias.t89 VGND 0.17882f
C6815 Vbias.n219 VGND 0.19501f
C6816 Vbias.n220 VGND 0.12932f
C6817 Vbias.t250 VGND 0.17882f
C6818 Vbias.n221 VGND 0.19501f
C6819 Vbias.n222 VGND 0.12932f
C6820 Vbias.n223 VGND 0.55831f
C6821 Vbias.t9 VGND 0.17882f
C6822 Vbias.n224 VGND 0.19466f
C6823 Vbias.t83 VGND 0.17882f
C6824 Vbias.n225 VGND 0.19501f
C6825 Vbias.n226 VGND 0.12932f
C6826 Vbias.t180 VGND 0.17882f
C6827 Vbias.n227 VGND 0.19501f
C6828 Vbias.n228 VGND 0.12932f
C6829 Vbias.t188 VGND 0.17882f
C6830 Vbias.n229 VGND 0.19501f
C6831 Vbias.n230 VGND 0.12932f
C6832 Vbias.t23 VGND 0.17882f
C6833 Vbias.n231 VGND 0.19501f
C6834 Vbias.n232 VGND 0.12932f
C6835 Vbias.t107 VGND 0.17882f
C6836 Vbias.n233 VGND 0.19501f
C6837 Vbias.n234 VGND 0.12932f
C6838 Vbias.t192 VGND 0.17882f
C6839 Vbias.n235 VGND 0.19501f
C6840 Vbias.n236 VGND 0.12932f
C6841 Vbias.t28 VGND 0.17882f
C6842 Vbias.n237 VGND 0.19501f
C6843 Vbias.n238 VGND 0.12932f
C6844 Vbias.t45 VGND 0.17882f
C6845 Vbias.n239 VGND 0.19501f
C6846 Vbias.n240 VGND 0.12932f
C6847 Vbias.t119 VGND 0.17882f
C6848 Vbias.n241 VGND 0.19501f
C6849 Vbias.n242 VGND 0.12932f
C6850 Vbias.t211 VGND 0.17882f
C6851 Vbias.n243 VGND 0.19501f
C6852 Vbias.n244 VGND 0.12932f
C6853 Vbias.t233 VGND 0.17882f
C6854 Vbias.n245 VGND 0.19501f
C6855 Vbias.n246 VGND 0.12932f
C6856 Vbias.t123 VGND 0.17882f
C6857 Vbias.n247 VGND 0.19501f
C6858 Vbias.n248 VGND 0.12932f
C6859 Vbias.t149 VGND 0.17882f
C6860 Vbias.n249 VGND 0.19501f
C6861 Vbias.n250 VGND 0.12932f
C6862 Vbias.t161 VGND 0.17882f
C6863 Vbias.n251 VGND 0.19501f
C6864 Vbias.n252 VGND 0.12932f
C6865 Vbias.t64 VGND 0.17882f
C6866 Vbias.n253 VGND 0.19501f
C6867 Vbias.n254 VGND 0.12932f
C6868 Vbias.n255 VGND 0.55831f
C6869 Vbias.t82 VGND 0.17882f
C6870 Vbias.n256 VGND 0.19466f
C6871 Vbias.t154 VGND 0.17882f
C6872 Vbias.n257 VGND 0.19501f
C6873 Vbias.n258 VGND 0.12932f
C6874 Vbias.t257 VGND 0.17882f
C6875 Vbias.n259 VGND 0.19501f
C6876 Vbias.n260 VGND 0.12932f
C6877 Vbias.t8 VGND 0.17882f
C6878 Vbias.n261 VGND 0.19501f
C6879 Vbias.n262 VGND 0.12932f
C6880 Vbias.t93 VGND 0.17882f
C6881 Vbias.n263 VGND 0.19501f
C6882 Vbias.n264 VGND 0.12932f
C6883 Vbias.t179 VGND 0.17882f
C6884 Vbias.n265 VGND 0.19501f
C6885 Vbias.n266 VGND 0.12932f
C6886 Vbias.t11 VGND 0.17882f
C6887 Vbias.n267 VGND 0.19501f
C6888 Vbias.n268 VGND 0.12932f
C6889 Vbias.t98 VGND 0.17882f
C6890 Vbias.n269 VGND 0.19501f
C6891 Vbias.n270 VGND 0.12932f
C6892 Vbias.t118 VGND 0.17882f
C6893 Vbias.n271 VGND 0.19501f
C6894 Vbias.n272 VGND 0.12932f
C6895 Vbias.t190 VGND 0.17882f
C6896 Vbias.n273 VGND 0.19501f
C6897 Vbias.n274 VGND 0.12932f
C6898 Vbias.t27 VGND 0.17882f
C6899 Vbias.n275 VGND 0.19501f
C6900 Vbias.n276 VGND 0.12932f
C6901 Vbias.t44 VGND 0.17882f
C6902 Vbias.n277 VGND 0.19501f
C6903 Vbias.n278 VGND 0.12932f
C6904 Vbias.t197 VGND 0.17882f
C6905 Vbias.n279 VGND 0.19501f
C6906 Vbias.n280 VGND 0.12932f
C6907 Vbias.t220 VGND 0.17882f
C6908 Vbias.n281 VGND 0.19501f
C6909 Vbias.n282 VGND 0.12932f
C6910 Vbias.t232 VGND 0.17882f
C6911 Vbias.n283 VGND 0.19501f
C6912 Vbias.n284 VGND 0.12932f
C6913 Vbias.t137 VGND 0.17882f
C6914 Vbias.n285 VGND 0.19501f
C6915 Vbias.n286 VGND 0.12932f
C6916 Vbias.n287 VGND 0.55831f
C6917 Vbias.t49 VGND 0.17882f
C6918 Vbias.n288 VGND 0.19466f
C6919 Vbias.t122 VGND 0.17882f
C6920 Vbias.n289 VGND 0.19501f
C6921 Vbias.n290 VGND 0.12932f
C6922 Vbias.t222 VGND 0.17882f
C6923 Vbias.n291 VGND 0.19501f
C6924 Vbias.n292 VGND 0.12932f
C6925 Vbias.t235 VGND 0.17882f
C6926 Vbias.n293 VGND 0.19501f
C6927 Vbias.n294 VGND 0.12932f
C6928 Vbias.t63 VGND 0.17882f
C6929 Vbias.n295 VGND 0.19501f
C6930 Vbias.n296 VGND 0.12932f
C6931 Vbias.t150 VGND 0.17882f
C6932 Vbias.n297 VGND 0.19501f
C6933 Vbias.n298 VGND 0.12932f
C6934 Vbias.t237 VGND 0.17882f
C6935 Vbias.n299 VGND 0.19501f
C6936 Vbias.n300 VGND 0.12932f
C6937 Vbias.t68 VGND 0.17882f
C6938 Vbias.n301 VGND 0.19501f
C6939 Vbias.n302 VGND 0.12932f
C6940 Vbias.t91 VGND 0.17882f
C6941 Vbias.n303 VGND 0.19501f
C6942 Vbias.n304 VGND 0.12932f
C6943 Vbias.t164 VGND 0.17882f
C6944 Vbias.n305 VGND 0.19501f
C6945 Vbias.n306 VGND 0.12932f
C6946 Vbias.t251 VGND 0.17882f
C6947 Vbias.n307 VGND 0.19501f
C6948 Vbias.n308 VGND 0.12932f
C6949 Vbias.t21 VGND 0.17882f
C6950 Vbias.n309 VGND 0.19501f
C6951 Vbias.n310 VGND 0.12932f
C6952 Vbias.t168 VGND 0.17882f
C6953 Vbias.n311 VGND 0.19501f
C6954 Vbias.n312 VGND 0.12932f
C6955 Vbias.t187 VGND 0.17882f
C6956 Vbias.n313 VGND 0.19501f
C6957 Vbias.n314 VGND 0.12932f
C6958 Vbias.t204 VGND 0.17882f
C6959 Vbias.n315 VGND 0.19501f
C6960 Vbias.n316 VGND 0.12932f
C6961 Vbias.t105 VGND 0.17882f
C6962 Vbias.n317 VGND 0.19501f
C6963 Vbias.n318 VGND 0.12932f
C6964 Vbias.n319 VGND 0.55831f
C6965 Vbias.t121 VGND 0.17882f
C6966 Vbias.n320 VGND 0.19466f
C6967 Vbias.t195 VGND 0.17882f
C6968 Vbias.n321 VGND 0.19501f
C6969 Vbias.n322 VGND 0.12932f
C6970 Vbias.t37 VGND 0.17882f
C6971 Vbias.n323 VGND 0.19501f
C6972 Vbias.n324 VGND 0.12932f
C6973 Vbias.t48 VGND 0.17882f
C6974 Vbias.n325 VGND 0.19501f
C6975 Vbias.n326 VGND 0.12932f
C6976 Vbias.t135 VGND 0.17882f
C6977 Vbias.n327 VGND 0.19501f
C6978 Vbias.n328 VGND 0.12932f
C6979 Vbias.t221 VGND 0.17882f
C6980 Vbias.n329 VGND 0.19501f
C6981 Vbias.n330 VGND 0.12932f
C6982 Vbias.t50 VGND 0.17882f
C6983 Vbias.n331 VGND 0.19501f
C6984 Vbias.n332 VGND 0.12932f
C6985 Vbias.t138 VGND 0.17882f
C6986 Vbias.n333 VGND 0.19501f
C6987 Vbias.n334 VGND 0.12932f
C6988 Vbias.t163 VGND 0.17882f
C6989 Vbias.n335 VGND 0.19501f
C6990 Vbias.n336 VGND 0.12932f
C6991 Vbias.t236 VGND 0.17882f
C6992 Vbias.n337 VGND 0.19501f
C6993 Vbias.n338 VGND 0.12932f
C6994 Vbias.t65 VGND 0.17882f
C6995 Vbias.n339 VGND 0.19501f
C6996 Vbias.n340 VGND 0.12932f
C6997 Vbias.t90 VGND 0.17882f
C6998 Vbias.n341 VGND 0.19501f
C6999 Vbias.n342 VGND 0.12932f
C7000 Vbias.t243 VGND 0.17882f
C7001 Vbias.n343 VGND 0.19501f
C7002 Vbias.n344 VGND 0.12932f
C7003 Vbias.t7 VGND 0.17882f
C7004 Vbias.n345 VGND 0.19501f
C7005 Vbias.n346 VGND 0.12932f
C7006 Vbias.t20 VGND 0.17882f
C7007 Vbias.n347 VGND 0.19501f
C7008 Vbias.n348 VGND 0.12932f
C7009 Vbias.t176 VGND 0.17882f
C7010 Vbias.n349 VGND 0.19501f
C7011 Vbias.n350 VGND 0.12932f
C7012 Vbias.n351 VGND 0.55831f
C7013 Vbias.t198 VGND 0.17882f
C7014 Vbias.n352 VGND 0.19466f
C7015 Vbias.t17 VGND 0.17882f
C7016 Vbias.n353 VGND 0.19501f
C7017 Vbias.n354 VGND 0.12932f
C7018 Vbias.t113 VGND 0.17882f
C7019 Vbias.n355 VGND 0.19501f
C7020 Vbias.n356 VGND 0.12932f
C7021 Vbias.t124 VGND 0.17882f
C7022 Vbias.n357 VGND 0.19501f
C7023 Vbias.n358 VGND 0.12932f
C7024 Vbias.t213 VGND 0.17882f
C7025 Vbias.n359 VGND 0.19501f
C7026 Vbias.n360 VGND 0.12932f
C7027 Vbias.t40 VGND 0.17882f
C7028 Vbias.n361 VGND 0.19501f
C7029 Vbias.n362 VGND 0.12932f
C7030 Vbias.t127 VGND 0.17882f
C7031 Vbias.n363 VGND 0.19501f
C7032 Vbias.n364 VGND 0.12932f
C7033 Vbias.t219 VGND 0.17882f
C7034 Vbias.n365 VGND 0.19501f
C7035 Vbias.n366 VGND 0.12932f
C7036 Vbias.t240 VGND 0.17882f
C7037 Vbias.n367 VGND 0.19501f
C7038 Vbias.n368 VGND 0.12932f
C7039 Vbias.t54 VGND 0.17882f
C7040 Vbias.n369 VGND 0.19501f
C7041 Vbias.n370 VGND 0.12932f
C7042 Vbias.t144 VGND 0.17882f
C7043 Vbias.n371 VGND 0.19501f
C7044 Vbias.n372 VGND 0.12932f
C7045 Vbias.t166 VGND 0.17882f
C7046 Vbias.n373 VGND 0.19501f
C7047 Vbias.n374 VGND 0.12932f
C7048 Vbias.t62 VGND 0.17882f
C7049 Vbias.n375 VGND 0.19501f
C7050 Vbias.n376 VGND 0.12932f
C7051 Vbias.t81 VGND 0.17882f
C7052 Vbias.n377 VGND 0.19501f
C7053 Vbias.n378 VGND 0.12932f
C7054 Vbias.t92 VGND 0.17882f
C7055 Vbias.n379 VGND 0.19501f
C7056 Vbias.n380 VGND 0.12932f
C7057 Vbias.t255 VGND 0.17882f
C7058 Vbias.n381 VGND 0.19501f
C7059 Vbias.n382 VGND 0.12932f
C7060 Vbias.n383 VGND 0.55831f
C7061 Vbias.t16 VGND 0.17882f
C7062 Vbias.n384 VGND 0.19466f
C7063 Vbias.t88 VGND 0.17882f
C7064 Vbias.n385 VGND 0.19501f
C7065 Vbias.n386 VGND 0.12932f
C7066 Vbias.t185 VGND 0.17882f
C7067 Vbias.n387 VGND 0.19501f
C7068 Vbias.n388 VGND 0.12932f
C7069 Vbias.t196 VGND 0.17882f
C7070 Vbias.n389 VGND 0.19501f
C7071 Vbias.n390 VGND 0.12932f
C7072 Vbias.t29 VGND 0.17882f
C7073 Vbias.n391 VGND 0.19501f
C7074 Vbias.n392 VGND 0.12932f
C7075 Vbias.t112 VGND 0.17882f
C7076 Vbias.n393 VGND 0.19501f
C7077 Vbias.n394 VGND 0.12932f
C7078 Vbias.t200 VGND 0.17882f
C7079 Vbias.n395 VGND 0.19501f
C7080 Vbias.n396 VGND 0.12932f
C7081 Vbias.t33 VGND 0.17882f
C7082 Vbias.n397 VGND 0.19501f
C7083 Vbias.n398 VGND 0.12932f
C7084 Vbias.t53 VGND 0.17882f
C7085 Vbias.n399 VGND 0.19501f
C7086 Vbias.n400 VGND 0.12932f
C7087 Vbias.t126 VGND 0.17882f
C7088 Vbias.n401 VGND 0.19501f
C7089 Vbias.n402 VGND 0.12932f
C7090 Vbias.t217 VGND 0.17882f
C7091 Vbias.n403 VGND 0.19501f
C7092 Vbias.n404 VGND 0.12932f
C7093 Vbias.t239 VGND 0.17882f
C7094 Vbias.n405 VGND 0.19501f
C7095 Vbias.n406 VGND 0.12932f
C7096 Vbias.t133 VGND 0.17882f
C7097 Vbias.n407 VGND 0.19501f
C7098 Vbias.n408 VGND 0.12932f
C7099 Vbias.t153 VGND 0.17882f
C7100 Vbias.n409 VGND 0.19501f
C7101 Vbias.n410 VGND 0.12932f
C7102 Vbias.t165 VGND 0.17882f
C7103 Vbias.n411 VGND 0.19501f
C7104 Vbias.n412 VGND 0.12932f
C7105 Vbias.t73 VGND 0.17882f
C7106 Vbias.n413 VGND 0.19501f
C7107 Vbias.n414 VGND 0.12932f
C7108 Vbias.n415 VGND 0.55831f
C7109 Vbias.t87 VGND 0.17882f
C7110 Vbias.n416 VGND 0.19466f
C7111 Vbias.t160 VGND 0.17882f
C7112 Vbias.n417 VGND 0.19501f
C7113 Vbias.n418 VGND 0.12932f
C7114 Vbias.t261 VGND 0.17882f
C7115 Vbias.n419 VGND 0.19501f
C7116 Vbias.n420 VGND 0.12932f
C7117 Vbias.t14 VGND 0.17882f
C7118 Vbias.n421 VGND 0.19501f
C7119 Vbias.n422 VGND 0.12932f
C7120 Vbias.t99 VGND 0.17882f
C7121 Vbias.n423 VGND 0.19501f
C7122 Vbias.n424 VGND 0.12932f
C7123 Vbias.t183 VGND 0.17882f
C7124 Vbias.n425 VGND 0.19501f
C7125 Vbias.n426 VGND 0.12932f
C7126 Vbias.t18 VGND 0.17882f
C7127 Vbias.n427 VGND 0.19501f
C7128 Vbias.n428 VGND 0.12932f
C7129 Vbias.t102 VGND 0.17882f
C7130 Vbias.n429 VGND 0.19501f
C7131 Vbias.n430 VGND 0.12932f
C7132 Vbias.t125 VGND 0.17882f
C7133 Vbias.n431 VGND 0.19501f
C7134 Vbias.n432 VGND 0.12932f
C7135 Vbias.t199 VGND 0.17882f
C7136 Vbias.n433 VGND 0.19501f
C7137 Vbias.n434 VGND 0.12932f
C7138 Vbias.t32 VGND 0.17882f
C7139 Vbias.n435 VGND 0.19501f
C7140 Vbias.n436 VGND 0.12932f
C7141 Vbias.t52 VGND 0.17882f
C7142 Vbias.n437 VGND 0.19501f
C7143 Vbias.n438 VGND 0.12932f
C7144 Vbias.t205 VGND 0.17882f
C7145 Vbias.n439 VGND 0.19501f
C7146 Vbias.n440 VGND 0.12932f
C7147 Vbias.t225 VGND 0.17882f
C7148 Vbias.n441 VGND 0.19501f
C7149 Vbias.n442 VGND 0.12932f
C7150 Vbias.t238 VGND 0.17882f
C7151 Vbias.n443 VGND 0.19501f
C7152 Vbias.n444 VGND 0.12932f
C7153 Vbias.t146 VGND 0.17882f
C7154 Vbias.n445 VGND 0.19501f
C7155 Vbias.n446 VGND 0.12932f
C7156 Vbias.n447 VGND 0.55831f
C7157 Vbias.t57 VGND 0.17882f
C7158 Vbias.n448 VGND 0.19466f
C7159 Vbias.t130 VGND 0.17882f
C7160 Vbias.n449 VGND 0.19501f
C7161 Vbias.n450 VGND 0.12932f
C7162 Vbias.t229 VGND 0.17882f
C7163 Vbias.n451 VGND 0.19501f
C7164 Vbias.n452 VGND 0.12932f
C7165 Vbias.t242 VGND 0.17882f
C7166 Vbias.n453 VGND 0.19501f
C7167 Vbias.n454 VGND 0.12932f
C7168 Vbias.t69 VGND 0.17882f
C7169 Vbias.n455 VGND 0.19501f
C7170 Vbias.n456 VGND 0.12932f
C7171 Vbias.t156 VGND 0.17882f
C7172 Vbias.n457 VGND 0.19501f
C7173 Vbias.n458 VGND 0.12932f
C7174 Vbias.t247 VGND 0.17882f
C7175 Vbias.n459 VGND 0.19501f
C7176 Vbias.n460 VGND 0.12932f
C7177 Vbias.t76 VGND 0.17882f
C7178 Vbias.n461 VGND 0.19501f
C7179 Vbias.n462 VGND 0.12932f
C7180 Vbias.t96 VGND 0.17882f
C7181 Vbias.n463 VGND 0.19501f
C7182 Vbias.n464 VGND 0.12932f
C7183 Vbias.t171 VGND 0.17882f
C7184 Vbias.n465 VGND 0.19501f
C7185 Vbias.n466 VGND 0.12932f
C7186 Vbias.t258 VGND 0.17882f
C7187 Vbias.n467 VGND 0.19501f
C7188 Vbias.n468 VGND 0.12932f
C7189 Vbias.t25 VGND 0.17882f
C7190 Vbias.n469 VGND 0.19501f
C7191 Vbias.n470 VGND 0.12932f
C7192 Vbias.t173 VGND 0.17882f
C7193 Vbias.n471 VGND 0.19501f
C7194 Vbias.n472 VGND 0.12932f
C7195 Vbias.t193 VGND 0.17882f
C7196 Vbias.n473 VGND 0.19501f
C7197 Vbias.n474 VGND 0.12932f
C7198 Vbias.t210 VGND 0.17882f
C7199 Vbias.n475 VGND 0.19501f
C7200 Vbias.n476 VGND 0.12932f
C7201 Vbias.t110 VGND 0.17882f
C7202 Vbias.n477 VGND 0.19501f
C7203 Vbias.n478 VGND 0.12932f
C7204 Vbias.n479 VGND 0.55831f
C7205 Vbias.t129 VGND 0.17882f
C7206 Vbias.n480 VGND 0.19466f
C7207 Vbias.t201 VGND 0.17882f
C7208 Vbias.n481 VGND 0.19501f
C7209 Vbias.n482 VGND 0.12932f
C7210 Vbias.t41 VGND 0.17882f
C7211 Vbias.n483 VGND 0.19501f
C7212 Vbias.n484 VGND 0.12932f
C7213 Vbias.t56 VGND 0.17882f
C7214 Vbias.n485 VGND 0.19501f
C7215 Vbias.n486 VGND 0.12932f
C7216 Vbias.t141 VGND 0.17882f
C7217 Vbias.n487 VGND 0.19501f
C7218 Vbias.n488 VGND 0.12932f
C7219 Vbias.t227 VGND 0.17882f
C7220 Vbias.n489 VGND 0.19501f
C7221 Vbias.n490 VGND 0.12932f
C7222 Vbias.t60 VGND 0.17882f
C7223 Vbias.n491 VGND 0.19501f
C7224 Vbias.n492 VGND 0.12932f
C7225 Vbias.t147 VGND 0.17882f
C7226 Vbias.n493 VGND 0.19501f
C7227 Vbias.n494 VGND 0.12932f
C7228 Vbias.t169 VGND 0.17882f
C7229 Vbias.n495 VGND 0.19501f
C7230 Vbias.n496 VGND 0.12932f
C7231 Vbias.t246 VGND 0.17882f
C7232 Vbias.n497 VGND 0.19501f
C7233 Vbias.n498 VGND 0.12932f
C7234 Vbias.t75 VGND 0.17882f
C7235 Vbias.n499 VGND 0.19501f
C7236 Vbias.n500 VGND 0.12932f
C7237 Vbias.t95 VGND 0.17882f
C7238 Vbias.n501 VGND 0.19501f
C7239 Vbias.n502 VGND 0.12932f
C7240 Vbias.t248 VGND 0.17882f
C7241 Vbias.n503 VGND 0.19501f
C7242 Vbias.n504 VGND 0.12932f
C7243 Vbias.t12 VGND 0.17882f
C7244 Vbias.n505 VGND 0.19501f
C7245 Vbias.n506 VGND 0.12932f
C7246 Vbias.t24 VGND 0.17882f
C7247 Vbias.n507 VGND 0.19501f
C7248 Vbias.n508 VGND 0.12932f
C7249 Vbias.t181 VGND 0.17882f
C7250 Vbias.n509 VGND 0.19501f
C7251 Vbias.n510 VGND 0.12932f
C7252 Vbias.n511 VGND 0.64934f
C7253 Vbias.t0 VGND 0.03654f
C7254 Vbias.t2 VGND 0.03654f
C7255 Vbias.n512 VGND 0.24617f
C7256 Vbias.t5 VGND 0.03654f
C7257 Vbias.t1 VGND 0.03654f
C7258 Vbias.n513 VGND 0.24617f
C7259 Vbias.n514 VGND 0.74304f
C7260 Vbias.t4 VGND 0.17043f
C7261 Vbias.t3 VGND 0.67015f
C7262 Vbias.n515 VGND 1.2407f
C7263 Vbias.n516 VGND 0.47721f
C7264 Vbias.n517 VGND 1.11739f
C7265 XA.Cn[2].t9 VGND 0.01169f
C7266 XA.Cn[2].t8 VGND 0.01169f
C7267 XA.Cn[2].n0 VGND 0.02361f
C7268 XA.Cn[2].t7 VGND 0.01169f
C7269 XA.Cn[2].t6 VGND 0.01169f
C7270 XA.Cn[2].n1 VGND 0.02762f
C7271 XA.Cn[2].n2 VGND 0.07732f
C7272 XA.Cn[2].n3 VGND 0.01731f
C7273 XA.Cn[2].n4 VGND 0.01731f
C7274 XA.Cn[2].n5 VGND 0.01731f
C7275 XA.Cn[2].n6 VGND 0.02884f
C7276 XA.Cn[2].n7 VGND 0.08243f
C7277 XA.Cn[2].n8 VGND 0.05096f
C7278 XA.Cn[2].n9 VGND 0.05751f
C7279 XA.Cn[2].t18 VGND 0.01012f
C7280 XA.Cn[2].n10 VGND 0.02261f
C7281 XA.Cn[2].n11 VGND 0.01292f
C7282 XA.Cn[2].n12 VGND 0.01571f
C7283 XA.Cn[2].t35 VGND 0.01012f
C7284 XA.Cn[2].n13 VGND 0.02261f
C7285 XA.Cn[2].n14 VGND 0.01292f
C7286 XA.Cn[2].n15 VGND 0.07465f
C7287 XA.Cn[2].t37 VGND 0.01012f
C7288 XA.Cn[2].n16 VGND 0.02261f
C7289 XA.Cn[2].n17 VGND 0.01292f
C7290 XA.Cn[2].n18 VGND 0.07465f
C7291 XA.Cn[2].t39 VGND 0.01012f
C7292 XA.Cn[2].n19 VGND 0.02261f
C7293 XA.Cn[2].n20 VGND 0.01292f
C7294 XA.Cn[2].n21 VGND 0.07465f
C7295 XA.Cn[2].t28 VGND 0.01012f
C7296 XA.Cn[2].n22 VGND 0.02261f
C7297 XA.Cn[2].n23 VGND 0.01292f
C7298 XA.Cn[2].n24 VGND 0.07465f
C7299 XA.Cn[2].t29 VGND 0.01012f
C7300 XA.Cn[2].n25 VGND 0.02261f
C7301 XA.Cn[2].n26 VGND 0.01292f
C7302 XA.Cn[2].n27 VGND 0.07465f
C7303 XA.Cn[2].t42 VGND 0.01012f
C7304 XA.Cn[2].n28 VGND 0.02261f
C7305 XA.Cn[2].n29 VGND 0.01292f
C7306 XA.Cn[2].n30 VGND 0.07465f
C7307 XA.Cn[2].t19 VGND 0.01012f
C7308 XA.Cn[2].n31 VGND 0.02261f
C7309 XA.Cn[2].n32 VGND 0.01292f
C7310 XA.Cn[2].n33 VGND 0.07465f
C7311 XA.Cn[2].t21 VGND 0.01012f
C7312 XA.Cn[2].n34 VGND 0.02261f
C7313 XA.Cn[2].n35 VGND 0.01292f
C7314 XA.Cn[2].n36 VGND 0.07465f
C7315 XA.Cn[2].t40 VGND 0.01012f
C7316 XA.Cn[2].n37 VGND 0.02261f
C7317 XA.Cn[2].n38 VGND 0.01292f
C7318 XA.Cn[2].n39 VGND 0.07465f
C7319 XA.Cn[2].t41 VGND 0.01012f
C7320 XA.Cn[2].n40 VGND 0.02261f
C7321 XA.Cn[2].n41 VGND 0.01292f
C7322 XA.Cn[2].n42 VGND 0.07465f
C7323 XA.Cn[2].t22 VGND 0.01012f
C7324 XA.Cn[2].n43 VGND 0.02261f
C7325 XA.Cn[2].n44 VGND 0.01292f
C7326 XA.Cn[2].n45 VGND 0.07465f
C7327 XA.Cn[2].t30 VGND 0.01012f
C7328 XA.Cn[2].n46 VGND 0.02261f
C7329 XA.Cn[2].n47 VGND 0.01292f
C7330 XA.Cn[2].n48 VGND 0.07465f
C7331 XA.Cn[2].t33 VGND 0.01012f
C7332 XA.Cn[2].n49 VGND 0.02261f
C7333 XA.Cn[2].n50 VGND 0.01292f
C7334 XA.Cn[2].n51 VGND 0.07465f
C7335 XA.Cn[2].t14 VGND 0.01012f
C7336 XA.Cn[2].n52 VGND 0.02261f
C7337 XA.Cn[2].n53 VGND 0.01292f
C7338 XA.Cn[2].n54 VGND 0.07465f
C7339 XA.Cn[2].t24 VGND 0.01012f
C7340 XA.Cn[2].n55 VGND 0.02261f
C7341 XA.Cn[2].n56 VGND 0.01292f
C7342 XA.Cn[2].n57 VGND 0.07465f
C7343 XA.Cn[2].n58 VGND 0.27153f
C7344 XA.Cn[2].n59 VGND 0.0441f
C7345 XA.Cn[2].n60 VGND 0.02447f
C7346 XA.Cn[4].t5 VGND 0.01194f
C7347 XA.Cn[4].t4 VGND 0.01194f
C7348 XA.Cn[4].n0 VGND 0.02411f
C7349 XA.Cn[4].t7 VGND 0.01194f
C7350 XA.Cn[4].t6 VGND 0.01194f
C7351 XA.Cn[4].n1 VGND 0.02821f
C7352 XA.Cn[4].n2 VGND 0.07897f
C7353 XA.Cn[4].n3 VGND 0.01768f
C7354 XA.Cn[4].n4 VGND 0.01768f
C7355 XA.Cn[4].n5 VGND 0.01768f
C7356 XA.Cn[4].n6 VGND 0.02946f
C7357 XA.Cn[4].n7 VGND 0.0842f
C7358 XA.Cn[4].n8 VGND 0.05205f
C7359 XA.Cn[4].n9 VGND 0.05874f
C7360 XA.Cn[4].t26 VGND 0.01034f
C7361 XA.Cn[4].n10 VGND 0.02309f
C7362 XA.Cn[4].n11 VGND 0.0132f
C7363 XA.Cn[4].n12 VGND 0.01605f
C7364 XA.Cn[4].t43 VGND 0.01034f
C7365 XA.Cn[4].n13 VGND 0.02309f
C7366 XA.Cn[4].n14 VGND 0.0132f
C7367 XA.Cn[4].n15 VGND 0.07625f
C7368 XA.Cn[4].t13 VGND 0.01034f
C7369 XA.Cn[4].n16 VGND 0.02309f
C7370 XA.Cn[4].n17 VGND 0.0132f
C7371 XA.Cn[4].n18 VGND 0.07625f
C7372 XA.Cn[4].t15 VGND 0.01034f
C7373 XA.Cn[4].n19 VGND 0.02309f
C7374 XA.Cn[4].n20 VGND 0.0132f
C7375 XA.Cn[4].n21 VGND 0.07625f
C7376 XA.Cn[4].t36 VGND 0.01034f
C7377 XA.Cn[4].n22 VGND 0.02309f
C7378 XA.Cn[4].n23 VGND 0.0132f
C7379 XA.Cn[4].n24 VGND 0.07625f
C7380 XA.Cn[4].t37 VGND 0.01034f
C7381 XA.Cn[4].n25 VGND 0.02309f
C7382 XA.Cn[4].n26 VGND 0.0132f
C7383 XA.Cn[4].n27 VGND 0.07625f
C7384 XA.Cn[4].t18 VGND 0.01034f
C7385 XA.Cn[4].n28 VGND 0.02309f
C7386 XA.Cn[4].n29 VGND 0.0132f
C7387 XA.Cn[4].n30 VGND 0.07625f
C7388 XA.Cn[4].t27 VGND 0.01034f
C7389 XA.Cn[4].n31 VGND 0.02309f
C7390 XA.Cn[4].n32 VGND 0.0132f
C7391 XA.Cn[4].n33 VGND 0.07625f
C7392 XA.Cn[4].t29 VGND 0.01034f
C7393 XA.Cn[4].n34 VGND 0.02309f
C7394 XA.Cn[4].n35 VGND 0.0132f
C7395 XA.Cn[4].n36 VGND 0.07625f
C7396 XA.Cn[4].t16 VGND 0.01034f
C7397 XA.Cn[4].n37 VGND 0.02309f
C7398 XA.Cn[4].n38 VGND 0.0132f
C7399 XA.Cn[4].n39 VGND 0.07625f
C7400 XA.Cn[4].t17 VGND 0.01034f
C7401 XA.Cn[4].n40 VGND 0.02309f
C7402 XA.Cn[4].n41 VGND 0.0132f
C7403 XA.Cn[4].n42 VGND 0.07625f
C7404 XA.Cn[4].t30 VGND 0.01034f
C7405 XA.Cn[4].n43 VGND 0.02309f
C7406 XA.Cn[4].n44 VGND 0.0132f
C7407 XA.Cn[4].n45 VGND 0.07625f
C7408 XA.Cn[4].t38 VGND 0.01034f
C7409 XA.Cn[4].n46 VGND 0.02309f
C7410 XA.Cn[4].n47 VGND 0.0132f
C7411 XA.Cn[4].n48 VGND 0.07625f
C7412 XA.Cn[4].t41 VGND 0.01034f
C7413 XA.Cn[4].n49 VGND 0.02309f
C7414 XA.Cn[4].n50 VGND 0.0132f
C7415 XA.Cn[4].n51 VGND 0.07625f
C7416 XA.Cn[4].t22 VGND 0.01034f
C7417 XA.Cn[4].n52 VGND 0.02309f
C7418 XA.Cn[4].n53 VGND 0.0132f
C7419 XA.Cn[4].n54 VGND 0.07625f
C7420 XA.Cn[4].t32 VGND 0.01034f
C7421 XA.Cn[4].n55 VGND 0.02309f
C7422 XA.Cn[4].n56 VGND 0.0132f
C7423 XA.Cn[4].n57 VGND 0.07625f
C7424 XA.Cn[4].n58 VGND 0.23757f
C7425 XA.Cn[4].n59 VGND 0.04514f
C7426 XA.Cn[4].n60 VGND 0.025f
C7427 XThR.Tn[5].t6 VGND 0.01808f
C7428 XThR.Tn[5].t7 VGND 0.01808f
C7429 XThR.Tn[5].n0 VGND 0.03649f
C7430 XThR.Tn[5].t5 VGND 0.01808f
C7431 XThR.Tn[5].t4 VGND 0.01808f
C7432 XThR.Tn[5].n1 VGND 0.04269f
C7433 XThR.Tn[5].n2 VGND 0.11952f
C7434 XThR.Tn[5].t11 VGND 0.01175f
C7435 XThR.Tn[5].t8 VGND 0.01175f
C7436 XThR.Tn[5].n3 VGND 0.02676f
C7437 XThR.Tn[5].t10 VGND 0.01175f
C7438 XThR.Tn[5].t9 VGND 0.01175f
C7439 XThR.Tn[5].n4 VGND 0.02676f
C7440 XThR.Tn[5].t0 VGND 0.01175f
C7441 XThR.Tn[5].t1 VGND 0.01175f
C7442 XThR.Tn[5].n5 VGND 0.04459f
C7443 XThR.Tn[5].t3 VGND 0.01175f
C7444 XThR.Tn[5].t2 VGND 0.01175f
C7445 XThR.Tn[5].n6 VGND 0.02676f
C7446 XThR.Tn[5].n7 VGND 0.12743f
C7447 XThR.Tn[5].n8 VGND 0.07877f
C7448 XThR.Tn[5].n9 VGND 0.0889f
C7449 XThR.Tn[5].t17 VGND 0.01413f
C7450 XThR.Tn[5].t72 VGND 0.01547f
C7451 XThR.Tn[5].n10 VGND 0.03778f
C7452 XThR.Tn[5].n11 VGND 0.07257f
C7453 XThR.Tn[5].t39 VGND 0.01413f
C7454 XThR.Tn[5].t26 VGND 0.01547f
C7455 XThR.Tn[5].n12 VGND 0.03778f
C7456 XThR.Tn[5].t13 VGND 0.01408f
C7457 XThR.Tn[5].t23 VGND 0.01542f
C7458 XThR.Tn[5].n13 VGND 0.03931f
C7459 XThR.Tn[5].n14 VGND 0.02761f
C7460 XThR.Tn[5].n16 VGND 0.08862f
C7461 XThR.Tn[5].t73 VGND 0.01413f
C7462 XThR.Tn[5].t66 VGND 0.01547f
C7463 XThR.Tn[5].n17 VGND 0.03778f
C7464 XThR.Tn[5].t48 VGND 0.01408f
C7465 XThR.Tn[5].t61 VGND 0.01542f
C7466 XThR.Tn[5].n18 VGND 0.03931f
C7467 XThR.Tn[5].n19 VGND 0.02761f
C7468 XThR.Tn[5].n21 VGND 0.08862f
C7469 XThR.Tn[5].t28 VGND 0.01413f
C7470 XThR.Tn[5].t21 VGND 0.01547f
C7471 XThR.Tn[5].n22 VGND 0.03778f
C7472 XThR.Tn[5].t65 VGND 0.01408f
C7473 XThR.Tn[5].t18 VGND 0.01542f
C7474 XThR.Tn[5].n23 VGND 0.03931f
C7475 XThR.Tn[5].n24 VGND 0.02761f
C7476 XThR.Tn[5].n26 VGND 0.08862f
C7477 XThR.Tn[5].t55 VGND 0.01413f
C7478 XThR.Tn[5].t51 VGND 0.01547f
C7479 XThR.Tn[5].n27 VGND 0.03778f
C7480 XThR.Tn[5].t33 VGND 0.01408f
C7481 XThR.Tn[5].t46 VGND 0.01542f
C7482 XThR.Tn[5].n28 VGND 0.03931f
C7483 XThR.Tn[5].n29 VGND 0.02761f
C7484 XThR.Tn[5].n31 VGND 0.08862f
C7485 XThR.Tn[5].t30 VGND 0.01413f
C7486 XThR.Tn[5].t22 VGND 0.01547f
C7487 XThR.Tn[5].n32 VGND 0.03778f
C7488 XThR.Tn[5].t67 VGND 0.01408f
C7489 XThR.Tn[5].t19 VGND 0.01542f
C7490 XThR.Tn[5].n33 VGND 0.03931f
C7491 XThR.Tn[5].n34 VGND 0.02761f
C7492 XThR.Tn[5].n36 VGND 0.08862f
C7493 XThR.Tn[5].t69 VGND 0.01413f
C7494 XThR.Tn[5].t40 VGND 0.01547f
C7495 XThR.Tn[5].n37 VGND 0.03778f
C7496 XThR.Tn[5].t43 VGND 0.01408f
C7497 XThR.Tn[5].t37 VGND 0.01542f
C7498 XThR.Tn[5].n38 VGND 0.03931f
C7499 XThR.Tn[5].n39 VGND 0.02761f
C7500 XThR.Tn[5].n41 VGND 0.08862f
C7501 XThR.Tn[5].t38 VGND 0.01413f
C7502 XThR.Tn[5].t32 VGND 0.01547f
C7503 XThR.Tn[5].n42 VGND 0.03778f
C7504 XThR.Tn[5].t14 VGND 0.01408f
C7505 XThR.Tn[5].t29 VGND 0.01542f
C7506 XThR.Tn[5].n43 VGND 0.03931f
C7507 XThR.Tn[5].n44 VGND 0.02761f
C7508 XThR.Tn[5].n46 VGND 0.08862f
C7509 XThR.Tn[5].t42 VGND 0.01413f
C7510 XThR.Tn[5].t49 VGND 0.01547f
C7511 XThR.Tn[5].n47 VGND 0.03778f
C7512 XThR.Tn[5].t16 VGND 0.01408f
C7513 XThR.Tn[5].t45 VGND 0.01542f
C7514 XThR.Tn[5].n48 VGND 0.03931f
C7515 XThR.Tn[5].n49 VGND 0.02761f
C7516 XThR.Tn[5].n51 VGND 0.08862f
C7517 XThR.Tn[5].t58 VGND 0.01413f
C7518 XThR.Tn[5].t68 VGND 0.01547f
C7519 XThR.Tn[5].n52 VGND 0.03778f
C7520 XThR.Tn[5].t36 VGND 0.01408f
C7521 XThR.Tn[5].t63 VGND 0.01542f
C7522 XThR.Tn[5].n53 VGND 0.03931f
C7523 XThR.Tn[5].n54 VGND 0.02761f
C7524 XThR.Tn[5].n56 VGND 0.08862f
C7525 XThR.Tn[5].t53 VGND 0.01413f
C7526 XThR.Tn[5].t24 VGND 0.01547f
C7527 XThR.Tn[5].n57 VGND 0.03778f
C7528 XThR.Tn[5].t25 VGND 0.01408f
C7529 XThR.Tn[5].t20 VGND 0.01542f
C7530 XThR.Tn[5].n58 VGND 0.03931f
C7531 XThR.Tn[5].n59 VGND 0.02761f
C7532 XThR.Tn[5].n61 VGND 0.08862f
C7533 XThR.Tn[5].t71 VGND 0.01413f
C7534 XThR.Tn[5].t60 VGND 0.01547f
C7535 XThR.Tn[5].n62 VGND 0.03778f
C7536 XThR.Tn[5].t44 VGND 0.01408f
C7537 XThR.Tn[5].t57 VGND 0.01542f
C7538 XThR.Tn[5].n63 VGND 0.03931f
C7539 XThR.Tn[5].n64 VGND 0.02761f
C7540 XThR.Tn[5].n66 VGND 0.08862f
C7541 XThR.Tn[5].t41 VGND 0.01413f
C7542 XThR.Tn[5].t35 VGND 0.01547f
C7543 XThR.Tn[5].n67 VGND 0.03778f
C7544 XThR.Tn[5].t15 VGND 0.01408f
C7545 XThR.Tn[5].t31 VGND 0.01542f
C7546 XThR.Tn[5].n68 VGND 0.03931f
C7547 XThR.Tn[5].n69 VGND 0.02761f
C7548 XThR.Tn[5].n71 VGND 0.08862f
C7549 XThR.Tn[5].t56 VGND 0.01413f
C7550 XThR.Tn[5].t52 VGND 0.01547f
C7551 XThR.Tn[5].n72 VGND 0.03778f
C7552 XThR.Tn[5].t34 VGND 0.01408f
C7553 XThR.Tn[5].t47 VGND 0.01542f
C7554 XThR.Tn[5].n73 VGND 0.03931f
C7555 XThR.Tn[5].n74 VGND 0.02761f
C7556 XThR.Tn[5].n76 VGND 0.08862f
C7557 XThR.Tn[5].t12 VGND 0.01413f
C7558 XThR.Tn[5].t70 VGND 0.01547f
C7559 XThR.Tn[5].n77 VGND 0.03778f
C7560 XThR.Tn[5].t50 VGND 0.01408f
C7561 XThR.Tn[5].t64 VGND 0.01542f
C7562 XThR.Tn[5].n78 VGND 0.03931f
C7563 XThR.Tn[5].n79 VGND 0.02761f
C7564 XThR.Tn[5].n81 VGND 0.08862f
C7565 XThR.Tn[5].t54 VGND 0.01413f
C7566 XThR.Tn[5].t62 VGND 0.01547f
C7567 XThR.Tn[5].n82 VGND 0.03778f
C7568 XThR.Tn[5].t27 VGND 0.01408f
C7569 XThR.Tn[5].t59 VGND 0.01542f
C7570 XThR.Tn[5].n83 VGND 0.03931f
C7571 XThR.Tn[5].n84 VGND 0.02761f
C7572 XThR.Tn[5].n86 VGND 0.08862f
C7573 XThR.Tn[5].n87 VGND 0.08053f
C7574 XThR.Tn[5].n88 VGND 0.15597f
C7575 XThR.Tn[5].n89 VGND 0.03783f
C7576 XThR.Tn[3].t5 VGND 0.01821f
C7577 XThR.Tn[3].t6 VGND 0.01821f
C7578 XThR.Tn[3].n0 VGND 0.03675f
C7579 XThR.Tn[3].t4 VGND 0.01821f
C7580 XThR.Tn[3].t7 VGND 0.01821f
C7581 XThR.Tn[3].n1 VGND 0.043f
C7582 XThR.Tn[3].n2 VGND 0.12037f
C7583 XThR.Tn[3].t11 VGND 0.01183f
C7584 XThR.Tn[3].t8 VGND 0.01183f
C7585 XThR.Tn[3].n3 VGND 0.02695f
C7586 XThR.Tn[3].t10 VGND 0.01183f
C7587 XThR.Tn[3].t9 VGND 0.01183f
C7588 XThR.Tn[3].n4 VGND 0.02695f
C7589 XThR.Tn[3].t3 VGND 0.01183f
C7590 XThR.Tn[3].t1 VGND 0.01183f
C7591 XThR.Tn[3].n5 VGND 0.02695f
C7592 XThR.Tn[3].t0 VGND 0.01183f
C7593 XThR.Tn[3].t2 VGND 0.01183f
C7594 XThR.Tn[3].n6 VGND 0.0449f
C7595 XThR.Tn[3].n7 VGND 0.12834f
C7596 XThR.Tn[3].n8 VGND 0.07933f
C7597 XThR.Tn[3].n9 VGND 0.08953f
C7598 XThR.Tn[3].t64 VGND 0.01423f
C7599 XThR.Tn[3].t57 VGND 0.01558f
C7600 XThR.Tn[3].n10 VGND 0.03805f
C7601 XThR.Tn[3].n11 VGND 0.07309f
C7602 XThR.Tn[3].t18 VGND 0.01423f
C7603 XThR.Tn[3].t70 VGND 0.01558f
C7604 XThR.Tn[3].n12 VGND 0.03805f
C7605 XThR.Tn[3].t24 VGND 0.01418f
C7606 XThR.Tn[3].t55 VGND 0.01553f
C7607 XThR.Tn[3].n13 VGND 0.03959f
C7608 XThR.Tn[3].n14 VGND 0.02781f
C7609 XThR.Tn[3].n16 VGND 0.08925f
C7610 XThR.Tn[3].t59 VGND 0.01423f
C7611 XThR.Tn[3].t49 VGND 0.01558f
C7612 XThR.Tn[3].n17 VGND 0.03805f
C7613 XThR.Tn[3].t62 VGND 0.01418f
C7614 XThR.Tn[3].t29 VGND 0.01553f
C7615 XThR.Tn[3].n18 VGND 0.03959f
C7616 XThR.Tn[3].n19 VGND 0.02781f
C7617 XThR.Tn[3].n21 VGND 0.08925f
C7618 XThR.Tn[3].t71 VGND 0.01423f
C7619 XThR.Tn[3].t67 VGND 0.01558f
C7620 XThR.Tn[3].n22 VGND 0.03805f
C7621 XThR.Tn[3].t12 VGND 0.01418f
C7622 XThR.Tn[3].t47 VGND 0.01553f
C7623 XThR.Tn[3].n23 VGND 0.03959f
C7624 XThR.Tn[3].n24 VGND 0.02781f
C7625 XThR.Tn[3].n26 VGND 0.08925f
C7626 XThR.Tn[3].t39 VGND 0.01423f
C7627 XThR.Tn[3].t33 VGND 0.01558f
C7628 XThR.Tn[3].n27 VGND 0.03805f
C7629 XThR.Tn[3].t42 VGND 0.01418f
C7630 XThR.Tn[3].t13 VGND 0.01553f
C7631 XThR.Tn[3].n28 VGND 0.03959f
C7632 XThR.Tn[3].n29 VGND 0.02781f
C7633 XThR.Tn[3].n31 VGND 0.08925f
C7634 XThR.Tn[3].t72 VGND 0.01423f
C7635 XThR.Tn[3].t68 VGND 0.01558f
C7636 XThR.Tn[3].n32 VGND 0.03805f
C7637 XThR.Tn[3].t16 VGND 0.01418f
C7638 XThR.Tn[3].t48 VGND 0.01553f
C7639 XThR.Tn[3].n33 VGND 0.03959f
C7640 XThR.Tn[3].n34 VGND 0.02781f
C7641 XThR.Tn[3].n36 VGND 0.08925f
C7642 XThR.Tn[3].t52 VGND 0.01423f
C7643 XThR.Tn[3].t20 VGND 0.01558f
C7644 XThR.Tn[3].n37 VGND 0.03805f
C7645 XThR.Tn[3].t56 VGND 0.01418f
C7646 XThR.Tn[3].t66 VGND 0.01553f
C7647 XThR.Tn[3].n38 VGND 0.03959f
C7648 XThR.Tn[3].n39 VGND 0.02781f
C7649 XThR.Tn[3].n41 VGND 0.08925f
C7650 XThR.Tn[3].t19 VGND 0.01423f
C7651 XThR.Tn[3].t14 VGND 0.01558f
C7652 XThR.Tn[3].n42 VGND 0.03805f
C7653 XThR.Tn[3].t23 VGND 0.01418f
C7654 XThR.Tn[3].t61 VGND 0.01553f
C7655 XThR.Tn[3].n43 VGND 0.03959f
C7656 XThR.Tn[3].n44 VGND 0.02781f
C7657 XThR.Tn[3].n46 VGND 0.08925f
C7658 XThR.Tn[3].t22 VGND 0.01423f
C7659 XThR.Tn[3].t31 VGND 0.01558f
C7660 XThR.Tn[3].n47 VGND 0.03805f
C7661 XThR.Tn[3].t28 VGND 0.01418f
C7662 XThR.Tn[3].t73 VGND 0.01553f
C7663 XThR.Tn[3].n48 VGND 0.03959f
C7664 XThR.Tn[3].n49 VGND 0.02781f
C7665 XThR.Tn[3].n51 VGND 0.08925f
C7666 XThR.Tn[3].t41 VGND 0.01423f
C7667 XThR.Tn[3].t51 VGND 0.01558f
C7668 XThR.Tn[3].n52 VGND 0.03805f
C7669 XThR.Tn[3].t45 VGND 0.01418f
C7670 XThR.Tn[3].t30 VGND 0.01553f
C7671 XThR.Tn[3].n53 VGND 0.03959f
C7672 XThR.Tn[3].n54 VGND 0.02781f
C7673 XThR.Tn[3].n56 VGND 0.08925f
C7674 XThR.Tn[3].t35 VGND 0.01423f
C7675 XThR.Tn[3].t69 VGND 0.01558f
C7676 XThR.Tn[3].n57 VGND 0.03805f
C7677 XThR.Tn[3].t37 VGND 0.01418f
C7678 XThR.Tn[3].t50 VGND 0.01553f
C7679 XThR.Tn[3].n58 VGND 0.03959f
C7680 XThR.Tn[3].n59 VGND 0.02781f
C7681 XThR.Tn[3].n61 VGND 0.08925f
C7682 XThR.Tn[3].t54 VGND 0.01423f
C7683 XThR.Tn[3].t44 VGND 0.01558f
C7684 XThR.Tn[3].n62 VGND 0.03805f
C7685 XThR.Tn[3].t58 VGND 0.01418f
C7686 XThR.Tn[3].t25 VGND 0.01553f
C7687 XThR.Tn[3].n63 VGND 0.03959f
C7688 XThR.Tn[3].n64 VGND 0.02781f
C7689 XThR.Tn[3].n66 VGND 0.08925f
C7690 XThR.Tn[3].t21 VGND 0.01423f
C7691 XThR.Tn[3].t17 VGND 0.01558f
C7692 XThR.Tn[3].n67 VGND 0.03805f
C7693 XThR.Tn[3].t26 VGND 0.01418f
C7694 XThR.Tn[3].t63 VGND 0.01553f
C7695 XThR.Tn[3].n68 VGND 0.03959f
C7696 XThR.Tn[3].n69 VGND 0.02781f
C7697 XThR.Tn[3].n71 VGND 0.08925f
C7698 XThR.Tn[3].t40 VGND 0.01423f
C7699 XThR.Tn[3].t34 VGND 0.01558f
C7700 XThR.Tn[3].n72 VGND 0.03805f
C7701 XThR.Tn[3].t43 VGND 0.01418f
C7702 XThR.Tn[3].t15 VGND 0.01553f
C7703 XThR.Tn[3].n73 VGND 0.03959f
C7704 XThR.Tn[3].n74 VGND 0.02781f
C7705 XThR.Tn[3].n76 VGND 0.08925f
C7706 XThR.Tn[3].t60 VGND 0.01423f
C7707 XThR.Tn[3].t53 VGND 0.01558f
C7708 XThR.Tn[3].n77 VGND 0.03805f
C7709 XThR.Tn[3].t65 VGND 0.01418f
C7710 XThR.Tn[3].t32 VGND 0.01553f
C7711 XThR.Tn[3].n78 VGND 0.03959f
C7712 XThR.Tn[3].n79 VGND 0.02781f
C7713 XThR.Tn[3].n81 VGND 0.08925f
C7714 XThR.Tn[3].t36 VGND 0.01423f
C7715 XThR.Tn[3].t46 VGND 0.01558f
C7716 XThR.Tn[3].n82 VGND 0.03805f
C7717 XThR.Tn[3].t38 VGND 0.01418f
C7718 XThR.Tn[3].t27 VGND 0.01553f
C7719 XThR.Tn[3].n83 VGND 0.03959f
C7720 XThR.Tn[3].n84 VGND 0.02781f
C7721 XThR.Tn[3].n86 VGND 0.08925f
C7722 XThR.Tn[3].n87 VGND 0.0811f
C7723 XThR.Tn[3].n88 VGND 0.17963f
C7724 XThR.Tn[3].n89 VGND 0.0381f
C7725 thermo15c_0.XTB4.Y.t4 VGND 0.02956f
C7726 thermo15c_0.XTB4.Y.t13 VGND 0.05016f
C7727 thermo15c_0.XTB4.Y.n0 VGND 0.05972f
C7728 thermo15c_0.XTB4.Y.t7 VGND 0.02956f
C7729 thermo15c_0.XTB4.Y.t17 VGND 0.05016f
C7730 thermo15c_0.XTB4.Y.n1 VGND 0.03074f
C7731 thermo15c_0.XTB4.Y.t10 VGND 0.02956f
C7732 thermo15c_0.XTB4.Y.t2 VGND 0.05016f
C7733 thermo15c_0.XTB4.Y.n2 VGND 0.06603f
C7734 thermo15c_0.XTB4.Y.t14 VGND 0.02956f
C7735 thermo15c_0.XTB4.Y.t3 VGND 0.05016f
C7736 thermo15c_0.XTB4.Y.n3 VGND 0.0613f
C7737 thermo15c_0.XTB4.Y.n4 VGND 0.03729f
C7738 thermo15c_0.XTB4.Y.n5 VGND 0.06174f
C7739 thermo15c_0.XTB4.Y.n6 VGND 0.02389f
C7740 thermo15c_0.XTB4.Y.n7 VGND 0.02916f
C7741 thermo15c_0.XTB4.Y.n8 VGND 0.06603f
C7742 thermo15c_0.XTB4.Y.n9 VGND 0.0331f
C7743 thermo15c_0.XTB4.Y.n10 VGND 0.06459f
C7744 thermo15c_0.XTB4.Y.t5 VGND 0.02956f
C7745 thermo15c_0.XTB4.Y.t16 VGND 0.05016f
C7746 thermo15c_0.XTB4.Y.n11 VGND 0.06761f
C7747 thermo15c_0.XTB4.Y.t9 VGND 0.02956f
C7748 thermo15c_0.XTB4.Y.t6 VGND 0.05016f
C7749 thermo15c_0.XTB4.Y.t15 VGND 0.02956f
C7750 thermo15c_0.XTB4.Y.t12 VGND 0.05016f
C7751 thermo15c_0.XTB4.Y.t11 VGND 0.02956f
C7752 thermo15c_0.XTB4.Y.t8 VGND 0.05016f
C7753 thermo15c_0.XTB4.Y.n12 VGND 0.08416f
C7754 thermo15c_0.XTB4.Y.n13 VGND 0.08889f
C7755 thermo15c_0.XTB4.Y.n14 VGND 0.03426f
C7756 thermo15c_0.XTB4.Y.n15 VGND 0.07234f
C7757 thermo15c_0.XTB4.Y.n16 VGND 0.0331f
C7758 thermo15c_0.XTB4.Y.n17 VGND 0.02701f
C7759 thermo15c_0.XTB4.Y.n18 VGND 0.63971f
C7760 thermo15c_0.XTB4.Y.n19 VGND 1.30917f
C7761 thermo15c_0.XTB4.Y.t1 VGND 0.06491f
C7762 thermo15c_0.XTB4.Y.n20 VGND 0.11223f
C7763 thermo15c_0.XTB4.Y.t0 VGND 0.12238f
C7764 thermo15c_0.XTB4.Y.n21 VGND 0.16166f
C7765 XA.Cn[0].t4 VGND 0.0118f
C7766 XA.Cn[0].t3 VGND 0.0118f
C7767 XA.Cn[0].n0 VGND 0.02383f
C7768 XA.Cn[0].t6 VGND 0.0118f
C7769 XA.Cn[0].t5 VGND 0.0118f
C7770 XA.Cn[0].n1 VGND 0.02788f
C7771 XA.Cn[0].n2 VGND 0.07804f
C7772 XA.Cn[0].n3 VGND 0.01747f
C7773 XA.Cn[0].n4 VGND 0.01747f
C7774 XA.Cn[0].n5 VGND 0.01747f
C7775 XA.Cn[0].n6 VGND 0.02911f
C7776 XA.Cn[0].n7 VGND 0.0832f
C7777 XA.Cn[0].n8 VGND 0.05143f
C7778 XA.Cn[0].n9 VGND 0.05805f
C7779 XA.Cn[0].t22 VGND 0.01022f
C7780 XA.Cn[0].n10 VGND 0.02282f
C7781 XA.Cn[0].n11 VGND 0.01304f
C7782 XA.Cn[0].n12 VGND 0.01586f
C7783 XA.Cn[0].t41 VGND 0.01022f
C7784 XA.Cn[0].n13 VGND 0.02282f
C7785 XA.Cn[0].n14 VGND 0.01304f
C7786 XA.Cn[0].n15 VGND 0.07535f
C7787 XA.Cn[0].t12 VGND 0.01022f
C7788 XA.Cn[0].n16 VGND 0.02282f
C7789 XA.Cn[0].n17 VGND 0.01304f
C7790 XA.Cn[0].n18 VGND 0.07535f
C7791 XA.Cn[0].t13 VGND 0.01022f
C7792 XA.Cn[0].n19 VGND 0.02282f
C7793 XA.Cn[0].n20 VGND 0.01304f
C7794 XA.Cn[0].n21 VGND 0.07535f
C7795 XA.Cn[0].t32 VGND 0.01022f
C7796 XA.Cn[0].n22 VGND 0.02282f
C7797 XA.Cn[0].n23 VGND 0.01304f
C7798 XA.Cn[0].n24 VGND 0.07535f
C7799 XA.Cn[0].t34 VGND 0.01022f
C7800 XA.Cn[0].n25 VGND 0.02282f
C7801 XA.Cn[0].n26 VGND 0.01304f
C7802 XA.Cn[0].n27 VGND 0.07535f
C7803 XA.Cn[0].t17 VGND 0.01022f
C7804 XA.Cn[0].n28 VGND 0.02282f
C7805 XA.Cn[0].n29 VGND 0.01304f
C7806 XA.Cn[0].n30 VGND 0.07535f
C7807 XA.Cn[0].t25 VGND 0.01022f
C7808 XA.Cn[0].n31 VGND 0.02282f
C7809 XA.Cn[0].n32 VGND 0.01304f
C7810 XA.Cn[0].n33 VGND 0.07535f
C7811 XA.Cn[0].t26 VGND 0.01022f
C7812 XA.Cn[0].n34 VGND 0.02282f
C7813 XA.Cn[0].n35 VGND 0.01304f
C7814 XA.Cn[0].n36 VGND 0.07535f
C7815 XA.Cn[0].t15 VGND 0.01022f
C7816 XA.Cn[0].n37 VGND 0.02282f
C7817 XA.Cn[0].n38 VGND 0.01304f
C7818 XA.Cn[0].n39 VGND 0.07535f
C7819 XA.Cn[0].t16 VGND 0.01022f
C7820 XA.Cn[0].n40 VGND 0.02282f
C7821 XA.Cn[0].n41 VGND 0.01304f
C7822 XA.Cn[0].n42 VGND 0.07535f
C7823 XA.Cn[0].t27 VGND 0.01022f
C7824 XA.Cn[0].n43 VGND 0.02282f
C7825 XA.Cn[0].n44 VGND 0.01304f
C7826 XA.Cn[0].n45 VGND 0.07535f
C7827 XA.Cn[0].t36 VGND 0.01022f
C7828 XA.Cn[0].n46 VGND 0.02282f
C7829 XA.Cn[0].n47 VGND 0.01304f
C7830 XA.Cn[0].n48 VGND 0.07535f
C7831 XA.Cn[0].t38 VGND 0.01022f
C7832 XA.Cn[0].n49 VGND 0.02282f
C7833 XA.Cn[0].n50 VGND 0.01304f
C7834 XA.Cn[0].n51 VGND 0.07535f
C7835 XA.Cn[0].t19 VGND 0.01022f
C7836 XA.Cn[0].n52 VGND 0.02282f
C7837 XA.Cn[0].n53 VGND 0.01304f
C7838 XA.Cn[0].n54 VGND 0.07535f
C7839 XA.Cn[0].t29 VGND 0.01022f
C7840 XA.Cn[0].n55 VGND 0.02282f
C7841 XA.Cn[0].n56 VGND 0.01304f
C7842 XA.Cn[0].n57 VGND 0.07535f
C7843 XA.Cn[0].n58 VGND 0.13474f
C7844 XA.Cn[0].n59 VGND 0.03416f
C7845 XA.Cn[0].n60 VGND 0.0247f
C7846 XA.Cn[13].n0 VGND 0.02342f
C7847 XA.Cn[13].n1 VGND 0.01878f
C7848 XA.Cn[13].n2 VGND 0.04331f
C7849 XA.Cn[13].t29 VGND 0.01145f
C7850 XA.Cn[13].t27 VGND 0.01251f
C7851 XA.Cn[13].n3 VGND 0.02793f
C7852 XA.Cn[13].n4 VGND 0.01596f
C7853 XA.Cn[13].n5 VGND 0.01941f
C7854 XA.Cn[13].t15 VGND 0.01145f
C7855 XA.Cn[13].t12 VGND 0.01251f
C7856 XA.Cn[13].n6 VGND 0.02793f
C7857 XA.Cn[13].n7 VGND 0.01596f
C7858 XA.Cn[13].n8 VGND 0.09223f
C7859 XA.Cn[13].t20 VGND 0.01145f
C7860 XA.Cn[13].t14 VGND 0.01251f
C7861 XA.Cn[13].n9 VGND 0.02793f
C7862 XA.Cn[13].n10 VGND 0.01596f
C7863 XA.Cn[13].n11 VGND 0.09223f
C7864 XA.Cn[13].t21 VGND 0.01145f
C7865 XA.Cn[13].t16 VGND 0.01251f
C7866 XA.Cn[13].n12 VGND 0.02793f
C7867 XA.Cn[13].n13 VGND 0.01596f
C7868 XA.Cn[13].n14 VGND 0.09223f
C7869 XA.Cn[13].t40 VGND 0.01145f
C7870 XA.Cn[13].t37 VGND 0.01251f
C7871 XA.Cn[13].n15 VGND 0.02793f
C7872 XA.Cn[13].n16 VGND 0.01596f
C7873 XA.Cn[13].n17 VGND 0.09223f
C7874 XA.Cn[13].t41 VGND 0.01145f
C7875 XA.Cn[13].t38 VGND 0.01251f
C7876 XA.Cn[13].n18 VGND 0.02793f
C7877 XA.Cn[13].n19 VGND 0.01596f
C7878 XA.Cn[13].n20 VGND 0.09223f
C7879 XA.Cn[13].t25 VGND 0.01145f
C7880 XA.Cn[13].t19 VGND 0.01251f
C7881 XA.Cn[13].n21 VGND 0.02793f
C7882 XA.Cn[13].n22 VGND 0.01596f
C7883 XA.Cn[13].n23 VGND 0.09223f
C7884 XA.Cn[13].t32 VGND 0.01145f
C7885 XA.Cn[13].t28 VGND 0.01251f
C7886 XA.Cn[13].n24 VGND 0.02793f
C7887 XA.Cn[13].n25 VGND 0.01596f
C7888 XA.Cn[13].n26 VGND 0.09223f
C7889 XA.Cn[13].t34 VGND 0.01145f
C7890 XA.Cn[13].t30 VGND 0.01251f
C7891 XA.Cn[13].n27 VGND 0.02793f
C7892 XA.Cn[13].n28 VGND 0.01596f
C7893 XA.Cn[13].n29 VGND 0.09223f
C7894 XA.Cn[13].t22 VGND 0.01145f
C7895 XA.Cn[13].t17 VGND 0.01251f
C7896 XA.Cn[13].n30 VGND 0.02793f
C7897 XA.Cn[13].n31 VGND 0.01596f
C7898 XA.Cn[13].n32 VGND 0.09223f
C7899 XA.Cn[13].t24 VGND 0.01145f
C7900 XA.Cn[13].t18 VGND 0.01251f
C7901 XA.Cn[13].n33 VGND 0.02793f
C7902 XA.Cn[13].n34 VGND 0.01596f
C7903 XA.Cn[13].n35 VGND 0.09223f
C7904 XA.Cn[13].t35 VGND 0.01145f
C7905 XA.Cn[13].t31 VGND 0.01251f
C7906 XA.Cn[13].n36 VGND 0.02793f
C7907 XA.Cn[13].n37 VGND 0.01596f
C7908 XA.Cn[13].n38 VGND 0.09223f
C7909 XA.Cn[13].t43 VGND 0.01145f
C7910 XA.Cn[13].t39 VGND 0.01251f
C7911 XA.Cn[13].n39 VGND 0.02793f
C7912 XA.Cn[13].n40 VGND 0.01596f
C7913 XA.Cn[13].n41 VGND 0.09223f
C7914 XA.Cn[13].t13 VGND 0.01145f
C7915 XA.Cn[13].t42 VGND 0.01251f
C7916 XA.Cn[13].n42 VGND 0.02793f
C7917 XA.Cn[13].n43 VGND 0.01596f
C7918 XA.Cn[13].n44 VGND 0.09223f
C7919 XA.Cn[13].t26 VGND 0.01145f
C7920 XA.Cn[13].t23 VGND 0.01251f
C7921 XA.Cn[13].n45 VGND 0.02793f
C7922 XA.Cn[13].n46 VGND 0.01596f
C7923 XA.Cn[13].n47 VGND 0.09223f
C7924 XA.Cn[13].t36 VGND 0.01145f
C7925 XA.Cn[13].t33 VGND 0.01251f
C7926 XA.Cn[13].n48 VGND 0.02793f
C7927 XA.Cn[13].n49 VGND 0.01596f
C7928 XA.Cn[13].n50 VGND 0.09223f
C7929 XA.Cn[13].n51 VGND 0.51097f
C7930 XA.Cn[13].n52 VGND 0.04181f
C7931 XA.Cn[13].t2 VGND 0.01445f
C7932 XA.Cn[13].t1 VGND 0.01445f
C7933 XA.Cn[13].n53 VGND 0.03122f
C7934 XA.Cn[13].t0 VGND 0.01445f
C7935 XA.Cn[13].t3 VGND 0.01445f
C7936 XA.Cn[13].n54 VGND 0.04921f
C7937 XA.Cn[13].n55 VGND 0.13032f
C7938 XA.Cn[13].t9 VGND 0.01445f
C7939 XA.Cn[13].t8 VGND 0.01445f
C7940 XA.Cn[13].n57 VGND 0.04387f
C7941 XA.Cn[13].t11 VGND 0.01445f
C7942 XA.Cn[13].t10 VGND 0.01445f
C7943 XA.Cn[13].n58 VGND 0.03212f
C7944 XA.Cn[13].n59 VGND 0.14294f
C7945 XA.Cn[12].n0 VGND 0.02348f
C7946 XA.Cn[12].n1 VGND 0.01883f
C7947 XA.Cn[12].n2 VGND 0.04736f
C7948 XA.Cn[12].t37 VGND 0.01148f
C7949 XA.Cn[12].t35 VGND 0.01254f
C7950 XA.Cn[12].n3 VGND 0.028f
C7951 XA.Cn[12].n4 VGND 0.016f
C7952 XA.Cn[12].n5 VGND 0.01946f
C7953 XA.Cn[12].t23 VGND 0.01148f
C7954 XA.Cn[12].t20 VGND 0.01254f
C7955 XA.Cn[12].n6 VGND 0.028f
C7956 XA.Cn[12].n7 VGND 0.016f
C7957 XA.Cn[12].n8 VGND 0.09245f
C7958 XA.Cn[12].t28 VGND 0.01148f
C7959 XA.Cn[12].t22 VGND 0.01254f
C7960 XA.Cn[12].n9 VGND 0.028f
C7961 XA.Cn[12].n10 VGND 0.016f
C7962 XA.Cn[12].n11 VGND 0.09245f
C7963 XA.Cn[12].t29 VGND 0.01148f
C7964 XA.Cn[12].t24 VGND 0.01254f
C7965 XA.Cn[12].n12 VGND 0.028f
C7966 XA.Cn[12].n13 VGND 0.016f
C7967 XA.Cn[12].n14 VGND 0.09245f
C7968 XA.Cn[12].t16 VGND 0.01148f
C7969 XA.Cn[12].t13 VGND 0.01254f
C7970 XA.Cn[12].n15 VGND 0.028f
C7971 XA.Cn[12].n16 VGND 0.016f
C7972 XA.Cn[12].n17 VGND 0.09245f
C7973 XA.Cn[12].t17 VGND 0.01148f
C7974 XA.Cn[12].t14 VGND 0.01254f
C7975 XA.Cn[12].n18 VGND 0.028f
C7976 XA.Cn[12].n19 VGND 0.016f
C7977 XA.Cn[12].n20 VGND 0.09245f
C7978 XA.Cn[12].t33 VGND 0.01148f
C7979 XA.Cn[12].t27 VGND 0.01254f
C7980 XA.Cn[12].n21 VGND 0.028f
C7981 XA.Cn[12].n22 VGND 0.016f
C7982 XA.Cn[12].n23 VGND 0.09245f
C7983 XA.Cn[12].t40 VGND 0.01148f
C7984 XA.Cn[12].t36 VGND 0.01254f
C7985 XA.Cn[12].n24 VGND 0.028f
C7986 XA.Cn[12].n25 VGND 0.016f
C7987 XA.Cn[12].n26 VGND 0.09245f
C7988 XA.Cn[12].t42 VGND 0.01148f
C7989 XA.Cn[12].t38 VGND 0.01254f
C7990 XA.Cn[12].n27 VGND 0.028f
C7991 XA.Cn[12].n28 VGND 0.016f
C7992 XA.Cn[12].n29 VGND 0.09245f
C7993 XA.Cn[12].t30 VGND 0.01148f
C7994 XA.Cn[12].t25 VGND 0.01254f
C7995 XA.Cn[12].n30 VGND 0.028f
C7996 XA.Cn[12].n31 VGND 0.016f
C7997 XA.Cn[12].n32 VGND 0.09245f
C7998 XA.Cn[12].t32 VGND 0.01148f
C7999 XA.Cn[12].t26 VGND 0.01254f
C8000 XA.Cn[12].n33 VGND 0.028f
C8001 XA.Cn[12].n34 VGND 0.016f
C8002 XA.Cn[12].n35 VGND 0.09245f
C8003 XA.Cn[12].t43 VGND 0.01148f
C8004 XA.Cn[12].t39 VGND 0.01254f
C8005 XA.Cn[12].n36 VGND 0.028f
C8006 XA.Cn[12].n37 VGND 0.016f
C8007 XA.Cn[12].n38 VGND 0.09245f
C8008 XA.Cn[12].t19 VGND 0.01148f
C8009 XA.Cn[12].t15 VGND 0.01254f
C8010 XA.Cn[12].n39 VGND 0.028f
C8011 XA.Cn[12].n40 VGND 0.016f
C8012 XA.Cn[12].n41 VGND 0.09245f
C8013 XA.Cn[12].t21 VGND 0.01148f
C8014 XA.Cn[12].t18 VGND 0.01254f
C8015 XA.Cn[12].n42 VGND 0.028f
C8016 XA.Cn[12].n43 VGND 0.016f
C8017 XA.Cn[12].n44 VGND 0.09245f
C8018 XA.Cn[12].t34 VGND 0.01148f
C8019 XA.Cn[12].t31 VGND 0.01254f
C8020 XA.Cn[12].n45 VGND 0.028f
C8021 XA.Cn[12].n46 VGND 0.016f
C8022 XA.Cn[12].n47 VGND 0.09245f
C8023 XA.Cn[12].t12 VGND 0.01148f
C8024 XA.Cn[12].t41 VGND 0.01254f
C8025 XA.Cn[12].n48 VGND 0.028f
C8026 XA.Cn[12].n49 VGND 0.016f
C8027 XA.Cn[12].n50 VGND 0.09245f
C8028 XA.Cn[12].n51 VGND 0.5067f
C8029 XA.Cn[12].n52 VGND 0.03519f
C8030 XA.Cn[12].t1 VGND 0.01448f
C8031 XA.Cn[12].t2 VGND 0.01448f
C8032 XA.Cn[12].n53 VGND 0.03129f
C8033 XA.Cn[12].t0 VGND 0.01448f
C8034 XA.Cn[12].t3 VGND 0.01448f
C8035 XA.Cn[12].n54 VGND 0.04762f
C8036 XA.Cn[12].n55 VGND 0.13232f
C8037 XA.Cn[12].n56 VGND 0.02081f
C8038 XA.Cn[12].t9 VGND 0.01448f
C8039 XA.Cn[12].t8 VGND 0.01448f
C8040 XA.Cn[12].n57 VGND 0.04397f
C8041 XA.Cn[12].t11 VGND 0.01448f
C8042 XA.Cn[12].t10 VGND 0.01448f
C8043 XA.Cn[12].n58 VGND 0.03219f
C8044 XA.Cn[12].n59 VGND 0.14328f
C8045 XA.Cn[11].t11 VGND 0.01474f
C8046 XA.Cn[11].t8 VGND 0.01474f
C8047 XA.Cn[11].n0 VGND 0.03186f
C8048 XA.Cn[11].t1 VGND 0.01474f
C8049 XA.Cn[11].t7 VGND 0.01474f
C8050 XA.Cn[11].n1 VGND 0.05022f
C8051 XA.Cn[11].n2 VGND 0.13299f
C8052 XA.Cn[11].t2 VGND 0.01474f
C8053 XA.Cn[11].t5 VGND 0.01474f
C8054 XA.Cn[11].n3 VGND 0.04477f
C8055 XA.Cn[11].t4 VGND 0.01474f
C8056 XA.Cn[11].t3 VGND 0.01474f
C8057 XA.Cn[11].n4 VGND 0.03278f
C8058 XA.Cn[11].n5 VGND 0.14588f
C8059 XA.Cn[11].t20 VGND 0.01169f
C8060 XA.Cn[11].t18 VGND 0.01277f
C8061 XA.Cn[11].n7 VGND 0.02851f
C8062 XA.Cn[11].n8 VGND 0.01629f
C8063 XA.Cn[11].n9 VGND 0.01981f
C8064 XA.Cn[11].t38 VGND 0.01169f
C8065 XA.Cn[11].t35 VGND 0.01277f
C8066 XA.Cn[11].n10 VGND 0.02851f
C8067 XA.Cn[11].n11 VGND 0.01629f
C8068 XA.Cn[11].n12 VGND 0.09412f
C8069 XA.Cn[11].t43 VGND 0.01169f
C8070 XA.Cn[11].t37 VGND 0.01277f
C8071 XA.Cn[11].n13 VGND 0.02851f
C8072 XA.Cn[11].n14 VGND 0.01629f
C8073 XA.Cn[11].n15 VGND 0.09412f
C8074 XA.Cn[11].t12 VGND 0.01169f
C8075 XA.Cn[11].t39 VGND 0.01277f
C8076 XA.Cn[11].n16 VGND 0.02851f
C8077 XA.Cn[11].n17 VGND 0.01629f
C8078 XA.Cn[11].n18 VGND 0.09412f
C8079 XA.Cn[11].t31 VGND 0.01169f
C8080 XA.Cn[11].t28 VGND 0.01277f
C8081 XA.Cn[11].n19 VGND 0.02851f
C8082 XA.Cn[11].n20 VGND 0.01629f
C8083 XA.Cn[11].n21 VGND 0.09412f
C8084 XA.Cn[11].t32 VGND 0.01169f
C8085 XA.Cn[11].t29 VGND 0.01277f
C8086 XA.Cn[11].n22 VGND 0.02851f
C8087 XA.Cn[11].n23 VGND 0.01629f
C8088 XA.Cn[11].n24 VGND 0.09412f
C8089 XA.Cn[11].t16 VGND 0.01169f
C8090 XA.Cn[11].t42 VGND 0.01277f
C8091 XA.Cn[11].n25 VGND 0.02851f
C8092 XA.Cn[11].n26 VGND 0.01629f
C8093 XA.Cn[11].n27 VGND 0.09412f
C8094 XA.Cn[11].t23 VGND 0.01169f
C8095 XA.Cn[11].t19 VGND 0.01277f
C8096 XA.Cn[11].n28 VGND 0.02851f
C8097 XA.Cn[11].n29 VGND 0.01629f
C8098 XA.Cn[11].n30 VGND 0.09412f
C8099 XA.Cn[11].t25 VGND 0.01169f
C8100 XA.Cn[11].t21 VGND 0.01277f
C8101 XA.Cn[11].n31 VGND 0.02851f
C8102 XA.Cn[11].n32 VGND 0.01629f
C8103 XA.Cn[11].n33 VGND 0.09412f
C8104 XA.Cn[11].t13 VGND 0.01169f
C8105 XA.Cn[11].t40 VGND 0.01277f
C8106 XA.Cn[11].n34 VGND 0.02851f
C8107 XA.Cn[11].n35 VGND 0.01629f
C8108 XA.Cn[11].n36 VGND 0.09412f
C8109 XA.Cn[11].t15 VGND 0.01169f
C8110 XA.Cn[11].t41 VGND 0.01277f
C8111 XA.Cn[11].n37 VGND 0.02851f
C8112 XA.Cn[11].n38 VGND 0.01629f
C8113 XA.Cn[11].n39 VGND 0.09412f
C8114 XA.Cn[11].t26 VGND 0.01169f
C8115 XA.Cn[11].t22 VGND 0.01277f
C8116 XA.Cn[11].n40 VGND 0.02851f
C8117 XA.Cn[11].n41 VGND 0.01629f
C8118 XA.Cn[11].n42 VGND 0.09412f
C8119 XA.Cn[11].t34 VGND 0.01169f
C8120 XA.Cn[11].t30 VGND 0.01277f
C8121 XA.Cn[11].n43 VGND 0.02851f
C8122 XA.Cn[11].n44 VGND 0.01629f
C8123 XA.Cn[11].n45 VGND 0.09412f
C8124 XA.Cn[11].t36 VGND 0.01169f
C8125 XA.Cn[11].t33 VGND 0.01277f
C8126 XA.Cn[11].n46 VGND 0.02851f
C8127 XA.Cn[11].n47 VGND 0.01629f
C8128 XA.Cn[11].n48 VGND 0.09412f
C8129 XA.Cn[11].t17 VGND 0.01169f
C8130 XA.Cn[11].t14 VGND 0.01277f
C8131 XA.Cn[11].n49 VGND 0.02851f
C8132 XA.Cn[11].n50 VGND 0.01629f
C8133 XA.Cn[11].n51 VGND 0.09412f
C8134 XA.Cn[11].t27 VGND 0.01169f
C8135 XA.Cn[11].t24 VGND 0.01277f
C8136 XA.Cn[11].n52 VGND 0.02851f
C8137 XA.Cn[11].n53 VGND 0.01629f
C8138 XA.Cn[11].n54 VGND 0.09412f
C8139 XA.Cn[11].n55 VGND 0.04302f
C8140 XA.Cn[11].n56 VGND 0.0239f
C8141 XA.Cn[11].n57 VGND 0.01917f
C8142 XA.Cn[11].n58 VGND 0.0442f
C8143 XA.Cn[9].n0 VGND 0.02381f
C8144 XA.Cn[9].n1 VGND 0.0191f
C8145 XA.Cn[9].n2 VGND 0.04403f
C8146 XA.Cn[9].t26 VGND 0.01164f
C8147 XA.Cn[9].t12 VGND 0.01272f
C8148 XA.Cn[9].n3 VGND 0.0284f
C8149 XA.Cn[9].n4 VGND 0.01623f
C8150 XA.Cn[9].n5 VGND 0.01974f
C8151 XA.Cn[9].t13 VGND 0.01164f
C8152 XA.Cn[9].t30 VGND 0.01272f
C8153 XA.Cn[9].n6 VGND 0.0284f
C8154 XA.Cn[9].n7 VGND 0.01623f
C8155 XA.Cn[9].n8 VGND 0.09378f
C8156 XA.Cn[9].t15 VGND 0.01164f
C8157 XA.Cn[9].t34 VGND 0.01272f
C8158 XA.Cn[9].n9 VGND 0.0284f
C8159 XA.Cn[9].n10 VGND 0.01623f
C8160 XA.Cn[9].n11 VGND 0.09378f
C8161 XA.Cn[9].t17 VGND 0.01164f
C8162 XA.Cn[9].t35 VGND 0.01272f
C8163 XA.Cn[9].n12 VGND 0.0284f
C8164 XA.Cn[9].n13 VGND 0.01623f
C8165 XA.Cn[9].n14 VGND 0.09378f
C8166 XA.Cn[9].t39 VGND 0.01164f
C8167 XA.Cn[9].t24 VGND 0.01272f
C8168 XA.Cn[9].n15 VGND 0.0284f
C8169 XA.Cn[9].n16 VGND 0.01623f
C8170 XA.Cn[9].n17 VGND 0.09378f
C8171 XA.Cn[9].t40 VGND 0.01164f
C8172 XA.Cn[9].t25 VGND 0.01272f
C8173 XA.Cn[9].n18 VGND 0.0284f
C8174 XA.Cn[9].n19 VGND 0.01623f
C8175 XA.Cn[9].n20 VGND 0.09378f
C8176 XA.Cn[9].t22 VGND 0.01164f
C8177 XA.Cn[9].t38 VGND 0.01272f
C8178 XA.Cn[9].n21 VGND 0.0284f
C8179 XA.Cn[9].n22 VGND 0.01623f
C8180 XA.Cn[9].n23 VGND 0.09378f
C8181 XA.Cn[9].t28 VGND 0.01164f
C8182 XA.Cn[9].t14 VGND 0.01272f
C8183 XA.Cn[9].n24 VGND 0.0284f
C8184 XA.Cn[9].n25 VGND 0.01623f
C8185 XA.Cn[9].n26 VGND 0.09378f
C8186 XA.Cn[9].t31 VGND 0.01164f
C8187 XA.Cn[9].t16 VGND 0.01272f
C8188 XA.Cn[9].n27 VGND 0.0284f
C8189 XA.Cn[9].n28 VGND 0.01623f
C8190 XA.Cn[9].n29 VGND 0.09378f
C8191 XA.Cn[9].t19 VGND 0.01164f
C8192 XA.Cn[9].t36 VGND 0.01272f
C8193 XA.Cn[9].n30 VGND 0.0284f
C8194 XA.Cn[9].n31 VGND 0.01623f
C8195 XA.Cn[9].n32 VGND 0.09378f
C8196 XA.Cn[9].t21 VGND 0.01164f
C8197 XA.Cn[9].t37 VGND 0.01272f
C8198 XA.Cn[9].n33 VGND 0.0284f
C8199 XA.Cn[9].n34 VGND 0.01623f
C8200 XA.Cn[9].n35 VGND 0.09378f
C8201 XA.Cn[9].t32 VGND 0.01164f
C8202 XA.Cn[9].t18 VGND 0.01272f
C8203 XA.Cn[9].n36 VGND 0.0284f
C8204 XA.Cn[9].n37 VGND 0.01623f
C8205 XA.Cn[9].n38 VGND 0.09378f
C8206 XA.Cn[9].t42 VGND 0.01164f
C8207 XA.Cn[9].t27 VGND 0.01272f
C8208 XA.Cn[9].n39 VGND 0.0284f
C8209 XA.Cn[9].n40 VGND 0.01623f
C8210 XA.Cn[9].n41 VGND 0.09378f
C8211 XA.Cn[9].t43 VGND 0.01164f
C8212 XA.Cn[9].t29 VGND 0.01272f
C8213 XA.Cn[9].n42 VGND 0.0284f
C8214 XA.Cn[9].n43 VGND 0.01623f
C8215 XA.Cn[9].n44 VGND 0.09378f
C8216 XA.Cn[9].t23 VGND 0.01164f
C8217 XA.Cn[9].t41 VGND 0.01272f
C8218 XA.Cn[9].n45 VGND 0.0284f
C8219 XA.Cn[9].n46 VGND 0.01623f
C8220 XA.Cn[9].n47 VGND 0.09378f
C8221 XA.Cn[9].t33 VGND 0.01164f
C8222 XA.Cn[9].t20 VGND 0.01272f
C8223 XA.Cn[9].n48 VGND 0.0284f
C8224 XA.Cn[9].n49 VGND 0.01623f
C8225 XA.Cn[9].n50 VGND 0.09378f
C8226 XA.Cn[9].n51 VGND 0.04286f
C8227 XA.Cn[9].t4 VGND 0.01469f
C8228 XA.Cn[9].t7 VGND 0.01469f
C8229 XA.Cn[9].n52 VGND 0.03174f
C8230 XA.Cn[9].t6 VGND 0.01469f
C8231 XA.Cn[9].t5 VGND 0.01469f
C8232 XA.Cn[9].n53 VGND 0.05003f
C8233 XA.Cn[9].n54 VGND 0.1325f
C8234 XA.Cn[9].t1 VGND 0.01469f
C8235 XA.Cn[9].t0 VGND 0.01469f
C8236 XA.Cn[9].n56 VGND 0.0446f
C8237 XA.Cn[9].t3 VGND 0.01469f
C8238 XA.Cn[9].t2 VGND 0.01469f
C8239 XA.Cn[9].n57 VGND 0.03266f
C8240 XA.Cn[9].n58 VGND 0.14534f
C8241 XA.Cn[5].t7 VGND 0.0121f
C8242 XA.Cn[5].t6 VGND 0.0121f
C8243 XA.Cn[5].n0 VGND 0.02443f
C8244 XA.Cn[5].t5 VGND 0.0121f
C8245 XA.Cn[5].t4 VGND 0.0121f
C8246 XA.Cn[5].n1 VGND 0.02858f
C8247 XA.Cn[5].n2 VGND 0.08573f
C8248 XA.Cn[5].n3 VGND 0.01791f
C8249 XA.Cn[5].n4 VGND 0.01791f
C8250 XA.Cn[5].n5 VGND 0.01791f
C8251 XA.Cn[5].n6 VGND 0.02985f
C8252 XA.Cn[5].n7 VGND 0.0853f
C8253 XA.Cn[5].n8 VGND 0.05273f
C8254 XA.Cn[5].n9 VGND 0.05951f
C8255 XA.Cn[5].t33 VGND 0.01048f
C8256 XA.Cn[5].n10 VGND 0.0234f
C8257 XA.Cn[5].n11 VGND 0.01337f
C8258 XA.Cn[5].n12 VGND 0.01626f
C8259 XA.Cn[5].t19 VGND 0.01048f
C8260 XA.Cn[5].n13 VGND 0.0234f
C8261 XA.Cn[5].n14 VGND 0.01337f
C8262 XA.Cn[5].n15 VGND 0.07725f
C8263 XA.Cn[5].t23 VGND 0.01048f
C8264 XA.Cn[5].n16 VGND 0.0234f
C8265 XA.Cn[5].n17 VGND 0.01337f
C8266 XA.Cn[5].n18 VGND 0.07725f
C8267 XA.Cn[5].t24 VGND 0.01048f
C8268 XA.Cn[5].n19 VGND 0.0234f
C8269 XA.Cn[5].n20 VGND 0.01337f
C8270 XA.Cn[5].n21 VGND 0.07725f
C8271 XA.Cn[5].t13 VGND 0.01048f
C8272 XA.Cn[5].n22 VGND 0.0234f
C8273 XA.Cn[5].n23 VGND 0.01337f
C8274 XA.Cn[5].n24 VGND 0.07725f
C8275 XA.Cn[5].t14 VGND 0.01048f
C8276 XA.Cn[5].n25 VGND 0.0234f
C8277 XA.Cn[5].n26 VGND 0.01337f
C8278 XA.Cn[5].n27 VGND 0.07725f
C8279 XA.Cn[5].t27 VGND 0.01048f
C8280 XA.Cn[5].n28 VGND 0.0234f
C8281 XA.Cn[5].n29 VGND 0.01337f
C8282 XA.Cn[5].n30 VGND 0.07725f
C8283 XA.Cn[5].t35 VGND 0.01048f
C8284 XA.Cn[5].n31 VGND 0.0234f
C8285 XA.Cn[5].n32 VGND 0.01337f
C8286 XA.Cn[5].n33 VGND 0.07725f
C8287 XA.Cn[5].t37 VGND 0.01048f
C8288 XA.Cn[5].n34 VGND 0.0234f
C8289 XA.Cn[5].n35 VGND 0.01337f
C8290 XA.Cn[5].n36 VGND 0.07725f
C8291 XA.Cn[5].t25 VGND 0.01048f
C8292 XA.Cn[5].n37 VGND 0.0234f
C8293 XA.Cn[5].n38 VGND 0.01337f
C8294 XA.Cn[5].n39 VGND 0.07725f
C8295 XA.Cn[5].t26 VGND 0.01048f
C8296 XA.Cn[5].n40 VGND 0.0234f
C8297 XA.Cn[5].n41 VGND 0.01337f
C8298 XA.Cn[5].n42 VGND 0.07725f
C8299 XA.Cn[5].t39 VGND 0.01048f
C8300 XA.Cn[5].n43 VGND 0.0234f
C8301 XA.Cn[5].n44 VGND 0.01337f
C8302 XA.Cn[5].n45 VGND 0.07725f
C8303 XA.Cn[5].t16 VGND 0.01048f
C8304 XA.Cn[5].n46 VGND 0.0234f
C8305 XA.Cn[5].n47 VGND 0.01337f
C8306 XA.Cn[5].n48 VGND 0.07725f
C8307 XA.Cn[5].t18 VGND 0.01048f
C8308 XA.Cn[5].n49 VGND 0.0234f
C8309 XA.Cn[5].n50 VGND 0.01337f
C8310 XA.Cn[5].n51 VGND 0.07725f
C8311 XA.Cn[5].t30 VGND 0.01048f
C8312 XA.Cn[5].n52 VGND 0.0234f
C8313 XA.Cn[5].n53 VGND 0.01337f
C8314 XA.Cn[5].n54 VGND 0.07725f
C8315 XA.Cn[5].t41 VGND 0.01048f
C8316 XA.Cn[5].n55 VGND 0.0234f
C8317 XA.Cn[5].n56 VGND 0.01337f
C8318 XA.Cn[5].n57 VGND 0.07725f
C8319 XA.Cn[5].n58 VGND 0.2186f
C8320 XA.Cn[5].n59 VGND 0.04035f
C8321 XThR.Tn[9].t0 VGND 0.01255f
C8322 XThR.Tn[9].t2 VGND 0.01255f
C8323 XThR.Tn[9].n0 VGND 0.0251f
C8324 XThR.Tn[9].t1 VGND 0.01255f
C8325 XThR.Tn[9].t3 VGND 0.01255f
C8326 XThR.Tn[9].n1 VGND 0.03131f
C8327 XThR.Tn[9].n2 VGND 0.06315f
C8328 XThR.Tn[9].t10 VGND 0.01931f
C8329 XThR.Tn[9].t8 VGND 0.01931f
C8330 XThR.Tn[9].n3 VGND 0.05863f
C8331 XThR.Tn[9].t11 VGND 0.01931f
C8332 XThR.Tn[9].t9 VGND 0.01931f
C8333 XThR.Tn[9].n4 VGND 0.04293f
C8334 XThR.Tn[9].n5 VGND 0.19519f
C8335 XThR.Tn[9].t6 VGND 0.01931f
C8336 XThR.Tn[9].t4 VGND 0.01931f
C8337 XThR.Tn[9].n6 VGND 0.04172f
C8338 XThR.Tn[9].t7 VGND 0.01931f
C8339 XThR.Tn[9].t5 VGND 0.01931f
C8340 XThR.Tn[9].n7 VGND 0.0635f
C8341 XThR.Tn[9].n8 VGND 0.17633f
C8342 XThR.Tn[9].n9 VGND 0.02361f
C8343 XThR.Tn[9].t17 VGND 0.01509f
C8344 XThR.Tn[9].t71 VGND 0.01653f
C8345 XThR.Tn[9].n10 VGND 0.04036f
C8346 XThR.Tn[9].n11 VGND 0.07752f
C8347 XThR.Tn[9].t35 VGND 0.01509f
C8348 XThR.Tn[9].t28 VGND 0.01653f
C8349 XThR.Tn[9].n12 VGND 0.04036f
C8350 XThR.Tn[9].t50 VGND 0.01504f
C8351 XThR.Tn[9].t19 VGND 0.01647f
C8352 XThR.Tn[9].n13 VGND 0.04199f
C8353 XThR.Tn[9].n14 VGND 0.0295f
C8354 XThR.Tn[9].n16 VGND 0.09466f
C8355 XThR.Tn[9].t72 VGND 0.01509f
C8356 XThR.Tn[9].t64 VGND 0.01653f
C8357 XThR.Tn[9].n17 VGND 0.04036f
C8358 XThR.Tn[9].t26 VGND 0.01504f
C8359 XThR.Tn[9].t59 VGND 0.01647f
C8360 XThR.Tn[9].n18 VGND 0.04199f
C8361 XThR.Tn[9].n19 VGND 0.0295f
C8362 XThR.Tn[9].n21 VGND 0.09466f
C8363 XThR.Tn[9].t29 VGND 0.01509f
C8364 XThR.Tn[9].t21 VGND 0.01653f
C8365 XThR.Tn[9].n22 VGND 0.04036f
C8366 XThR.Tn[9].t41 VGND 0.01504f
C8367 XThR.Tn[9].t15 VGND 0.01647f
C8368 XThR.Tn[9].n23 VGND 0.04199f
C8369 XThR.Tn[9].n24 VGND 0.0295f
C8370 XThR.Tn[9].n26 VGND 0.09466f
C8371 XThR.Tn[9].t56 VGND 0.01509f
C8372 XThR.Tn[9].t46 VGND 0.01653f
C8373 XThR.Tn[9].n27 VGND 0.04036f
C8374 XThR.Tn[9].t73 VGND 0.01504f
C8375 XThR.Tn[9].t42 VGND 0.01647f
C8376 XThR.Tn[9].n28 VGND 0.04199f
C8377 XThR.Tn[9].n29 VGND 0.0295f
C8378 XThR.Tn[9].n31 VGND 0.09466f
C8379 XThR.Tn[9].t31 VGND 0.01509f
C8380 XThR.Tn[9].t23 VGND 0.01653f
C8381 XThR.Tn[9].n32 VGND 0.04036f
C8382 XThR.Tn[9].t44 VGND 0.01504f
C8383 XThR.Tn[9].t16 VGND 0.01647f
C8384 XThR.Tn[9].n33 VGND 0.04199f
C8385 XThR.Tn[9].n34 VGND 0.0295f
C8386 XThR.Tn[9].n36 VGND 0.09466f
C8387 XThR.Tn[9].t67 VGND 0.01509f
C8388 XThR.Tn[9].t37 VGND 0.01653f
C8389 XThR.Tn[9].n37 VGND 0.04036f
C8390 XThR.Tn[9].t20 VGND 0.01504f
C8391 XThR.Tn[9].t33 VGND 0.01647f
C8392 XThR.Tn[9].n38 VGND 0.04199f
C8393 XThR.Tn[9].n39 VGND 0.0295f
C8394 XThR.Tn[9].n41 VGND 0.09466f
C8395 XThR.Tn[9].t36 VGND 0.01509f
C8396 XThR.Tn[9].t32 VGND 0.01653f
C8397 XThR.Tn[9].n42 VGND 0.04036f
C8398 XThR.Tn[9].t51 VGND 0.01504f
C8399 XThR.Tn[9].t25 VGND 0.01647f
C8400 XThR.Tn[9].n43 VGND 0.04199f
C8401 XThR.Tn[9].n44 VGND 0.0295f
C8402 XThR.Tn[9].n46 VGND 0.09466f
C8403 XThR.Tn[9].t39 VGND 0.01509f
C8404 XThR.Tn[9].t45 VGND 0.01653f
C8405 XThR.Tn[9].n47 VGND 0.04036f
C8406 XThR.Tn[9].t55 VGND 0.01504f
C8407 XThR.Tn[9].t40 VGND 0.01647f
C8408 XThR.Tn[9].n48 VGND 0.04199f
C8409 XThR.Tn[9].n49 VGND 0.0295f
C8410 XThR.Tn[9].n51 VGND 0.09466f
C8411 XThR.Tn[9].t58 VGND 0.01509f
C8412 XThR.Tn[9].t66 VGND 0.01653f
C8413 XThR.Tn[9].n52 VGND 0.04036f
C8414 XThR.Tn[9].t13 VGND 0.01504f
C8415 XThR.Tn[9].t60 VGND 0.01647f
C8416 XThR.Tn[9].n53 VGND 0.04199f
C8417 XThR.Tn[9].n54 VGND 0.0295f
C8418 XThR.Tn[9].n56 VGND 0.09466f
C8419 XThR.Tn[9].t48 VGND 0.01509f
C8420 XThR.Tn[9].t24 VGND 0.01653f
C8421 XThR.Tn[9].n57 VGND 0.04036f
C8422 XThR.Tn[9].t65 VGND 0.01504f
C8423 XThR.Tn[9].t18 VGND 0.01647f
C8424 XThR.Tn[9].n58 VGND 0.04199f
C8425 XThR.Tn[9].n59 VGND 0.0295f
C8426 XThR.Tn[9].n61 VGND 0.09466f
C8427 XThR.Tn[9].t70 VGND 0.01509f
C8428 XThR.Tn[9].t62 VGND 0.01653f
C8429 XThR.Tn[9].n62 VGND 0.04036f
C8430 XThR.Tn[9].t22 VGND 0.01504f
C8431 XThR.Tn[9].t52 VGND 0.01647f
C8432 XThR.Tn[9].n63 VGND 0.04199f
C8433 XThR.Tn[9].n64 VGND 0.0295f
C8434 XThR.Tn[9].n66 VGND 0.09466f
C8435 XThR.Tn[9].t38 VGND 0.01509f
C8436 XThR.Tn[9].t34 VGND 0.01653f
C8437 XThR.Tn[9].n67 VGND 0.04036f
C8438 XThR.Tn[9].t53 VGND 0.01504f
C8439 XThR.Tn[9].t27 VGND 0.01647f
C8440 XThR.Tn[9].n68 VGND 0.04199f
C8441 XThR.Tn[9].n69 VGND 0.0295f
C8442 XThR.Tn[9].n71 VGND 0.09466f
C8443 XThR.Tn[9].t57 VGND 0.01509f
C8444 XThR.Tn[9].t47 VGND 0.01653f
C8445 XThR.Tn[9].n72 VGND 0.04036f
C8446 XThR.Tn[9].t12 VGND 0.01504f
C8447 XThR.Tn[9].t43 VGND 0.01647f
C8448 XThR.Tn[9].n73 VGND 0.04199f
C8449 XThR.Tn[9].n74 VGND 0.0295f
C8450 XThR.Tn[9].n76 VGND 0.09466f
C8451 XThR.Tn[9].t14 VGND 0.01509f
C8452 XThR.Tn[9].t69 VGND 0.01653f
C8453 XThR.Tn[9].n77 VGND 0.04036f
C8454 XThR.Tn[9].t30 VGND 0.01504f
C8455 XThR.Tn[9].t61 VGND 0.01647f
C8456 XThR.Tn[9].n78 VGND 0.04199f
C8457 XThR.Tn[9].n79 VGND 0.0295f
C8458 XThR.Tn[9].n81 VGND 0.09466f
C8459 XThR.Tn[9].t49 VGND 0.01509f
C8460 XThR.Tn[9].t63 VGND 0.01653f
C8461 XThR.Tn[9].n82 VGND 0.04036f
C8462 XThR.Tn[9].t68 VGND 0.01504f
C8463 XThR.Tn[9].t54 VGND 0.01647f
C8464 XThR.Tn[9].n83 VGND 0.04199f
C8465 XThR.Tn[9].n84 VGND 0.0295f
C8466 XThR.Tn[9].n86 VGND 0.09466f
C8467 XThR.Tn[9].n87 VGND 0.08603f
C8468 XThR.Tn[9].n88 VGND 0.27907f
C8469 XA.Cn[6].n0 VGND 0.0301f
C8470 XA.Cn[6].n1 VGND 0.01807f
C8471 XA.Cn[6].n2 VGND 0.08604f
C8472 XA.Cn[6].n3 VGND 0.01807f
C8473 XA.Cn[6].n4 VGND 0.05319f
C8474 XA.Cn[6].n5 VGND 0.01807f
C8475 XA.Cn[6].n6 VGND 0.06003f
C8476 XA.Cn[6].t26 VGND 0.01057f
C8477 XA.Cn[6].n7 VGND 0.0236f
C8478 XA.Cn[6].n8 VGND 0.01349f
C8479 XA.Cn[6].n9 VGND 0.0164f
C8480 XA.Cn[6].t13 VGND 0.01057f
C8481 XA.Cn[6].n10 VGND 0.0236f
C8482 XA.Cn[6].n11 VGND 0.01349f
C8483 XA.Cn[6].n12 VGND 0.07792f
C8484 XA.Cn[6].t17 VGND 0.01057f
C8485 XA.Cn[6].n13 VGND 0.0236f
C8486 XA.Cn[6].n14 VGND 0.01349f
C8487 XA.Cn[6].n15 VGND 0.07792f
C8488 XA.Cn[6].t18 VGND 0.01057f
C8489 XA.Cn[6].n16 VGND 0.0236f
C8490 XA.Cn[6].n17 VGND 0.01349f
C8491 XA.Cn[6].n18 VGND 0.07792f
C8492 XA.Cn[6].t37 VGND 0.01057f
C8493 XA.Cn[6].n19 VGND 0.0236f
C8494 XA.Cn[6].n20 VGND 0.01349f
C8495 XA.Cn[6].n21 VGND 0.07792f
C8496 XA.Cn[6].t38 VGND 0.01057f
C8497 XA.Cn[6].n22 VGND 0.0236f
C8498 XA.Cn[6].n23 VGND 0.01349f
C8499 XA.Cn[6].n24 VGND 0.07792f
C8500 XA.Cn[6].t22 VGND 0.01057f
C8501 XA.Cn[6].n25 VGND 0.0236f
C8502 XA.Cn[6].n26 VGND 0.01349f
C8503 XA.Cn[6].n27 VGND 0.07792f
C8504 XA.Cn[6].t29 VGND 0.01057f
C8505 XA.Cn[6].n28 VGND 0.0236f
C8506 XA.Cn[6].n29 VGND 0.01349f
C8507 XA.Cn[6].n30 VGND 0.07792f
C8508 XA.Cn[6].t31 VGND 0.01057f
C8509 XA.Cn[6].n31 VGND 0.0236f
C8510 XA.Cn[6].n32 VGND 0.01349f
C8511 XA.Cn[6].n33 VGND 0.07792f
C8512 XA.Cn[6].t19 VGND 0.01057f
C8513 XA.Cn[6].n34 VGND 0.0236f
C8514 XA.Cn[6].n35 VGND 0.01349f
C8515 XA.Cn[6].n36 VGND 0.07792f
C8516 XA.Cn[6].t21 VGND 0.01057f
C8517 XA.Cn[6].n37 VGND 0.0236f
C8518 XA.Cn[6].n38 VGND 0.01349f
C8519 XA.Cn[6].n39 VGND 0.07792f
C8520 XA.Cn[6].t32 VGND 0.01057f
C8521 XA.Cn[6].n40 VGND 0.0236f
C8522 XA.Cn[6].n41 VGND 0.01349f
C8523 XA.Cn[6].n42 VGND 0.07792f
C8524 XA.Cn[6].t41 VGND 0.01057f
C8525 XA.Cn[6].n43 VGND 0.0236f
C8526 XA.Cn[6].n44 VGND 0.01349f
C8527 XA.Cn[6].n45 VGND 0.07792f
C8528 XA.Cn[6].t43 VGND 0.01057f
C8529 XA.Cn[6].n46 VGND 0.0236f
C8530 XA.Cn[6].n47 VGND 0.01349f
C8531 XA.Cn[6].n48 VGND 0.07792f
C8532 XA.Cn[6].t24 VGND 0.01057f
C8533 XA.Cn[6].n49 VGND 0.0236f
C8534 XA.Cn[6].n50 VGND 0.01349f
C8535 XA.Cn[6].n51 VGND 0.07792f
C8536 XA.Cn[6].t34 VGND 0.01057f
C8537 XA.Cn[6].n52 VGND 0.0236f
C8538 XA.Cn[6].n53 VGND 0.01349f
C8539 XA.Cn[6].n54 VGND 0.07792f
C8540 XA.Cn[6].n55 VGND 0.20284f
C8541 XA.Cn[6].n56 VGND 0.04609f
C8542 XA.Cn[6].t1 VGND 0.01221f
C8543 XA.Cn[6].t0 VGND 0.01221f
C8544 XA.Cn[6].n57 VGND 0.02883f
C8545 XA.Cn[6].t3 VGND 0.01221f
C8546 XA.Cn[6].t2 VGND 0.01221f
C8547 XA.Cn[6].n58 VGND 0.02464f
C8548 XA.Cn[6].n59 VGND 0.0807f
C8549 XA.Cn[6].n60 VGND 0.02554f
C8550 thermo15c_0.XTBN.Y.n0 VGND 0.01531f
C8551 thermo15c_0.XTBN.Y.t50 VGND 0.01024f
C8552 thermo15c_0.XTBN.Y.t18 VGND 0.01024f
C8553 thermo15c_0.XTBN.Y.n1 VGND 0.01477f
C8554 thermo15c_0.XTBN.Y.t120 VGND 0.01024f
C8555 thermo15c_0.XTBN.Y.t114 VGND 0.01024f
C8556 thermo15c_0.XTBN.Y.n3 VGND 0.0138f
C8557 thermo15c_0.XTBN.Y.n5 VGND 0.01477f
C8558 thermo15c_0.XTBN.Y.n10 VGND 0.02164f
C8559 thermo15c_0.XTBN.Y.t79 VGND 0.01024f
C8560 thermo15c_0.XTBN.Y.t36 VGND 0.01024f
C8561 thermo15c_0.XTBN.Y.n13 VGND 0.01477f
C8562 thermo15c_0.XTBN.Y.t26 VGND 0.01024f
C8563 thermo15c_0.XTBN.Y.t21 VGND 0.01024f
C8564 thermo15c_0.XTBN.Y.n15 VGND 0.0138f
C8565 thermo15c_0.XTBN.Y.n17 VGND 0.01477f
C8566 thermo15c_0.XTBN.Y.n22 VGND 0.02164f
C8567 thermo15c_0.XTBN.Y.n25 VGND 0.11789f
C8568 thermo15c_0.XTBN.Y.t106 VGND 0.01024f
C8569 thermo15c_0.XTBN.Y.t70 VGND 0.01024f
C8570 thermo15c_0.XTBN.Y.n26 VGND 0.01477f
C8571 thermo15c_0.XTBN.Y.t56 VGND 0.01024f
C8572 thermo15c_0.XTBN.Y.t48 VGND 0.01024f
C8573 thermo15c_0.XTBN.Y.n28 VGND 0.0138f
C8574 thermo15c_0.XTBN.Y.n30 VGND 0.01477f
C8575 thermo15c_0.XTBN.Y.n35 VGND 0.02164f
C8576 thermo15c_0.XTBN.Y.n38 VGND 0.07443f
C8577 thermo15c_0.XTBN.Y.t39 VGND 0.01024f
C8578 thermo15c_0.XTBN.Y.t122 VGND 0.01024f
C8579 thermo15c_0.XTBN.Y.n39 VGND 0.01477f
C8580 thermo15c_0.XTBN.Y.t109 VGND 0.01024f
C8581 thermo15c_0.XTBN.Y.t102 VGND 0.01024f
C8582 thermo15c_0.XTBN.Y.n41 VGND 0.0138f
C8583 thermo15c_0.XTBN.Y.n43 VGND 0.01477f
C8584 thermo15c_0.XTBN.Y.n48 VGND 0.02164f
C8585 thermo15c_0.XTBN.Y.n51 VGND 0.07443f
C8586 thermo15c_0.XTBN.Y.t47 VGND 0.01024f
C8587 thermo15c_0.XTBN.Y.t17 VGND 0.01024f
C8588 thermo15c_0.XTBN.Y.n52 VGND 0.01477f
C8589 thermo15c_0.XTBN.Y.t116 VGND 0.01024f
C8590 thermo15c_0.XTBN.Y.t111 VGND 0.01024f
C8591 thermo15c_0.XTBN.Y.n54 VGND 0.0138f
C8592 thermo15c_0.XTBN.Y.n56 VGND 0.01477f
C8593 thermo15c_0.XTBN.Y.n61 VGND 0.02164f
C8594 thermo15c_0.XTBN.Y.n64 VGND 0.07443f
C8595 thermo15c_0.XTBN.Y.t101 VGND 0.01024f
C8596 thermo15c_0.XTBN.Y.t63 VGND 0.01024f
C8597 thermo15c_0.XTBN.Y.n65 VGND 0.01477f
C8598 thermo15c_0.XTBN.Y.t52 VGND 0.01024f
C8599 thermo15c_0.XTBN.Y.t44 VGND 0.01024f
C8600 thermo15c_0.XTBN.Y.n67 VGND 0.0138f
C8601 thermo15c_0.XTBN.Y.n69 VGND 0.01477f
C8602 thermo15c_0.XTBN.Y.n74 VGND 0.02164f
C8603 thermo15c_0.XTBN.Y.n77 VGND 0.07443f
C8604 thermo15c_0.XTBN.Y.t25 VGND 0.01024f
C8605 thermo15c_0.XTBN.Y.t100 VGND 0.01024f
C8606 thermo15c_0.XTBN.Y.n78 VGND 0.01477f
C8607 thermo15c_0.XTBN.Y.t93 VGND 0.01024f
C8608 thermo15c_0.XTBN.Y.t90 VGND 0.01024f
C8609 thermo15c_0.XTBN.Y.n80 VGND 0.0138f
C8610 thermo15c_0.XTBN.Y.n82 VGND 0.01477f
C8611 thermo15c_0.XTBN.Y.n87 VGND 0.02164f
C8612 thermo15c_0.XTBN.Y.n90 VGND 0.06646f
C8613 thermo15c_0.XTBN.Y.t46 VGND 0.01024f
C8614 thermo15c_0.XTBN.Y.t6 VGND 0.01024f
C8615 thermo15c_0.XTBN.Y.n92 VGND 0.01243f
C8616 thermo15c_0.XTBN.Y.t12 VGND 0.01024f
C8617 thermo15c_0.XTBN.Y.n93 VGND 0.01348f
C8618 thermo15c_0.XTBN.Y.n95 VGND 0.01252f
C8619 thermo15c_0.XTBN.Y.n98 VGND 0.01348f
C8620 thermo15c_0.XTBN.Y.t54 VGND 0.01024f
C8621 thermo15c_0.XTBN.Y.n99 VGND 0.01227f
C8622 thermo15c_0.XTBN.Y.n101 VGND 0.01009f
C8623 thermo15c_0.XTBN.Y.t38 VGND 0.01024f
C8624 thermo15c_0.XTBN.Y.t113 VGND 0.01024f
C8625 thermo15c_0.XTBN.Y.n103 VGND 0.01243f
C8626 thermo15c_0.XTBN.Y.t119 VGND 0.01024f
C8627 thermo15c_0.XTBN.Y.n104 VGND 0.01348f
C8628 thermo15c_0.XTBN.Y.n106 VGND 0.01252f
C8629 thermo15c_0.XTBN.Y.n109 VGND 0.01348f
C8630 thermo15c_0.XTBN.Y.t42 VGND 0.01024f
C8631 thermo15c_0.XTBN.Y.n110 VGND 0.01227f
C8632 thermo15c_0.XTBN.Y.n113 VGND 0.11256f
C8633 thermo15c_0.XTBN.Y.t30 VGND 0.01024f
C8634 thermo15c_0.XTBN.Y.t98 VGND 0.01024f
C8635 thermo15c_0.XTBN.Y.n115 VGND 0.01243f
C8636 thermo15c_0.XTBN.Y.t103 VGND 0.01024f
C8637 thermo15c_0.XTBN.Y.n116 VGND 0.01348f
C8638 thermo15c_0.XTBN.Y.n118 VGND 0.01252f
C8639 thermo15c_0.XTBN.Y.n121 VGND 0.01348f
C8640 thermo15c_0.XTBN.Y.t34 VGND 0.01024f
C8641 thermo15c_0.XTBN.Y.n122 VGND 0.01227f
C8642 thermo15c_0.XTBN.Y.n125 VGND 0.07521f
C8643 thermo15c_0.XTBN.Y.t96 VGND 0.01024f
C8644 thermo15c_0.XTBN.Y.t51 VGND 0.01024f
C8645 thermo15c_0.XTBN.Y.n127 VGND 0.01243f
C8646 thermo15c_0.XTBN.Y.t58 VGND 0.01024f
C8647 thermo15c_0.XTBN.Y.n128 VGND 0.01348f
C8648 thermo15c_0.XTBN.Y.n130 VGND 0.01252f
C8649 thermo15c_0.XTBN.Y.n133 VGND 0.01348f
C8650 thermo15c_0.XTBN.Y.t99 VGND 0.01024f
C8651 thermo15c_0.XTBN.Y.n134 VGND 0.01227f
C8652 thermo15c_0.XTBN.Y.n137 VGND 0.07521f
C8653 thermo15c_0.XTBN.Y.t88 VGND 0.01024f
C8654 thermo15c_0.XTBN.Y.t37 VGND 0.01024f
C8655 thermo15c_0.XTBN.Y.n139 VGND 0.01243f
C8656 thermo15c_0.XTBN.Y.t40 VGND 0.01024f
C8657 thermo15c_0.XTBN.Y.n140 VGND 0.01348f
C8658 thermo15c_0.XTBN.Y.n142 VGND 0.01252f
C8659 thermo15c_0.XTBN.Y.n145 VGND 0.01348f
C8660 thermo15c_0.XTBN.Y.t91 VGND 0.01024f
C8661 thermo15c_0.XTBN.Y.n146 VGND 0.01227f
C8662 thermo15c_0.XTBN.Y.n149 VGND 0.07534f
C8663 thermo15c_0.XTBN.Y.t7 VGND 0.01024f
C8664 thermo15c_0.XTBN.Y.t81 VGND 0.01024f
C8665 thermo15c_0.XTBN.Y.n151 VGND 0.01243f
C8666 thermo15c_0.XTBN.Y.t86 VGND 0.01024f
C8667 thermo15c_0.XTBN.Y.n152 VGND 0.01348f
C8668 thermo15c_0.XTBN.Y.n154 VGND 0.01252f
C8669 thermo15c_0.XTBN.Y.n157 VGND 0.01348f
C8670 thermo15c_0.XTBN.Y.t13 VGND 0.01024f
C8671 thermo15c_0.XTBN.Y.n158 VGND 0.01227f
C8672 thermo15c_0.XTBN.Y.n161 VGND 0.07521f
C8673 thermo15c_0.XTBN.Y.t23 VGND 0.01024f
C8674 thermo15c_0.XTBN.Y.t95 VGND 0.01024f
C8675 thermo15c_0.XTBN.Y.n163 VGND 0.01243f
C8676 thermo15c_0.XTBN.Y.t97 VGND 0.01024f
C8677 thermo15c_0.XTBN.Y.n164 VGND 0.01348f
C8678 thermo15c_0.XTBN.Y.n166 VGND 0.01252f
C8679 thermo15c_0.XTBN.Y.n169 VGND 0.01348f
C8680 thermo15c_0.XTBN.Y.t28 VGND 0.01024f
C8681 thermo15c_0.XTBN.Y.n170 VGND 0.01227f
C8682 thermo15c_0.XTBN.Y.n173 VGND 0.08751f
C8683 thermo15c_0.XTBN.Y.n174 VGND 0.11019f
C8684 thermo15c_0.XTBN.Y.t75 VGND 0.01024f
C8685 thermo15c_0.XTBN.Y.t33 VGND 0.01024f
C8686 thermo15c_0.XTBN.Y.n175 VGND 0.01477f
C8687 thermo15c_0.XTBN.Y.t27 VGND 0.01024f
C8688 thermo15c_0.XTBN.Y.n176 VGND 0.02293f
C8689 thermo15c_0.XTBN.Y.n181 VGND 0.01477f
C8690 thermo15c_0.XTBN.Y.t9 VGND 0.01024f
C8691 thermo15c_0.XTBN.Y.n182 VGND 0.0138f
C8692 thermo15c_0.XTBN.Y.n186 VGND 0.11129f
C8693 thermo15c_0.XTBN.Y.n187 VGND 0.02169f
C8694 thermo15c_0.XTBN.Y.n191 VGND 0.01513f
C8695 thermo15c_0.XTBN.Y.n192 VGND 0.0307f
C8696 XThR.Tn[12].t11 VGND 0.01931f
C8697 XThR.Tn[12].t9 VGND 0.01931f
C8698 XThR.Tn[12].n0 VGND 0.05864f
C8699 XThR.Tn[12].t8 VGND 0.01931f
C8700 XThR.Tn[12].t10 VGND 0.01931f
C8701 XThR.Tn[12].n1 VGND 0.04293f
C8702 XThR.Tn[12].n2 VGND 0.1952f
C8703 XThR.Tn[12].t6 VGND 0.01931f
C8704 XThR.Tn[12].t4 VGND 0.01931f
C8705 XThR.Tn[12].n3 VGND 0.04172f
C8706 XThR.Tn[12].t7 VGND 0.01931f
C8707 XThR.Tn[12].t5 VGND 0.01931f
C8708 XThR.Tn[12].n4 VGND 0.06351f
C8709 XThR.Tn[12].n5 VGND 0.17633f
C8710 XThR.Tn[12].t36 VGND 0.01509f
C8711 XThR.Tn[12].t28 VGND 0.01653f
C8712 XThR.Tn[12].n7 VGND 0.04036f
C8713 XThR.Tn[12].n8 VGND 0.07753f
C8714 XThR.Tn[12].t53 VGND 0.01509f
C8715 XThR.Tn[12].t43 VGND 0.01653f
C8716 XThR.Tn[12].n9 VGND 0.04036f
C8717 XThR.Tn[12].t71 VGND 0.01504f
C8718 XThR.Tn[12].t21 VGND 0.01647f
C8719 XThR.Tn[12].n10 VGND 0.04199f
C8720 XThR.Tn[12].n11 VGND 0.0295f
C8721 XThR.Tn[12].n13 VGND 0.09466f
C8722 XThR.Tn[12].t30 VGND 0.01509f
C8723 XThR.Tn[12].t20 VGND 0.01653f
C8724 XThR.Tn[12].n14 VGND 0.04036f
C8725 XThR.Tn[12].t49 VGND 0.01504f
C8726 XThR.Tn[12].t60 VGND 0.01647f
C8727 XThR.Tn[12].n15 VGND 0.04199f
C8728 XThR.Tn[12].n16 VGND 0.0295f
C8729 XThR.Tn[12].n18 VGND 0.09466f
C8730 XThR.Tn[12].t45 VGND 0.01509f
C8731 XThR.Tn[12].t38 VGND 0.01653f
C8732 XThR.Tn[12].n19 VGND 0.04036f
C8733 XThR.Tn[12].t63 VGND 0.01504f
C8734 XThR.Tn[12].t15 VGND 0.01647f
C8735 XThR.Tn[12].n20 VGND 0.04199f
C8736 XThR.Tn[12].n21 VGND 0.0295f
C8737 XThR.Tn[12].n23 VGND 0.09466f
C8738 XThR.Tn[12].t70 VGND 0.01509f
C8739 XThR.Tn[12].t66 VGND 0.01653f
C8740 XThR.Tn[12].n24 VGND 0.04036f
C8741 XThR.Tn[12].t33 VGND 0.01504f
C8742 XThR.Tn[12].t46 VGND 0.01647f
C8743 XThR.Tn[12].n25 VGND 0.04199f
C8744 XThR.Tn[12].n26 VGND 0.0295f
C8745 XThR.Tn[12].n28 VGND 0.09466f
C8746 XThR.Tn[12].t48 VGND 0.01509f
C8747 XThR.Tn[12].t39 VGND 0.01653f
C8748 XThR.Tn[12].n29 VGND 0.04036f
C8749 XThR.Tn[12].t64 VGND 0.01504f
C8750 XThR.Tn[12].t17 VGND 0.01647f
C8751 XThR.Tn[12].n30 VGND 0.04199f
C8752 XThR.Tn[12].n31 VGND 0.0295f
C8753 XThR.Tn[12].n33 VGND 0.09466f
C8754 XThR.Tn[12].t23 VGND 0.01509f
C8755 XThR.Tn[12].t56 VGND 0.01653f
C8756 XThR.Tn[12].n34 VGND 0.04036f
C8757 XThR.Tn[12].t41 VGND 0.01504f
C8758 XThR.Tn[12].t37 VGND 0.01647f
C8759 XThR.Tn[12].n35 VGND 0.04199f
C8760 XThR.Tn[12].n36 VGND 0.0295f
C8761 XThR.Tn[12].n38 VGND 0.09466f
C8762 XThR.Tn[12].t54 VGND 0.01509f
C8763 XThR.Tn[12].t51 VGND 0.01653f
C8764 XThR.Tn[12].n39 VGND 0.04036f
C8765 XThR.Tn[12].t72 VGND 0.01504f
C8766 XThR.Tn[12].t29 VGND 0.01647f
C8767 XThR.Tn[12].n40 VGND 0.04199f
C8768 XThR.Tn[12].n41 VGND 0.0295f
C8769 XThR.Tn[12].n43 VGND 0.09466f
C8770 XThR.Tn[12].t59 VGND 0.01509f
C8771 XThR.Tn[12].t65 VGND 0.01653f
C8772 XThR.Tn[12].n44 VGND 0.04036f
C8773 XThR.Tn[12].t14 VGND 0.01504f
C8774 XThR.Tn[12].t44 VGND 0.01647f
C8775 XThR.Tn[12].n45 VGND 0.04199f
C8776 XThR.Tn[12].n46 VGND 0.0295f
C8777 XThR.Tn[12].n48 VGND 0.09466f
C8778 XThR.Tn[12].t12 VGND 0.01509f
C8779 XThR.Tn[12].t22 VGND 0.01653f
C8780 XThR.Tn[12].n49 VGND 0.04036f
C8781 XThR.Tn[12].t35 VGND 0.01504f
C8782 XThR.Tn[12].t61 VGND 0.01647f
C8783 XThR.Tn[12].n50 VGND 0.04199f
C8784 XThR.Tn[12].n51 VGND 0.0295f
C8785 XThR.Tn[12].n53 VGND 0.09466f
C8786 XThR.Tn[12].t68 VGND 0.01509f
C8787 XThR.Tn[12].t40 VGND 0.01653f
C8788 XThR.Tn[12].n54 VGND 0.04036f
C8789 XThR.Tn[12].t26 VGND 0.01504f
C8790 XThR.Tn[12].t19 VGND 0.01647f
C8791 XThR.Tn[12].n55 VGND 0.04199f
C8792 XThR.Tn[12].n56 VGND 0.0295f
C8793 XThR.Tn[12].n58 VGND 0.09466f
C8794 XThR.Tn[12].t25 VGND 0.01509f
C8795 XThR.Tn[12].t16 VGND 0.01653f
C8796 XThR.Tn[12].n59 VGND 0.04036f
C8797 XThR.Tn[12].t42 VGND 0.01504f
C8798 XThR.Tn[12].t55 VGND 0.01647f
C8799 XThR.Tn[12].n60 VGND 0.04199f
C8800 XThR.Tn[12].n61 VGND 0.0295f
C8801 XThR.Tn[12].n63 VGND 0.09466f
C8802 XThR.Tn[12].t57 VGND 0.01509f
C8803 XThR.Tn[12].t52 VGND 0.01653f
C8804 XThR.Tn[12].n64 VGND 0.04036f
C8805 XThR.Tn[12].t13 VGND 0.01504f
C8806 XThR.Tn[12].t31 VGND 0.01647f
C8807 XThR.Tn[12].n65 VGND 0.04199f
C8808 XThR.Tn[12].n66 VGND 0.0295f
C8809 XThR.Tn[12].n68 VGND 0.09466f
C8810 XThR.Tn[12].t73 VGND 0.01509f
C8811 XThR.Tn[12].t67 VGND 0.01653f
C8812 XThR.Tn[12].n69 VGND 0.04036f
C8813 XThR.Tn[12].t34 VGND 0.01504f
C8814 XThR.Tn[12].t47 VGND 0.01647f
C8815 XThR.Tn[12].n70 VGND 0.04199f
C8816 XThR.Tn[12].n71 VGND 0.0295f
C8817 XThR.Tn[12].n73 VGND 0.09466f
C8818 XThR.Tn[12].t32 VGND 0.01509f
C8819 XThR.Tn[12].t24 VGND 0.01653f
C8820 XThR.Tn[12].n74 VGND 0.04036f
C8821 XThR.Tn[12].t50 VGND 0.01504f
C8822 XThR.Tn[12].t62 VGND 0.01647f
C8823 XThR.Tn[12].n75 VGND 0.04199f
C8824 XThR.Tn[12].n76 VGND 0.0295f
C8825 XThR.Tn[12].n78 VGND 0.09466f
C8826 XThR.Tn[12].t69 VGND 0.01509f
C8827 XThR.Tn[12].t18 VGND 0.01653f
C8828 XThR.Tn[12].n79 VGND 0.04036f
C8829 XThR.Tn[12].t27 VGND 0.01504f
C8830 XThR.Tn[12].t58 VGND 0.01647f
C8831 XThR.Tn[12].n80 VGND 0.04199f
C8832 XThR.Tn[12].n81 VGND 0.0295f
C8833 XThR.Tn[12].n83 VGND 0.09466f
C8834 XThR.Tn[12].n84 VGND 0.08603f
C8835 XThR.Tn[12].n85 VGND 0.29341f
C8836 XThR.Tn[12].t2 VGND 0.01255f
C8837 XThR.Tn[12].t0 VGND 0.01255f
C8838 XThR.Tn[12].n86 VGND 0.0251f
C8839 XThR.Tn[12].t3 VGND 0.01255f
C8840 XThR.Tn[12].t1 VGND 0.01255f
C8841 XThR.Tn[12].n87 VGND 0.03131f
C8842 XThR.Tn[12].n88 VGND 0.05789f
C8843 XThR.Tn[14].t8 VGND 0.0197f
C8844 XThR.Tn[14].t9 VGND 0.0197f
C8845 XThR.Tn[14].n0 VGND 0.0598f
C8846 XThR.Tn[14].t10 VGND 0.0197f
C8847 XThR.Tn[14].t11 VGND 0.0197f
C8848 XThR.Tn[14].n1 VGND 0.04378f
C8849 XThR.Tn[14].n2 VGND 0.19909f
C8850 XThR.Tn[14].t6 VGND 0.0128f
C8851 XThR.Tn[14].t7 VGND 0.0128f
C8852 XThR.Tn[14].n3 VGND 0.03193f
C8853 XThR.Tn[14].t4 VGND 0.0128f
C8854 XThR.Tn[14].t5 VGND 0.0128f
C8855 XThR.Tn[14].n4 VGND 0.02561f
C8856 XThR.Tn[14].n5 VGND 0.05904f
C8857 XThR.Tn[14].t69 VGND 0.01539f
C8858 XThR.Tn[14].t62 VGND 0.01686f
C8859 XThR.Tn[14].n6 VGND 0.04116f
C8860 XThR.Tn[14].n7 VGND 0.07907f
C8861 XThR.Tn[14].t24 VGND 0.01539f
C8862 XThR.Tn[14].t13 VGND 0.01686f
C8863 XThR.Tn[14].n8 VGND 0.04116f
C8864 XThR.Tn[14].t28 VGND 0.01534f
C8865 XThR.Tn[14].t60 VGND 0.0168f
C8866 XThR.Tn[14].n9 VGND 0.04283f
C8867 XThR.Tn[14].n10 VGND 0.03009f
C8868 XThR.Tn[14].n12 VGND 0.09655f
C8869 XThR.Tn[14].t64 VGND 0.01539f
C8870 XThR.Tn[14].t54 VGND 0.01686f
C8871 XThR.Tn[14].n13 VGND 0.04116f
C8872 XThR.Tn[14].t67 VGND 0.01534f
C8873 XThR.Tn[14].t34 VGND 0.0168f
C8874 XThR.Tn[14].n14 VGND 0.04283f
C8875 XThR.Tn[14].n15 VGND 0.03009f
C8876 XThR.Tn[14].n17 VGND 0.09655f
C8877 XThR.Tn[14].t14 VGND 0.01539f
C8878 XThR.Tn[14].t72 VGND 0.01686f
C8879 XThR.Tn[14].n18 VGND 0.04116f
C8880 XThR.Tn[14].t17 VGND 0.01534f
C8881 XThR.Tn[14].t52 VGND 0.0168f
C8882 XThR.Tn[14].n19 VGND 0.04283f
C8883 XThR.Tn[14].n20 VGND 0.03009f
C8884 XThR.Tn[14].n22 VGND 0.09655f
C8885 XThR.Tn[14].t44 VGND 0.01539f
C8886 XThR.Tn[14].t38 VGND 0.01686f
C8887 XThR.Tn[14].n23 VGND 0.04116f
C8888 XThR.Tn[14].t47 VGND 0.01534f
C8889 XThR.Tn[14].t18 VGND 0.0168f
C8890 XThR.Tn[14].n24 VGND 0.04283f
C8891 XThR.Tn[14].n25 VGND 0.03009f
C8892 XThR.Tn[14].n27 VGND 0.09655f
C8893 XThR.Tn[14].t15 VGND 0.01539f
C8894 XThR.Tn[14].t73 VGND 0.01686f
C8895 XThR.Tn[14].n28 VGND 0.04116f
C8896 XThR.Tn[14].t21 VGND 0.01534f
C8897 XThR.Tn[14].t53 VGND 0.0168f
C8898 XThR.Tn[14].n29 VGND 0.04283f
C8899 XThR.Tn[14].n30 VGND 0.03009f
C8900 XThR.Tn[14].n32 VGND 0.09655f
C8901 XThR.Tn[14].t57 VGND 0.01539f
C8902 XThR.Tn[14].t25 VGND 0.01686f
C8903 XThR.Tn[14].n33 VGND 0.04116f
C8904 XThR.Tn[14].t61 VGND 0.01534f
C8905 XThR.Tn[14].t71 VGND 0.0168f
C8906 XThR.Tn[14].n34 VGND 0.04283f
C8907 XThR.Tn[14].n35 VGND 0.03009f
C8908 XThR.Tn[14].n37 VGND 0.09655f
C8909 XThR.Tn[14].t23 VGND 0.01539f
C8910 XThR.Tn[14].t19 VGND 0.01686f
C8911 XThR.Tn[14].n38 VGND 0.04116f
C8912 XThR.Tn[14].t29 VGND 0.01534f
C8913 XThR.Tn[14].t66 VGND 0.0168f
C8914 XThR.Tn[14].n39 VGND 0.04283f
C8915 XThR.Tn[14].n40 VGND 0.03009f
C8916 XThR.Tn[14].n42 VGND 0.09655f
C8917 XThR.Tn[14].t27 VGND 0.01539f
C8918 XThR.Tn[14].t36 VGND 0.01686f
C8919 XThR.Tn[14].n43 VGND 0.04116f
C8920 XThR.Tn[14].t33 VGND 0.01534f
C8921 XThR.Tn[14].t16 VGND 0.0168f
C8922 XThR.Tn[14].n44 VGND 0.04283f
C8923 XThR.Tn[14].n45 VGND 0.03009f
C8924 XThR.Tn[14].n47 VGND 0.09655f
C8925 XThR.Tn[14].t46 VGND 0.01539f
C8926 XThR.Tn[14].t56 VGND 0.01686f
C8927 XThR.Tn[14].n48 VGND 0.04116f
C8928 XThR.Tn[14].t50 VGND 0.01534f
C8929 XThR.Tn[14].t35 VGND 0.0168f
C8930 XThR.Tn[14].n49 VGND 0.04283f
C8931 XThR.Tn[14].n50 VGND 0.03009f
C8932 XThR.Tn[14].n52 VGND 0.09655f
C8933 XThR.Tn[14].t40 VGND 0.01539f
C8934 XThR.Tn[14].t12 VGND 0.01686f
C8935 XThR.Tn[14].n53 VGND 0.04116f
C8936 XThR.Tn[14].t42 VGND 0.01534f
C8937 XThR.Tn[14].t55 VGND 0.0168f
C8938 XThR.Tn[14].n54 VGND 0.04283f
C8939 XThR.Tn[14].n55 VGND 0.03009f
C8940 XThR.Tn[14].n57 VGND 0.09655f
C8941 XThR.Tn[14].t59 VGND 0.01539f
C8942 XThR.Tn[14].t49 VGND 0.01686f
C8943 XThR.Tn[14].n58 VGND 0.04116f
C8944 XThR.Tn[14].t63 VGND 0.01534f
C8945 XThR.Tn[14].t30 VGND 0.0168f
C8946 XThR.Tn[14].n59 VGND 0.04283f
C8947 XThR.Tn[14].n60 VGND 0.03009f
C8948 XThR.Tn[14].n62 VGND 0.09655f
C8949 XThR.Tn[14].t26 VGND 0.01539f
C8950 XThR.Tn[14].t22 VGND 0.01686f
C8951 XThR.Tn[14].n63 VGND 0.04116f
C8952 XThR.Tn[14].t31 VGND 0.01534f
C8953 XThR.Tn[14].t68 VGND 0.0168f
C8954 XThR.Tn[14].n64 VGND 0.04283f
C8955 XThR.Tn[14].n65 VGND 0.03009f
C8956 XThR.Tn[14].n67 VGND 0.09655f
C8957 XThR.Tn[14].t45 VGND 0.01539f
C8958 XThR.Tn[14].t39 VGND 0.01686f
C8959 XThR.Tn[14].n68 VGND 0.04116f
C8960 XThR.Tn[14].t48 VGND 0.01534f
C8961 XThR.Tn[14].t20 VGND 0.0168f
C8962 XThR.Tn[14].n69 VGND 0.04283f
C8963 XThR.Tn[14].n70 VGND 0.03009f
C8964 XThR.Tn[14].n72 VGND 0.09655f
C8965 XThR.Tn[14].t65 VGND 0.01539f
C8966 XThR.Tn[14].t58 VGND 0.01686f
C8967 XThR.Tn[14].n73 VGND 0.04116f
C8968 XThR.Tn[14].t70 VGND 0.01534f
C8969 XThR.Tn[14].t37 VGND 0.0168f
C8970 XThR.Tn[14].n74 VGND 0.04283f
C8971 XThR.Tn[14].n75 VGND 0.03009f
C8972 XThR.Tn[14].n77 VGND 0.09655f
C8973 XThR.Tn[14].t41 VGND 0.01539f
C8974 XThR.Tn[14].t51 VGND 0.01686f
C8975 XThR.Tn[14].n78 VGND 0.04116f
C8976 XThR.Tn[14].t43 VGND 0.01534f
C8977 XThR.Tn[14].t32 VGND 0.0168f
C8978 XThR.Tn[14].n79 VGND 0.04283f
C8979 XThR.Tn[14].n80 VGND 0.03009f
C8980 XThR.Tn[14].n82 VGND 0.09655f
C8981 XThR.Tn[14].n83 VGND 0.08774f
C8982 XThR.Tn[14].n84 VGND 0.35247f
C8983 XThR.Tn[14].t2 VGND 0.0197f
C8984 XThR.Tn[14].t3 VGND 0.0197f
C8985 XThR.Tn[14].n85 VGND 0.04256f
C8986 XThR.Tn[14].t0 VGND 0.0197f
C8987 XThR.Tn[14].t1 VGND 0.0197f
C8988 XThR.Tn[14].n86 VGND 0.06477f
C8989 XThR.Tn[14].n87 VGND 0.17985f
C8990 XThR.Tn[6].t7 VGND 0.01813f
C8991 XThR.Tn[6].t4 VGND 0.01813f
C8992 XThR.Tn[6].n0 VGND 0.0366f
C8993 XThR.Tn[6].t6 VGND 0.01813f
C8994 XThR.Tn[6].t5 VGND 0.01813f
C8995 XThR.Tn[6].n1 VGND 0.04282f
C8996 XThR.Tn[6].n2 VGND 0.12845f
C8997 XThR.Tn[6].t8 VGND 0.01179f
C8998 XThR.Tn[6].t9 VGND 0.01179f
C8999 XThR.Tn[6].n3 VGND 0.02684f
C9000 XThR.Tn[6].t11 VGND 0.01179f
C9001 XThR.Tn[6].t10 VGND 0.01179f
C9002 XThR.Tn[6].n4 VGND 0.02684f
C9003 XThR.Tn[6].t0 VGND 0.01179f
C9004 XThR.Tn[6].t1 VGND 0.01179f
C9005 XThR.Tn[6].n5 VGND 0.04472f
C9006 XThR.Tn[6].t3 VGND 0.01179f
C9007 XThR.Tn[6].t2 VGND 0.01179f
C9008 XThR.Tn[6].n6 VGND 0.02684f
C9009 XThR.Tn[6].n7 VGND 0.12781f
C9010 XThR.Tn[6].n8 VGND 0.07901f
C9011 XThR.Tn[6].n9 VGND 0.08917f
C9012 XThR.Tn[6].t62 VGND 0.01417f
C9013 XThR.Tn[6].t56 VGND 0.01552f
C9014 XThR.Tn[6].n10 VGND 0.03789f
C9015 XThR.Tn[6].n11 VGND 0.07279f
C9016 XThR.Tn[6].t20 VGND 0.01417f
C9017 XThR.Tn[6].t72 VGND 0.01552f
C9018 XThR.Tn[6].n12 VGND 0.03789f
C9019 XThR.Tn[6].t36 VGND 0.01412f
C9020 XThR.Tn[6].t68 VGND 0.01547f
C9021 XThR.Tn[6].n13 VGND 0.03943f
C9022 XThR.Tn[6].n14 VGND 0.0277f
C9023 XThR.Tn[6].n16 VGND 0.08888f
C9024 XThR.Tn[6].t57 VGND 0.01417f
C9025 XThR.Tn[6].t49 VGND 0.01552f
C9026 XThR.Tn[6].n17 VGND 0.03789f
C9027 XThR.Tn[6].t14 VGND 0.01412f
C9028 XThR.Tn[6].t45 VGND 0.01547f
C9029 XThR.Tn[6].n18 VGND 0.03943f
C9030 XThR.Tn[6].n19 VGND 0.0277f
C9031 XThR.Tn[6].n21 VGND 0.08888f
C9032 XThR.Tn[6].t73 VGND 0.01417f
C9033 XThR.Tn[6].t66 VGND 0.01552f
C9034 XThR.Tn[6].n22 VGND 0.03789f
C9035 XThR.Tn[6].t26 VGND 0.01412f
C9036 XThR.Tn[6].t63 VGND 0.01547f
C9037 XThR.Tn[6].n23 VGND 0.03943f
C9038 XThR.Tn[6].n24 VGND 0.0277f
C9039 XThR.Tn[6].n26 VGND 0.08888f
C9040 XThR.Tn[6].t35 VGND 0.01417f
C9041 XThR.Tn[6].t31 VGND 0.01552f
C9042 XThR.Tn[6].n27 VGND 0.03789f
C9043 XThR.Tn[6].t59 VGND 0.01412f
C9044 XThR.Tn[6].t27 VGND 0.01547f
C9045 XThR.Tn[6].n28 VGND 0.03943f
C9046 XThR.Tn[6].n29 VGND 0.0277f
C9047 XThR.Tn[6].n31 VGND 0.08888f
C9048 XThR.Tn[6].t13 VGND 0.01417f
C9049 XThR.Tn[6].t67 VGND 0.01552f
C9050 XThR.Tn[6].n32 VGND 0.03789f
C9051 XThR.Tn[6].t29 VGND 0.01412f
C9052 XThR.Tn[6].t64 VGND 0.01547f
C9053 XThR.Tn[6].n33 VGND 0.03943f
C9054 XThR.Tn[6].n34 VGND 0.0277f
C9055 XThR.Tn[6].n36 VGND 0.08888f
C9056 XThR.Tn[6].t51 VGND 0.01417f
C9057 XThR.Tn[6].t22 VGND 0.01552f
C9058 XThR.Tn[6].n37 VGND 0.03789f
C9059 XThR.Tn[6].t70 VGND 0.01412f
C9060 XThR.Tn[6].t19 VGND 0.01547f
C9061 XThR.Tn[6].n38 VGND 0.03943f
C9062 XThR.Tn[6].n39 VGND 0.0277f
C9063 XThR.Tn[6].n41 VGND 0.08888f
C9064 XThR.Tn[6].t21 VGND 0.01417f
C9065 XThR.Tn[6].t17 VGND 0.01552f
C9066 XThR.Tn[6].n42 VGND 0.03789f
C9067 XThR.Tn[6].t37 VGND 0.01412f
C9068 XThR.Tn[6].t12 VGND 0.01547f
C9069 XThR.Tn[6].n43 VGND 0.03943f
C9070 XThR.Tn[6].n44 VGND 0.0277f
C9071 XThR.Tn[6].n46 VGND 0.08888f
C9072 XThR.Tn[6].t24 VGND 0.01417f
C9073 XThR.Tn[6].t30 VGND 0.01552f
C9074 XThR.Tn[6].n47 VGND 0.03789f
C9075 XThR.Tn[6].t43 VGND 0.01412f
C9076 XThR.Tn[6].t25 VGND 0.01547f
C9077 XThR.Tn[6].n48 VGND 0.03943f
C9078 XThR.Tn[6].n49 VGND 0.0277f
C9079 XThR.Tn[6].n51 VGND 0.08888f
C9080 XThR.Tn[6].t40 VGND 0.01417f
C9081 XThR.Tn[6].t50 VGND 0.01552f
C9082 XThR.Tn[6].n52 VGND 0.03789f
C9083 XThR.Tn[6].t61 VGND 0.01412f
C9084 XThR.Tn[6].t47 VGND 0.01547f
C9085 XThR.Tn[6].n53 VGND 0.03943f
C9086 XThR.Tn[6].n54 VGND 0.0277f
C9087 XThR.Tn[6].n56 VGND 0.08888f
C9088 XThR.Tn[6].t33 VGND 0.01417f
C9089 XThR.Tn[6].t69 VGND 0.01552f
C9090 XThR.Tn[6].n57 VGND 0.03789f
C9091 XThR.Tn[6].t54 VGND 0.01412f
C9092 XThR.Tn[6].t65 VGND 0.01547f
C9093 XThR.Tn[6].n58 VGND 0.03943f
C9094 XThR.Tn[6].n59 VGND 0.0277f
C9095 XThR.Tn[6].n61 VGND 0.08888f
C9096 XThR.Tn[6].t53 VGND 0.01417f
C9097 XThR.Tn[6].t44 VGND 0.01552f
C9098 XThR.Tn[6].n62 VGND 0.03789f
C9099 XThR.Tn[6].t71 VGND 0.01412f
C9100 XThR.Tn[6].t39 VGND 0.01547f
C9101 XThR.Tn[6].n63 VGND 0.03943f
C9102 XThR.Tn[6].n64 VGND 0.0277f
C9103 XThR.Tn[6].n66 VGND 0.08888f
C9104 XThR.Tn[6].t23 VGND 0.01417f
C9105 XThR.Tn[6].t18 VGND 0.01552f
C9106 XThR.Tn[6].n67 VGND 0.03789f
C9107 XThR.Tn[6].t41 VGND 0.01412f
C9108 XThR.Tn[6].t15 VGND 0.01547f
C9109 XThR.Tn[6].n68 VGND 0.03943f
C9110 XThR.Tn[6].n69 VGND 0.0277f
C9111 XThR.Tn[6].n71 VGND 0.08888f
C9112 XThR.Tn[6].t38 VGND 0.01417f
C9113 XThR.Tn[6].t32 VGND 0.01552f
C9114 XThR.Tn[6].n72 VGND 0.03789f
C9115 XThR.Tn[6].t60 VGND 0.01412f
C9116 XThR.Tn[6].t28 VGND 0.01547f
C9117 XThR.Tn[6].n73 VGND 0.03943f
C9118 XThR.Tn[6].n74 VGND 0.0277f
C9119 XThR.Tn[6].n76 VGND 0.08888f
C9120 XThR.Tn[6].t58 VGND 0.01417f
C9121 XThR.Tn[6].t52 VGND 0.01552f
C9122 XThR.Tn[6].n77 VGND 0.03789f
C9123 XThR.Tn[6].t16 VGND 0.01412f
C9124 XThR.Tn[6].t48 VGND 0.01547f
C9125 XThR.Tn[6].n78 VGND 0.03943f
C9126 XThR.Tn[6].n79 VGND 0.0277f
C9127 XThR.Tn[6].n81 VGND 0.08888f
C9128 XThR.Tn[6].t34 VGND 0.01417f
C9129 XThR.Tn[6].t46 VGND 0.01552f
C9130 XThR.Tn[6].n82 VGND 0.03789f
C9131 XThR.Tn[6].t55 VGND 0.01412f
C9132 XThR.Tn[6].t42 VGND 0.01547f
C9133 XThR.Tn[6].n83 VGND 0.03943f
C9134 XThR.Tn[6].n84 VGND 0.0277f
C9135 XThR.Tn[6].n86 VGND 0.08888f
C9136 XThR.Tn[6].n87 VGND 0.08078f
C9137 XThR.Tn[6].n88 VGND 0.13446f
C9138 XA.Cn[10].n0 VGND 0.02345f
C9139 XA.Cn[10].n1 VGND 0.0188f
C9140 XA.Cn[10].n2 VGND 0.0473f
C9141 XA.Cn[10].t38 VGND 0.01146f
C9142 XA.Cn[10].t36 VGND 0.01252f
C9143 XA.Cn[10].n3 VGND 0.02796f
C9144 XA.Cn[10].n4 VGND 0.01598f
C9145 XA.Cn[10].n5 VGND 0.01943f
C9146 XA.Cn[10].t24 VGND 0.01146f
C9147 XA.Cn[10].t21 VGND 0.01252f
C9148 XA.Cn[10].n6 VGND 0.02796f
C9149 XA.Cn[10].n7 VGND 0.01598f
C9150 XA.Cn[10].n8 VGND 0.09232f
C9151 XA.Cn[10].t29 VGND 0.01146f
C9152 XA.Cn[10].t23 VGND 0.01252f
C9153 XA.Cn[10].n9 VGND 0.02796f
C9154 XA.Cn[10].n10 VGND 0.01598f
C9155 XA.Cn[10].n11 VGND 0.09232f
C9156 XA.Cn[10].t30 VGND 0.01146f
C9157 XA.Cn[10].t25 VGND 0.01252f
C9158 XA.Cn[10].n12 VGND 0.02796f
C9159 XA.Cn[10].n13 VGND 0.01598f
C9160 XA.Cn[10].n14 VGND 0.09232f
C9161 XA.Cn[10].t17 VGND 0.01146f
C9162 XA.Cn[10].t14 VGND 0.01252f
C9163 XA.Cn[10].n15 VGND 0.02796f
C9164 XA.Cn[10].n16 VGND 0.01598f
C9165 XA.Cn[10].n17 VGND 0.09232f
C9166 XA.Cn[10].t18 VGND 0.01146f
C9167 XA.Cn[10].t15 VGND 0.01252f
C9168 XA.Cn[10].n18 VGND 0.02796f
C9169 XA.Cn[10].n19 VGND 0.01598f
C9170 XA.Cn[10].n20 VGND 0.09232f
C9171 XA.Cn[10].t34 VGND 0.01146f
C9172 XA.Cn[10].t28 VGND 0.01252f
C9173 XA.Cn[10].n21 VGND 0.02796f
C9174 XA.Cn[10].n22 VGND 0.01598f
C9175 XA.Cn[10].n23 VGND 0.09232f
C9176 XA.Cn[10].t41 VGND 0.01146f
C9177 XA.Cn[10].t37 VGND 0.01252f
C9178 XA.Cn[10].n24 VGND 0.02796f
C9179 XA.Cn[10].n25 VGND 0.01598f
C9180 XA.Cn[10].n26 VGND 0.09232f
C9181 XA.Cn[10].t43 VGND 0.01146f
C9182 XA.Cn[10].t39 VGND 0.01252f
C9183 XA.Cn[10].n27 VGND 0.02796f
C9184 XA.Cn[10].n28 VGND 0.01598f
C9185 XA.Cn[10].n29 VGND 0.09232f
C9186 XA.Cn[10].t31 VGND 0.01146f
C9187 XA.Cn[10].t26 VGND 0.01252f
C9188 XA.Cn[10].n30 VGND 0.02796f
C9189 XA.Cn[10].n31 VGND 0.01598f
C9190 XA.Cn[10].n32 VGND 0.09232f
C9191 XA.Cn[10].t33 VGND 0.01146f
C9192 XA.Cn[10].t27 VGND 0.01252f
C9193 XA.Cn[10].n33 VGND 0.02796f
C9194 XA.Cn[10].n34 VGND 0.01598f
C9195 XA.Cn[10].n35 VGND 0.09232f
C9196 XA.Cn[10].t12 VGND 0.01146f
C9197 XA.Cn[10].t40 VGND 0.01252f
C9198 XA.Cn[10].n36 VGND 0.02796f
C9199 XA.Cn[10].n37 VGND 0.01598f
C9200 XA.Cn[10].n38 VGND 0.09232f
C9201 XA.Cn[10].t20 VGND 0.01146f
C9202 XA.Cn[10].t16 VGND 0.01252f
C9203 XA.Cn[10].n39 VGND 0.02796f
C9204 XA.Cn[10].n40 VGND 0.01598f
C9205 XA.Cn[10].n41 VGND 0.09232f
C9206 XA.Cn[10].t22 VGND 0.01146f
C9207 XA.Cn[10].t19 VGND 0.01252f
C9208 XA.Cn[10].n42 VGND 0.02796f
C9209 XA.Cn[10].n43 VGND 0.01598f
C9210 XA.Cn[10].n44 VGND 0.09232f
C9211 XA.Cn[10].t35 VGND 0.01146f
C9212 XA.Cn[10].t32 VGND 0.01252f
C9213 XA.Cn[10].n45 VGND 0.02796f
C9214 XA.Cn[10].n46 VGND 0.01598f
C9215 XA.Cn[10].n47 VGND 0.09232f
C9216 XA.Cn[10].t13 VGND 0.01146f
C9217 XA.Cn[10].t42 VGND 0.01252f
C9218 XA.Cn[10].n48 VGND 0.02796f
C9219 XA.Cn[10].n49 VGND 0.01598f
C9220 XA.Cn[10].n50 VGND 0.09232f
C9221 XA.Cn[10].n51 VGND 0.46113f
C9222 XA.Cn[10].n52 VGND 0.03515f
C9223 XA.Cn[10].t2 VGND 0.01446f
C9224 XA.Cn[10].t8 VGND 0.01446f
C9225 XA.Cn[10].n53 VGND 0.03125f
C9226 XA.Cn[10].t9 VGND 0.01446f
C9227 XA.Cn[10].t1 VGND 0.01446f
C9228 XA.Cn[10].n54 VGND 0.04756f
C9229 XA.Cn[10].n55 VGND 0.13215f
C9230 XA.Cn[10].n56 VGND 0.02078f
C9231 XA.Cn[10].t5 VGND 0.01446f
C9232 XA.Cn[10].t4 VGND 0.01446f
C9233 XA.Cn[10].n57 VGND 0.03215f
C9234 XA.Cn[10].t11 VGND 0.01446f
C9235 XA.Cn[10].t0 VGND 0.01446f
C9236 XA.Cn[10].n58 VGND 0.04391f
C9237 XA.Cn[10].n59 VGND 0.14309f
C9238 Iout.n0 VGND 0.22972f
C9239 Iout.n1 VGND 1.20114f
C9240 Iout.n2 VGND 0.22972f
C9241 Iout.n3 VGND 0.22972f
C9242 Iout.t144 VGND 0.02212f
C9243 Iout.n4 VGND 0.04919f
C9244 Iout.n5 VGND 0.19431f
C9245 Iout.n6 VGND 0.22972f
C9246 Iout.n7 VGND 1.20114f
C9247 Iout.n8 VGND 0.22972f
C9248 Iout.t170 VGND 0.02212f
C9249 Iout.n9 VGND 0.04919f
C9250 Iout.n10 VGND 0.19431f
C9251 Iout.n11 VGND 0.22972f
C9252 Iout.n12 VGND 1.20114f
C9253 Iout.n13 VGND 0.22972f
C9254 Iout.t11 VGND 0.02212f
C9255 Iout.n14 VGND 0.04919f
C9256 Iout.n15 VGND 0.19431f
C9257 Iout.n16 VGND 0.22972f
C9258 Iout.n17 VGND 1.20114f
C9259 Iout.n18 VGND 0.22972f
C9260 Iout.t56 VGND 0.02212f
C9261 Iout.n19 VGND 0.04919f
C9262 Iout.n20 VGND 0.19431f
C9263 Iout.n21 VGND 0.47625f
C9264 Iout.t223 VGND 0.02212f
C9265 Iout.n22 VGND 0.04919f
C9266 Iout.n23 VGND 0.28657f
C9267 Iout.n24 VGND 0.22972f
C9268 Iout.n25 VGND 0.22972f
C9269 Iout.n26 VGND 0.22972f
C9270 Iout.n27 VGND 0.22972f
C9271 Iout.n28 VGND 0.22972f
C9272 Iout.n29 VGND 0.22972f
C9273 Iout.n30 VGND 0.22972f
C9274 Iout.n31 VGND 0.22972f
C9275 Iout.n32 VGND 0.22972f
C9276 Iout.n33 VGND 0.22972f
C9277 Iout.n34 VGND 0.22972f
C9278 Iout.n35 VGND 0.22972f
C9279 Iout.n36 VGND 0.22972f
C9280 Iout.n37 VGND 0.22972f
C9281 Iout.t61 VGND 0.02212f
C9282 Iout.n38 VGND 0.04919f
C9283 Iout.n39 VGND 0.02502f
C9284 Iout.n40 VGND 0.22972f
C9285 Iout.n41 VGND 0.04584f
C9286 Iout.t103 VGND 0.02212f
C9287 Iout.n42 VGND 0.04919f
C9288 Iout.n43 VGND 0.02502f
C9289 Iout.t241 VGND 0.02212f
C9290 Iout.n44 VGND 0.04919f
C9291 Iout.n45 VGND 0.02502f
C9292 Iout.n46 VGND 0.22972f
C9293 Iout.t185 VGND 0.02212f
C9294 Iout.n47 VGND 0.04919f
C9295 Iout.n48 VGND 0.02502f
C9296 Iout.n49 VGND 0.22972f
C9297 Iout.t77 VGND 0.02212f
C9298 Iout.n50 VGND 0.04919f
C9299 Iout.n51 VGND 0.02502f
C9300 Iout.n52 VGND 0.22972f
C9301 Iout.t159 VGND 0.02212f
C9302 Iout.n53 VGND 0.04919f
C9303 Iout.n54 VGND 0.02502f
C9304 Iout.n55 VGND 0.22972f
C9305 Iout.t39 VGND 0.02212f
C9306 Iout.n56 VGND 0.04919f
C9307 Iout.n57 VGND 0.02502f
C9308 Iout.n58 VGND 0.22972f
C9309 Iout.t101 VGND 0.02212f
C9310 Iout.n59 VGND 0.04919f
C9311 Iout.n60 VGND 0.02502f
C9312 Iout.n61 VGND 0.22972f
C9313 Iout.t240 VGND 0.02212f
C9314 Iout.n62 VGND 0.04919f
C9315 Iout.n63 VGND 0.02502f
C9316 Iout.n64 VGND 0.22972f
C9317 Iout.t202 VGND 0.02212f
C9318 Iout.n65 VGND 0.04919f
C9319 Iout.n66 VGND 0.02502f
C9320 Iout.n67 VGND 0.22972f
C9321 Iout.t250 VGND 0.02212f
C9322 Iout.n68 VGND 0.04919f
C9323 Iout.n69 VGND 0.02502f
C9324 Iout.n70 VGND 0.22972f
C9325 Iout.t59 VGND 0.02212f
C9326 Iout.n71 VGND 0.04919f
C9327 Iout.n72 VGND 0.02502f
C9328 Iout.n73 VGND 0.22972f
C9329 Iout.t32 VGND 0.02212f
C9330 Iout.n74 VGND 0.04919f
C9331 Iout.n75 VGND 0.02502f
C9332 Iout.n76 VGND 0.22972f
C9333 Iout.t171 VGND 0.02212f
C9334 Iout.n77 VGND 0.04919f
C9335 Iout.n78 VGND 0.02502f
C9336 Iout.n79 VGND 0.22972f
C9337 Iout.n80 VGND 0.22972f
C9338 Iout.t118 VGND 0.02212f
C9339 Iout.n81 VGND 0.04919f
C9340 Iout.n82 VGND 0.02502f
C9341 Iout.n83 VGND 0.22972f
C9342 Iout.n84 VGND 0.04584f
C9343 Iout.t81 VGND 0.02212f
C9344 Iout.n85 VGND 0.04919f
C9345 Iout.n86 VGND 0.02502f
C9346 Iout.t208 VGND 0.02212f
C9347 Iout.n87 VGND 0.04919f
C9348 Iout.n88 VGND 0.02502f
C9349 Iout.n89 VGND 0.22972f
C9350 Iout.t215 VGND 0.02212f
C9351 Iout.n90 VGND 0.04919f
C9352 Iout.n91 VGND 0.02502f
C9353 Iout.n92 VGND 0.22972f
C9354 Iout.t134 VGND 0.02212f
C9355 Iout.n93 VGND 0.04919f
C9356 Iout.n94 VGND 0.02502f
C9357 Iout.n95 VGND 0.22972f
C9358 Iout.t74 VGND 0.02212f
C9359 Iout.n96 VGND 0.04919f
C9360 Iout.n97 VGND 0.02502f
C9361 Iout.n98 VGND 0.22972f
C9362 Iout.t141 VGND 0.02212f
C9363 Iout.n99 VGND 0.04919f
C9364 Iout.n100 VGND 0.02502f
C9365 Iout.n101 VGND 0.22972f
C9366 Iout.t149 VGND 0.02212f
C9367 Iout.n102 VGND 0.04919f
C9368 Iout.n103 VGND 0.02502f
C9369 Iout.n104 VGND 0.22972f
C9370 Iout.t104 VGND 0.02212f
C9371 Iout.n105 VGND 0.04919f
C9372 Iout.n106 VGND 0.02502f
C9373 Iout.n107 VGND 0.22972f
C9374 Iout.t29 VGND 0.02212f
C9375 Iout.n108 VGND 0.04919f
C9376 Iout.n109 VGND 0.02502f
C9377 Iout.n110 VGND 0.22972f
C9378 Iout.t122 VGND 0.02212f
C9379 Iout.n111 VGND 0.04919f
C9380 Iout.n112 VGND 0.02502f
C9381 Iout.n113 VGND 0.22972f
C9382 Iout.t130 VGND 0.02212f
C9383 Iout.n114 VGND 0.04919f
C9384 Iout.n115 VGND 0.02502f
C9385 Iout.n116 VGND 0.22972f
C9386 Iout.t82 VGND 0.02212f
C9387 Iout.n117 VGND 0.04919f
C9388 Iout.n118 VGND 0.02502f
C9389 Iout.n119 VGND 0.22972f
C9390 Iout.t0 VGND 0.02212f
C9391 Iout.n120 VGND 0.04919f
C9392 Iout.n121 VGND 0.02502f
C9393 Iout.n122 VGND 0.04584f
C9394 Iout.t150 VGND 0.02212f
C9395 Iout.n123 VGND 0.04919f
C9396 Iout.n124 VGND 0.02502f
C9397 Iout.n125 VGND 0.22972f
C9398 Iout.n126 VGND 0.22972f
C9399 Iout.t152 VGND 0.02212f
C9400 Iout.n127 VGND 0.04919f
C9401 Iout.n128 VGND 0.02502f
C9402 Iout.n129 VGND 0.04584f
C9403 Iout.t210 VGND 0.02212f
C9404 Iout.n130 VGND 0.04919f
C9405 Iout.n131 VGND 0.02502f
C9406 Iout.n132 VGND 0.22972f
C9407 Iout.t47 VGND 0.02212f
C9408 Iout.n133 VGND 0.04919f
C9409 Iout.n134 VGND 0.02502f
C9410 Iout.n135 VGND 0.04584f
C9411 Iout.t230 VGND 0.02212f
C9412 Iout.n136 VGND 0.04919f
C9413 Iout.n137 VGND 0.02502f
C9414 Iout.n138 VGND 0.22972f
C9415 Iout.n139 VGND 0.22972f
C9416 Iout.t253 VGND 0.02212f
C9417 Iout.n140 VGND 0.04919f
C9418 Iout.n141 VGND 0.02502f
C9419 Iout.n142 VGND 0.04584f
C9420 Iout.t9 VGND 0.02212f
C9421 Iout.n143 VGND 0.04919f
C9422 Iout.n144 VGND 0.02502f
C9423 Iout.n145 VGND 0.13561f
C9424 Iout.t217 VGND 0.02212f
C9425 Iout.n146 VGND 0.04919f
C9426 Iout.n147 VGND 0.02502f
C9427 Iout.n148 VGND 0.04584f
C9428 Iout.t102 VGND 0.02212f
C9429 Iout.n149 VGND 0.04919f
C9430 Iout.n150 VGND 0.02502f
C9431 Iout.n151 VGND 0.22972f
C9432 Iout.n152 VGND 0.13561f
C9433 Iout.n153 VGND 0.22972f
C9434 Iout.n154 VGND 0.22972f
C9435 Iout.n155 VGND 0.22972f
C9436 Iout.t94 VGND 0.02212f
C9437 Iout.n156 VGND 0.04919f
C9438 Iout.n157 VGND 0.02502f
C9439 Iout.n158 VGND 0.22972f
C9440 Iout.n159 VGND 0.22972f
C9441 Iout.n160 VGND 0.22972f
C9442 Iout.n161 VGND 0.22972f
C9443 Iout.n162 VGND 0.22972f
C9444 Iout.n163 VGND 0.22972f
C9445 Iout.n164 VGND 0.22972f
C9446 Iout.n165 VGND 0.22972f
C9447 Iout.n166 VGND 0.22972f
C9448 Iout.n167 VGND 0.22972f
C9449 Iout.t251 VGND 0.02212f
C9450 Iout.n168 VGND 0.04919f
C9451 Iout.n169 VGND 0.02502f
C9452 Iout.n170 VGND 0.22972f
C9453 Iout.n171 VGND 0.04584f
C9454 Iout.t212 VGND 0.02212f
C9455 Iout.n172 VGND 0.04919f
C9456 Iout.n173 VGND 0.02502f
C9457 Iout.t188 VGND 0.02212f
C9458 Iout.n174 VGND 0.04919f
C9459 Iout.n175 VGND 0.02502f
C9460 Iout.n176 VGND 0.22972f
C9461 Iout.t129 VGND 0.02212f
C9462 Iout.n177 VGND 0.04919f
C9463 Iout.n178 VGND 0.02502f
C9464 Iout.n179 VGND 0.22972f
C9465 Iout.t84 VGND 0.02212f
C9466 Iout.n180 VGND 0.04919f
C9467 Iout.n181 VGND 0.02502f
C9468 Iout.n182 VGND 0.22972f
C9469 Iout.t14 VGND 0.02212f
C9470 Iout.n183 VGND 0.04919f
C9471 Iout.n184 VGND 0.02502f
C9472 Iout.n185 VGND 0.22972f
C9473 Iout.t51 VGND 0.02212f
C9474 Iout.n186 VGND 0.04919f
C9475 Iout.n187 VGND 0.02502f
C9476 Iout.n188 VGND 0.22972f
C9477 Iout.t18 VGND 0.02212f
C9478 Iout.n189 VGND 0.04919f
C9479 Iout.n190 VGND 0.02502f
C9480 Iout.n191 VGND 0.13561f
C9481 Iout.t175 VGND 0.02212f
C9482 Iout.n192 VGND 0.04919f
C9483 Iout.n193 VGND 0.02502f
C9484 Iout.n194 VGND 0.04584f
C9485 Iout.t234 VGND 0.02212f
C9486 Iout.n195 VGND 0.04919f
C9487 Iout.n196 VGND 0.02502f
C9488 Iout.n197 VGND 0.13561f
C9489 Iout.n198 VGND 0.04584f
C9490 Iout.t143 VGND 0.02212f
C9491 Iout.n199 VGND 0.04919f
C9492 Iout.n200 VGND 0.02502f
C9493 Iout.n201 VGND 0.04584f
C9494 Iout.t75 VGND 0.02212f
C9495 Iout.n202 VGND 0.04919f
C9496 Iout.n203 VGND 0.02502f
C9497 Iout.n204 VGND 0.13561f
C9498 Iout.n205 VGND 0.04584f
C9499 Iout.t187 VGND 0.02212f
C9500 Iout.n206 VGND 0.04919f
C9501 Iout.n207 VGND 0.02502f
C9502 Iout.n208 VGND 0.13561f
C9503 Iout.n209 VGND 0.04584f
C9504 Iout.t44 VGND 0.02212f
C9505 Iout.n210 VGND 0.04919f
C9506 Iout.n211 VGND 0.02502f
C9507 Iout.n212 VGND 0.13561f
C9508 Iout.n213 VGND 0.04584f
C9509 Iout.t6 VGND 0.02212f
C9510 Iout.n214 VGND 0.04919f
C9511 Iout.n215 VGND 0.02502f
C9512 Iout.n216 VGND 0.13561f
C9513 Iout.n217 VGND 0.04584f
C9514 Iout.t52 VGND 0.02212f
C9515 Iout.n218 VGND 0.04919f
C9516 Iout.n219 VGND 0.02502f
C9517 Iout.n220 VGND 0.13561f
C9518 Iout.n221 VGND 0.04584f
C9519 Iout.t115 VGND 0.02212f
C9520 Iout.n222 VGND 0.04919f
C9521 Iout.n223 VGND 0.02502f
C9522 Iout.n224 VGND 0.13561f
C9523 Iout.n225 VGND 0.04584f
C9524 Iout.t116 VGND 0.02212f
C9525 Iout.n226 VGND 0.04919f
C9526 Iout.n227 VGND 0.02502f
C9527 Iout.n228 VGND 0.04584f
C9528 Iout.n229 VGND 0.13561f
C9529 Iout.n230 VGND 0.22972f
C9530 Iout.n231 VGND 0.04584f
C9531 Iout.t199 VGND 0.02212f
C9532 Iout.n232 VGND 0.04919f
C9533 Iout.n233 VGND 0.02502f
C9534 Iout.n234 VGND 0.04584f
C9535 Iout.t196 VGND 0.02212f
C9536 Iout.n235 VGND 0.04919f
C9537 Iout.n236 VGND 0.02502f
C9538 Iout.n237 VGND 0.04584f
C9539 Iout.t89 VGND 0.02212f
C9540 Iout.n238 VGND 0.04919f
C9541 Iout.n239 VGND 0.02502f
C9542 Iout.n240 VGND 0.04584f
C9543 Iout.t88 VGND 0.02212f
C9544 Iout.n241 VGND 0.04919f
C9545 Iout.n242 VGND 0.02502f
C9546 Iout.n243 VGND 0.04584f
C9547 Iout.t254 VGND 0.02212f
C9548 Iout.n244 VGND 0.04919f
C9549 Iout.n245 VGND 0.02502f
C9550 Iout.n246 VGND 0.04584f
C9551 Iout.t20 VGND 0.02212f
C9552 Iout.n247 VGND 0.04919f
C9553 Iout.n248 VGND 0.02502f
C9554 Iout.n249 VGND 0.04584f
C9555 Iout.t19 VGND 0.02212f
C9556 Iout.n250 VGND 0.04919f
C9557 Iout.n251 VGND 0.02502f
C9558 Iout.t72 VGND 0.02212f
C9559 Iout.n252 VGND 0.04919f
C9560 Iout.n253 VGND 0.02502f
C9561 Iout.n254 VGND 0.04584f
C9562 Iout.t5 VGND 0.02212f
C9563 Iout.n255 VGND 0.04919f
C9564 Iout.n256 VGND 0.02502f
C9565 Iout.n257 VGND 0.04584f
C9566 Iout.n258 VGND 0.22972f
C9567 Iout.t169 VGND 0.02212f
C9568 Iout.n259 VGND 0.04919f
C9569 Iout.n260 VGND 0.02502f
C9570 Iout.n261 VGND 0.04584f
C9571 Iout.n262 VGND 0.22972f
C9572 Iout.n263 VGND 0.22972f
C9573 Iout.n264 VGND 0.04584f
C9574 Iout.t41 VGND 0.02212f
C9575 Iout.n265 VGND 0.04919f
C9576 Iout.n266 VGND 0.02502f
C9577 Iout.n267 VGND 0.04584f
C9578 Iout.n268 VGND 0.22972f
C9579 Iout.n269 VGND 0.22972f
C9580 Iout.n270 VGND 0.04584f
C9581 Iout.t93 VGND 0.02212f
C9582 Iout.n271 VGND 0.04919f
C9583 Iout.n272 VGND 0.02502f
C9584 Iout.n273 VGND 0.04584f
C9585 Iout.n274 VGND 0.22972f
C9586 Iout.n275 VGND 0.22972f
C9587 Iout.n276 VGND 0.04584f
C9588 Iout.t62 VGND 0.02212f
C9589 Iout.n277 VGND 0.04919f
C9590 Iout.n278 VGND 0.02502f
C9591 Iout.n279 VGND 0.04584f
C9592 Iout.n280 VGND 0.22972f
C9593 Iout.n281 VGND 0.22972f
C9594 Iout.n282 VGND 0.04584f
C9595 Iout.t3 VGND 0.02212f
C9596 Iout.n283 VGND 0.04919f
C9597 Iout.n284 VGND 0.02502f
C9598 Iout.n285 VGND 0.04584f
C9599 Iout.n286 VGND 0.22972f
C9600 Iout.n287 VGND 0.22972f
C9601 Iout.n288 VGND 0.04584f
C9602 Iout.t165 VGND 0.02212f
C9603 Iout.n289 VGND 0.04919f
C9604 Iout.n290 VGND 0.02502f
C9605 Iout.n291 VGND 0.04584f
C9606 Iout.n292 VGND 0.22972f
C9607 Iout.n293 VGND 0.22972f
C9608 Iout.n294 VGND 0.04584f
C9609 Iout.t58 VGND 0.02212f
C9610 Iout.n295 VGND 0.04919f
C9611 Iout.n296 VGND 0.02502f
C9612 Iout.n297 VGND 0.04584f
C9613 Iout.n298 VGND 0.22972f
C9614 Iout.n299 VGND 0.22972f
C9615 Iout.n300 VGND 0.04584f
C9616 Iout.t55 VGND 0.02212f
C9617 Iout.n301 VGND 0.04919f
C9618 Iout.n302 VGND 0.02502f
C9619 Iout.n303 VGND 0.04584f
C9620 Iout.n304 VGND 0.22972f
C9621 Iout.t121 VGND 0.02212f
C9622 Iout.n305 VGND 0.04919f
C9623 Iout.n306 VGND 0.02502f
C9624 Iout.n307 VGND 0.04584f
C9625 Iout.t136 VGND 0.02212f
C9626 Iout.n308 VGND 0.04919f
C9627 Iout.n309 VGND 0.02502f
C9628 Iout.n310 VGND 0.04584f
C9629 Iout.t168 VGND 0.02212f
C9630 Iout.n311 VGND 0.04919f
C9631 Iout.n312 VGND 0.02502f
C9632 Iout.n313 VGND 0.04584f
C9633 Iout.t239 VGND 0.02212f
C9634 Iout.n314 VGND 0.04919f
C9635 Iout.n315 VGND 0.02502f
C9636 Iout.n316 VGND 0.04584f
C9637 Iout.t109 VGND 0.02212f
C9638 Iout.n317 VGND 0.04919f
C9639 Iout.n318 VGND 0.02502f
C9640 Iout.n319 VGND 0.04584f
C9641 Iout.t139 VGND 0.02212f
C9642 Iout.n320 VGND 0.04919f
C9643 Iout.n321 VGND 0.02502f
C9644 Iout.n322 VGND 0.04584f
C9645 Iout.t200 VGND 0.02212f
C9646 Iout.n323 VGND 0.04919f
C9647 Iout.n324 VGND 0.02502f
C9648 Iout.n325 VGND 0.04584f
C9649 Iout.t133 VGND 0.02212f
C9650 Iout.n326 VGND 0.04919f
C9651 Iout.n327 VGND 0.02502f
C9652 Iout.n328 VGND 0.04584f
C9653 Iout.t22 VGND 0.02212f
C9654 Iout.n329 VGND 0.04919f
C9655 Iout.n330 VGND 0.02502f
C9656 Iout.n331 VGND 0.04584f
C9657 Iout.n332 VGND 0.22972f
C9658 Iout.t227 VGND 0.02212f
C9659 Iout.n333 VGND 0.04919f
C9660 Iout.n334 VGND 0.02502f
C9661 Iout.n335 VGND 0.04584f
C9662 Iout.t117 VGND 0.02212f
C9663 Iout.n336 VGND 0.04919f
C9664 Iout.n337 VGND 0.02502f
C9665 Iout.n338 VGND 0.04584f
C9666 Iout.t157 VGND 0.02212f
C9667 Iout.n339 VGND 0.04919f
C9668 Iout.n340 VGND 0.02502f
C9669 Iout.n341 VGND 0.04584f
C9670 Iout.t194 VGND 0.02212f
C9671 Iout.n342 VGND 0.04919f
C9672 Iout.n343 VGND 0.02502f
C9673 Iout.n344 VGND 0.04584f
C9674 Iout.t123 VGND 0.02212f
C9675 Iout.n345 VGND 0.04919f
C9676 Iout.n346 VGND 0.02502f
C9677 Iout.n347 VGND 0.04584f
C9678 Iout.t191 VGND 0.02212f
C9679 Iout.n348 VGND 0.04919f
C9680 Iout.n349 VGND 0.02502f
C9681 Iout.n350 VGND 0.04584f
C9682 Iout.t78 VGND 0.02212f
C9683 Iout.n351 VGND 0.04919f
C9684 Iout.n352 VGND 0.02502f
C9685 Iout.n353 VGND 0.04584f
C9686 Iout.t131 VGND 0.02212f
C9687 Iout.n354 VGND 0.04919f
C9688 Iout.n355 VGND 0.02502f
C9689 Iout.n356 VGND 0.04584f
C9690 Iout.t192 VGND 0.02212f
C9691 Iout.n357 VGND 0.04919f
C9692 Iout.n358 VGND 0.02502f
C9693 Iout.n359 VGND 0.04584f
C9694 Iout.t110 VGND 0.02212f
C9695 Iout.n360 VGND 0.04919f
C9696 Iout.n361 VGND 0.02502f
C9697 Iout.n362 VGND 0.04584f
C9698 Iout.t229 VGND 0.02212f
C9699 Iout.n363 VGND 0.04919f
C9700 Iout.n364 VGND 0.02502f
C9701 Iout.n365 VGND 0.04584f
C9702 Iout.t90 VGND 0.02212f
C9703 Iout.n366 VGND 0.04919f
C9704 Iout.n367 VGND 0.02502f
C9705 Iout.n368 VGND 0.04584f
C9706 Iout.n369 VGND 0.22972f
C9707 Iout.t28 VGND 0.02212f
C9708 Iout.n370 VGND 0.04919f
C9709 Iout.n371 VGND 0.02502f
C9710 Iout.n372 VGND 0.04584f
C9711 Iout.n373 VGND 0.22972f
C9712 Iout.n374 VGND 0.22972f
C9713 Iout.n375 VGND 0.04584f
C9714 Iout.t43 VGND 0.02212f
C9715 Iout.n376 VGND 0.04919f
C9716 Iout.n377 VGND 0.02502f
C9717 Iout.t235 VGND 0.02212f
C9718 Iout.n378 VGND 0.04919f
C9719 Iout.n379 VGND 0.02502f
C9720 Iout.n380 VGND 0.04584f
C9721 Iout.n381 VGND 0.22972f
C9722 Iout.n382 VGND 0.22972f
C9723 Iout.n383 VGND 0.04584f
C9724 Iout.t178 VGND 0.02212f
C9725 Iout.n384 VGND 0.04919f
C9726 Iout.n385 VGND 0.02502f
C9727 Iout.t38 VGND 0.02212f
C9728 Iout.n386 VGND 0.04919f
C9729 Iout.n387 VGND 0.02502f
C9730 Iout.n388 VGND 0.04584f
C9731 Iout.n389 VGND 0.22972f
C9732 Iout.n390 VGND 0.22972f
C9733 Iout.n391 VGND 0.04584f
C9734 Iout.t111 VGND 0.02212f
C9735 Iout.n392 VGND 0.04919f
C9736 Iout.n393 VGND 0.02502f
C9737 Iout.t154 VGND 0.02212f
C9738 Iout.n394 VGND 0.04919f
C9739 Iout.n395 VGND 0.02502f
C9740 Iout.n396 VGND 0.04584f
C9741 Iout.n397 VGND 0.22972f
C9742 Iout.n398 VGND 0.22972f
C9743 Iout.n399 VGND 0.04584f
C9744 Iout.t120 VGND 0.02212f
C9745 Iout.n400 VGND 0.04919f
C9746 Iout.n401 VGND 0.02502f
C9747 Iout.t7 VGND 0.02212f
C9748 Iout.n402 VGND 0.04919f
C9749 Iout.n403 VGND 0.02502f
C9750 Iout.n404 VGND 0.04584f
C9751 Iout.n405 VGND 0.22972f
C9752 Iout.n406 VGND 0.22972f
C9753 Iout.n407 VGND 0.04584f
C9754 Iout.t8 VGND 0.02212f
C9755 Iout.n408 VGND 0.04919f
C9756 Iout.n409 VGND 0.02502f
C9757 Iout.t180 VGND 0.02212f
C9758 Iout.n410 VGND 0.04919f
C9759 Iout.n411 VGND 0.02502f
C9760 Iout.n412 VGND 0.04584f
C9761 Iout.n413 VGND 0.22972f
C9762 Iout.n414 VGND 0.22972f
C9763 Iout.n415 VGND 0.04584f
C9764 Iout.t45 VGND 0.02212f
C9765 Iout.n416 VGND 0.04919f
C9766 Iout.n417 VGND 0.02502f
C9767 Iout.t70 VGND 0.02212f
C9768 Iout.n418 VGND 0.04919f
C9769 Iout.n419 VGND 0.02502f
C9770 Iout.n420 VGND 0.04584f
C9771 Iout.n421 VGND 0.22972f
C9772 Iout.n422 VGND 0.22972f
C9773 Iout.n423 VGND 0.04584f
C9774 Iout.t206 VGND 0.02212f
C9775 Iout.n424 VGND 0.04919f
C9776 Iout.n425 VGND 0.02502f
C9777 Iout.t203 VGND 0.02212f
C9778 Iout.n426 VGND 0.04919f
C9779 Iout.n427 VGND 0.02502f
C9780 Iout.n428 VGND 0.04584f
C9781 Iout.n429 VGND 0.22972f
C9782 Iout.n430 VGND 0.22972f
C9783 Iout.n431 VGND 0.04584f
C9784 Iout.t164 VGND 0.02212f
C9785 Iout.n432 VGND 0.04919f
C9786 Iout.n433 VGND 0.02502f
C9787 Iout.t189 VGND 0.02212f
C9788 Iout.n434 VGND 0.04919f
C9789 Iout.n435 VGND 0.02502f
C9790 Iout.n436 VGND 0.22972f
C9791 Iout.n437 VGND 0.04584f
C9792 Iout.t233 VGND 0.02212f
C9793 Iout.n438 VGND 0.04919f
C9794 Iout.n439 VGND 0.02502f
C9795 Iout.n440 VGND 0.04584f
C9796 Iout.t176 VGND 0.02212f
C9797 Iout.n441 VGND 0.04919f
C9798 Iout.n442 VGND 0.02502f
C9799 Iout.n443 VGND 0.04584f
C9800 Iout.n444 VGND 0.22972f
C9801 Iout.n445 VGND 0.22972f
C9802 Iout.n446 VGND 0.04584f
C9803 Iout.t218 VGND 0.02212f
C9804 Iout.n447 VGND 0.04919f
C9805 Iout.n448 VGND 0.02502f
C9806 Iout.t63 VGND 0.02212f
C9807 Iout.n449 VGND 0.04919f
C9808 Iout.n450 VGND 0.02502f
C9809 Iout.n451 VGND 0.04584f
C9810 Iout.t65 VGND 0.02212f
C9811 Iout.n452 VGND 0.04919f
C9812 Iout.n453 VGND 0.02502f
C9813 Iout.n454 VGND 0.04584f
C9814 Iout.n455 VGND 0.22972f
C9815 Iout.n456 VGND 0.22972f
C9816 Iout.n457 VGND 0.04584f
C9817 Iout.t126 VGND 0.02212f
C9818 Iout.n458 VGND 0.04919f
C9819 Iout.n459 VGND 0.02502f
C9820 Iout.t177 VGND 0.02212f
C9821 Iout.n460 VGND 0.04919f
C9822 Iout.n461 VGND 0.02502f
C9823 Iout.n462 VGND 0.04584f
C9824 Iout.t232 VGND 0.02212f
C9825 Iout.n463 VGND 0.04919f
C9826 Iout.n464 VGND 0.02502f
C9827 Iout.n465 VGND 0.04584f
C9828 Iout.n466 VGND 0.22972f
C9829 Iout.n467 VGND 0.22972f
C9830 Iout.n468 VGND 0.04584f
C9831 Iout.t153 VGND 0.02212f
C9832 Iout.n469 VGND 0.04919f
C9833 Iout.n470 VGND 0.02502f
C9834 Iout.n471 VGND 0.04584f
C9835 Iout.t221 VGND 0.02212f
C9836 Iout.n472 VGND 0.04919f
C9837 Iout.n473 VGND 0.02502f
C9838 Iout.n474 VGND 0.04584f
C9839 Iout.n475 VGND 0.22972f
C9840 Iout.n476 VGND 0.22972f
C9841 Iout.n477 VGND 0.04584f
C9842 Iout.t247 VGND 0.02212f
C9843 Iout.n478 VGND 0.04919f
C9844 Iout.n479 VGND 0.02502f
C9845 Iout.t156 VGND 0.02212f
C9846 Iout.n480 VGND 0.04919f
C9847 Iout.n481 VGND 0.02502f
C9848 Iout.n482 VGND 0.04584f
C9849 Iout.t57 VGND 0.02212f
C9850 Iout.n483 VGND 0.04919f
C9851 Iout.n484 VGND 0.02502f
C9852 Iout.n485 VGND 0.04584f
C9853 Iout.n486 VGND 0.22972f
C9854 Iout.n487 VGND 0.22972f
C9855 Iout.n488 VGND 0.04584f
C9856 Iout.t30 VGND 0.02212f
C9857 Iout.n489 VGND 0.04919f
C9858 Iout.n490 VGND 0.02502f
C9859 Iout.t91 VGND 0.02212f
C9860 Iout.n491 VGND 0.04919f
C9861 Iout.n492 VGND 0.02502f
C9862 Iout.n493 VGND 0.04584f
C9863 Iout.t207 VGND 0.02212f
C9864 Iout.n494 VGND 0.04919f
C9865 Iout.n495 VGND 0.02502f
C9866 Iout.n496 VGND 0.04584f
C9867 Iout.n497 VGND 0.22972f
C9868 Iout.n498 VGND 0.13561f
C9869 Iout.n499 VGND 0.04584f
C9870 Iout.t98 VGND 0.02212f
C9871 Iout.n500 VGND 0.04919f
C9872 Iout.n501 VGND 0.02502f
C9873 Iout.n502 VGND 0.13561f
C9874 Iout.n503 VGND 0.04584f
C9875 Iout.t246 VGND 0.02212f
C9876 Iout.n504 VGND 0.04919f
C9877 Iout.n505 VGND 0.02502f
C9878 Iout.n506 VGND 0.04584f
C9879 Iout.t76 VGND 0.02212f
C9880 Iout.n507 VGND 0.04919f
C9881 Iout.n508 VGND 0.02502f
C9882 Iout.t138 VGND 0.02212f
C9883 Iout.n509 VGND 0.04919f
C9884 Iout.n510 VGND 0.02502f
C9885 Iout.n511 VGND 0.13561f
C9886 Iout.n512 VGND 0.04584f
C9887 Iout.t4 VGND 0.02212f
C9888 Iout.n513 VGND 0.04919f
C9889 Iout.n514 VGND 0.02502f
C9890 Iout.n515 VGND 0.04584f
C9891 Iout.n516 VGND 0.13561f
C9892 Iout.n517 VGND 0.22972f
C9893 Iout.n518 VGND 0.04584f
C9894 Iout.t27 VGND 0.02212f
C9895 Iout.n519 VGND 0.04919f
C9896 Iout.n520 VGND 0.02502f
C9897 Iout.n521 VGND 0.04584f
C9898 Iout.n522 VGND 0.22972f
C9899 Iout.n523 VGND 0.22972f
C9900 Iout.n524 VGND 0.04584f
C9901 Iout.t112 VGND 0.02212f
C9902 Iout.n525 VGND 0.04919f
C9903 Iout.n526 VGND 0.02502f
C9904 Iout.n527 VGND 0.04584f
C9905 Iout.n528 VGND 0.22972f
C9906 Iout.n529 VGND 0.22972f
C9907 Iout.n530 VGND 0.04584f
C9908 Iout.t50 VGND 0.02212f
C9909 Iout.n531 VGND 0.04919f
C9910 Iout.n532 VGND 0.02502f
C9911 Iout.n533 VGND 0.04584f
C9912 Iout.t46 VGND 0.02212f
C9913 Iout.n534 VGND 0.04919f
C9914 Iout.n535 VGND 0.02502f
C9915 Iout.t140 VGND 0.02212f
C9916 Iout.n536 VGND 0.04919f
C9917 Iout.n537 VGND 0.02502f
C9918 Iout.n538 VGND 0.04584f
C9919 Iout.n539 VGND 0.22972f
C9920 Iout.n540 VGND 0.22972f
C9921 Iout.n541 VGND 0.04584f
C9922 Iout.t209 VGND 0.02212f
C9923 Iout.n542 VGND 0.04919f
C9924 Iout.n543 VGND 0.02502f
C9925 Iout.n544 VGND 0.04584f
C9926 Iout.n545 VGND 0.22972f
C9927 Iout.n546 VGND 0.22972f
C9928 Iout.n547 VGND 0.04584f
C9929 Iout.t242 VGND 0.02212f
C9930 Iout.n548 VGND 0.04919f
C9931 Iout.n549 VGND 0.02502f
C9932 Iout.n550 VGND 0.04584f
C9933 Iout.n551 VGND 0.22972f
C9934 Iout.n552 VGND 0.22972f
C9935 Iout.n553 VGND 0.04584f
C9936 Iout.t53 VGND 0.02212f
C9937 Iout.n554 VGND 0.04919f
C9938 Iout.n555 VGND 0.02502f
C9939 Iout.n556 VGND 0.04584f
C9940 Iout.t119 VGND 0.02212f
C9941 Iout.n557 VGND 0.04919f
C9942 Iout.n558 VGND 0.02502f
C9943 Iout.t220 VGND 0.02212f
C9944 Iout.n559 VGND 0.04919f
C9945 Iout.n560 VGND 0.02502f
C9946 Iout.n561 VGND 0.04584f
C9947 Iout.n562 VGND 0.22972f
C9948 Iout.t92 VGND 0.02212f
C9949 Iout.n563 VGND 0.04919f
C9950 Iout.n564 VGND 0.02502f
C9951 Iout.n565 VGND 0.04584f
C9952 Iout.n566 VGND 0.22972f
C9953 Iout.n567 VGND 0.22972f
C9954 Iout.n568 VGND 0.04584f
C9955 Iout.t24 VGND 0.02212f
C9956 Iout.n569 VGND 0.04919f
C9957 Iout.n570 VGND 0.02502f
C9958 Iout.n571 VGND 0.04584f
C9959 Iout.n572 VGND 0.22972f
C9960 Iout.t16 VGND 0.02212f
C9961 Iout.n573 VGND 0.04919f
C9962 Iout.n574 VGND 0.02502f
C9963 Iout.n575 VGND 0.04584f
C9964 Iout.t193 VGND 0.02212f
C9965 Iout.n576 VGND 0.04919f
C9966 Iout.n577 VGND 0.02502f
C9967 Iout.n578 VGND 0.04584f
C9968 Iout.n579 VGND 0.22972f
C9969 Iout.n580 VGND 0.22972f
C9970 Iout.n581 VGND 0.04584f
C9971 Iout.t181 VGND 0.02212f
C9972 Iout.n582 VGND 0.04919f
C9973 Iout.n583 VGND 0.02502f
C9974 Iout.n584 VGND 0.04584f
C9975 Iout.n585 VGND 0.22972f
C9976 Iout.n586 VGND 0.22972f
C9977 Iout.n587 VGND 0.04584f
C9978 Iout.t40 VGND 0.02212f
C9979 Iout.n588 VGND 0.04919f
C9980 Iout.n589 VGND 0.02502f
C9981 Iout.n590 VGND 0.04584f
C9982 Iout.n591 VGND 0.22972f
C9983 Iout.n592 VGND 0.22972f
C9984 Iout.n593 VGND 0.04584f
C9985 Iout.t127 VGND 0.02212f
C9986 Iout.n594 VGND 0.04919f
C9987 Iout.n595 VGND 0.02502f
C9988 Iout.n596 VGND 0.04584f
C9989 Iout.n597 VGND 0.22972f
C9990 Iout.n598 VGND 0.22972f
C9991 Iout.n599 VGND 0.04584f
C9992 Iout.t172 VGND 0.02212f
C9993 Iout.n600 VGND 0.04919f
C9994 Iout.n601 VGND 0.02502f
C9995 Iout.n602 VGND 0.04584f
C9996 Iout.n603 VGND 0.22972f
C9997 Iout.n604 VGND 0.22972f
C9998 Iout.n605 VGND 0.04584f
C9999 Iout.t147 VGND 0.02212f
C10000 Iout.n606 VGND 0.04919f
C10001 Iout.n607 VGND 0.02502f
C10002 Iout.n608 VGND 0.04584f
C10003 Iout.n609 VGND 0.22972f
C10004 Iout.n610 VGND 0.22972f
C10005 Iout.n611 VGND 0.04584f
C10006 Iout.t173 VGND 0.02212f
C10007 Iout.n612 VGND 0.04919f
C10008 Iout.n613 VGND 0.02502f
C10009 Iout.n614 VGND 0.04584f
C10010 Iout.n615 VGND 0.22972f
C10011 Iout.n616 VGND 0.22972f
C10012 Iout.n617 VGND 0.04584f
C10013 Iout.t99 VGND 0.02212f
C10014 Iout.n618 VGND 0.04919f
C10015 Iout.n619 VGND 0.02502f
C10016 Iout.n620 VGND 0.04584f
C10017 Iout.n621 VGND 0.22972f
C10018 Iout.n622 VGND 0.22972f
C10019 Iout.n623 VGND 0.04584f
C10020 Iout.t255 VGND 0.02212f
C10021 Iout.n624 VGND 0.04919f
C10022 Iout.n625 VGND 0.02502f
C10023 Iout.n626 VGND 0.04584f
C10024 Iout.n627 VGND 0.22972f
C10025 Iout.n628 VGND 0.22972f
C10026 Iout.n629 VGND 0.04584f
C10027 Iout.t248 VGND 0.02212f
C10028 Iout.n630 VGND 0.04919f
C10029 Iout.n631 VGND 0.02502f
C10030 Iout.n632 VGND 0.04584f
C10031 Iout.n633 VGND 0.22972f
C10032 Iout.n634 VGND 0.22972f
C10033 Iout.n635 VGND 0.04584f
C10034 Iout.t64 VGND 0.02212f
C10035 Iout.n636 VGND 0.04919f
C10036 Iout.n637 VGND 0.02502f
C10037 Iout.n638 VGND 0.04584f
C10038 Iout.n639 VGND 0.22972f
C10039 Iout.n640 VGND 0.22972f
C10040 Iout.n641 VGND 0.04584f
C10041 Iout.t237 VGND 0.02212f
C10042 Iout.n642 VGND 0.04919f
C10043 Iout.n643 VGND 0.02502f
C10044 Iout.n644 VGND 0.04584f
C10045 Iout.n645 VGND 0.22972f
C10046 Iout.n646 VGND 0.22972f
C10047 Iout.n647 VGND 0.04584f
C10048 Iout.t34 VGND 0.02212f
C10049 Iout.n648 VGND 0.04919f
C10050 Iout.n649 VGND 0.02502f
C10051 Iout.n650 VGND 0.04584f
C10052 Iout.n651 VGND 0.22972f
C10053 Iout.n652 VGND 0.22972f
C10054 Iout.n653 VGND 0.04584f
C10055 Iout.t211 VGND 0.02212f
C10056 Iout.n654 VGND 0.04919f
C10057 Iout.n655 VGND 0.02502f
C10058 Iout.n656 VGND 0.04584f
C10059 Iout.t87 VGND 0.02212f
C10060 Iout.n657 VGND 0.04919f
C10061 Iout.n658 VGND 0.02502f
C10062 Iout.n659 VGND 0.04584f
C10063 Iout.t95 VGND 0.02212f
C10064 Iout.n660 VGND 0.04919f
C10065 Iout.n661 VGND 0.02502f
C10066 Iout.n662 VGND 0.04584f
C10067 Iout.t23 VGND 0.02212f
C10068 Iout.n663 VGND 0.04919f
C10069 Iout.n664 VGND 0.02502f
C10070 Iout.n665 VGND 0.04584f
C10071 Iout.t83 VGND 0.02212f
C10072 Iout.n666 VGND 0.04919f
C10073 Iout.n667 VGND 0.02502f
C10074 Iout.n668 VGND 0.04584f
C10075 Iout.t214 VGND 0.02212f
C10076 Iout.n669 VGND 0.04919f
C10077 Iout.n670 VGND 0.02502f
C10078 Iout.n671 VGND 0.04584f
C10079 Iout.t160 VGND 0.02212f
C10080 Iout.n672 VGND 0.04919f
C10081 Iout.n673 VGND 0.02502f
C10082 Iout.n674 VGND 0.04584f
C10083 Iout.t151 VGND 0.02212f
C10084 Iout.n675 VGND 0.04919f
C10085 Iout.n676 VGND 0.02502f
C10086 Iout.n677 VGND 0.04584f
C10087 Iout.t213 VGND 0.02212f
C10088 Iout.n678 VGND 0.04919f
C10089 Iout.n679 VGND 0.02502f
C10090 Iout.n680 VGND 0.04584f
C10091 Iout.t15 VGND 0.02212f
C10092 Iout.n681 VGND 0.04919f
C10093 Iout.n682 VGND 0.02502f
C10094 Iout.n683 VGND 0.04584f
C10095 Iout.t10 VGND 0.02212f
C10096 Iout.n684 VGND 0.04919f
C10097 Iout.n685 VGND 0.02502f
C10098 Iout.n686 VGND 0.04584f
C10099 Iout.t36 VGND 0.02212f
C10100 Iout.n687 VGND 0.04919f
C10101 Iout.n688 VGND 0.02502f
C10102 Iout.n689 VGND 0.04584f
C10103 Iout.t25 VGND 0.02212f
C10104 Iout.n690 VGND 0.04919f
C10105 Iout.n691 VGND 0.02502f
C10106 Iout.t179 VGND 0.02212f
C10107 Iout.n692 VGND 0.04919f
C10108 Iout.n693 VGND 0.02502f
C10109 Iout.n694 VGND 0.04584f
C10110 Iout.t163 VGND 0.02212f
C10111 Iout.n695 VGND 0.04919f
C10112 Iout.n696 VGND 0.02502f
C10113 Iout.n697 VGND 0.04584f
C10114 Iout.n698 VGND 0.22972f
C10115 Iout.t226 VGND 0.02212f
C10116 Iout.n699 VGND 0.04919f
C10117 Iout.n700 VGND 0.02502f
C10118 Iout.n701 VGND 0.04584f
C10119 Iout.n702 VGND 0.22972f
C10120 Iout.n703 VGND 0.22972f
C10121 Iout.n704 VGND 0.04584f
C10122 Iout.t190 VGND 0.02212f
C10123 Iout.n705 VGND 0.04919f
C10124 Iout.n706 VGND 0.02502f
C10125 Iout.n707 VGND 0.04584f
C10126 Iout.n708 VGND 0.22972f
C10127 Iout.n709 VGND 0.22972f
C10128 Iout.n710 VGND 0.04584f
C10129 Iout.t161 VGND 0.02212f
C10130 Iout.n711 VGND 0.04919f
C10131 Iout.n712 VGND 0.02502f
C10132 Iout.n713 VGND 0.04584f
C10133 Iout.n714 VGND 0.22972f
C10134 Iout.n715 VGND 0.22972f
C10135 Iout.n716 VGND 0.04584f
C10136 Iout.t132 VGND 0.02212f
C10137 Iout.n717 VGND 0.04919f
C10138 Iout.n718 VGND 0.02502f
C10139 Iout.n719 VGND 0.04584f
C10140 Iout.n720 VGND 0.22972f
C10141 Iout.n721 VGND 0.22972f
C10142 Iout.n722 VGND 0.04584f
C10143 Iout.t13 VGND 0.02212f
C10144 Iout.n723 VGND 0.04919f
C10145 Iout.n724 VGND 0.02502f
C10146 Iout.n725 VGND 0.04584f
C10147 Iout.n726 VGND 0.22972f
C10148 Iout.n727 VGND 0.22972f
C10149 Iout.n728 VGND 0.04584f
C10150 Iout.t204 VGND 0.02212f
C10151 Iout.n729 VGND 0.04919f
C10152 Iout.n730 VGND 0.02502f
C10153 Iout.n731 VGND 0.04584f
C10154 Iout.n732 VGND 0.22972f
C10155 Iout.n733 VGND 0.22972f
C10156 Iout.n734 VGND 0.04584f
C10157 Iout.t48 VGND 0.02212f
C10158 Iout.n735 VGND 0.04919f
C10159 Iout.n736 VGND 0.02502f
C10160 Iout.n737 VGND 0.04584f
C10161 Iout.n738 VGND 0.22972f
C10162 Iout.n739 VGND 0.22972f
C10163 Iout.n740 VGND 0.04584f
C10164 Iout.t114 VGND 0.02212f
C10165 Iout.n741 VGND 0.04919f
C10166 Iout.n742 VGND 0.02502f
C10167 Iout.n743 VGND 0.04584f
C10168 Iout.n744 VGND 0.22972f
C10169 Iout.n745 VGND 0.22972f
C10170 Iout.n746 VGND 0.04584f
C10171 Iout.t66 VGND 0.02212f
C10172 Iout.n747 VGND 0.04919f
C10173 Iout.n748 VGND 0.02502f
C10174 Iout.n749 VGND 0.04584f
C10175 Iout.n750 VGND 0.22972f
C10176 Iout.n751 VGND 0.22972f
C10177 Iout.n752 VGND 0.04584f
C10178 Iout.t184 VGND 0.02212f
C10179 Iout.n753 VGND 0.04919f
C10180 Iout.n754 VGND 0.02502f
C10181 Iout.n755 VGND 0.04584f
C10182 Iout.n756 VGND 0.22972f
C10183 Iout.n757 VGND 0.22972f
C10184 Iout.n758 VGND 0.04584f
C10185 Iout.t33 VGND 0.02212f
C10186 Iout.n759 VGND 0.04919f
C10187 Iout.n760 VGND 0.02502f
C10188 Iout.n761 VGND 0.04584f
C10189 Iout.n762 VGND 0.22972f
C10190 Iout.n763 VGND 0.22972f
C10191 Iout.n764 VGND 0.04584f
C10192 Iout.t71 VGND 0.02212f
C10193 Iout.n765 VGND 0.04919f
C10194 Iout.n766 VGND 0.02502f
C10195 Iout.n767 VGND 0.04584f
C10196 Iout.n768 VGND 0.22972f
C10197 Iout.n769 VGND 0.22972f
C10198 Iout.n770 VGND 0.04584f
C10199 Iout.t219 VGND 0.02212f
C10200 Iout.n771 VGND 0.04919f
C10201 Iout.n772 VGND 0.02502f
C10202 Iout.n773 VGND 0.04584f
C10203 Iout.n774 VGND 0.22972f
C10204 Iout.n775 VGND 0.22972f
C10205 Iout.n776 VGND 0.04584f
C10206 Iout.t201 VGND 0.02212f
C10207 Iout.n777 VGND 0.04919f
C10208 Iout.n778 VGND 0.02502f
C10209 Iout.n779 VGND 0.04584f
C10210 Iout.n780 VGND 0.22972f
C10211 Iout.t228 VGND 0.02212f
C10212 Iout.n781 VGND 0.04919f
C10213 Iout.n782 VGND 0.02502f
C10214 Iout.n783 VGND 0.04584f
C10215 Iout.t142 VGND 0.02212f
C10216 Iout.n784 VGND 0.04919f
C10217 Iout.n785 VGND 0.02502f
C10218 Iout.n786 VGND 0.04584f
C10219 Iout.t245 VGND 0.02212f
C10220 Iout.n787 VGND 0.04919f
C10221 Iout.n788 VGND 0.02502f
C10222 Iout.n789 VGND 0.04584f
C10223 Iout.t146 VGND 0.02212f
C10224 Iout.n790 VGND 0.04919f
C10225 Iout.n791 VGND 0.02502f
C10226 Iout.n792 VGND 0.04584f
C10227 Iout.t231 VGND 0.02212f
C10228 Iout.n793 VGND 0.04919f
C10229 Iout.n794 VGND 0.02502f
C10230 Iout.n795 VGND 0.04584f
C10231 Iout.t155 VGND 0.02212f
C10232 Iout.n796 VGND 0.04919f
C10233 Iout.n797 VGND 0.02502f
C10234 Iout.n798 VGND 0.04584f
C10235 Iout.t100 VGND 0.02212f
C10236 Iout.n799 VGND 0.04919f
C10237 Iout.n800 VGND 0.02502f
C10238 Iout.n801 VGND 0.04584f
C10239 Iout.t26 VGND 0.02212f
C10240 Iout.n802 VGND 0.04919f
C10241 Iout.n803 VGND 0.02502f
C10242 Iout.n804 VGND 0.04584f
C10243 Iout.t183 VGND 0.02212f
C10244 Iout.n805 VGND 0.04919f
C10245 Iout.n806 VGND 0.02502f
C10246 Iout.n807 VGND 0.04584f
C10247 Iout.t195 VGND 0.02212f
C10248 Iout.n808 VGND 0.04919f
C10249 Iout.n809 VGND 0.02502f
C10250 Iout.n810 VGND 0.04584f
C10251 Iout.t162 VGND 0.02212f
C10252 Iout.n811 VGND 0.04919f
C10253 Iout.n812 VGND 0.02502f
C10254 Iout.n813 VGND 0.04584f
C10255 Iout.t73 VGND 0.02212f
C10256 Iout.n814 VGND 0.04919f
C10257 Iout.n815 VGND 0.02502f
C10258 Iout.n816 VGND 0.04584f
C10259 Iout.t49 VGND 0.02212f
C10260 Iout.n817 VGND 0.04919f
C10261 Iout.n818 VGND 0.02502f
C10262 Iout.n819 VGND 0.04584f
C10263 Iout.t69 VGND 0.02212f
C10264 Iout.n820 VGND 0.04919f
C10265 Iout.n821 VGND 0.02502f
C10266 Iout.n822 VGND 0.04584f
C10267 Iout.t174 VGND 0.02212f
C10268 Iout.n823 VGND 0.04919f
C10269 Iout.n824 VGND 0.02502f
C10270 Iout.n825 VGND 0.04584f
C10271 Iout.n826 VGND 0.22972f
C10272 Iout.t182 VGND 0.02212f
C10273 Iout.n827 VGND 0.04919f
C10274 Iout.n828 VGND 0.02502f
C10275 Iout.n829 VGND 0.07841f
C10276 Iout.n830 VGND 0.47625f
C10277 Iout.n831 VGND 0.04584f
C10278 Iout.t205 VGND 0.02212f
C10279 Iout.n832 VGND 0.04919f
C10280 Iout.n833 VGND 0.02502f
C10281 Iout.t60 VGND 0.02212f
C10282 Iout.n834 VGND 0.04919f
C10283 Iout.n835 VGND 0.02502f
C10284 Iout.n836 VGND 0.04584f
C10285 Iout.n837 VGND 0.47625f
C10286 Iout.n838 VGND 0.07841f
C10287 Iout.t128 VGND 0.02212f
C10288 Iout.n839 VGND 0.04919f
C10289 Iout.n840 VGND 0.02502f
C10290 Iout.t197 VGND 0.02212f
C10291 Iout.n841 VGND 0.04919f
C10292 Iout.n842 VGND 0.02502f
C10293 Iout.n843 VGND 0.07841f
C10294 Iout.n844 VGND 0.47625f
C10295 Iout.n845 VGND 0.04584f
C10296 Iout.t96 VGND 0.02212f
C10297 Iout.n846 VGND 0.04919f
C10298 Iout.n847 VGND 0.02502f
C10299 Iout.t166 VGND 0.02212f
C10300 Iout.n848 VGND 0.04919f
C10301 Iout.n849 VGND 0.02502f
C10302 Iout.n850 VGND 0.04584f
C10303 Iout.n851 VGND 0.47625f
C10304 Iout.n852 VGND 0.07841f
C10305 Iout.t135 VGND 0.02212f
C10306 Iout.n853 VGND 0.04919f
C10307 Iout.n854 VGND 0.02502f
C10308 Iout.t158 VGND 0.02212f
C10309 Iout.n855 VGND 0.04919f
C10310 Iout.n856 VGND 0.02502f
C10311 Iout.n857 VGND 0.07841f
C10312 Iout.n858 VGND 0.47625f
C10313 Iout.n859 VGND 0.04584f
C10314 Iout.t31 VGND 0.02212f
C10315 Iout.n860 VGND 0.04919f
C10316 Iout.n861 VGND 0.02502f
C10317 Iout.t107 VGND 0.02212f
C10318 Iout.n862 VGND 0.04919f
C10319 Iout.n863 VGND 0.02502f
C10320 Iout.n864 VGND 0.04584f
C10321 Iout.n865 VGND 0.47625f
C10322 Iout.n866 VGND 0.07841f
C10323 Iout.t252 VGND 0.02212f
C10324 Iout.n867 VGND 0.04919f
C10325 Iout.n868 VGND 0.02502f
C10326 Iout.t35 VGND 0.02212f
C10327 Iout.n869 VGND 0.04919f
C10328 Iout.n870 VGND 0.02502f
C10329 Iout.n871 VGND 0.07841f
C10330 Iout.n872 VGND 0.47625f
C10331 Iout.n873 VGND 0.04584f
C10332 Iout.t249 VGND 0.02212f
C10333 Iout.n874 VGND 0.04919f
C10334 Iout.n875 VGND 0.02502f
C10335 Iout.t108 VGND 0.02212f
C10336 Iout.n876 VGND 0.04919f
C10337 Iout.n877 VGND 0.02502f
C10338 Iout.n878 VGND 0.04584f
C10339 Iout.n879 VGND 0.47625f
C10340 Iout.n880 VGND 0.07841f
C10341 Iout.t238 VGND 0.02212f
C10342 Iout.n881 VGND 0.04919f
C10343 Iout.n882 VGND 0.02502f
C10344 Iout.t2 VGND 0.02212f
C10345 Iout.n883 VGND 0.04919f
C10346 Iout.n884 VGND 0.02502f
C10347 Iout.n885 VGND 0.07841f
C10348 Iout.n886 VGND 0.47625f
C10349 Iout.n887 VGND 0.04584f
C10350 Iout.t243 VGND 0.02212f
C10351 Iout.n888 VGND 0.04919f
C10352 Iout.n889 VGND 0.02502f
C10353 Iout.t225 VGND 0.02212f
C10354 Iout.n890 VGND 0.04919f
C10355 Iout.n891 VGND 0.02502f
C10356 Iout.n892 VGND 0.04584f
C10357 Iout.n893 VGND 0.47625f
C10358 Iout.n894 VGND 0.07841f
C10359 Iout.t216 VGND 0.02212f
C10360 Iout.n895 VGND 0.04919f
C10361 Iout.n896 VGND 0.02502f
C10362 Iout.t113 VGND 0.02212f
C10363 Iout.n897 VGND 0.04919f
C10364 Iout.n898 VGND 0.02502f
C10365 Iout.n899 VGND 0.07841f
C10366 Iout.n900 VGND 0.47625f
C10367 Iout.n901 VGND 0.04584f
C10368 Iout.t86 VGND 0.02212f
C10369 Iout.n902 VGND 0.04919f
C10370 Iout.n903 VGND 0.02502f
C10371 Iout.t148 VGND 0.02212f
C10372 Iout.n904 VGND 0.04919f
C10373 Iout.n905 VGND 0.02502f
C10374 Iout.n906 VGND 0.04584f
C10375 Iout.n907 VGND 0.47625f
C10376 Iout.n908 VGND 0.07841f
C10377 Iout.t244 VGND 0.02212f
C10378 Iout.n909 VGND 0.04919f
C10379 Iout.n910 VGND 0.02502f
C10380 Iout.t68 VGND 0.02212f
C10381 Iout.n911 VGND 0.04919f
C10382 Iout.n912 VGND 0.02502f
C10383 Iout.n913 VGND 0.07841f
C10384 Iout.n914 VGND 0.47625f
C10385 Iout.n915 VGND 0.04584f
C10386 Iout.t167 VGND 0.02212f
C10387 Iout.n916 VGND 0.04919f
C10388 Iout.n917 VGND 0.02502f
C10389 Iout.t12 VGND 0.02212f
C10390 Iout.n918 VGND 0.04919f
C10391 Iout.n919 VGND 0.02502f
C10392 Iout.n920 VGND 0.04584f
C10393 Iout.n921 VGND 0.47625f
C10394 Iout.n922 VGND 0.07841f
C10395 Iout.t80 VGND 0.02212f
C10396 Iout.n923 VGND 0.04919f
C10397 Iout.n924 VGND 0.02502f
C10398 Iout.n925 VGND 0.07841f
C10399 Iout.t124 VGND 0.02212f
C10400 Iout.n926 VGND 0.04919f
C10401 Iout.n927 VGND 0.02502f
C10402 Iout.n928 VGND 0.07841f
C10403 Iout.n929 VGND 0.47625f
C10404 Iout.n930 VGND 0.04584f
C10405 Iout.t1 VGND 0.02212f
C10406 Iout.n931 VGND 0.04919f
C10407 Iout.n932 VGND 0.02502f
C10408 Iout.n933 VGND 0.04584f
C10409 Iout.t17 VGND 0.02212f
C10410 Iout.n934 VGND 0.04919f
C10411 Iout.n935 VGND 0.19431f
C10412 Iout.n936 VGND 2.54526f
C10413 Iout.n937 VGND 1.20114f
C10414 Iout.t79 VGND 0.02212f
C10415 Iout.n938 VGND 0.04919f
C10416 Iout.n939 VGND 0.19431f
C10417 Iout.n940 VGND 0.04584f
C10418 Iout.n941 VGND 0.22972f
C10419 Iout.n942 VGND 0.22972f
C10420 Iout.n943 VGND 0.04584f
C10421 Iout.t54 VGND 0.02212f
C10422 Iout.n944 VGND 0.04919f
C10423 Iout.n945 VGND 0.02502f
C10424 Iout.n946 VGND 0.04584f
C10425 Iout.n947 VGND 0.22972f
C10426 Iout.n948 VGND 0.22972f
C10427 Iout.n949 VGND 0.04584f
C10428 Iout.t198 VGND 0.02212f
C10429 Iout.n950 VGND 0.04919f
C10430 Iout.n951 VGND 0.02502f
C10431 Iout.n952 VGND 0.04584f
C10432 Iout.t224 VGND 0.02212f
C10433 Iout.n953 VGND 0.04919f
C10434 Iout.n954 VGND 0.19431f
C10435 Iout.n955 VGND 1.20114f
C10436 Iout.n956 VGND 1.20114f
C10437 Iout.t42 VGND 0.02212f
C10438 Iout.n957 VGND 0.04919f
C10439 Iout.n958 VGND 0.19431f
C10440 Iout.n959 VGND 0.04584f
C10441 Iout.n960 VGND 0.22972f
C10442 Iout.n961 VGND 0.22972f
C10443 Iout.n962 VGND 0.04584f
C10444 Iout.t97 VGND 0.02212f
C10445 Iout.n963 VGND 0.04919f
C10446 Iout.n964 VGND 0.02502f
C10447 Iout.n965 VGND 0.04584f
C10448 Iout.n966 VGND 0.22972f
C10449 Iout.n967 VGND 0.22972f
C10450 Iout.n968 VGND 0.04584f
C10451 Iout.t236 VGND 0.02212f
C10452 Iout.n969 VGND 0.04919f
C10453 Iout.n970 VGND 0.02502f
C10454 Iout.n971 VGND 0.04584f
C10455 Iout.t145 VGND 0.02212f
C10456 Iout.n972 VGND 0.04919f
C10457 Iout.n973 VGND 0.19431f
C10458 Iout.n974 VGND 1.20114f
C10459 Iout.n975 VGND 1.20114f
C10460 Iout.t106 VGND 0.02212f
C10461 Iout.n976 VGND 0.04919f
C10462 Iout.n977 VGND 0.19431f
C10463 Iout.n978 VGND 0.04584f
C10464 Iout.n979 VGND 0.22972f
C10465 Iout.n980 VGND 0.22972f
C10466 Iout.n981 VGND 0.04584f
C10467 Iout.t137 VGND 0.02212f
C10468 Iout.n982 VGND 0.04919f
C10469 Iout.n983 VGND 0.02502f
C10470 Iout.n984 VGND 0.04584f
C10471 Iout.n985 VGND 0.22972f
C10472 Iout.n986 VGND 0.22972f
C10473 Iout.n987 VGND 0.04584f
C10474 Iout.t85 VGND 0.02212f
C10475 Iout.n988 VGND 0.04919f
C10476 Iout.n989 VGND 0.02502f
C10477 Iout.n990 VGND 0.04584f
C10478 Iout.t125 VGND 0.02212f
C10479 Iout.n991 VGND 0.04919f
C10480 Iout.n992 VGND 0.19431f
C10481 Iout.n993 VGND 1.20114f
C10482 Iout.n994 VGND 1.20114f
C10483 Iout.t21 VGND 0.02212f
C10484 Iout.n995 VGND 0.04919f
C10485 Iout.n996 VGND 0.19431f
C10486 Iout.n997 VGND 0.04584f
C10487 Iout.n998 VGND 0.22972f
C10488 Iout.n999 VGND 0.22972f
C10489 Iout.n1000 VGND 0.04584f
C10490 Iout.t186 VGND 0.02212f
C10491 Iout.n1001 VGND 0.04919f
C10492 Iout.n1002 VGND 0.02502f
C10493 Iout.n1003 VGND 0.04584f
C10494 Iout.n1004 VGND 0.22972f
C10495 Iout.n1005 VGND 0.22972f
C10496 Iout.n1006 VGND 0.04584f
C10497 Iout.t67 VGND 0.02212f
C10498 Iout.n1007 VGND 0.04919f
C10499 Iout.n1008 VGND 0.02502f
C10500 Iout.n1009 VGND 0.04584f
C10501 Iout.t105 VGND 0.02212f
C10502 Iout.n1010 VGND 0.04919f
C10503 Iout.n1011 VGND 0.19431f
C10504 Iout.n1012 VGND 1.20114f
C10505 Iout.n1013 VGND 1.07853f
C10506 Iout.t37 VGND 0.02212f
C10507 Iout.n1014 VGND 0.04919f
C10508 Iout.n1015 VGND 0.19431f
C10509 Iout.n1016 VGND 0.04584f
C10510 Iout.n1017 VGND 0.22972f
C10511 Iout.n1018 VGND 0.13561f
C10512 Iout.n1019 VGND 0.04584f
C10513 Iout.t222 VGND 0.02212f
C10514 Iout.n1020 VGND 0.04919f
C10515 Iout.n1021 VGND 0.19431f
C10516 Iout.n1022 VGND 0.22314f
C10517 VPWR.n0 VGND 0.03466f
C10518 VPWR.t1837 VGND 0.21918f
C10519 VPWR.t1126 VGND 0.09699f
C10520 VPWR.t387 VGND 0.27964f
C10521 VPWR.t366 VGND 0.10581f
C10522 VPWR.t1759 VGND 0.10581f
C10523 VPWR.t1325 VGND 0.10581f
C10524 VPWR.t140 VGND 0.10581f
C10525 VPWR.t262 VGND 0.10581f
C10526 VPWR.t258 VGND 0.10581f
C10527 VPWR.t1727 VGND 0.07432f
C10528 VPWR.n1 VGND 0.13503f
C10529 VPWR.n2 VGND 0.07145f
C10530 VPWR.t1127 VGND 0.04227f
C10531 VPWR.t1728 VGND 0.0106f
C10532 VPWR.t259 VGND 0.0106f
C10533 VPWR.n4 VGND 0.02326f
C10534 VPWR.t263 VGND 0.0106f
C10535 VPWR.t141 VGND 0.0106f
C10536 VPWR.n5 VGND 0.02322f
C10537 VPWR.n6 VGND 0.0477f
C10538 VPWR.n7 VGND 0.13446f
C10539 VPWR.n8 VGND 0.04257f
C10540 VPWR.n9 VGND 0.03127f
C10541 VPWR.n10 VGND 0.05604f
C10542 VPWR.n12 VGND 0.01206f
C10543 VPWR.n13 VGND 0.01413f
C10544 VPWR.n14 VGND 0.02072f
C10545 VPWR.n15 VGND 0.06272f
C10546 VPWR.t1838 VGND 0.04226f
C10547 VPWR.n17 VGND 0.05435f
C10548 VPWR.n18 VGND 0.2482f
C10549 VPWR.n19 VGND 0.72374f
C10550 VPWR.n20 VGND 0.23558f
C10551 VPWR.n21 VGND 0.75117f
C10552 VPWR.n22 VGND 0.1027f
C10553 VPWR.n23 VGND 0.02214f
C10554 VPWR.n24 VGND 0.05881f
C10555 VPWR.n25 VGND 0.02214f
C10556 VPWR.n26 VGND 0.11837f
C10557 VPWR.n27 VGND 0.02214f
C10558 VPWR.n28 VGND 0.09431f
C10559 VPWR.n29 VGND 0.02214f
C10560 VPWR.n30 VGND 0.09431f
C10561 VPWR.n31 VGND 0.02214f
C10562 VPWR.n32 VGND 0.09431f
C10563 VPWR.n33 VGND 0.02214f
C10564 VPWR.n34 VGND 0.09431f
C10565 VPWR.n35 VGND 0.02214f
C10566 VPWR.n36 VGND 0.09431f
C10567 VPWR.n37 VGND 0.02214f
C10568 VPWR.n38 VGND 0.09431f
C10569 VPWR.n39 VGND 0.02214f
C10570 VPWR.n40 VGND 0.09431f
C10571 VPWR.n41 VGND 0.02214f
C10572 VPWR.n42 VGND 0.09431f
C10573 VPWR.n43 VGND 0.02214f
C10574 VPWR.n44 VGND 0.09431f
C10575 VPWR.n45 VGND 0.02214f
C10576 VPWR.n46 VGND 0.09431f
C10577 VPWR.n47 VGND 0.02214f
C10578 VPWR.n48 VGND 0.09431f
C10579 VPWR.n49 VGND 0.02214f
C10580 VPWR.n50 VGND 0.09431f
C10581 VPWR.n51 VGND 0.02214f
C10582 VPWR.n52 VGND 0.09431f
C10583 VPWR.n53 VGND 0.02214f
C10584 VPWR.n54 VGND 0.10211f
C10585 VPWR.n55 VGND 0.08525f
C10586 VPWR.t711 VGND 0.02464f
C10587 VPWR.t816 VGND 0.02189f
C10588 VPWR.n56 VGND 0.06768f
C10589 VPWR.t579 VGND 0.06817f
C10590 VPWR.t586 VGND 0.02464f
C10591 VPWR.t580 VGND 0.02189f
C10592 VPWR.n57 VGND 0.06768f
C10593 VPWR.n58 VGND 0.02542f
C10594 VPWR.n59 VGND 0.10289f
C10595 VPWR.n60 VGND 0.10289f
C10596 VPWR.n61 VGND 0.02542f
C10597 VPWR.t567 VGND 0.02464f
C10598 VPWR.t940 VGND 0.02189f
C10599 VPWR.n62 VGND 0.06768f
C10600 VPWR.t806 VGND 0.06817f
C10601 VPWR.t717 VGND 0.02464f
C10602 VPWR.t807 VGND 0.02189f
C10603 VPWR.n63 VGND 0.06768f
C10604 VPWR.n64 VGND 0.02542f
C10605 VPWR.n65 VGND 0.10289f
C10606 VPWR.n66 VGND 0.10289f
C10607 VPWR.n67 VGND 0.02542f
C10608 VPWR.t687 VGND 0.02464f
C10609 VPWR.t679 VGND 0.02189f
C10610 VPWR.n68 VGND 0.06768f
C10611 VPWR.t660 VGND 0.06817f
C10612 VPWR.t943 VGND 0.02464f
C10613 VPWR.t661 VGND 0.02189f
C10614 VPWR.n69 VGND 0.06768f
C10615 VPWR.n70 VGND 0.02542f
C10616 VPWR.n71 VGND 0.10289f
C10617 VPWR.n72 VGND 0.10289f
C10618 VPWR.n73 VGND 0.02542f
C10619 VPWR.t813 VGND 0.02464f
C10620 VPWR.t894 VGND 0.02189f
C10621 VPWR.n74 VGND 0.06768f
C10622 VPWR.t783 VGND 0.06817f
C10623 VPWR.t797 VGND 0.02464f
C10624 VPWR.t784 VGND 0.02189f
C10625 VPWR.n75 VGND 0.06768f
C10626 VPWR.n76 VGND 0.02542f
C10627 VPWR.n77 VGND 0.10289f
C10628 VPWR.n78 VGND 0.10289f
C10629 VPWR.n79 VGND 0.02542f
C10630 VPWR.t637 VGND 0.02464f
C10631 VPWR.t656 VGND 0.02189f
C10632 VPWR.n80 VGND 0.06768f
C10633 VPWR.t620 VGND 0.06817f
C10634 VPWR.t916 VGND 0.02464f
C10635 VPWR.t621 VGND 0.02189f
C10636 VPWR.n81 VGND 0.06768f
C10637 VPWR.n82 VGND 0.02542f
C10638 VPWR.n83 VGND 0.10289f
C10639 VPWR.n84 VGND 0.10289f
C10640 VPWR.n85 VGND 0.02542f
C10641 VPWR.t760 VGND 0.02464f
C10642 VPWR.t897 VGND 0.02189f
C10643 VPWR.n86 VGND 0.06768f
C10644 VPWR.t741 VGND 0.06817f
C10645 VPWR.t751 VGND 0.02464f
C10646 VPWR.t742 VGND 0.02189f
C10647 VPWR.n87 VGND 0.06768f
C10648 VPWR.n88 VGND 0.02542f
C10649 VPWR.n89 VGND 0.10289f
C10650 VPWR.n90 VGND 0.10289f
C10651 VPWR.n91 VGND 0.02542f
C10652 VPWR.t640 VGND 0.02464f
C10653 VPWR.t634 VGND 0.02189f
C10654 VPWR.n92 VGND 0.06768f
C10655 VPWR.t871 VGND 0.06817f
C10656 VPWR.t875 VGND 0.02464f
C10657 VPWR.t872 VGND 0.02189f
C10658 VPWR.n93 VGND 0.06768f
C10659 VPWR.n94 VGND 0.02542f
C10660 VPWR.n95 VGND 0.10289f
C10661 VPWR.n96 VGND 0.10289f
C10662 VPWR.n97 VGND 0.02542f
C10663 VPWR.t763 VGND 0.02464f
C10664 VPWR.t854 VGND 0.02189f
C10665 VPWR.n98 VGND 0.06768f
C10666 VPWR.t617 VGND 0.10732f
C10667 VPWR.t593 VGND 0.05805f
C10668 VPWR.t724 VGND 0.06817f
C10669 VPWR.t618 VGND 0.02464f
C10670 VPWR.t725 VGND 0.02189f
C10671 VPWR.n99 VGND 0.06768f
C10672 VPWR.n100 VGND 0.02213f
C10673 VPWR.n101 VGND 0.02429f
C10674 VPWR.n103 VGND 0.01347f
C10675 VPWR.n104 VGND 0.02213f
C10676 VPWR.n105 VGND 0.02429f
C10677 VPWR.n106 VGND 0.02304f
C10678 VPWR.n107 VGND 0.01456f
C10679 VPWR.n108 VGND 0.02047f
C10680 VPWR.n109 VGND 0.02084f
C10681 VPWR.n110 VGND 0.01313f
C10682 VPWR.n112 VGND 0.01347f
C10683 VPWR.n113 VGND 0.01963f
C10684 VPWR.n114 VGND 0.02213f
C10685 VPWR.n115 VGND 0.02429f
C10686 VPWR.n116 VGND 0.02304f
C10687 VPWR.n117 VGND 0.02731f
C10688 VPWR.n119 VGND 0.02047f
C10689 VPWR.n120 VGND 0.02084f
C10690 VPWR.n121 VGND 0.01313f
C10691 VPWR.n123 VGND 0.01347f
C10692 VPWR.n124 VGND 0.01879f
C10693 VPWR.n125 VGND 0.02213f
C10694 VPWR.n126 VGND 0.02429f
C10695 VPWR.n127 VGND 0.02304f
C10696 VPWR.n128 VGND 0.02731f
C10697 VPWR.n130 VGND 0.02047f
C10698 VPWR.n131 VGND 0.02084f
C10699 VPWR.n132 VGND 0.01313f
C10700 VPWR.n134 VGND 0.01347f
C10701 VPWR.n135 VGND 0.01763f
C10702 VPWR.n136 VGND 0.1565f
C10703 VPWR.n137 VGND 0.02213f
C10704 VPWR.n138 VGND 0.02429f
C10705 VPWR.n139 VGND 0.02304f
C10706 VPWR.n140 VGND 0.02731f
C10707 VPWR.n142 VGND 0.02047f
C10708 VPWR.n143 VGND 0.02084f
C10709 VPWR.n144 VGND 0.01313f
C10710 VPWR.n146 VGND 0.01347f
C10711 VPWR.n147 VGND 0.01763f
C10712 VPWR.n148 VGND 0.13004f
C10713 VPWR.n149 VGND 0.02213f
C10714 VPWR.n150 VGND 0.02429f
C10715 VPWR.n151 VGND 0.02304f
C10716 VPWR.n152 VGND 0.02731f
C10717 VPWR.n154 VGND 0.02047f
C10718 VPWR.n155 VGND 0.02084f
C10719 VPWR.n156 VGND 0.01313f
C10720 VPWR.n158 VGND 0.01347f
C10721 VPWR.n159 VGND 0.01763f
C10722 VPWR.n160 VGND 0.13004f
C10723 VPWR.n161 VGND 0.02213f
C10724 VPWR.n162 VGND 0.02429f
C10725 VPWR.n163 VGND 0.02304f
C10726 VPWR.n164 VGND 0.02731f
C10727 VPWR.n166 VGND 0.02047f
C10728 VPWR.n167 VGND 0.02084f
C10729 VPWR.n168 VGND 0.01313f
C10730 VPWR.n170 VGND 0.01347f
C10731 VPWR.n171 VGND 0.01763f
C10732 VPWR.n172 VGND 0.13004f
C10733 VPWR.n173 VGND 0.02213f
C10734 VPWR.n174 VGND 0.02429f
C10735 VPWR.n175 VGND 0.02304f
C10736 VPWR.n176 VGND 0.02731f
C10737 VPWR.n178 VGND 0.02047f
C10738 VPWR.n179 VGND 0.02084f
C10739 VPWR.n180 VGND 0.01313f
C10740 VPWR.n182 VGND 0.01347f
C10741 VPWR.n183 VGND 0.01763f
C10742 VPWR.n184 VGND 0.13004f
C10743 VPWR.n185 VGND 0.02213f
C10744 VPWR.n186 VGND 0.02429f
C10745 VPWR.n187 VGND 0.02304f
C10746 VPWR.n188 VGND 0.02731f
C10747 VPWR.n190 VGND 0.02047f
C10748 VPWR.n191 VGND 0.02084f
C10749 VPWR.n192 VGND 0.01313f
C10750 VPWR.n194 VGND 0.01347f
C10751 VPWR.n195 VGND 0.01763f
C10752 VPWR.n196 VGND 0.13004f
C10753 VPWR.n197 VGND 0.02213f
C10754 VPWR.n198 VGND 0.02429f
C10755 VPWR.n199 VGND 0.02304f
C10756 VPWR.n200 VGND 0.02731f
C10757 VPWR.n202 VGND 0.02047f
C10758 VPWR.n203 VGND 0.02084f
C10759 VPWR.n204 VGND 0.01313f
C10760 VPWR.n206 VGND 0.01347f
C10761 VPWR.n207 VGND 0.01763f
C10762 VPWR.n208 VGND 0.13004f
C10763 VPWR.n209 VGND 0.02213f
C10764 VPWR.n210 VGND 0.02429f
C10765 VPWR.n211 VGND 0.02304f
C10766 VPWR.n212 VGND 0.02731f
C10767 VPWR.n214 VGND 0.02047f
C10768 VPWR.n215 VGND 0.02084f
C10769 VPWR.n216 VGND 0.01313f
C10770 VPWR.n218 VGND 0.01347f
C10771 VPWR.n219 VGND 0.01763f
C10772 VPWR.n220 VGND 0.13004f
C10773 VPWR.n221 VGND 0.02213f
C10774 VPWR.n222 VGND 0.02429f
C10775 VPWR.n223 VGND 0.02304f
C10776 VPWR.n224 VGND 0.02731f
C10777 VPWR.n226 VGND 0.02047f
C10778 VPWR.n227 VGND 0.02084f
C10779 VPWR.n228 VGND 0.01313f
C10780 VPWR.n230 VGND 0.01347f
C10781 VPWR.n231 VGND 0.01763f
C10782 VPWR.n232 VGND 0.13004f
C10783 VPWR.n233 VGND 0.02213f
C10784 VPWR.n234 VGND 0.02429f
C10785 VPWR.n235 VGND 0.02304f
C10786 VPWR.n236 VGND 0.02731f
C10787 VPWR.n238 VGND 0.02047f
C10788 VPWR.n239 VGND 0.02084f
C10789 VPWR.n240 VGND 0.01313f
C10790 VPWR.n242 VGND 0.01347f
C10791 VPWR.n243 VGND 0.01763f
C10792 VPWR.n244 VGND 0.13004f
C10793 VPWR.n245 VGND 0.02213f
C10794 VPWR.n246 VGND 0.02429f
C10795 VPWR.n247 VGND 0.02304f
C10796 VPWR.n248 VGND 0.02731f
C10797 VPWR.n250 VGND 0.02047f
C10798 VPWR.n251 VGND 0.02084f
C10799 VPWR.n252 VGND 0.01313f
C10800 VPWR.n254 VGND 0.01347f
C10801 VPWR.n255 VGND 0.01763f
C10802 VPWR.n256 VGND 0.13004f
C10803 VPWR.n257 VGND 0.02213f
C10804 VPWR.n258 VGND 0.02429f
C10805 VPWR.n259 VGND 0.02304f
C10806 VPWR.n260 VGND 0.02731f
C10807 VPWR.n262 VGND 0.02047f
C10808 VPWR.n263 VGND 0.02084f
C10809 VPWR.n264 VGND 0.01313f
C10810 VPWR.n266 VGND 0.01347f
C10811 VPWR.n267 VGND 0.01763f
C10812 VPWR.n268 VGND 0.13004f
C10813 VPWR.n269 VGND 0.02213f
C10814 VPWR.n270 VGND 0.02429f
C10815 VPWR.n271 VGND 0.02304f
C10816 VPWR.n272 VGND 0.02731f
C10817 VPWR.n274 VGND 0.02047f
C10818 VPWR.n275 VGND 0.02084f
C10819 VPWR.n276 VGND 0.01313f
C10820 VPWR.n278 VGND 0.01347f
C10821 VPWR.n279 VGND 0.01763f
C10822 VPWR.n280 VGND 0.13004f
C10823 VPWR.n281 VGND 0.17544f
C10824 VPWR.n282 VGND 0.01763f
C10825 VPWR.n283 VGND 0.01313f
C10826 VPWR.n284 VGND 0.02047f
C10827 VPWR.n285 VGND 0.02084f
C10828 VPWR.n287 VGND 0.02304f
C10829 VPWR.n288 VGND 0.02731f
C10830 VPWR.n289 VGND 0.02542f
C10831 VPWR.t1464 VGND 0.02464f
C10832 VPWR.t990 VGND 0.02189f
C10833 VPWR.n290 VGND 0.06768f
C10834 VPWR.t1463 VGND 0.10732f
C10835 VPWR.t1253 VGND 0.05805f
C10836 VPWR.t989 VGND 0.06817f
C10837 VPWR.t195 VGND 0.02464f
C10838 VPWR.t924 VGND 0.02189f
C10839 VPWR.n291 VGND 0.06768f
C10840 VPWR.n292 VGND 0.01329f
C10841 VPWR.n293 VGND 0.05634f
C10842 VPWR.t923 VGND 0.0986f
C10843 VPWR.t1591 VGND 0.05805f
C10844 VPWR.t194 VGND 0.08842f
C10845 VPWR.t530 VGND 0.02464f
C10846 VPWR.t1628 VGND 0.02189f
C10847 VPWR.n294 VGND 0.06768f
C10848 VPWR.n295 VGND 0.01329f
C10849 VPWR.n297 VGND 0.08003f
C10850 VPWR.t1627 VGND 0.06817f
C10851 VPWR.t1915 VGND 0.05805f
C10852 VPWR.t529 VGND 0.08842f
C10853 VPWR.t287 VGND 0.02464f
C10854 VPWR.t1427 VGND 0.02189f
C10855 VPWR.n298 VGND 0.06768f
C10856 VPWR.n299 VGND 0.01329f
C10857 VPWR.n301 VGND 0.08003f
C10858 VPWR.t1426 VGND 0.06817f
C10859 VPWR.t1710 VGND 0.05805f
C10860 VPWR.t286 VGND 0.08842f
C10861 VPWR.t38 VGND 0.02464f
C10862 VPWR.t165 VGND 0.02189f
C10863 VPWR.n302 VGND 0.06768f
C10864 VPWR.n303 VGND 0.01329f
C10865 VPWR.n305 VGND 0.08003f
C10866 VPWR.t164 VGND 0.06817f
C10867 VPWR.t1711 VGND 0.05805f
C10868 VPWR.t37 VGND 0.08842f
C10869 VPWR.t1515 VGND 0.02464f
C10870 VPWR.t969 VGND 0.02189f
C10871 VPWR.n306 VGND 0.06768f
C10872 VPWR.n307 VGND 0.01329f
C10873 VPWR.n309 VGND 0.08003f
C10874 VPWR.t968 VGND 0.06817f
C10875 VPWR.t1254 VGND 0.05805f
C10876 VPWR.t1514 VGND 0.08842f
C10877 VPWR.t383 VGND 0.02464f
C10878 VPWR.t1748 VGND 0.02189f
C10879 VPWR.n310 VGND 0.06768f
C10880 VPWR.n311 VGND 0.01329f
C10881 VPWR.n313 VGND 0.08003f
C10882 VPWR.t1747 VGND 0.06817f
C10883 VPWR.t1255 VGND 0.05805f
C10884 VPWR.t382 VGND 0.08842f
C10885 VPWR.t1041 VGND 0.02464f
C10886 VPWR.t408 VGND 0.02189f
C10887 VPWR.n314 VGND 0.06768f
C10888 VPWR.n315 VGND 0.01329f
C10889 VPWR.n317 VGND 0.08003f
C10890 VPWR.t407 VGND 0.06817f
C10891 VPWR.t1589 VGND 0.05805f
C10892 VPWR.t1040 VGND 0.08842f
C10893 VPWR.t273 VGND 0.02464f
C10894 VPWR.t319 VGND 0.02189f
C10895 VPWR.n318 VGND 0.06768f
C10896 VPWR.n319 VGND 0.01329f
C10897 VPWR.n321 VGND 0.08003f
C10898 VPWR.t318 VGND 0.06817f
C10899 VPWR.t1592 VGND 0.05805f
C10900 VPWR.t272 VGND 0.08842f
C10901 VPWR.t1862 VGND 0.02464f
C10902 VPWR.t249 VGND 0.02189f
C10903 VPWR.n322 VGND 0.06768f
C10904 VPWR.n323 VGND 0.01329f
C10905 VPWR.n325 VGND 0.08003f
C10906 VPWR.t248 VGND 0.06817f
C10907 VPWR.t1251 VGND 0.05805f
C10908 VPWR.t1861 VGND 0.08842f
C10909 VPWR.t1483 VGND 0.02464f
C10910 VPWR.t1868 VGND 0.02189f
C10911 VPWR.n326 VGND 0.06768f
C10912 VPWR.n327 VGND 0.01329f
C10913 VPWR.n329 VGND 0.08003f
C10914 VPWR.t1867 VGND 0.06817f
C10915 VPWR.t1587 VGND 0.05805f
C10916 VPWR.t1482 VGND 0.08842f
C10917 VPWR.t1529 VGND 0.02464f
C10918 VPWR.t1258 VGND 0.02189f
C10919 VPWR.n330 VGND 0.06768f
C10920 VPWR.n331 VGND 0.01329f
C10921 VPWR.n333 VGND 0.08003f
C10922 VPWR.t1257 VGND 0.06817f
C10923 VPWR.t1588 VGND 0.05805f
C10924 VPWR.t1528 VGND 0.08842f
C10925 VPWR.t1047 VGND 0.02464f
C10926 VPWR.t112 VGND 0.02189f
C10927 VPWR.n334 VGND 0.06768f
C10928 VPWR.n335 VGND 0.01329f
C10929 VPWR.n337 VGND 0.08003f
C10930 VPWR.t111 VGND 0.06817f
C10931 VPWR.t1252 VGND 0.05805f
C10932 VPWR.t1046 VGND 0.08842f
C10933 VPWR.t1164 VGND 0.02464f
C10934 VPWR.t1081 VGND 0.02189f
C10935 VPWR.n338 VGND 0.06768f
C10936 VPWR.n339 VGND 0.01329f
C10937 VPWR.n341 VGND 0.08003f
C10938 VPWR.t1080 VGND 0.06817f
C10939 VPWR.t1256 VGND 0.05805f
C10940 VPWR.t1163 VGND 0.08842f
C10941 VPWR.t1715 VGND 0.02464f
C10942 VPWR.t1140 VGND 0.02189f
C10943 VPWR.n342 VGND 0.06768f
C10944 VPWR.n343 VGND 0.01329f
C10945 VPWR.n345 VGND 0.08003f
C10946 VPWR.t1139 VGND 0.06817f
C10947 VPWR.t1914 VGND 0.05805f
C10948 VPWR.t1714 VGND 0.08842f
C10949 VPWR.t1622 VGND 0.02464f
C10950 VPWR.t1545 VGND 0.02189f
C10951 VPWR.n346 VGND 0.06768f
C10952 VPWR.n347 VGND 0.01329f
C10953 VPWR.n349 VGND 0.08003f
C10954 VPWR.t1544 VGND 0.06817f
C10955 VPWR.t1590 VGND 0.05805f
C10956 VPWR.t1621 VGND 0.08842f
C10957 VPWR.n350 VGND 0.08003f
C10958 VPWR.n352 VGND 0.01329f
C10959 VPWR.n353 VGND 0.10289f
C10960 VPWR.n354 VGND 0.74646f
C10961 VPWR.n355 VGND 0.10289f
C10962 VPWR.t1458 VGND 0.02464f
C10963 VPWR.t64 VGND 0.02189f
C10964 VPWR.n356 VGND 0.06768f
C10965 VPWR.t1457 VGND 0.10732f
C10966 VPWR.t1877 VGND 0.05805f
C10967 VPWR.t63 VGND 0.06817f
C10968 VPWR.t1548 VGND 0.08842f
C10969 VPWR.t986 VGND 0.02464f
C10970 VPWR.t1531 VGND 0.02189f
C10971 VPWR.n357 VGND 0.06768f
C10972 VPWR.n358 VGND 0.10289f
C10973 VPWR.n359 VGND 0.10289f
C10974 VPWR.t1549 VGND 0.02464f
C10975 VPWR.t1132 VGND 0.02189f
C10976 VPWR.n360 VGND 0.06768f
C10977 VPWR.t99 VGND 0.05805f
C10978 VPWR.t1131 VGND 0.06817f
C10979 VPWR.t1054 VGND 0.08842f
C10980 VPWR.t1156 VGND 0.02464f
C10981 VPWR.t1073 VGND 0.02189f
C10982 VPWR.n361 VGND 0.06768f
C10983 VPWR.n362 VGND 0.10289f
C10984 VPWR.n363 VGND 0.10289f
C10985 VPWR.t1055 VGND 0.02464f
C10986 VPWR.t1604 VGND 0.02189f
C10987 VPWR.n364 VGND 0.06768f
C10988 VPWR.t1876 VGND 0.05805f
C10989 VPWR.t1603 VGND 0.06817f
C10990 VPWR.t1261 VGND 0.08842f
C10991 VPWR.t116 VGND 0.02464f
C10992 VPWR.t1268 VGND 0.02189f
C10993 VPWR.n365 VGND 0.06768f
C10994 VPWR.n366 VGND 0.10289f
C10995 VPWR.n367 VGND 0.10289f
C10996 VPWR.t1262 VGND 0.02464f
C10997 VPWR.t1690 VGND 0.02189f
C10998 VPWR.n368 VGND 0.06768f
C10999 VPWR.t1878 VGND 0.05805f
C11000 VPWR.t1689 VGND 0.06817f
C11001 VPWR.t278 VGND 0.08842f
C11002 VPWR.t1872 VGND 0.02464f
C11003 VPWR.t955 VGND 0.02189f
C11004 VPWR.n369 VGND 0.06768f
C11005 VPWR.n370 VGND 0.10289f
C11006 VPWR.n371 VGND 0.10289f
C11007 VPWR.t279 VGND 0.02464f
C11008 VPWR.t1112 VGND 0.02189f
C11009 VPWR.n372 VGND 0.06768f
C11010 VPWR.t1874 VGND 0.05805f
C11011 VPWR.t1111 VGND 0.06817f
C11012 VPWR.t403 VGND 0.08842f
C11013 VPWR.t323 VGND 0.02464f
C11014 VPWR.t414 VGND 0.02189f
C11015 VPWR.n373 VGND 0.06768f
C11016 VPWR.n374 VGND 0.10289f
C11017 VPWR.n375 VGND 0.10289f
C11018 VPWR.t404 VGND 0.02464f
C11019 VPWR.t199 VGND 0.02189f
C11020 VPWR.n376 VGND 0.06768f
C11021 VPWR.t1720 VGND 0.05805f
C11022 VPWR.t198 VGND 0.06817f
C11023 VPWR.t964 VGND 0.08842f
C11024 VPWR.t1752 VGND 0.02464f
C11025 VPWR.t496 VGND 0.02189f
C11026 VPWR.n377 VGND 0.06768f
C11027 VPWR.n378 VGND 0.10289f
C11028 VPWR.n379 VGND 0.10289f
C11029 VPWR.t965 VGND 0.02464f
C11030 VPWR.t177 VGND 0.02189f
C11031 VPWR.n380 VGND 0.06768f
C11032 VPWR.t102 VGND 0.05805f
C11033 VPWR.t176 VGND 0.06817f
C11034 VPWR.t1422 VGND 0.08842f
C11035 VPWR.t293 VGND 0.02464f
C11036 VPWR.t1433 VGND 0.02189f
C11037 VPWR.n381 VGND 0.06768f
C11038 VPWR.n382 VGND 0.10289f
C11039 VPWR.n383 VGND 0.10289f
C11040 VPWR.t1423 VGND 0.02464f
C11041 VPWR.t1640 VGND 0.02189f
C11042 VPWR.n384 VGND 0.06768f
C11043 VPWR.t100 VGND 0.05805f
C11044 VPWR.t1639 VGND 0.06817f
C11045 VPWR.t394 VGND 0.02464f
C11046 VPWR.t881 VGND 0.02189f
C11047 VPWR.n385 VGND 0.06768f
C11048 VPWR.t187 VGND 0.02464f
C11049 VPWR.t602 VGND 0.02189f
C11050 VPWR.n386 VGND 0.06768f
C11051 VPWR.t1467 VGND 0.10732f
C11052 VPWR.t123 VGND 0.05805f
C11053 VPWR.t1617 VGND 0.06817f
C11054 VPWR.t1468 VGND 0.02464f
C11055 VPWR.t1618 VGND 0.02189f
C11056 VPWR.n387 VGND 0.06768f
C11057 VPWR.n388 VGND 0.01329f
C11058 VPWR.n390 VGND 0.08003f
C11059 VPWR.t312 VGND 0.08842f
C11060 VPWR.t980 VGND 0.05805f
C11061 VPWR.t1708 VGND 0.06817f
C11062 VPWR.t313 VGND 0.02464f
C11063 VPWR.t1709 VGND 0.02189f
C11064 VPWR.n391 VGND 0.06768f
C11065 VPWR.n392 VGND 0.01329f
C11066 VPWR.n394 VGND 0.08003f
C11067 VPWR.t1611 VGND 0.08842f
C11068 VPWR.t1323 VGND 0.05805f
C11069 VPWR.t1149 VGND 0.06817f
C11070 VPWR.t1612 VGND 0.02464f
C11071 VPWR.t1150 VGND 0.02189f
C11072 VPWR.n395 VGND 0.06768f
C11073 VPWR.n396 VGND 0.01329f
C11074 VPWR.n398 VGND 0.08003f
C11075 VPWR.t1173 VGND 0.08842f
C11076 VPWR.t1322 VGND 0.05805f
C11077 VPWR.t1058 VGND 0.06817f
C11078 VPWR.t1174 VGND 0.02464f
C11079 VPWR.t1059 VGND 0.02189f
C11080 VPWR.n399 VGND 0.06768f
C11081 VPWR.n400 VGND 0.01329f
C11082 VPWR.n402 VGND 0.08003f
C11083 VPWR.t1410 VGND 0.08842f
C11084 VPWR.t122 VGND 0.05805f
C11085 VPWR.t1318 VGND 0.06817f
C11086 VPWR.t1411 VGND 0.02464f
C11087 VPWR.t1319 VGND 0.02189f
C11088 VPWR.n403 VGND 0.06768f
C11089 VPWR.n404 VGND 0.01329f
C11090 VPWR.n406 VGND 0.08003f
C11091 VPWR.t1524 VGND 0.08842f
C11092 VPWR.t1704 VGND 0.05805f
C11093 VPWR.t1281 VGND 0.06817f
C11094 VPWR.t1525 VGND 0.02464f
C11095 VPWR.t1282 VGND 0.02189f
C11096 VPWR.n407 VGND 0.06768f
C11097 VPWR.n408 VGND 0.01329f
C11098 VPWR.n410 VGND 0.08003f
C11099 VPWR.t1275 VGND 0.08842f
C11100 VPWR.t1703 VGND 0.05805f
C11101 VPWR.t1857 VGND 0.06817f
C11102 VPWR.t1276 VGND 0.02464f
C11103 VPWR.t1858 VGND 0.02189f
C11104 VPWR.n411 VGND 0.06768f
C11105 VPWR.n412 VGND 0.01329f
C11106 VPWR.n414 VGND 0.08003f
C11107 VPWR.t234 VGND 0.08842f
C11108 VPWR.t121 VGND 0.05805f
C11109 VPWR.t535 VGND 0.06817f
C11110 VPWR.t235 VGND 0.02464f
C11111 VPWR.t536 VGND 0.02189f
C11112 VPWR.n415 VGND 0.06768f
C11113 VPWR.n416 VGND 0.01329f
C11114 VPWR.n418 VGND 0.08003f
C11115 VPWR.t242 VGND 0.08842f
C11116 VPWR.t120 VGND 0.05805f
C11117 VPWR.t981 VGND 0.06817f
C11118 VPWR.t243 VGND 0.02464f
C11119 VPWR.t982 VGND 0.02189f
C11120 VPWR.n419 VGND 0.06768f
C11121 VPWR.n420 VGND 0.01329f
C11122 VPWR.n422 VGND 0.08003f
C11123 VPWR.t134 VGND 0.08842f
C11124 VPWR.t1705 VGND 0.05805f
C11125 VPWR.t378 VGND 0.06817f
C11126 VPWR.t135 VGND 0.02464f
C11127 VPWR.t379 VGND 0.02189f
C11128 VPWR.n423 VGND 0.06768f
C11129 VPWR.n424 VGND 0.01329f
C11130 VPWR.n426 VGND 0.08003f
C11131 VPWR.t360 VGND 0.08842f
C11132 VPWR.t1321 VGND 0.05805f
C11133 VPWR.t1510 VGND 0.06817f
C11134 VPWR.t361 VGND 0.02464f
C11135 VPWR.t1511 VGND 0.02189f
C11136 VPWR.n427 VGND 0.06768f
C11137 VPWR.n428 VGND 0.01329f
C11138 VPWR.n430 VGND 0.08003f
C11139 VPWR.t1122 VGND 0.08842f
C11140 VPWR.t1320 VGND 0.05805f
C11141 VPWR.t1843 VGND 0.06817f
C11142 VPWR.t1123 VGND 0.02464f
C11143 VPWR.t1844 VGND 0.02189f
C11144 VPWR.n431 VGND 0.06768f
C11145 VPWR.n432 VGND 0.01329f
C11146 VPWR.n434 VGND 0.08003f
C11147 VPWR.t1540 VGND 0.08842f
C11148 VPWR.t1702 VGND 0.05805f
C11149 VPWR.t298 VGND 0.06817f
C11150 VPWR.t1541 VGND 0.02464f
C11151 VPWR.t299 VGND 0.02189f
C11152 VPWR.n435 VGND 0.06768f
C11153 VPWR.n436 VGND 0.01329f
C11154 VPWR.n438 VGND 0.08003f
C11155 VPWR.t53 VGND 0.08842f
C11156 VPWR.t1701 VGND 0.05805f
C11157 VPWR.t974 VGND 0.06817f
C11158 VPWR.t54 VGND 0.02464f
C11159 VPWR.t975 VGND 0.02189f
C11160 VPWR.n439 VGND 0.06768f
C11161 VPWR.n440 VGND 0.01329f
C11162 VPWR.n442 VGND 0.08003f
C11163 VPWR.t489 VGND 0.08842f
C11164 VPWR.t1324 VGND 0.05805f
C11165 VPWR.t397 VGND 0.06817f
C11166 VPWR.t490 VGND 0.02464f
C11167 VPWR.t398 VGND 0.02189f
C11168 VPWR.n443 VGND 0.06768f
C11169 VPWR.n444 VGND 0.01329f
C11170 VPWR.n446 VGND 0.08003f
C11171 VPWR.t186 VGND 0.08842f
C11172 VPWR.t119 VGND 0.05805f
C11173 VPWR.t601 VGND 0.0986f
C11174 VPWR.n447 VGND 0.05634f
C11175 VPWR.n448 VGND 0.01329f
C11176 VPWR.n449 VGND 0.10289f
C11177 VPWR.n450 VGND 0.75117f
C11178 VPWR.n451 VGND 0.10289f
C11179 VPWR.t5 VGND 0.02464f
C11180 VPWR.t714 VGND 0.02189f
C11181 VPWR.n452 VGND 0.06768f
C11182 VPWR.t188 VGND 0.06817f
C11183 VPWR.t1207 VGND 0.02464f
C11184 VPWR.t189 VGND 0.02189f
C11185 VPWR.n453 VGND 0.06768f
C11186 VPWR.n454 VGND 0.10289f
C11187 VPWR.n455 VGND 0.10289f
C11188 VPWR.t183 VGND 0.02464f
C11189 VPWR.t1083 VGND 0.02189f
C11190 VPWR.n456 VGND 0.06768f
C11191 VPWR.t280 VGND 0.06817f
C11192 VPWR.t1900 VGND 0.02464f
C11193 VPWR.t281 VGND 0.02189f
C11194 VPWR.n457 VGND 0.06768f
C11195 VPWR.n458 VGND 0.10289f
C11196 VPWR.n459 VGND 0.10289f
C11197 VPWR.t1736 VGND 0.02464f
C11198 VPWR.t1887 VGND 0.02189f
C11199 VPWR.n460 VGND 0.06768f
C11200 VPWR.t451 VGND 0.06817f
C11201 VPWR.t448 VGND 0.02464f
C11202 VPWR.t452 VGND 0.02189f
C11203 VPWR.n461 VGND 0.06768f
C11204 VPWR.n462 VGND 0.10289f
C11205 VPWR.n463 VGND 0.10289f
C11206 VPWR.t562 VGND 0.02464f
C11207 VPWR.t353 VGND 0.02189f
C11208 VPWR.n464 VGND 0.06768f
C11209 VPWR.t1219 VGND 0.06817f
C11210 VPWR.t1385 VGND 0.02464f
C11211 VPWR.t1220 VGND 0.02189f
C11212 VPWR.n465 VGND 0.06768f
C11213 VPWR.n466 VGND 0.10289f
C11214 VPWR.n467 VGND 0.10289f
C11215 VPWR.t221 VGND 0.02464f
C11216 VPWR.t169 VGND 0.02189f
C11217 VPWR.n468 VGND 0.06768f
C11218 VPWR.t224 VGND 0.06817f
C11219 VPWR.t1290 VGND 0.02464f
C11220 VPWR.t225 VGND 0.02189f
C11221 VPWR.n469 VGND 0.06768f
C11222 VPWR.n470 VGND 0.10289f
C11223 VPWR.n471 VGND 0.10289f
C11224 VPWR.t1580 VGND 0.02464f
C11225 VPWR.t1342 VGND 0.02189f
C11226 VPWR.n472 VGND 0.06768f
C11227 VPWR.t1304 VGND 0.06817f
C11228 VPWR.t147 VGND 0.02464f
C11229 VPWR.t1305 VGND 0.02189f
C11230 VPWR.n473 VGND 0.06768f
C11231 VPWR.n474 VGND 0.10289f
C11232 VPWR.n475 VGND 0.10289f
C11233 VPWR.t1190 VGND 0.02464f
C11234 VPWR.t1413 VGND 0.02189f
C11235 VPWR.n476 VGND 0.06768f
C11236 VPWR.t1167 VGND 0.06817f
C11237 VPWR.t129 VGND 0.02464f
C11238 VPWR.t1168 VGND 0.02189f
C11239 VPWR.n477 VGND 0.06768f
C11240 VPWR.n478 VGND 0.10289f
C11241 VPWR.n479 VGND 0.10289f
C11242 VPWR.t86 VGND 0.02464f
C11243 VPWR.t509 VGND 0.02189f
C11244 VPWR.n480 VGND 0.06768f
C11245 VPWR.t1476 VGND 0.10732f
C11246 VPWR.t1677 VGND 0.05805f
C11247 VPWR.t461 VGND 0.06817f
C11248 VPWR.t1477 VGND 0.02464f
C11249 VPWR.t462 VGND 0.02189f
C11250 VPWR.n481 VGND 0.06768f
C11251 VPWR.t1466 VGND 0.02464f
C11252 VPWR.t988 VGND 0.02189f
C11253 VPWR.n482 VGND 0.06768f
C11254 VPWR.t1465 VGND 0.10732f
C11255 VPWR.t1911 VGND 0.05805f
C11256 VPWR.t987 VGND 0.06817f
C11257 VPWR.t193 VGND 0.02464f
C11258 VPWR.t932 VGND 0.02189f
C11259 VPWR.n483 VGND 0.06768f
C11260 VPWR.n484 VGND 0.01329f
C11261 VPWR.n485 VGND 0.05634f
C11262 VPWR.t931 VGND 0.0986f
C11263 VPWR.t19 VGND 0.05805f
C11264 VPWR.t192 VGND 0.08842f
C11265 VPWR.t528 VGND 0.02464f
C11266 VPWR.t400 VGND 0.02189f
C11267 VPWR.n486 VGND 0.06768f
C11268 VPWR.n487 VGND 0.01329f
C11269 VPWR.n489 VGND 0.08003f
C11270 VPWR.t399 VGND 0.06817f
C11271 VPWR.t1847 VGND 0.05805f
C11272 VPWR.t527 VGND 0.08842f
C11273 VPWR.t283 VGND 0.02464f
C11274 VPWR.t1425 VGND 0.02189f
C11275 VPWR.n490 VGND 0.06768f
C11276 VPWR.n491 VGND 0.01329f
C11277 VPWR.n493 VGND 0.08003f
C11278 VPWR.t1424 VGND 0.06817f
C11279 VPWR.t30 VGND 0.05805f
C11280 VPWR.t282 VGND 0.08842f
C11281 VPWR.t36 VGND 0.02464f
C11282 VPWR.t161 VGND 0.02189f
C11283 VPWR.n494 VGND 0.06768f
C11284 VPWR.n495 VGND 0.01329f
C11285 VPWR.n497 VGND 0.08003f
C11286 VPWR.t160 VGND 0.06817f
C11287 VPWR.t31 VGND 0.05805f
C11288 VPWR.t35 VGND 0.08842f
C11289 VPWR.t1513 VGND 0.02464f
C11290 VPWR.t967 VGND 0.02189f
C11291 VPWR.n498 VGND 0.06768f
C11292 VPWR.n499 VGND 0.01329f
C11293 VPWR.n501 VGND 0.08003f
C11294 VPWR.t966 VGND 0.06817f
C11295 VPWR.t1912 VGND 0.05805f
C11296 VPWR.t1512 VGND 0.08842f
C11297 VPWR.t381 VGND 0.02464f
C11298 VPWR.t1744 VGND 0.02189f
C11299 VPWR.n502 VGND 0.06768f
C11300 VPWR.n503 VGND 0.01329f
C11301 VPWR.n505 VGND 0.08003f
C11302 VPWR.t1743 VGND 0.06817f
C11303 VPWR.t1913 VGND 0.05805f
C11304 VPWR.t380 VGND 0.08842f
C11305 VPWR.t1039 VGND 0.02464f
C11306 VPWR.t406 VGND 0.02189f
C11307 VPWR.n506 VGND 0.06768f
C11308 VPWR.n507 VGND 0.01329f
C11309 VPWR.n509 VGND 0.08003f
C11310 VPWR.t405 VGND 0.06817f
C11311 VPWR.t34 VGND 0.05805f
C11312 VPWR.t1038 VGND 0.08842f
C11313 VPWR.t500 VGND 0.02464f
C11314 VPWR.t1043 VGND 0.02189f
C11315 VPWR.n510 VGND 0.06768f
C11316 VPWR.n511 VGND 0.01329f
C11317 VPWR.n513 VGND 0.08003f
C11318 VPWR.t1042 VGND 0.06817f
C11319 VPWR.t20 VGND 0.05805f
C11320 VPWR.t499 VGND 0.08842f
C11321 VPWR.t1860 VGND 0.02464f
C11322 VPWR.t271 VGND 0.02189f
C11323 VPWR.n514 VGND 0.06768f
C11324 VPWR.n515 VGND 0.01329f
C11325 VPWR.n517 VGND 0.08003f
C11326 VPWR.t270 VGND 0.06817f
C11327 VPWR.t1909 VGND 0.05805f
C11328 VPWR.t1859 VGND 0.08842f
C11329 VPWR.t1481 VGND 0.02464f
C11330 VPWR.t1864 VGND 0.02189f
C11331 VPWR.n518 VGND 0.06768f
C11332 VPWR.n519 VGND 0.01329f
C11333 VPWR.n521 VGND 0.08003f
C11334 VPWR.t1863 VGND 0.06817f
C11335 VPWR.t32 VGND 0.05805f
C11336 VPWR.t1480 VGND 0.08842f
C11337 VPWR.t1527 VGND 0.02464f
C11338 VPWR.t1485 VGND 0.02189f
C11339 VPWR.n522 VGND 0.06768f
C11340 VPWR.n523 VGND 0.01329f
C11341 VPWR.n525 VGND 0.08003f
C11342 VPWR.t1484 VGND 0.06817f
C11343 VPWR.t33 VGND 0.05805f
C11344 VPWR.t1526 VGND 0.08842f
C11345 VPWR.t1045 VGND 0.02464f
C11346 VPWR.t108 VGND 0.02189f
C11347 VPWR.n526 VGND 0.06768f
C11348 VPWR.n527 VGND 0.01329f
C11349 VPWR.n529 VGND 0.08003f
C11350 VPWR.t107 VGND 0.06817f
C11351 VPWR.t1910 VGND 0.05805f
C11352 VPWR.t1044 VGND 0.08842f
C11353 VPWR.t1166 VGND 0.02464f
C11354 VPWR.t1079 VGND 0.02189f
C11355 VPWR.n530 VGND 0.06768f
C11356 VPWR.n531 VGND 0.01329f
C11357 VPWR.n533 VGND 0.08003f
C11358 VPWR.t1078 VGND 0.06817f
C11359 VPWR.t1845 VGND 0.05805f
C11360 VPWR.t1165 VGND 0.08842f
C11361 VPWR.t1713 VGND 0.02464f
C11362 VPWR.t1142 VGND 0.02189f
C11363 VPWR.n534 VGND 0.06768f
C11364 VPWR.n535 VGND 0.01329f
C11365 VPWR.n537 VGND 0.08003f
C11366 VPWR.t1141 VGND 0.06817f
C11367 VPWR.t1846 VGND 0.05805f
C11368 VPWR.t1712 VGND 0.08842f
C11369 VPWR.t1620 VGND 0.02464f
C11370 VPWR.t1717 VGND 0.02189f
C11371 VPWR.n538 VGND 0.06768f
C11372 VPWR.n539 VGND 0.01329f
C11373 VPWR.n541 VGND 0.08003f
C11374 VPWR.t1716 VGND 0.06817f
C11375 VPWR.t18 VGND 0.05805f
C11376 VPWR.t1619 VGND 0.08842f
C11377 VPWR.n542 VGND 0.08003f
C11378 VPWR.n544 VGND 0.01329f
C11379 VPWR.n545 VGND 0.10289f
C11380 VPWR.n546 VGND 0.74646f
C11381 VPWR.n547 VGND 0.10289f
C11382 VPWR.t1452 VGND 0.02464f
C11383 VPWR.t1108 VGND 0.02189f
C11384 VPWR.n548 VGND 0.06768f
C11385 VPWR.t1451 VGND 0.10732f
C11386 VPWR.t347 VGND 0.05805f
C11387 VPWR.t1107 VGND 0.06817f
C11388 VPWR.t1647 VGND 0.08842f
C11389 VPWR.t558 VGND 0.02464f
C11390 VPWR.t1656 VGND 0.02189f
C11391 VPWR.n549 VGND 0.06768f
C11392 VPWR.n550 VGND 0.10289f
C11393 VPWR.n551 VGND 0.10289f
C11394 VPWR.t1648 VGND 0.02464f
C11395 VPWR.t1182 VGND 0.02189f
C11396 VPWR.n552 VGND 0.06768f
C11397 VPWR.t1439 VGND 0.05805f
C11398 VPWR.t1181 VGND 0.06817f
C11399 VPWR.t1068 VGND 0.08842f
C11400 VPWR.t1144 VGND 0.02464f
C11401 VPWR.t1024 VGND 0.02189f
C11402 VPWR.n553 VGND 0.06768f
C11403 VPWR.n554 VGND 0.10289f
C11404 VPWR.n555 VGND 0.10289f
C11405 VPWR.t1069 VGND 0.02464f
C11406 VPWR.t1563 VGND 0.02189f
C11407 VPWR.n556 VGND 0.06768f
C11408 VPWR.t346 VGND 0.05805f
C11409 VPWR.t1562 VGND 0.06817f
C11410 VPWR.t1496 VGND 0.08842f
C11411 VPWR.t1555 VGND 0.02464f
C11412 VPWR.t1505 VGND 0.02189f
C11413 VPWR.n557 VGND 0.06768f
C11414 VPWR.n558 VGND 0.10289f
C11415 VPWR.n559 VGND 0.10289f
C11416 VPWR.t1497 VGND 0.02464f
C11417 VPWR.t217 VGND 0.02189f
C11418 VPWR.n560 VGND 0.06768f
C11419 VPWR.t1680 VGND 0.05805f
C11420 VPWR.t216 VGND 0.06817f
C11421 VPWR.t250 VGND 0.08842f
C11422 VPWR.t1698 VGND 0.02464f
C11423 VPWR.t1402 VGND 0.02189f
C11424 VPWR.n561 VGND 0.06768f
C11425 VPWR.n562 VGND 0.10289f
C11426 VPWR.n563 VGND 0.10289f
C11427 VPWR.t251 VGND 0.02464f
C11428 VPWR.t74 VGND 0.02189f
C11429 VPWR.n564 VGND 0.06768f
C11430 VPWR.t344 VGND 0.05805f
C11431 VPWR.t73 VGND 0.06817f
C11432 VPWR.t435 VGND 0.08842f
C11433 VPWR.t523 VGND 0.02464f
C11434 VPWR.t444 VGND 0.02189f
C11435 VPWR.n565 VGND 0.06768f
C11436 VPWR.n566 VGND 0.10289f
C11437 VPWR.n567 VGND 0.10289f
C11438 VPWR.t436 VGND 0.02464f
C11439 VPWR.t484 VGND 0.02189f
C11440 VPWR.n568 VGND 0.06768f
C11441 VPWR.t1437 VGND 0.05805f
C11442 VPWR.t483 VGND 0.06817f
C11443 VPWR.t1441 VGND 0.08842f
C11444 VPWR.t476 VGND 0.02464f
C11445 VPWR.t1896 VGND 0.02189f
C11446 VPWR.n569 VGND 0.06768f
C11447 VPWR.n570 VGND 0.10289f
C11448 VPWR.n571 VGND 0.10289f
C11449 VPWR.t1442 VGND 0.02464f
C11450 VPWR.t46 VGND 0.02189f
C11451 VPWR.n572 VGND 0.06768f
C11452 VPWR.t1679 VGND 0.05805f
C11453 VPWR.t45 VGND 0.06817f
C11454 VPWR.t1568 VGND 0.08842f
C11455 VPWR.t167 VGND 0.02464f
C11456 VPWR.t1203 VGND 0.02189f
C11457 VPWR.n573 VGND 0.06768f
C11458 VPWR.n574 VGND 0.10289f
C11459 VPWR.n575 VGND 0.10289f
C11460 VPWR.t1569 VGND 0.02464f
C11461 VPWR.t203 VGND 0.02189f
C11462 VPWR.n576 VGND 0.06768f
C11463 VPWR.t1440 VGND 0.05805f
C11464 VPWR.t202 VGND 0.06817f
C11465 VPWR.t1636 VGND 0.02464f
C11466 VPWR.t781 VGND 0.02189f
C11467 VPWR.n577 VGND 0.06768f
C11468 VPWR.t390 VGND 0.02464f
C11469 VPWR.t889 VGND 0.02189f
C11470 VPWR.n578 VGND 0.06768f
C11471 VPWR.t1459 VGND 0.10732f
C11472 VPWR.t433 VGND 0.05805f
C11473 VPWR.t993 VGND 0.06817f
C11474 VPWR.t1460 VGND 0.02464f
C11475 VPWR.t994 VGND 0.02189f
C11476 VPWR.n579 VGND 0.06768f
C11477 VPWR.n580 VGND 0.01329f
C11478 VPWR.n582 VGND 0.08003f
C11479 VPWR.t983 VGND 0.08842f
C11480 VPWR.t428 VGND 0.05805f
C11481 VPWR.t314 VGND 0.06817f
C11482 VPWR.t984 VGND 0.02464f
C11483 VPWR.t315 VGND 0.02189f
C11484 VPWR.n583 VGND 0.06768f
C11485 VPWR.n584 VGND 0.01329f
C11486 VPWR.n586 VGND 0.08003f
C11487 VPWR.t1546 VGND 0.08842f
C11488 VPWR.t470 VGND 0.05805f
C11489 VPWR.t1133 VGND 0.06817f
C11490 VPWR.t1547 VGND 0.02464f
C11491 VPWR.t1134 VGND 0.02189f
C11492 VPWR.n587 VGND 0.06768f
C11493 VPWR.n588 VGND 0.01329f
C11494 VPWR.n590 VGND 0.08003f
C11495 VPWR.t1157 VGND 0.08842f
C11496 VPWR.t469 VGND 0.05805f
C11497 VPWR.t1070 VGND 0.06817f
C11498 VPWR.t1158 VGND 0.02464f
C11499 VPWR.t1071 VGND 0.02189f
C11500 VPWR.n591 VGND 0.06768f
C11501 VPWR.n592 VGND 0.01329f
C11502 VPWR.n594 VGND 0.08003f
C11503 VPWR.t1050 VGND 0.08842f
C11504 VPWR.t432 VGND 0.05805f
C11505 VPWR.t1601 VGND 0.06817f
C11506 VPWR.t1051 VGND 0.02464f
C11507 VPWR.t1602 VGND 0.02189f
C11508 VPWR.n595 VGND 0.06768f
C11509 VPWR.n596 VGND 0.01329f
C11510 VPWR.n598 VGND 0.08003f
C11511 VPWR.t113 VGND 0.08842f
C11512 VPWR.t426 VGND 0.05805f
C11513 VPWR.t1265 VGND 0.06817f
C11514 VPWR.t114 VGND 0.02464f
C11515 VPWR.t1266 VGND 0.02189f
C11516 VPWR.n599 VGND 0.06768f
C11517 VPWR.n600 VGND 0.01329f
C11518 VPWR.n602 VGND 0.08003f
C11519 VPWR.t1259 VGND 0.08842f
C11520 VPWR.t425 VGND 0.05805f
C11521 VPWR.t1687 VGND 0.06817f
C11522 VPWR.t1260 VGND 0.02464f
C11523 VPWR.t1688 VGND 0.02189f
C11524 VPWR.n603 VGND 0.06768f
C11525 VPWR.n604 VGND 0.01329f
C11526 VPWR.n606 VGND 0.08003f
C11527 VPWR.t1869 VGND 0.08842f
C11528 VPWR.t431 VGND 0.05805f
C11529 VPWR.t256 VGND 0.06817f
C11530 VPWR.t1870 VGND 0.02464f
C11531 VPWR.t257 VGND 0.02189f
C11532 VPWR.n607 VGND 0.06768f
C11533 VPWR.n608 VGND 0.01329f
C11534 VPWR.n610 VGND 0.08003f
C11535 VPWR.t276 VGND 0.08842f
C11536 VPWR.t430 VGND 0.05805f
C11537 VPWR.t326 VGND 0.06817f
C11538 VPWR.t277 VGND 0.02464f
C11539 VPWR.t327 VGND 0.02189f
C11540 VPWR.n611 VGND 0.06768f
C11541 VPWR.n612 VGND 0.01329f
C11542 VPWR.n614 VGND 0.08003f
C11543 VPWR.t320 VGND 0.08842f
C11544 VPWR.t427 VGND 0.05805f
C11545 VPWR.t411 VGND 0.06817f
C11546 VPWR.t321 VGND 0.02464f
C11547 VPWR.t412 VGND 0.02189f
C11548 VPWR.n615 VGND 0.06768f
C11549 VPWR.n616 VGND 0.01329f
C11550 VPWR.n618 VGND 0.08003f
C11551 VPWR.t401 VGND 0.08842f
C11552 VPWR.t468 VGND 0.05805f
C11553 VPWR.t1755 VGND 0.06817f
C11554 VPWR.t402 VGND 0.02464f
C11555 VPWR.t1756 VGND 0.02189f
C11556 VPWR.n619 VGND 0.06768f
C11557 VPWR.n620 VGND 0.01329f
C11558 VPWR.n622 VGND 0.08003f
C11559 VPWR.t1749 VGND 0.08842f
C11560 VPWR.t434 VGND 0.05805f
C11561 VPWR.t493 VGND 0.06817f
C11562 VPWR.t1750 VGND 0.02464f
C11563 VPWR.t494 VGND 0.02189f
C11564 VPWR.n623 VGND 0.06768f
C11565 VPWR.n624 VGND 0.01329f
C11566 VPWR.n626 VGND 0.08003f
C11567 VPWR.t962 VGND 0.08842f
C11568 VPWR.t424 VGND 0.05805f
C11569 VPWR.t174 VGND 0.06817f
C11570 VPWR.t963 VGND 0.02464f
C11571 VPWR.t175 VGND 0.02189f
C11572 VPWR.n627 VGND 0.06768f
C11573 VPWR.n628 VGND 0.01329f
C11574 VPWR.n630 VGND 0.08003f
C11575 VPWR.t290 VGND 0.08842f
C11576 VPWR.t423 VGND 0.05805f
C11577 VPWR.t1430 VGND 0.06817f
C11578 VPWR.t291 VGND 0.02464f
C11579 VPWR.t1431 VGND 0.02189f
C11580 VPWR.n631 VGND 0.06768f
C11581 VPWR.n632 VGND 0.01329f
C11582 VPWR.n634 VGND 0.08003f
C11583 VPWR.t1420 VGND 0.08842f
C11584 VPWR.t422 VGND 0.05805f
C11585 VPWR.t1637 VGND 0.06817f
C11586 VPWR.t1421 VGND 0.02464f
C11587 VPWR.t1638 VGND 0.02189f
C11588 VPWR.n635 VGND 0.06768f
C11589 VPWR.n636 VGND 0.01329f
C11590 VPWR.n638 VGND 0.08003f
C11591 VPWR.t389 VGND 0.08842f
C11592 VPWR.t429 VGND 0.05805f
C11593 VPWR.t888 VGND 0.0986f
C11594 VPWR.n639 VGND 0.05634f
C11595 VPWR.n640 VGND 0.01329f
C11596 VPWR.n641 VGND 0.10289f
C11597 VPWR.n642 VGND 0.75117f
C11598 VPWR.n643 VGND 0.10289f
C11599 VPWR.t207 VGND 0.02464f
C11600 VPWR.t615 VGND 0.02189f
C11601 VPWR.n644 VGND 0.06768f
C11602 VPWR.t391 VGND 0.06817f
C11603 VPWR.t486 VGND 0.02464f
C11604 VPWR.t392 VGND 0.02189f
C11605 VPWR.n645 VGND 0.06768f
C11606 VPWR.n646 VGND 0.10289f
C11607 VPWR.n647 VGND 0.10289f
C11608 VPWR.t50 VGND 0.02464f
C11609 VPWR.t492 VGND 0.02189f
C11610 VPWR.n648 VGND 0.06768f
C11611 VPWR.t294 VGND 0.06817f
C11612 VPWR.t1537 VGND 0.02464f
C11613 VPWR.t295 VGND 0.02189f
C11614 VPWR.n649 VGND 0.06768f
C11615 VPWR.n650 VGND 0.10289f
C11616 VPWR.n651 VGND 0.10289f
C11617 VPWR.t1119 VGND 0.02464f
C11618 VPWR.t1840 VGND 0.02189f
C11619 VPWR.n652 VGND 0.06768f
C11620 VPWR.t1124 VGND 0.06817f
C11621 VPWR.t357 VGND 0.02464f
C11622 VPWR.t1125 VGND 0.02189f
C11623 VPWR.n653 VGND 0.06768f
C11624 VPWR.n654 VGND 0.10289f
C11625 VPWR.n655 VGND 0.10289f
C11626 VPWR.t131 VGND 0.02464f
C11627 VPWR.t363 VGND 0.02189f
C11628 VPWR.n656 VGND 0.06768f
C11629 VPWR.t136 VGND 0.06817f
C11630 VPWR.t1406 VGND 0.02464f
C11631 VPWR.t137 VGND 0.02189f
C11632 VPWR.n657 VGND 0.06768f
C11633 VPWR.n658 VGND 0.10289f
C11634 VPWR.n659 VGND 0.10289f
C11635 VPWR.t231 VGND 0.02464f
C11636 VPWR.t532 VGND 0.02189f
C11637 VPWR.n660 VGND 0.06768f
C11638 VPWR.t236 VGND 0.06817f
C11639 VPWR.t1272 VGND 0.02464f
C11640 VPWR.t237 VGND 0.02189f
C11641 VPWR.n661 VGND 0.06768f
C11642 VPWR.n662 VGND 0.10289f
C11643 VPWR.n663 VGND 0.10289f
C11644 VPWR.t1521 VGND 0.02464f
C11645 VPWR.t1278 VGND 0.02189f
C11646 VPWR.n664 VGND 0.06768f
C11647 VPWR.t1314 VGND 0.06817f
C11648 VPWR.t1028 VGND 0.02464f
C11649 VPWR.t1315 VGND 0.02189f
C11650 VPWR.n665 VGND 0.06768f
C11651 VPWR.n666 VGND 0.10289f
C11652 VPWR.n667 VGND 0.10289f
C11653 VPWR.t1180 VGND 0.02464f
C11654 VPWR.t1053 VGND 0.02189f
C11655 VPWR.n668 VGND 0.06768f
C11656 VPWR.t1153 VGND 0.06817f
C11657 VPWR.t1608 VGND 0.02464f
C11658 VPWR.t1154 VGND 0.02189f
C11659 VPWR.n669 VGND 0.06768f
C11660 VPWR.n670 VGND 0.10289f
C11661 VPWR.n671 VGND 0.10289f
C11662 VPWR.t309 VGND 0.02464f
C11663 VPWR.t1614 VGND 0.02189f
C11664 VPWR.n672 VGND 0.06768f
C11665 VPWR.t1471 VGND 0.10732f
C11666 VPWR.t1089 VGND 0.05805f
C11667 VPWR.t995 VGND 0.06817f
C11668 VPWR.t1472 VGND 0.02464f
C11669 VPWR.t996 VGND 0.02189f
C11670 VPWR.n673 VGND 0.06768f
C11671 VPWR.t1479 VGND 0.02464f
C11672 VPWR.t90 VGND 0.02189f
C11673 VPWR.n674 VGND 0.06768f
C11674 VPWR.t1478 VGND 0.10732f
C11675 VPWR.t467 VGND 0.05805f
C11676 VPWR.t89 VGND 0.06817f
C11677 VPWR.t1646 VGND 0.02464f
C11678 VPWR.t722 VGND 0.02189f
C11679 VPWR.n675 VGND 0.06768f
C11680 VPWR.n676 VGND 0.01329f
C11681 VPWR.n677 VGND 0.05634f
C11682 VPWR.t721 VGND 0.0986f
C11683 VPWR.t1096 VGND 0.05805f
C11684 VPWR.t1645 VGND 0.08842f
C11685 VPWR.t1205 VGND 0.02464f
C11686 VPWR.t185 VGND 0.02189f
C11687 VPWR.n678 VGND 0.06768f
C11688 VPWR.n679 VGND 0.01329f
C11689 VPWR.n681 VGND 0.08003f
C11690 VPWR.t184 VGND 0.06817f
C11691 VPWR.t1197 VGND 0.05805f
C11692 VPWR.t1204 VGND 0.08842f
C11693 VPWR.t181 VGND 0.02464f
C11694 VPWR.t1584 VGND 0.02189f
C11695 VPWR.n682 VGND 0.06768f
C11696 VPWR.n683 VGND 0.01329f
C11697 VPWR.n685 VGND 0.08003f
C11698 VPWR.t1583 VGND 0.06817f
C11699 VPWR.t1198 VGND 0.05805f
C11700 VPWR.t180 VGND 0.08842f
C11701 VPWR.t1898 VGND 0.02464f
C11702 VPWR.t56 VGND 0.02189f
C11703 VPWR.n686 VGND 0.06768f
C11704 VPWR.n687 VGND 0.01329f
C11705 VPWR.n689 VGND 0.08003f
C11706 VPWR.t55 VGND 0.06817f
C11707 VPWR.t1199 VGND 0.05805f
C11708 VPWR.t1897 VGND 0.08842f
C11709 VPWR.t1734 VGND 0.02464f
C11710 VPWR.t1883 VGND 0.02189f
C11711 VPWR.n690 VGND 0.06768f
C11712 VPWR.n691 VGND 0.01329f
C11713 VPWR.n693 VGND 0.08003f
C11714 VPWR.t1882 VGND 0.06817f
C11715 VPWR.t1098 VGND 0.05805f
C11716 VPWR.t1733 VGND 0.08842f
C11717 VPWR.t446 VGND 0.02464f
C11718 VPWR.t1738 VGND 0.02189f
C11719 VPWR.n694 VGND 0.06768f
C11720 VPWR.n695 VGND 0.01329f
C11721 VPWR.n697 VGND 0.08003f
C11722 VPWR.t1737 VGND 0.06817f
C11723 VPWR.t1099 VGND 0.05805f
C11724 VPWR.t445 VGND 0.08842f
C11725 VPWR.t560 VGND 0.02464f
C11726 VPWR.t349 VGND 0.02189f
C11727 VPWR.n698 VGND 0.06768f
C11728 VPWR.n699 VGND 0.01329f
C11729 VPWR.n701 VGND 0.08003f
C11730 VPWR.t348 VGND 0.06817f
C11731 VPWR.t1673 VGND 0.05805f
C11732 VPWR.t559 VGND 0.08842f
C11733 VPWR.t959 VGND 0.02464f
C11734 VPWR.t564 VGND 0.02189f
C11735 VPWR.n702 VGND 0.06768f
C11736 VPWR.n703 VGND 0.01329f
C11737 VPWR.n705 VGND 0.08003f
C11738 VPWR.t563 VGND 0.06817f
C11739 VPWR.t1097 VGND 0.05805f
C11740 VPWR.t958 VGND 0.08842f
C11741 VPWR.t953 VGND 0.02464f
C11742 VPWR.t245 VGND 0.02189f
C11743 VPWR.n706 VGND 0.06768f
C11744 VPWR.n707 VGND 0.01329f
C11745 VPWR.n709 VGND 0.08003f
C11746 VPWR.t244 VGND 0.06817f
C11747 VPWR.t465 VGND 0.05805f
C11748 VPWR.t952 VGND 0.08842f
C11749 VPWR.t1288 VGND 0.02464f
C11750 VPWR.t223 VGND 0.02189f
C11751 VPWR.n710 VGND 0.06768f
C11752 VPWR.n711 VGND 0.01329f
C11753 VPWR.n713 VGND 0.08003f
C11754 VPWR.t222 VGND 0.06817f
C11755 VPWR.t1671 VGND 0.05805f
C11756 VPWR.t1287 VGND 0.08842f
C11757 VPWR.t1578 VGND 0.02464f
C11758 VPWR.t1292 VGND 0.02189f
C11759 VPWR.n714 VGND 0.06768f
C11760 VPWR.n715 VGND 0.01329f
C11761 VPWR.n717 VGND 0.08003f
C11762 VPWR.t1291 VGND 0.06817f
C11763 VPWR.t1672 VGND 0.05805f
C11764 VPWR.t1577 VGND 0.08842f
C11765 VPWR.t145 VGND 0.02464f
C11766 VPWR.t1303 VGND 0.02189f
C11767 VPWR.n718 VGND 0.06768f
C11768 VPWR.n719 VGND 0.01329f
C11769 VPWR.n721 VGND 0.08003f
C11770 VPWR.t1302 VGND 0.06817f
C11771 VPWR.t466 VGND 0.05805f
C11772 VPWR.t144 VGND 0.08842f
C11773 VPWR.t1192 VGND 0.02464f
C11774 VPWR.t1409 VGND 0.02189f
C11775 VPWR.n722 VGND 0.06768f
C11776 VPWR.n723 VGND 0.01329f
C11777 VPWR.n725 VGND 0.08003f
C11778 VPWR.t1408 VGND 0.06817f
C11779 VPWR.t1100 VGND 0.05805f
C11780 VPWR.t1191 VGND 0.08842f
C11781 VPWR.t127 VGND 0.02464f
C11782 VPWR.t1170 VGND 0.02189f
C11783 VPWR.n726 VGND 0.06768f
C11784 VPWR.n727 VGND 0.01329f
C11785 VPWR.n729 VGND 0.08003f
C11786 VPWR.t1169 VGND 0.06817f
C11787 VPWR.t1196 VGND 0.05805f
C11788 VPWR.t126 VGND 0.08842f
C11789 VPWR.t1110 VGND 0.02464f
C11790 VPWR.t507 VGND 0.02189f
C11791 VPWR.n730 VGND 0.06768f
C11792 VPWR.n731 VGND 0.01329f
C11793 VPWR.n733 VGND 0.08003f
C11794 VPWR.t506 VGND 0.06817f
C11795 VPWR.t1674 VGND 0.05805f
C11796 VPWR.t1109 VGND 0.08842f
C11797 VPWR.n734 VGND 0.08003f
C11798 VPWR.n736 VGND 0.01329f
C11799 VPWR.n737 VGND 0.10289f
C11800 VPWR.n738 VGND 0.74646f
C11801 VPWR.n739 VGND 0.10289f
C11802 VPWR.t1475 VGND 0.02464f
C11803 VPWR.t464 VGND 0.02189f
C11804 VPWR.n740 VGND 0.06768f
C11805 VPWR.t1474 VGND 0.10732f
C11806 VPWR.t1250 VGND 0.05805f
C11807 VPWR.t463 VGND 0.06817f
C11808 VPWR.t510 VGND 0.08842f
C11809 VPWR.t460 VGND 0.02464f
C11810 VPWR.t513 VGND 0.02189f
C11811 VPWR.n741 VGND 0.06768f
C11812 VPWR.n742 VGND 0.10289f
C11813 VPWR.n743 VGND 0.10289f
C11814 VPWR.t511 VGND 0.02464f
C11815 VPWR.t1162 VGND 0.02189f
C11816 VPWR.n744 VGND 0.06768f
C11817 VPWR.t1006 VGND 0.05805f
C11818 VPWR.t1161 VGND 0.06817f
C11819 VPWR.t148 VGND 0.08842f
C11820 VPWR.t1186 VGND 0.02464f
C11821 VPWR.t1415 VGND 0.02189f
C11822 VPWR.n745 VGND 0.06768f
C11823 VPWR.n746 VGND 0.10289f
C11824 VPWR.n747 VGND 0.10289f
C11825 VPWR.t149 VGND 0.02464f
C11826 VPWR.t1309 VGND 0.02189f
C11827 VPWR.n748 VGND 0.06768f
C11828 VPWR.t1249 VGND 0.05805f
C11829 VPWR.t1308 VGND 0.06817f
C11830 VPWR.t1343 VGND 0.08842f
C11831 VPWR.t1307 VGND 0.02464f
C11832 VPWR.t1346 VGND 0.02189f
C11833 VPWR.n749 VGND 0.06768f
C11834 VPWR.n750 VGND 0.10289f
C11835 VPWR.n751 VGND 0.10289f
C11836 VPWR.t1344 VGND 0.02464f
C11837 VPWR.t229 VGND 0.02189f
C11838 VPWR.n752 VGND 0.06768f
C11839 VPWR.t1010 VGND 0.05805f
C11840 VPWR.t228 VGND 0.06817f
C11841 VPWR.t1386 VGND 0.08842f
C11842 VPWR.t227 VGND 0.02464f
C11843 VPWR.t502 VGND 0.02189f
C11844 VPWR.n753 VGND 0.06768f
C11845 VPWR.n754 VGND 0.10289f
C11846 VPWR.n755 VGND 0.10289f
C11847 VPWR.t1387 VGND 0.02464f
C11848 VPWR.t1224 VGND 0.02189f
C11849 VPWR.n756 VGND 0.06768f
C11850 VPWR.t1247 VGND 0.05805f
C11851 VPWR.t1223 VGND 0.06817f
C11852 VPWR.t350 VGND 0.08842f
C11853 VPWR.t1222 VGND 0.02464f
C11854 VPWR.t355 VGND 0.02189f
C11855 VPWR.n757 VGND 0.06768f
C11856 VPWR.n758 VGND 0.10289f
C11857 VPWR.n759 VGND 0.10289f
C11858 VPWR.t351 VGND 0.02464f
C11859 VPWR.t1851 VGND 0.02189f
C11860 VPWR.n760 VGND 0.06768f
C11861 VPWR.t1004 VGND 0.05805f
C11862 VPWR.t1850 VGND 0.06817f
C11863 VPWR.t1884 VGND 0.08842f
C11864 VPWR.t1849 VGND 0.02464f
C11865 VPWR.t1535 VGND 0.02189f
C11866 VPWR.n761 VGND 0.06768f
C11867 VPWR.n762 VGND 0.10289f
C11868 VPWR.n763 VGND 0.10289f
C11869 VPWR.t1885 VGND 0.02464f
C11870 VPWR.t285 VGND 0.02189f
C11871 VPWR.n764 VGND 0.06768f
C11872 VPWR.t1009 VGND 0.05805f
C11873 VPWR.t284 VGND 0.06817f
C11874 VPWR.t1585 VGND 0.08842f
C11875 VPWR.t40 VGND 0.02464f
C11876 VPWR.t1085 VGND 0.02189f
C11877 VPWR.n765 VGND 0.06768f
C11878 VPWR.n766 VGND 0.10289f
C11879 VPWR.n767 VGND 0.10289f
C11880 VPWR.t1586 VGND 0.02464f
C11881 VPWR.t191 VGND 0.02189f
C11882 VPWR.n768 VGND 0.06768f
C11883 VPWR.t1007 VGND 0.05805f
C11884 VPWR.t190 VGND 0.06817f
C11885 VPWR.t7 VGND 0.02464f
C11886 VPWR.t682 VGND 0.02189f
C11887 VPWR.n769 VGND 0.06768f
C11888 VPWR.t1632 VGND 0.02464f
C11889 VPWR.t787 VGND 0.02189f
C11890 VPWR.n770 VGND 0.06768f
C11891 VPWR.t1453 VGND 0.10732f
C11892 VPWR.t1340 VGND 0.05805f
C11893 VPWR.t1105 VGND 0.06817f
C11894 VPWR.t1454 VGND 0.02464f
C11895 VPWR.t1106 VGND 0.02189f
C11896 VPWR.n771 VGND 0.06768f
C11897 VPWR.n772 VGND 0.01329f
C11898 VPWR.n774 VGND 0.08003f
C11899 VPWR.t555 VGND 0.08842f
C11900 VPWR.t1335 VGND 0.05805f
C11901 VPWR.t1651 VGND 0.06817f
C11902 VPWR.t556 VGND 0.02464f
C11903 VPWR.t1652 VGND 0.02189f
C11904 VPWR.n775 VGND 0.06768f
C11905 VPWR.n776 VGND 0.01329f
C11906 VPWR.n778 VGND 0.08003f
C11907 VPWR.t516 VGND 0.08842f
C11908 VPWR.t1380 VGND 0.05805f
C11909 VPWR.t1175 VGND 0.06817f
C11910 VPWR.t517 VGND 0.02464f
C11911 VPWR.t1176 VGND 0.02189f
C11912 VPWR.n779 VGND 0.06768f
C11913 VPWR.n780 VGND 0.01329f
C11914 VPWR.n782 VGND 0.08003f
C11915 VPWR.t1145 VGND 0.08842f
C11916 VPWR.t1379 VGND 0.05805f
C11917 VPWR.t152 VGND 0.06817f
C11918 VPWR.t1146 VGND 0.02464f
C11919 VPWR.t153 VGND 0.02189f
C11920 VPWR.n783 VGND 0.06768f
C11921 VPWR.n784 VGND 0.01329f
C11922 VPWR.n786 VGND 0.08003f
C11923 VPWR.t1064 VGND 0.08842f
C11924 VPWR.t1339 VGND 0.05805f
C11925 VPWR.t1558 VGND 0.06817f
C11926 VPWR.t1065 VGND 0.02464f
C11927 VPWR.t1559 VGND 0.02189f
C11928 VPWR.n787 VGND 0.06768f
C11929 VPWR.n788 VGND 0.01329f
C11930 VPWR.n790 VGND 0.08003f
C11931 VPWR.t1552 VGND 0.08842f
C11932 VPWR.t1333 VGND 0.05805f
C11933 VPWR.t1500 VGND 0.06817f
C11934 VPWR.t1553 VGND 0.02464f
C11935 VPWR.t1501 VGND 0.02189f
C11936 VPWR.n791 VGND 0.06768f
C11937 VPWR.n792 VGND 0.01329f
C11938 VPWR.n794 VGND 0.08003f
C11939 VPWR.t1494 VGND 0.08842f
C11940 VPWR.t1332 VGND 0.05805f
C11941 VPWR.t212 VGND 0.06817f
C11942 VPWR.t1495 VGND 0.02464f
C11943 VPWR.t213 VGND 0.02189f
C11944 VPWR.n795 VGND 0.06768f
C11945 VPWR.n796 VGND 0.01329f
C11946 VPWR.n798 VGND 0.08003f
C11947 VPWR.t1695 VGND 0.08842f
C11948 VPWR.t1338 VGND 0.05805f
C11949 VPWR.t1399 VGND 0.06817f
C11950 VPWR.t1696 VGND 0.02464f
C11951 VPWR.t1400 VGND 0.02189f
C11952 VPWR.n799 VGND 0.06768f
C11953 VPWR.n800 VGND 0.01329f
C11954 VPWR.n802 VGND 0.08003f
C11955 VPWR.t246 VGND 0.08842f
C11956 VPWR.t1337 VGND 0.05805f
C11957 VPWR.t69 VGND 0.06817f
C11958 VPWR.t247 VGND 0.02464f
C11959 VPWR.t70 VGND 0.02189f
C11960 VPWR.n803 VGND 0.06768f
C11961 VPWR.n804 VGND 0.01329f
C11962 VPWR.n806 VGND 0.08003f
C11963 VPWR.t520 VGND 0.08842f
C11964 VPWR.t1334 VGND 0.05805f
C11965 VPWR.t441 VGND 0.06817f
C11966 VPWR.t521 VGND 0.02464f
C11967 VPWR.t442 VGND 0.02189f
C11968 VPWR.n807 VGND 0.06768f
C11969 VPWR.n808 VGND 0.01329f
C11970 VPWR.n810 VGND 0.08003f
C11971 VPWR.t374 VGND 0.08842f
C11972 VPWR.t1378 VGND 0.05805f
C11973 VPWR.t479 VGND 0.06817f
C11974 VPWR.t375 VGND 0.02464f
C11975 VPWR.t480 VGND 0.02189f
C11976 VPWR.n811 VGND 0.06768f
C11977 VPWR.n812 VGND 0.01329f
C11978 VPWR.n814 VGND 0.08003f
C11979 VPWR.t473 VGND 0.08842f
C11980 VPWR.t1377 VGND 0.05805f
C11981 VPWR.t1447 VGND 0.06817f
C11982 VPWR.t474 VGND 0.02464f
C11983 VPWR.t1448 VGND 0.02189f
C11984 VPWR.n815 VGND 0.06768f
C11985 VPWR.n816 VGND 0.01329f
C11986 VPWR.n818 VGND 0.08003f
C11987 VPWR.t1359 VGND 0.08842f
C11988 VPWR.t1383 VGND 0.05805f
C11989 VPWR.t43 VGND 0.06817f
C11990 VPWR.t1360 VGND 0.02464f
C11991 VPWR.t44 VGND 0.02189f
C11992 VPWR.n819 VGND 0.06768f
C11993 VPWR.n820 VGND 0.01329f
C11994 VPWR.n822 VGND 0.08003f
C11995 VPWR.t162 VGND 0.08842f
C11996 VPWR.t1382 VGND 0.05805f
C11997 VPWR.t1200 VGND 0.06817f
C11998 VPWR.t163 VGND 0.02464f
C11999 VPWR.t1201 VGND 0.02189f
C12000 VPWR.n823 VGND 0.06768f
C12001 VPWR.n824 VGND 0.01329f
C12002 VPWR.n826 VGND 0.08003f
C12003 VPWR.t1566 VGND 0.08842f
C12004 VPWR.t1381 VGND 0.05805f
C12005 VPWR.t10 VGND 0.06817f
C12006 VPWR.t1567 VGND 0.02464f
C12007 VPWR.t11 VGND 0.02189f
C12008 VPWR.n827 VGND 0.06768f
C12009 VPWR.n828 VGND 0.01329f
C12010 VPWR.n830 VGND 0.08003f
C12011 VPWR.t1631 VGND 0.08842f
C12012 VPWR.t1336 VGND 0.05805f
C12013 VPWR.t786 VGND 0.0986f
C12014 VPWR.n831 VGND 0.05634f
C12015 VPWR.n832 VGND 0.01329f
C12016 VPWR.n833 VGND 0.10289f
C12017 VPWR.n834 VGND 0.75117f
C12018 VPWR.n835 VGND 0.10289f
C12019 VPWR.t209 VGND 0.02464f
C12020 VPWR.t610 VGND 0.02189f
C12021 VPWR.n836 VGND 0.06768f
C12022 VPWR.t395 VGND 0.06817f
C12023 VPWR.t488 VGND 0.02464f
C12024 VPWR.t396 VGND 0.02189f
C12025 VPWR.n837 VGND 0.06768f
C12026 VPWR.n838 VGND 0.10289f
C12027 VPWR.n839 VGND 0.10289f
C12028 VPWR.t52 VGND 0.02464f
C12029 VPWR.t973 VGND 0.02189f
C12030 VPWR.n840 VGND 0.06768f
C12031 VPWR.t296 VGND 0.06817f
C12032 VPWR.t1539 VGND 0.02464f
C12033 VPWR.t297 VGND 0.02189f
C12034 VPWR.n841 VGND 0.06768f
C12035 VPWR.n842 VGND 0.10289f
C12036 VPWR.n843 VGND 0.10289f
C12037 VPWR.t1121 VGND 0.02464f
C12038 VPWR.t1842 VGND 0.02189f
C12039 VPWR.n844 VGND 0.06768f
C12040 VPWR.t1508 VGND 0.06817f
C12041 VPWR.t359 VGND 0.02464f
C12042 VPWR.t1509 VGND 0.02189f
C12043 VPWR.n845 VGND 0.06768f
C12044 VPWR.n846 VGND 0.10289f
C12045 VPWR.n847 VGND 0.10289f
C12046 VPWR.t133 VGND 0.02464f
C12047 VPWR.t377 VGND 0.02189f
C12048 VPWR.n848 VGND 0.06768f
C12049 VPWR.t138 VGND 0.06817f
C12050 VPWR.t241 VGND 0.02464f
C12051 VPWR.t139 VGND 0.02189f
C12052 VPWR.n849 VGND 0.06768f
C12053 VPWR.n850 VGND 0.10289f
C12054 VPWR.n851 VGND 0.10289f
C12055 VPWR.t233 VGND 0.02464f
C12056 VPWR.t534 VGND 0.02189f
C12057 VPWR.n852 VGND 0.06768f
C12058 VPWR.t238 VGND 0.06817f
C12059 VPWR.t1274 VGND 0.02464f
C12060 VPWR.t239 VGND 0.02189f
C12061 VPWR.n853 VGND 0.06768f
C12062 VPWR.n854 VGND 0.10289f
C12063 VPWR.n855 VGND 0.10289f
C12064 VPWR.t1523 VGND 0.02464f
C12065 VPWR.t1280 VGND 0.02189f
C12066 VPWR.n856 VGND 0.06768f
C12067 VPWR.t1316 VGND 0.06817f
C12068 VPWR.t1061 VGND 0.02464f
C12069 VPWR.t1317 VGND 0.02189f
C12070 VPWR.n857 VGND 0.06768f
C12071 VPWR.n858 VGND 0.10289f
C12072 VPWR.n859 VGND 0.10289f
C12073 VPWR.t1178 VGND 0.02464f
C12074 VPWR.t1057 VGND 0.02189f
C12075 VPWR.n860 VGND 0.06768f
C12076 VPWR.t1151 VGND 0.06817f
C12077 VPWR.t1610 VGND 0.02464f
C12078 VPWR.t1152 VGND 0.02189f
C12079 VPWR.n861 VGND 0.06768f
C12080 VPWR.n862 VGND 0.10289f
C12081 VPWR.n863 VGND 0.10289f
C12082 VPWR.t311 VGND 0.02464f
C12083 VPWR.t1707 VGND 0.02189f
C12084 VPWR.n864 VGND 0.06768f
C12085 VPWR.t1469 VGND 0.10732f
C12086 VPWR.t1002 VGND 0.05805f
C12087 VPWR.t1615 VGND 0.06817f
C12088 VPWR.t1470 VGND 0.02464f
C12089 VPWR.t1616 VGND 0.02189f
C12090 VPWR.n865 VGND 0.06768f
C12091 VPWR.t1456 VGND 0.02464f
C12092 VPWR.t1104 VGND 0.02189f
C12093 VPWR.n866 VGND 0.06768f
C12094 VPWR.t1455 VGND 0.10732f
C12095 VPWR.t1396 VGND 0.05805f
C12096 VPWR.t1103 VGND 0.06817f
C12097 VPWR.t1630 VGND 0.02464f
C12098 VPWR.t794 VGND 0.02189f
C12099 VPWR.n867 VGND 0.06768f
C12100 VPWR.n868 VGND 0.01329f
C12101 VPWR.n869 VGND 0.05634f
C12102 VPWR.t793 VGND 0.0986f
C12103 VPWR.t1392 VGND 0.05805f
C12104 VPWR.t1629 VGND 0.08842f
C12105 VPWR.t1565 VGND 0.02464f
C12106 VPWR.t9 VGND 0.02189f
C12107 VPWR.n870 VGND 0.06768f
C12108 VPWR.n871 VGND 0.01329f
C12109 VPWR.n873 VGND 0.08003f
C12110 VPWR.t8 VGND 0.06817f
C12111 VPWR.t1920 VGND 0.05805f
C12112 VPWR.t1564 VGND 0.08842f
C12113 VPWR.t159 VGND 0.02464f
C12114 VPWR.t106 VGND 0.02189f
C12115 VPWR.n874 VGND 0.06768f
C12116 VPWR.n875 VGND 0.01329f
C12117 VPWR.n877 VGND 0.08003f
C12118 VPWR.t105 VGND 0.06817f
C12119 VPWR.t57 VGND 0.05805f
C12120 VPWR.t158 VGND 0.08842f
C12121 VPWR.t1358 VGND 0.02464f
C12122 VPWR.t42 VGND 0.02189f
C12123 VPWR.n878 VGND 0.06768f
C12124 VPWR.n879 VGND 0.01329f
C12125 VPWR.n881 VGND 0.08003f
C12126 VPWR.t41 VGND 0.06817f
C12127 VPWR.t58 VGND 0.05805f
C12128 VPWR.t1357 VGND 0.08842f
C12129 VPWR.t472 VGND 0.02464f
C12130 VPWR.t1446 VGND 0.02189f
C12131 VPWR.n882 VGND 0.06768f
C12132 VPWR.n883 VGND 0.01329f
C12133 VPWR.n885 VGND 0.08003f
C12134 VPWR.t1445 VGND 0.06817f
C12135 VPWR.t1916 VGND 0.05805f
C12136 VPWR.t471 VGND 0.08842f
C12137 VPWR.t373 VGND 0.02464f
C12138 VPWR.t478 VGND 0.02189f
C12139 VPWR.n886 VGND 0.06768f
C12140 VPWR.n887 VGND 0.01329f
C12141 VPWR.n889 VGND 0.08003f
C12142 VPWR.t477 VGND 0.06817f
C12143 VPWR.t1917 VGND 0.05805f
C12144 VPWR.t372 VGND 0.08842f
C12145 VPWR.t519 VGND 0.02464f
C12146 VPWR.t440 VGND 0.02189f
C12147 VPWR.n890 VGND 0.06768f
C12148 VPWR.n891 VGND 0.01329f
C12149 VPWR.n893 VGND 0.08003f
C12150 VPWR.t439 VGND 0.06817f
C12151 VPWR.t61 VGND 0.05805f
C12152 VPWR.t518 VGND 0.08842f
C12153 VPWR.t269 VGND 0.02464f
C12154 VPWR.t68 VGND 0.02189f
C12155 VPWR.n894 VGND 0.06768f
C12156 VPWR.n895 VGND 0.01329f
C12157 VPWR.n897 VGND 0.08003f
C12158 VPWR.t67 VGND 0.06817f
C12159 VPWR.t1393 VGND 0.05805f
C12160 VPWR.t268 VGND 0.08842f
C12161 VPWR.t1694 VGND 0.02464f
C12162 VPWR.t1398 VGND 0.02189f
C12163 VPWR.n898 VGND 0.06768f
C12164 VPWR.n899 VGND 0.01329f
C12165 VPWR.n901 VGND 0.08003f
C12166 VPWR.t1397 VGND 0.06817f
C12167 VPWR.t1394 VGND 0.05805f
C12168 VPWR.t1693 VGND 0.08842f
C12169 VPWR.t1493 VGND 0.02464f
C12170 VPWR.t211 VGND 0.02189f
C12171 VPWR.n902 VGND 0.06768f
C12172 VPWR.n903 VGND 0.01329f
C12173 VPWR.n905 VGND 0.08003f
C12174 VPWR.t210 VGND 0.06817f
C12175 VPWR.t59 VGND 0.05805f
C12176 VPWR.t1492 VGND 0.08842f
C12177 VPWR.t1700 VGND 0.02464f
C12178 VPWR.t1499 VGND 0.02189f
C12179 VPWR.n906 VGND 0.06768f
C12180 VPWR.n907 VGND 0.01329f
C12181 VPWR.n909 VGND 0.08003f
C12182 VPWR.t1498 VGND 0.06817f
C12183 VPWR.t60 VGND 0.05805f
C12184 VPWR.t1699 VGND 0.08842f
C12185 VPWR.t1063 VGND 0.02464f
C12186 VPWR.t1557 VGND 0.02189f
C12187 VPWR.n910 VGND 0.06768f
C12188 VPWR.n911 VGND 0.01329f
C12189 VPWR.n913 VGND 0.08003f
C12190 VPWR.t1556 VGND 0.06817f
C12191 VPWR.t1395 VGND 0.05805f
C12192 VPWR.t1062 VGND 0.08842f
C12193 VPWR.t1148 VGND 0.02464f
C12194 VPWR.t151 VGND 0.02189f
C12195 VPWR.n914 VGND 0.06768f
C12196 VPWR.n915 VGND 0.01329f
C12197 VPWR.n917 VGND 0.08003f
C12198 VPWR.t150 VGND 0.06817f
C12199 VPWR.t1918 VGND 0.05805f
C12200 VPWR.t1147 VGND 0.08842f
C12201 VPWR.t515 VGND 0.02464f
C12202 VPWR.t1184 VGND 0.02189f
C12203 VPWR.n918 VGND 0.06768f
C12204 VPWR.n919 VGND 0.01329f
C12205 VPWR.n921 VGND 0.08003f
C12206 VPWR.t1183 VGND 0.06817f
C12207 VPWR.t1919 VGND 0.05805f
C12208 VPWR.t514 VGND 0.08842f
C12209 VPWR.t554 VGND 0.02464f
C12210 VPWR.t1650 VGND 0.02189f
C12211 VPWR.n922 VGND 0.06768f
C12212 VPWR.n923 VGND 0.01329f
C12213 VPWR.n925 VGND 0.08003f
C12214 VPWR.t1649 VGND 0.06817f
C12215 VPWR.t62 VGND 0.05805f
C12216 VPWR.t553 VGND 0.08842f
C12217 VPWR.n926 VGND 0.08003f
C12218 VPWR.n928 VGND 0.01329f
C12219 VPWR.n929 VGND 0.10289f
C12220 VPWR.n930 VGND 0.74646f
C12221 VPWR.n931 VGND 0.10289f
C12222 VPWR.t1462 VGND 0.02464f
C12223 VPWR.t992 VGND 0.02189f
C12224 VPWR.n932 VGND 0.06768f
C12225 VPWR.t1461 VGND 0.10732f
C12226 VPWR.t1921 VGND 0.05805f
C12227 VPWR.t991 VGND 0.06817f
C12228 VPWR.t1542 VGND 0.08842f
C12229 VPWR.t17 VGND 0.02464f
C12230 VPWR.t1551 VGND 0.02189f
C12231 VPWR.n933 VGND 0.06768f
C12232 VPWR.n934 VGND 0.10289f
C12233 VPWR.n935 VGND 0.10289f
C12234 VPWR.t1543 VGND 0.02464f
C12235 VPWR.t1136 VGND 0.02189f
C12236 VPWR.n936 VGND 0.06768f
C12237 VPWR.t1925 VGND 0.05805f
C12238 VPWR.t1135 VGND 0.06817f
C12239 VPWR.t1048 VGND 0.08842f
C12240 VPWR.t1160 VGND 0.02464f
C12241 VPWR.t1067 VGND 0.02189f
C12242 VPWR.n937 VGND 0.06768f
C12243 VPWR.n938 VGND 0.10289f
C12244 VPWR.n939 VGND 0.10289f
C12245 VPWR.t1049 VGND 0.02464f
C12246 VPWR.t118 VGND 0.02189f
C12247 VPWR.n940 VGND 0.06768f
C12248 VPWR.t29 VGND 0.05805f
C12249 VPWR.t117 VGND 0.06817f
C12250 VPWR.t1486 VGND 0.08842f
C12251 VPWR.t110 VGND 0.02464f
C12252 VPWR.t1264 VGND 0.02189f
C12253 VPWR.n941 VGND 0.06768f
C12254 VPWR.n942 VGND 0.10289f
C12255 VPWR.n943 VGND 0.10289f
C12256 VPWR.t1487 VGND 0.02464f
C12257 VPWR.t1686 VGND 0.02189f
C12258 VPWR.n944 VGND 0.06768f
C12259 VPWR.t1329 VGND 0.05805f
C12260 VPWR.t1685 VGND 0.06817f
C12261 VPWR.t274 VGND 0.08842f
C12262 VPWR.t1866 VGND 0.02464f
C12263 VPWR.t253 VGND 0.02189f
C12264 VPWR.n945 VGND 0.06768f
C12265 VPWR.n946 VGND 0.10289f
C12266 VPWR.n947 VGND 0.10289f
C12267 VPWR.t275 VGND 0.02464f
C12268 VPWR.t325 VGND 0.02189f
C12269 VPWR.n948 VGND 0.06768f
C12270 VPWR.t27 VGND 0.05805f
C12271 VPWR.t324 VGND 0.06817f
C12272 VPWR.t384 VGND 0.08842f
C12273 VPWR.t317 VGND 0.02464f
C12274 VPWR.t410 VGND 0.02189f
C12275 VPWR.n949 VGND 0.06768f
C12276 VPWR.n950 VGND 0.10289f
C12277 VPWR.n951 VGND 0.10289f
C12278 VPWR.t385 VGND 0.02464f
C12279 VPWR.t1754 VGND 0.02189f
C12280 VPWR.n952 VGND 0.06768f
C12281 VPWR.t1923 VGND 0.05805f
C12282 VPWR.t1753 VGND 0.06817f
C12283 VPWR.t960 VGND 0.08842f
C12284 VPWR.t1746 VGND 0.02464f
C12285 VPWR.t971 VGND 0.02189f
C12286 VPWR.n953 VGND 0.06768f
C12287 VPWR.n954 VGND 0.10289f
C12288 VPWR.n955 VGND 0.10289f
C12289 VPWR.t961 VGND 0.02464f
C12290 VPWR.t171 VGND 0.02189f
C12291 VPWR.n956 VGND 0.06768f
C12292 VPWR.t1328 VGND 0.05805f
C12293 VPWR.t170 VGND 0.06817f
C12294 VPWR.t1418 VGND 0.08842f
C12295 VPWR.t289 VGND 0.02464f
C12296 VPWR.t1429 VGND 0.02189f
C12297 VPWR.n957 VGND 0.06768f
C12298 VPWR.n958 VGND 0.10289f
C12299 VPWR.n959 VGND 0.10289f
C12300 VPWR.t1419 VGND 0.02464f
C12301 VPWR.t1634 VGND 0.02189f
C12302 VPWR.n960 VGND 0.06768f
C12303 VPWR.t1326 VGND 0.05805f
C12304 VPWR.t1633 VGND 0.06817f
C12305 VPWR.t197 VGND 0.02464f
C12306 VPWR.t902 VGND 0.02189f
C12307 VPWR.n961 VGND 0.06768f
C12308 VPWR.t1642 VGND 0.02464f
C12309 VPWR.t754 VGND 0.02189f
C12310 VPWR.n962 VGND 0.06768f
C12311 VPWR.t1449 VGND 0.10732f
C12312 VPWR.t1626 VGND 0.05805f
C12313 VPWR.t87 VGND 0.06817f
C12314 VPWR.t1450 VGND 0.02464f
C12315 VPWR.t88 VGND 0.02189f
C12316 VPWR.n963 VGND 0.06768f
C12317 VPWR.n964 VGND 0.01329f
C12318 VPWR.n966 VGND 0.08003f
C12319 VPWR.t1101 VGND 0.08842f
C12320 VPWR.t1625 VGND 0.05805f
C12321 VPWR.t124 VGND 0.06817f
C12322 VPWR.t1102 VGND 0.02464f
C12323 VPWR.t125 VGND 0.02189f
C12324 VPWR.n967 VGND 0.06768f
C12325 VPWR.n968 VGND 0.01329f
C12326 VPWR.n970 VGND 0.08003f
C12327 VPWR.t1653 VGND 0.08842f
C12328 VPWR.t84 VGND 0.05805f
C12329 VPWR.t1171 VGND 0.06817f
C12330 VPWR.t1654 VGND 0.02464f
C12331 VPWR.t1172 VGND 0.02189f
C12332 VPWR.n971 VGND 0.06768f
C12333 VPWR.n972 VGND 0.01329f
C12334 VPWR.n974 VGND 0.08003f
C12335 VPWR.t1137 VGND 0.08842f
C12336 VPWR.t83 VGND 0.05805f
C12337 VPWR.t1025 VGND 0.06817f
C12338 VPWR.t1138 VGND 0.02464f
C12339 VPWR.t1026 VGND 0.02189f
C12340 VPWR.n975 VGND 0.06768f
C12341 VPWR.n976 VGND 0.01329f
C12342 VPWR.n978 VGND 0.08003f
C12343 VPWR.t1074 VGND 0.08842f
C12344 VPWR.t80 VGND 0.05805f
C12345 VPWR.t1575 VGND 0.06817f
C12346 VPWR.t1075 VGND 0.02464f
C12347 VPWR.t1576 VGND 0.02189f
C12348 VPWR.n979 VGND 0.06768f
C12349 VPWR.n980 VGND 0.01329f
C12350 VPWR.n982 VGND 0.08003f
C12351 VPWR.t1560 VGND 0.08842f
C12352 VPWR.t1623 VGND 0.05805f
C12353 VPWR.t1285 VGND 0.06817f
C12354 VPWR.t1561 VGND 0.02464f
C12355 VPWR.t1286 VGND 0.02189f
C12356 VPWR.n983 VGND 0.06768f
C12357 VPWR.n984 VGND 0.01329f
C12358 VPWR.n986 VGND 0.08003f
C12359 VPWR.t1502 VGND 0.08842f
C12360 VPWR.t1660 VGND 0.05805f
C12361 VPWR.t218 VGND 0.06817f
C12362 VPWR.t1503 VGND 0.02464f
C12363 VPWR.t219 VGND 0.02189f
C12364 VPWR.n987 VGND 0.06768f
C12365 VPWR.n988 VGND 0.01329f
C12366 VPWR.n990 VGND 0.08003f
C12367 VPWR.t214 VGND 0.08842f
C12368 VPWR.t79 VGND 0.05805f
C12369 VPWR.t1403 VGND 0.06817f
C12370 VPWR.t215 VGND 0.02464f
C12371 VPWR.t1404 VGND 0.02189f
C12372 VPWR.n991 VGND 0.06768f
C12373 VPWR.n992 VGND 0.01329f
C12374 VPWR.n994 VGND 0.08003f
C12375 VPWR.t254 VGND 0.08842f
C12376 VPWR.t78 VGND 0.05805f
C12377 VPWR.t75 VGND 0.06817f
C12378 VPWR.t255 VGND 0.02464f
C12379 VPWR.t76 VGND 0.02189f
C12380 VPWR.n995 VGND 0.06768f
C12381 VPWR.n996 VGND 0.01329f
C12382 VPWR.n998 VGND 0.08003f
C12383 VPWR.t71 VGND 0.08842f
C12384 VPWR.t1624 VGND 0.05805f
C12385 VPWR.t449 VGND 0.06817f
C12386 VPWR.t72 VGND 0.02464f
C12387 VPWR.t450 VGND 0.02189f
C12388 VPWR.n999 VGND 0.06768f
C12389 VPWR.n1000 VGND 0.01329f
C12390 VPWR.n1002 VGND 0.08003f
C12391 VPWR.t437 VGND 0.08842f
C12392 VPWR.t82 VGND 0.05805f
C12393 VPWR.t1731 VGND 0.06817f
C12394 VPWR.t438 VGND 0.02464f
C12395 VPWR.t1732 VGND 0.02189f
C12396 VPWR.n1003 VGND 0.06768f
C12397 VPWR.n1004 VGND 0.01329f
C12398 VPWR.n1006 VGND 0.08003f
C12399 VPWR.t481 VGND 0.08842f
C12400 VPWR.t81 VGND 0.05805f
C12401 VPWR.t1901 VGND 0.06817f
C12402 VPWR.t482 VGND 0.02464f
C12403 VPWR.t1902 VGND 0.02189f
C12404 VPWR.n1007 VGND 0.06768f
C12405 VPWR.n1008 VGND 0.01329f
C12406 VPWR.n1010 VGND 0.08003f
C12407 VPWR.t1443 VGND 0.08842f
C12408 VPWR.t1659 VGND 0.05805f
C12409 VPWR.t47 VGND 0.06817f
C12410 VPWR.t1444 VGND 0.02464f
C12411 VPWR.t48 VGND 0.02189f
C12412 VPWR.n1011 VGND 0.06768f
C12413 VPWR.n1012 VGND 0.01329f
C12414 VPWR.n1014 VGND 0.08003f
C12415 VPWR.t172 VGND 0.08842f
C12416 VPWR.t1658 VGND 0.05805f
C12417 VPWR.t1581 VGND 0.06817f
C12418 VPWR.t173 VGND 0.02464f
C12419 VPWR.t1582 VGND 0.02189f
C12420 VPWR.n1015 VGND 0.06768f
C12421 VPWR.n1016 VGND 0.01329f
C12422 VPWR.n1018 VGND 0.08003f
C12423 VPWR.t103 VGND 0.08842f
C12424 VPWR.t1657 VGND 0.05805f
C12425 VPWR.t204 VGND 0.06817f
C12426 VPWR.t104 VGND 0.02464f
C12427 VPWR.t205 VGND 0.02189f
C12428 VPWR.n1019 VGND 0.06768f
C12429 VPWR.n1020 VGND 0.01329f
C12430 VPWR.n1022 VGND 0.08003f
C12431 VPWR.t1641 VGND 0.08842f
C12432 VPWR.t77 VGND 0.05805f
C12433 VPWR.t753 VGND 0.0986f
C12434 VPWR.n1023 VGND 0.05634f
C12435 VPWR.n1024 VGND 0.01329f
C12436 VPWR.n1025 VGND 0.10289f
C12437 VPWR.n1026 VGND 4.32396f
C12438 VPWR.n1027 VGND 0.04856f
C12439 VPWR.n1028 VGND -0.0138f
C12440 VPWR.n1029 VGND 0.0225f
C12441 VPWR.t757 VGND 0.01981f
C12442 VPWR.n1031 VGND 0.04233f
C12443 VPWR.t865 VGND 0.02189f
C12444 VPWR.n1032 VGND 0.0347f
C12445 VPWR.t1643 VGND 0.06817f
C12446 VPWR.n1033 VGND 0.0225f
C12447 VPWR.t649 VGND 0.01981f
C12448 VPWR.n1035 VGND 0.04233f
C12449 VPWR.t1644 VGND 0.02189f
C12450 VPWR.n1036 VGND 0.0347f
C12451 VPWR.n1037 VGND -0.0138f
C12452 VPWR.n1038 VGND 0.04856f
C12453 VPWR.n1039 VGND 0.02048f
C12454 VPWR.n1040 VGND 0.01403f
C12455 VPWR.n1041 VGND 0.04617f
C12456 VPWR.n1042 VGND 0.07207f
C12457 VPWR.n1043 VGND 0.04023f
C12458 VPWR.n1044 VGND 0.04856f
C12459 VPWR.n1045 VGND -0.0138f
C12460 VPWR.n1046 VGND 0.0225f
C12461 VPWR.t735 VGND 0.01981f
C12462 VPWR.n1048 VGND 0.04233f
C12463 VPWR.t498 VGND 0.02189f
C12464 VPWR.n1049 VGND 0.0347f
C12465 VPWR.t497 VGND 0.06817f
C12466 VPWR.t598 VGND 0.08842f
C12467 VPWR.n1050 VGND 0.0225f
C12468 VPWR.t776 VGND 0.01981f
C12469 VPWR.n1052 VGND 0.04233f
C12470 VPWR.t179 VGND 0.02189f
C12471 VPWR.n1053 VGND 0.0347f
C12472 VPWR.n1055 VGND 0.14325f
C12473 VPWR.n1056 VGND 0.06176f
C12474 VPWR.n1057 VGND 0.02542f
C12475 VPWR.t829 VGND 0.02464f
C12476 VPWR.t821 VGND 0.02189f
C12477 VPWR.n1058 VGND 0.06768f
C12478 VPWR.t820 VGND 0.06817f
C12479 VPWR.t576 VGND 0.08842f
C12480 VPWR.t857 VGND 0.02464f
C12481 VPWR.t849 VGND 0.02189f
C12482 VPWR.n1059 VGND 0.06768f
C12483 VPWR.t577 VGND 0.02464f
C12484 VPWR.t700 VGND 0.02189f
C12485 VPWR.n1061 VGND 0.06768f
C12486 VPWR.t572 VGND 0.05805f
C12487 VPWR.t699 VGND 0.0986f
C12488 VPWR.n1062 VGND 0.05631f
C12489 VPWR.n1063 VGND 0.01256f
C12490 VPWR.n1064 VGND 0.02213f
C12491 VPWR.n1065 VGND 0.02429f
C12492 VPWR.n1067 VGND 0.01347f
C12493 VPWR.n1068 VGND 0.13004f
C12494 VPWR.n1069 VGND 0.02213f
C12495 VPWR.n1070 VGND 0.02429f
C12496 VPWR.n1071 VGND 0.01268f
C12497 VPWR.n1074 VGND 0.01268f
C12498 VPWR.n1076 VGND 0.02047f
C12499 VPWR.n1077 VGND 0.02084f
C12500 VPWR.n1078 VGND 0.01347f
C12501 VPWR.n1079 VGND 0.13004f
C12502 VPWR.n1080 VGND 0.02213f
C12503 VPWR.n1081 VGND 0.02429f
C12504 VPWR.n1082 VGND 0.01268f
C12505 VPWR.n1084 VGND 0.01268f
C12506 VPWR.n1086 VGND 0.02047f
C12507 VPWR.n1087 VGND 0.02084f
C12508 VPWR.n1088 VGND 0.01347f
C12509 VPWR.n1089 VGND 0.13004f
C12510 VPWR.n1090 VGND 0.02213f
C12511 VPWR.n1091 VGND 0.02429f
C12512 VPWR.n1092 VGND 0.01268f
C12513 VPWR.n1094 VGND 0.01268f
C12514 VPWR.n1096 VGND 0.02047f
C12515 VPWR.n1097 VGND 0.02084f
C12516 VPWR.n1098 VGND 0.01347f
C12517 VPWR.n1099 VGND 0.13004f
C12518 VPWR.n1100 VGND 0.02213f
C12519 VPWR.n1101 VGND 0.02429f
C12520 VPWR.n1102 VGND 0.01268f
C12521 VPWR.n1104 VGND 0.01268f
C12522 VPWR.n1106 VGND 0.02047f
C12523 VPWR.n1107 VGND 0.02084f
C12524 VPWR.n1108 VGND 0.01347f
C12525 VPWR.n1109 VGND 0.01963f
C12526 VPWR.n1110 VGND 0.02213f
C12527 VPWR.n1111 VGND 0.02429f
C12528 VPWR.n1112 VGND 0.01347f
C12529 VPWR.n1114 VGND 0.02304f
C12530 VPWR.n1115 VGND 0.01456f
C12531 VPWR.n1116 VGND 0.02047f
C12532 VPWR.n1117 VGND 0.02084f
C12533 VPWR.n1118 VGND 0.01313f
C12534 VPWR.n1119 VGND 0.02213f
C12535 VPWR.n1120 VGND 0.02429f
C12536 VPWR.t878 VGND 0.02464f
C12537 VPWR.t596 VGND 0.02189f
C12538 VPWR.n1122 VGND 0.06768f
C12539 VPWR.t877 VGND 0.10732f
C12540 VPWR.t867 VGND 0.05805f
C12541 VPWR.t595 VGND 0.06817f
C12542 VPWR.t747 VGND 0.08842f
C12543 VPWR.t646 VGND 0.02464f
C12544 VPWR.t732 VGND 0.02189f
C12545 VPWR.n1123 VGND 0.06768f
C12546 VPWR.n1125 VGND 0.02304f
C12547 VPWR.n1126 VGND 0.02731f
C12548 VPWR.n1127 VGND 0.02542f
C12549 VPWR.n1128 VGND 0.10289f
C12550 VPWR.n1130 VGND 0.01329f
C12551 VPWR.n1131 VGND 0.04856f
C12552 VPWR.n1132 VGND 0.04023f
C12553 VPWR.n1133 VGND 0.02048f
C12554 VPWR.n1134 VGND 0.01403f
C12555 VPWR.n1135 VGND 0.04617f
C12556 VPWR.n1136 VGND 0.07207f
C12557 VPWR.n1137 VGND 0.04856f
C12558 VPWR.n1138 VGND 0.04856f
C12559 VPWR.n1139 VGND 0.04856f
C12560 VPWR.n1140 VGND 0.04856f
C12561 VPWR.n1141 VGND 0.04856f
C12562 VPWR.n1142 VGND 0.04856f
C12563 VPWR.n1143 VGND 0.04023f
C12564 VPWR.n1145 VGND -0.0138f
C12565 VPWR.n1146 VGND 0.0225f
C12566 VPWR.t862 VGND 0.01981f
C12567 VPWR.n1148 VGND 0.04233f
C12568 VPWR.t416 VGND 0.02189f
C12569 VPWR.n1149 VGND 0.0347f
C12570 VPWR.t415 VGND 0.06817f
C12571 VPWR.t607 VGND 0.05805f
C12572 VPWR.t734 VGND 0.08842f
C12573 VPWR.n1150 VGND 0.0225f
C12574 VPWR.t605 VGND 0.01981f
C12575 VPWR.n1152 VGND 0.04233f
C12576 VPWR.t201 VGND 0.02189f
C12577 VPWR.n1153 VGND 0.0347f
C12578 VPWR.n1156 VGND 0.0225f
C12579 VPWR.t846 VGND 0.01981f
C12580 VPWR.n1158 VGND 0.04233f
C12581 VPWR.t1114 VGND 0.02189f
C12582 VPWR.n1159 VGND 0.0347f
C12583 VPWR.t956 VGND 0.06817f
C12584 VPWR.n1160 VGND 0.0225f
C12585 VPWR.t705 VGND 0.01981f
C12586 VPWR.n1162 VGND 0.04233f
C12587 VPWR.t957 VGND 0.02189f
C12588 VPWR.n1163 VGND 0.0347f
C12589 VPWR.n1166 VGND 0.0225f
C12590 VPWR.t583 VGND 0.01981f
C12591 VPWR.n1168 VGND 0.04233f
C12592 VPWR.t1692 VGND 0.02189f
C12593 VPWR.n1169 VGND 0.0347f
C12594 VPWR.t1762 VGND 0.06817f
C12595 VPWR.n1170 VGND 0.0225f
C12596 VPWR.t832 VGND 0.01981f
C12597 VPWR.n1172 VGND 0.04233f
C12598 VPWR.t1763 VGND 0.02189f
C12599 VPWR.n1173 VGND 0.0347f
C12600 VPWR.n1176 VGND 0.02304f
C12601 VPWR.n1177 VGND 0.02731f
C12602 VPWR.n1178 VGND 0.02542f
C12603 VPWR.t631 VGND 0.02464f
C12604 VPWR.t626 VGND 0.02189f
C12605 VPWR.n1179 VGND 0.06768f
C12606 VPWR.t737 VGND 0.05805f
C12607 VPWR.t744 VGND 0.06817f
C12608 VPWR.t748 VGND 0.02464f
C12609 VPWR.t745 VGND 0.02189f
C12610 VPWR.n1180 VGND 0.06768f
C12611 VPWR.n1182 VGND 0.08003f
C12612 VPWR.t912 VGND 0.08842f
C12613 VPWR.t778 VGND 0.05805f
C12614 VPWR.t904 VGND 0.06817f
C12615 VPWR.t913 VGND 0.02464f
C12616 VPWR.t905 VGND 0.02189f
C12617 VPWR.n1183 VGND 0.06768f
C12618 VPWR.n1185 VGND 0.08003f
C12619 VPWR.t630 VGND 0.08842f
C12620 VPWR.t886 VGND 0.05805f
C12621 VPWR.t625 VGND 0.06817f
C12622 VPWR.t702 VGND 0.05805f
C12623 VPWR.t828 VGND 0.08842f
C12624 VPWR.t591 VGND 0.02464f
C12625 VPWR.t692 VGND 0.02189f
C12626 VPWR.n1186 VGND 0.06768f
C12627 VPWR.n1188 VGND 0.08003f
C12628 VPWR.t691 VGND 0.06817f
C12629 VPWR.t676 VGND 0.05805f
C12630 VPWR.t590 VGND 0.08842f
C12631 VPWR.t570 VGND 0.02464f
C12632 VPWR.t948 VGND 0.02189f
C12633 VPWR.n1189 VGND 0.06768f
C12634 VPWR.n1191 VGND 0.08003f
C12635 VPWR.t947 VGND 0.06817f
C12636 VPWR.t826 VGND 0.05805f
C12637 VPWR.t569 VGND 0.08842f
C12638 VPWR.t824 VGND 0.02464f
C12639 VPWR.t929 VGND 0.02189f
C12640 VPWR.n1192 VGND 0.06768f
C12641 VPWR.n1194 VGND 0.02304f
C12642 VPWR.n1195 VGND 0.02731f
C12643 VPWR.n1196 VGND 0.02542f
C12644 VPWR.n1197 VGND 0.01268f
C12645 VPWR.n1199 VGND 0.08003f
C12646 VPWR.t928 VGND 0.06817f
C12647 VPWR.t804 VGND 0.05805f
C12648 VPWR.t823 VGND 0.08842f
C12649 VPWR.t697 VGND 0.02464f
C12650 VPWR.t770 VGND 0.02189f
C12651 VPWR.n1200 VGND 0.06768f
C12652 VPWR.n1202 VGND 0.08003f
C12653 VPWR.t769 VGND 0.06817f
C12654 VPWR.t651 VGND 0.05805f
C12655 VPWR.t696 VGND 0.08842f
C12656 VPWR.t671 VGND 0.02464f
C12657 VPWR.t666 VGND 0.02189f
C12658 VPWR.n1203 VGND 0.06768f
C12659 VPWR.n1205 VGND 0.08003f
C12660 VPWR.t665 VGND 0.06817f
C12661 VPWR.t934 VGND 0.05805f
C12662 VPWR.t670 VGND 0.08842f
C12663 VPWR.t910 VGND 0.02464f
C12664 VPWR.t921 VGND 0.02189f
C12665 VPWR.n1206 VGND 0.06768f
C12666 VPWR.n1208 VGND 0.02304f
C12667 VPWR.n1209 VGND 0.02731f
C12668 VPWR.n1210 VGND 0.02542f
C12669 VPWR.n1211 VGND 0.01268f
C12670 VPWR.n1213 VGND 0.08003f
C12671 VPWR.t920 VGND 0.06817f
C12672 VPWR.t891 VGND 0.05805f
C12673 VPWR.t909 VGND 0.08842f
C12674 VPWR.t802 VGND 0.02464f
C12675 VPWR.t884 VGND 0.02189f
C12676 VPWR.n1214 VGND 0.06768f
C12677 VPWR.n1216 VGND 0.08003f
C12678 VPWR.t883 VGND 0.06817f
C12679 VPWR.t668 VGND 0.05805f
C12680 VPWR.t801 VGND 0.08842f
C12681 VPWR.t643 VGND 0.02464f
C12682 VPWR.t773 VGND 0.02189f
C12683 VPWR.n1217 VGND 0.06768f
C12684 VPWR.n1219 VGND 0.08003f
C12685 VPWR.t772 VGND 0.06817f
C12686 VPWR.t653 VGND 0.05805f
C12687 VPWR.t642 VGND 0.08842f
C12688 VPWR.n1220 VGND 0.08003f
C12689 VPWR.n1222 VGND 0.01268f
C12690 VPWR.n1224 VGND 0.0225f
C12691 VPWR.t810 VGND 0.01981f
C12692 VPWR.n1226 VGND 0.04233f
C12693 VPWR.t1606 VGND 0.02189f
C12694 VPWR.n1227 VGND 0.0347f
C12695 VPWR.t673 VGND 0.10732f
C12696 VPWR.t658 VGND 0.05805f
C12697 VPWR.t65 VGND 0.06817f
C12698 VPWR.n1228 VGND 0.0225f
C12699 VPWR.t674 VGND 0.01981f
C12700 VPWR.n1230 VGND 0.04233f
C12701 VPWR.t66 VGND 0.02189f
C12702 VPWR.n1231 VGND 0.0347f
C12703 VPWR.n1232 VGND -0.0138f
C12704 VPWR.n1233 VGND 0.03466f
C12705 VPWR.t417 VGND 0.72151f
C12706 VPWR.n1234 VGND 0.39351f
C12707 VPWR.t364 VGND 0.72151f
C12708 VPWR.n1235 VGND 0.30604f
C12709 VPWR.n1236 VGND 0.21505f
C12710 VPWR.t1129 VGND 0.04227f
C12711 VPWR.t1434 VGND 0.0106f
C12712 VPWR.t1194 VGND 0.0106f
C12713 VPWR.n1238 VGND 0.02326f
C12714 VPWR.t1195 VGND 0.0106f
C12715 VPWR.t1013 VGND 0.0106f
C12716 VPWR.n1239 VGND 0.02322f
C12717 VPWR.t1597 VGND 0.0106f
C12718 VPWR.t1596 VGND 0.0106f
C12719 VPWR.n1240 VGND 0.02322f
C12720 VPWR.n1241 VGND 0.07706f
C12721 VPWR.n1242 VGND 0.13446f
C12722 VPWR.n1243 VGND 0.04257f
C12723 VPWR.n1244 VGND 0.03127f
C12724 VPWR.t1593 VGND 0.0106f
C12725 VPWR.t1598 VGND 0.0106f
C12726 VPWR.n1245 VGND 0.02326f
C12727 VPWR.n1246 VGND 0.09541f
C12728 VPWR.n1248 VGND 0.01206f
C12729 VPWR.n1249 VGND 0.01413f
C12730 VPWR.n1250 VGND 0.02072f
C12731 VPWR.t1128 VGND 0.04227f
C12732 VPWR.n1251 VGND 0.11136f
C12733 VPWR.t1739 VGND 0.04226f
C12734 VPWR.t1208 VGND 0.04226f
C12735 VPWR.n1253 VGND 0.09943f
C12736 VPWR.n1254 VGND 0.2482f
C12737 VPWR.n1255 VGND 1.21348f
C12738 VPWR.n1256 VGND 0.03466f
C12739 VPWR.t335 VGND 0.72151f
C12740 VPWR.n1257 VGND 0.39351f
C12741 VPWR.t154 VGND 0.72151f
C12742 VPWR.n1258 VGND 0.30604f
C12743 VPWR.n1259 VGND 0.21698f
C12744 VPWR.t341 VGND 0.0106f
C12745 VPWR.t339 VGND 0.0106f
C12746 VPWR.n1261 VGND 0.02326f
C12747 VPWR.t338 VGND 0.0106f
C12748 VPWR.t336 VGND 0.0106f
C12749 VPWR.n1262 VGND 0.02322f
C12750 VPWR.t1300 VGND 0.0106f
C12751 VPWR.t1301 VGND 0.0106f
C12752 VPWR.n1263 VGND 0.02322f
C12753 VPWR.n1264 VGND 0.07706f
C12754 VPWR.n1265 VGND 0.13446f
C12755 VPWR.n1266 VGND 0.04257f
C12756 VPWR.n1267 VGND 0.03127f
C12757 VPWR.t155 VGND 0.0106f
C12758 VPWR.t157 VGND 0.0106f
C12759 VPWR.n1268 VGND 0.02326f
C12760 VPWR.n1269 VGND 0.09541f
C12761 VPWR.n1271 VGND 0.01206f
C12762 VPWR.n1272 VGND 0.01413f
C12763 VPWR.n1273 VGND 0.02034f
C12764 VPWR.t1130 VGND 0.04221f
C12765 VPWR.n1275 VGND 0.04512f
C12766 VPWR.t1836 VGND 0.0423f
C12767 VPWR.n1277 VGND 0.06737f
C12768 VPWR.n1278 VGND 0.2482f
C12769 VPWR.n1279 VGND 1.21348f
C12770 VPWR.n1280 VGND 0.03466f
C12771 VPWR.t302 VGND 0.72151f
C12772 VPWR.n1281 VGND 0.39351f
C12773 VPWR.t1029 VGND 0.72151f
C12774 VPWR.n1282 VGND 0.30604f
C12775 VPWR.n1283 VGND 0.21698f
C12776 VPWR.t1354 VGND 0.0106f
C12777 VPWR.t1352 VGND 0.0106f
C12778 VPWR.n1285 VGND 0.02326f
C12779 VPWR.t1351 VGND 0.0106f
C12780 VPWR.t1350 VGND 0.0106f
C12781 VPWR.n1286 VGND 0.02322f
C12782 VPWR.t1030 VGND 0.0106f
C12783 VPWR.t1037 VGND 0.0106f
C12784 VPWR.n1287 VGND 0.02322f
C12785 VPWR.n1288 VGND 0.07706f
C12786 VPWR.n1289 VGND 0.13446f
C12787 VPWR.n1290 VGND 0.04257f
C12788 VPWR.n1291 VGND 0.03127f
C12789 VPWR.t1034 VGND 0.0106f
C12790 VPWR.t1031 VGND 0.0106f
C12791 VPWR.n1292 VGND 0.02326f
C12792 VPWR.n1293 VGND 0.09541f
C12793 VPWR.n1295 VGND 0.01206f
C12794 VPWR.n1296 VGND 0.01413f
C12795 VPWR.n1297 VGND 0.02034f
C12796 VPWR.n1298 VGND 0.01034f
C12797 VPWR.t1740 VGND 0.0423f
C12798 VPWR.t1209 VGND 0.0423f
C12799 VPWR.n1300 VGND 0.12493f
C12800 VPWR.n1301 VGND 0.2482f
C12801 VPWR.n1302 VGND 1.21348f
C12802 VPWR.t977 VGND 0.04223f
C12803 VPWR.t951 VGND 0.0423f
C12804 VPWR.t979 VGND 0.04194f
C12805 VPWR.n1303 VGND 0.10875f
C12806 VPWR.t307 VGND 0.04146f
C12807 VPWR.n1304 VGND 0.0501f
C12808 VPWR.n1305 VGND 0.03466f
C12809 VPWR.t1730 VGND 0.03991f
C12810 VPWR.n1306 VGND 0.03796f
C12811 VPWR.t265 VGND 0.0106f
C12812 VPWR.t1765 VGND 0.0106f
C12813 VPWR.n1307 VGND 0.02315f
C12814 VPWR.t1758 VGND 0.03708f
C12815 VPWR.n1308 VGND 0.05562f
C12816 VPWR.n1309 VGND 0.03466f
C12817 VPWR.t304 VGND 0.04225f
C12818 VPWR.n1310 VGND 0.05319f
C12819 VPWR.n1311 VGND 0.02034f
C12820 VPWR.n1312 VGND 0.03466f
C12821 VPWR.t1767 VGND 0.0106f
C12822 VPWR.t1294 VGND 0.0106f
C12823 VPWR.n1314 VGND 0.02315f
C12824 VPWR.n1315 VGND 0.03393f
C12825 VPWR.n1317 VGND 0.02599f
C12826 VPWR.n1318 VGND 0.02599f
C12827 VPWR.n1319 VGND 0.03466f
C12828 VPWR.t261 VGND 0.0106f
C12829 VPWR.t143 VGND 0.0106f
C12830 VPWR.n1321 VGND 0.02315f
C12831 VPWR.n1322 VGND 0.02666f
C12832 VPWR.t419 VGND 0.0106f
C12833 VPWR.t1116 VGND 0.0106f
C12834 VPWR.n1323 VGND 0.02315f
C12835 VPWR.n1324 VGND 0.02946f
C12836 VPWR.n1326 VGND 0.03146f
C12837 VPWR.n1327 VGND 0.01187f
C12838 VPWR.t524 VGND 0.03554f
C12839 VPWR.t976 VGND 0.07996f
C12840 VPWR.t950 VGND 0.09329f
C12841 VPWR.t978 VGND 0.17324f
C12842 VPWR.t303 VGND 0.09321f
C12843 VPWR.t1293 VGND 0.10581f
C12844 VPWR.t1766 VGND 0.10287f
C12845 VPWR.t1764 VGND 0.16452f
C12846 VPWR.t264 VGND 0.13993f
C12847 VPWR.t1757 VGND 0.09329f
C12848 VPWR.t142 VGND 0.09329f
C12849 VPWR.t1115 VGND 0.09329f
C12850 VPWR.t260 VGND 0.09329f
C12851 VPWR.t418 VGND 0.09329f
C12852 VPWR.t1729 VGND 0.09329f
C12853 VPWR.t306 VGND 0.09217f
C12854 VPWR.n1329 VGND 0.31703f
C12855 VPWR.n1330 VGND 0.12882f
C12856 VPWR.n1331 VGND 0.01413f
C12857 VPWR.n1332 VGND 0.02599f
C12858 VPWR.n1333 VGND 0.03127f
C12859 VPWR.n1335 VGND 0.04701f
C12860 VPWR.n1336 VGND 0.23407f
C12861 VPWR.n1337 VGND 1.21348f
C12862 VPWR.t1516 VGND 0.04155f
C12863 VPWR.t1906 VGND 0.04143f
C12864 VPWR.t949 VGND 0.04226f
C12865 VPWR.n1338 VGND 0.05889f
C12866 VPWR.t1718 VGND 0.04034f
C12867 VPWR.t1599 VGND 0.04034f
C12868 VPWR.n1339 VGND 0.07319f
C12869 VPWR.n1340 VGND 0.03466f
C12870 VPWR.n1342 VGND 0.03466f
C12871 VPWR.t1435 VGND 0.0106f
C12872 VPWR.t1312 VGND 0.0106f
C12873 VPWR.n1343 VGND 0.02315f
C12874 VPWR.t1600 VGND 0.0106f
C12875 VPWR.t365 VGND 0.0106f
C12876 VPWR.n1344 VGND 0.02315f
C12877 VPWR.n1345 VGND 0.04717f
C12878 VPWR.t368 VGND 0.04225f
C12879 VPWR.t1295 VGND 0.04225f
C12880 VPWR.n1346 VGND 0.09738f
C12881 VPWR.n1347 VGND 0.02034f
C12882 VPWR.n1348 VGND 0.03466f
C12883 VPWR.t1297 VGND 0.0106f
C12884 VPWR.t1760 VGND 0.0106f
C12885 VPWR.n1350 VGND 0.02315f
C12886 VPWR.t386 VGND 0.0106f
C12887 VPWR.t22 VGND 0.0106f
C12888 VPWR.n1351 VGND 0.02315f
C12889 VPWR.n1352 VGND 0.05331f
C12890 VPWR.n1354 VGND 0.03466f
C12891 VPWR.n1355 VGND 0.03466f
C12892 VPWR.n1356 VGND 0.03466f
C12893 VPWR.t1014 VGND 0.0106f
C12894 VPWR.t1193 VGND 0.0106f
C12895 VPWR.n1358 VGND 0.02315f
C12896 VPWR.t1595 VGND 0.0106f
C12897 VPWR.t1594 VGND 0.0106f
C12898 VPWR.n1359 VGND 0.02315f
C12899 VPWR.n1360 VGND 0.04717f
C12900 VPWR.n1363 VGND 0.03466f
C12901 VPWR.n1364 VGND 0.02599f
C12902 VPWR.t367 VGND 0.72151f
C12903 VPWR.n1366 VGND 0.39351f
C12904 VPWR.t21 VGND 0.72151f
C12905 VPWR.n1367 VGND 0.30604f
C12906 VPWR.n1368 VGND 0.21505f
C12907 VPWR.n1369 VGND 0.01413f
C12908 VPWR.n1370 VGND 0.02599f
C12909 VPWR.n1371 VGND 0.03146f
C12910 VPWR.n1373 VGND 0.04309f
C12911 VPWR.n1374 VGND 0.05837f
C12912 VPWR.n1375 VGND 0.23388f
C12913 VPWR.n1376 VGND 1.21348f
C12914 VPWR.t1225 VGND 0.04221f
C12915 VPWR.t1 VGND 0.04221f
C12916 VPWR.n1377 VGND 0.01034f
C12917 VPWR.t337 VGND 0.04034f
C12918 VPWR.t156 VGND 0.04034f
C12919 VPWR.n1378 VGND 0.07319f
C12920 VPWR.n1379 VGND 0.03466f
C12921 VPWR.n1381 VGND 0.03466f
C12922 VPWR.t342 VGND 0.0106f
C12923 VPWR.t369 VGND 0.0106f
C12924 VPWR.n1382 VGND 0.02315f
C12925 VPWR.t1889 VGND 0.0106f
C12926 VPWR.t1296 VGND 0.0106f
C12927 VPWR.n1383 VGND 0.02315f
C12928 VPWR.n1384 VGND 0.04717f
C12929 VPWR.t1310 VGND 0.04225f
C12930 VPWR.t421 VGND 0.04225f
C12931 VPWR.n1385 VGND 0.09738f
C12932 VPWR.n1386 VGND 0.02034f
C12933 VPWR.n1387 VGND 0.03466f
C12934 VPWR.t388 VGND 0.0106f
C12935 VPWR.t24 VGND 0.0106f
C12936 VPWR.n1389 VGND 0.02315f
C12937 VPWR.t1311 VGND 0.0106f
C12938 VPWR.t1299 VGND 0.0106f
C12939 VPWR.n1390 VGND 0.02315f
C12940 VPWR.n1391 VGND 0.05331f
C12941 VPWR.n1393 VGND 0.03466f
C12942 VPWR.n1394 VGND 0.03466f
C12943 VPWR.n1395 VGND 0.03466f
C12944 VPWR.t343 VGND 0.0106f
C12945 VPWR.t340 VGND 0.0106f
C12946 VPWR.n1397 VGND 0.02315f
C12947 VPWR.t1888 VGND 0.0106f
C12948 VPWR.t1890 VGND 0.0106f
C12949 VPWR.n1398 VGND 0.02315f
C12950 VPWR.n1399 VGND 0.04717f
C12951 VPWR.n1402 VGND 0.03466f
C12952 VPWR.n1403 VGND 0.02599f
C12953 VPWR.t23 VGND 0.72151f
C12954 VPWR.n1405 VGND 0.39351f
C12955 VPWR.t0 VGND 0.72151f
C12956 VPWR.n1406 VGND 0.30604f
C12957 VPWR.n1407 VGND 0.21698f
C12958 VPWR.n1408 VGND 0.01413f
C12959 VPWR.n1409 VGND 0.02599f
C12960 VPWR.n1410 VGND 0.03146f
C12961 VPWR.n1412 VGND 0.08532f
C12962 VPWR.n1413 VGND 0.23765f
C12963 VPWR.n1414 VGND 1.21348f
C12964 VPWR.t1353 VGND 0.04034f
C12965 VPWR.t1032 VGND 0.04034f
C12966 VPWR.n1415 VGND 0.07319f
C12967 VPWR.n1416 VGND 0.03466f
C12968 VPWR.n1418 VGND 0.03466f
C12969 VPWR.t1348 VGND 0.0106f
C12970 VPWR.t1313 VGND 0.0106f
C12971 VPWR.n1419 VGND 0.02315f
C12972 VPWR.t1033 VGND 0.0106f
C12973 VPWR.t301 VGND 0.0106f
C12974 VPWR.n1420 VGND 0.02315f
C12975 VPWR.n1421 VGND 0.04717f
C12976 VPWR.t371 VGND 0.04225f
C12977 VPWR.t1117 VGND 0.04225f
C12978 VPWR.n1422 VGND 0.09738f
C12979 VPWR.n1423 VGND 0.02034f
C12980 VPWR.n1424 VGND 0.03466f
C12981 VPWR.t1298 VGND 0.0106f
C12982 VPWR.t1761 VGND 0.0106f
C12983 VPWR.n1426 VGND 0.02315f
C12984 VPWR.t305 VGND 0.0106f
C12985 VPWR.t420 VGND 0.0106f
C12986 VPWR.n1427 VGND 0.02315f
C12987 VPWR.n1428 VGND 0.05331f
C12988 VPWR.n1430 VGND 0.03466f
C12989 VPWR.n1431 VGND 0.03466f
C12990 VPWR.n1432 VGND 0.03466f
C12991 VPWR.t1349 VGND 0.0106f
C12992 VPWR.t1347 VGND 0.0106f
C12993 VPWR.n1434 VGND 0.02315f
C12994 VPWR.t1036 VGND 0.0106f
C12995 VPWR.t1035 VGND 0.0106f
C12996 VPWR.n1435 VGND 0.02315f
C12997 VPWR.n1436 VGND 0.04717f
C12998 VPWR.n1439 VGND 0.03466f
C12999 VPWR.n1440 VGND 0.02599f
C13000 VPWR.t370 VGND 0.55347f
C13001 VPWR.n1442 VGND 0.31666f
C13002 VPWR.t300 VGND 0.55347f
C13003 VPWR.n1443 VGND 0.24813f
C13004 VPWR.n1444 VGND 0.20802f
C13005 VPWR.n1445 VGND 0.31801f
C13006 VPWR.n1446 VGND 4.62393f
C13007 VPWR.n1447 VGND 6.76927f
C13008 VPWR.n1448 VGND 0.06176f
C13009 VPWR.n1449 VGND 0.81338f
C13010 VPWR.n1450 VGND 0.74646f
C13011 VPWR.n1451 VGND 0.04794f
C13012 VPWR.n1452 VGND 0.04023f
C13013 VPWR.n1453 VGND 0.02048f
C13014 VPWR.n1454 VGND 0.01403f
C13015 VPWR.n1455 VGND 0.04617f
C13016 VPWR.n1456 VGND 0.0574f
C13017 VPWR.n1457 VGND 0.06785f
C13018 VPWR.n1458 VGND 0.02048f
C13019 VPWR.n1459 VGND 0.01403f
C13020 VPWR.n1460 VGND 0.04617f
C13021 VPWR.n1461 VGND 0.07207f
C13022 VPWR.n1462 VGND 0.06785f
C13023 VPWR.n1463 VGND 0.04856f
C13024 VPWR.n1464 VGND 0.04023f
C13025 VPWR.n1465 VGND 0.10289f
C13026 VPWR.n1466 VGND 0.01329f
C13027 VPWR.n1468 VGND 0.08003f
C13028 VPWR.t834 VGND 0.08842f
C13029 VPWR.t789 VGND 0.05805f
C13030 VPWR.t1532 VGND 0.06817f
C13031 VPWR.n1469 VGND 0.0225f
C13032 VPWR.t835 VGND 0.01981f
C13033 VPWR.n1471 VGND 0.04233f
C13034 VPWR.t1533 VGND 0.02189f
C13035 VPWR.n1472 VGND 0.0347f
C13036 VPWR.n1473 VGND 0.01329f
C13037 VPWR.n1475 VGND 0.08003f
C13038 VPWR.t936 VGND 0.08842f
C13039 VPWR.t918 VGND 0.05805f
C13040 VPWR.t1187 VGND 0.06817f
C13041 VPWR.n1476 VGND 0.0225f
C13042 VPWR.t937 VGND 0.01981f
C13043 VPWR.n1478 VGND 0.04233f
C13044 VPWR.t1188 VGND 0.02189f
C13045 VPWR.n1479 VGND 0.0347f
C13046 VPWR.n1481 VGND 0.08003f
C13047 VPWR.t707 VGND 0.08842f
C13048 VPWR.t574 VGND 0.05805f
C13049 VPWR.t1076 VGND 0.06817f
C13050 VPWR.n1482 VGND 0.0225f
C13051 VPWR.t708 VGND 0.01981f
C13052 VPWR.n1484 VGND 0.04233f
C13053 VPWR.t1077 VGND 0.02189f
C13054 VPWR.n1485 VGND 0.0347f
C13055 VPWR.n1487 VGND 0.06176f
C13056 VPWR.n1488 VGND -0.0138f
C13057 VPWR.n1489 VGND 0.10289f
C13058 VPWR.n1490 VGND 0.01329f
C13059 VPWR.n1492 VGND 0.08003f
C13060 VPWR.t809 VGND 0.08842f
C13061 VPWR.t684 VGND 0.05805f
C13062 VPWR.t1605 VGND 0.06817f
C13063 VPWR.t839 VGND 0.05805f
C13064 VPWR.t831 VGND 0.08842f
C13065 VPWR.n1493 VGND 0.08003f
C13066 VPWR.n1495 VGND 0.01329f
C13067 VPWR.n1496 VGND 0.04023f
C13068 VPWR.n1497 VGND 0.10289f
C13069 VPWR.n1498 VGND -0.0138f
C13070 VPWR.n1499 VGND 0.06176f
C13071 VPWR.n1500 VGND 0.06176f
C13072 VPWR.n1501 VGND -0.0138f
C13073 VPWR.n1502 VGND 0.04023f
C13074 VPWR.n1503 VGND 0.10289f
C13075 VPWR.n1504 VGND 0.01329f
C13076 VPWR.n1506 VGND 0.08003f
C13077 VPWR.t582 VGND 0.08842f
C13078 VPWR.t841 VGND 0.05805f
C13079 VPWR.t1691 VGND 0.06817f
C13080 VPWR.t689 VGND 0.05805f
C13081 VPWR.t704 VGND 0.08842f
C13082 VPWR.n1507 VGND 0.08003f
C13083 VPWR.n1509 VGND 0.01329f
C13084 VPWR.n1510 VGND 0.04023f
C13085 VPWR.n1511 VGND 0.10289f
C13086 VPWR.n1512 VGND -0.0138f
C13087 VPWR.n1513 VGND 0.06176f
C13088 VPWR.n1514 VGND 0.06176f
C13089 VPWR.n1515 VGND -0.0138f
C13090 VPWR.n1516 VGND 0.04023f
C13091 VPWR.n1517 VGND 0.10289f
C13092 VPWR.n1518 VGND 0.01329f
C13093 VPWR.n1520 VGND 0.08003f
C13094 VPWR.t845 VGND 0.08842f
C13095 VPWR.t719 VGND 0.05805f
C13096 VPWR.t1113 VGND 0.06817f
C13097 VPWR.t837 VGND 0.05805f
C13098 VPWR.t861 VGND 0.08842f
C13099 VPWR.n1521 VGND 0.08003f
C13100 VPWR.n1523 VGND 0.01329f
C13101 VPWR.n1524 VGND 0.04023f
C13102 VPWR.n1525 VGND 0.10289f
C13103 VPWR.n1526 VGND -0.0138f
C13104 VPWR.n1527 VGND 0.06176f
C13105 VPWR.n1528 VGND 0.06176f
C13106 VPWR.n1529 VGND 0.06176f
C13107 VPWR.n1530 VGND 0.06176f
C13108 VPWR.n1531 VGND -0.0138f
C13109 VPWR.n1532 VGND 0.10289f
C13110 VPWR.n1533 VGND 0.01329f
C13111 VPWR.n1535 VGND 0.08003f
C13112 VPWR.t200 VGND 0.06817f
C13113 VPWR.t588 VGND 0.05805f
C13114 VPWR.t604 VGND 0.08842f
C13115 VPWR.n1536 VGND 0.08003f
C13116 VPWR.n1538 VGND 0.01329f
C13117 VPWR.n1539 VGND 0.10289f
C13118 VPWR.n1540 VGND 0.04023f
C13119 VPWR.n1541 VGND 0.04856f
C13120 VPWR.n1542 VGND 0.06785f
C13121 VPWR.n1543 VGND 0.02048f
C13122 VPWR.n1544 VGND 0.01403f
C13123 VPWR.n1545 VGND 0.04617f
C13124 VPWR.n1546 VGND 0.07207f
C13125 VPWR.n1547 VGND 0.06785f
C13126 VPWR.n1548 VGND 0.02048f
C13127 VPWR.n1549 VGND 0.01403f
C13128 VPWR.n1550 VGND 0.04617f
C13129 VPWR.n1551 VGND 0.07207f
C13130 VPWR.n1552 VGND 0.06785f
C13131 VPWR.n1553 VGND 0.02048f
C13132 VPWR.n1554 VGND 0.01403f
C13133 VPWR.n1555 VGND 0.04617f
C13134 VPWR.n1556 VGND 0.07207f
C13135 VPWR.n1557 VGND 0.06785f
C13136 VPWR.n1558 VGND 0.02048f
C13137 VPWR.n1559 VGND 0.01403f
C13138 VPWR.n1560 VGND 0.04617f
C13139 VPWR.n1561 VGND 0.07207f
C13140 VPWR.n1562 VGND 0.06785f
C13141 VPWR.n1563 VGND 0.02048f
C13142 VPWR.n1564 VGND 0.01403f
C13143 VPWR.n1565 VGND 0.04617f
C13144 VPWR.n1566 VGND 0.07207f
C13145 VPWR.n1567 VGND 0.06785f
C13146 VPWR.n1568 VGND 0.02048f
C13147 VPWR.n1569 VGND 0.01403f
C13148 VPWR.n1570 VGND 0.04617f
C13149 VPWR.n1571 VGND 0.07207f
C13150 VPWR.n1572 VGND 0.06785f
C13151 VPWR.n1573 VGND 0.02048f
C13152 VPWR.n1574 VGND 0.01403f
C13153 VPWR.n1575 VGND 0.04617f
C13154 VPWR.n1576 VGND 0.07207f
C13155 VPWR.n1577 VGND 0.06785f
C13156 VPWR.n1578 VGND 0.02048f
C13157 VPWR.n1579 VGND 0.01403f
C13158 VPWR.n1580 VGND 0.04617f
C13159 VPWR.n1581 VGND 0.07207f
C13160 VPWR.n1582 VGND 0.06785f
C13161 VPWR.n1583 VGND 0.04856f
C13162 VPWR.n1584 VGND 0.04023f
C13163 VPWR.n1585 VGND 0.10289f
C13164 VPWR.n1586 VGND -0.0138f
C13165 VPWR.n1587 VGND 0.06176f
C13166 VPWR.n1588 VGND 0.06176f
C13167 VPWR.n1589 VGND -0.0138f
C13168 VPWR.n1591 VGND 0.01268f
C13169 VPWR.n1593 VGND 0.08003f
C13170 VPWR.t731 VGND 0.06817f
C13171 VPWR.t612 VGND 0.05805f
C13172 VPWR.t645 VGND 0.08842f
C13173 VPWR.n1594 VGND 0.08003f
C13174 VPWR.n1596 VGND 0.01268f
C13175 VPWR.n1597 VGND 0.02542f
C13176 VPWR.n1598 VGND 0.02304f
C13177 VPWR.n1599 VGND 0.02731f
C13178 VPWR.n1601 VGND 0.02047f
C13179 VPWR.n1602 VGND 0.02084f
C13180 VPWR.n1603 VGND 0.01313f
C13181 VPWR.n1605 VGND 0.01347f
C13182 VPWR.n1606 VGND 0.01763f
C13183 VPWR.n1607 VGND 0.17544f
C13184 VPWR.n1608 VGND 0.13004f
C13185 VPWR.n1609 VGND 0.01763f
C13186 VPWR.n1610 VGND 0.01313f
C13187 VPWR.n1611 VGND 0.02213f
C13188 VPWR.n1612 VGND 0.02429f
C13189 VPWR.n1613 VGND 0.02542f
C13190 VPWR.n1614 VGND 0.02304f
C13191 VPWR.n1615 VGND 0.02731f
C13192 VPWR.n1617 VGND 0.02047f
C13193 VPWR.n1618 VGND 0.02084f
C13194 VPWR.n1619 VGND 0.01347f
C13195 VPWR.n1620 VGND 0.01763f
C13196 VPWR.n1621 VGND 0.01313f
C13197 VPWR.n1622 VGND 0.02213f
C13198 VPWR.n1623 VGND 0.02429f
C13199 VPWR.n1624 VGND 0.02542f
C13200 VPWR.n1625 VGND 0.02304f
C13201 VPWR.n1626 VGND 0.02731f
C13202 VPWR.n1628 VGND 0.02047f
C13203 VPWR.n1629 VGND 0.02084f
C13204 VPWR.n1630 VGND 0.01313f
C13205 VPWR.n1632 VGND 0.01347f
C13206 VPWR.n1633 VGND 0.01763f
C13207 VPWR.n1634 VGND 0.13004f
C13208 VPWR.n1635 VGND 0.13004f
C13209 VPWR.n1636 VGND 0.01763f
C13210 VPWR.n1637 VGND 0.01313f
C13211 VPWR.n1638 VGND 0.02213f
C13212 VPWR.n1639 VGND 0.02429f
C13213 VPWR.n1640 VGND 0.02542f
C13214 VPWR.n1641 VGND 0.02304f
C13215 VPWR.n1642 VGND 0.02731f
C13216 VPWR.n1644 VGND 0.02047f
C13217 VPWR.n1645 VGND 0.02084f
C13218 VPWR.n1646 VGND 0.01347f
C13219 VPWR.n1647 VGND 0.01763f
C13220 VPWR.n1648 VGND 0.01313f
C13221 VPWR.n1649 VGND 0.02213f
C13222 VPWR.n1650 VGND 0.02429f
C13223 VPWR.n1651 VGND 0.02542f
C13224 VPWR.n1652 VGND 0.02304f
C13225 VPWR.n1653 VGND 0.02731f
C13226 VPWR.n1655 VGND 0.02047f
C13227 VPWR.n1656 VGND 0.02084f
C13228 VPWR.n1657 VGND 0.01313f
C13229 VPWR.n1659 VGND 0.01347f
C13230 VPWR.n1660 VGND 0.01763f
C13231 VPWR.n1661 VGND 0.13004f
C13232 VPWR.n1662 VGND 0.13004f
C13233 VPWR.n1663 VGND 0.01763f
C13234 VPWR.n1664 VGND 0.01313f
C13235 VPWR.n1665 VGND 0.02213f
C13236 VPWR.n1666 VGND 0.02429f
C13237 VPWR.n1667 VGND 0.02542f
C13238 VPWR.n1668 VGND 0.02304f
C13239 VPWR.n1669 VGND 0.02731f
C13240 VPWR.n1671 VGND 0.02047f
C13241 VPWR.n1672 VGND 0.02084f
C13242 VPWR.n1673 VGND 0.01347f
C13243 VPWR.n1674 VGND 0.01763f
C13244 VPWR.n1675 VGND 0.01313f
C13245 VPWR.n1676 VGND 0.02213f
C13246 VPWR.n1677 VGND 0.02429f
C13247 VPWR.n1678 VGND 0.02542f
C13248 VPWR.n1679 VGND 0.02304f
C13249 VPWR.n1680 VGND 0.02731f
C13250 VPWR.n1682 VGND 0.02047f
C13251 VPWR.n1683 VGND 0.02084f
C13252 VPWR.n1684 VGND 0.01313f
C13253 VPWR.n1686 VGND 0.01347f
C13254 VPWR.n1687 VGND 0.01763f
C13255 VPWR.n1688 VGND 0.13004f
C13256 VPWR.n1689 VGND 0.13004f
C13257 VPWR.n1690 VGND 0.01763f
C13258 VPWR.n1691 VGND 0.01313f
C13259 VPWR.n1692 VGND 0.02213f
C13260 VPWR.n1693 VGND 0.02429f
C13261 VPWR.n1694 VGND 0.02542f
C13262 VPWR.n1695 VGND 0.02304f
C13263 VPWR.n1696 VGND 0.02731f
C13264 VPWR.n1698 VGND 0.02047f
C13265 VPWR.n1699 VGND 0.02084f
C13266 VPWR.n1700 VGND 0.01347f
C13267 VPWR.n1701 VGND 0.01763f
C13268 VPWR.n1702 VGND 0.01313f
C13269 VPWR.n1703 VGND 0.02213f
C13270 VPWR.n1704 VGND 0.02429f
C13271 VPWR.n1705 VGND 0.02542f
C13272 VPWR.n1706 VGND 0.02304f
C13273 VPWR.n1707 VGND 0.02731f
C13274 VPWR.n1709 VGND 0.02047f
C13275 VPWR.n1710 VGND 0.02084f
C13276 VPWR.n1711 VGND 0.01313f
C13277 VPWR.n1713 VGND 0.01347f
C13278 VPWR.n1714 VGND 0.01763f
C13279 VPWR.n1715 VGND 0.13004f
C13280 VPWR.n1716 VGND 0.02213f
C13281 VPWR.n1717 VGND 0.02429f
C13282 VPWR.n1718 VGND 0.02304f
C13283 VPWR.n1719 VGND 0.02731f
C13284 VPWR.n1721 VGND 0.02047f
C13285 VPWR.n1722 VGND 0.02084f
C13286 VPWR.n1723 VGND 0.01313f
C13287 VPWR.n1725 VGND 0.01347f
C13288 VPWR.n1726 VGND 0.01763f
C13289 VPWR.n1727 VGND 0.1565f
C13290 VPWR.n1728 VGND 0.01879f
C13291 VPWR.n1729 VGND 0.01313f
C13292 VPWR.n1730 VGND 0.02047f
C13293 VPWR.n1731 VGND 0.02084f
C13294 VPWR.n1733 VGND 0.02304f
C13295 VPWR.n1734 VGND 0.02731f
C13296 VPWR.n1735 VGND 0.02542f
C13297 VPWR.n1737 VGND 0.01268f
C13298 VPWR.n1739 VGND 0.08003f
C13299 VPWR.t848 VGND 0.06817f
C13300 VPWR.t727 VGND 0.05805f
C13301 VPWR.t856 VGND 0.08842f
C13302 VPWR.n1740 VGND 0.08003f
C13303 VPWR.n1742 VGND 0.01268f
C13304 VPWR.n1744 VGND 0.04023f
C13305 VPWR.n1745 VGND 0.0225f
C13306 VPWR.t599 VGND 0.01981f
C13307 VPWR.n1747 VGND 0.04233f
C13308 VPWR.t1417 VGND 0.02189f
C13309 VPWR.n1748 VGND 0.0347f
C13310 VPWR.t869 VGND 0.05805f
C13311 VPWR.t1416 VGND 0.06817f
C13312 VPWR.t907 VGND 0.05805f
C13313 VPWR.t648 VGND 0.08842f
C13314 VPWR.n1749 VGND 0.08003f
C13315 VPWR.n1751 VGND 0.01329f
C13316 VPWR.n1752 VGND 0.10289f
C13317 VPWR.n1753 VGND -0.0138f
C13318 VPWR.n1754 VGND 0.06176f
C13319 VPWR.n1755 VGND 0.06176f
C13320 VPWR.n1756 VGND -0.0138f
C13321 VPWR.n1757 VGND 0.10289f
C13322 VPWR.n1758 VGND 0.01329f
C13323 VPWR.n1760 VGND 0.08003f
C13324 VPWR.t178 VGND 0.06817f
C13325 VPWR.t851 VGND 0.05805f
C13326 VPWR.t775 VGND 0.08842f
C13327 VPWR.n1761 VGND 0.08003f
C13328 VPWR.n1763 VGND 0.01329f
C13329 VPWR.n1764 VGND 0.10289f
C13330 VPWR.n1765 VGND 0.04023f
C13331 VPWR.n1766 VGND 0.04856f
C13332 VPWR.n1767 VGND 0.06785f
C13333 VPWR.n1768 VGND 0.02048f
C13334 VPWR.n1769 VGND 0.01403f
C13335 VPWR.n1770 VGND 0.04617f
C13336 VPWR.n1771 VGND 0.07207f
C13337 VPWR.n1772 VGND 0.06785f
C13338 VPWR.n1773 VGND 0.02048f
C13339 VPWR.n1774 VGND 0.01403f
C13340 VPWR.n1775 VGND 0.04617f
C13341 VPWR.n1776 VGND 0.07207f
C13342 VPWR.n1777 VGND 0.02048f
C13343 VPWR.n1778 VGND 0.01403f
C13344 VPWR.n1779 VGND 0.04616f
C13345 VPWR.n1780 VGND 0.038f
C13346 VPWR.n1781 VGND 0.02048f
C13347 VPWR.n1782 VGND 0.01403f
C13348 VPWR.n1783 VGND 0.04617f
C13349 VPWR.n1784 VGND 0.07207f
C13350 VPWR.n1785 VGND 0.06785f
C13351 VPWR.n1786 VGND 0.04856f
C13352 VPWR.n1787 VGND 0.04023f
C13353 VPWR.n1788 VGND 0.10289f
C13354 VPWR.n1789 VGND 0.01329f
C13355 VPWR.n1791 VGND 0.08003f
C13356 VPWR.t756 VGND 0.08842f
C13357 VPWR.t739 VGND 0.05805f
C13358 VPWR.t864 VGND 0.0986f
C13359 VPWR.n1792 VGND 0.05634f
C13360 VPWR.n1793 VGND 0.01329f
C13361 VPWR.n1794 VGND 0.10289f
C13362 VPWR.n1795 VGND 0.12172f
C13363 VPWR.n1796 VGND 0.75117f
C13364 VPWR.n1797 VGND 0.06176f
C13365 VPWR.n1798 VGND 0.06176f
C13366 VPWR.n1799 VGND 0.06176f
C13367 VPWR.n1800 VGND 0.06176f
C13368 VPWR.n1801 VGND 0.06176f
C13369 VPWR.n1802 VGND 0.06176f
C13370 VPWR.n1803 VGND 0.06176f
C13371 VPWR.n1804 VGND 0.06176f
C13372 VPWR.n1805 VGND 0.06176f
C13373 VPWR.n1806 VGND 0.06176f
C13374 VPWR.n1807 VGND 0.06176f
C13375 VPWR.n1808 VGND 0.06176f
C13376 VPWR.n1809 VGND 0.06176f
C13377 VPWR.n1810 VGND 0.06176f
C13378 VPWR.n1811 VGND 0.06176f
C13379 VPWR.n1812 VGND 0.14325f
C13380 VPWR.n1813 VGND 0.75117f
C13381 VPWR.n1814 VGND 0.75117f
C13382 VPWR.n1815 VGND 0.14325f
C13383 VPWR.n1816 VGND 0.10289f
C13384 VPWR.n1817 VGND 0.01329f
C13385 VPWR.n1818 VGND 0.05634f
C13386 VPWR.t901 VGND 0.0986f
C13387 VPWR.t26 VGND 0.05805f
C13388 VPWR.t196 VGND 0.08842f
C13389 VPWR.n1819 VGND 0.08003f
C13390 VPWR.n1821 VGND 0.01329f
C13391 VPWR.n1822 VGND 0.10289f
C13392 VPWR.n1823 VGND 0.06176f
C13393 VPWR.n1824 VGND 0.06176f
C13394 VPWR.n1825 VGND 0.10289f
C13395 VPWR.n1826 VGND 0.01329f
C13396 VPWR.n1828 VGND 0.08003f
C13397 VPWR.t1428 VGND 0.06817f
C13398 VPWR.t1327 VGND 0.05805f
C13399 VPWR.t288 VGND 0.08842f
C13400 VPWR.n1829 VGND 0.08003f
C13401 VPWR.n1831 VGND 0.01329f
C13402 VPWR.n1832 VGND 0.10289f
C13403 VPWR.n1833 VGND 0.06176f
C13404 VPWR.n1834 VGND 0.06176f
C13405 VPWR.n1835 VGND 0.10289f
C13406 VPWR.n1836 VGND 0.01329f
C13407 VPWR.n1838 VGND 0.08003f
C13408 VPWR.t970 VGND 0.06817f
C13409 VPWR.t1922 VGND 0.05805f
C13410 VPWR.t1745 VGND 0.08842f
C13411 VPWR.n1839 VGND 0.08003f
C13412 VPWR.n1841 VGND 0.01329f
C13413 VPWR.n1842 VGND 0.10289f
C13414 VPWR.n1843 VGND 0.06176f
C13415 VPWR.n1844 VGND 0.06176f
C13416 VPWR.n1845 VGND 0.10289f
C13417 VPWR.n1846 VGND 0.01329f
C13418 VPWR.n1848 VGND 0.08003f
C13419 VPWR.t409 VGND 0.06817f
C13420 VPWR.t1331 VGND 0.05805f
C13421 VPWR.t316 VGND 0.08842f
C13422 VPWR.n1849 VGND 0.08003f
C13423 VPWR.n1851 VGND 0.01329f
C13424 VPWR.n1852 VGND 0.10289f
C13425 VPWR.n1853 VGND 0.06176f
C13426 VPWR.n1854 VGND 0.06176f
C13427 VPWR.n1855 VGND 0.10289f
C13428 VPWR.n1856 VGND 0.01329f
C13429 VPWR.n1858 VGND 0.08003f
C13430 VPWR.t252 VGND 0.06817f
C13431 VPWR.t28 VGND 0.05805f
C13432 VPWR.t1865 VGND 0.08842f
C13433 VPWR.n1859 VGND 0.08003f
C13434 VPWR.n1861 VGND 0.01329f
C13435 VPWR.n1862 VGND 0.10289f
C13436 VPWR.n1863 VGND 0.06176f
C13437 VPWR.n1864 VGND 0.06176f
C13438 VPWR.n1865 VGND 0.10289f
C13439 VPWR.n1866 VGND 0.01329f
C13440 VPWR.n1868 VGND 0.08003f
C13441 VPWR.t1263 VGND 0.06817f
C13442 VPWR.t1330 VGND 0.05805f
C13443 VPWR.t109 VGND 0.08842f
C13444 VPWR.n1869 VGND 0.08003f
C13445 VPWR.n1871 VGND 0.01329f
C13446 VPWR.n1872 VGND 0.10289f
C13447 VPWR.n1873 VGND 0.06176f
C13448 VPWR.n1874 VGND 0.06176f
C13449 VPWR.n1875 VGND 0.10289f
C13450 VPWR.n1876 VGND 0.01329f
C13451 VPWR.n1878 VGND 0.08003f
C13452 VPWR.t1066 VGND 0.06817f
C13453 VPWR.t1924 VGND 0.05805f
C13454 VPWR.t1159 VGND 0.08842f
C13455 VPWR.n1879 VGND 0.08003f
C13456 VPWR.n1881 VGND 0.01329f
C13457 VPWR.n1882 VGND 0.10289f
C13458 VPWR.n1883 VGND 0.06176f
C13459 VPWR.n1884 VGND 0.06176f
C13460 VPWR.n1885 VGND 0.10289f
C13461 VPWR.n1886 VGND 0.01329f
C13462 VPWR.n1888 VGND 0.08003f
C13463 VPWR.t1550 VGND 0.06817f
C13464 VPWR.t25 VGND 0.05805f
C13465 VPWR.t16 VGND 0.08842f
C13466 VPWR.n1889 VGND 0.08003f
C13467 VPWR.n1891 VGND 0.01329f
C13468 VPWR.n1892 VGND 0.10289f
C13469 VPWR.n1893 VGND 0.06176f
C13470 VPWR.n1894 VGND 0.74646f
C13471 VPWR.n1895 VGND 0.14325f
C13472 VPWR.n1896 VGND 0.06176f
C13473 VPWR.n1897 VGND 0.06176f
C13474 VPWR.n1898 VGND 0.06176f
C13475 VPWR.n1899 VGND 0.06176f
C13476 VPWR.n1900 VGND 0.06176f
C13477 VPWR.n1901 VGND 0.06176f
C13478 VPWR.n1902 VGND 0.06176f
C13479 VPWR.n1903 VGND 0.06176f
C13480 VPWR.n1904 VGND 0.06176f
C13481 VPWR.n1905 VGND 0.06176f
C13482 VPWR.n1906 VGND 0.06176f
C13483 VPWR.n1907 VGND 0.06176f
C13484 VPWR.n1908 VGND 0.06176f
C13485 VPWR.n1909 VGND 0.06176f
C13486 VPWR.n1910 VGND 0.06176f
C13487 VPWR.n1911 VGND 0.74646f
C13488 VPWR.n1912 VGND 0.74646f
C13489 VPWR.n1913 VGND 0.06176f
C13490 VPWR.n1914 VGND 0.10289f
C13491 VPWR.n1915 VGND 0.01329f
C13492 VPWR.n1917 VGND 0.08003f
C13493 VPWR.t310 VGND 0.08842f
C13494 VPWR.t997 VGND 0.05805f
C13495 VPWR.t1706 VGND 0.06817f
C13496 VPWR.t331 VGND 0.05805f
C13497 VPWR.t1609 VGND 0.08842f
C13498 VPWR.n1918 VGND 0.08003f
C13499 VPWR.n1920 VGND 0.01329f
C13500 VPWR.n1921 VGND 0.10289f
C13501 VPWR.n1922 VGND 0.06176f
C13502 VPWR.n1923 VGND 0.06176f
C13503 VPWR.n1924 VGND 0.10289f
C13504 VPWR.n1925 VGND 0.01329f
C13505 VPWR.n1927 VGND 0.08003f
C13506 VPWR.t1177 VGND 0.08842f
C13507 VPWR.t330 VGND 0.05805f
C13508 VPWR.t1056 VGND 0.06817f
C13509 VPWR.t1001 VGND 0.05805f
C13510 VPWR.t1060 VGND 0.08842f
C13511 VPWR.n1928 VGND 0.08003f
C13512 VPWR.n1930 VGND 0.01329f
C13513 VPWR.n1931 VGND 0.10289f
C13514 VPWR.n1932 VGND 0.06176f
C13515 VPWR.n1933 VGND 0.06176f
C13516 VPWR.n1934 VGND 0.10289f
C13517 VPWR.n1935 VGND 0.01329f
C13518 VPWR.n1937 VGND 0.08003f
C13519 VPWR.t1522 VGND 0.08842f
C13520 VPWR.t1904 VGND 0.05805f
C13521 VPWR.t1279 VGND 0.06817f
C13522 VPWR.t1903 VGND 0.05805f
C13523 VPWR.t1273 VGND 0.08842f
C13524 VPWR.n1938 VGND 0.08003f
C13525 VPWR.n1940 VGND 0.01329f
C13526 VPWR.n1941 VGND 0.10289f
C13527 VPWR.n1942 VGND 0.06176f
C13528 VPWR.n1943 VGND 0.06176f
C13529 VPWR.n1944 VGND 0.10289f
C13530 VPWR.n1945 VGND 0.01329f
C13531 VPWR.n1947 VGND 0.08003f
C13532 VPWR.t232 VGND 0.08842f
C13533 VPWR.t1000 VGND 0.05805f
C13534 VPWR.t533 VGND 0.06817f
C13535 VPWR.t999 VGND 0.05805f
C13536 VPWR.t240 VGND 0.08842f
C13537 VPWR.n1948 VGND 0.08003f
C13538 VPWR.n1950 VGND 0.01329f
C13539 VPWR.n1951 VGND 0.10289f
C13540 VPWR.n1952 VGND 0.06176f
C13541 VPWR.n1953 VGND 0.06176f
C13542 VPWR.n1954 VGND 0.10289f
C13543 VPWR.n1955 VGND 0.01329f
C13544 VPWR.n1957 VGND 0.08003f
C13545 VPWR.t132 VGND 0.08842f
C13546 VPWR.t1905 VGND 0.05805f
C13547 VPWR.t376 VGND 0.06817f
C13548 VPWR.t329 VGND 0.05805f
C13549 VPWR.t358 VGND 0.08842f
C13550 VPWR.n1958 VGND 0.08003f
C13551 VPWR.n1960 VGND 0.01329f
C13552 VPWR.n1961 VGND 0.10289f
C13553 VPWR.n1962 VGND 0.06176f
C13554 VPWR.n1963 VGND 0.06176f
C13555 VPWR.n1964 VGND 0.10289f
C13556 VPWR.n1965 VGND 0.01329f
C13557 VPWR.n1967 VGND 0.08003f
C13558 VPWR.t1120 VGND 0.08842f
C13559 VPWR.t328 VGND 0.05805f
C13560 VPWR.t1841 VGND 0.06817f
C13561 VPWR.t334 VGND 0.05805f
C13562 VPWR.t1538 VGND 0.08842f
C13563 VPWR.n1968 VGND 0.08003f
C13564 VPWR.n1970 VGND 0.01329f
C13565 VPWR.n1971 VGND 0.10289f
C13566 VPWR.n1972 VGND 0.06176f
C13567 VPWR.n1973 VGND 0.06176f
C13568 VPWR.n1974 VGND 0.10289f
C13569 VPWR.n1975 VGND 0.01329f
C13570 VPWR.n1977 VGND 0.08003f
C13571 VPWR.t51 VGND 0.08842f
C13572 VPWR.t333 VGND 0.05805f
C13573 VPWR.t972 VGND 0.06817f
C13574 VPWR.t332 VGND 0.05805f
C13575 VPWR.t487 VGND 0.08842f
C13576 VPWR.n1978 VGND 0.08003f
C13577 VPWR.n1980 VGND 0.01329f
C13578 VPWR.n1981 VGND 0.10289f
C13579 VPWR.n1982 VGND 0.06176f
C13580 VPWR.n1983 VGND 0.06176f
C13581 VPWR.n1984 VGND 0.10289f
C13582 VPWR.n1985 VGND 0.01329f
C13583 VPWR.n1987 VGND 0.08003f
C13584 VPWR.t208 VGND 0.08842f
C13585 VPWR.t998 VGND 0.05805f
C13586 VPWR.t609 VGND 0.0986f
C13587 VPWR.n1988 VGND 0.05634f
C13588 VPWR.n1989 VGND 0.01329f
C13589 VPWR.n1990 VGND 0.10289f
C13590 VPWR.n1991 VGND 0.14325f
C13591 VPWR.n1992 VGND 0.75117f
C13592 VPWR.n1993 VGND 0.06176f
C13593 VPWR.n1994 VGND 0.06176f
C13594 VPWR.n1995 VGND 0.06176f
C13595 VPWR.n1996 VGND 0.06176f
C13596 VPWR.n1997 VGND 0.06176f
C13597 VPWR.n1998 VGND 0.06176f
C13598 VPWR.n1999 VGND 0.06176f
C13599 VPWR.n2000 VGND 0.06176f
C13600 VPWR.n2001 VGND 0.06176f
C13601 VPWR.n2002 VGND 0.06176f
C13602 VPWR.n2003 VGND 0.06176f
C13603 VPWR.n2004 VGND 0.06176f
C13604 VPWR.n2005 VGND 0.06176f
C13605 VPWR.n2006 VGND 0.06176f
C13606 VPWR.n2007 VGND 0.06176f
C13607 VPWR.n2008 VGND 0.14325f
C13608 VPWR.n2009 VGND 0.75117f
C13609 VPWR.n2010 VGND 0.75117f
C13610 VPWR.n2011 VGND 0.14325f
C13611 VPWR.n2012 VGND 0.10289f
C13612 VPWR.n2013 VGND 0.01329f
C13613 VPWR.n2014 VGND 0.05634f
C13614 VPWR.t681 VGND 0.0986f
C13615 VPWR.t1246 VGND 0.05805f
C13616 VPWR.t6 VGND 0.08842f
C13617 VPWR.n2015 VGND 0.08003f
C13618 VPWR.n2017 VGND 0.01329f
C13619 VPWR.n2018 VGND 0.10289f
C13620 VPWR.n2019 VGND 0.06176f
C13621 VPWR.n2020 VGND 0.06176f
C13622 VPWR.n2021 VGND 0.10289f
C13623 VPWR.n2022 VGND 0.01329f
C13624 VPWR.n2024 VGND 0.08003f
C13625 VPWR.t1084 VGND 0.06817f
C13626 VPWR.t1008 VGND 0.05805f
C13627 VPWR.t39 VGND 0.08842f
C13628 VPWR.n2025 VGND 0.08003f
C13629 VPWR.n2027 VGND 0.01329f
C13630 VPWR.n2028 VGND 0.10289f
C13631 VPWR.n2029 VGND 0.06176f
C13632 VPWR.n2030 VGND 0.06176f
C13633 VPWR.n2031 VGND 0.10289f
C13634 VPWR.n2032 VGND 0.01329f
C13635 VPWR.n2034 VGND 0.08003f
C13636 VPWR.t1534 VGND 0.06817f
C13637 VPWR.t1003 VGND 0.05805f
C13638 VPWR.t1848 VGND 0.08842f
C13639 VPWR.n2035 VGND 0.08003f
C13640 VPWR.n2037 VGND 0.01329f
C13641 VPWR.n2038 VGND 0.10289f
C13642 VPWR.n2039 VGND 0.06176f
C13643 VPWR.n2040 VGND 0.06176f
C13644 VPWR.n2041 VGND 0.10289f
C13645 VPWR.n2042 VGND 0.01329f
C13646 VPWR.n2044 VGND 0.08003f
C13647 VPWR.t354 VGND 0.06817f
C13648 VPWR.t1570 VGND 0.05805f
C13649 VPWR.t1221 VGND 0.08842f
C13650 VPWR.n2045 VGND 0.08003f
C13651 VPWR.n2047 VGND 0.01329f
C13652 VPWR.n2048 VGND 0.10289f
C13653 VPWR.n2049 VGND 0.06176f
C13654 VPWR.n2050 VGND 0.06176f
C13655 VPWR.n2051 VGND 0.10289f
C13656 VPWR.n2052 VGND 0.01329f
C13657 VPWR.n2054 VGND 0.08003f
C13658 VPWR.t501 VGND 0.06817f
C13659 VPWR.t1248 VGND 0.05805f
C13660 VPWR.t226 VGND 0.08842f
C13661 VPWR.n2055 VGND 0.08003f
C13662 VPWR.n2057 VGND 0.01329f
C13663 VPWR.n2058 VGND 0.10289f
C13664 VPWR.n2059 VGND 0.06176f
C13665 VPWR.n2060 VGND 0.06176f
C13666 VPWR.n2061 VGND 0.10289f
C13667 VPWR.n2062 VGND 0.01329f
C13668 VPWR.n2064 VGND 0.08003f
C13669 VPWR.t1345 VGND 0.06817f
C13670 VPWR.t1011 VGND 0.05805f
C13671 VPWR.t1306 VGND 0.08842f
C13672 VPWR.n2065 VGND 0.08003f
C13673 VPWR.n2067 VGND 0.01329f
C13674 VPWR.n2068 VGND 0.10289f
C13675 VPWR.n2069 VGND 0.06176f
C13676 VPWR.n2070 VGND 0.06176f
C13677 VPWR.n2071 VGND 0.10289f
C13678 VPWR.n2072 VGND 0.01329f
C13679 VPWR.n2074 VGND 0.08003f
C13680 VPWR.t1414 VGND 0.06817f
C13681 VPWR.t1005 VGND 0.05805f
C13682 VPWR.t1185 VGND 0.08842f
C13683 VPWR.n2075 VGND 0.08003f
C13684 VPWR.n2077 VGND 0.01329f
C13685 VPWR.n2078 VGND 0.10289f
C13686 VPWR.n2079 VGND 0.06176f
C13687 VPWR.n2080 VGND 0.06176f
C13688 VPWR.n2081 VGND 0.10289f
C13689 VPWR.n2082 VGND 0.01329f
C13690 VPWR.n2084 VGND 0.08003f
C13691 VPWR.t512 VGND 0.06817f
C13692 VPWR.t1571 VGND 0.05805f
C13693 VPWR.t459 VGND 0.08842f
C13694 VPWR.n2085 VGND 0.08003f
C13695 VPWR.n2087 VGND 0.01329f
C13696 VPWR.n2088 VGND 0.10289f
C13697 VPWR.n2089 VGND 0.06176f
C13698 VPWR.n2090 VGND 0.74646f
C13699 VPWR.n2091 VGND 0.14325f
C13700 VPWR.n2092 VGND 0.06176f
C13701 VPWR.n2093 VGND 0.06176f
C13702 VPWR.n2094 VGND 0.06176f
C13703 VPWR.n2095 VGND 0.06176f
C13704 VPWR.n2096 VGND 0.06176f
C13705 VPWR.n2097 VGND 0.06176f
C13706 VPWR.n2098 VGND 0.06176f
C13707 VPWR.n2099 VGND 0.06176f
C13708 VPWR.n2100 VGND 0.06176f
C13709 VPWR.n2101 VGND 0.06176f
C13710 VPWR.n2102 VGND 0.06176f
C13711 VPWR.n2103 VGND 0.06176f
C13712 VPWR.n2104 VGND 0.06176f
C13713 VPWR.n2105 VGND 0.06176f
C13714 VPWR.n2106 VGND 0.06176f
C13715 VPWR.n2107 VGND 0.74646f
C13716 VPWR.n2108 VGND 0.74646f
C13717 VPWR.n2109 VGND 0.06176f
C13718 VPWR.n2110 VGND 0.10289f
C13719 VPWR.n2111 VGND 0.01329f
C13720 VPWR.n2113 VGND 0.08003f
C13721 VPWR.t308 VGND 0.08842f
C13722 VPWR.t1090 VGND 0.05805f
C13723 VPWR.t1613 VGND 0.06817f
C13724 VPWR.t1517 VGND 0.05805f
C13725 VPWR.t1607 VGND 0.08842f
C13726 VPWR.n2114 VGND 0.08003f
C13727 VPWR.n2116 VGND 0.01329f
C13728 VPWR.n2117 VGND 0.10289f
C13729 VPWR.n2118 VGND 0.06176f
C13730 VPWR.n2119 VGND 0.06176f
C13731 VPWR.n2120 VGND 0.10289f
C13732 VPWR.n2121 VGND 0.01329f
C13733 VPWR.n2123 VGND 0.08003f
C13734 VPWR.t1179 VGND 0.08842f
C13735 VPWR.t505 VGND 0.05805f
C13736 VPWR.t1052 VGND 0.06817f
C13737 VPWR.t1088 VGND 0.05805f
C13738 VPWR.t1027 VGND 0.08842f
C13739 VPWR.n2124 VGND 0.08003f
C13740 VPWR.n2126 VGND 0.01329f
C13741 VPWR.n2127 VGND 0.10289f
C13742 VPWR.n2128 VGND 0.06176f
C13743 VPWR.n2129 VGND 0.06176f
C13744 VPWR.n2130 VGND 0.10289f
C13745 VPWR.n2131 VGND 0.01329f
C13746 VPWR.n2133 VGND 0.08003f
C13747 VPWR.t1520 VGND 0.08842f
C13748 VPWR.t97 VGND 0.05805f
C13749 VPWR.t1277 VGND 0.06817f
C13750 VPWR.t96 VGND 0.05805f
C13751 VPWR.t1271 VGND 0.08842f
C13752 VPWR.n2134 VGND 0.08003f
C13753 VPWR.n2136 VGND 0.01329f
C13754 VPWR.n2137 VGND 0.10289f
C13755 VPWR.n2138 VGND 0.06176f
C13756 VPWR.n2139 VGND 0.06176f
C13757 VPWR.n2140 VGND 0.10289f
C13758 VPWR.n2141 VGND 0.01329f
C13759 VPWR.n2143 VGND 0.08003f
C13760 VPWR.t230 VGND 0.08842f
C13761 VPWR.t1087 VGND 0.05805f
C13762 VPWR.t531 VGND 0.06817f
C13763 VPWR.t1086 VGND 0.05805f
C13764 VPWR.t1405 VGND 0.08842f
C13765 VPWR.n2144 VGND 0.08003f
C13766 VPWR.n2146 VGND 0.01329f
C13767 VPWR.n2147 VGND 0.10289f
C13768 VPWR.n2148 VGND 0.06176f
C13769 VPWR.n2149 VGND 0.06176f
C13770 VPWR.n2150 VGND 0.10289f
C13771 VPWR.n2151 VGND 0.01329f
C13772 VPWR.n2153 VGND 0.08003f
C13773 VPWR.t130 VGND 0.08842f
C13774 VPWR.t98 VGND 0.05805f
C13775 VPWR.t362 VGND 0.06817f
C13776 VPWR.t504 VGND 0.05805f
C13777 VPWR.t356 VGND 0.08842f
C13778 VPWR.n2154 VGND 0.08003f
C13779 VPWR.n2156 VGND 0.01329f
C13780 VPWR.n2157 VGND 0.10289f
C13781 VPWR.n2158 VGND 0.06176f
C13782 VPWR.n2159 VGND 0.06176f
C13783 VPWR.n2160 VGND 0.10289f
C13784 VPWR.n2161 VGND 0.01329f
C13785 VPWR.n2163 VGND 0.08003f
C13786 VPWR.t1118 VGND 0.08842f
C13787 VPWR.t503 VGND 0.05805f
C13788 VPWR.t1839 VGND 0.06817f
C13789 VPWR.t95 VGND 0.05805f
C13790 VPWR.t1536 VGND 0.08842f
C13791 VPWR.n2164 VGND 0.08003f
C13792 VPWR.n2166 VGND 0.01329f
C13793 VPWR.n2167 VGND 0.10289f
C13794 VPWR.n2168 VGND 0.06176f
C13795 VPWR.n2169 VGND 0.06176f
C13796 VPWR.n2170 VGND 0.10289f
C13797 VPWR.n2171 VGND 0.01329f
C13798 VPWR.n2173 VGND 0.08003f
C13799 VPWR.t49 VGND 0.08842f
C13800 VPWR.t1519 VGND 0.05805f
C13801 VPWR.t491 VGND 0.06817f
C13802 VPWR.t1518 VGND 0.05805f
C13803 VPWR.t485 VGND 0.08842f
C13804 VPWR.n2174 VGND 0.08003f
C13805 VPWR.n2176 VGND 0.01329f
C13806 VPWR.n2177 VGND 0.10289f
C13807 VPWR.n2178 VGND 0.06176f
C13808 VPWR.n2179 VGND 0.06176f
C13809 VPWR.n2180 VGND 0.10289f
C13810 VPWR.n2181 VGND 0.01329f
C13811 VPWR.n2183 VGND 0.08003f
C13812 VPWR.t206 VGND 0.08842f
C13813 VPWR.t1091 VGND 0.05805f
C13814 VPWR.t614 VGND 0.0986f
C13815 VPWR.n2184 VGND 0.05634f
C13816 VPWR.n2185 VGND 0.01329f
C13817 VPWR.n2186 VGND 0.10289f
C13818 VPWR.n2187 VGND 0.14325f
C13819 VPWR.n2188 VGND 0.75117f
C13820 VPWR.n2189 VGND 0.06176f
C13821 VPWR.n2190 VGND 0.06176f
C13822 VPWR.n2191 VGND 0.06176f
C13823 VPWR.n2192 VGND 0.06176f
C13824 VPWR.n2193 VGND 0.06176f
C13825 VPWR.n2194 VGND 0.06176f
C13826 VPWR.n2195 VGND 0.06176f
C13827 VPWR.n2196 VGND 0.06176f
C13828 VPWR.n2197 VGND 0.06176f
C13829 VPWR.n2198 VGND 0.06176f
C13830 VPWR.n2199 VGND 0.06176f
C13831 VPWR.n2200 VGND 0.06176f
C13832 VPWR.n2201 VGND 0.06176f
C13833 VPWR.n2202 VGND 0.06176f
C13834 VPWR.n2203 VGND 0.06176f
C13835 VPWR.n2204 VGND 0.14325f
C13836 VPWR.n2205 VGND 0.75117f
C13837 VPWR.n2206 VGND 0.75117f
C13838 VPWR.n2207 VGND 0.14325f
C13839 VPWR.n2208 VGND 0.10289f
C13840 VPWR.n2209 VGND 0.01329f
C13841 VPWR.n2210 VGND 0.05634f
C13842 VPWR.t780 VGND 0.0986f
C13843 VPWR.t1684 VGND 0.05805f
C13844 VPWR.t1635 VGND 0.08842f
C13845 VPWR.n2211 VGND 0.08003f
C13846 VPWR.n2213 VGND 0.01329f
C13847 VPWR.n2214 VGND 0.10289f
C13848 VPWR.n2215 VGND 0.06176f
C13849 VPWR.n2216 VGND 0.06176f
C13850 VPWR.n2217 VGND 0.10289f
C13851 VPWR.n2218 VGND 0.01329f
C13852 VPWR.n2220 VGND 0.08003f
C13853 VPWR.t1202 VGND 0.06817f
C13854 VPWR.t1678 VGND 0.05805f
C13855 VPWR.t166 VGND 0.08842f
C13856 VPWR.n2221 VGND 0.08003f
C13857 VPWR.n2223 VGND 0.01329f
C13858 VPWR.n2224 VGND 0.10289f
C13859 VPWR.n2225 VGND 0.06176f
C13860 VPWR.n2226 VGND 0.06176f
C13861 VPWR.n2227 VGND 0.10289f
C13862 VPWR.n2228 VGND 0.01329f
C13863 VPWR.n2230 VGND 0.08003f
C13864 VPWR.t1895 VGND 0.06817f
C13865 VPWR.t1436 VGND 0.05805f
C13866 VPWR.t475 VGND 0.08842f
C13867 VPWR.n2231 VGND 0.08003f
C13868 VPWR.n2233 VGND 0.01329f
C13869 VPWR.n2234 VGND 0.10289f
C13870 VPWR.n2235 VGND 0.06176f
C13871 VPWR.n2236 VGND 0.06176f
C13872 VPWR.n2237 VGND 0.10289f
C13873 VPWR.n2238 VGND 0.01329f
C13874 VPWR.n2240 VGND 0.08003f
C13875 VPWR.t443 VGND 0.06817f
C13876 VPWR.t1682 VGND 0.05805f
C13877 VPWR.t522 VGND 0.08842f
C13878 VPWR.n2241 VGND 0.08003f
C13879 VPWR.n2243 VGND 0.01329f
C13880 VPWR.n2244 VGND 0.10289f
C13881 VPWR.n2245 VGND 0.06176f
C13882 VPWR.n2246 VGND 0.06176f
C13883 VPWR.n2247 VGND 0.10289f
C13884 VPWR.n2248 VGND 0.01329f
C13885 VPWR.n2250 VGND 0.08003f
C13886 VPWR.t1401 VGND 0.06817f
C13887 VPWR.t345 VGND 0.05805f
C13888 VPWR.t1697 VGND 0.08842f
C13889 VPWR.n2251 VGND 0.08003f
C13890 VPWR.n2253 VGND 0.01329f
C13891 VPWR.n2254 VGND 0.10289f
C13892 VPWR.n2255 VGND 0.06176f
C13893 VPWR.n2256 VGND 0.06176f
C13894 VPWR.n2257 VGND 0.10289f
C13895 VPWR.n2258 VGND 0.01329f
C13896 VPWR.n2260 VGND 0.08003f
C13897 VPWR.t1504 VGND 0.06817f
C13898 VPWR.t1681 VGND 0.05805f
C13899 VPWR.t1554 VGND 0.08842f
C13900 VPWR.n2261 VGND 0.08003f
C13901 VPWR.n2263 VGND 0.01329f
C13902 VPWR.n2264 VGND 0.10289f
C13903 VPWR.n2265 VGND 0.06176f
C13904 VPWR.n2266 VGND 0.06176f
C13905 VPWR.n2267 VGND 0.10289f
C13906 VPWR.n2268 VGND 0.01329f
C13907 VPWR.n2270 VGND 0.08003f
C13908 VPWR.t1023 VGND 0.06817f
C13909 VPWR.t1438 VGND 0.05805f
C13910 VPWR.t1143 VGND 0.08842f
C13911 VPWR.n2271 VGND 0.08003f
C13912 VPWR.n2273 VGND 0.01329f
C13913 VPWR.n2274 VGND 0.10289f
C13914 VPWR.n2275 VGND 0.06176f
C13915 VPWR.n2276 VGND 0.06176f
C13916 VPWR.n2277 VGND 0.10289f
C13917 VPWR.n2278 VGND 0.01329f
C13918 VPWR.n2280 VGND 0.08003f
C13919 VPWR.t1655 VGND 0.06817f
C13920 VPWR.t1683 VGND 0.05805f
C13921 VPWR.t557 VGND 0.08842f
C13922 VPWR.n2281 VGND 0.08003f
C13923 VPWR.n2283 VGND 0.01329f
C13924 VPWR.n2284 VGND 0.10289f
C13925 VPWR.n2285 VGND 0.06176f
C13926 VPWR.n2286 VGND 0.74646f
C13927 VPWR.n2287 VGND 0.14325f
C13928 VPWR.n2288 VGND 0.06176f
C13929 VPWR.n2289 VGND 0.06176f
C13930 VPWR.n2290 VGND 0.06176f
C13931 VPWR.n2291 VGND 0.06176f
C13932 VPWR.n2292 VGND 0.06176f
C13933 VPWR.n2293 VGND 0.06176f
C13934 VPWR.n2294 VGND 0.06176f
C13935 VPWR.n2295 VGND 0.06176f
C13936 VPWR.n2296 VGND 0.06176f
C13937 VPWR.n2297 VGND 0.06176f
C13938 VPWR.n2298 VGND 0.06176f
C13939 VPWR.n2299 VGND 0.06176f
C13940 VPWR.n2300 VGND 0.06176f
C13941 VPWR.n2301 VGND 0.06176f
C13942 VPWR.n2302 VGND 0.06176f
C13943 VPWR.n2303 VGND 0.74646f
C13944 VPWR.n2304 VGND 0.74646f
C13945 VPWR.n2305 VGND 0.06176f
C13946 VPWR.n2306 VGND 0.10289f
C13947 VPWR.n2307 VGND 0.01329f
C13948 VPWR.n2309 VGND 0.08003f
C13949 VPWR.t85 VGND 0.08842f
C13950 VPWR.t1572 VGND 0.05805f
C13951 VPWR.t508 VGND 0.06817f
C13952 VPWR.t1855 VGND 0.05805f
C13953 VPWR.t128 VGND 0.08842f
C13954 VPWR.n2310 VGND 0.08003f
C13955 VPWR.n2312 VGND 0.01329f
C13956 VPWR.n2313 VGND 0.10289f
C13957 VPWR.n2314 VGND 0.06176f
C13958 VPWR.n2315 VGND 0.06176f
C13959 VPWR.n2316 VGND 0.10289f
C13960 VPWR.n2317 VGND 0.01329f
C13961 VPWR.n2319 VGND 0.08003f
C13962 VPWR.t1189 VGND 0.08842f
C13963 VPWR.t1854 VGND 0.05805f
C13964 VPWR.t1412 VGND 0.06817f
C13965 VPWR.t1676 VGND 0.05805f
C13966 VPWR.t146 VGND 0.08842f
C13967 VPWR.n2320 VGND 0.08003f
C13968 VPWR.n2322 VGND 0.01329f
C13969 VPWR.n2323 VGND 0.10289f
C13970 VPWR.n2324 VGND 0.06176f
C13971 VPWR.n2325 VGND 0.06176f
C13972 VPWR.n2326 VGND 0.10289f
C13973 VPWR.n2327 VGND 0.01329f
C13974 VPWR.n2329 VGND 0.08003f
C13975 VPWR.t1579 VGND 0.08842f
C13976 VPWR.t1725 VGND 0.05805f
C13977 VPWR.t1341 VGND 0.06817f
C13978 VPWR.t1724 VGND 0.05805f
C13979 VPWR.t1289 VGND 0.08842f
C13980 VPWR.n2330 VGND 0.08003f
C13981 VPWR.n2332 VGND 0.01329f
C13982 VPWR.n2333 VGND 0.10289f
C13983 VPWR.n2334 VGND 0.06176f
C13984 VPWR.n2335 VGND 0.06176f
C13985 VPWR.n2336 VGND 0.10289f
C13986 VPWR.n2337 VGND 0.01329f
C13987 VPWR.n2339 VGND 0.08003f
C13988 VPWR.t220 VGND 0.08842f
C13989 VPWR.t1675 VGND 0.05805f
C13990 VPWR.t168 VGND 0.06817f
C13991 VPWR.t1574 VGND 0.05805f
C13992 VPWR.t1384 VGND 0.08842f
C13993 VPWR.n2340 VGND 0.08003f
C13994 VPWR.n2342 VGND 0.01329f
C13995 VPWR.n2343 VGND 0.10289f
C13996 VPWR.n2344 VGND 0.06176f
C13997 VPWR.n2345 VGND 0.06176f
C13998 VPWR.n2346 VGND 0.10289f
C13999 VPWR.n2347 VGND 0.01329f
C14000 VPWR.n2349 VGND 0.08003f
C14001 VPWR.t561 VGND 0.08842f
C14002 VPWR.t1726 VGND 0.05805f
C14003 VPWR.t352 VGND 0.06817f
C14004 VPWR.t1853 VGND 0.05805f
C14005 VPWR.t447 VGND 0.08842f
C14006 VPWR.n2350 VGND 0.08003f
C14007 VPWR.n2352 VGND 0.01329f
C14008 VPWR.n2353 VGND 0.10289f
C14009 VPWR.n2354 VGND 0.06176f
C14010 VPWR.n2355 VGND 0.06176f
C14011 VPWR.n2356 VGND 0.10289f
C14012 VPWR.n2357 VGND 0.01329f
C14013 VPWR.n2359 VGND 0.08003f
C14014 VPWR.t1735 VGND 0.08842f
C14015 VPWR.t1852 VGND 0.05805f
C14016 VPWR.t1886 VGND 0.06817f
C14017 VPWR.t1723 VGND 0.05805f
C14018 VPWR.t1899 VGND 0.08842f
C14019 VPWR.n2360 VGND 0.08003f
C14020 VPWR.n2362 VGND 0.01329f
C14021 VPWR.n2363 VGND 0.10289f
C14022 VPWR.n2364 VGND 0.06176f
C14023 VPWR.n2365 VGND 0.06176f
C14024 VPWR.n2366 VGND 0.10289f
C14025 VPWR.n2367 VGND 0.01329f
C14026 VPWR.n2369 VGND 0.08003f
C14027 VPWR.t182 VGND 0.08842f
C14028 VPWR.t1722 VGND 0.05805f
C14029 VPWR.t1082 VGND 0.06817f
C14030 VPWR.t1856 VGND 0.05805f
C14031 VPWR.t1206 VGND 0.08842f
C14032 VPWR.n2370 VGND 0.08003f
C14033 VPWR.n2372 VGND 0.01329f
C14034 VPWR.n2373 VGND 0.10289f
C14035 VPWR.n2374 VGND 0.06176f
C14036 VPWR.n2375 VGND 0.06176f
C14037 VPWR.n2376 VGND 0.10289f
C14038 VPWR.n2377 VGND 0.01329f
C14039 VPWR.n2379 VGND 0.08003f
C14040 VPWR.t4 VGND 0.08842f
C14041 VPWR.t1573 VGND 0.05805f
C14042 VPWR.t713 VGND 0.0986f
C14043 VPWR.n2380 VGND 0.05634f
C14044 VPWR.n2381 VGND 0.01329f
C14045 VPWR.n2382 VGND 0.10289f
C14046 VPWR.n2383 VGND 0.14325f
C14047 VPWR.n2384 VGND 0.75117f
C14048 VPWR.n2385 VGND 0.06176f
C14049 VPWR.n2386 VGND 0.06176f
C14050 VPWR.n2387 VGND 0.06176f
C14051 VPWR.n2388 VGND 0.06176f
C14052 VPWR.n2389 VGND 0.06176f
C14053 VPWR.n2390 VGND 0.06176f
C14054 VPWR.n2391 VGND 0.06176f
C14055 VPWR.n2392 VGND 0.06176f
C14056 VPWR.n2393 VGND 0.06176f
C14057 VPWR.n2394 VGND 0.06176f
C14058 VPWR.n2395 VGND 0.06176f
C14059 VPWR.n2396 VGND 0.06176f
C14060 VPWR.n2397 VGND 0.06176f
C14061 VPWR.n2398 VGND 0.06176f
C14062 VPWR.n2399 VGND 0.06176f
C14063 VPWR.n2400 VGND 0.14325f
C14064 VPWR.n2401 VGND 0.75117f
C14065 VPWR.n2402 VGND 0.75117f
C14066 VPWR.n2403 VGND 0.14325f
C14067 VPWR.n2404 VGND 0.10289f
C14068 VPWR.n2405 VGND 0.01329f
C14069 VPWR.n2406 VGND 0.05634f
C14070 VPWR.t880 VGND 0.0986f
C14071 VPWR.t1873 VGND 0.05805f
C14072 VPWR.t393 VGND 0.08842f
C14073 VPWR.n2407 VGND 0.08003f
C14074 VPWR.n2409 VGND 0.01329f
C14075 VPWR.n2410 VGND 0.10289f
C14076 VPWR.n2411 VGND 0.06176f
C14077 VPWR.n2412 VGND 0.06176f
C14078 VPWR.n2413 VGND 0.10289f
C14079 VPWR.n2414 VGND 0.01329f
C14080 VPWR.n2416 VGND 0.08003f
C14081 VPWR.t1432 VGND 0.06817f
C14082 VPWR.t101 VGND 0.05805f
C14083 VPWR.t292 VGND 0.08842f
C14084 VPWR.n2417 VGND 0.08003f
C14085 VPWR.n2419 VGND 0.01329f
C14086 VPWR.n2420 VGND 0.10289f
C14087 VPWR.n2421 VGND 0.06176f
C14088 VPWR.n2422 VGND 0.06176f
C14089 VPWR.n2423 VGND 0.10289f
C14090 VPWR.n2424 VGND 0.01329f
C14091 VPWR.n2426 VGND 0.08003f
C14092 VPWR.t495 VGND 0.06817f
C14093 VPWR.t1719 VGND 0.05805f
C14094 VPWR.t1751 VGND 0.08842f
C14095 VPWR.n2427 VGND 0.08003f
C14096 VPWR.n2429 VGND 0.01329f
C14097 VPWR.n2430 VGND 0.10289f
C14098 VPWR.n2431 VGND 0.06176f
C14099 VPWR.n2432 VGND 0.06176f
C14100 VPWR.n2433 VGND 0.10289f
C14101 VPWR.n2434 VGND 0.01329f
C14102 VPWR.n2436 VGND 0.08003f
C14103 VPWR.t413 VGND 0.06817f
C14104 VPWR.t1880 VGND 0.05805f
C14105 VPWR.t322 VGND 0.08842f
C14106 VPWR.n2437 VGND 0.08003f
C14107 VPWR.n2439 VGND 0.01329f
C14108 VPWR.n2440 VGND 0.10289f
C14109 VPWR.n2441 VGND 0.06176f
C14110 VPWR.n2442 VGND 0.06176f
C14111 VPWR.n2443 VGND 0.10289f
C14112 VPWR.n2444 VGND 0.01329f
C14113 VPWR.n2446 VGND 0.08003f
C14114 VPWR.t954 VGND 0.06817f
C14115 VPWR.t1875 VGND 0.05805f
C14116 VPWR.t1871 VGND 0.08842f
C14117 VPWR.n2447 VGND 0.08003f
C14118 VPWR.n2449 VGND 0.01329f
C14119 VPWR.n2450 VGND 0.10289f
C14120 VPWR.n2451 VGND 0.06176f
C14121 VPWR.n2452 VGND 0.06176f
C14122 VPWR.n2453 VGND 0.10289f
C14123 VPWR.n2454 VGND 0.01329f
C14124 VPWR.n2456 VGND 0.08003f
C14125 VPWR.t1267 VGND 0.06817f
C14126 VPWR.t1879 VGND 0.05805f
C14127 VPWR.t115 VGND 0.08842f
C14128 VPWR.n2457 VGND 0.08003f
C14129 VPWR.n2459 VGND 0.01329f
C14130 VPWR.n2460 VGND 0.10289f
C14131 VPWR.n2461 VGND 0.06176f
C14132 VPWR.n2462 VGND 0.06176f
C14133 VPWR.n2463 VGND 0.10289f
C14134 VPWR.n2464 VGND 0.01329f
C14135 VPWR.n2466 VGND 0.08003f
C14136 VPWR.t1072 VGND 0.06817f
C14137 VPWR.t1721 VGND 0.05805f
C14138 VPWR.t1155 VGND 0.08842f
C14139 VPWR.n2467 VGND 0.08003f
C14140 VPWR.n2469 VGND 0.01329f
C14141 VPWR.n2470 VGND 0.10289f
C14142 VPWR.n2471 VGND 0.06176f
C14143 VPWR.n2472 VGND 0.06176f
C14144 VPWR.n2473 VGND 0.10289f
C14145 VPWR.n2474 VGND 0.01329f
C14146 VPWR.n2476 VGND 0.08003f
C14147 VPWR.t1530 VGND 0.06817f
C14148 VPWR.t1881 VGND 0.05805f
C14149 VPWR.t985 VGND 0.08842f
C14150 VPWR.n2477 VGND 0.08003f
C14151 VPWR.n2479 VGND 0.01329f
C14152 VPWR.n2480 VGND 0.10289f
C14153 VPWR.n2481 VGND 0.06176f
C14154 VPWR.n2482 VGND 0.74646f
C14155 VPWR.n2483 VGND 0.14325f
C14156 VPWR.n2484 VGND 0.06176f
C14157 VPWR.n2485 VGND 0.06176f
C14158 VPWR.n2486 VGND 0.06176f
C14159 VPWR.n2487 VGND 0.06176f
C14160 VPWR.n2488 VGND 0.06176f
C14161 VPWR.n2489 VGND 0.06176f
C14162 VPWR.n2490 VGND 0.06176f
C14163 VPWR.n2491 VGND 0.06176f
C14164 VPWR.n2492 VGND 0.06176f
C14165 VPWR.n2493 VGND 0.06176f
C14166 VPWR.n2494 VGND 0.06176f
C14167 VPWR.n2495 VGND 0.06176f
C14168 VPWR.n2496 VGND 0.06176f
C14169 VPWR.n2497 VGND 0.06176f
C14170 VPWR.n2498 VGND 0.06176f
C14171 VPWR.n2499 VGND 0.74646f
C14172 VPWR.n2500 VGND 0.42248f
C14173 VPWR.n2501 VGND 0.06176f
C14174 VPWR.n2502 VGND 0.064f
C14175 VPWR.n2504 VGND 0.01268f
C14176 VPWR.n2506 VGND 0.08003f
C14177 VPWR.t762 VGND 0.08842f
C14178 VPWR.t729 VGND 0.05805f
C14179 VPWR.t853 VGND 0.06817f
C14180 VPWR.t859 VGND 0.05805f
C14181 VPWR.t874 VGND 0.08842f
C14182 VPWR.n2507 VGND 0.08003f
C14183 VPWR.n2509 VGND 0.01268f
C14184 VPWR.n2511 VGND 0.064f
C14185 VPWR.n2512 VGND 0.06176f
C14186 VPWR.n2513 VGND 0.06176f
C14187 VPWR.n2514 VGND 0.064f
C14188 VPWR.n2516 VGND 0.01268f
C14189 VPWR.n2518 VGND 0.08003f
C14190 VPWR.t639 VGND 0.08842f
C14191 VPWR.t899 VGND 0.05805f
C14192 VPWR.t633 VGND 0.06817f
C14193 VPWR.t623 VGND 0.05805f
C14194 VPWR.t750 VGND 0.08842f
C14195 VPWR.n2519 VGND 0.08003f
C14196 VPWR.n2521 VGND 0.01268f
C14197 VPWR.n2523 VGND 0.064f
C14198 VPWR.n2524 VGND 0.06176f
C14199 VPWR.n2525 VGND 0.06176f
C14200 VPWR.n2526 VGND 0.064f
C14201 VPWR.n2528 VGND 0.01268f
C14202 VPWR.n2530 VGND 0.08003f
C14203 VPWR.t759 VGND 0.08842f
C14204 VPWR.t767 VGND 0.05805f
C14205 VPWR.t896 VGND 0.06817f
C14206 VPWR.t791 VGND 0.05805f
C14207 VPWR.t915 VGND 0.08842f
C14208 VPWR.n2531 VGND 0.08003f
C14209 VPWR.n2533 VGND 0.01268f
C14210 VPWR.n2535 VGND 0.064f
C14211 VPWR.n2536 VGND 0.06176f
C14212 VPWR.n2537 VGND 0.06176f
C14213 VPWR.n2538 VGND 0.064f
C14214 VPWR.n2540 VGND 0.01268f
C14215 VPWR.n2542 VGND 0.08003f
C14216 VPWR.t636 VGND 0.08842f
C14217 VPWR.t628 VGND 0.05805f
C14218 VPWR.t655 VGND 0.06817f
C14219 VPWR.t663 VGND 0.05805f
C14220 VPWR.t796 VGND 0.08842f
C14221 VPWR.n2543 VGND 0.08003f
C14222 VPWR.n2545 VGND 0.01268f
C14223 VPWR.n2547 VGND 0.064f
C14224 VPWR.n2548 VGND 0.06176f
C14225 VPWR.n2549 VGND 0.06176f
C14226 VPWR.n2550 VGND 0.064f
C14227 VPWR.n2552 VGND 0.01268f
C14228 VPWR.n2554 VGND 0.08003f
C14229 VPWR.t812 VGND 0.08842f
C14230 VPWR.t765 VGND 0.05805f
C14231 VPWR.t893 VGND 0.06817f
C14232 VPWR.t926 VGND 0.05805f
C14233 VPWR.t942 VGND 0.08842f
C14234 VPWR.n2555 VGND 0.08003f
C14235 VPWR.n2557 VGND 0.01268f
C14236 VPWR.n2559 VGND 0.064f
C14237 VPWR.n2560 VGND 0.06176f
C14238 VPWR.n2561 VGND 0.06176f
C14239 VPWR.n2562 VGND 0.064f
C14240 VPWR.n2564 VGND 0.01268f
C14241 VPWR.n2566 VGND 0.08003f
C14242 VPWR.t686 VGND 0.08842f
C14243 VPWR.t945 VGND 0.05805f
C14244 VPWR.t678 VGND 0.06817f
C14245 VPWR.t799 VGND 0.05805f
C14246 VPWR.t716 VGND 0.08842f
C14247 VPWR.n2567 VGND 0.08003f
C14248 VPWR.n2569 VGND 0.01268f
C14249 VPWR.n2571 VGND 0.064f
C14250 VPWR.n2572 VGND 0.06176f
C14251 VPWR.n2573 VGND 0.06176f
C14252 VPWR.n2574 VGND 0.064f
C14253 VPWR.n2576 VGND 0.01268f
C14254 VPWR.n2578 VGND 0.08003f
C14255 VPWR.t566 VGND 0.08842f
C14256 VPWR.t818 VGND 0.05805f
C14257 VPWR.t939 VGND 0.06817f
C14258 VPWR.t843 VGND 0.05805f
C14259 VPWR.t585 VGND 0.08842f
C14260 VPWR.n2579 VGND 0.08003f
C14261 VPWR.n2581 VGND 0.01268f
C14262 VPWR.n2583 VGND 0.064f
C14263 VPWR.n2584 VGND 0.06176f
C14264 VPWR.n2585 VGND 0.06176f
C14265 VPWR.n2586 VGND 0.064f
C14266 VPWR.n2588 VGND 0.01268f
C14267 VPWR.n2590 VGND 0.08003f
C14268 VPWR.t710 VGND 0.08842f
C14269 VPWR.t694 VGND 0.05805f
C14270 VPWR.t815 VGND 0.0986f
C14271 VPWR.n2591 VGND 0.05631f
C14272 VPWR.n2592 VGND 0.01256f
C14273 VPWR.n2594 VGND 0.08026f
C14274 VPWR.n2595 VGND 0.14325f
C14275 VPWR.n2596 VGND 1.96905f
C14276 VPWR.n2597 VGND 0.80188f
C14277 VPWR.n2598 VGND 0.33599f
C14278 VPWR.t540 VGND 0.04034f
C14279 VPWR.t1017 VGND 0.04034f
C14280 VPWR.n2599 VGND 0.07319f
C14281 VPWR.n2600 VGND 0.03466f
C14282 VPWR.t538 VGND 0.0106f
C14283 VPWR.t546 VGND 0.0106f
C14284 VPWR.n2601 VGND 0.02274f
C14285 VPWR.t1022 VGND 0.0106f
C14286 VPWR.t1016 VGND 0.0106f
C14287 VPWR.n2602 VGND 0.02274f
C14288 VPWR.n2604 VGND 0.03466f
C14289 VPWR.t1828 VGND 0.0106f
C14290 VPWR.t1809 VGND 0.0106f
C14291 VPWR.n2605 VGND 0.02274f
C14292 VPWR.t1792 VGND 0.0106f
C14293 VPWR.t1798 VGND 0.0106f
C14294 VPWR.n2606 VGND 0.02274f
C14295 VPWR.t1805 VGND 0.04225f
C14296 VPWR.t1784 VGND 0.04225f
C14297 VPWR.n2607 VGND 0.09744f
C14298 VPWR.n2608 VGND 0.03127f
C14299 VPWR.n2609 VGND 0.01007f
C14300 VPWR.n2610 VGND 0.04572f
C14301 VPWR.t1786 VGND 0.0106f
C14302 VPWR.t544 VGND 0.0106f
C14303 VPWR.n2612 VGND 0.02274f
C14304 VPWR.t1804 VGND 0.0106f
C14305 VPWR.t1020 VGND 0.0106f
C14306 VPWR.n2613 VGND 0.02274f
C14307 VPWR.n2614 VGND 0.04572f
C14308 VPWR.n2615 VGND 0.01054f
C14309 VPWR.n2616 VGND 0.03466f
C14310 VPWR.n2617 VGND 0.03466f
C14311 VPWR.n2618 VGND 0.03466f
C14312 VPWR.n2620 VGND 0.04572f
C14313 VPWR.n2623 VGND 0.03466f
C14314 VPWR.n2624 VGND 0.02599f
C14315 VPWR.t1783 VGND 0.1266f
C14316 VPWR.t1791 VGND 0.18657f
C14317 VPWR.t1797 VGND 0.18657f
C14318 VPWR.t1785 VGND 0.18657f
C14319 VPWR.t543 VGND 0.18657f
C14320 VPWR.t537 VGND 0.18657f
C14321 VPWR.t545 VGND 0.18657f
C14322 VPWR.t539 VGND 0.41537f
C14323 VPWR.n2626 VGND 0.45337f
C14324 VPWR.n2627 VGND 0.01319f
C14325 VPWR.n2628 VGND 0.7952f
C14326 VPWR.n2629 VGND 0.03466f
C14327 VPWR.t1781 VGND 0.1266f
C14328 VPWR.t1794 VGND 0.18657f
C14329 VPWR.t1768 VGND 0.18657f
C14330 VPWR.t1820 VGND 0.18657f
C14331 VPWR.t1238 VGND 0.18657f
C14332 VPWR.t1230 VGND 0.18657f
C14333 VPWR.t1242 VGND 0.18657f
C14334 VPWR.t1234 VGND 0.30651f
C14335 VPWR.t525 VGND 0.32539f
C14336 VPWR.n2630 VGND 0.45918f
C14337 VPWR.n2631 VGND 0.13062f
C14338 VPWR.n2632 VGND 0.03466f
C14339 VPWR.t1490 VGND 0.0106f
C14340 VPWR.t1269 VGND 0.0106f
C14341 VPWR.n2633 VGND 0.02274f
C14342 VPWR.t1231 VGND 0.0106f
C14343 VPWR.t1243 VGND 0.0106f
C14344 VPWR.n2634 VGND 0.02274f
C14345 VPWR.n2635 VGND 0.04572f
C14346 VPWR.n2636 VGND 0.03466f
C14347 VPWR.t1831 VGND 0.0106f
C14348 VPWR.t1270 VGND 0.0106f
C14349 VPWR.n2637 VGND 0.02274f
C14350 VPWR.t1821 VGND 0.0106f
C14351 VPWR.t1239 VGND 0.0106f
C14352 VPWR.n2638 VGND 0.02274f
C14353 VPWR.t1782 VGND 0.04225f
C14354 VPWR.t1830 VGND 0.04225f
C14355 VPWR.n2640 VGND 0.09744f
C14356 VPWR.t1813 VGND 0.0106f
C14357 VPWR.t1788 VGND 0.0106f
C14358 VPWR.n2641 VGND 0.02274f
C14359 VPWR.t1795 VGND 0.0106f
C14360 VPWR.t1769 VGND 0.0106f
C14361 VPWR.n2642 VGND 0.02274f
C14362 VPWR.n2643 VGND 0.04572f
C14363 VPWR.n2644 VGND 0.01007f
C14364 VPWR.n2645 VGND 0.03127f
C14365 VPWR.n2646 VGND 0.03466f
C14366 VPWR.n2647 VGND 0.03466f
C14367 VPWR.n2648 VGND 0.01054f
C14368 VPWR.n2649 VGND 0.04572f
C14369 VPWR.n2652 VGND 0.03466f
C14370 VPWR.n2653 VGND 0.03466f
C14371 VPWR.t1489 VGND 0.04034f
C14372 VPWR.t1235 VGND 0.04034f
C14373 VPWR.n2656 VGND 0.07319f
C14374 VPWR.n2658 VGND 0.02599f
C14375 VPWR.n2659 VGND 0.01319f
C14376 VPWR.n2660 VGND 0.02599f
C14377 VPWR.n2661 VGND 0.01034f
C14378 VPWR.t1012 VGND 0.04221f
C14379 VPWR.t526 VGND 0.04221f
C14380 VPWR.n2663 VGND 0.08532f
C14381 VPWR.n2664 VGND 0.02411f
C14382 VPWR.n2665 VGND 1.21026f
C14383 VPWR.n2666 VGND 0.03466f
C14384 VPWR.t1742 VGND 0.04143f
C14385 VPWR.t1815 VGND 0.1266f
C14386 VPWR.t1772 VGND 0.18657f
C14387 VPWR.t1822 VGND 0.18657f
C14388 VPWR.t1799 VGND 0.18657f
C14389 VPWR.t2 VGND 0.18657f
C14390 VPWR.t1506 VGND 0.18657f
C14391 VPWR.t1244 VGND 0.18657f
C14392 VPWR.t1226 VGND 0.30651f
C14393 VPWR.t1907 VGND 0.11772f
C14394 VPWR.t1741 VGND 0.09329f
C14395 VPWR.t457 VGND 0.20767f
C14396 VPWR.n2667 VGND 0.40698f
C14397 VPWR.n2668 VGND 0.12868f
C14398 VPWR.n2669 VGND 0.03466f
C14399 VPWR.t1665 VGND 0.0106f
C14400 VPWR.t1669 VGND 0.0106f
C14401 VPWR.n2670 VGND 0.02274f
C14402 VPWR.t1507 VGND 0.0106f
C14403 VPWR.t1245 VGND 0.0106f
C14404 VPWR.n2671 VGND 0.02274f
C14405 VPWR.n2672 VGND 0.04572f
C14406 VPWR.n2673 VGND 0.03466f
C14407 VPWR.t1817 VGND 0.0106f
C14408 VPWR.t1668 VGND 0.0106f
C14409 VPWR.n2674 VGND 0.02274f
C14410 VPWR.t1800 VGND 0.0106f
C14411 VPWR.t3 VGND 0.0106f
C14412 VPWR.n2675 VGND 0.02274f
C14413 VPWR.t1829 VGND 0.04225f
C14414 VPWR.t1816 VGND 0.04225f
C14415 VPWR.n2677 VGND 0.09744f
C14416 VPWR.t1789 VGND 0.0106f
C14417 VPWR.t1835 VGND 0.0106f
C14418 VPWR.n2678 VGND 0.02274f
C14419 VPWR.t1773 VGND 0.0106f
C14420 VPWR.t1823 VGND 0.0106f
C14421 VPWR.n2679 VGND 0.02274f
C14422 VPWR.n2680 VGND 0.04572f
C14423 VPWR.n2681 VGND 0.01007f
C14424 VPWR.n2682 VGND 0.03127f
C14425 VPWR.n2683 VGND 0.03466f
C14426 VPWR.n2684 VGND 0.03466f
C14427 VPWR.n2685 VGND 0.01054f
C14428 VPWR.n2686 VGND 0.04572f
C14429 VPWR.n2689 VGND 0.03466f
C14430 VPWR.n2690 VGND 0.03466f
C14431 VPWR.t1666 VGND 0.04034f
C14432 VPWR.t1227 VGND 0.04034f
C14433 VPWR.n2693 VGND 0.07319f
C14434 VPWR.n2695 VGND 0.02599f
C14435 VPWR.n2696 VGND 0.01319f
C14436 VPWR.n2697 VGND 0.02599f
C14437 VPWR.t458 VGND 0.04226f
C14438 VPWR.n2698 VGND 0.05889f
C14439 VPWR.n2700 VGND 0.04309f
C14440 VPWR.t1908 VGND 0.04154f
C14441 VPWR.n2701 VGND 0.05384f
C14442 VPWR.n2702 VGND 0.02053f
C14443 VPWR.n2703 VGND 1.21026f
C14444 VPWR.n2704 VGND 0.03466f
C14445 VPWR.t1818 VGND 0.0718f
C14446 VPWR.t1776 VGND 0.10581f
C14447 VPWR.t1824 VGND 0.10287f
C14448 VPWR.t1802 VGND 0.16452f
C14449 VPWR.t1369 VGND 0.13993f
C14450 VPWR.t1806 VGND 0.09329f
C14451 VPWR.t1363 VGND 0.09329f
C14452 VPWR.t1778 VGND 0.09329f
C14453 VPWR.t1371 VGND 0.09329f
C14454 VPWR.t1810 VGND 0.09329f
C14455 VPWR.t1365 VGND 0.09329f
C14456 VPWR.t1833 VGND 0.12993f
C14457 VPWR.t1407 VGND 0.0733f
C14458 VPWR.t1891 VGND 0.07996f
C14459 VPWR.t455 VGND 0.09329f
C14460 VPWR.t1893 VGND 0.17324f
C14461 VPWR.n2705 VGND 0.27927f
C14462 VPWR.n2706 VGND 0.12882f
C14463 VPWR.t1894 VGND 0.04194f
C14464 VPWR.n2707 VGND 0.03466f
C14465 VPWR.t1834 VGND 0.04146f
C14466 VPWR.t1366 VGND 0.03991f
C14467 VPWR.t1779 VGND 0.0106f
C14468 VPWR.t1811 VGND 0.0106f
C14469 VPWR.n2708 VGND 0.02274f
C14470 VPWR.t1364 VGND 0.0106f
C14471 VPWR.t1372 VGND 0.0106f
C14472 VPWR.n2709 VGND 0.02274f
C14473 VPWR.n2710 VGND 0.02593f
C14474 VPWR.n2711 VGND 0.03466f
C14475 VPWR.t1803 VGND 0.0106f
C14476 VPWR.t1370 VGND 0.0106f
C14477 VPWR.n2712 VGND 0.02274f
C14478 VPWR.t1819 VGND 0.04225f
C14479 VPWR.n2714 VGND 0.05325f
C14480 VPWR.t1777 VGND 0.0106f
C14481 VPWR.t1825 VGND 0.0106f
C14482 VPWR.n2715 VGND 0.02274f
C14483 VPWR.n2716 VGND 0.02593f
C14484 VPWR.n2717 VGND 0.01007f
C14485 VPWR.n2718 VGND 0.03127f
C14486 VPWR.n2719 VGND 0.03466f
C14487 VPWR.n2720 VGND 0.03466f
C14488 VPWR.n2721 VGND 0.01054f
C14489 VPWR.n2722 VGND 0.02533f
C14490 VPWR.t1807 VGND 0.03708f
C14491 VPWR.n2723 VGND 0.02956f
C14492 VPWR.n2725 VGND 0.03466f
C14493 VPWR.n2726 VGND 0.03466f
C14494 VPWR.n2727 VGND 0.02873f
C14495 VPWR.n2729 VGND 0.03803f
C14496 VPWR.n2730 VGND 0.0501f
C14497 VPWR.n2732 VGND 0.02053f
C14498 VPWR.n2733 VGND 0.01319f
C14499 VPWR.n2734 VGND 0.02599f
C14500 VPWR.t456 VGND 0.0423f
C14501 VPWR.n2735 VGND 0.10875f
C14502 VPWR.t1892 VGND 0.04223f
C14503 VPWR.n2737 VGND 0.04701f
C14504 VPWR.n2738 VGND 0.02034f
C14505 VPWR.n2739 VGND 1.21026f
C14506 VPWR.n2740 VGND 0.03127f
C14507 VPWR.t1812 VGND 0.49308f
C14508 VPWR.t1771 VGND 0.18657f
C14509 VPWR.t1801 VGND 0.18657f
C14510 VPWR.t1775 VGND 0.18657f
C14511 VPWR.t547 VGND 0.18657f
C14512 VPWR.t541 VGND 0.18657f
C14513 VPWR.t549 VGND 0.18657f
C14514 VPWR.t551 VGND 0.1688f
C14515 VPWR.t1390 VGND 0.40868f
C14516 VPWR.t1212 VGND 0.11327f
C14517 VPWR.n2741 VGND 0.24485f
C14518 VPWR.n2742 VGND 0.13062f
C14519 VPWR.t548 VGND 0.0106f
C14520 VPWR.t542 VGND 0.0106f
C14521 VPWR.n2743 VGND 0.02322f
C14522 VPWR.t1019 VGND 0.0106f
C14523 VPWR.t1018 VGND 0.0106f
C14524 VPWR.n2744 VGND 0.02322f
C14525 VPWR.n2745 VGND 0.08815f
C14526 VPWR.n2746 VGND 0.07146f
C14527 VPWR.t550 VGND 0.0106f
C14528 VPWR.t552 VGND 0.0106f
C14529 VPWR.n2747 VGND 0.02326f
C14530 VPWR.t1021 VGND 0.0106f
C14531 VPWR.t1015 VGND 0.0106f
C14532 VPWR.n2748 VGND 0.02326f
C14533 VPWR.n2749 VGND 0.09662f
C14534 VPWR.n2751 VGND 0.27909f
C14535 VPWR.n2752 VGND 0.01319f
C14536 VPWR.n2753 VGND 0.01206f
C14537 VPWR.n2754 VGND 0.01034f
C14538 VPWR.t1661 VGND 0.0423f
C14539 VPWR.t1391 VGND 0.0423f
C14540 VPWR.n2756 VGND 0.12493f
C14541 VPWR.n2757 VGND 0.02599f
C14542 VPWR.n2758 VGND 1.21026f
C14543 VPWR.n2759 VGND 0.03127f
C14544 VPWR.t1793 VGND 0.49308f
C14545 VPWR.t1826 VGND 0.18657f
C14546 VPWR.t1780 VGND 0.18657f
C14547 VPWR.t1827 VGND 0.18657f
C14548 VPWR.t1228 VGND 0.18657f
C14549 VPWR.t1240 VGND 0.18657f
C14550 VPWR.t1232 VGND 0.18657f
C14551 VPWR.t1236 VGND 0.1688f
C14552 VPWR.t14 VGND 0.36315f
C14553 VPWR.t1214 VGND 0.07996f
C14554 VPWR.t1218 VGND 0.07885f
C14555 VPWR.n2760 VGND 0.24374f
C14556 VPWR.n2761 VGND 0.13062f
C14557 VPWR.t1284 VGND 0.0106f
C14558 VPWR.t1488 VGND 0.0106f
C14559 VPWR.n2762 VGND 0.02322f
C14560 VPWR.t1229 VGND 0.0106f
C14561 VPWR.t1241 VGND 0.0106f
C14562 VPWR.n2763 VGND 0.02322f
C14563 VPWR.n2764 VGND 0.08815f
C14564 VPWR.n2765 VGND 0.07146f
C14565 VPWR.t1283 VGND 0.0106f
C14566 VPWR.t1491 VGND 0.0106f
C14567 VPWR.n2766 VGND 0.02326f
C14568 VPWR.t1233 VGND 0.0106f
C14569 VPWR.t1237 VGND 0.0106f
C14570 VPWR.n2767 VGND 0.02326f
C14571 VPWR.n2768 VGND 0.09662f
C14572 VPWR.n2770 VGND 0.27909f
C14573 VPWR.n2771 VGND 0.01319f
C14574 VPWR.n2772 VGND 0.01187f
C14575 VPWR.t1215 VGND 0.04221f
C14576 VPWR.n2774 VGND 0.04512f
C14577 VPWR.t15 VGND 0.0423f
C14578 VPWR.n2776 VGND 0.06737f
C14579 VPWR.n2777 VGND 0.02599f
C14580 VPWR.n2778 VGND 1.21026f
C14581 VPWR.n2779 VGND 0.03164f
C14582 VPWR.t1774 VGND 0.49308f
C14583 VPWR.t1787 VGND 0.18657f
C14584 VPWR.t1814 VGND 0.18657f
C14585 VPWR.t1790 VGND 0.18657f
C14586 VPWR.t1092 VGND 0.18657f
C14587 VPWR.t1355 VGND 0.18657f
C14588 VPWR.t91 VGND 0.18657f
C14589 VPWR.t453 VGND 0.1688f
C14590 VPWR.t1388 VGND 0.38647f
C14591 VPWR.t1210 VGND 0.13327f
C14592 VPWR.n2780 VGND 0.24262f
C14593 VPWR.n2781 VGND 0.12868f
C14594 VPWR.t1213 VGND 0.04227f
C14595 VPWR.t1670 VGND 0.0106f
C14596 VPWR.t1667 VGND 0.0106f
C14597 VPWR.n2782 VGND 0.02322f
C14598 VPWR.t1093 VGND 0.0106f
C14599 VPWR.t1356 VGND 0.0106f
C14600 VPWR.n2783 VGND 0.02322f
C14601 VPWR.n2784 VGND 0.08815f
C14602 VPWR.n2785 VGND 0.07146f
C14603 VPWR.t1663 VGND 0.0106f
C14604 VPWR.t1664 VGND 0.0106f
C14605 VPWR.n2786 VGND 0.02326f
C14606 VPWR.t92 VGND 0.0106f
C14607 VPWR.t454 VGND 0.0106f
C14608 VPWR.n2787 VGND 0.02326f
C14609 VPWR.n2788 VGND 0.09662f
C14610 VPWR.n2790 VGND 0.27909f
C14611 VPWR.n2791 VGND 0.01319f
C14612 VPWR.n2792 VGND 0.01168f
C14613 VPWR.t1211 VGND 0.04227f
C14614 VPWR.n2793 VGND 0.11136f
C14615 VPWR.t1662 VGND 0.04226f
C14616 VPWR.t1389 VGND 0.04226f
C14617 VPWR.n2795 VGND 0.09943f
C14618 VPWR.n2796 VGND 0.02599f
C14619 VPWR.n2797 VGND 1.21026f
C14620 VPWR.n2798 VGND 0.03164f
C14621 VPWR.t13 VGND 0.04226f
C14622 VPWR.n2799 VGND 0.01168f
C14623 VPWR.t1217 VGND 0.04227f
C14624 VPWR.n2800 VGND 0.01319f
C14625 VPWR.t1808 VGND 0.27964f
C14626 VPWR.t1832 VGND 0.10581f
C14627 VPWR.t1796 VGND 0.10581f
C14628 VPWR.t1770 VGND 0.10581f
C14629 VPWR.t1367 VGND 0.10581f
C14630 VPWR.t1361 VGND 0.10581f
C14631 VPWR.t1373 VGND 0.10581f
C14632 VPWR.t1375 VGND 0.09573f
C14633 VPWR.t12 VGND 0.21918f
C14634 VPWR.t1216 VGND 0.07558f
C14635 VPWR.n2801 VGND 0.13503f
C14636 VPWR.t1374 VGND 0.0106f
C14637 VPWR.t1376 VGND 0.0106f
C14638 VPWR.n2802 VGND 0.02326f
C14639 VPWR.n2803 VGND 0.05725f
C14640 VPWR.t1368 VGND 0.0106f
C14641 VPWR.t1362 VGND 0.0106f
C14642 VPWR.n2804 VGND 0.02421f
C14643 VPWR.n2805 VGND 0.12927f
C14644 VPWR.n2806 VGND 0.27909f
C14645 VPWR.n2808 VGND 0.07145f
C14646 VPWR.n2809 VGND 0.06272f
C14647 VPWR.n2811 VGND 0.05435f
C14648 VPWR.n2812 VGND 0.02599f
C14649 VPWR.n2813 VGND 1.76121f
C14650 VPWR.n2814 VGND 1.42636f
C14651 VPWR.t267 VGND 0.02149f
C14652 VPWR.n2815 VGND 0.09631f
C14653 VPWR.n2816 VGND 0.21199f
C14654 VPWR.n2817 VGND 0.0559f
C14655 VPWR.n2818 VGND 0.02655f
C14656 VPWR.n2819 VGND 0.03242f
C14657 VPWR.n2820 VGND 0.06571f
C14658 VPWR.n2821 VGND 0.08566f
C14659 VPWR.n2822 VGND 0.06571f
C14660 VPWR.t93 VGND 2.0669f
C14661 VPWR.t266 VGND 0.65281f
C14662 VPWR.n2823 VGND 0.08633f
C14663 VPWR.n2824 VGND 0.34157f
C14664 VPWR.t94 VGND 0.02148f
C14665 VPWR.n2825 VGND 0.1315f
C14666 VPWR.n2826 VGND 0.01328f
C14667 VPWR.n2827 VGND 0.07245f
C14668 VPWR.n2828 VGND 0.06504f
C14669 VPWR.n2829 VGND 0.08633f
C14670 VPWR.n2830 VGND 0.05437f
C14671 VPWR.t1473 VGND 0.02148f
C14672 VPWR.n2831 VGND 0.1315f
C14673 VPWR.n2832 VGND 0.01328f
C14674 VPWR.n2833 VGND 0.08633f
C14675 VPWR.n2834 VGND 0.0565f
C14676 VPWR.n2835 VGND 0.06443f
C14677 VPWR.n2836 VGND 1.23519f
C14678 VPWR.n2837 VGND 0.06443f
C14679 VPWR.n2838 VGND 0.0565f
C14680 VPWR.n2839 VGND 0.08633f
C14681 VPWR.n2840 VGND 0.07238f
C14682 VPWR.n2841 VGND 0.05987f
C14683 VPWR.n2842 VGND 0.74248f
C14684 VPWR.n2843 VGND 0.04672f
C14685 VPWR.n2844 VGND 0.06535f
C14686 VPWR.n2845 VGND 0.04543f
C14687 VPWR.n2846 VGND 0.01328f
C14688 VPWR.n2847 VGND 0.04672f
C14689 VPWR.n2848 VGND 0.03587f
C14690 VPWR.n2849 VGND 0.12835f
C14691 VPWR.n2850 VGND 0.05056f
C14692 VPWR.n2851 VGND 0.03242f
C14693 VPWR.t1094 VGND 0.25559f
C14694 VPWR.n2852 VGND 0.05987f
C14695 VPWR.n2853 VGND 0.07238f
C14696 VPWR.n2854 VGND 0.02655f
C14697 VPWR.n2855 VGND 1.49593f
C14698 VPWR.n2856 VGND 0.02655f
C14699 VPWR.n2857 VGND 0.02655f
C14700 VPWR.n2858 VGND 0.06598f
C14701 VPWR.n2859 VGND 0.03622f
C14702 VPWR.n2860 VGND 0.28054f
C14703 VPWR.n2861 VGND 0.23083f
C14704 VPWR.t1095 VGND 0.02147f
C14705 VPWR.n2862 VGND 0.16245f
C14706 VPWR.n2863 VGND 2.5721f
C14707 XThR.Tn[2].t7 VGND 0.01796f
C14708 XThR.Tn[2].t4 VGND 0.01796f
C14709 XThR.Tn[2].n0 VGND 0.03626f
C14710 XThR.Tn[2].t6 VGND 0.01796f
C14711 XThR.Tn[2].t5 VGND 0.01796f
C14712 XThR.Tn[2].n1 VGND 0.04242f
C14713 XThR.Tn[2].n2 VGND 0.12726f
C14714 XThR.Tn[2].t10 VGND 0.01168f
C14715 XThR.Tn[2].t11 VGND 0.01168f
C14716 XThR.Tn[2].n3 VGND 0.02659f
C14717 XThR.Tn[2].t9 VGND 0.01168f
C14718 XThR.Tn[2].t8 VGND 0.01168f
C14719 XThR.Tn[2].n4 VGND 0.02659f
C14720 XThR.Tn[2].t1 VGND 0.01168f
C14721 XThR.Tn[2].t2 VGND 0.01168f
C14722 XThR.Tn[2].n5 VGND 0.0443f
C14723 XThR.Tn[2].t0 VGND 0.01168f
C14724 XThR.Tn[2].t3 VGND 0.01168f
C14725 XThR.Tn[2].n6 VGND 0.02659f
C14726 XThR.Tn[2].n7 VGND 0.12662f
C14727 XThR.Tn[2].n8 VGND 0.07828f
C14728 XThR.Tn[2].n9 VGND 0.08834f
C14729 XThR.Tn[2].t21 VGND 0.01404f
C14730 XThR.Tn[2].t14 VGND 0.01537f
C14731 XThR.Tn[2].n10 VGND 0.03754f
C14732 XThR.Tn[2].n11 VGND 0.07211f
C14733 XThR.Tn[2].t40 VGND 0.01404f
C14734 XThR.Tn[2].t31 VGND 0.01537f
C14735 XThR.Tn[2].n12 VGND 0.03754f
C14736 XThR.Tn[2].t55 VGND 0.01399f
C14737 XThR.Tn[2].t66 VGND 0.01532f
C14738 XThR.Tn[2].n13 VGND 0.03906f
C14739 XThR.Tn[2].n14 VGND 0.02744f
C14740 XThR.Tn[2].n16 VGND 0.08806f
C14741 XThR.Tn[2].t15 VGND 0.01404f
C14742 XThR.Tn[2].t67 VGND 0.01537f
C14743 XThR.Tn[2].n17 VGND 0.03754f
C14744 XThR.Tn[2].t30 VGND 0.01399f
C14745 XThR.Tn[2].t43 VGND 0.01532f
C14746 XThR.Tn[2].n18 VGND 0.03906f
C14747 XThR.Tn[2].n19 VGND 0.02744f
C14748 XThR.Tn[2].n21 VGND 0.08806f
C14749 XThR.Tn[2].t32 VGND 0.01404f
C14750 XThR.Tn[2].t23 VGND 0.01537f
C14751 XThR.Tn[2].n22 VGND 0.03754f
C14752 XThR.Tn[2].t47 VGND 0.01399f
C14753 XThR.Tn[2].t60 VGND 0.01532f
C14754 XThR.Tn[2].n23 VGND 0.03906f
C14755 XThR.Tn[2].n24 VGND 0.02744f
C14756 XThR.Tn[2].n26 VGND 0.08806f
C14757 XThR.Tn[2].t58 VGND 0.01404f
C14758 XThR.Tn[2].t50 VGND 0.01537f
C14759 XThR.Tn[2].n27 VGND 0.03754f
C14760 XThR.Tn[2].t16 VGND 0.01399f
C14761 XThR.Tn[2].t28 VGND 0.01532f
C14762 XThR.Tn[2].n28 VGND 0.03906f
C14763 XThR.Tn[2].n29 VGND 0.02744f
C14764 XThR.Tn[2].n31 VGND 0.08806f
C14765 XThR.Tn[2].t34 VGND 0.01404f
C14766 XThR.Tn[2].t25 VGND 0.01537f
C14767 XThR.Tn[2].n32 VGND 0.03754f
C14768 XThR.Tn[2].t48 VGND 0.01399f
C14769 XThR.Tn[2].t62 VGND 0.01532f
C14770 XThR.Tn[2].n33 VGND 0.03906f
C14771 XThR.Tn[2].n34 VGND 0.02744f
C14772 XThR.Tn[2].n36 VGND 0.08806f
C14773 XThR.Tn[2].t70 VGND 0.01404f
C14774 XThR.Tn[2].t41 VGND 0.01537f
C14775 XThR.Tn[2].n37 VGND 0.03754f
C14776 XThR.Tn[2].t22 VGND 0.01399f
C14777 XThR.Tn[2].t20 VGND 0.01532f
C14778 XThR.Tn[2].n38 VGND 0.03906f
C14779 XThR.Tn[2].n39 VGND 0.02744f
C14780 XThR.Tn[2].n41 VGND 0.08806f
C14781 XThR.Tn[2].t39 VGND 0.01404f
C14782 XThR.Tn[2].t35 VGND 0.01537f
C14783 XThR.Tn[2].n42 VGND 0.03754f
C14784 XThR.Tn[2].t54 VGND 0.01399f
C14785 XThR.Tn[2].t12 VGND 0.01532f
C14786 XThR.Tn[2].n43 VGND 0.03906f
C14787 XThR.Tn[2].n44 VGND 0.02744f
C14788 XThR.Tn[2].n46 VGND 0.08806f
C14789 XThR.Tn[2].t44 VGND 0.01404f
C14790 XThR.Tn[2].t49 VGND 0.01537f
C14791 XThR.Tn[2].n47 VGND 0.03754f
C14792 XThR.Tn[2].t57 VGND 0.01399f
C14793 XThR.Tn[2].t27 VGND 0.01532f
C14794 XThR.Tn[2].n48 VGND 0.03906f
C14795 XThR.Tn[2].n49 VGND 0.02744f
C14796 XThR.Tn[2].n51 VGND 0.08806f
C14797 XThR.Tn[2].t61 VGND 0.01404f
C14798 XThR.Tn[2].t69 VGND 0.01537f
C14799 XThR.Tn[2].n52 VGND 0.03754f
C14800 XThR.Tn[2].t18 VGND 0.01399f
C14801 XThR.Tn[2].t45 VGND 0.01532f
C14802 XThR.Tn[2].n53 VGND 0.03906f
C14803 XThR.Tn[2].n54 VGND 0.02744f
C14804 XThR.Tn[2].n56 VGND 0.08806f
C14805 XThR.Tn[2].t52 VGND 0.01404f
C14806 XThR.Tn[2].t26 VGND 0.01537f
C14807 XThR.Tn[2].n57 VGND 0.03754f
C14808 XThR.Tn[2].t68 VGND 0.01399f
C14809 XThR.Tn[2].t63 VGND 0.01532f
C14810 XThR.Tn[2].n58 VGND 0.03906f
C14811 XThR.Tn[2].n59 VGND 0.02744f
C14812 XThR.Tn[2].n61 VGND 0.08806f
C14813 XThR.Tn[2].t73 VGND 0.01404f
C14814 XThR.Tn[2].t64 VGND 0.01537f
C14815 XThR.Tn[2].n62 VGND 0.03754f
C14816 XThR.Tn[2].t24 VGND 0.01399f
C14817 XThR.Tn[2].t37 VGND 0.01532f
C14818 XThR.Tn[2].n63 VGND 0.03906f
C14819 XThR.Tn[2].n64 VGND 0.02744f
C14820 XThR.Tn[2].n66 VGND 0.08806f
C14821 XThR.Tn[2].t42 VGND 0.01404f
C14822 XThR.Tn[2].t36 VGND 0.01537f
C14823 XThR.Tn[2].n67 VGND 0.03754f
C14824 XThR.Tn[2].t56 VGND 0.01399f
C14825 XThR.Tn[2].t13 VGND 0.01532f
C14826 XThR.Tn[2].n68 VGND 0.03906f
C14827 XThR.Tn[2].n69 VGND 0.02744f
C14828 XThR.Tn[2].n71 VGND 0.08806f
C14829 XThR.Tn[2].t59 VGND 0.01404f
C14830 XThR.Tn[2].t51 VGND 0.01537f
C14831 XThR.Tn[2].n72 VGND 0.03754f
C14832 XThR.Tn[2].t17 VGND 0.01399f
C14833 XThR.Tn[2].t29 VGND 0.01532f
C14834 XThR.Tn[2].n73 VGND 0.03906f
C14835 XThR.Tn[2].n74 VGND 0.02744f
C14836 XThR.Tn[2].n76 VGND 0.08806f
C14837 XThR.Tn[2].t19 VGND 0.01404f
C14838 XThR.Tn[2].t72 VGND 0.01537f
C14839 XThR.Tn[2].n77 VGND 0.03754f
C14840 XThR.Tn[2].t33 VGND 0.01399f
C14841 XThR.Tn[2].t46 VGND 0.01532f
C14842 XThR.Tn[2].n78 VGND 0.03906f
C14843 XThR.Tn[2].n79 VGND 0.02744f
C14844 XThR.Tn[2].n81 VGND 0.08806f
C14845 XThR.Tn[2].t53 VGND 0.01404f
C14846 XThR.Tn[2].t65 VGND 0.01537f
C14847 XThR.Tn[2].n82 VGND 0.03754f
C14848 XThR.Tn[2].t71 VGND 0.01399f
C14849 XThR.Tn[2].t38 VGND 0.01532f
C14850 XThR.Tn[2].n83 VGND 0.03906f
C14851 XThR.Tn[2].n84 VGND 0.02744f
C14852 XThR.Tn[2].n86 VGND 0.08806f
C14853 XThR.Tn[2].n87 VGND 0.08002f
C14854 XThR.Tn[2].n88 VGND 0.17341f
.ends

