* NGSPICE file created from csdac255_parax.ext - technology: sky130A

.subckt csdac255_parax Iout VPWR VGND Vbias data[0] data[1] data[2] data[3] data[4]
+ data[5] data[6] data[7] bias[0] bias[1] bias[2]
X0 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout VGND.t1712 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1 VPWR.t830 XThR.Tn[2].t12 XA.XIR[3].XIC[8].icell.PUM VPWR.t829 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2 XA.XIR[12].XIC[10].icell.SM XA.XIR[12].XIC[10].icell.Ien Iout.t225 VGND.t2232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X3 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1721 VPWR.t1723 VPWR.t1722 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X4 VGND.t298 XThC.Tn[10].t12 XA.XIR[4].XIC[10].icell.PDM VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X5 VGND.t450 XThR.XTBN.Y.t4 a_n997_2667# VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t1255 XThR.Tn[6].t12 XA.XIR[7].XIC[8].icell.PUM VPWR.t1254 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X7 XA.XIR[14].XIC[5].icell.Ien XThR.Tn[14].t12 VPWR.t162 VPWR.t161 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X8 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12].t12 XA.XIR[12].XIC[6].icell.Ien VGND.t1501 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X9 XThC.Tn[6].t11 XThC.XTBN.Y.t4 VGND.t485 VGND.t484 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1926 VGND.t1653 VGND.t1652 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X11 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[9].t12 VGND.t785 VGND.t784 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X12 VGND.t486 XThC.XTBN.Y.t5 XThC.Tn[5].t11 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 XA.XIR[15].XIC[9].icell.PUM XThC.Tn[9].t12 XA.XIR[15].XIC[9].icell.Ien VPWR.t26 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X14 XA.XIR[9].XIC[0].icell.SM XA.XIR[9].XIC[0].icell.Ien Iout.t76 VGND.t720 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X15 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[12].t13 VGND.t1503 VGND.t1502 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X16 VGND.t2433 XThC.Tn[11].t12 XA.XIR[12].XIC[11].icell.PDM VGND.t2432 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X17 XA.XIR[12].XIC[1].icell.SM XA.XIR[12].XIC[1].icell.Ien Iout.t213 VGND.t2093 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X18 XA.XIR[8].XIC[12].icell.SM XA.XIR[8].XIC[12].icell.Ien Iout.t43 VGND.t249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X19 XThC.Tn[12].t7 XThC.XTB5.Y VPWR.t417 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 XA.XIR[8].XIC_15.icell.PDM VPWR.t1927 VGND.t1655 VGND.t1654 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X21 XA.XIR[7].XIC[13].icell.SM XA.XIR[7].XIC[13].icell.Ien Iout.t227 VGND.t2370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X22 XA.XIR[14].XIC[13].icell.PUM XThC.Tn[13].t12 XA.XIR[14].XIC[13].icell.Ien VPWR.t998 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X23 a_2979_9615# XThC.XTBN.Y.t6 XThC.Tn[0].t3 VPWR.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1719 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1720 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X25 XA.XIR[10].XIC[14].icell.SM XA.XIR[10].XIC[14].icell.Ien Iout.t188 VGND.t1602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X26 a_4861_9615# XThC.XTB4.Y.t2 VPWR.t1845 VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_5949_9615# XThC.XTBN.Y.t7 XThC.Tn[5].t7 VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6].t13 XA.XIR[6].XIC[10].icell.Ien VGND.t2120 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X29 XA.XIR[0].XIC[4].icell.PDM VGND.t1904 VGND.t1906 VGND.t1905 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X30 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[3].t12 VGND.t2227 VGND.t2226 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X31 XThR.Tn[5].t11 XThR.XTBN.Y.t5 a_n1049_5611# VPWR.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 XThC.Tn[4].t3 XThC.XTB5.Y VGND.t567 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND.t487 XThC.XTBN.Y.t8 XThC.Tn[2].t8 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 XThR.XTB2.Y XThR.XTB6.A VPWR.t46 VPWR.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[6].t14 VGND.t2122 VGND.t2121 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X36 XA.XIR[6].XIC[11].icell.SM XA.XIR[6].XIC[11].icell.Ien Iout.t244 VGND.t2485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X37 VGND.t2685 XThC.Tn[2].t12 XA.XIR[12].XIC[2].icell.PDM VGND.t2684 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X38 VPWR.t1718 VPWR.t1716 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1717 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X39 VGND.t1657 VPWR.t1928 XA.XIR[7].XIC_dummy_left.icell.PDM VGND.t1656 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X40 VPWR.t1331 XThR.Tn[3].t13 XA.XIR[4].XIC[11].icell.PUM VPWR.t1330 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X41 VGND.t2390 Vbias.t6 XA.XIR[14].XIC[11].icell.SM VGND.t2389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X42 XA.XIR[2].XIC[1].icell.PUM XThC.Tn[1].t12 XA.XIR[2].XIC[1].icell.Ien VPWR.t940 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X43 VGND.t2134 XThC.Tn[3].t12 XA.XIR[15].XIC[3].icell.PDM VGND.t2133 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X44 VGND.t1659 VPWR.t1929 XA.XIR[10].XIC_15.icell.PDM VGND.t1658 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X45 VPWR.t1114 XThR.Tn[10].t12 XA.XIR[11].XIC[9].icell.PUM VPWR.t1113 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X46 XA.XIR[0].XIC[14].icell.PUM XThC.Tn[14].t12 XA.XIR[0].XIC[14].icell.Ien VPWR.t1836 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X47 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1713 VPWR.t1715 VPWR.t1714 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X48 a_7651_9569# XThC.XTB1.Y.t3 XThC.Tn[8].t3 VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 VGND.t2392 Vbias.t7 XA.XIR[2].XIC[5].icell.SM VGND.t2391 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X50 XA.XIR[1].XIC[6].icell.Ien XThR.Tn[1].t12 VPWR.t1138 VPWR.t1137 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X51 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t3 VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 VGND.t2475 XThC.Tn[4].t12 XA.XIR[2].XIC[4].icell.PDM VGND.t2474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X53 XThC.XTB5.Y XThC.XTB7.B VGND.t1140 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 XThC.Tn[7].t7 XThC.XTBN.Y.t9 VPWR.t331 VPWR.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X55 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[9].t13 VGND.t787 VGND.t786 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X56 VGND.t1558 XThR.XTB7.Y XThR.Tn[6].t3 VGND.t1557 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X57 XA.XIR[4].XIC[7].icell.Ien XThR.Tn[4].t12 VPWR.t719 VPWR.t718 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X58 VPWR.t310 XThR.XTBN.Y.t6 XThR.Tn[9].t11 VPWR.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 XThR.XTB7.Y XThR.XTB7.A VGND.t1196 VGND.t1195 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 XA.XIR[3].XIC[8].icell.Ien XThR.Tn[3].t14 VPWR.t1333 VPWR.t1332 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X61 VPWR.t1335 XThR.Tn[3].t15 XA.XIR[4].XIC[2].icell.PUM VPWR.t1334 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X62 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[12].t14 VGND.t1505 VGND.t1504 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X63 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[1].t13 XA.XIR[1].XIC[9].icell.Ien VGND.t1962 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X64 VPWR.t828 XThR.Tn[2].t13 XA.XIR[3].XIC[3].icell.PUM VPWR.t827 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X65 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout VGND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X66 VPWR.t1257 XThR.Tn[6].t15 XA.XIR[7].XIC[3].icell.PUM VPWR.t1256 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X67 VPWR.t1712 VPWR.t1710 XA.XIR[2].XIC_15.icell.PUM VPWR.t1711 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X68 a_6243_9615# XThC.XTB7.Y VPWR.t918 VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X69 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11].t12 XA.XIR[11].XIC[14].icell.Ien VGND.t1907 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X70 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11].t13 XA.XIR[11].XIC[8].icell.Ien VGND.t1908 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X71 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[3].t16 VGND.t2229 VGND.t2228 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X72 XThR.Tn[7].t7 XThR.XTBN.Y.t7 VPWR.t312 VPWR.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[0].t12 VGND.t2165 VGND.t2164 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X74 a_8963_9569# XThC.XTBN.Y.t10 VGND.t489 VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X75 VGND.t2394 Vbias.t8 XA.XIR[12].XIC[7].icell.SM VGND.t2393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X76 VGND.t569 XThC.Tn[6].t12 XA.XIR[12].XIC[6].icell.PDM VGND.t568 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X77 XA.XIR[6].XIC[9].icell.SM XA.XIR[6].XIC[9].icell.Ien Iout.t128 VGND.t1166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X78 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout VGND.t1181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X79 XA.XIR[3].XIC[11].icell.SM XA.XIR[3].XIC[11].icell.Ien Iout.t113 VGND.t1105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X80 VGND.t1661 VPWR.t1930 XA.XIR[4].XIC_dummy_left.icell.PDM VGND.t1660 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X81 VGND.t452 XThR.XTBN.Y.t8 XThR.Tn[5].t7 VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 VGND.t2396 Vbias.t9 XA.XIR[15].XIC[8].icell.SM VGND.t2395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X83 VGND.t2398 Vbias.t10 XA.XIR[14].XIC[9].icell.SM VGND.t2397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X84 VGND.t147 XThC.Tn[7].t8 XA.XIR[15].XIC[7].icell.PDM VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X85 VGND.t2435 XThC.Tn[11].t13 XA.XIR[6].XIC[11].icell.PDM VGND.t2434 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X86 VGND.t1409 XThC.Tn[1].t13 XA.XIR[3].XIC[1].icell.PDM VGND.t1408 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X87 XA.XIR[4].XIC[11].icell.Ien XThR.Tn[4].t13 VPWR.t721 VPWR.t720 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X88 VPWR.t129 XThR.XTB6.Y a_n1049_5611# VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X89 XA.XIR[14].XIC[6].icell.PUM XThC.Tn[6].t13 XA.XIR[14].XIC[6].icell.Ien VPWR.t418 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X90 VGND.t2400 Vbias.t11 XA.XIR[9].XIC[7].icell.SM VGND.t2399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X91 VGND.t2687 XThC.Tn[2].t13 XA.XIR[6].XIC[2].icell.PDM VGND.t2686 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X92 XA.XIR[11].XIC[9].icell.Ien XThR.Tn[11].t14 VPWR.t1079 VPWR.t1078 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X93 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t1931 XA.XIR[6].XIC_dummy_left.icell.Ien VGND.t1662 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X94 VGND.t1457 Vbias.t1 Vbias.t2 VGND.t1456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X95 a_n1049_7787# XThR.XTB2.Y VPWR.t932 VPWR.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X96 VGND.t23 XThC.Tn[9].t13 XA.XIR[14].XIC[9].icell.PDM VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X97 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8].t12 XA.XIR[8].XIC[11].icell.Ien VGND.t1224 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X98 VGND.t2402 Vbias.t12 XA.XIR[2].XIC[0].icell.SM VGND.t2401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X99 XA.XIR[1].XIC[1].icell.Ien XThR.Tn[1].t14 VPWR.t1140 VPWR.t1139 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X100 XA.XIR[13].XIC[4].icell.PUM XThC.Tn[4].t13 XA.XIR[13].XIC[4].icell.Ien VPWR.t1848 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X101 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1708 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1709 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X102 VGND.t2404 Vbias.t13 XA.XIR[0].XIC[13].icell.SM VGND.t2403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X103 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[0].t13 VGND.t2167 VGND.t2166 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X104 XA.XIR[4].XIC[2].icell.Ien XThR.Tn[4].t14 VPWR.t723 VPWR.t722 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X105 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[8].t13 VGND.t1226 VGND.t1225 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X106 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[8].t14 VGND.t1228 VGND.t1227 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X107 XA.XIR[3].XIC[3].icell.Ien XThR.Tn[3].t17 VPWR.t1337 VPWR.t1336 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X108 VGND.t2501 XThC.Tn[12].t12 XA.XIR[0].XIC[12].icell.PDM VGND.t2500 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X109 VPWR.t1768 XThC.XTB3.Y.t3 a_4067_9615# VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[1].t15 XA.XIR[1].XIC[4].icell.Ien VGND.t1963 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X111 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5].t12 XA.XIR[5].XIC[1].icell.Ien VGND.t2052 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X112 VPWR.t134 data[4].t0 a_n1335_4229# VPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X113 XA.XIR[2].XIC_15.icell.Ien XThR.Tn[2].t14 VPWR.t826 VPWR.t825 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X114 XA.XIR[3].XIC[9].icell.SM XA.XIR[3].XIC[9].icell.Ien Iout.t182 VGND.t1521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X115 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9].t14 XA.XIR[9].XIC[1].icell.Ien VGND.t788 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X116 VGND.t454 XThR.XTBN.Y.t9 XThR.Tn[7].t3 VGND.t453 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X117 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[4].t15 XA.XIR[4].XIC[5].icell.Ien VGND.t166 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X118 a_n1319_5317# XThR.XTB7.A VPWR.t836 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X119 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8].t15 XA.XIR[8].XIC[2].icell.Ien VGND.t1110 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X120 VPWR.t36 XThR.Tn[13].t12 XA.XIR[14].XIC[14].icell.PUM VPWR.t35 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X121 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11].t15 XA.XIR[11].XIC[3].icell.Ien VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X122 XA.XIR[7].XIC[8].icell.PUM XThC.Tn[8].t12 XA.XIR[7].XIC[8].icell.Ien VPWR.t1167 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X123 XThC.Tn[9].t7 XThC.XTB2.Y VPWR.t56 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X124 XA.XIR[15].XIC[4].icell.Ien VPWR.t1705 VPWR.t1707 VPWR.t1706 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X125 VGND.t2406 Vbias.t14 XA.XIR[12].XIC[2].icell.SM VGND.t2405 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X126 XA.XIR[6].XIC[4].icell.SM XA.XIR[6].XIC[4].icell.Ien Iout.t69 VGND.t646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X127 VGND.t2408 Vbias.t15 XA.XIR[11].XIC_15.icell.SM VGND.t2407 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X128 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1702 VPWR.t1704 VPWR.t1703 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X129 XThC.Tn[5].t10 XThC.XTBN.Y.t11 VGND.t490 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X130 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout VGND.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X131 VGND.t2410 Vbias.t16 XA.XIR[15].XIC[3].icell.SM VGND.t2409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X132 VGND.t270 Vbias.t17 XA.XIR[14].XIC[4].icell.SM VGND.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X133 VGND.t571 XThC.Tn[6].t14 XA.XIR[6].XIC[6].icell.PDM VGND.t570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X134 VPWR.t727 XThR.Tn[8].t16 XA.XIR[9].XIC[4].icell.PUM VPWR.t726 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X135 VPWR.t964 XThR.Tn[12].t15 XA.XIR[13].XIC[12].icell.PUM VPWR.t963 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X136 VGND.t1903 VGND.t1901 XA.XIR[13].XIC_dummy_right.icell.SM VGND.t1902 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X137 XThR.Tn[9].t3 XThR.XTB2.Y a_n997_3755# VGND.t1402 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X138 XThC.Tn[0].t2 XThC.XTBN.Y.t12 a_2979_9615# VPWR.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X139 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1932 VGND.t1664 VGND.t1663 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X140 XThC.Tn[5].t6 XThC.XTBN.Y.t13 a_5949_9615# VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X141 VGND.t566 XThC.XTB5.Y XThC.Tn[4].t2 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X142 XA.XIR[14].XIC[1].icell.PUM XThC.Tn[1].t14 XA.XIR[14].XIC[1].icell.Ien VPWR.t941 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X143 VGND.t272 Vbias.t18 XA.XIR[9].XIC[2].icell.SM VGND.t271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X144 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t3 VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X145 XA.XIR[13].XIC[0].icell.PUM XThC.Tn[0].t12 XA.XIR[13].XIC[0].icell.Ien VPWR.t1873 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X146 XThC.Tn[7].t3 XThC.XTBN.Y.t14 VGND.t492 VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X147 XThC.Tn[2].t7 XThC.XTBN.Y.t15 VGND.t493 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X148 VGND.t300 XThC.Tn[10].t13 XA.XIR[0].XIC[10].icell.PDM VGND.t299 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X149 a_n997_1579# XThR.XTBN.Y.t10 VGND.t456 VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X150 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[5].t13 VGND.t2054 VGND.t2053 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X151 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[5].t14 VGND.t2056 VGND.t2055 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X152 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1700 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1701 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X153 XA.XIR[9].XIC[14].icell.SM XA.XIR[9].XIC[14].icell.Ien Iout.t170 VGND.t1485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X154 VGND.t2477 XThC.Tn[4].t14 XA.XIR[14].XIC[4].icell.PDM VGND.t2476 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X155 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8].t17 XA.XIR[8].XIC[6].icell.Ien VGND.t1111 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X156 XA.XIR[1].XIC[7].icell.PUM XThC.Tn[7].t9 XA.XIR[1].XIC[7].icell.Ien VPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X157 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[6].t16 VGND.t2124 VGND.t2123 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X158 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[1].t16 VGND.t1965 VGND.t1964 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X159 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11].t16 XA.XIR[11].XIC[7].icell.Ien VGND.t1334 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X160 XA.XIR[4].XIC[8].icell.PUM XThC.Tn[8].t13 XA.XIR[4].XIC[8].icell.Ien VPWR.t1168 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X161 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[8].t18 VGND.t1113 VGND.t1112 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X162 XA.XIR[0].XIC_15.icell.SM XA.XIR[0].XIC_15.icell.Ien Iout.t48 VGND.t370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X163 XA.XIR[4].XIC[12].icell.SM XA.XIR[4].XIC[12].icell.Ien Iout.t247 VGND.t2502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X164 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[13].t13 VGND.t41 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X165 XA.XIR[11].XIC[12].icell.PUM XThC.Tn[12].t13 XA.XIR[11].XIC[12].icell.Ien VPWR.t1856 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X166 XA.XIR[12].XIC[4].icell.Ien XThR.Tn[12].t16 VPWR.t966 VPWR.t965 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X167 XA.XIR[3].XIC[4].icell.SM XA.XIR[3].XIC[4].icell.Ien Iout.t137 VGND.t1193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X168 XA.XIR[15].XIC[0].icell.Ien VPWR.t1697 VPWR.t1699 VPWR.t1698 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X169 VGND.t274 Vbias.t19 XA.XIR[8].XIC_15.icell.SM VGND.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X170 VGND.t129 XThC.Tn[14].t13 XA.XIR[8].XIC[14].icell.PDM VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X171 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1694 VPWR.t1696 VPWR.t1695 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X172 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[4].t16 XA.XIR[4].XIC[0].icell.Ien VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X173 VGND.t2045 XThC.Tn[8].t14 XA.XIR[8].XIC[8].icell.PDM VGND.t2044 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X174 XA.XIR[14].XIC[14].icell.Ien XThR.Tn[14].t13 VPWR.t164 VPWR.t163 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X175 VGND.t494 XThC.XTBN.Y.t16 XThC.Tn[1].t11 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X176 VGND.t276 Vbias.t20 XA.XIR[1].XIC[5].icell.SM VGND.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X177 VPWR.t968 XThR.Tn[12].t17 XA.XIR[13].XIC[10].icell.PUM VPWR.t967 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X178 XA.XIR[7].XIC[3].icell.PUM XThC.Tn[3].t13 XA.XIR[7].XIC[3].icell.Ien VPWR.t1266 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X179 XA.XIR[2].XIC_15.icell.PUM VPWR.t1692 XA.XIR[2].XIC_15.icell.Ien VPWR.t1693 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X180 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[2].t15 XA.XIR[2].XIC[13].icell.Ien VGND.t1160 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X181 VPWR.t584 XThR.Tn[9].t15 XA.XIR[10].XIC[12].icell.PUM VPWR.t583 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X182 VPWR.t729 XThR.Tn[8].t19 XA.XIR[9].XIC[0].icell.PUM VPWR.t728 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X183 VGND.t278 Vbias.t21 XA.XIR[4].XIC[6].icell.SM VGND.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X184 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1933 VGND.t1666 VGND.t1665 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X185 VPWR.t1691 VPWR.t1689 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1690 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X186 VPWR.t333 XThC.XTBN.Y.t17 XThC.Tn[10].t0 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X187 VGND.t457 XThR.XTBN.Y.t11 XThR.Tn[3].t11 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X188 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[2].t16 VGND.t1159 VGND.t1158 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X189 XA.XIR[6].XIC[8].icell.Ien XThR.Tn[6].t17 VPWR.t1259 VPWR.t1258 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X190 XThR.Tn[0].t7 XThR.XTBN.Y.t12 a_n1049_8581# VPWR.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X191 XA.XIR[13].XIC[12].icell.Ien XThR.Tn[13].t14 VPWR.t38 VPWR.t37 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X192 XA.XIR[13].XIC[7].icell.SM XA.XIR[13].XIC[7].icell.Ien Iout.t114 VGND.t1106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X193 VPWR.t1077 VGND.t2688 XA.XIR[0].XIC[8].icell.PUM VPWR.t1076 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X194 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10].t13 XA.XIR[10].XIC[14].icell.Ien VGND.t1949 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X195 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10].t14 XA.XIR[10].XIC[8].icell.Ien VGND.t1950 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X196 XThC.Tn[12].t6 XThC.XTB5.Y VPWR.t416 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 XA.XIR[1].XIC[11].icell.PUM XThC.Tn[11].t14 XA.XIR[1].XIC[11].icell.Ien VPWR.t662 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X198 XThR.Tn[11].t11 XThR.XTBN.Y.t13 VPWR.t314 VPWR.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 XA.XIR[0].XIC[7].icell.Ien XThR.Tn[0].t14 VPWR.t1296 VPWR.t1295 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X200 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[2].t17 VGND.t1157 VGND.t1156 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X201 XA.XIR[8].XIC[9].icell.PUM XThC.Tn[9].t14 XA.XIR[8].XIC[9].icell.Ien VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X202 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[8].t20 VGND.t1115 VGND.t1114 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X203 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout VGND.t2079 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X204 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[5].t15 VGND.t751 VGND.t750 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X205 VGND.t910 XThC.Tn[11].t15 XA.XIR[5].XIC[11].icell.PDM VGND.t909 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X206 XA.XIR[11].XIC[10].icell.PUM XThC.Tn[10].t14 XA.XIR[11].XIC[10].icell.Ien VPWR.t167 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X207 XThR.Tn[2].t6 XThR.XTBN.Y.t14 VGND.t459 VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X208 VGND.t912 XThC.Tn[11].t16 XA.XIR[9].XIC[11].icell.PDM VGND.t911 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X209 VGND.t1900 VGND.t1898 XA.XIR[13].XIC_dummy_left.icell.SM VGND.t1899 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X210 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12].t18 VPWR.t970 VPWR.t969 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X211 XA.XIR[1].XIC[2].icell.PUM XThC.Tn[2].t14 XA.XIR[1].XIC[2].icell.Ien VPWR.t1925 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X212 VPWR.t315 XThR.XTBN.Y.t15 XThR.Tn[12].t11 VPWR.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X213 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[1].t17 VGND.t1967 VGND.t1966 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X214 XThC.XTB7.A data[0].t0 VPWR.t746 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X215 VPWR.t586 XThR.Tn[9].t16 XA.XIR[10].XIC[10].icell.PUM VPWR.t585 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X216 XA.XIR[4].XIC[3].icell.PUM XThC.Tn[3].t14 XA.XIR[4].XIC[3].icell.Ien VPWR.t1267 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X217 VGND.t280 Vbias.t22 XA.XIR[4].XIC[10].icell.SM VGND.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X218 XA.XIR[0].XIC[13].icell.PDM VGND.t1895 VGND.t1897 VGND.t1896 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X219 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[13].t15 VGND.t43 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X220 VGND.t1668 VPWR.t1934 XA.XIR[0].XIC_dummy_left.icell.PDM VGND.t1667 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X221 VGND.t1423 XThC.Tn[2].t15 XA.XIR[5].XIC[2].icell.PDM VGND.t1422 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X222 VGND.t282 Vbias.t23 XA.XIR[11].XIC[8].icell.SM VGND.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X223 XThC.Tn[9].t3 XThC.XTB2.Y a_7875_9569# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X224 VGND.t2374 XThC.Tn[5].t12 XA.XIR[1].XIC[5].icell.PDM VGND.t2373 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X225 XA.XIR[10].XIC[9].icell.Ien XThR.Tn[10].t15 VPWR.t1116 VPWR.t1115 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X226 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1935 VGND.t1670 VGND.t1669 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X227 VGND.t1425 XThC.Tn[2].t16 XA.XIR[9].XIC[2].icell.PDM VGND.t1424 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X228 VGND.t2136 XThC.Tn[3].t15 XA.XIR[8].XIC[3].icell.PDM VGND.t2135 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X229 VGND.t1672 VPWR.t1936 XA.XIR[3].XIC_15.icell.PDM VGND.t1671 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X230 a_n1319_5611# XThR.XTB6.A VPWR.t44 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X231 XA.XIR[13].XIC[10].icell.Ien XThR.Tn[13].t16 VPWR.t40 VPWR.t39 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X232 VGND.t460 XThR.XTBN.Y.t16 a_n997_3979# VGND.t360 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X233 XA.XIR[15].XIC_15.icell.SM XA.XIR[15].XIC_15.icell.Ien Iout.t174 VGND.t1490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X234 VPWR.t390 XThC.XTBN.Y.t18 XThC.Tn[14].t11 VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X235 VGND.t284 Vbias.t24 XA.XIR[1].XIC[0].icell.SM VGND.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X236 VPWR.t972 XThR.Tn[12].t19 XA.XIR[13].XIC[5].icell.PUM VPWR.t971 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X237 XA.XIR[12].XIC[4].icell.PUM XThC.Tn[4].t15 XA.XIR[12].XIC[4].icell.Ien VPWR.t1849 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X238 VGND.t286 Vbias.t25 XA.XIR[4].XIC[1].icell.SM VGND.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X239 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7].t8 XA.XIR[7].XIC[14].icell.Ien VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X240 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7].t9 XA.XIR[7].XIC[8].icell.Ien VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X241 XA.XIR[0].XIC[11].icell.Ien XThR.Tn[0].t15 VPWR.t1017 VPWR.t1016 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X242 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[2].t18 VGND.t1155 VGND.t1154 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X243 XA.XIR[6].XIC[3].icell.Ien XThR.Tn[6].t18 VPWR.t1261 VPWR.t1260 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X244 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14].t14 XA.XIR[14].XIC[12].icell.Ien VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X245 XA.XIR[11].XIC[6].icell.SM XA.XIR[11].XIC[6].icell.Ien Iout.t175 VGND.t1491 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X246 XA.XIR[1].XIC_15.icell.Ien XThR.Tn[1].t18 VPWR.t1893 VPWR.t1892 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X247 VGND.t288 Vbias.t26 XA.XIR[2].XIC[14].icell.SM VGND.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X248 VGND.t1567 XThC.Tn[13].t13 XA.XIR[2].XIC[13].icell.PDM VGND.t1566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X249 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[5].t16 VGND.t753 VGND.t752 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X250 VPWR.t476 XThR.XTB4.Y a_n1049_6699# VPWR.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X251 VGND.t1674 VPWR.t1937 XA.XIR[15].XIC_dummy_right.icell.PDM VGND.t1673 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X252 XA.XIR[13].XIC[2].icell.SM XA.XIR[13].XIC[2].icell.Ien Iout.t26 VGND.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X253 VPWR.t1075 VGND.t2689 XA.XIR[0].XIC[3].icell.PUM VPWR.t1074 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X254 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10].t16 XA.XIR[10].XIC[3].icell.Ien VGND.t1951 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X255 VPWR.t764 XThC.XTB6.Y a_5949_9615# VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X256 VPWR.t1095 XThR.XTB1.Y a_n1049_8581# VPWR.t1094 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X257 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5].t17 XA.XIR[5].XIC_15.icell.Ien VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X258 VPWR.t920 XThR.Tn[11].t17 XA.XIR[12].XIC[7].icell.PUM VPWR.t919 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X259 XA.XIR[0].XIC[2].icell.Ien XThR.Tn[0].t16 VPWR.t1019 VPWR.t1018 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X260 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9].t17 XA.XIR[9].XIC_15.icell.Ien VGND.t789 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X261 XA.XIR[0].XIC[8].icell.SM XA.XIR[0].XIC[8].icell.Ien Iout.t25 VGND.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X262 VGND.t290 Vbias.t27 XA.XIR[5].XIC[7].icell.SM VGND.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X263 XA.XIR[11].XIC[5].icell.PUM XThC.Tn[5].t13 XA.XIR[11].XIC[5].icell.Ien VPWR.t1773 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X264 VGND.t573 XThC.Tn[6].t15 XA.XIR[5].XIC[6].icell.PDM VGND.t572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X265 VGND.t1929 XThR.XTB7.B a_n1335_8107# VGND.t1923 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X266 VPWR.t66 XThR.Tn[7].t10 XA.XIR[8].XIC[4].icell.PUM VPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X267 XA.XIR[0].XIC[5].icell.PDM XThR.Tn[0].t17 XA.XIR[0].XIC[5].icell.Ien VGND.t1593 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X268 VPWR.t1688 VPWR.t1686 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1687 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X269 VGND.t575 XThC.Tn[6].t16 XA.XIR[9].XIC[6].icell.PDM VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X270 VGND.t292 Vbias.t28 XA.XIR[8].XIC[8].icell.SM VGND.t291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X271 XA.XIR[7].XIC[9].icell.Ien XThR.Tn[7].t11 VPWR.t68 VPWR.t67 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X272 XThC.XTB4.Y.t1 XThC.XTB7.B VPWR.t744 VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X273 VGND.t1894 VGND.t1892 XA.XIR[12].XIC_dummy_right.icell.SM VGND.t1893 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X274 VGND.t149 XThC.Tn[7].t10 XA.XIR[8].XIC[7].icell.PDM VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X275 VPWR.t1685 VPWR.t1683 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1684 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X276 XThR.Tn[2].t10 XThR.XTB3.Y VGND.t870 VGND.t652 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X277 VGND.t461 XThR.XTBN.Y.t17 a_n997_2891# VGND.t376 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X278 VPWR.t588 XThR.Tn[9].t18 XA.XIR[10].XIC[5].icell.PUM VPWR.t587 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X279 XA.XIR[5].XIC[5].icell.SM XA.XIR[5].XIC[5].icell.Ien Iout.t164 VGND.t1387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X280 VPWR.t756 XThR.XTB5.Y XThR.Tn[12].t7 VPWR.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X281 XA.XIR[12].XIC[0].icell.PUM XThC.Tn[0].t13 XA.XIR[12].XIC[0].icell.Ien VPWR.t1874 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X282 VGND.t2519 XThC.Tn[0].t14 XA.XIR[1].XIC[0].icell.PDM VGND.t2518 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X283 VGND.t816 Vbias.t29 XA.XIR[11].XIC[3].icell.SM VGND.t815 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X284 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14].t15 XA.XIR[14].XIC[10].icell.Ien VGND.t294 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X285 XA.XIR[11].XIC[10].icell.SM XA.XIR[11].XIC[10].icell.Ien Iout.t72 VGND.t662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X286 VGND.t463 XThR.XTBN.Y.t18 XThR.Tn[6].t11 VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X287 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[11].t18 VGND.t1336 VGND.t1335 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X288 VPWR.t316 XThR.XTBN.Y.t19 XThR.Tn[9].t10 VPWR.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X289 XA.XIR[8].XIC[6].icell.SM XA.XIR[8].XIC[6].icell.Ien Iout.t70 VGND.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X290 XA.XIR[13].XIC[5].icell.Ien XThR.Tn[13].t17 VPWR.t42 VPWR.t41 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X291 VGND.t1891 VGND.t1889 XA.XIR[9].XIC_dummy_right.icell.SM VGND.t1890 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X292 XA.XIR[14].XIC_15.icell.PUM VPWR.t1681 XA.XIR[14].XIC_15.icell.Ien VPWR.t1682 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X293 a_n997_715# XThR.XTBN.Y.t20 VGND.t465 VGND.t464 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X294 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10].t17 XA.XIR[10].XIC[7].icell.Ien VGND.t1952 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X295 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7].t12 XA.XIR[7].XIC[3].icell.Ien VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X296 XThC.Tn[1].t10 XThC.XTBN.Y.t19 VGND.t547 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X297 VPWR.t922 XThR.Tn[11].t19 XA.XIR[12].XIC[11].icell.PUM VPWR.t921 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X298 XA.XIR[6].XIC[4].icell.PUM XThC.Tn[4].t16 XA.XIR[6].XIC[4].icell.Ien VPWR.t1850 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X299 XThR.Tn[14].t7 XThR.XTB7.Y VPWR.t994 VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X300 XA.XIR[10].XIC[12].icell.PUM XThC.Tn[12].t14 XA.XIR[10].XIC[12].icell.Ien VPWR.t605 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X301 XA.XIR[2].XIC[5].icell.SM XA.XIR[2].XIC[5].icell.Ien Iout.t41 VGND.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X302 XA.XIR[11].XIC[1].icell.SM XA.XIR[11].XIC[1].icell.Ien Iout.t206 VGND.t2077 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X303 XA.XIR[7].XIC_15.icell.PDM VPWR.t1938 VGND.t1676 VGND.t1675 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X304 XA.XIR[6].XIC[13].icell.SM XA.XIR[6].XIC[13].icell.Ien Iout.t29 VGND.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X305 XA.XIR[13].XIC[13].icell.PUM XThC.Tn[13].t14 XA.XIR[13].XIC[13].icell.Ien VPWR.t975 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X306 VGND.t818 Vbias.t30 XA.XIR[15].XIC[12].icell.SM VGND.t817 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X307 VGND.t820 Vbias.t31 XA.XIR[14].XIC[13].icell.SM VGND.t819 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X308 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[2].t19 XA.XIR[2].XIC[1].icell.Ien VGND.t1153 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X309 VPWR.t70 XThR.Tn[7].t13 XA.XIR[8].XIC[0].icell.PUM VPWR.t69 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X310 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[1].t19 XA.XIR[1].XIC[13].icell.Ien VGND.t2650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X311 VPWR.t755 XThR.XTB5.Y a_n1049_6405# VPWR.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X312 VPWR.t924 XThR.Tn[11].t20 XA.XIR[12].XIC[2].icell.PUM VPWR.t923 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X313 XThR.XTB7.B data[6].t0 VPWR.t840 VPWR.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X314 XA.XIR[0].XIC[8].icell.PUM XThC.Tn[8].t15 XA.XIR[0].XIC[8].icell.Ien VPWR.t1169 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X315 VPWR.t1846 XThC.XTB4.Y.t3 a_4861_9615# VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X316 XA.XIR[0].XIC[3].icell.SM XA.XIR[0].XIC[3].icell.Ien Iout.t60 VGND.t558 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X317 VGND.t822 Vbias.t32 XA.XIR[5].XIC[2].icell.SM VGND.t821 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X318 XA.XIR[8].XIC[4].icell.Ien XThR.Tn[8].t21 VPWR.t731 VPWR.t730 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X319 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1678 VPWR.t1680 VPWR.t1679 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X320 VGND.t1401 XThR.XTB2.Y XThR.Tn[1].t3 VGND.t1400 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X321 XA.XIR[0].XIC[0].icell.PDM XThR.Tn[0].t18 XA.XIR[0].XIC[0].icell.Ien VGND.t1594 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X322 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[11].t21 VGND.t1338 VGND.t1337 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X323 XA.XIR[12].XIC[7].icell.SM XA.XIR[12].XIC[7].icell.Ien Iout.t34 VGND.t205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X324 XThR.XTB7.A data[4].t1 a_n1331_2891# VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X325 XA.XIR[8].XIC[10].icell.SM XA.XIR[8].XIC[10].icell.Ien Iout.t249 VGND.t2504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X326 VGND.t824 Vbias.t33 XA.XIR[8].XIC[3].icell.SM VGND.t823 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X327 XA.XIR[15].XIC[13].icell.Ien VPWR.t1675 VPWR.t1677 VPWR.t1676 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X328 XA.XIR[15].XIC[8].icell.SM XA.XIR[15].XIC[8].icell.Ien Iout.t107 VGND.t1074 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X329 VPWR.t554 XThR.Tn[5].t18 XA.XIR[6].XIC[12].icell.PUM VPWR.t553 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X330 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1939 XA.XIR[11].XIC_dummy_right.icell.Ien VGND.t1677 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X331 VPWR.t1895 XThR.Tn[8].t22 XA.XIR[9].XIC[13].icell.PUM VPWR.t1894 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X332 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7].t14 XA.XIR[7].XIC[7].icell.Ien VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X333 a_n1049_7787# XThR.XTBN.Y.t21 XThR.Tn[1].t7 VPWR.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X334 XA.XIR[5].XIC[0].icell.SM XA.XIR[5].XIC[0].icell.Ien Iout.t219 VGND.t2220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X335 XA.XIR[10].XIC[10].icell.PUM XThC.Tn[10].t15 XA.XIR[10].XIC[10].icell.Ien VPWR.t168 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X336 VGND.t549 XThC.XTBN.Y.t20 XThC.Tn[4].t11 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X337 XA.XIR[6].XIC[0].icell.PUM XThC.Tn[0].t15 XA.XIR[6].XIC[0].icell.Ien VPWR.t1875 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X338 XA.XIR[8].XIC[1].icell.SM XA.XIR[8].XIC[1].icell.Ien Iout.t71 VGND.t661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X339 XA.XIR[3].XIC[13].icell.SM XA.XIR[3].XIC[13].icell.Ien Iout.t198 VGND.t1938 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X340 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1673 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1674 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X341 VGND.t1888 VGND.t1886 XA.XIR[12].XIC_dummy_left.icell.SM VGND.t1887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X342 XThC.XTB5.A data[1].t0 a_7331_10587# VPWR.t1232 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X343 VGND.t331 data[1].t1 a_8739_10571# VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X344 XA.XIR[0].XIC[1].icell.PDM VGND.t1883 VGND.t1885 VGND.t1884 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X345 VPWR.t931 XThR.XTB2.Y XThR.Tn[9].t7 VPWR.t650 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X346 VGND.t2455 XThR.XTBN.Y.t22 XThR.Tn[7].t2 VGND.t2454 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X347 VGND.t1507 XThC.Tn[13].t15 XA.XIR[14].XIC[13].icell.PDM VGND.t1506 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X348 XA.XIR[2].XIC[0].icell.SM XA.XIR[2].XIC[0].icell.Ien Iout.t129 VGND.t1167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X349 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1940 XA.XIR[14].XIC_dummy_left.icell.Ien VGND.t1678 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X350 XThR.Tn[13].t11 XThR.XTBN.Y.t23 VPWR.t1830 VPWR.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X351 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[10].t18 VGND.t2464 VGND.t2463 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X352 XA.XIR[14].XIC_15.icell.SM XA.XIR[14].XIC_15.icell.Ien Iout.t142 VGND.t1209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X353 VGND.t826 Vbias.t34 XA.XIR[10].XIC[11].icell.SM VGND.t825 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X354 VGND.t1882 VGND.t1880 XA.XIR[9].XIC_dummy_left.icell.SM VGND.t1881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X355 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8].t23 VPWR.t1897 VPWR.t1896 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X356 VPWR.t824 XThR.Tn[2].t20 XA.XIR[3].XIC[9].icell.PUM VPWR.t823 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X357 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1670 VPWR.t1672 VPWR.t1671 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X358 XA.XIR[12].XIC[13].icell.Ien XThR.Tn[12].t20 VPWR.t974 VPWR.t973 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X359 VPWR.t1858 XThR.Tn[6].t19 XA.XIR[7].XIC[9].icell.PUM VPWR.t1857 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X360 XA.XIR[0].XIC[3].icell.PUM XThC.Tn[3].t16 XA.XIR[0].XIC[3].icell.Ien VPWR.t1268 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X361 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1667 VPWR.t1669 VPWR.t1668 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X362 VPWR.t556 XThR.Tn[5].t19 XA.XIR[6].XIC[10].icell.PUM VPWR.t555 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X363 VGND.t611 XThC.Tn[1].t15 XA.XIR[2].XIC[1].icell.PDM VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X364 VGND.t218 XThR.XTB6.Y XThR.Tn[5].t3 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X365 XA.XIR[13].XIC[6].icell.PUM XThC.Tn[6].t17 XA.XIR[13].XIC[6].icell.Ien VPWR.t419 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X366 XThR.Tn[9].t2 XThR.XTB2.Y a_n997_3755# VGND.t1399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X367 VGND.t828 Vbias.t35 XA.XIR[1].XIC[14].icell.SM VGND.t827 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X368 XThR.XTB6.Y XThR.XTB6.A VGND.t58 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X369 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t1941 VGND.t1680 VGND.t1679 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X370 XA.XIR[12].XIC[2].icell.SM XA.XIR[12].XIC[2].icell.Ien Iout.t4 VGND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X371 a_n997_1579# XThR.XTBN.Y.t24 VGND.t2456 VGND.t398 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X372 VGND.t25 XThC.Tn[9].t15 XA.XIR[13].XIC[9].icell.PDM VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X373 XA.XIR[15].XIC[3].icell.SM XA.XIR[15].XIC[3].icell.Ien Iout.t10 VGND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X374 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[3].t18 XA.XIR[3].XIC[14].icell.Ien VGND.t2230 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X375 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[3].t19 XA.XIR[3].XIC[8].icell.Ien VGND.t2231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X376 VPWR.t166 XThR.Tn[14].t16 XA.XIR[15].XIC[7].icell.PUM VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X377 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1665 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1666 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X378 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout VGND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X379 VPWR.t882 XThR.Tn[13].t18 XA.XIR[14].XIC[8].icell.PUM VPWR.t881 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X380 XA.XIR[10].XIC[5].icell.PUM XThC.Tn[5].t14 XA.XIR[10].XIC[5].icell.Ien VPWR.t1774 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X381 XA.XIR[15].XIC[6].icell.Ien VPWR.t1662 VPWR.t1664 VPWR.t1663 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X382 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t1942 VGND.t1682 VGND.t1681 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X383 VGND.t830 Vbias.t36 XA.XIR[10].XIC[9].icell.SM VGND.t829 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X384 VPWR.t536 XThR.Tn[12].t21 XA.XIR[13].XIC[14].icell.PUM VPWR.t535 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X385 VPWR.t1899 XThR.Tn[8].t24 XA.XIR[9].XIC[6].icell.PUM VPWR.t1898 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X386 XA.XIR[15].XIC[9].icell.PDM VPWR.t1943 XA.XIR[15].XIC[9].icell.Ien VGND.t1683 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X387 XA.XIR[3].XIC[9].icell.Ien XThR.Tn[3].t20 VPWR.t1339 VPWR.t1338 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X388 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[10].t19 VGND.t2466 VGND.t2465 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X389 XA.XIR[15].XIC[12].icell.PDM XThR.Tn[14].t17 VGND.t296 VGND.t295 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X390 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1944 VGND.t1685 VGND.t1684 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X391 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[13].t19 VGND.t1258 VGND.t1257 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X392 VPWR.t192 XThR.XTBN.A XThR.XTBN.Y.t3 VPWR.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X393 VPWR.t558 XThR.Tn[5].t20 XA.XIR[6].XIC[5].icell.PUM VPWR.t557 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X394 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[4].t17 XA.XIR[4].XIC[11].icell.Ien VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X395 XA.XIR[5].XIC[4].icell.PUM XThC.Tn[4].t17 XA.XIR[5].XIC[4].icell.Ien VPWR.t1851 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X396 VPWR.t868 XThR.Tn[14].t18 XA.XIR[15].XIC[11].icell.PUM VPWR.t867 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X397 XA.XIR[1].XIC[5].icell.SM XA.XIR[1].XIC[5].icell.Ien Iout.t96 VGND.t881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X398 XA.XIR[13].XIC[1].icell.PUM XThC.Tn[1].t16 XA.XIR[13].XIC[1].icell.Ien VPWR.t456 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X399 XA.XIR[9].XIC[4].icell.PUM XThC.Tn[4].t18 XA.XIR[9].XIC[4].icell.Ien VPWR.t670 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X400 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1660 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1661 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X401 a_3523_10575# XThC.XTB7.B VGND.t1139 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X402 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[4].t18 VGND.t170 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X403 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[4].t19 VGND.t172 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X404 XA.XIR[12].XIC[13].icell.PUM XThC.Tn[13].t16 XA.XIR[12].XIC[13].icell.Ien VPWR.t976 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X405 XA.XIR[4].XIC[6].icell.SM XA.XIR[4].XIC[6].icell.Ien Iout.t152 VGND.t1262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X406 XA.XIR[11].XIC[14].icell.PUM XThC.Tn[14].t14 XA.XIR[11].XIC[14].icell.Ien VPWR.t87 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X407 VPWR.t392 XThC.XTBN.Y.t21 XThC.Tn[13].t11 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[1].t20 XA.XIR[1].XIC[1].icell.Ien VGND.t2651 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X409 VGND.t832 Vbias.t37 XA.XIR[13].XIC[5].icell.SM VGND.t831 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X410 VGND.t927 XThC.Tn[4].t19 XA.XIR[13].XIC[4].icell.PDM VGND.t926 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X411 XA.XIR[12].XIC[6].icell.Ien XThR.Tn[12].t22 VPWR.t538 VPWR.t537 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X412 XThC.Tn[5].t3 XThC.XTB6.Y VGND.t1177 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 XThC.Tn[4].t1 XThC.XTB5.Y VGND.t565 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X414 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[4].t20 XA.XIR[4].XIC[2].icell.Ien VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X415 VGND.t1687 VPWR.t1945 XA.XIR[8].XIC_dummy_right.icell.PDM VGND.t1686 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X416 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[3].t21 XA.XIR[3].XIC[3].icell.Ien VGND.t980 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X417 XA.XIR[14].XIC[8].icell.Ien XThR.Tn[14].t19 VPWR.t870 VPWR.t869 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X418 VPWR.t872 XThR.Tn[14].t20 XA.XIR[15].XIC[2].icell.PUM VPWR.t871 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X419 XA.XIR[2].XIC_15.icell.PDM XThR.Tn[2].t21 XA.XIR[2].XIC_15.icell.Ien VGND.t2493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X420 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t3 VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X421 VPWR.t884 XThR.Tn[13].t20 XA.XIR[14].XIC[3].icell.PUM VPWR.t883 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X422 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12].t23 XA.XIR[12].XIC[9].icell.Ien VGND.t724 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X423 VPWR.t590 XThR.Tn[9].t19 XA.XIR[10].XIC[14].icell.PUM VPWR.t589 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X424 XA.XIR[15].XIC[1].icell.Ien VPWR.t1657 VPWR.t1659 VPWR.t1658 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X425 VGND.t834 Vbias.t38 XA.XIR[11].XIC[12].icell.SM VGND.t833 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X426 VGND.t836 Vbias.t39 XA.XIR[7].XIC_15.icell.SM VGND.t835 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X427 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1654 VPWR.t1656 VPWR.t1655 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X428 VGND.t131 XThC.Tn[14].t15 XA.XIR[7].XIC[14].icell.PDM VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X429 VGND.t739 XThC.Tn[8].t16 XA.XIR[7].XIC[8].icell.PDM VGND.t738 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X430 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t2 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X431 XThC.Tn[4].t10 XThC.XTBN.Y.t22 VGND.t550 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X432 VPWR.t1021 XThR.Tn[0].t19 XA.XIR[1].XIC[4].icell.PUM VPWR.t1020 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X433 a_n1049_5317# XThR.XTB7.Y VPWR.t993 VPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X434 XA.XIR[13].XIC[14].icell.Ien XThR.Tn[13].t21 VPWR.t886 VPWR.t885 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X435 XA.XIR[14].XIC[8].icell.SM XA.XIR[14].XIC[8].icell.Ien Iout.t6 VGND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X436 XA.XIR[15].XIC[10].icell.PDM XThR.Tn[14].t21 VGND.t1244 VGND.t1243 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X437 VGND.t838 Vbias.t40 XA.XIR[10].XIC[4].icell.SM VGND.t837 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X438 VGND.t1879 VGND.t1877 XA.XIR[5].XIC_dummy_right.icell.SM VGND.t1878 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X439 VPWR.t1901 XThR.Tn[8].t25 XA.XIR[9].XIC[1].icell.PUM VPWR.t1900 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X440 VPWR.t113 XThR.Tn[4].t21 XA.XIR[5].XIC[4].icell.PUM VPWR.t112 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X441 XThC.XTB6.Y XThC.XTB7.B VGND.t1138 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X442 VPWR.t1653 VPWR.t1651 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1652 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X443 XA.XIR[15].XIC[4].icell.PDM VPWR.t1946 XA.XIR[15].XIC[4].icell.Ien VGND.t1688 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X444 VPWR.t72 XThR.Tn[7].t15 XA.XIR[8].XIC[13].icell.PUM VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X445 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t1947 XA.XIR[10].XIC_dummy_right.icell.Ien VGND.t1689 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X446 a_6243_9615# XThC.XTBN.Y.t23 XThC.Tn[6].t7 VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X447 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout VGND.t942 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X448 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[1].t21 VGND.t2653 VGND.t2652 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X449 XA.XIR[5].XIC[0].icell.PUM XThC.Tn[0].t16 XA.XIR[5].XIC[0].icell.Ien VPWR.t1876 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X450 XA.XIR[4].XIC[10].icell.SM XA.XIR[4].XIC[10].icell.Ien Iout.t228 VGND.t2372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X451 XA.XIR[9].XIC[0].icell.PUM XThC.Tn[0].t17 XA.XIR[9].XIC[0].icell.Ien VPWR.t1877 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X452 XThC.Tn[13].t7 XThC.XTB6.Y VPWR.t763 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X453 XA.XIR[5].XIC[14].icell.SM XA.XIR[5].XIC[14].icell.Ien Iout.t8 VGND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X454 VGND.t552 XThC.XTBN.Y.t24 XThC.Tn[0].t7 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X455 XThR.Tn[3].t7 XThR.XTBN.Y.t25 a_n1049_6699# VPWR.t1831 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X456 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[4].t22 XA.XIR[4].XIC[6].icell.Ien VGND.t871 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X457 VGND.t613 XThC.Tn[1].t17 XA.XIR[14].XIC[1].icell.PDM VGND.t612 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X458 VGND.t659 XThR.XTB4.Y XThR.Tn[3].t3 VGND.t658 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X459 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[3].t22 XA.XIR[3].XIC[7].icell.Ien VGND.t981 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X460 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[1].t22 VGND.t2655 VGND.t2654 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X461 XA.XIR[7].XIC[9].icell.PUM XThC.Tn[9].t16 XA.XIR[7].XIC[9].icell.Ien VPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X462 XA.XIR[1].XIC[0].icell.SM XA.XIR[1].XIC[0].icell.Ien Iout.t11 VGND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X463 XA.XIR[3].XIC[12].icell.PUM XThC.Tn[12].t15 XA.XIR[3].XIC[12].icell.Ien VPWR.t606 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X464 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[4].t23 VGND.t873 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X465 XA.XIR[0].XIC[12].icell.SM XA.XIR[0].XIC[12].icell.Ien Iout.t67 VGND.t644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X466 XA.XIR[0].XIC_15.icell.PDM VPWR.t1948 VGND.t1691 VGND.t1690 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X467 XA.XIR[4].XIC[1].icell.SM XA.XIR[4].XIC[1].icell.Ien Iout.t153 VGND.t1266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X468 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[9].t20 VGND.t791 VGND.t790 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X469 VGND.t621 Vbias.t41 XA.XIR[13].XIC[0].icell.SM VGND.t620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X470 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12].t24 VPWR.t540 VPWR.t539 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X471 XA.XIR[6].XIC[13].icell.PUM XThC.Tn[13].t17 XA.XIR[6].XIC[13].icell.Ien VPWR.t977 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X472 VGND.t623 Vbias.t42 XA.XIR[8].XIC[12].icell.SM VGND.t622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X473 XA.XIR[2].XIC[14].icell.SM XA.XIR[2].XIC[14].icell.Ien Iout.t3 VGND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X474 XThR.Tn[11].t7 XThR.XTB4.Y VPWR.t474 VPWR.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X475 VGND.t741 XThC.Tn[8].t17 XA.XIR[4].XIC[8].icell.PDM VGND.t740 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X476 VGND.t133 XThC.Tn[14].t16 XA.XIR[4].XIC[14].icell.PDM VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X477 XThC.Tn[14].t3 XThC.XTB7.Y a_10915_9569# VGND.t1308 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X478 VPWR.t1023 XThR.Tn[0].t20 XA.XIR[1].XIC[0].icell.PUM VPWR.t1022 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X479 XA.XIR[14].XIC[3].icell.Ien XThR.Tn[14].t22 VPWR.t874 VPWR.t873 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X480 VGND.t802 XThC.Tn[12].t16 XA.XIR[11].XIC[12].icell.PDM VGND.t801 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X481 VPWR.t655 XThR.Tn[4].t24 XA.XIR[5].XIC[0].icell.PUM VPWR.t654 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X482 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12].t25 XA.XIR[12].XIC[4].icell.Ien VGND.t725 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X483 XA.XIR[12].XIC[6].icell.PUM XThC.Tn[6].t18 XA.XIR[12].XIC[6].icell.Ien VPWR.t420 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X484 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t1949 XA.XIR[7].XIC_dummy_right.icell.Ien VGND.t1692 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X485 VPWR.t1650 VPWR.t1648 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1649 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X486 XA.XIR[15].XIC[7].icell.PUM XThC.Tn[7].t11 XA.XIR[15].XIC[7].icell.Ien VPWR.t101 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X487 VGND.t2472 XThC.XTB4.Y.t4 XThC.Tn[3].t11 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X488 VPWR.t55 XThC.XTB2.Y XThC.Tn[9].t6 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X489 XA.XIR[5].XIC[12].icell.Ien XThR.Tn[5].t21 VPWR.t560 VPWR.t559 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X490 VGND.t2440 XThC.Tn[3].t17 XA.XIR[7].XIC[3].icell.PDM VGND.t2439 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X491 VGND.t625 Vbias.t43 XA.XIR[6].XIC[11].icell.SM VGND.t624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X492 VGND.t1694 VPWR.t1950 XA.XIR[2].XIC_15.icell.PDM VGND.t1693 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X493 VPWR.t754 XThR.XTB5.Y XThR.Tn[12].t6 VPWR.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 VGND.t27 XThC.Tn[9].t17 XA.XIR[12].XIC[9].icell.PDM VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X495 XA.XIR[14].XIC[3].icell.SM XA.XIR[14].XIC[3].icell.Ien Iout.t5 VGND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X496 XA.XIR[9].XIC[12].icell.Ien XThR.Tn[9].t21 VPWR.t592 VPWR.t591 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X497 XA.XIR[8].XIC[13].icell.Ien XThR.Tn[8].t26 VPWR.t1903 VPWR.t1902 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X498 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout VGND.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X499 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6].t20 XA.XIR[6].XIC[14].icell.Ien VGND.t2507 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X500 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6].t21 XA.XIR[6].XIC[8].icell.Ien VGND.t2508 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X501 VPWR.t992 XThR.XTB7.Y XThR.Tn[14].t6 VPWR.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X502 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[1].t23 VGND.t2657 VGND.t2656 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X503 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13].t22 XA.XIR[13].XIC[12].icell.Ien VGND.t1259 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X504 XA.XIR[4].XIC[9].icell.PUM XThC.Tn[9].t18 XA.XIR[4].XIC[9].icell.Ien VPWR.t29 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X505 XThR.Tn[8].t3 XThR.XTB1.Y a_n997_3979# VGND.t1402 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X506 XA.XIR[3].XIC[10].icell.PUM XThC.Tn[10].t16 XA.XIR[3].XIC[10].icell.Ien VPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X507 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[4].t25 VGND.t875 VGND.t874 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X508 VGND.t914 XThC.Tn[11].t17 XA.XIR[1].XIC[11].icell.PDM VGND.t913 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X509 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1951 VGND.t1696 VGND.t1695 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X510 VPWR.t74 XThR.Tn[7].t16 XA.XIR[8].XIC[6].icell.PUM VPWR.t73 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X511 VPWR.t269 data[2].t0 XThC.XTB7.B VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X512 VGND.t1876 VGND.t1874 XA.XIR[5].XIC_dummy_left.icell.SM VGND.t1875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X513 VPWR.t1838 XThR.Tn[10].t20 XA.XIR[11].XIC[7].icell.PUM VPWR.t1837 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X514 VGND.t302 XThC.Tn[10].t17 XA.XIR[11].XIC[10].icell.PDM VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X515 XThC.Tn[13].t2 XThC.XTB6.Y a_10051_9569# VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X516 XThR.Tn[4].t7 XThR.XTBN.Y.t26 a_n1049_6405# VPWR.t1831 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X517 XThR.XTB5.Y XThR.XTB7.B a_n1319_6405# VPWR.t1104 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X518 VGND.t627 Vbias.t44 XA.XIR[4].XIC[7].icell.SM VGND.t626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X519 XThC.Tn[8].t11 XThC.XTBN.Y.t25 VPWR.t394 VPWR.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X520 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[13].t23 VGND.t1261 VGND.t1260 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X521 XA.XIR[15].XIC[11].icell.PUM XThC.Tn[11].t18 XA.XIR[15].XIC[11].icell.Ien VPWR.t663 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X522 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[9].t22 VGND.t581 VGND.t580 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X523 a_n1335_4229# data[5].t0 XThR.XTB5.A VPWR.t1235 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X524 VGND.t1427 XThC.Tn[2].t17 XA.XIR[1].XIC[2].icell.PDM VGND.t1426 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X525 VGND.t629 Vbias.t45 XA.XIR[7].XIC[8].icell.SM VGND.t628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X526 XA.XIR[6].XIC[9].icell.Ien XThR.Tn[6].t22 VPWR.t1860 VPWR.t1859 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X527 XA.XIR[5].XIC[10].icell.Ien XThR.Tn[5].t22 VPWR.t562 VPWR.t561 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X528 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[12].t26 VGND.t727 VGND.t726 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X529 VGND.t151 XThC.Tn[7].t12 XA.XIR[7].XIC[7].icell.PDM VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X530 VGND.t631 Vbias.t46 XA.XIR[6].XIC[9].icell.SM VGND.t630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X531 VGND.t633 Vbias.t47 XA.XIR[3].XIC[11].icell.SM VGND.t632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X532 XThC.Tn[8].t2 XThC.XTB1.Y.t4 a_7651_9569# VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X533 XThC.Tn[13].t10 XThC.XTBN.Y.t26 VPWR.t395 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X534 VGND.t2442 XThC.Tn[3].t18 XA.XIR[4].XIC[3].icell.PDM VGND.t2441 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X535 XA.XIR[9].XIC[10].icell.Ien XThR.Tn[9].t23 VPWR.t426 VPWR.t425 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X536 XA.XIR[7].XIC_15.icell.SM XA.XIR[7].XIC_15.icell.Ien Iout.t233 VGND.t2436 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X537 XA.XIR[15].XIC[12].icell.SM XA.XIR[15].XIC[12].icell.Ien Iout.t234 VGND.t2437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X538 VPWR.t1073 VGND.t2690 XA.XIR[0].XIC[9].icell.PUM VPWR.t1072 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X539 VGND.t1176 XThC.XTB6.Y XThC.Tn[5].t2 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X540 XA.XIR[12].XIC[1].icell.PUM XThC.Tn[1].t18 XA.XIR[12].XIC[1].icell.Ien VPWR.t457 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X541 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1645 VPWR.t1647 VPWR.t1646 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X542 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[3].t23 VGND.t983 VGND.t982 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X543 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[3].t24 VGND.t985 VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X544 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13].t24 XA.XIR[13].XIC[10].icell.Ien VGND.t1263 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X545 XA.XIR[15].XIC[2].icell.PUM XThC.Tn[2].t18 XA.XIR[15].XIC[2].icell.Ien VPWR.t946 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X546 XA.XIR[6].XIC[6].icell.PUM XThC.Tn[6].t19 XA.XIR[6].XIC[6].icell.Ien VPWR.t421 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X547 XA.XIR[10].XIC[14].icell.PUM XThC.Tn[14].t17 XA.XIR[10].XIC[14].icell.Ien VPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X548 VGND.t635 Vbias.t48 XA.XIR[12].XIC[5].icell.SM VGND.t634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X549 VGND.t929 XThC.Tn[4].t20 XA.XIR[12].XIC[4].icell.PDM VGND.t928 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X550 a_n1049_5611# XThR.XTB6.Y VPWR.t127 VPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X551 XA.XIR[13].XIC_15.icell.PUM VPWR.t1643 XA.XIR[13].XIC_15.icell.Ien VPWR.t1644 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X552 XThR.Tn[10].t3 XThR.XTB3.Y a_n997_2891# VGND.t651 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X553 VGND.t637 Vbias.t49 XA.XIR[15].XIC[6].icell.SM VGND.t636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X554 XA.XIR[0].XIC[11].icell.PDM XThR.Tn[0].t21 XA.XIR[0].XIC[11].icell.Ien VGND.t1595 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X555 VGND.t2376 XThC.Tn[5].t15 XA.XIR[15].XIC[5].icell.PDM VGND.t2375 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X556 VGND.t29 XThC.Tn[9].t19 XA.XIR[6].XIC[9].icell.PDM VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X557 VPWR.t397 XThC.XTBN.Y.t27 XThC.Tn[7].t6 VPWR.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X558 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6].t23 XA.XIR[6].XIC[3].icell.Ien VGND.t2509 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X559 XA.XIR[1].XIC_15.icell.PDM XThR.Tn[1].t24 XA.XIR[1].XIC_15.icell.Ien VGND.t2658 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X560 VPWR.t1840 XThR.Tn[10].t21 XA.XIR[11].XIC[11].icell.PUM VPWR.t1839 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X561 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1641 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1642 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X562 VPWR.t930 XThR.XTB2.Y XThR.Tn[9].t6 VPWR.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X563 VPWR.t1071 VGND.t2691 Vbias.t5 VPWR.t668 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X564 XThC.Tn[6].t6 XThC.XTBN.Y.t28 a_6243_9615# VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X565 XA.XIR[3].XIC[5].icell.PUM XThC.Tn[5].t16 XA.XIR[3].XIC[5].icell.Ien VPWR.t1775 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X566 VGND.t639 Vbias.t50 XA.XIR[9].XIC[5].icell.SM VGND.t638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X567 XA.XIR[8].XIC[6].icell.Ien XThR.Tn[8].t27 VPWR.t1905 VPWR.t1904 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X568 VGND.t577 XThC.Tn[6].t20 XA.XIR[1].XIC[6].icell.PDM VGND.t576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X569 VPWR.t680 XThR.Tn[3].t25 XA.XIR[4].XIC[4].icell.PUM VPWR.t679 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X570 VPWR.t570 XThR.Tn[7].t17 XA.XIR[8].XIC[1].icell.PUM VPWR.t569 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X571 XA.XIR[0].XIC[2].icell.PDM XThR.Tn[0].t22 XA.XIR[0].XIC[2].icell.Ien VGND.t1278 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X572 XA.XIR[11].XIC[7].icell.Ien XThR.Tn[11].t22 VPWR.t1807 VPWR.t1806 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X573 VGND.t641 Vbias.t51 XA.XIR[3].XIC[9].icell.SM VGND.t640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X574 VGND.t153 XThC.Tn[7].t13 XA.XIR[4].XIC[7].icell.PDM VGND.t152 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X575 XA.XIR[15].XIC_15.icell.Ien VPWR.t1638 VPWR.t1640 VPWR.t1639 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X576 VPWR.t1842 XThR.Tn[10].t22 XA.XIR[11].XIC[2].icell.PUM VPWR.t1841 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X577 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout VGND.t2487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X578 VPWR.t564 XThR.Tn[5].t23 XA.XIR[6].XIC[14].icell.PUM VPWR.t563 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X579 a_n1049_7493# XThR.XTBN.Y.t27 XThR.Tn[2].t11 VPWR.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X580 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8].t28 XA.XIR[8].XIC[9].icell.Ien VGND.t2659 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X581 XThC.Tn[0].t6 XThC.XTBN.Y.t29 VGND.t553 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X582 VGND.t643 Vbias.t52 XA.XIR[4].XIC[2].icell.SM VGND.t642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X583 VPWR.t1637 VPWR.t1635 XA.XIR[9].XIC_15.icell.PUM VPWR.t1636 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X584 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[0].t23 VGND.t1280 VGND.t1279 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X585 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[0].t24 VGND.t1282 VGND.t1281 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X586 VGND.t1459 Vbias.t53 XA.XIR[7].XIC[3].icell.SM VGND.t1458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X587 a_4067_9615# XThC.XTBN.Y.t30 XThC.Tn[2].t4 VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X588 XThR.Tn[0].t3 XThR.XTB1.Y VGND.t1913 VGND.t1394 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X589 VGND.t2457 XThR.XTBN.Y.t28 XThR.Tn[5].t6 VGND.t404 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X590 XA.XIR[11].XIC[7].icell.SM XA.XIR[11].XIC[7].icell.Ien Iout.t123 VGND.t1129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X591 XA.XIR[5].XIC[5].icell.Ien XThR.Tn[5].t24 VPWR.t1171 VPWR.t1170 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X592 VGND.t1461 Vbias.t54 XA.XIR[6].XIC[4].icell.SM VGND.t1460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X593 XThR.Tn[14].t3 XThR.XTB7.Y a_n997_715# VGND.t1556 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X594 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[12].t27 VGND.t729 VGND.t728 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X595 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[7].t18 VGND.t772 VGND.t771 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X596 VGND.t1463 Vbias.t55 XA.XIR[15].XIC[10].icell.SM VGND.t1462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X597 XA.XIR[9].XIC[5].icell.Ien XThR.Tn[9].t24 VPWR.t428 VPWR.t427 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X598 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[10].t23 VGND.t2468 VGND.t2467 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X599 XA.XIR[10].XIC[11].icell.SM XA.XIR[10].XIC[11].icell.Ien Iout.t216 VGND.t2102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X600 VGND.t1698 VPWR.t1952 XA.XIR[11].XIC_dummy_left.icell.PDM VGND.t1697 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X601 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6].t24 XA.XIR[6].XIC[7].icell.Ien VGND.t2510 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X602 VGND.t2458 XThR.XTBN.Y.t29 XThR.Tn[4].t11 VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X603 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[3].t26 VGND.t987 VGND.t986 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X604 XA.XIR[6].XIC[1].icell.PUM XThC.Tn[1].t19 XA.XIR[6].XIC[1].icell.Ien VPWR.t458 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X605 VGND.t1700 VPWR.t1953 XA.XIR[14].XIC_15.icell.PDM VGND.t1699 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X606 a_8963_9569# XThC.XTB4.Y.t5 XThC.Tn[11].t10 VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X607 XA.XIR[5].XIC[13].icell.PUM XThC.Tn[13].t18 XA.XIR[5].XIC[13].icell.Ien VPWR.t978 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X608 VGND.t1465 Vbias.t56 XA.XIR[12].XIC[0].icell.SM VGND.t1464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X609 XA.XIR[1].XIC[14].icell.SM XA.XIR[1].XIC[14].icell.Ien Iout.t126 VGND.t1141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X610 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1633 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1634 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X611 XA.XIR[9].XIC[13].icell.PUM XThC.Tn[13].t19 XA.XIR[9].XIC[13].icell.Ien VPWR.t979 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X612 VGND.t1467 Vbias.t57 XA.XIR[15].XIC[1].icell.SM VGND.t1466 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X613 XA.XIR[0].XIC[6].icell.PDM XThR.Tn[0].t25 XA.XIR[0].XIC[6].icell.Ien VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X614 VGND.t931 XThC.Tn[4].t21 XA.XIR[6].XIC[4].icell.PDM VGND.t930 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X615 VGND.t2521 XThC.Tn[0].t18 XA.XIR[15].XIC[0].icell.PDM VGND.t2520 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X616 VGND.t1469 Vbias.t58 XA.XIR[10].XIC[13].icell.SM VGND.t1468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X617 XA.XIR[11].XIC[11].icell.Ien XThR.Tn[11].t23 VPWR.t1809 VPWR.t1808 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X618 VGND.t804 XThC.Tn[12].t17 XA.XIR[10].XIC[12].icell.PDM VGND.t803 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X619 VPWR.t682 XThR.Tn[3].t27 XA.XIR[4].XIC[0].icell.PUM VPWR.t681 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X620 VGND.t1471 Vbias.t59 XA.XIR[13].XIC[14].icell.SM VGND.t1470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X621 XA.XIR[12].XIC_15.icell.Ien XThR.Tn[12].t28 VPWR.t542 VPWR.t541 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X622 VGND.t554 XThC.XTBN.Y.t31 a_8739_9569# VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X623 VGND.t1509 XThC.Tn[13].t20 XA.XIR[13].XIC[13].icell.PDM VGND.t1508 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X624 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t1954 XA.XIR[13].XIC_dummy_left.icell.Ien VGND.t1701 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X625 VPWR.t669 bias[0].t0 Vbias.t3 VPWR.t668 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X626 VGND.t1473 Vbias.t60 XA.XIR[9].XIC[0].icell.SM VGND.t1472 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X627 XA.XIR[4].XIC[4].icell.Ien XThR.Tn[4].t26 VPWR.t657 VPWR.t656 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X628 XA.XIR[8].XIC[1].icell.Ien XThR.Tn[8].t29 VPWR.t1106 VPWR.t1105 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X629 VGND.t1475 Vbias.t61 XA.XIR[0].XIC_15.icell.SM VGND.t1474 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X630 VGND.t743 XThC.Tn[8].t18 XA.XIR[0].XIC[8].icell.PDM VGND.t742 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X631 VGND.t135 XThC.Tn[14].t18 XA.XIR[0].XIC[14].icell.PDM VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X632 XA.XIR[11].XIC[2].icell.Ien XThR.Tn[11].t24 VPWR.t1811 VPWR.t1810 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X633 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[7].t19 VGND.t774 VGND.t773 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X634 XA.XIR[8].XIC[7].icell.SM XA.XIR[8].XIC[7].icell.Ien Iout.t203 VGND.t1994 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X635 a_9827_9569# XThC.XTBN.Y.t32 VGND.t555 VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X636 VGND.t1477 Vbias.t62 XA.XIR[3].XIC[4].icell.SM VGND.t1476 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X637 XA.XIR[7].XIC[8].icell.SM XA.XIR[7].XIC[8].icell.Ien Iout.t207 VGND.t2078 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X638 VPWR.t256 XThR.Tn[1].t25 XA.XIR[2].XIC[12].icell.PUM VPWR.t255 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X639 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8].t30 XA.XIR[8].XIC[4].icell.Ien VGND.t1930 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X640 VPWR.t910 XThR.Tn[0].t26 XA.XIR[1].XIC[13].icell.PUM VPWR.t909 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X641 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t1955 XA.XIR[3].XIC_dummy_right.icell.Ien VGND.t1702 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X642 XA.XIR[10].XIC[9].icell.SM XA.XIR[10].XIC[9].icell.Ien Iout.t232 VGND.t2388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X643 VPWR.t659 XThR.Tn[4].t27 XA.XIR[5].XIC[13].icell.PUM VPWR.t658 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X644 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11].t25 XA.XIR[11].XIC[5].icell.Ien VGND.t2421 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X645 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[3].t28 VGND.t989 VGND.t988 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X646 VPWR.t1632 VPWR.t1630 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1631 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X647 XA.XIR[15].XIC[13].icell.PDM VPWR.t1956 XA.XIR[15].XIC[13].icell.Ien VGND.t1703 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X648 VGND.t1522 XThC.XTB1.Y.t5 XThC.Tn[0].t8 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[0].t27 VGND.t1285 VGND.t1284 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X650 XA.XIR[11].XIC[2].icell.SM XA.XIR[11].XIC[2].icell.Ien Iout.t83 VGND.t766 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X651 XThR.XTB7.A data[5].t1 VPWR.t1234 VPWR.t1233 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X652 VGND.t304 XThC.Tn[10].t18 XA.XIR[10].XIC[10].icell.PDM VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X653 VPWR.t544 XThR.Tn[12].t29 XA.XIR[13].XIC[8].icell.PUM VPWR.t543 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X654 VGND.t2084 XThC.XTBN.A XThC.XTBN.Y.t1 VGND.t2083 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X655 XA.XIR[0].XIC[9].icell.PUM XThC.Tn[9].t20 XA.XIR[0].XIC[9].icell.Ien VPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X656 VPWR.t1103 XThR.XTB7.B XThR.XTB1.Y VPWR.t1102 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X657 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t2 VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X658 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[2].t22 VGND.t2492 VGND.t2491 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X659 XA.XIR[4].XIC[0].icell.Ien XThR.Tn[4].t28 VPWR.t661 VPWR.t660 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X660 XA.XIR[14].XIC[12].icell.SM XA.XIR[14].XIC[12].icell.Ien Iout.t124 VGND.t1130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X661 XA.XIR[14].XIC_15.icell.PDM VPWR.t1957 VGND.t1705 VGND.t1704 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X662 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1627 VPWR.t1629 VPWR.t1628 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X663 XA.XIR[13].XIC[5].icell.SM XA.XIR[13].XIC[5].icell.Ien Iout.t82 VGND.t765 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X664 VPWR.t258 XThR.Tn[1].t26 XA.XIR[2].XIC[10].icell.PUM VPWR.t257 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X665 XA.XIR[5].XIC[6].icell.PUM XThC.Tn[6].t21 XA.XIR[5].XIC[6].icell.Ien VPWR.t422 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X666 XThC.Tn[7].t5 XThC.XTBN.Y.t33 VPWR.t934 VPWR.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X667 VGND.t1928 XThR.XTB7.B a_n1335_7243# VGND.t1927 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X668 XA.XIR[9].XIC[6].icell.PUM XThC.Tn[6].t22 XA.XIR[9].XIC[6].icell.Ien VPWR.t423 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X669 XA.XIR[8].XIC[7].icell.PUM XThC.Tn[7].t14 XA.XIR[8].XIC[7].icell.Ien VPWR.t565 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X670 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[0].t28 VGND.t1287 VGND.t1286 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X671 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1958 VGND.t1707 VGND.t1706 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X672 XA.XIR[12].XIC_15.icell.PUM VPWR.t1625 XA.XIR[12].XIC_15.icell.Ien VPWR.t1626 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X673 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[8].t31 VGND.t1932 VGND.t1931 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X674 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12].t30 XA.XIR[12].XIC[13].icell.Ien VGND.t730 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X675 VGND.t2444 XThC.Tn[3].t19 XA.XIR[0].XIC[3].icell.PDM VGND.t2443 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X676 XA.XIR[11].XIC[8].icell.PUM XThC.Tn[8].t19 XA.XIR[11].XIC[8].icell.Ien VPWR.t547 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X677 VGND.t31 XThC.Tn[9].t21 XA.XIR[5].XIC[9].icell.PDM VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X678 XA.XIR[8].XIC[2].icell.SM XA.XIR[8].XIC[2].icell.Ien Iout.t192 VGND.t1909 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X679 XA.XIR[2].XIC[12].icell.Ien XThR.Tn[2].t23 VPWR.t822 VPWR.t821 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X680 XA.XIR[7].XIC[3].icell.SM XA.XIR[7].XIC[3].icell.Ien Iout.t24 VGND.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X681 XThC.Tn[11].t11 XThC.XTB4.Y.t6 VPWR.t1847 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X682 VGND.t2170 XThC.Tn[9].t22 XA.XIR[9].XIC[9].icell.PDM VGND.t2169 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X683 XA.XIR[10].XIC[4].icell.SM XA.XIR[10].XIC[4].icell.Ien Iout.t85 VGND.t782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X684 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1622 VPWR.t1624 VPWR.t1623 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X685 a_n997_1803# XThR.XTBN.Y.t30 VGND.t2459 VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X686 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11].t26 XA.XIR[11].XIC[0].icell.Ien VGND.t2422 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X687 XThR.Tn[3].t6 XThR.XTBN.Y.t31 a_n1049_6699# VPWR.t1832 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X688 VPWR.t430 XThR.Tn[9].t25 XA.XIR[10].XIC[8].icell.PUM VPWR.t429 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X689 VGND.t2460 XThR.XTBN.Y.t32 XThR.Tn[3].t10 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X690 VGND.t1479 Vbias.t63 XA.XIR[11].XIC[6].icell.SM VGND.t1478 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X691 XA.XIR[10].XIC[7].icell.Ien XThR.Tn[10].t24 VPWR.t1844 VPWR.t1843 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X692 VGND.t2276 VPWR.t1959 XA.XIR[7].XIC_dummy_right.icell.PDM VGND.t2275 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X693 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1960 VGND.t2278 VGND.t2277 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X694 XThC.Tn[2].t3 XThC.XTBN.Y.t34 a_4067_9615# VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X695 VPWR.t898 XThR.Tn[0].t29 XA.XIR[1].XIC[6].icell.PUM VPWR.t897 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X696 XA.XIR[13].XIC[8].icell.Ien XThR.Tn[13].t25 VPWR.t888 VPWR.t887 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X697 VPWR.t400 XThR.Tn[4].t29 XA.XIR[5].XIC[6].icell.PUM VPWR.t399 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X698 VPWR.t546 XThR.Tn[12].t31 XA.XIR[13].XIC[3].icell.PUM VPWR.t545 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X699 XThR.Tn[11].t6 XThR.XTB4.Y VPWR.t472 VPWR.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X700 VPWR.t1621 VPWR.t1619 XA.XIR[8].XIC_15.icell.PUM VPWR.t1620 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X701 VPWR.t54 XThC.XTB2.Y a_3773_9615# VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X702 a_n1049_8581# XThR.XTB1.Y VPWR.t1093 VPWR.t1092 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X703 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1617 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1618 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X704 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[2].t24 VGND.t2490 VGND.t2489 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X705 XA.XIR[8].XIC[11].icell.PUM XThC.Tn[11].t19 XA.XIR[8].XIC[11].icell.Ien VPWR.t664 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X706 VGND.t1481 Vbias.t64 XA.XIR[0].XIC[8].icell.SM VGND.t1480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X707 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[10].t25 VGND.t2470 VGND.t2469 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X708 VGND.t756 XThC.Tn[7].t15 XA.XIR[0].XIC[7].icell.PDM VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X709 VGND.t1873 VGND.t1871 XA.XIR[4].XIC_dummy_right.icell.SM VGND.t1872 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X710 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[5].t25 VGND.t2047 VGND.t2046 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X711 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[9].t26 VGND.t583 VGND.t582 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X712 XA.XIR[9].XIC[11].icell.SM XA.XIR[9].XIC[11].icell.Ien Iout.t191 VGND.t1711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X713 XA.XIR[2].XIC[10].icell.Ien XThR.Tn[2].t25 VPWR.t808 VPWR.t807 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X714 XA.XIR[13].XIC[0].icell.SM XA.XIR[13].XIC[0].icell.Ien Iout.t33 VGND.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X715 VGND.t2280 VPWR.t1961 XA.XIR[10].XIC_dummy_left.icell.PDM VGND.t2279 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X716 VPWR.t82 XThC.XTB6.A a_5949_10571# VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X717 VPWR.t260 XThR.Tn[1].t27 XA.XIR[2].XIC[5].icell.PUM VPWR.t259 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X718 XA.XIR[1].XIC[4].icell.PUM XThC.Tn[4].t22 XA.XIR[1].XIC[4].icell.Ien VPWR.t671 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X719 XA.XIR[5].XIC[1].icell.PUM XThC.Tn[1].t20 XA.XIR[5].XIC[1].icell.Ien VPWR.t459 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X720 VGND.t869 XThR.XTB3.Y XThR.Tn[2].t9 VGND.t649 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X721 VPWR.t890 XThR.Tn[13].t26 XA.XIR[14].XIC[9].icell.PUM VPWR.t889 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X722 XA.XIR[9].XIC[1].icell.PUM XThC.Tn[1].t21 XA.XIR[9].XIC[1].icell.Ien VPWR.t460 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X723 XA.XIR[8].XIC[2].icell.PUM XThC.Tn[2].t19 XA.XIR[8].XIC[2].icell.Ien VPWR.t947 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X724 XA.XIR[3].XIC[14].icell.PUM XThC.Tn[14].t19 XA.XIR[3].XIC[14].icell.Ien VPWR.t89 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X725 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[8].t32 VGND.t1934 VGND.t1933 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X726 XA.XIR[0].XIC[6].icell.SM XA.XIR[0].XIC[6].icell.Ien Iout.t220 VGND.t2221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X727 XThC.XTBN.Y.t3 XThC.XTBN.A VPWR.t1201 VPWR.t1200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X728 VGND.t2021 Vbias.t65 XA.XIR[5].XIC[5].icell.SM VGND.t2020 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X729 XA.XIR[11].XIC[3].icell.PUM XThC.Tn[3].t20 XA.XIR[11].XIC[3].icell.Ien VPWR.t1820 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X730 VGND.t933 XThC.Tn[4].t23 XA.XIR[5].XIC[4].icell.PDM VGND.t932 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X731 VGND.t2023 Vbias.t66 XA.XIR[11].XIC[10].icell.SM VGND.t2022 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X732 XA.XIR[10].XIC[11].icell.Ien XThR.Tn[10].t26 VPWR.t1825 VPWR.t1824 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X733 XThR.Tn[8].t2 XThR.XTB1.Y a_n997_3979# VGND.t1399 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X734 XA.XIR[6].XIC_15.icell.PUM VPWR.t1615 XA.XIR[6].XIC_15.icell.Ien VPWR.t1616 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X735 VGND.t615 XThC.Tn[1].t22 XA.XIR[13].XIC[1].icell.PDM VGND.t614 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X736 VGND.t2025 Vbias.t67 XA.XIR[12].XIC[14].icell.SM VGND.t2024 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X737 VGND.t935 XThC.Tn[4].t24 XA.XIR[9].XIC[4].icell.PDM VGND.t934 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X738 VGND.t2027 Vbias.t68 XA.XIR[8].XIC[6].icell.SM VGND.t2026 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X739 XA.XIR[7].XIC[7].icell.Ien XThR.Tn[7].t20 VPWR.t572 VPWR.t571 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X740 VGND.t2282 VPWR.t1962 XA.XIR[4].XIC_dummy_right.icell.PDM VGND.t2281 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X741 VGND.t2378 XThC.Tn[5].t17 XA.XIR[8].XIC[5].icell.PDM VGND.t2377 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X742 VGND.t1511 XThC.Tn[13].t21 XA.XIR[12].XIC[13].icell.PDM VGND.t1510 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X743 VGND.t1403 XThC.XTBN.Y.t35 a_9827_9569# VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X744 XA.XIR[2].XIC[12].icell.PUM XThC.Tn[12].t18 XA.XIR[2].XIC[12].icell.Ien VPWR.t607 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X745 VPWR.t432 XThR.Tn[9].t27 XA.XIR[10].XIC[3].icell.PUM VPWR.t431 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X746 VPWR.t917 XThC.XTB7.Y XThC.Tn[14].t7 VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X747 XThR.Tn[4].t6 XThR.XTBN.Y.t33 a_n1049_6405# VPWR.t1832 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X748 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14].t23 XA.XIR[14].XIC[8].icell.Ien VGND.t1245 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X749 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14].t24 XA.XIR[14].XIC[14].icell.Ien VGND.t1246 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X750 VGND.t2029 Vbias.t69 XA.XIR[11].XIC[1].icell.SM VGND.t2028 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X751 XA.XIR[10].XIC[2].icell.Ien XThR.Tn[10].t27 VPWR.t1827 VPWR.t1826 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X752 VGND.t2031 Vbias.t70 XA.XIR[7].XIC[12].icell.SM VGND.t2030 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X753 VPWR.t470 XThR.XTB4.Y a_n1049_6699# VPWR.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X754 XA.XIR[5].XIC[14].icell.Ien XThR.Tn[5].t26 VPWR.t1173 VPWR.t1172 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X755 VGND.t2033 Vbias.t71 XA.XIR[6].XIC[13].icell.SM VGND.t2032 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X756 VPWR.t900 XThR.Tn[0].t30 XA.XIR[1].XIC[1].icell.PUM VPWR.t899 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X757 XA.XIR[13].XIC[3].icell.Ien XThR.Tn[13].t27 VPWR.t892 VPWR.t891 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X758 XA.XIR[9].XIC[14].icell.Ien XThR.Tn[9].t28 VPWR.t434 VPWR.t433 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X759 VGND.t2035 Vbias.t72 XA.XIR[9].XIC[14].icell.SM VGND.t2034 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X760 VPWR.t402 XThR.Tn[4].t30 XA.XIR[5].XIC[1].icell.PUM VPWR.t401 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X761 XA.XIR[9].XIC[9].icell.SM XA.XIR[9].XIC[9].icell.Ien Iout.t156 VGND.t1277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X762 XA.XIR[8].XIC_15.icell.Ien XThR.Tn[8].t33 VPWR.t1108 VPWR.t1107 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X763 XA.XIR[15].XIC[1].icell.PDM VPWR.t1963 XA.XIR[15].XIC[1].icell.Ien VGND.t2283 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X764 VPWR.t684 XThR.Tn[3].t29 XA.XIR[4].XIC[13].icell.PUM VPWR.t683 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X765 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10].t28 XA.XIR[10].XIC[5].icell.Ien VGND.t2449 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X766 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1964 XA.XIR[6].XIC_dummy_right.icell.Ien VGND.t2284 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X767 XA.XIR[0].XIC[4].icell.Ien XThR.Tn[0].t31 VPWR.t902 VPWR.t901 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X768 XA.XIR[1].XIC[0].icell.PUM XThC.Tn[0].t19 XA.XIR[1].XIC[0].icell.Ien VPWR.t1878 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X769 VGND.t2037 Vbias.t73 XA.XIR[0].XIC[3].icell.SM VGND.t2036 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X770 XA.XIR[4].XIC[7].icell.SM XA.XIR[4].XIC[7].icell.Ien Iout.t173 VGND.t1489 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X771 XA.XIR[0].XIC[10].icell.SM XA.XIR[0].XIC[10].icell.Ien Iout.t157 VGND.t1288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X772 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[5].t27 VGND.t2049 VGND.t2048 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X773 XA.XIR[2].XIC[5].icell.Ien XThR.Tn[2].t26 VPWR.t820 VPWR.t819 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X774 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout VGND.t800 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X775 VGND.t2039 Vbias.t74 XA.XIR[8].XIC[10].icell.SM VGND.t2038 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X776 VPWR.t1834 XThR.XTBN.Y.t34 XThR.Tn[8].t11 VPWR.t1833 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X777 XA.XIR[7].XIC[11].icell.Ien XThR.Tn[7].t21 VPWR.t574 VPWR.t573 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X778 XThR.Tn[10].t2 XThR.XTB3.Y a_n997_2891# VGND.t648 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X779 XA.XIR[14].XIC[9].icell.Ien XThR.Tn[14].t25 VPWR.t876 VPWR.t875 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X780 XA.XIR[2].XIC[10].icell.PUM XThC.Tn[10].t19 XA.XIR[2].XIC[10].icell.Ien VPWR.t170 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X781 XThC.XTB3.Y.t0 XThC.XTB7.B VPWR.t743 VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X782 XA.XIR[0].XIC[1].icell.SM XA.XIR[0].XIC[1].icell.Ien Iout.t241 VGND.t2482 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X783 VGND.t2041 Vbias.t75 XA.XIR[5].XIC[0].icell.SM VGND.t2040 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X784 VGND.t1870 VGND.t1868 XA.XIR[4].XIC_dummy_left.icell.SM VGND.t1869 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X785 VGND.t2043 Vbias.t76 XA.XIR[8].XIC[1].icell.SM VGND.t2042 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X786 VPWR.t80 XThC.XTB6.A XThC.XTB2.Y VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X787 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[11].t27 VGND.t2424 VGND.t2423 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X788 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[11].t28 VGND.t2426 VGND.t2425 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X789 XA.XIR[12].XIC[5].icell.SM XA.XIR[12].XIC[5].icell.Ien Iout.t242 VGND.t2483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X790 XA.XIR[7].XIC[2].icell.Ien XThR.Tn[7].t22 VPWR.t576 VPWR.t575 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X791 VGND.t1605 Vbias.t77 XA.XIR[3].XIC[13].icell.SM VGND.t1604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X792 VGND.t2523 XThC.Tn[0].t20 XA.XIR[8].XIC[0].icell.PDM VGND.t2522 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X793 VGND.t806 XThC.Tn[12].t19 XA.XIR[3].XIC[12].icell.PDM VGND.t805 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X794 XThR.XTB3.Y XThR.XTB7.A VPWR.t835 VPWR.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X795 XA.XIR[15].XIC[6].icell.SM XA.XIR[15].XIC[6].icell.Ien Iout.t32 VGND.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X796 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12].t32 XA.XIR[12].XIC[1].icell.Ien VGND.t731 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X797 VGND.t1513 XThC.Tn[13].t22 XA.XIR[6].XIC[13].icell.PDM VGND.t1512 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X798 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7].t23 XA.XIR[7].XIC[5].icell.Ien VGND.t775 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X799 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1965 VGND.t2286 VGND.t2285 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X800 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t2 VGND.t1555 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X801 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14].t26 XA.XIR[14].XIC[3].icell.Ien VGND.t1247 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X802 XA.XIR[10].XIC[8].icell.PUM XThC.Tn[8].t20 XA.XIR[10].XIC[8].icell.Ien VPWR.t548 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X803 XA.XIR[1].XIC[12].icell.Ien XThR.Tn[1].t28 VPWR.t262 VPWR.t261 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X804 VGND.t1607 Vbias.t78 XA.XIR[2].XIC[11].icell.SM VGND.t1606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X805 XA.XIR[6].XIC_15.icell.SM XA.XIR[6].XIC_15.icell.Ien Iout.t18 VGND.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X806 XA.XIR[0].XIC[0].icell.Ien XThR.Tn[0].t32 VPWR.t904 VPWR.t903 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X807 XThR.Tn[0].t11 XThR.XTBN.Y.t35 VGND.t2461 VGND.t442 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X808 VPWR.t753 XThR.XTB5.Y a_n1049_6405# VPWR.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X809 XA.XIR[4].XIC[13].icell.Ien XThR.Tn[4].t31 VPWR.t404 VPWR.t403 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X810 VGND.t1609 Vbias.t79 XA.XIR[14].XIC_15.icell.SM VGND.t1608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X811 XA.XIR[9].XIC[4].icell.SM XA.XIR[9].XIC[4].icell.Ien Iout.t100 VGND.t925 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X812 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10].t29 XA.XIR[10].XIC[0].icell.Ien VGND.t2450 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X813 XThC.Tn[10].t9 XThC.XTB3.Y.t4 VPWR.t1769 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X814 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5].t28 XA.XIR[5].XIC[12].icell.Ien VGND.t2050 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X815 VPWR.t1835 XThR.XTBN.Y.t36 XThR.Tn[10].t11 VPWR.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X816 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout VGND.t1295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X817 VPWR.t97 XThR.Tn[11].t29 XA.XIR[12].XIC[4].icell.PUM VPWR.t96 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X818 VPWR.t935 XThC.XTBN.Y.t36 XThC.Tn[13].t9 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X819 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9].t29 XA.XIR[9].XIC[12].icell.Ien VGND.t584 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X820 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8].t34 XA.XIR[8].XIC[13].icell.Ien VGND.t1935 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X821 a_3773_9615# XThC.XTB2.Y VPWR.t53 VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X822 XThC.Tn[5].t1 XThC.XTB6.Y VGND.t1175 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X823 XA.XIR[4].XIC[2].icell.SM XA.XIR[4].XIC[2].icell.Ien Iout.t202 VGND.t1942 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X824 XThC.Tn[2].t10 XThC.XTB3.Y.t5 VGND.t2266 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X825 VPWR.t686 XThR.Tn[3].t30 XA.XIR[4].XIC[6].icell.PUM VPWR.t685 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X826 VPWR.t818 XThR.Tn[2].t27 XA.XIR[3].XIC[7].icell.PUM VPWR.t817 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X827 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[12].t33 VGND.t733 VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X828 VGND.t306 XThC.Tn[10].t20 XA.XIR[3].XIC[10].icell.PDM VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X829 VPWR.t1862 XThR.Tn[6].t25 XA.XIR[7].XIC[7].icell.PUM VPWR.t1861 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X830 XA.XIR[15].XIC[10].icell.SM XA.XIR[15].XIC[10].icell.Ien Iout.t38 VGND.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X831 VPWR.t1175 XThR.Tn[5].t29 XA.XIR[6].XIC[8].icell.PUM VPWR.t1174 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X832 VGND.t2462 XThR.XTBN.Y.t37 a_n997_3755# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X833 XA.XIR[2].XIC[5].icell.PUM XThC.Tn[5].t18 XA.XIR[2].XIC[5].icell.Ien VPWR.t1776 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X834 VPWR.t982 XThC.XTB1.Y.t6 a_2979_9615# VPWR.t981 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X835 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[9].t30 VGND.t586 VGND.t585 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X836 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1966 VGND.t2288 VGND.t2287 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X837 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14].t27 XA.XIR[14].XIC[7].icell.Ien VGND.t1248 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X838 XA.XIR[1].XIC[10].icell.Ien XThR.Tn[1].t29 VPWR.t264 VPWR.t263 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X839 VGND.t1611 Vbias.t80 XA.XIR[2].XIC[9].icell.SM VGND.t1610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X840 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[12].t34 VGND.t735 VGND.t734 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X841 XA.XIR[12].XIC[0].icell.SM XA.XIR[12].XIC[0].icell.Ien Iout.t62 VGND.t560 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X842 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[11].t30 VGND.t139 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X843 XA.XIR[3].XIC_15.icell.SM XA.XIR[3].XIC_15.icell.Ien Iout.t78 VGND.t746 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X844 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout VGND.t466 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X845 XA.XIR[7].XIC[12].icell.SM XA.XIR[7].XIC[12].icell.Ien Iout.t118 VGND.t1124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X846 XA.XIR[14].XIC[12].icell.PUM XThC.Tn[12].t20 XA.XIR[14].XIC[12].icell.Ien VPWR.t608 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X847 XA.XIR[15].XIC[1].icell.SM XA.XIR[15].XIC[1].icell.Ien Iout.t224 VGND.t2225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X848 VGND.t916 XThC.Tn[11].t20 XA.XIR[15].XIC[11].icell.PDM VGND.t915 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X849 XA.XIR[11].XIC_15.icell.PDM VPWR.t1967 VGND.t2290 VGND.t2289 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X850 XA.XIR[10].XIC[13].icell.SM XA.XIR[10].XIC[13].icell.Ien Iout.t171 VGND.t1486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X851 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5].t30 XA.XIR[5].XIC[10].icell.Ien VGND.t2051 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X852 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7].t24 XA.XIR[7].XIC[0].icell.Ien VGND.t1142 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X853 XA.XIR[13].XIC[14].icell.SM XA.XIR[13].XIC[14].icell.Ien Iout.t7 VGND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X854 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9].t31 XA.XIR[9].XIC[10].icell.Ien VGND.t587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X855 XA.XIR[10].XIC[3].icell.PUM XThC.Tn[3].t21 XA.XIR[10].XIC[3].icell.Ien VPWR.t1821 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X856 a_5155_9615# XThC.XTB5.Y VPWR.t415 VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X857 XA.XIR[5].XIC_15.icell.PUM VPWR.t1613 XA.XIR[5].XIC_15.icell.Ien VPWR.t1614 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X858 VPWR.t99 XThR.Tn[11].t31 XA.XIR[12].XIC[0].icell.PUM VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X859 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[6].t26 VGND.t2512 VGND.t2511 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X860 a_n1049_7493# XThR.XTB3.Y VPWR.t653 VPWR.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X861 VGND.t617 XThC.Tn[1].t23 XA.XIR[12].XIC[1].icell.PDM VGND.t616 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X862 XA.XIR[9].XIC_15.icell.PUM VPWR.t1611 XA.XIR[9].XIC_15.icell.Ien VPWR.t1612 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X863 VGND.t1429 XThC.Tn[2].t20 XA.XIR[15].XIC[2].icell.PDM VGND.t1428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X864 VPWR.t816 XThR.Tn[2].t28 XA.XIR[3].XIC[11].icell.PUM VPWR.t815 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X865 VPWR.t1864 XThR.Tn[6].t27 XA.XIR[7].XIC[11].icell.PUM VPWR.t1863 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X866 VGND.t2292 VPWR.t1968 XA.XIR[13].XIC_15.icell.PDM VGND.t2291 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X867 XThC.Tn[8].t7 XThC.XTB1.Y.t7 VPWR.t984 VPWR.t983 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X868 Vbias.t0 bias[2].t0 VPWR.t194 VPWR.t193 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X869 XA.XIR[4].XIC[6].icell.Ien XThR.Tn[4].t32 VPWR.t406 VPWR.t405 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X870 XA.XIR[3].XIC[7].icell.Ien XThR.Tn[3].t31 VPWR.t688 VPWR.t687 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X871 VGND.t1165 XThR.XTB5.Y XThR.Tn[4].t3 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X872 a_5155_9615# XThC.XTBN.Y.t37 XThC.Tn[4].t7 VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X873 VGND.t2294 VPWR.t1969 XA.XIR[0].XIC_dummy_right.icell.PDM VGND.t2293 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X874 VPWR.t633 XThR.Tn[3].t32 XA.XIR[4].XIC[1].icell.PUM VPWR.t632 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X875 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[12].t35 VGND.t737 VGND.t736 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X876 VPWR.t814 XThR.Tn[2].t29 XA.XIR[3].XIC[2].icell.PUM VPWR.t813 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X877 XThR.XTB5.Y XThR.XTB5.A VGND.t1191 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X878 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[11].t32 VGND.t141 VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X879 VPWR.t1866 XThR.Tn[6].t28 XA.XIR[7].XIC[2].icell.PUM VPWR.t1865 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X880 VPWR.t266 XThR.Tn[1].t30 XA.XIR[2].XIC[14].icell.PUM VPWR.t265 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X881 VPWR.t1177 XThR.Tn[5].t31 XA.XIR[6].XIC[3].icell.PUM VPWR.t1176 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X882 XA.XIR[14].XIC[10].icell.PUM XThC.Tn[10].t21 XA.XIR[14].XIC[10].icell.Ien VPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X883 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout VGND.t1488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X884 VPWR.t1610 VPWR.t1608 XA.XIR[1].XIC_15.icell.PUM VPWR.t1609 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X885 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[4].t33 XA.XIR[4].XIC[9].icell.Ien VGND.t562 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X886 VPWR.t1607 VPWR.t1605 XA.XIR[5].XIC_15.icell.PUM VPWR.t1606 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X887 XA.XIR[15].XIC_15.icell.PDM VPWR.t1970 XA.XIR[15].XIC_15.icell.Ien VGND.t2295 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X888 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[6].t29 VGND.t2514 VGND.t2513 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X889 XA.XIR[1].XIC[5].icell.Ien XThR.Tn[1].t31 VPWR.t268 VPWR.t267 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X890 VGND.t1613 Vbias.t81 XA.XIR[2].XIC[4].icell.SM VGND.t1612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X891 XA.XIR[6].XIC[8].icell.SM XA.XIR[6].XIC[8].icell.Ien Iout.t172 VGND.t1487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X892 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[2].t30 VGND.t714 VGND.t713 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X893 VGND.t1615 Vbias.t82 XA.XIR[15].XIC[7].icell.SM VGND.t1614 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X894 VGND.t2297 VPWR.t1971 XA.XIR[3].XIC_dummy_left.icell.PDM VGND.t2296 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X895 VGND.t1617 Vbias.t83 XA.XIR[14].XIC[8].icell.SM VGND.t1616 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X896 VGND.t579 XThC.Tn[6].t23 XA.XIR[15].XIC[6].icell.PDM VGND.t578 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X897 VPWR.t1604 VPWR.t1602 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1603 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X898 XThC.Tn[14].t2 XThC.XTB7.Y a_10915_9569# VGND.t1307 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X899 XThC.XTB3.Y.t1 XThC.XTB7.A a_4387_10575# VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X900 a_n997_1803# XThR.XTBN.Y.t38 VGND.t399 VGND.t398 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X901 XA.XIR[1].XIC[13].icell.PUM XThC.Tn[13].t23 XA.XIR[1].XIC[13].icell.Ien VPWR.t980 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X902 XA.XIR[3].XIC[11].icell.Ien XThR.Tn[3].t33 VPWR.t635 VPWR.t634 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X903 XA.XIR[15].XIC[14].icell.PDM XThR.Tn[14].t28 VGND.t1250 VGND.t1249 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X904 a_3773_9615# XThC.XTBN.Y.t38 XThC.Tn[1].t7 VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X905 VGND.t2058 XThC.Tn[1].t24 XA.XIR[6].XIC[1].icell.PDM VGND.t2057 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X906 XA.XIR[14].XIC[6].icell.SM XA.XIR[14].XIC[6].icell.Ien Iout.t36 VGND.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X907 XA.XIR[15].XIC[8].icell.PDM XThR.Tn[14].t29 VGND.t1252 VGND.t1251 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X908 VGND.t1619 Vbias.t84 XA.XIR[5].XIC[14].icell.SM VGND.t1618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X909 VGND.t1515 XThC.Tn[13].t24 XA.XIR[5].XIC[13].icell.PDM VGND.t1514 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X910 VPWR.t552 XThC.XTB5.A XThC.XTB1.Y.t0 VPWR.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X911 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1972 XA.XIR[5].XIC_dummy_left.icell.Ien VGND.t2298 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X912 VGND.t1517 XThC.Tn[13].t25 XA.XIR[9].XIC[13].icell.PDM VGND.t1516 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X913 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t1973 XA.XIR[9].XIC_dummy_left.icell.Ien VGND.t2299 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X914 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[1].t32 VGND.t1184 VGND.t1183 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X915 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11].t33 XA.XIR[11].XIC[11].icell.Ien VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X916 VGND.t1621 Vbias.t85 XA.XIR[1].XIC[11].icell.SM VGND.t1620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X917 XA.XIR[4].XIC[1].icell.Ien XThR.Tn[4].t34 VPWR.t408 VPWR.t407 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X918 VGND.t1623 Vbias.t86 XA.XIR[0].XIC[12].icell.SM VGND.t1622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X919 XA.XIR[3].XIC[2].icell.Ien XThR.Tn[3].t34 VPWR.t637 VPWR.t636 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X920 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12].t36 XA.XIR[12].XIC_15.icell.Ien VGND.t2153 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X921 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1600 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1601 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X922 XA.XIR[2].XIC[14].icell.Ien XThR.Tn[2].t31 VPWR.t812 VPWR.t811 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X923 XA.XIR[3].XIC[8].icell.SM XA.XIR[3].XIC[8].icell.Ien Iout.t138 VGND.t1197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X924 VGND.t2267 XThC.XTB3.Y.t6 XThC.Tn[2].t11 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X925 XA.XIR[14].XIC[5].icell.PUM XThC.Tn[5].t19 XA.XIR[14].XIC[5].icell.Ien VPWR.t1777 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X926 a_8739_9569# XThC.XTB3.Y.t7 XThC.Tn[10].t10 VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X927 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8].t35 XA.XIR[8].XIC[1].icell.Ien VGND.t1936 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X928 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[4].t35 XA.XIR[4].XIC[4].icell.Ien VGND.t563 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X929 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[3].t35 XA.XIR[3].XIC[5].icell.Ien VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X930 a_n1319_6405# XThR.XTB5.A VPWR.t834 VPWR.t833 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X931 VPWR.t878 XThR.Tn[14].t30 XA.XIR[15].XIC[4].icell.PUM VPWR.t877 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X932 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11].t34 XA.XIR[11].XIC[2].icell.Ien VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X933 XA.XIR[7].XIC[7].icell.PUM XThC.Tn[7].t16 XA.XIR[7].XIC[7].icell.Ien VPWR.t566 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X934 VPWR.t1599 VPWR.t1597 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1598 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X935 XA.XIR[6].XIC[3].icell.SM XA.XIR[6].XIC[3].icell.Ien Iout.t103 VGND.t940 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X936 a_2979_9615# XThC.XTB1.Y.t8 VPWR.t986 VPWR.t985 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X937 XA.XIR[0].XIC[13].icell.Ien XThR.Tn[0].t33 VPWR.t906 VPWR.t905 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X938 VGND.t1625 Vbias.t87 XA.XIR[15].XIC[2].icell.SM VGND.t1624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X939 VGND.t1627 Vbias.t88 XA.XIR[14].XIC[3].icell.SM VGND.t1626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X940 XThR.Tn[12].t10 XThR.XTBN.Y.t39 VPWR.t271 VPWR.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X941 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout VGND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X942 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1594 VPWR.t1596 VPWR.t1595 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X943 XA.XIR[14].XIC[10].icell.SM XA.XIR[14].XIC[10].icell.Ien Iout.t111 VGND.t1103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X944 XThC.Tn[11].t4 XThC.XTBN.Y.t39 VPWR.t936 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X945 VGND.t239 data[4].t2 XThR.XTB5.A VGND.t238 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X946 XThR.XTBN.Y.t1 XThR.XTBN.A VGND.t329 VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X947 VGND.t2249 data[3].t0 XThC.XTBN.A VGND.t2248 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X948 VGND.t1016 Vbias.t89 XA.XIR[1].XIC[9].icell.SM VGND.t1015 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X949 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1974 VGND.t2301 VGND.t2300 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X950 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[8].t36 VGND.t707 VGND.t706 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X951 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t3 VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X952 XA.XIR[15].XIC[3].icell.PDM XThR.Tn[14].t31 VGND.t1254 VGND.t1253 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X953 XA.XIR[14].XIC[1].icell.SM XA.XIR[14].XIC[1].icell.Ien Iout.t179 VGND.t1518 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X954 XA.XIR[10].XIC_15.icell.PDM VPWR.t1975 VGND.t2303 VGND.t2302 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X955 XA.XIR[9].XIC[13].icell.SM XA.XIR[9].XIC[13].icell.Ien Iout.t195 VGND.t1916 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X956 a_n997_2667# XThR.XTBN.Y.t40 VGND.t400 VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X957 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1592 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1593 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X958 XA.XIR[12].XIC[14].icell.SM XA.XIR[12].XIC[14].icell.Ien Iout.t139 VGND.t1198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X959 XA.XIR[1].XIC[6].icell.PUM XThC.Tn[6].t24 XA.XIR[1].XIC[6].icell.Ien VPWR.t424 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X960 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[1].t33 VGND.t1186 VGND.t1185 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X961 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11].t35 XA.XIR[11].XIC[6].icell.Ien VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X962 XA.XIR[7].XIC[11].icell.PUM XThC.Tn[11].t21 XA.XIR[7].XIC[11].icell.Ien VPWR.t665 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X963 XA.XIR[4].XIC[7].icell.PUM XThC.Tn[7].t17 XA.XIR[4].XIC[7].icell.Ien VPWR.t567 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X964 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[4].t36 VGND.t693 VGND.t692 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X965 VPWR.t880 XThR.Tn[14].t32 XA.XIR[15].XIC[0].icell.PUM VPWR.t879 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X966 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[8].t37 VGND.t709 VGND.t708 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X967 XA.XIR[3].XIC[8].icell.PUM XThC.Tn[8].t21 XA.XIR[3].XIC[8].icell.Ien VPWR.t549 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X968 VGND.t2172 XThC.Tn[9].t23 XA.XIR[1].XIC[9].icell.PDM VGND.t2171 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X969 XA.XIR[3].XIC[3].icell.SM XA.XIR[3].XIC[3].icell.Ien Iout.t94 VGND.t879 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X970 XThC.Tn[4].t6 XThC.XTBN.Y.t40 a_5155_9615# VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X971 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[3].t36 XA.XIR[3].XIC[0].icell.Ien VGND.t855 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X972 VGND.t2305 VPWR.t1976 XA.XIR[12].XIC_15.icell.PDM VGND.t2304 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X973 VPWR.t1280 XThR.Tn[12].t37 XA.XIR[13].XIC[9].icell.PUM VPWR.t1279 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X974 VPWR.t273 XThR.XTBN.Y.t41 XThR.Tn[8].t10 VPWR.t272 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X975 VGND.t137 XThC.Tn[14].t20 XA.XIR[11].XIC[14].icell.PDM VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X976 VGND.t745 XThC.Tn[8].t22 XA.XIR[11].XIC[8].icell.PDM VGND.t744 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X977 XA.XIR[7].XIC[2].icell.PUM XThC.Tn[2].t21 XA.XIR[7].XIC[2].icell.Ien VPWR.t948 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X978 XA.XIR[2].XIC[14].icell.PUM XThC.Tn[14].t21 XA.XIR[2].XIC[14].icell.Ien VPWR.t304 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X979 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1589 VPWR.t1591 VPWR.t1590 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X980 a_7651_9569# XThC.XTB1.Y.t9 XThC.Tn[8].t1 VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X981 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[2].t32 XA.XIR[2].XIC[12].icell.Ien VGND.t2497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X982 VGND.t1018 Vbias.t90 XA.XIR[4].XIC[5].icell.SM VGND.t1017 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X983 VPWR.t414 XThC.XTB5.Y XThC.Tn[12].t5 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X984 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t1977 XA.XIR[14].XIC_dummy_right.icell.Ien VGND.t2306 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X985 VPWR.t1795 XThR.Tn[11].t36 XA.XIR[12].XIC[13].icell.PUM VPWR.t1794 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X986 VPWR.t1588 VPWR.t1586 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1587 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X987 VGND.t1020 Vbias.t91 XA.XIR[7].XIC[6].icell.SM VGND.t1019 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X988 XA.XIR[6].XIC[7].icell.Ien XThR.Tn[6].t30 VPWR.t1868 VPWR.t1867 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X989 XA.XIR[5].XIC[8].icell.Ien XThR.Tn[5].t32 VPWR.t1179 VPWR.t1178 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X990 VGND.t2380 XThC.Tn[5].t20 XA.XIR[7].XIC[5].icell.PDM VGND.t2379 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X991 VGND.t402 XThR.XTBN.Y.t42 XThR.Tn[1].t11 VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X992 XA.XIR[15].XIC[7].icell.PDM XThR.Tn[14].t33 VGND.t1256 VGND.t1255 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X993 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[5].t33 VGND.t1986 VGND.t1985 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X994 XA.XIR[9].XIC[8].icell.Ien XThR.Tn[9].t32 VPWR.t436 VPWR.t435 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X995 VPWR.t1070 VGND.t2692 XA.XIR[0].XIC[7].icell.PUM VPWR.t1069 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X996 VPWR.t1585 VPWR.t1583 XA.XIR[4].XIC_15.icell.PUM VPWR.t1584 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X997 XA.XIR[0].XIC[6].icell.Ien XThR.Tn[0].t34 VPWR.t908 VPWR.t907 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X998 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13].t28 XA.XIR[13].XIC[14].icell.Ien VGND.t1264 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X999 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13].t29 XA.XIR[13].XIC[8].icell.Ien VGND.t1265 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1000 VGND.t1022 Vbias.t92 XA.XIR[1].XIC[4].icell.SM VGND.t1021 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1001 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[2].t33 VGND.t2496 VGND.t2495 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1002 XThR.Tn[6].t2 XThR.XTB7.Y VGND.t1554 VGND.t1553 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1003 a_9827_9569# XThC.XTBN.Y.t41 VGND.t1404 VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1004 XA.XIR[4].XIC[11].icell.PUM XThC.Tn[11].t22 XA.XIR[4].XIC[11].icell.Ien VPWR.t666 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1005 XThR.Tn[9].t9 XThR.XTBN.Y.t43 VPWR.t275 VPWR.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1006 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[8].t38 VGND.t711 VGND.t710 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1007 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[5].t34 VGND.t1988 VGND.t1987 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1008 XA.XIR[11].XIC[9].icell.PUM XThC.Tn[9].t24 XA.XIR[11].XIC[9].icell.Ien VPWR.t1297 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1009 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout VGND.t557 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1010 XA.XIR[5].XIC[11].icell.SM XA.XIR[5].XIC[11].icell.Ien Iout.t199 VGND.t1939 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1011 XA.XIR[0].XIC[9].icell.PDM XThR.Tn[0].t35 XA.XIR[0].XIC[9].icell.Ien VGND.t1275 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1012 XThC.Tn[1].t6 XThC.XTBN.Y.t42 a_3773_9615# VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1013 VGND.t918 XThC.Tn[11].t23 XA.XIR[8].XIC[11].icell.PDM VGND.t917 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1014 XThR.Tn[0].t10 XThR.XTBN.Y.t44 VGND.t403 VGND.t356 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1015 XThC.Tn[13].t1 XThC.XTB6.Y a_10051_9569# VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1016 XA.XIR[1].XIC[1].icell.PUM XThC.Tn[1].t25 XA.XIR[1].XIC[1].icell.Ien VPWR.t1180 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1017 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[2].t34 XA.XIR[2].XIC[10].icell.Ien VGND.t2494 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1018 XA.XIR[4].XIC[2].icell.PUM XThC.Tn[2].t22 XA.XIR[4].XIC[2].icell.Ien VPWR.t949 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1019 VPWR.t277 XThR.XTBN.Y.t45 XThR.Tn[10].t10 VPWR.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1020 VPWR.t438 XThR.Tn[9].t33 XA.XIR[10].XIC[9].icell.PUM VPWR.t437 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1021 XA.XIR[3].XIC[3].icell.PUM XThC.Tn[3].t22 XA.XIR[3].XIC[3].icell.Ien VPWR.t1822 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1022 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[4].t37 VGND.t695 VGND.t694 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1023 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1580 VPWR.t1582 VPWR.t1581 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1024 XA.XIR[0].XIC[12].icell.PDM VGND.t1865 VGND.t1867 VGND.t1866 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1025 VGND.t937 XThC.Tn[4].t25 XA.XIR[1].XIC[4].icell.PDM VGND.t936 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1026 VGND.t2060 XThC.Tn[1].t26 XA.XIR[5].XIC[1].icell.PDM VGND.t2059 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1027 VGND.t1024 Vbias.t93 XA.XIR[11].XIC[7].icell.SM VGND.t1023 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1028 VGND.t1026 Vbias.t94 XA.XIR[7].XIC[10].icell.SM VGND.t1025 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1029 XA.XIR[6].XIC[11].icell.Ien XThR.Tn[6].t31 VPWR.t1870 VPWR.t1869 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1030 VPWR.t916 XThC.XTB7.Y a_6243_9615# VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1031 XA.XIR[2].XIC[11].icell.SM XA.XIR[2].XIC[11].icell.Ien Iout.t121 VGND.t1127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1032 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1978 VGND.t2308 VGND.t2307 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1033 VGND.t2062 XThC.Tn[1].t27 XA.XIR[9].XIC[1].icell.PDM VGND.t2061 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1034 VGND.t2382 XThC.Tn[5].t21 XA.XIR[4].XIC[5].icell.PDM VGND.t2381 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1035 XA.XIR[13].XIC[9].icell.Ien XThR.Tn[13].t30 VPWR.t21 VPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1036 VGND.t1431 XThC.Tn[2].t23 XA.XIR[8].XIC[2].icell.PDM VGND.t1430 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1037 VPWR.t1068 VGND.t2693 XA.XIR[0].XIC[11].icell.PUM VPWR.t1067 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1038 VGND.t2446 XThC.Tn[3].t23 XA.XIR[11].XIC[3].icell.PDM VGND.t2445 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1039 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10].t30 XA.XIR[10].XIC[11].icell.Ien VGND.t2451 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1040 VGND.t2310 VPWR.t1979 XA.XIR[6].XIC_15.icell.PDM VGND.t2309 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1041 VGND.t1405 XThC.XTBN.Y.t43 a_8963_9569# VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1042 VGND.t1028 Vbias.t95 XA.XIR[4].XIC[0].icell.SM VGND.t1027 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1043 XA.XIR[15].XIC[4].icell.PUM XThC.Tn[4].t26 XA.XIR[15].XIC[4].icell.Ien VPWR.t672 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1044 VPWR.t1091 XThR.XTB1.Y XThR.Tn[8].t7 VPWR.t1090 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1045 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1578 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1579 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1046 VGND.t1030 Vbias.t96 XA.XIR[7].XIC[1].icell.SM VGND.t1029 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1047 VGND.t1032 Vbias.t97 XA.XIR[2].XIC[13].icell.SM VGND.t1031 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1048 XA.XIR[6].XIC[2].icell.Ien XThR.Tn[6].t32 VPWR.t1872 VPWR.t1871 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1049 XA.XIR[11].XIC[5].icell.SM XA.XIR[11].XIC[5].icell.Ien Iout.t105 VGND.t943 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1050 VGND.t2525 XThC.Tn[0].t21 XA.XIR[7].XIC[0].icell.PDM VGND.t2524 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1051 XA.XIR[1].XIC[14].icell.Ien XThR.Tn[1].t34 VPWR.t766 VPWR.t765 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1052 XA.XIR[5].XIC[3].icell.Ien XThR.Tn[5].t35 VPWR.t1162 VPWR.t1161 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1053 VGND.t808 XThC.Tn[12].t21 XA.XIR[2].XIC[12].icell.PDM VGND.t807 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1054 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[5].t36 VGND.t1990 VGND.t1989 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1055 XThR.XTBN.A data[7].t0 VPWR.t739 VPWR.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1056 XA.XIR[9].XIC[3].icell.Ien XThR.Tn[9].t34 VPWR.t440 VPWR.t439 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1057 XA.XIR[4].XIC_15.icell.Ien XThR.Tn[4].t38 VPWR.t506 VPWR.t505 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1058 XA.XIR[5].XIC[9].icell.SM XA.XIR[5].XIC[9].icell.Ien Iout.t90 VGND.t866 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1059 a_6243_10571# XThC.XTB7.B XThC.XTB7.Y VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1060 VPWR.t1066 VGND.t2694 XA.XIR[0].XIC[2].icell.PUM VPWR.t1065 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1061 VPWR.t929 XThR.XTB2.Y a_n1049_7787# VPWR.t646 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1062 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10].t31 XA.XIR[10].XIC[2].icell.Ien VGND.t2452 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1063 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6].t33 XA.XIR[6].XIC[5].icell.Ien VGND.t2515 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1064 XA.XIR[0].XIC[1].icell.Ien XThR.Tn[0].t36 VPWR.t894 VPWR.t893 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1065 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13].t31 XA.XIR[13].XIC[3].icell.Ien VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1066 VPWR.t1797 XThR.Tn[11].t37 XA.XIR[12].XIC[6].icell.PUM VPWR.t1796 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1067 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8].t39 XA.XIR[8].XIC_15.icell.Ien VGND.t712 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1068 XA.XIR[0].XIC[7].icell.SM XA.XIR[0].XIC[7].icell.Ien Iout.t50 VGND.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1069 XA.XIR[0].XIC[10].icell.PDM VGND.t1862 VGND.t1864 VGND.t1863 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1070 XA.XIR[0].XIC[4].icell.PDM XThR.Tn[0].t37 XA.XIR[0].XIC[4].icell.Ien VGND.t1267 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1071 VGND.t1034 Vbias.t98 XA.XIR[8].XIC[7].icell.SM VGND.t1033 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1072 a_n1049_7493# XThR.XTBN.Y.t46 XThR.Tn[2].t4 VPWR.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1073 XA.XIR[2].XIC[9].icell.SM XA.XIR[2].XIC[9].icell.Ien Iout.t27 VGND.t165 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1074 VGND.t510 XThC.Tn[6].t25 XA.XIR[8].XIC[6].icell.PDM VGND.t509 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1075 XThC.Tn[8].t6 XThC.XTB1.Y.t10 VPWR.t1193 VPWR.t1192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1076 VPWR.t1829 XThR.Tn[10].t32 XA.XIR[11].XIC[4].icell.PUM VPWR.t1828 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1077 VPWR.t1577 VPWR.t1575 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1576 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1078 VGND.t1861 VGND.t1859 XA.XIR[15].XIC_dummy_right.icell.SM VGND.t1860 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1079 VGND.t758 XThC.Tn[7].t18 XA.XIR[11].XIC[7].icell.PDM VGND.t757 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1080 XThR.Tn[0].t2 XThR.XTB1.Y VGND.t1912 VGND.t1391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1081 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7].t25 XA.XIR[7].XIC[11].icell.Ien VGND.t1143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1082 VGND.t1036 Vbias.t99 XA.XIR[11].XIC[2].icell.SM VGND.t1035 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1083 XA.XIR[15].XIC[0].icell.PUM XThC.Tn[0].t22 XA.XIR[15].XIC[0].icell.Ien VPWR.t1879 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1084 VPWR.t651 XThR.XTB3.Y XThR.Tn[10].t7 VPWR.t650 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1085 VGND.t308 XThC.Tn[10].t22 XA.XIR[2].XIC[10].icell.PDM VGND.t307 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1086 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[7].t26 VGND.t1145 VGND.t1144 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1087 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[7].t27 VGND.t1147 VGND.t1146 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1088 XA.XIR[8].XIC[5].icell.SM XA.XIR[8].XIC[5].icell.Ien Iout.t143 VGND.t1210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1089 VPWR.t52 XThC.XTB2.Y a_3773_9615# VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1090 VGND.t2527 XThC.Tn[0].t23 XA.XIR[4].XIC[0].icell.PDM VGND.t2526 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1091 VGND.t405 XThR.XTBN.Y.t47 XThR.Tn[4].t10 VGND.t404 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1092 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1573 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1574 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1093 XA.XIR[7].XIC[6].icell.SM XA.XIR[7].XIC[6].icell.Ien Iout.t93 VGND.t878 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1094 XA.XIR[14].XIC[14].icell.PUM XThC.Tn[14].t22 XA.XIR[14].XIC[14].icell.Ien VPWR.t305 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1095 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10].t33 XA.XIR[10].XIC[6].icell.Ien VGND.t2453 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1096 VPWR.t937 XThC.XTBN.Y.t44 XThC.Tn[9].t11 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1097 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t1980 XA.XIR[2].XIC_dummy_left.icell.Ien VGND.t2311 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1098 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7].t28 XA.XIR[7].XIC[2].icell.Ien VGND.t1148 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1099 VGND.t1406 XThC.XTBN.Y.t45 XThC.Tn[5].t9 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1100 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[3].t37 VGND.t857 VGND.t856 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1101 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13].t32 XA.XIR[13].XIC[7].icell.Ien VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1102 XA.XIR[11].XIC[0].icell.SM XA.XIR[11].XIC[0].icell.Ien Iout.t254 VGND.t2660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1103 XA.XIR[6].XIC[12].icell.SM XA.XIR[6].XIC[12].icell.Ien Iout.t229 VGND.t2385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1104 VGND.t407 XThR.XTBN.Y.t48 a_n997_1579# VGND.t406 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1105 XA.XIR[13].XIC[12].icell.PUM XThC.Tn[12].t22 XA.XIR[13].XIC[12].icell.Ien VPWR.t609 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1106 XA.XIR[5].XIC[4].icell.SM XA.XIR[5].XIC[4].icell.Ien Iout.t236 VGND.t2471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1107 VGND.t1038 Vbias.t100 XA.XIR[14].XIC[12].icell.SM VGND.t1037 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1108 VGND.t992 Vbias.t101 XA.XIR[10].XIC_15.icell.SM VGND.t991 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1109 a_2979_9615# XThC.XTBN.Y.t46 XThC.Tn[0].t1 VPWR.t938 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1110 VGND.t445 XThC.Tn[14].t23 XA.XIR[10].XIC[14].icell.PDM VGND.t444 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1111 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6].t34 XA.XIR[6].XIC[0].icell.Ien VGND.t2516 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1112 VGND.t2203 XThC.Tn[8].t23 XA.XIR[10].XIC[8].icell.PDM VGND.t2202 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1113 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[1].t35 XA.XIR[1].XIC[12].icell.Ien VGND.t1187 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1114 VPWR.t1799 XThR.Tn[11].t38 XA.XIR[12].XIC[1].icell.PUM VPWR.t1798 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1115 XA.XIR[0].XIC[7].icell.PUM XThC.Tn[7].t19 XA.XIR[0].XIC[7].icell.Ien VPWR.t568 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1116 XThC.Tn[12].t2 XThC.XTB5.Y a_9827_9569# VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1117 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[4].t39 XA.XIR[4].XIC[13].icell.Ien VGND.t696 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1118 VPWR.t522 XThR.Tn[10].t34 XA.XIR[11].XIC[0].icell.PUM VPWR.t521 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1119 XThR.XTB6.A data[5].t2 VPWR.t1853 VPWR.t1852 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1120 XA.XIR[0].XIC[2].icell.SM XA.XIR[0].XIC[2].icell.Ien Iout.t166 VGND.t1389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1121 VPWR.t1572 VPWR.t1570 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1571 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1122 XThR.Tn[14].t1 XThR.XTB7.Y a_n997_715# VGND.t1552 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1123 VPWR.t1003 XThR.Tn[14].t34 XA.XIR[15].XIC[13].icell.PUM VPWR.t1002 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1124 a_n1049_5317# XThR.XTBN.Y.t49 XThR.Tn[6].t7 VPWR.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1125 XA.XIR[11].XIC[4].icell.Ien XThR.Tn[11].t39 VPWR.t1801 VPWR.t1800 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1126 VGND.t994 Vbias.t102 XA.XIR[8].XIC[2].icell.SM VGND.t993 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1127 XA.XIR[2].XIC[4].icell.SM XA.XIR[2].XIC[4].icell.Ien Iout.t201 VGND.t1941 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1128 XA.XIR[15].XIC[12].icell.Ien VPWR.t1567 VPWR.t1569 VPWR.t1568 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1129 XA.XIR[7].XIC[10].icell.SM XA.XIR[7].XIC[10].icell.Ien Iout.t162 VGND.t1294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1130 XA.XIR[15].XIC[7].icell.SM XA.XIR[15].XIC[7].icell.Ien Iout.t1 VGND.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1131 VPWR.t768 XThR.Tn[1].t36 XA.XIR[2].XIC[8].icell.PUM VPWR.t767 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1132 VPWR.t516 XThR.Tn[8].t40 XA.XIR[9].XIC[12].icell.PUM VPWR.t515 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1133 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7].t29 XA.XIR[7].XIC[6].icell.Ien VGND.t1149 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1134 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1981 VGND.t2313 VGND.t2312 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1135 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[0].t38 VGND.t1269 VGND.t1268 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1136 XA.XIR[10].XIC[9].icell.PUM XThC.Tn[9].t25 XA.XIR[10].XIC[9].icell.Ien VPWR.t1298 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1137 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[7].t30 VGND.t1151 VGND.t1150 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1138 XA.XIR[8].XIC[0].icell.SM XA.XIR[8].XIC[0].icell.Ien Iout.t150 VGND.t1241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1139 XA.XIR[3].XIC[12].icell.SM XA.XIR[3].XIC[12].icell.Ien Iout.t12 VGND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1140 XA.XIR[3].XIC_15.icell.PDM VPWR.t1982 VGND.t2315 VGND.t2314 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1141 XA.XIR[13].XIC[10].icell.PUM XThC.Tn[10].t23 XA.XIR[13].XIC[10].icell.Ien VPWR.t172 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1142 XA.XIR[7].XIC[1].icell.SM XA.XIR[7].XIC[1].icell.Ien Iout.t204 VGND.t1995 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1143 a_6243_9615# XThC.XTB7.Y VPWR.t915 VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1144 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1565 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1566 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1145 VGND.t1858 VGND.t1856 XA.XIR[15].XIC_dummy_left.icell.SM VGND.t1857 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1146 XThC.Tn[10].t4 XThC.XTBN.Y.t47 VPWR.t939 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1147 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[1].t37 XA.XIR[1].XIC[10].icell.Ien VGND.t1188 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1148 XA.XIR[0].XIC[11].icell.PUM XThC.Tn[11].t24 XA.XIR[0].XIC[11].icell.Ien VPWR.t667 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1149 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[3].t38 VGND.t859 VGND.t858 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1150 VGND.t810 XThC.Tn[12].t23 XA.XIR[14].XIC[12].icell.PDM VGND.t809 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1151 XA.XIR[1].XIC_15.icell.PUM VPWR.t1563 XA.XIR[1].XIC_15.icell.Ien VPWR.t1564 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1152 XThC.Tn[10].t11 XThC.XTB3.Y.t8 a_8739_9569# VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1153 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[1].t38 VGND.t1190 VGND.t1189 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1154 VGND.t1306 XThC.XTB7.Y XThC.Tn[6].t3 VGND.t1305 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1155 XA.XIR[1].XIC[11].icell.SM XA.XIR[1].XIC[11].icell.Ien Iout.t73 VGND.t663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1156 VGND.t2317 VPWR.t1983 XA.XIR[2].XIC_dummy_left.icell.PDM VGND.t2316 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1157 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1984 VGND.t2319 VGND.t2318 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1158 XThR.Tn[11].t10 XThR.XTBN.Y.t50 VPWR.t280 VPWR.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1159 VGND.t2448 XThC.Tn[3].t24 XA.XIR[10].XIC[3].icell.PDM VGND.t2447 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1160 VPWR.t952 XThC.XTBN.Y.t48 XThC.Tn[12].t11 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1161 VGND.t2321 VPWR.t1985 XA.XIR[5].XIC_15.icell.PDM VGND.t2320 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1162 XA.XIR[15].XIC[10].icell.Ien VPWR.t1560 VPWR.t1562 VPWR.t1561 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1163 VGND.t996 Vbias.t103 XA.XIR[13].XIC[11].icell.SM VGND.t995 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1164 XA.XIR[12].XIC[12].icell.Ien XThR.Tn[12].t38 VPWR.t1282 VPWR.t1281 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1165 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11].t40 VPWR.t1803 VPWR.t1802 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1166 VGND.t2323 VPWR.t1986 XA.XIR[9].XIC_15.icell.PDM VGND.t2322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1167 VPWR.t1164 XThR.Tn[5].t37 XA.XIR[6].XIC[9].icell.PUM VPWR.t1163 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1168 XA.XIR[0].XIC[2].icell.PUM XThC.Tn[2].t24 XA.XIR[0].XIC[2].icell.Ien VPWR.t1269 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1169 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1557 VPWR.t1559 VPWR.t1558 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1170 VPWR.t518 XThR.Tn[8].t41 XA.XIR[9].XIC[10].icell.PUM VPWR.t517 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1171 VGND.t998 Vbias.t104 XA.XIR[1].XIC[13].icell.SM VGND.t997 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1172 VGND.t1000 Vbias.t105 XA.XIR[0].XIC[6].icell.SM VGND.t999 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1173 VGND.t2384 XThC.Tn[5].t22 XA.XIR[0].XIC[5].icell.PDM VGND.t2383 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1174 VGND.t1002 Vbias.t106 XA.XIR[4].XIC[14].icell.SM VGND.t1001 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1175 VGND.t2499 XThC.XTB7.A XThC.XTB7.Y VGND.t2498 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1176 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[7].t31 VGND.t1215 VGND.t1214 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1177 XA.XIR[2].XIC[8].icell.Ien XThR.Tn[2].t35 VPWR.t810 VPWR.t809 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1178 VPWR.t1130 XThR.Tn[1].t39 XA.XIR[2].XIC[3].icell.PUM VPWR.t1129 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1179 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t2 VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1180 XA.XIR[15].XIC[2].icell.SM XA.XIR[15].XIC[2].icell.Ien Iout.t235 VGND.t2438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1181 a_n997_2667# XThR.XTBN.Y.t51 VGND.t409 VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1182 VPWR.t1005 XThR.Tn[14].t35 XA.XIR[15].XIC[6].icell.PUM VPWR.t1004 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1183 VPWR.t23 XThR.Tn[13].t33 XA.XIR[14].XIC[7].icell.PUM VPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1184 a_7875_9569# XThC.XTBN.Y.t49 VGND.t1446 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1185 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[0].t39 VGND.t1271 VGND.t1270 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1186 VGND.t310 XThC.Tn[10].t24 XA.XIR[14].XIC[10].icell.PDM VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1187 VGND.t411 XThR.XTBN.Y.t52 a_n997_3979# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1188 XA.XIR[0].XIC_15.icell.Ien XThR.Tn[0].t40 VPWR.t896 VPWR.t895 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1189 XA.XIR[1].XIC[9].icell.SM XA.XIR[1].XIC[9].icell.Ien Iout.t104 VGND.t941 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1190 XA.XIR[13].XIC[5].icell.PUM XThC.Tn[5].t23 XA.XIR[13].XIC[5].icell.Ien VPWR.t859 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1191 XThC.Tn[14].t10 XThC.XTBN.Y.t50 VPWR.t953 VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1192 a_n1049_6699# XThR.XTB4.Y VPWR.t468 VPWR.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1193 a_4861_9615# XThC.XTBN.Y.t51 XThC.Tn[3].t3 VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1194 VGND.t1004 Vbias.t107 XA.XIR[10].XIC[8].icell.SM VGND.t1003 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1195 VGND.t760 XThC.Tn[7].t20 XA.XIR[10].XIC[7].icell.PDM VGND.t759 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1196 VGND.t1006 Vbias.t108 XA.XIR[13].XIC[9].icell.SM VGND.t1005 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1197 XA.XIR[12].XIC[10].icell.Ien XThR.Tn[12].t39 VPWR.t1284 VPWR.t1283 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1198 XThC.Tn[2].t0 XThC.XTB3.Y.t9 VGND.t851 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1199 XThC.Tn[9].t10 XThC.XTBN.Y.t52 VPWR.t954 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1200 XThC.Tn[5].t8 XThC.XTBN.Y.t53 VGND.t1447 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1201 a_n1335_8107# XThR.XTB6.A XThR.XTB2.Y VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1202 VGND.t1008 Vbias.t109 XA.XIR[0].XIC[10].icell.SM VGND.t1007 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1203 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[13].t34 VGND.t18 VGND.t17 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1204 VGND.t840 XThC.Tn[13].t26 XA.XIR[1].XIC[13].icell.PDM VGND.t839 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1205 XA.XIR[15].XIC[5].icell.Ien VPWR.t1554 VPWR.t1556 VPWR.t1555 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1206 VGND.t1855 VGND.t1853 XA.XIR[11].XIC_dummy_right.icell.SM VGND.t1854 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1207 VPWR.t1195 XThC.XTB1.Y.t11 a_2979_9615# VPWR.t1194 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1208 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1987 XA.XIR[1].XIC_dummy_left.icell.Ien VGND.t2324 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1209 XThC.Tn[0].t0 XThC.XTBN.Y.t54 a_2979_9615# VPWR.t955 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1210 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[3].t39 XA.XIR[3].XIC[11].icell.Ien VGND.t860 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1211 VPWR.t520 XThR.Tn[8].t42 XA.XIR[9].XIC[5].icell.PUM VPWR.t519 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1212 VPWR.t25 XThR.Tn[13].t35 XA.XIR[14].XIC[11].icell.PUM VPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1213 XThR.Tn[12].t5 XThR.XTB5.Y VPWR.t752 VPWR.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1214 XA.XIR[8].XIC[4].icell.PUM XThC.Tn[4].t27 XA.XIR[8].XIC[4].icell.Ien VPWR.t83 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1215 XA.XIR[12].XIC[12].icell.PUM XThC.Tn[12].t24 XA.XIR[12].XIC[12].icell.Ien VPWR.t610 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1216 VGND.t1010 Vbias.t110 XA.XIR[0].XIC[1].icell.SM VGND.t1009 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1217 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1552 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1553 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1218 XA.XIR[4].XIC[5].icell.SM XA.XIR[4].XIC[5].icell.Ien Iout.t86 VGND.t783 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1219 VGND.t945 XThC.Tn[0].t24 XA.XIR[0].XIC[0].icell.PDM VGND.t944 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1220 XThR.Tn[6].t10 XThR.XTBN.Y.t53 VGND.t413 VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1221 a_n1049_5611# XThR.XTBN.Y.t54 XThR.Tn[5].t10 VPWR.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1222 XA.XIR[15].XIC[13].icell.PUM XThC.Tn[13].t27 XA.XIR[15].XIC[13].icell.Ien VPWR.t622 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1223 VGND.t388 XThR.XTBN.Y.t55 a_n997_2891# VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1224 VGND.t1926 XThR.XTB7.B XThR.XTB7.Y VGND.t1925 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1225 XA.XIR[2].XIC[3].icell.Ien XThR.Tn[2].t36 VPWR.t806 VPWR.t805 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1226 XA.XIR[11].XIC[14].icell.SM XA.XIR[11].XIC[14].icell.Ien Iout.t135 VGND.t1182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1227 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[4].t40 XA.XIR[4].XIC[1].icell.Ien VGND.t697 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1228 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[3].t40 XA.XIR[3].XIC[2].icell.Ien VGND.t861 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1229 XA.XIR[14].XIC[7].icell.Ien XThR.Tn[14].t36 VPWR.t1007 VPWR.t1006 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1230 VPWR.t1009 XThR.Tn[14].t37 XA.XIR[15].XIC[1].icell.PUM VPWR.t1008 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1231 VGND.t2326 VPWR.t1988 XA.XIR[11].XIC_dummy_right.icell.PDM VGND.t2325 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1232 XA.XIR[2].XIC[8].icell.PUM XThC.Tn[8].t24 XA.XIR[2].XIC[8].icell.Ien VPWR.t1313 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1233 VPWR.t9 XThR.Tn[13].t36 XA.XIR[14].XIC[2].icell.PUM VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1234 a_n997_2667# XThR.XTB4.Y XThR.Tn[11].t3 VGND.t657 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1235 VPWR.t1551 VPWR.t1549 XA.XIR[12].XIC_15.icell.PUM VPWR.t1550 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1236 XA.XIR[1].XIC[4].icell.SM XA.XIR[1].XIC[4].icell.Ien Iout.t35 VGND.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1237 XA.XIR[10].XIC[4].icell.Ien XThR.Tn[10].t35 VPWR.t524 VPWR.t523 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1238 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1546 VPWR.t1548 VPWR.t1547 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1239 VGND.t1012 Vbias.t111 XA.XIR[6].XIC_15.icell.SM VGND.t1011 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1240 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout VGND.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1241 XA.XIR[14].XIC[7].icell.SM XA.XIR[14].XIC[7].icell.Ien Iout.t122 VGND.t1128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1242 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[13].t37 VGND.t6 VGND.t5 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1243 VGND.t1014 Vbias.t112 XA.XIR[10].XIC[3].icell.SM VGND.t1013 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1244 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1543 VPWR.t1545 VPWR.t1544 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1245 VGND.t1448 XThC.XTBN.Y.t55 XThC.Tn[1].t9 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1246 a_n1049_6405# XThR.XTB5.Y VPWR.t751 VPWR.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1247 VGND.t179 Vbias.t113 XA.XIR[13].XIC[4].icell.SM VGND.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1248 XA.XIR[12].XIC[5].icell.Ien XThR.Tn[12].t40 VPWR.t1286 VPWR.t1285 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1249 VPWR.t842 XThR.Tn[7].t32 XA.XIR[8].XIC[12].icell.PUM VPWR.t841 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1250 XA.XIR[0].XIC[13].icell.PDM XThR.Tn[0].t41 XA.XIR[0].XIC[13].icell.Ien VGND.t1272 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1251 VGND.t1852 VGND.t1850 XA.XIR[8].XIC_dummy_right.icell.SM VGND.t1851 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1252 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1989 XA.XIR[13].XIC_dummy_right.icell.Ien VGND.t2327 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1253 VGND.t2329 VPWR.t1990 XA.XIR[14].XIC_dummy_left.icell.PDM VGND.t2328 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1254 VPWR.t526 XThR.Tn[10].t36 XA.XIR[11].XIC[13].icell.PUM VPWR.t525 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1255 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[4].t41 VGND.t699 VGND.t698 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1256 XA.XIR[12].XIC[10].icell.PUM XThC.Tn[10].t25 XA.XIR[12].XIC[10].icell.Ien VPWR.t173 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1257 VPWR.t1089 XThR.XTB1.Y XThR.Tn[8].t6 VPWR.t1088 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1258 XA.XIR[8].XIC[0].icell.PUM XThC.Tn[0].t25 XA.XIR[8].XIC[0].icell.Ien VPWR.t673 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1259 XA.XIR[5].XIC[13].icell.SM XA.XIR[5].XIC[13].icell.Ien Iout.t81 VGND.t761 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1260 VPWR.t244 XThR.XTBN.Y.t56 XThR.Tn[7].t6 VPWR.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1261 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1541 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1542 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1262 VGND.t68 XThC.XTB2.Y XThC.Tn[1].t3 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1263 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1539 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1540 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1264 XA.XIR[8].XIC[14].icell.SM XA.XIR[8].XIC[14].icell.Ien Iout.t212 VGND.t2090 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1265 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[3].t41 XA.XIR[3].XIC[6].icell.Ien VGND.t862 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1266 XThC.Tn[12].t10 XThC.XTBN.Y.t56 VPWR.t956 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1267 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[1].t40 VGND.t1959 VGND.t1958 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1268 XA.XIR[14].XIC[11].icell.Ien XThR.Tn[14].t38 VPWR.t1011 VPWR.t1010 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1269 VGND.t1398 XThR.XTB2.Y XThR.Tn[1].t2 VGND.t1397 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1270 XThR.Tn[1].t6 XThR.XTBN.Y.t57 a_n1049_7787# VPWR.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1271 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[4].t42 VGND.t701 VGND.t700 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1272 XA.XIR[4].XIC[0].icell.SM XA.XIR[4].XIC[0].icell.Ien Iout.t130 VGND.t1172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1273 XA.XIR[6].XIC[12].icell.PUM XThC.Tn[12].t25 XA.XIR[6].XIC[12].icell.Ien VPWR.t611 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1274 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[12].t41 VGND.t2155 VGND.t2154 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1275 VGND.t920 XThC.Tn[11].t25 XA.XIR[7].XIC[11].icell.PDM VGND.t919 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1276 XA.XIR[2].XIC[13].icell.SM XA.XIR[2].XIC[13].icell.Ien Iout.t248 VGND.t2503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1277 XA.XIR[7].XIC[4].icell.Ien XThR.Tn[7].t33 VPWR.t844 VPWR.t843 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1278 VGND.t181 Vbias.t114 XA.XIR[3].XIC_15.icell.SM VGND.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1279 VGND.t183 Vbias.t115 XA.XIR[12].XIC[11].icell.SM VGND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1280 VGND.t1849 VGND.t1847 XA.XIR[11].XIC_dummy_left.icell.SM VGND.t1848 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1281 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10].t37 VPWR.t528 VPWR.t527 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1282 VGND.t2205 XThC.Tn[8].t25 XA.XIR[3].XIC[8].icell.PDM VGND.t2204 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1283 VGND.t447 XThC.Tn[14].t24 XA.XIR[3].XIC[14].icell.PDM VGND.t446 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1284 XA.XIR[14].XIC[2].icell.Ien XThR.Tn[14].t39 VPWR.t1013 VPWR.t1012 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1285 XThR.Tn[9].t5 XThR.XTB2.Y VPWR.t928 VPWR.t644 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1286 XThR.Tn[7].t1 XThR.XTBN.Y.t58 VGND.t390 VGND.t389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1287 VPWR.t745 data[1].t2 XThC.XTB6.A VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1288 XA.XIR[2].XIC[3].icell.PUM XThC.Tn[3].t25 XA.XIR[2].XIC[3].icell.Ien VPWR.t1823 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1289 VPWR.t846 XThR.Tn[7].t34 XA.XIR[8].XIC[10].icell.PUM VPWR.t845 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1290 XA.XIR[15].XIC[6].icell.PUM XThC.Tn[6].t26 XA.XIR[15].XIC[6].icell.Ien VPWR.t348 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1291 VPWR.t1538 VPWR.t1536 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1537 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1292 VGND.t1449 XThC.XTBN.Y.t57 a_7875_9569# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1293 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14].t40 XA.XIR[14].XIC[5].icell.Ien VGND.t1580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1294 VPWR.t246 XThR.XTBN.Y.t59 XThR.Tn[13].t10 VPWR.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1295 XA.XIR[1].XIC[8].icell.Ien XThR.Tn[1].t41 VPWR.t1132 VPWR.t1131 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1296 VPWR.t1535 VPWR.t1533 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1534 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1297 VGND.t2138 XThC.Tn[2].t25 XA.XIR[7].XIC[2].icell.PDM VGND.t2137 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1298 a_8739_10571# data[0].t1 XThC.XTB7.A VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1299 XA.XIR[14].XIC[2].icell.SM XA.XIR[14].XIC[2].icell.Ien Iout.t87 VGND.t852 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1300 VGND.t185 Vbias.t116 XA.XIR[9].XIC[11].icell.SM VGND.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1301 VPWR.t649 XThR.XTB3.Y XThR.Tn[10].t6 VPWR.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1302 XA.XIR[8].XIC[12].icell.Ien XThR.Tn[8].t43 VPWR.t103 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1303 VGND.t2174 XThC.Tn[9].t26 XA.XIR[15].XIC[9].icell.PDM VGND.t2173 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1304 XThC.Tn[3].t2 XThC.XTBN.Y.t58 a_4861_9615# VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1305 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5].t38 XA.XIR[5].XIC[8].icell.Ien VGND.t1991 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1306 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5].t39 XA.XIR[5].XIC[14].icell.Ien VGND.t1992 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1307 XA.XIR[11].XIC[13].icell.Ien XThR.Tn[11].t41 VPWR.t1805 VPWR.t1804 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1308 XThR.Tn[5].t2 XThR.XTB6.Y VGND.t214 VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1309 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9].t35 XA.XIR[9].XIC[14].icell.Ien VGND.t588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1310 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9].t36 XA.XIR[9].XIC[8].icell.Ien VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1311 VPWR.t1101 XThR.XTB7.B XThR.XTB4.Y VPWR.t1100 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1312 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout VGND.t1217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1313 XA.XIR[3].XIC[9].icell.PUM XThC.Tn[9].t27 XA.XIR[3].XIC[9].icell.Ien VPWR.t1299 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1314 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[4].t43 VGND.t2211 VGND.t2210 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1315 XA.XIR[12].XIC[5].icell.PUM XThC.Tn[5].t24 XA.XIR[12].XIC[5].icell.Ien VPWR.t860 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1316 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1991 VGND.t2331 VGND.t2330 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1317 XA.XIR[6].XIC[10].icell.PUM XThC.Tn[10].t26 XA.XIR[6].XIC[10].icell.Ien VPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1318 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout VGND.t883 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1319 VGND.t187 Vbias.t117 XA.XIR[12].XIC[9].icell.SM VGND.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1320 VGND.t922 XThC.Tn[11].t26 XA.XIR[4].XIC[11].icell.PDM VGND.t921 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1321 VPWR.t530 XThR.Tn[10].t38 XA.XIR[11].XIC[6].icell.PUM VPWR.t529 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1322 VGND.t1846 VGND.t1844 XA.XIR[8].XIC_dummy_left.icell.SM VGND.t1845 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1323 XA.XIR[7].XIC[0].icell.Ien XThR.Tn[7].t35 VPWR.t848 VPWR.t847 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1324 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t0 VGND.t1551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1325 VGND.t2064 XThC.Tn[1].t28 XA.XIR[1].XIC[1].icell.PDM VGND.t2063 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1326 VGND.t189 Vbias.t118 XA.XIR[7].XIC[7].icell.SM VGND.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1327 XA.XIR[5].XIC[9].icell.Ien XThR.Tn[5].t40 VPWR.t1166 VPWR.t1165 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1328 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[12].t42 VGND.t2157 VGND.t2156 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1329 VGND.t512 XThC.Tn[6].t27 XA.XIR[7].XIC[6].icell.PDM VGND.t511 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1330 VGND.t191 Vbias.t119 XA.XIR[6].XIC[8].icell.SM VGND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1331 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[11].t42 VGND.t2420 VGND.t2419 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1332 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t1992 VGND.t2333 VGND.t2332 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1333 VGND.t2140 XThC.Tn[2].t26 XA.XIR[4].XIC[2].icell.PDM VGND.t2139 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1334 XA.XIR[9].XIC[9].icell.Ien XThR.Tn[9].t37 VPWR.t335 VPWR.t334 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1335 VGND.t605 XThC.Tn[3].t26 XA.XIR[3].XIC[3].icell.PDM VGND.t604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1336 XA.XIR[14].XIC[8].icell.PUM XThC.Tn[8].t26 XA.XIR[14].XIC[8].icell.Ien VPWR.t1314 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1337 VGND.t193 Vbias.t120 XA.XIR[9].XIC[9].icell.SM VGND.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1338 XA.XIR[8].XIC[10].icell.Ien XThR.Tn[8].t44 VPWR.t105 VPWR.t104 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1339 XA.XIR[10].XIC_15.icell.SM XA.XIR[10].XIC_15.icell.Ien Iout.t148 VGND.t1218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1340 VPWR.t850 XThR.Tn[7].t36 XA.XIR[8].XIC[5].icell.PUM VPWR.t849 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1341 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6].t35 XA.XIR[6].XIC[11].icell.Ien VGND.t2517 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1342 XA.XIR[15].XIC[1].icell.PUM XThC.Tn[1].t29 XA.XIR[15].XIC[1].icell.Ien VPWR.t1181 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1343 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14].t41 XA.XIR[14].XIC[0].icell.Ien VGND.t1581 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1344 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[6].t36 VGND.t2238 VGND.t2237 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1345 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[6].t37 VGND.t2240 VGND.t2239 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1346 XA.XIR[1].XIC[3].icell.Ien XThR.Tn[1].t42 VPWR.t1134 VPWR.t1133 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1347 XA.XIR[6].XIC[6].icell.SM XA.XIR[6].XIC[6].icell.Ien Iout.t57 VGND.t496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1348 XA.XIR[13].XIC[14].icell.PUM XThC.Tn[14].t25 XA.XIR[13].XIC[14].icell.Ien VPWR.t306 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1349 VGND.t195 Vbias.t121 XA.XIR[15].XIC[5].icell.SM VGND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1350 VGND.t197 Vbias.t122 XA.XIR[14].XIC[6].icell.SM VGND.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1351 VGND.t117 XThC.Tn[4].t28 XA.XIR[15].XIC[4].icell.PDM VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1352 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6].t38 XA.XIR[6].XIC[2].icell.Ien VGND.t2241 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1353 VGND.t2335 VPWR.t1993 XA.XIR[10].XIC_dummy_right.icell.PDM VGND.t2334 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1354 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5].t41 XA.XIR[5].XIC[3].icell.Ien VGND.t1993 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1355 XThC.Tn[1].t8 XThC.XTBN.Y.t59 VGND.t1450 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1356 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9].t38 XA.XIR[9].XIC[3].icell.Ien VGND.t501 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1357 XA.XIR[4].XIC_15.icell.PDM XThR.Tn[4].t44 XA.XIR[4].XIC_15.icell.Ien VGND.t2212 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1358 VPWR.t1532 VPWR.t1530 XA.XIR[15].XIC_15.icell.PUM VPWR.t1531 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1359 XA.XIR[6].XIC[5].icell.PUM XThC.Tn[5].t25 XA.XIR[6].XIC[5].icell.Ien VPWR.t861 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1360 XA.XIR[0].XIC[1].icell.PDM XThR.Tn[0].t42 XA.XIR[0].XIC[1].icell.Ien VGND.t1273 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1361 XA.XIR[11].XIC[6].icell.Ien XThR.Tn[11].t43 VPWR.t1156 VPWR.t1155 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1362 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t1 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1363 VPWR.t804 XThR.Tn[2].t37 XA.XIR[3].XIC[4].icell.PUM VPWR.t803 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1364 VGND.t199 Vbias.t123 XA.XIR[3].XIC[8].icell.SM VGND.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1365 VGND.t514 XThC.Tn[6].t28 XA.XIR[4].XIC[6].icell.PDM VGND.t513 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1366 XA.XIR[15].XIC[14].icell.Ien VPWR.t1527 VPWR.t1529 VPWR.t1528 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1367 VGND.t201 Vbias.t124 XA.XIR[12].XIC[4].icell.SM VGND.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1368 VPWR.t532 XThR.Tn[10].t39 XA.XIR[11].XIC[1].icell.PUM VPWR.t531 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1369 VGND.t1201 XThC.Tn[7].t21 XA.XIR[3].XIC[7].icell.PDM VGND.t1200 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1370 VPWR.t1731 XThR.Tn[6].t39 XA.XIR[7].XIC[4].icell.PUM VPWR.t1730 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1371 VPWR.t1523 VPWR.t1521 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1522 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1372 XThR.Tn[13].t1 XThR.XTB6.Y a_n997_1579# VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1373 a_n1049_8581# XThR.XTBN.Y.t60 XThR.Tn[0].t6 VPWR.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1374 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout VGND.t2075 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1375 VPWR.t107 XThR.Tn[8].t45 XA.XIR[9].XIC[14].icell.PUM VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1376 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11].t44 XA.XIR[11].XIC[9].icell.Ien VGND.t1980 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1377 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[3].t42 VGND.t864 VGND.t863 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1378 VGND.t1629 Vbias.t125 XA.XIR[7].XIC[2].icell.SM VGND.t1628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1379 VGND.t1631 Vbias.t126 XA.XIR[6].XIC[3].icell.SM VGND.t1630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1380 XA.XIR[6].XIC[10].icell.SM XA.XIR[6].XIC[10].icell.Ien Iout.t88 VGND.t853 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1381 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[11].t45 VGND.t1982 VGND.t1981 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1382 XA.XIR[3].XIC[6].icell.SM XA.XIR[3].XIC[6].icell.Ien Iout.t20 VGND.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1383 XA.XIR[14].XIC[3].icell.PUM XThC.Tn[3].t27 XA.XIR[14].XIC[3].icell.Ien VPWR.t450 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1384 VGND.t1633 Vbias.t127 XA.XIR[9].XIC[4].icell.SM VGND.t1632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1385 XA.XIR[8].XIC[5].icell.Ien XThR.Tn[8].t46 VPWR.t109 VPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1386 VGND.t1635 Vbias.t128 XA.XIR[14].XIC[10].icell.SM VGND.t1634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1387 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[10].t40 VGND.t722 VGND.t721 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1388 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6].t40 XA.XIR[6].XIC[6].icell.Ien VGND.t2242 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1389 VGND.t1577 data[2].t1 XThC.XTB7.B VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1390 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5].t42 XA.XIR[5].XIC[7].icell.Ien VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1391 VGND.t392 XThR.XTBN.Y.t61 XThR.Tn[2].t3 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1392 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[3].t43 VGND.t1738 VGND.t1737 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1393 XA.XIR[13].XIC[11].icell.SM XA.XIR[13].XIC[11].icell.Ien Iout.t214 VGND.t2098 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1394 a_n1049_5317# XThR.XTB7.Y VPWR.t991 VPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1395 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9].t39 XA.XIR[9].XIC[7].icell.Ien VGND.t502 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1396 VGND.t1451 XThC.XTBN.Y.t60 XThC.Tn[4].t9 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1397 XA.XIR[5].XIC[12].icell.PUM XThC.Tn[12].t26 XA.XIR[5].XIC[12].icell.Ien VPWR.t1883 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1398 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[6].t41 VGND.t2244 VGND.t2243 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1399 XA.XIR[2].XIC_15.icell.PDM VPWR.t1994 VGND.t2337 VGND.t2336 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1400 XA.XIR[6].XIC[1].icell.SM XA.XIR[6].XIC[1].icell.Ien Iout.t55 VGND.t470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1401 XA.XIR[1].XIC[13].icell.SM XA.XIR[1].XIC[13].icell.Ien Iout.t177 VGND.t1493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1402 XA.XIR[9].XIC[12].icell.PUM XThC.Tn[12].t27 XA.XIR[9].XIC[12].icell.Ien VPWR.t1884 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1403 VGND.t1637 Vbias.t129 XA.XIR[15].XIC[0].icell.SM VGND.t1636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1404 XA.XIR[8].XIC[13].icell.PUM XThC.Tn[13].t28 XA.XIR[8].XIC[13].icell.Ien VPWR.t623 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1405 VGND.t1639 Vbias.t130 XA.XIR[14].XIC[1].icell.SM VGND.t1638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1406 VGND.t1641 Vbias.t131 XA.XIR[10].XIC[12].icell.SM VGND.t1640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1407 XA.XIR[4].XIC[14].icell.SM XA.XIR[4].XIC[14].icell.Ien Iout.t255 VGND.t2661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1408 XThR.Tn[3].t2 XThR.XTB4.Y VGND.t656 VGND.t655 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1409 VGND.t1643 Vbias.t132 XA.XIR[13].XIC[13].icell.SM VGND.t1642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1410 VPWR.t802 XThR.Tn[2].t38 XA.XIR[3].XIC[0].icell.PUM VPWR.t801 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1411 VGND.t2539 XThC.Tn[12].t28 XA.XIR[13].XIC[12].icell.PDM VGND.t2538 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1412 XA.XIR[12].XIC[14].icell.Ien XThR.Tn[12].t43 VPWR.t1288 VPWR.t1287 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1413 VPWR.t1733 XThR.Tn[6].t42 XA.XIR[7].XIC[0].icell.PUM VPWR.t1732 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1414 VPWR.t914 XThC.XTB7.Y a_6243_9615# VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1415 VPWR.t762 XThC.XTB6.Y XThC.Tn[13].t6 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1416 VPWR.t1526 VPWR.t1524 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1525 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1417 VGND.t990 data[1].t3 XThC.XTB5.A VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1418 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[0].t43 VGND.t2663 VGND.t2662 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1419 XA.XIR[3].XIC[4].icell.Ien XThR.Tn[3].t44 VPWR.t1032 VPWR.t1031 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1420 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[8].t47 VGND.t156 VGND.t155 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1421 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11].t46 VPWR.t1158 VPWR.t1157 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1422 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1518 VPWR.t1520 VPWR.t1519 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1423 VGND.t1645 Vbias.t133 XA.XIR[3].XIC[3].icell.SM VGND.t1644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1424 XA.XIR[7].XIC[7].icell.SM XA.XIR[7].XIC[7].icell.Ien Iout.t205 VGND.t2076 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1425 XA.XIR[3].XIC[10].icell.SM XA.XIR[3].XIC[10].icell.Ien Iout.t46 VGND.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1426 XA.XIR[10].XIC[13].icell.Ien XThR.Tn[10].t41 VPWR.t534 VPWR.t533 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1427 VPWR.t1907 XThR.Tn[0].t44 XA.XIR[1].XIC[12].icell.PUM VPWR.t1906 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1428 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[10].t42 VGND.t345 VGND.t344 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1429 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout VGND.t884 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1430 XA.XIR[10].XIC[8].icell.SM XA.XIR[10].XIC[8].icell.Ien Iout.t223 VGND.t2224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1431 VGND.t1453 XThC.XTBN.Y.t61 XThC.Tn[7].t2 VGND.t1452 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1432 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[3].t45 VGND.t1740 VGND.t1739 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1433 VPWR.t1317 XThR.Tn[4].t45 XA.XIR[5].XIC[12].icell.PUM VPWR.t1316 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1434 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11].t47 XA.XIR[11].XIC[4].icell.Ien VGND.t1983 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1435 XA.XIR[13].XIC[9].icell.SM XA.XIR[13].XIC[9].icell.Ien Iout.t196 VGND.t1917 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1436 XA.XIR[15].XIC[12].icell.PDM VPWR.t1995 XA.XIR[15].XIC[12].icell.Ien VGND.t2338 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1437 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[0].t45 VGND.t2665 VGND.t2664 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1438 XA.XIR[5].XIC[10].icell.PUM XThC.Tn[10].t27 XA.XIR[5].XIC[10].icell.Ien VPWR.t175 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1439 XThR.Tn[12].t4 XThR.XTB5.Y VPWR.t750 VPWR.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1440 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[6].t43 VGND.t2246 VGND.t2245 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1441 a_10915_9569# XThC.XTBN.Y.t62 VGND.t1455 VGND.t1454 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1442 XA.XIR[3].XIC[1].icell.SM XA.XIR[3].XIC[1].icell.Ien Iout.t215 VGND.t2099 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1443 XA.XIR[9].XIC[10].icell.PUM XThC.Tn[10].t28 XA.XIR[9].XIC[10].icell.Ien VPWR.t1304 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1444 XThR.Tn[6].t9 XThR.XTBN.Y.t62 VGND.t394 VGND.t393 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1445 VPWR.t1290 XThR.Tn[12].t44 XA.XIR[13].XIC[7].icell.PUM VPWR.t1289 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1446 XThC.Tn[3].t10 XThC.XTB4.Y.t7 VGND.t2473 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1447 XThC.Tn[9].t5 XThC.XTB2.Y VPWR.t51 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1448 VGND.t2184 XThC.Tn[10].t29 XA.XIR[13].XIC[10].icell.PDM VGND.t2183 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1449 a_n997_2667# XThR.XTB4.Y XThR.Tn[11].t2 VGND.t654 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1450 VGND.t424 XThC.Tn[11].t27 XA.XIR[0].XIC[11].icell.PDM VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1451 XA.XIR[15].XIC[5].icell.PDM XThR.Tn[14].t42 VGND.t1583 VGND.t1582 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1452 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[5].t43 VGND.t75 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1453 VGND.t1647 Vbias.t134 XA.XIR[5].XIC[11].icell.SM VGND.t1646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1454 XA.XIR[3].XIC[0].icell.Ien XThR.Tn[3].t46 VPWR.t1034 VPWR.t1033 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1455 XA.XIR[9].XIC_15.icell.SM XA.XIR[9].XIC_15.icell.Ien Iout.t167 VGND.t1390 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1456 VGND.t2340 VPWR.t1996 XA.XIR[1].XIC_15.icell.PDM VGND.t2339 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1457 VPWR.t1136 XThR.Tn[1].t43 XA.XIR[2].XIC[9].icell.PUM VPWR.t1135 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1458 VPWR.t1909 XThR.Tn[0].t46 XA.XIR[1].XIC[10].icell.PUM VPWR.t1908 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1459 XA.XIR[7].XIC[13].icell.Ien XThR.Tn[7].t37 VPWR.t852 VPWR.t851 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1460 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1515 VPWR.t1517 VPWR.t1516 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1461 VPWR.t1319 XThR.Tn[4].t46 XA.XIR[5].XIC[10].icell.PUM VPWR.t1318 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1462 XA.XIR[15].XIC[10].icell.PDM VPWR.t1997 XA.XIR[15].XIC[10].icell.Ien VGND.t2341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1463 XA.XIR[12].XIC[14].icell.PUM XThC.Tn[14].t26 XA.XIR[12].XIC[14].icell.Ien VPWR.t307 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1464 XA.XIR[8].XIC[6].icell.PUM XThC.Tn[6].t29 XA.XIR[8].XIC[6].icell.Ien VPWR.t349 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1465 VGND.t1924 XThR.XTB7.B a_n1335_8331# VGND.t1923 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1466 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[0].t47 VGND.t2667 VGND.t2666 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1467 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12].t45 XA.XIR[12].XIC[12].icell.Ien VGND.t2158 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1468 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[8].t48 VGND.t158 VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1469 VGND.t2142 XThC.Tn[2].t27 XA.XIR[0].XIC[2].icell.PDM VGND.t2141 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1470 XA.XIR[11].XIC[7].icell.PUM XThC.Tn[7].t22 XA.XIR[11].XIC[7].icell.Ien VPWR.t837 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1471 VPWR.t1764 XThC.XTBN.Y.t63 XThC.Tn[9].t9 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1472 XA.XIR[15].XIC_15.icell.PUM VPWR.t1513 XA.XIR[15].XIC_15.icell.Ien VPWR.t1514 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1473 XA.XIR[7].XIC[2].icell.SM XA.XIR[7].XIC[2].icell.Ien Iout.t243 VGND.t2484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1474 a_10051_9569# XThC.XTBN.Y.t64 VGND.t2254 VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1475 VGND.t2176 XThC.Tn[9].t28 XA.XIR[8].XIC[9].icell.PDM VGND.t2175 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1476 XA.XIR[10].XIC[3].icell.SM XA.XIR[10].XIC[3].icell.Ien Iout.t146 VGND.t1213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1477 VPWR.t249 XThR.XTBN.Y.t63 XThR.Tn[7].t5 VPWR.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1478 VPWR.t1292 XThR.Tn[12].t46 XA.XIR[13].XIC[11].icell.PUM VPWR.t1291 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1479 XA.XIR[7].XIC[4].icell.PUM XThC.Tn[4].t29 XA.XIR[7].XIC[4].icell.Ien VPWR.t84 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1480 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1511 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1512 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1481 XA.XIR[13].XIC[4].icell.SM XA.XIR[13].XIC[4].icell.Ien Iout.t222 VGND.t2223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1482 VPWR.t337 XThR.Tn[9].t40 XA.XIR[10].XIC[7].icell.PUM VPWR.t336 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1483 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[2].t39 XA.XIR[2].XIC[8].icell.Ien VGND.t717 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1484 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[2].t40 XA.XIR[2].XIC[14].icell.Ien VGND.t716 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1485 XThC.Tn[11].t5 XThC.XTB4.Y.t8 VPWR.t1028 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1486 VGND.t395 XThR.XTBN.Y.t64 XThR.Tn[1].t10 VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1487 XThR.Tn[1].t5 XThR.XTBN.Y.t65 a_n1049_7787# VPWR.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1488 a_7651_9569# XThC.XTBN.Y.t65 VGND.t2255 VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1489 XA.XIR[5].XIC[5].icell.PUM XThC.Tn[5].t26 XA.XIR[5].XIC[5].icell.Ien VPWR.t862 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1490 VGND.t1649 Vbias.t135 XA.XIR[11].XIC[5].icell.SM VGND.t1648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1491 XA.XIR[10].XIC[6].icell.Ien XThR.Tn[10].t43 VPWR.t217 VPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1492 XA.XIR[9].XIC[5].icell.PUM XThC.Tn[5].t27 XA.XIR[9].XIC[5].icell.Ien VPWR.t863 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1493 XA.XIR[13].XIC[7].icell.Ien XThR.Tn[13].t38 VPWR.t11 VPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1494 VGND.t1651 Vbias.t136 XA.XIR[5].XIC[9].icell.SM VGND.t1650 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1495 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t1998 VGND.t2343 VGND.t2342 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1496 VPWR.t1294 XThR.Tn[12].t47 XA.XIR[13].XIC[2].icell.PUM VPWR.t1293 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1497 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout VGND.t1407 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1498 VPWR.t285 XThR.Tn[7].t38 XA.XIR[8].XIC[14].icell.PUM VPWR.t284 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1499 XA.XIR[0].XIC_15.icell.PDM XThR.Tn[0].t48 XA.XIR[0].XIC_15.icell.Ien VGND.t2668 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1500 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10].t44 XA.XIR[10].XIC[9].icell.Ien VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1501 XThR.Tn[6].t1 XThR.XTB7.Y VGND.t1550 VGND.t1549 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1502 a_n1049_5611# XThR.XTB6.Y VPWR.t125 VPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1503 XThR.Tn[9].t4 XThR.XTB2.Y VPWR.t927 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1504 VPWR.t1510 VPWR.t1508 XA.XIR[11].XIC_15.icell.PUM VPWR.t1509 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1505 VGND.t1997 Vbias.t137 XA.XIR[0].XIC[7].icell.SM VGND.t1996 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1506 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12].t48 XA.XIR[12].XIC[10].icell.Ien VGND.t2159 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1507 XThC.Tn[4].t8 XThC.XTBN.Y.t66 VGND.t2256 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1508 VGND.t516 XThC.Tn[6].t30 XA.XIR[0].XIC[6].icell.PDM VGND.t515 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1509 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[5].t44 VGND.t77 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1510 XA.XIR[15].XIC[0].icell.PDM XThR.Tn[14].t43 VGND.t1585 VGND.t1584 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1511 XA.XIR[11].XIC[11].icell.PUM XThC.Tn[11].t28 XA.XIR[11].XIC[11].icell.Ien VPWR.t290 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1512 VPWR.t252 XThR.XTBN.Y.t66 XThR.Tn[13].t9 VPWR.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1513 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[9].t41 VGND.t504 VGND.t503 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1514 XA.XIR[2].XIC[9].icell.Ien XThR.Tn[2].t41 VPWR.t800 VPWR.t799 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1515 VGND.t1843 VGND.t1841 XA.XIR[7].XIC_dummy_right.icell.SM VGND.t1842 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1516 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[12].t49 VGND.t2161 VGND.t2160 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1517 XA.XIR[12].XIC[11].icell.SM XA.XIR[12].XIC[11].icell.Ien Iout.t28 VGND.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1518 VPWR.t1911 XThR.Tn[0].t49 XA.XIR[1].XIC[5].icell.PUM VPWR.t1910 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1519 VGND.t2345 VPWR.t1999 XA.XIR[13].XIC_dummy_left.icell.PDM VGND.t2344 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1520 VPWR.t1321 XThR.Tn[4].t47 XA.XIR[5].XIC[5].icell.PUM VPWR.t1320 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1521 VPWR.t339 XThR.Tn[9].t42 XA.XIR[10].XIC[11].icell.PUM VPWR.t338 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1522 XA.XIR[8].XIC[1].icell.PUM XThC.Tn[1].t30 XA.XIR[8].XIC[1].icell.Ien VPWR.t1182 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1523 XA.XIR[4].XIC[4].icell.PUM XThC.Tn[4].t30 XA.XIR[4].XIC[4].icell.Ien VPWR.t85 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1524 VGND.t1911 XThR.XTB1.Y XThR.Tn[0].t1 VGND.t1400 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1525 XA.XIR[0].XIC[5].icell.SM XA.XIR[0].XIC[5].icell.Ien Iout.t221 VGND.t2222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1526 XThR.Tn[5].t5 XThR.XTBN.Y.t67 VGND.t396 VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1527 XA.XIR[7].XIC[0].icell.PUM XThC.Tn[0].t26 XA.XIR[7].XIC[0].icell.Ien VPWR.t674 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1528 XA.XIR[0].XIC[8].icell.PDM VGND.t1838 VGND.t1840 VGND.t1839 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1529 XA.XIR[0].XIC[14].icell.PDM VGND.t1835 VGND.t1837 VGND.t1836 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1530 VGND.t1922 XThR.XTB7.B XThR.XTB6.Y VGND.t1920 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 XA.XIR[11].XIC[2].icell.PUM XThC.Tn[2].t28 XA.XIR[11].XIC[2].icell.Ien VPWR.t1270 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1532 XA.XIR[6].XIC[14].icell.PUM XThC.Tn[14].t27 XA.XIR[6].XIC[14].icell.Ien VPWR.t308 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1533 VGND.t2257 XThC.XTBN.Y.t67 XThC.Tn[0].t5 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1534 VGND.t1999 Vbias.t138 XA.XIR[8].XIC[5].icell.SM VGND.t1998 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1535 XA.XIR[7].XIC[6].icell.Ien XThR.Tn[7].t39 VPWR.t287 VPWR.t286 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1536 XA.XIR[13].XIC[11].icell.Ien XThR.Tn[13].t39 VPWR.t13 VPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1537 VGND.t2001 Vbias.t139 XA.XIR[12].XIC[13].icell.SM VGND.t2000 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1538 VGND.t119 XThC.Tn[4].t31 XA.XIR[8].XIC[4].icell.PDM VGND.t118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1539 VGND.t2347 VPWR.t2000 XA.XIR[3].XIC_dummy_right.icell.PDM VGND.t2346 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1540 VGND.t2541 XThC.Tn[12].t29 XA.XIR[12].XIC[12].icell.PDM VGND.t2540 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1541 VGND.t2258 XThC.XTBN.Y.t68 XThC.Tn[3].t7 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1542 VGND.t2003 Vbias.t140 XA.XIR[15].XIC[14].icell.SM VGND.t2002 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1543 VGND.t1230 XThC.Tn[5].t28 XA.XIR[11].XIC[5].icell.PDM VGND.t1229 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1544 VGND.t842 XThC.Tn[13].t29 XA.XIR[15].XIC[13].icell.PDM VGND.t841 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1545 VPWR.t341 XThR.Tn[9].t43 XA.XIR[10].XIC[2].icell.PUM VPWR.t340 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1546 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[2].t42 XA.XIR[2].XIC[3].icell.Ien VGND.t715 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1547 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t2001 XA.XIR[15].XIC_dummy_left.icell.Ien VGND.t2348 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1548 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7].t40 XA.XIR[7].XIC[9].icell.Ien VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1549 XThC.Tn[7].t1 XThC.XTBN.Y.t69 VGND.t2260 VGND.t2259 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1550 VPWR.t1765 XThC.XTBN.Y.t70 XThC.Tn[12].t9 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1551 VGND.t2005 Vbias.t141 XA.XIR[11].XIC[0].icell.SM VGND.t2004 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1552 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10].t45 VPWR.t219 VPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1553 XA.XIR[6].XIC[4].icell.Ien XThR.Tn[6].t44 VPWR.t1735 VPWR.t1734 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1554 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1505 VPWR.t1507 VPWR.t1506 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1555 VGND.t2007 Vbias.t142 XA.XIR[2].XIC_15.icell.SM VGND.t2006 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1556 VGND.t2009 Vbias.t143 XA.XIR[6].XIC[12].icell.SM VGND.t2008 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1557 VGND.t2207 XThC.Tn[8].t27 XA.XIR[2].XIC[8].icell.PDM VGND.t2206 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1558 VGND.t449 XThC.Tn[14].t28 XA.XIR[2].XIC[14].icell.PDM VGND.t448 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1559 VPWR.t926 XThR.XTB2.Y a_n1049_7787# VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1560 XA.XIR[13].XIC[2].icell.Ien XThR.Tn[13].t40 VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1561 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[9].t44 VGND.t506 VGND.t505 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1562 VGND.t2011 Vbias.t144 XA.XIR[5].XIC[4].icell.SM VGND.t2010 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1563 VGND.t2013 Vbias.t145 XA.XIR[9].XIC[13].icell.SM VGND.t2012 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1564 XA.XIR[9].XIC[8].icell.SM XA.XIR[9].XIC[8].icell.Ien Iout.t59 VGND.t499 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1565 XA.XIR[8].XIC[14].icell.Ien XThR.Tn[8].t49 VPWR.t111 VPWR.t110 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1566 VGND.t2262 XThC.XTBN.Y.t71 a_10915_9569# VGND.t2261 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1567 VPWR.t1064 VGND.t2695 XA.XIR[0].XIC[4].icell.PUM VPWR.t1063 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1568 VPWR.t1036 XThR.Tn[3].t47 XA.XIR[4].XIC[12].icell.PUM VPWR.t1035 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1569 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10].t46 XA.XIR[10].XIC[4].icell.Ien VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1570 VPWR.t798 XThR.Tn[2].t43 XA.XIR[3].XIC[13].icell.PUM VPWR.t797 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1571 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t2002 XA.XIR[5].XIC_dummy_right.icell.Ien VGND.t2349 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1572 XA.XIR[12].XIC[9].icell.SM XA.XIR[12].XIC[9].icell.Ien Iout.t116 VGND.t1116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1573 XA.XIR[11].XIC_15.icell.Ien XThR.Tn[11].t48 VPWR.t1160 VPWR.t1159 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1574 XThC.Tn[11].t6 XThC.XTB4.Y.t9 a_8963_9569# VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1575 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13].t41 XA.XIR[13].XIC[5].icell.Ien VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1576 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t2003 XA.XIR[9].XIC_dummy_right.icell.Ien VGND.t2350 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1577 VPWR.t1737 XThR.Tn[6].t45 XA.XIR[7].XIC[13].icell.PUM VPWR.t1736 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1578 VGND.t1709 XThC.XTB4.Y.t10 XThC.Tn[3].t9 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1579 VGND.t2015 Vbias.t146 XA.XIR[0].XIC[2].icell.SM VGND.t2014 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1580 XThR.Tn[14].t11 XThR.XTBN.Y.t68 VPWR.t254 VPWR.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1581 XA.XIR[4].XIC[0].icell.PUM XThC.Tn[0].t27 XA.XIR[4].XIC[0].icell.Ien VPWR.t675 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1582 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1503 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1504 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1583 a_7875_9569# XThC.XTBN.Y.t72 VGND.t2263 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1584 VPWR.t123 XThR.XTB6.Y XThR.Tn[13].t7 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1585 VGND.t2186 XThC.Tn[10].t30 XA.XIR[12].XIC[10].icell.PDM VGND.t2185 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1586 XA.XIR[2].XIC[9].icell.PUM XThC.Tn[9].t29 XA.XIR[2].XIC[9].icell.Ien VPWR.t1300 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1587 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[2].t44 XA.XIR[2].XIC[7].icell.Ien VGND.t718 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1588 XA.XIR[0].XIC[0].icell.SM XA.XIR[0].XIC[0].icell.Ien Iout.t141 VGND.t1208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1589 XA.XIR[0].XIC[3].icell.PDM VGND.t1832 VGND.t1834 VGND.t1833 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1590 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t2004 XA.XIR[12].XIC_dummy_left.icell.Ien VGND.t2351 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1591 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14].t44 XA.XIR[14].XIC[11].icell.Ien VGND.t1586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1592 XThC.Tn[11].t7 XThC.XTB4.Y.t11 a_8963_9569# VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1593 VGND.t2017 Vbias.t147 XA.XIR[8].XIC[0].icell.SM VGND.t2016 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1594 XA.XIR[7].XIC[1].icell.Ien XThR.Tn[7].t41 VPWR.t289 VPWR.t288 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1595 VGND.t2019 Vbias.t148 XA.XIR[3].XIC[12].icell.SM VGND.t2018 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1596 XA.XIR[6].XIC[0].icell.Ien XThR.Tn[6].t46 VPWR.t1739 VPWR.t1738 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1597 VGND.t1831 VGND.t1829 XA.XIR[7].XIC_dummy_left.icell.SM VGND.t1830 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1598 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1501 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1502 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1599 XThC.Tn[0].t9 XThC.XTB1.Y.t12 VGND.t2072 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1600 XA.XIR[15].XIC[5].icell.SM XA.XIR[15].XIC[5].icell.Ien Iout.t95 VGND.t880 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1601 VGND.t2264 XThC.XTBN.Y.t73 a_10051_9569# VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1602 VGND.t947 XThC.Tn[0].t28 XA.XIR[11].XIC[0].icell.PDM VGND.t946 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1603 VPWR.t1038 XThR.Tn[3].t48 XA.XIR[4].XIC[10].icell.PUM VPWR.t1037 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1604 VGND.t2543 XThC.Tn[12].t30 XA.XIR[6].XIC[12].icell.PDM VGND.t2542 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1605 XThR.XTB1.Y XThR.XTB5.A VPWR.t832 VPWR.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1606 VPWR.t1062 VGND.t2696 XA.XIR[0].XIC[0].icell.PUM VPWR.t1061 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1607 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7].t42 XA.XIR[7].XIC[4].icell.Ien VGND.t418 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1608 XThR.Tn[13].t0 XThR.XTB6.Y a_n997_1579# VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1609 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14].t45 XA.XIR[14].XIC[2].icell.Ien VGND.t1587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1610 XA.XIR[10].XIC[7].icell.PUM XThC.Tn[7].t23 XA.XIR[10].XIC[7].icell.Ien VPWR.t838 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1611 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2005 VGND.t2353 VGND.t2352 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1612 VGND.t607 XThC.Tn[3].t28 XA.XIR[2].XIC[3].icell.PDM VGND.t606 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1613 XA.XIR[13].XIC[8].icell.PUM XThC.Tn[8].t28 XA.XIR[13].XIC[8].icell.Ien VPWR.t1315 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1614 VGND.t2265 XThC.XTBN.Y.t74 a_7651_9569# VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1615 XA.XIR[4].XIC[12].icell.Ien XThR.Tn[4].t48 VPWR.t1323 VPWR.t1322 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1616 XA.XIR[9].XIC[3].icell.SM XA.XIR[9].XIC[3].icell.Ien Iout.t61 VGND.t559 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1617 XThC.XTBN.Y.t0 XThC.XTBN.A VGND.t2082 VGND.t2081 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1618 XA.XIR[3].XIC[13].icell.Ien XThR.Tn[3].t49 VPWR.t1040 VPWR.t1039 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1619 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1498 VPWR.t1500 VPWR.t1499 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1620 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[1].t44 XA.XIR[1].XIC[14].icell.Ien VGND.t1960 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1621 XA.XIR[12].XIC[4].icell.SM XA.XIR[12].XIC[4].icell.Ien Iout.t136 VGND.t1192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1622 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[1].t45 XA.XIR[1].XIC[8].icell.Ien VGND.t1961 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1623 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout VGND.t1171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1624 a_n1335_7243# XThR.XTB7.A XThR.XTB3.Y VGND.t1194 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1625 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13].t42 XA.XIR[13].XIC[0].icell.Ien VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1626 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8].t50 XA.XIR[8].XIC[12].icell.Ien VGND.t776 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1627 XA.XIR[0].XIC[7].icell.PDM VGND.t1826 VGND.t1828 VGND.t1827 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1628 a_n1049_5317# XThR.XTBN.Y.t69 XThR.Tn[6].t6 VPWR.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1629 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11].t49 XA.XIR[11].XIC[13].icell.Ien VGND.t1984 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1630 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2006 VGND.t2355 VGND.t2354 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1631 a_4067_9615# XThC.XTB3.Y.t10 VPWR.t628 VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1632 VPWR.t1767 XThC.XTBN.Y.t75 XThC.Tn[7].t4 VPWR.t1766 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1633 VPWR.t796 XThR.Tn[2].t45 XA.XIR[3].XIC[6].icell.PUM VPWR.t795 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1634 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[11].t50 VGND.t1973 VGND.t1972 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1635 XA.XIR[15].XIC[8].icell.Ien VPWR.t1495 VPWR.t1497 VPWR.t1496 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1636 VPWR.t1741 XThR.Tn[6].t47 XA.XIR[7].XIC[6].icell.PUM VPWR.t1740 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1637 VGND.t471 XThR.XTBN.Y.t70 a_n997_1803# VGND.t406 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1638 VPWR.t58 XThR.Tn[5].t45 XA.XIR[6].XIC[7].icell.PUM VPWR.t57 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1639 XThR.Tn[3].t9 XThR.XTBN.Y.t71 VGND.t472 VGND.t342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1640 VGND.t2188 XThC.Tn[10].t31 XA.XIR[6].XIC[10].icell.PDM VGND.t2187 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1641 VPWR.t578 XThR.Tn[8].t51 XA.XIR[9].XIC[8].icell.PUM VPWR.t577 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1642 VPWR.t1029 XThC.XTB4.Y.t12 XThC.Tn[11].t8 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14].t46 XA.XIR[14].XIC[6].icell.Ien VGND.t1588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1644 XA.XIR[10].XIC[11].icell.PUM XThC.Tn[11].t29 XA.XIR[10].XIC[11].icell.Ien VPWR.t291 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1645 VGND.t1340 Vbias.t149 XA.XIR[2].XIC[8].icell.SM VGND.t1339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1646 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[12].t50 VGND.t2163 VGND.t2162 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1647 XA.XIR[1].XIC[9].icell.Ien XThR.Tn[1].t46 VPWR.t508 VPWR.t507 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1648 VGND.t1203 XThC.Tn[7].t24 XA.XIR[2].XIC[7].icell.PDM VGND.t1202 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1649 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[11].t51 VGND.t1975 VGND.t1974 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1650 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[7].t43 VGND.t420 VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1651 XA.XIR[4].XIC[10].icell.Ien XThR.Tn[4].t49 VPWR.t1325 VPWR.t1324 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1652 XA.XIR[15].XIC[0].icell.SM XA.XIR[15].XIC[0].icell.Ien Iout.t79 VGND.t747 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1653 VGND.t2357 VPWR.t2007 XA.XIR[12].XIC_dummy_left.icell.PDM VGND.t2356 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1654 XThC.Tn[0].t4 XThC.XTBN.Y.t76 VGND.t1432 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1655 XA.XIR[10].XIC[12].icell.SM XA.XIR[10].XIC[12].icell.Ien Iout.t40 VGND.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1656 VPWR.t1042 XThR.Tn[3].t50 XA.XIR[4].XIC[5].icell.PUM VPWR.t1041 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1657 XA.XIR[13].XIC[13].icell.SM XA.XIR[13].XIC[13].icell.Ien Iout.t185 VGND.t1578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1658 XThC.Tn[3].t6 XThC.XTBN.Y.t77 VGND.t1433 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1659 VGND.t2209 XThC.Tn[8].t29 XA.XIR[14].XIC[8].icell.PDM VGND.t2208 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1660 VGND.t1079 XThC.Tn[14].t29 XA.XIR[14].XIC[14].icell.PDM VGND.t1078 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1661 XA.XIR[10].XIC[2].icell.PUM XThC.Tn[2].t29 XA.XIR[10].XIC[2].icell.Ien VPWR.t1271 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1662 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8].t52 XA.XIR[8].XIC[10].icell.Ien VGND.t777 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1663 XA.XIR[5].XIC[14].icell.PUM XThC.Tn[14].t30 XA.XIR[5].XIC[14].icell.Ien VPWR.t699 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1664 XA.XIR[13].XIC[3].icell.PUM XThC.Tn[3].t29 XA.XIR[13].XIC[3].icell.Ien VPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1665 XA.XIR[9].XIC[14].icell.PUM XThC.Tn[14].t31 XA.XIR[9].XIC[14].icell.Ien VPWR.t700 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1666 XA.XIR[8].XIC_15.icell.PUM VPWR.t1493 XA.XIR[8].XIC_15.icell.Ien VPWR.t1494 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1667 a_n1049_8581# XThR.XTB1.Y VPWR.t1087 VPWR.t1086 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1668 VGND.t2066 XThC.Tn[1].t31 XA.XIR[15].XIC[1].icell.PDM VGND.t2065 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1669 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[8].t53 VGND.t779 VGND.t778 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1670 VPWR.t1492 VPWR.t1490 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1491 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1671 VGND.t1342 Vbias.t150 XA.XIR[10].XIC[6].icell.SM VGND.t1341 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1672 VGND.t1232 XThC.Tn[5].t29 XA.XIR[10].XIC[5].icell.PDM VGND.t1231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1673 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[1].t47 XA.XIR[1].XIC[3].icell.Ien VGND.t702 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1674 XA.XIR[12].XIC[8].icell.Ien XThR.Tn[12].t51 VPWR.t1237 VPWR.t1236 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1675 VPWR.t60 XThR.Tn[5].t46 XA.XIR[6].XIC[11].icell.PUM VPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1676 XA.XIR[0].XIC[4].icell.PUM XThC.Tn[4].t32 XA.XIR[0].XIC[4].icell.Ien VPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1677 VGND.t1344 Vbias.t151 XA.XIR[1].XIC_15.icell.SM VGND.t1343 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1678 XA.XIR[7].XIC[13].icell.PUM XThC.Tn[13].t30 XA.XIR[7].XIC[13].icell.Ien VPWR.t624 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1679 XThC.XTB1.Y.t1 XThC.XTB5.A a_3299_10575# VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1680 XA.XIR[3].XIC[6].icell.Ien XThR.Tn[3].t51 VPWR.t1044 VPWR.t1043 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1681 VPWR.t794 XThR.Tn[2].t46 XA.XIR[3].XIC[1].icell.PUM VPWR.t793 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1682 VGND.t868 XThR.XTB3.Y XThR.Tn[2].t8 VGND.t658 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1683 XA.XIR[15].XIC[3].icell.Ien VPWR.t1487 VPWR.t1489 VPWR.t1488 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1684 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[11].t52 VGND.t1977 VGND.t1976 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1685 VGND.t1346 Vbias.t152 XA.XIR[11].XIC[14].icell.SM VGND.t1345 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1686 XA.XIR[10].XIC_15.icell.Ien XThR.Tn[10].t47 VPWR.t221 VPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1687 XA.XIR[14].XIC[9].icell.PUM XThC.Tn[9].t30 XA.XIR[14].XIC[9].icell.Ien VPWR.t1301 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1688 VPWR.t1743 XThR.Tn[6].t48 XA.XIR[7].XIC[1].icell.PUM VPWR.t1742 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1689 VPWR.t62 XThR.Tn[5].t47 XA.XIR[6].XIC[2].icell.PUM VPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1690 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout VGND.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1691 VPWR.t613 XThR.Tn[0].t50 XA.XIR[1].XIC[14].icell.PUM VPWR.t612 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1692 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[3].t52 XA.XIR[3].XIC[9].icell.Ien VGND.t1741 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1693 VPWR.t1185 XThR.Tn[4].t50 XA.XIR[5].XIC[14].icell.PUM VPWR.t1184 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1694 VPWR.t580 XThR.Tn[8].t54 XA.XIR[9].XIC[3].icell.PUM VPWR.t579 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1695 VGND.t1435 XThC.XTBN.Y.t78 XThC.Tn[6].t10 VGND.t1434 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1696 VGND.t1348 Vbias.t153 XA.XIR[2].XIC[3].icell.SM VGND.t1347 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1697 XA.XIR[6].XIC[7].icell.SM XA.XIR[6].XIC[7].icell.Ien Iout.t132 VGND.t1178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1698 XThC.Tn[10].t1 XThC.XTB3.Y.t11 VPWR.t629 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1699 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[7].t44 VGND.t422 VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1700 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[2].t47 VGND.t1061 VGND.t1060 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1701 XA.XIR[4].XIC[5].icell.Ien XThR.Tn[4].t51 VPWR.t1187 VPWR.t1186 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1702 VGND.t1825 VGND.t1823 XA.XIR[0].XIC_dummy_right.icell.SM VGND.t1824 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1703 VGND.t1350 Vbias.t154 XA.XIR[14].XIC[7].icell.SM VGND.t1349 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1704 VGND.t1352 Vbias.t155 XA.XIR[10].XIC[10].icell.SM VGND.t1351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1705 XThC.Tn[14].t6 XThC.XTB7.Y VPWR.t913 VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1706 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[5].t48 VGND.t79 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1707 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[1].t48 XA.XIR[1].XIC[7].icell.Ien VGND.t703 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1708 VGND.t2359 VPWR.t2008 XA.XIR[6].XIC_dummy_left.icell.PDM VGND.t2358 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1709 VGND.t2073 XThC.XTB1.Y.t13 XThC.Tn[0].t10 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1710 VGND.t609 XThC.Tn[3].t30 XA.XIR[14].XIC[3].icell.PDM VGND.t608 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1711 XA.XIR[0].XIC[0].icell.PUM XThC.Tn[0].t29 XA.XIR[0].XIC[0].icell.Ien VPWR.t676 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1712 XA.XIR[1].XIC[12].icell.PUM XThC.Tn[12].t31 XA.XIR[1].XIC[12].icell.Ien VPWR.t1885 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1713 XA.XIR[4].XIC[13].icell.PUM XThC.Tn[13].t31 XA.XIR[4].XIC[13].icell.Ien VPWR.t625 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1714 VGND.t1354 Vbias.t156 XA.XIR[10].XIC[1].icell.SM VGND.t1353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1715 XThR.Tn[8].t9 XThR.XTBN.Y.t72 VPWR.t323 VPWR.t322 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1716 XA.XIR[0].XIC[14].icell.SM XA.XIR[0].XIC[14].icell.Ien Iout.t133 VGND.t1179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1717 VGND.t1356 Vbias.t157 XA.XIR[5].XIC[13].icell.SM VGND.t1355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1718 XA.XIR[14].XIC[5].icell.SM XA.XIR[14].XIC[5].icell.Ien Iout.t183 VGND.t1565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1719 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[13].t43 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1720 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[13].t44 VGND.t12 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1721 VGND.t949 XThC.Tn[0].t30 XA.XIR[10].XIC[0].icell.PDM VGND.t948 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1722 VGND.t2545 XThC.Tn[12].t32 XA.XIR[5].XIC[12].icell.PDM VGND.t2544 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1723 XA.XIR[12].XIC[3].icell.Ien XThR.Tn[12].t52 VPWR.t1239 VPWR.t1238 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1724 VGND.t2547 XThC.Tn[12].t33 XA.XIR[9].XIC[12].icell.PDM VGND.t2546 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1725 VGND.t1358 Vbias.t158 XA.XIR[8].XIC[14].icell.SM VGND.t1357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1726 XA.XIR[7].XIC_15.icell.Ien XThR.Tn[7].t45 VPWR.t733 VPWR.t732 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1727 VGND.t844 XThC.Tn[13].t32 XA.XIR[8].XIC[13].icell.PDM VGND.t843 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1728 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t2009 XA.XIR[8].XIC_dummy_left.icell.Ien VGND.t2360 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1729 a_n1049_5611# XThR.XTBN.Y.t73 XThR.Tn[5].t9 VPWR.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1730 XA.XIR[3].XIC[1].icell.Ien XThR.Tn[3].t53 VPWR.t1046 VPWR.t1045 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1731 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[4].t52 VGND.t2068 VGND.t2067 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1732 XA.XIR[12].XIC[8].icell.PUM XThC.Tn[8].t30 XA.XIR[12].XIC[8].icell.Ien VPWR.t689 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1733 VGND.t1360 Vbias.t159 XA.XIR[4].XIC[11].icell.SM VGND.t1359 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1734 XA.XIR[3].XIC[7].icell.SM XA.XIR[3].XIC[7].icell.Ien Iout.t9 VGND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1735 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[2].t48 VGND.t1059 VGND.t1058 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1736 XThR.XTBN.A data[7].t1 VGND.t2101 VGND.t2100 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1737 XA.XIR[6].XIC[13].icell.Ien XThR.Tn[6].t49 VPWR.t1745 VPWR.t1744 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1738 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[3].t54 XA.XIR[3].XIC[4].icell.Ien VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1739 XThC.Tn[14].t5 XThC.XTB7.Y VPWR.t912 VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1740 VPWR.t17 XThR.Tn[13].t45 XA.XIR[14].XIC[4].icell.PUM VPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1741 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11].t53 XA.XIR[11].XIC[1].icell.Ien VGND.t1978 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1742 XA.XIR[7].XIC[6].icell.PUM XThC.Tn[6].t31 XA.XIR[7].XIC[6].icell.Ien VPWR.t350 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1743 VPWR.t1060 VGND.t2697 XA.XIR[0].XIC[13].icell.PUM VPWR.t1059 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1744 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2010 XA.XIR[2].XIC_dummy_right.icell.Ien VGND.t2361 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1745 VGND.t1205 XThC.Tn[7].t25 XA.XIR[14].XIC[7].icell.PDM VGND.t1204 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1746 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10].t48 XA.XIR[10].XIC[13].icell.Ien VGND.t348 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1747 XThC.XTB2.Y XThC.XTB7.B VPWR.t742 VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1748 XA.XIR[1].XIC[10].icell.PUM XThC.Tn[10].t32 XA.XIR[1].XIC[10].icell.Ien VPWR.t1305 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1749 XA.XIR[6].XIC[2].icell.SM XA.XIR[6].XIC[2].icell.Ien Iout.t160 VGND.t1291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1750 XA.XIR[0].XIC[12].icell.Ien XThR.Tn[0].t51 VPWR.t615 VPWR.t614 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1751 XThR.Tn[5].t4 XThR.XTBN.Y.t74 VGND.t473 VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1752 VGND.t2178 XThC.Tn[9].t31 XA.XIR[7].XIC[9].icell.PDM VGND.t2177 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1753 XA.XIR[15].XIC[11].icell.PDM XThR.Tn[14].t47 VGND.t1590 VGND.t1589 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1754 VGND.t1362 Vbias.t160 XA.XIR[14].XIC[2].icell.SM VGND.t1361 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1755 VGND.t2190 XThC.Tn[10].t33 XA.XIR[5].XIC[10].icell.PDM VGND.t2189 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1756 XThR.Tn[10].t9 XThR.XTBN.Y.t75 VPWR.t324 VPWR.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1757 VPWR.t735 XThR.Tn[7].t46 XA.XIR[8].XIC[8].icell.PUM VPWR.t734 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1758 VGND.t2192 XThC.Tn[10].t34 XA.XIR[9].XIC[10].icell.PDM VGND.t2191 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1759 a_5949_9615# XThC.XTB6.Y VPWR.t761 VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1760 VGND.t91 Vbias.t161 XA.XIR[1].XIC[8].icell.SM VGND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1761 VGND.t93 Vbias.t162 XA.XIR[4].XIC[9].icell.SM VGND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1762 XA.XIR[14].XIC[0].icell.SM XA.XIR[14].XIC[0].icell.Ien Iout.t115 VGND.t1109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1763 XA.XIR[15].XIC[2].icell.PDM XThR.Tn[14].t48 VGND.t1592 VGND.t1591 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1764 VPWR.t630 XThC.XTB3.Y.t12 XThC.Tn[10].t2 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1765 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[13].t46 VGND.t14 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1766 VGND.t1822 VGND.t1820 XA.XIR[0].XIC_dummy_left.icell.SM VGND.t1821 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1767 XA.XIR[5].XIC_15.icell.SM XA.XIR[5].XIC_15.icell.Ien Iout.t193 VGND.t1914 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1768 XA.XIR[9].XIC[12].icell.SM XA.XIR[9].XIC[12].icell.Ien Iout.t178 VGND.t1500 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1769 XThC.Tn[13].t8 XThC.XTBN.Y.t79 VPWR.t950 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1770 XA.XIR[13].XIC_15.icell.PDM VPWR.t2011 VGND.t2363 VGND.t2362 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1771 a_n997_3755# XThR.XTBN.Y.t76 VGND.t474 VGND.t383 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1772 XA.XIR[12].XIC[13].icell.SM XA.XIR[12].XIC[13].icell.Ien Iout.t0 VGND.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1773 VPWR.t325 XThR.XTBN.Y.t77 XThR.Tn[14].t10 VPWR.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 XA.XIR[15].XIC[14].icell.SM XA.XIR[15].XIC[14].icell.Ien Iout.t98 VGND.t923 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1775 XA.XIR[4].XIC[6].icell.PUM XThC.Tn[6].t32 XA.XIR[4].XIC[6].icell.Ien VPWR.t351 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1776 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[8].t55 VGND.t781 VGND.t780 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1777 XA.XIR[3].XIC[7].icell.PUM XThC.Tn[7].t26 XA.XIR[3].XIC[7].icell.Ien VPWR.t839 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1778 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[4].t53 VGND.t2070 VGND.t2069 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1779 XA.XIR[12].XIC[3].icell.PUM XThC.Tn[3].t31 XA.XIR[12].XIC[3].icell.Ien VPWR.t452 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1780 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2012 VGND.t2365 VGND.t2364 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1781 VPWR.t19 XThR.Tn[13].t47 XA.XIR[14].XIC[0].icell.PUM VPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1782 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7].t47 XA.XIR[7].XIC[13].icell.Ien VGND.t1117 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1783 XA.XIR[0].XIC[10].icell.Ien XThR.Tn[0].t52 VPWR.t617 VPWR.t616 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1784 XA.XIR[3].XIC[2].icell.SM XA.XIR[3].XIC[2].icell.Ien Iout.t119 VGND.t1125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1785 XA.XIR[6].XIC[8].icell.PUM XThC.Tn[8].t31 XA.XIR[6].XIC[8].icell.Ien VPWR.t690 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1786 XA.XIR[11].XIC[11].icell.SM XA.XIR[11].XIC[11].icell.Ien Iout.t108 VGND.t1075 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1787 XThR.Tn[7].t0 XThR.XTBN.Y.t78 VGND.t476 VGND.t475 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1788 XA.XIR[2].XIC_15.icell.SM XA.XIR[2].XIC_15.icell.Ien Iout.t161 VGND.t1293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1789 VPWR.t1486 VPWR.t1484 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1485 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1790 VGND.t2180 XThC.Tn[9].t32 XA.XIR[4].XIC[9].icell.PDM VGND.t2179 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1791 XA.XIR[14].XIC[4].icell.Ien XThR.Tn[14].t49 VPWR.t1015 VPWR.t1014 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1792 XA.XIR[7].XIC[1].icell.PUM XThC.Tn[1].t32 XA.XIR[7].XIC[1].icell.Ien VPWR.t1183 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1793 VGND.t2367 VPWR.t2013 XA.XIR[15].XIC_15.icell.PDM VGND.t2366 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1794 XThC.XTB4.Y.t0 XThC.XTB7.B VGND.t1137 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1795 VPWR.t121 XThR.XTB6.Y XThR.Tn[13].t6 VPWR.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VPWR.t647 XThR.XTB3.Y a_n1049_7493# VPWR.t646 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1797 XA.XIR[1].XIC[5].icell.PUM XThC.Tn[5].t30 XA.XIR[1].XIC[5].icell.Ien VPWR.t864 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1798 VPWR.t1152 XThR.Tn[11].t54 XA.XIR[12].XIC[12].icell.PUM VPWR.t1151 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1799 VGND.t95 Vbias.t163 XA.XIR[7].XIC[5].icell.SM VGND.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1800 XA.XIR[6].XIC[6].icell.Ien XThR.Tn[6].t50 VPWR.t1747 VPWR.t1746 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1801 XA.XIR[5].XIC[7].icell.Ien XThR.Tn[5].t49 VPWR.t64 VPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1802 VPWR.t136 data[4].t3 XThR.XTB7.A VPWR.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1803 VGND.t121 XThC.Tn[4].t33 XA.XIR[7].XIC[4].icell.PDM VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1804 VGND.t97 Vbias.t164 XA.XIR[6].XIC[6].icell.SM VGND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1805 VGND.t2369 VPWR.t2014 XA.XIR[2].XIC_dummy_right.icell.PDM VGND.t2368 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1806 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2015 VGND.t2560 VGND.t2559 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1807 XA.XIR[15].XIC[6].icell.PDM XThR.Tn[14].t50 VGND.t333 VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1808 XThC.Tn[6].t9 XThC.XTBN.Y.t80 VGND.t1437 VGND.t1436 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1809 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[13].t48 VGND.t34 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1810 XA.XIR[9].XIC[7].icell.Ien XThR.Tn[9].t45 VPWR.t343 VPWR.t342 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1811 XA.XIR[8].XIC[8].icell.Ien XThR.Tn[8].t56 VPWR.t582 VPWR.t581 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1812 VPWR.t1058 VGND.t2698 XA.XIR[0].XIC[6].icell.PUM VPWR.t1057 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1813 VPWR.t148 XThR.Tn[3].t55 XA.XIR[4].XIC[14].icell.PUM VPWR.t147 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1814 XThR.Tn[5].t1 XThR.XTB6.Y VGND.t210 VGND.t209 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1815 VPWR.t737 XThR.Tn[7].t48 XA.XIR[8].XIC[3].icell.PUM VPWR.t736 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1816 VPWR.t413 XThC.XTB5.Y a_5155_9615# VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1817 VPWR.t1483 VPWR.t1481 XA.XIR[3].XIC_15.icell.PUM VPWR.t1482 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1818 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6].t51 XA.XIR[6].XIC[9].icell.Ien VGND.t2247 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1819 VPWR.t1480 VPWR.t1478 XA.XIR[7].XIC_15.icell.PUM VPWR.t1479 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1820 VGND.t99 Vbias.t165 XA.XIR[1].XIC[3].icell.SM VGND.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1821 XA.XIR[3].XIC[11].icell.PUM XThC.Tn[11].t30 XA.XIR[3].XIC[11].icell.Ien VPWR.t292 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1822 XThR.Tn[4].t2 XThR.XTB5.Y VGND.t1164 VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1823 a_4861_9615# XThC.XTB4.Y.t13 VPWR.t1030 VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1824 a_5949_9615# XThC.XTBN.Y.t81 XThC.Tn[5].t5 VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1825 VGND.t101 Vbias.t166 XA.XIR[4].XIC[4].icell.SM VGND.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1826 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[5].t50 VGND.t81 VGND.t80 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1827 VGND.t2562 VPWR.t2016 XA.XIR[5].XIC_dummy_left.icell.PDM VGND.t2561 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1828 XA.XIR[11].XIC[9].icell.SM XA.XIR[11].XIC[9].icell.Ien Iout.t51 VGND.t373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1829 VGND.t1438 XThC.XTBN.Y.t82 XThC.Tn[2].t6 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1830 VGND.t2564 VPWR.t2017 XA.XIR[9].XIC_dummy_left.icell.PDM VGND.t2563 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1831 XA.XIR[8].XIC[11].icell.SM XA.XIR[8].XIC[11].icell.Ien Iout.t208 VGND.t2080 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1832 VPWR.t1197 XThC.XTB1.Y.t14 XThC.Tn[8].t5 VPWR.t1196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1833 VGND.t426 XThC.Tn[11].t31 XA.XIR[11].XIC[11].icell.PDM VGND.t425 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1834 a_5155_10571# XThC.XTB7.B XThC.XTB5.Y VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1835 a_10915_9569# XThC.XTBN.Y.t83 VGND.t1440 VGND.t1439 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1836 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14].t51 VPWR.t196 VPWR.t195 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1837 XA.XIR[4].XIC[1].icell.PUM XThC.Tn[1].t33 XA.XIR[4].XIC[1].icell.Ien VPWR.t1920 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1838 XA.XIR[3].XIC[2].icell.PUM XThC.Tn[2].t30 XA.XIR[3].XIC[2].icell.Ien VPWR.t1272 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1839 VPWR.t1154 XThR.Tn[11].t55 XA.XIR[12].XIC[10].icell.PUM VPWR.t1153 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1840 XA.XIR[0].XIC[5].icell.Ien XThR.Tn[0].t53 VPWR.t619 VPWR.t618 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1841 XA.XIR[6].XIC[3].icell.PUM XThC.Tn[3].t32 XA.XIR[6].XIC[3].icell.Ien VPWR.t453 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1842 VGND.t103 Vbias.t167 XA.XIR[6].XIC[10].icell.SM VGND.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1843 XA.XIR[5].XIC[11].icell.Ien XThR.Tn[5].t51 VPWR.t1813 VPWR.t1812 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1844 XThC.Tn[3].t8 XThC.XTB4.Y.t14 VGND.t1710 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1845 VGND.t105 Vbias.t168 XA.XIR[3].XIC[6].icell.SM VGND.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1846 VGND.t123 XThC.Tn[4].t34 XA.XIR[4].XIC[4].icell.PDM VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1847 VGND.t2677 XThC.Tn[1].t34 XA.XIR[8].XIC[1].icell.PDM VGND.t2676 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1848 VGND.t1234 XThC.Tn[5].t31 XA.XIR[3].XIC[5].icell.PDM VGND.t1233 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1849 XA.XIR[9].XIC[11].icell.Ien XThR.Tn[9].t46 VPWR.t345 VPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1850 VGND.t2144 XThC.Tn[2].t31 XA.XIR[11].XIC[2].icell.PDM VGND.t2143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1851 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[3].t56 VGND.t258 VGND.t257 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1852 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13].t49 XA.XIR[13].XIC[11].icell.Ien VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1853 XThR.Tn[3].t8 XThR.XTBN.Y.t79 VGND.t477 VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1854 XA.XIR[0].XIC[13].icell.PUM XThC.Tn[13].t33 XA.XIR[0].XIC[13].icell.Ien VPWR.t626 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1855 XA.XIR[6].XIC[1].icell.Ien XThR.Tn[6].t52 VPWR.t1749 VPWR.t1748 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1856 VGND.t107 Vbias.t169 XA.XIR[7].XIC[0].icell.SM VGND.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1857 VGND.t109 Vbias.t170 XA.XIR[2].XIC[12].icell.SM VGND.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1858 XA.XIR[5].XIC[2].icell.Ien XThR.Tn[5].t52 VPWR.t1815 VPWR.t1814 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1859 VGND.t111 Vbias.t171 XA.XIR[6].XIC[1].icell.SM VGND.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1860 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1476 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1477 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1861 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t1 VGND.t1304 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1862 XA.XIR[9].XIC[2].icell.Ien XThR.Tn[9].t47 VPWR.t347 VPWR.t346 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1863 a_4387_10575# XThC.XTB7.B VGND.t1135 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1864 XA.XIR[4].XIC[14].icell.Ien XThR.Tn[4].t54 VPWR.t1189 VPWR.t1188 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1865 XA.XIR[5].XIC[8].icell.SM XA.XIR[5].XIC[8].icell.Ien Iout.t194 VGND.t1915 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1866 XA.XIR[8].XIC[3].icell.Ien XThR.Tn[8].t57 VPWR.t854 VPWR.t853 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1867 VPWR.t1056 VGND.t2699 XA.XIR[0].XIC[1].icell.PUM VPWR.t1055 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1868 XA.XIR[3].XIC_15.icell.Ien XThR.Tn[3].t57 VPWR.t150 VPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1869 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10].t49 XA.XIR[10].XIC[1].icell.Ien VGND.t349 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1870 XA.XIR[8].XIC[9].icell.SM XA.XIR[8].XIC[9].icell.Ien Iout.t42 VGND.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1871 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6].t53 XA.XIR[6].XIC[4].icell.Ien VGND.t665 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1872 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t2018 XA.XIR[1].XIC_dummy_right.icell.Ien VGND.t2565 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1873 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5].t53 XA.XIR[5].XIC[5].icell.Ien VGND.t2427 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1874 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13].t50 XA.XIR[13].XIC[2].icell.Ien VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1875 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9].t48 XA.XIR[9].XIC[5].icell.Ien VGND.t507 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1876 a_10051_9569# XThC.XTBN.Y.t84 VGND.t1441 VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1877 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11].t56 XA.XIR[11].XIC_15.icell.Ien VGND.t1979 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1878 XThC.XTB1.Y.t2 XThC.XTB7.B VPWR.t741 VPWR.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1879 a_n1049_6699# XThR.XTBN.Y.t80 XThR.Tn[3].t5 VPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1880 XA.XIR[2].XIC[8].icell.SM XA.XIR[2].XIC[8].icell.Ien Iout.t210 VGND.t2088 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1881 XA.XIR[11].XIC[4].icell.SM XA.XIR[11].XIC[4].icell.Ien Iout.t109 VGND.t1076 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1882 VGND.t113 Vbias.t172 XA.XIR[3].XIC[10].icell.SM VGND.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1883 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1473 VPWR.t1475 VPWR.t1474 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1884 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout VGND.t1292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1885 a_n1049_8581# XThR.XTBN.Y.t81 XThR.Tn[0].t5 VPWR.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1886 a_7651_9569# XThC.XTBN.Y.t85 VGND.t1442 VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1887 VGND.t1819 VGND.t1817 XA.XIR[14].XIC_dummy_right.icell.SM VGND.t1818 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1888 VGND.t518 XThC.Tn[6].t33 XA.XIR[11].XIC[6].icell.PDM VGND.t517 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1889 VPWR.t1855 XThC.XTB7.A a_6243_10571# VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1890 VPWR.t1472 VPWR.t1470 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1471 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1891 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[0].t54 VGND.t812 VGND.t811 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1892 VPWR.t1142 XThR.Tn[11].t57 XA.XIR[12].XIC[5].icell.PUM VPWR.t1141 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1893 XThC.Tn[10].t3 XThC.XTB3.Y.t13 a_8739_9569# VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1894 VGND.t1364 Vbias.t173 XA.XIR[3].XIC[1].icell.SM VGND.t1363 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1895 XA.XIR[7].XIC[5].icell.SM XA.XIR[7].XIC[5].icell.Ien Iout.t47 VGND.t268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1896 VGND.t951 XThC.Tn[0].t31 XA.XIR[3].XIC[0].icell.PDM VGND.t950 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1897 VGND.t375 XThR.XTBN.Y.t82 XThR.Tn[2].t1 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1898 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[10].t50 VGND.t1089 VGND.t1088 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1899 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[10].t51 VGND.t1091 VGND.t1090 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1900 XA.XIR[10].XIC[6].icell.SM XA.XIR[10].XIC[6].icell.Ien Iout.t231 VGND.t2387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1901 XThR.XTB5.A data[5].t3 VGND.t1170 VGND.t1169 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1902 XA.XIR[14].XIC[14].icell.SM XA.XIR[14].XIC[14].icell.Ien Iout.t125 VGND.t1131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1903 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1468 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1469 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1904 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[3].t58 VGND.t260 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1905 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7].t49 XA.XIR[7].XIC[1].icell.Ien VGND.t1118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1906 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13].t51 XA.XIR[13].XIC[6].icell.Ien VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1907 XThR.Tn[12].t9 XThR.XTBN.Y.t83 VPWR.t236 VPWR.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1908 VGND.t2567 VPWR.t2019 XA.XIR[14].XIC_dummy_right.icell.PDM VGND.t2566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1909 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[6].t54 VGND.t667 VGND.t666 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1910 XA.XIR[5].XIC[8].icell.PUM XThC.Tn[8].t32 XA.XIR[5].XIC[8].icell.Ien VPWR.t691 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1911 XThR.Tn[12].t1 XThR.XTB5.Y a_n997_1803# VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1912 XA.XIR[1].XIC_15.icell.SM XA.XIR[1].XIC_15.icell.Ien Iout.t181 VGND.t1520 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1913 XA.XIR[9].XIC[8].icell.PUM XThC.Tn[8].t33 XA.XIR[9].XIC[8].icell.Ien VPWR.t692 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1914 XThR.Tn[3].t1 XThR.XTB4.Y VGND.t653 VGND.t652 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1915 XA.XIR[5].XIC[3].icell.SM XA.XIR[5].XIC[3].icell.Ien Iout.t120 VGND.t1126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1916 VGND.t377 XThR.XTBN.Y.t84 a_n997_2667# VGND.t376 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1917 XA.XIR[9].XIC_15.icell.PDM VPWR.t2020 VGND.t2569 VGND.t2568 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1918 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5].t54 XA.XIR[5].XIC[0].icell.Ien VGND.t2428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1919 XA.XIR[8].XIC[4].icell.SM XA.XIR[8].XIC[4].icell.Ien Iout.t92 VGND.t877 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1920 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout VGND.t764 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1921 VGND.t1366 Vbias.t174 XA.XIR[13].XIC_15.icell.SM VGND.t1365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1922 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1465 VPWR.t1467 VPWR.t1466 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1923 XA.XIR[0].XIC[6].icell.PUM XThC.Tn[6].t34 XA.XIR[0].XIC[6].icell.Ien VPWR.t352 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1924 VGND.t1081 XThC.Tn[14].t32 XA.XIR[13].XIC[14].icell.PDM VGND.t1080 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1925 VGND.t1050 XThC.Tn[8].t34 XA.XIR[13].XIC[8].icell.PDM VGND.t1049 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1926 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9].t49 XA.XIR[9].XIC[0].icell.Ien VGND.t508 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1927 a_5155_9615# XThC.XTB5.Y VPWR.t412 VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1928 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[4].t55 XA.XIR[4].XIC[12].icell.Ien VGND.t2071 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1929 VPWR.t411 XThC.XTB5.Y XThC.Tn[12].t4 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1930 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[3].t59 XA.XIR[3].XIC[13].icell.Ien VGND.t261 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1931 VPWR.t198 XThR.Tn[14].t52 XA.XIR[15].XIC[12].icell.PUM VPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1932 XA.XIR[7].XIC_15.icell.PUM VPWR.t1463 XA.XIR[7].XIC_15.icell.Ien VPWR.t1464 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1933 VPWR.t32 XThR.Tn[13].t52 XA.XIR[14].XIC[13].icell.PUM VPWR.t31 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1934 VPWR.t1462 VPWR.t1460 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1461 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1935 VGND.t2182 XThC.Tn[9].t33 XA.XIR[0].XIC[9].icell.PDM VGND.t2181 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1936 XThC.Tn[5].t4 XThC.XTBN.Y.t86 a_5949_9615# VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1937 XA.XIR[2].XIC[3].icell.SM XA.XIR[2].XIC[3].icell.Ien Iout.t252 VGND.t2648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1938 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[7].t50 VGND.t1120 VGND.t1119 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1939 VGND.t564 XThC.XTB5.Y XThC.Tn[4].t0 VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1940 a_n1049_6405# XThR.XTBN.Y.t85 XThR.Tn[4].t5 VPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1941 VPWR.t510 XThR.Tn[1].t49 XA.XIR[2].XIC[7].icell.PUM VPWR.t509 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1942 VPWR.t621 XThR.Tn[0].t55 XA.XIR[1].XIC[8].icell.PUM VPWR.t620 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1943 XA.XIR[10].XIC[10].icell.SM XA.XIR[10].XIC[10].icell.Ien Iout.t158 VGND.t1289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1944 XThC.Tn[2].t5 XThC.XTBN.Y.t87 VGND.t365 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1945 VPWR.t1191 XThR.Tn[4].t56 XA.XIR[5].XIC[8].icell.PUM VPWR.t1190 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1946 XA.XIR[15].XIC[14].icell.PDM VPWR.t2021 XA.XIR[15].XIC[14].icell.Ien VGND.t2570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1947 XA.XIR[15].XIC[8].icell.PDM VPWR.t2022 XA.XIR[15].XIC[8].icell.Ien VGND.t2571 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1948 a_5155_9615# XThC.XTBN.Y.t88 XThC.Tn[4].t5 VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1949 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[0].t56 VGND.t814 VGND.t813 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1950 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[7].t51 VGND.t1122 VGND.t1121 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1951 XA.XIR[13].XIC[9].icell.PUM XThC.Tn[9].t34 XA.XIR[13].XIC[9].icell.Ien VPWR.t1302 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1952 XA.XIR[7].XIC[0].icell.SM XA.XIR[7].XIC[0].icell.Ien Iout.t56 VGND.t495 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1953 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout VGND.t1077 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1954 VPWR.t1099 XThR.XTB7.B XThR.XTB2.Y VPWR.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1955 XThC.Tn[8].t0 XThC.XTB1.Y.t15 a_7651_9569# VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1956 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[10].t52 VGND.t1093 VGND.t1092 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1957 VGND.t428 XThC.Tn[11].t32 XA.XIR[10].XIC[11].icell.PDM VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1958 XA.XIR[10].XIC[1].icell.SM XA.XIR[10].XIC[1].icell.Ien Iout.t65 VGND.t618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1959 XA.XIR[6].XIC_15.icell.PDM VPWR.t2023 VGND.t2573 VGND.t2572 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1960 VGND.t749 XThC.XTB5.A XThC.XTB5.Y VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1961 VGND.t1816 VGND.t1814 XA.XIR[14].XIC_dummy_left.icell.SM VGND.t1815 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1962 VGND.t1548 XThR.XTB7.Y XThR.Tn[6].t0 VGND.t1547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1963 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[4].t57 XA.XIR[4].XIC[10].icell.Ien VGND.t1953 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1964 XA.XIR[1].XIC[14].icell.PUM XThC.Tn[14].t33 XA.XIR[1].XIC[14].icell.Ien VPWR.t701 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1965 XA.XIR[5].XIC[3].icell.PUM XThC.Tn[3].t33 XA.XIR[5].XIC[3].icell.Ien VPWR.t454 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1966 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[6].t55 VGND.t669 VGND.t668 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1967 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[1].t50 VGND.t705 VGND.t704 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1968 VPWR.t200 XThR.Tn[14].t53 XA.XIR[15].XIC[10].icell.PUM VPWR.t199 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1969 XA.XIR[9].XIC[3].icell.PUM XThC.Tn[3].t34 XA.XIR[9].XIC[3].icell.Ien VPWR.t455 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1970 XA.XIR[4].XIC_15.icell.PUM VPWR.t1458 XA.XIR[4].XIC_15.icell.Ien VPWR.t1459 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1971 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[4].t58 VGND.t1955 VGND.t1954 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1972 XA.XIR[4].XIC[11].icell.SM XA.XIR[4].XIC[11].icell.Ien Iout.t145 VGND.t1212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1973 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2024 VGND.t2575 VGND.t2574 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1974 XA.XIR[15].XIC[9].icell.Ien VPWR.t1455 VPWR.t1457 VPWR.t1456 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1975 VGND.t2146 XThC.Tn[2].t32 XA.XIR[10].XIC[2].icell.PDM VGND.t2145 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1976 XThR.Tn[9].t8 XThR.XTBN.Y.t86 VPWR.t238 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1977 VGND.t367 XThC.XTBN.Y.t89 a_9827_9569# VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1978 XA.XIR[0].XIC[1].icell.PUM XThC.Tn[1].t35 XA.XIR[0].XIC[1].icell.Ien VPWR.t1921 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1979 VPWR.t512 XThR.Tn[1].t51 XA.XIR[2].XIC[11].icell.PUM VPWR.t511 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1980 VGND.t224 XThC.Tn[3].t35 XA.XIR[13].XIC[3].icell.PDM VGND.t223 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1981 VGND.t2577 VPWR.t2025 XA.XIR[8].XIC_15.icell.PDM VGND.t2576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1982 VPWR.t856 XThR.Tn[8].t58 XA.XIR[9].XIC[9].icell.PUM VPWR.t855 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1983 VGND.t1368 Vbias.t175 XA.XIR[1].XIC[12].icell.SM VGND.t1367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1984 XA.XIR[14].XIC[13].icell.Ien XThR.Tn[14].t54 VPWR.t202 VPWR.t201 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1985 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1452 VPWR.t1454 VPWR.t1453 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1986 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12].t53 XA.XIR[12].XIC[14].icell.Ien VGND.t2112 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1987 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1450 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1451 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1988 XThC.Tn[0].t11 XThC.XTB1.Y.t16 VGND.t2074 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1989 VGND.t1370 Vbias.t176 XA.XIR[0].XIC[5].icell.SM VGND.t1369 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1990 VGND.t1372 Vbias.t177 XA.XIR[4].XIC[13].icell.SM VGND.t1371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1991 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12].t54 XA.XIR[12].XIC[8].icell.Ien VGND.t2113 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1992 VGND.t125 XThC.Tn[4].t35 XA.XIR[0].XIC[4].icell.PDM VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1993 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t0 VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1994 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[7].t52 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1995 XA.XIR[2].XIC[7].icell.Ien XThR.Tn[2].t49 VPWR.t792 VPWR.t791 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1996 VGND.t1374 Vbias.t178 XA.XIR[7].XIC[14].icell.SM VGND.t1373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1997 XA.XIR[6].XIC_15.icell.Ien XThR.Tn[6].t56 VPWR.t486 VPWR.t485 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1998 VPWR.t514 XThR.Tn[1].t52 XA.XIR[2].XIC[2].icell.PUM VPWR.t513 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1999 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[10].t53 VGND.t1095 VGND.t1094 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2000 VGND.t846 XThC.Tn[13].t34 XA.XIR[7].XIC[13].icell.PDM VGND.t845 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2001 VPWR.t958 XThR.Tn[0].t57 XA.XIR[1].XIC[3].icell.PUM VPWR.t957 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2002 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout VGND.t556 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2003 XThR.Tn[14].t9 XThR.XTBN.Y.t87 VPWR.t240 VPWR.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2004 VPWR.t1122 XThR.Tn[4].t59 XA.XIR[5].XIC[3].icell.PUM VPWR.t1121 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2005 VPWR.t1449 VPWR.t1447 XA.XIR[0].XIC_15.icell.PUM VPWR.t1448 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2006 VPWR.t34 XThR.Tn[13].t53 XA.XIR[14].XIC[6].icell.PUM VPWR.t33 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2007 XA.XIR[15].XIC[3].icell.PDM VPWR.t2026 XA.XIR[15].XIC[3].icell.Ien VGND.t2578 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2008 a_n997_3755# XThR.XTBN.Y.t88 VGND.t379 VGND.t378 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2009 XThR.Tn[8].t5 XThR.XTB1.Y VPWR.t1085 VPWR.t1084 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2010 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10].t54 XA.XIR[10].XIC_15.icell.Ien VGND.t1096 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2011 XA.XIR[0].XIC[14].icell.Ien XThR.Tn[0].t58 VPWR.t960 VPWR.t959 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2012 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[1].t53 VGND.t251 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2013 XA.XIR[1].XIC[8].icell.SM XA.XIR[1].XIC[8].icell.Ien Iout.t147 VGND.t1216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2014 VGND.t1376 Vbias.t179 XA.XIR[10].XIC[7].icell.SM VGND.t1375 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2015 a_n1049_7787# XThR.XTB2.Y VPWR.t925 VPWR.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2016 XA.XIR[4].XIC[9].icell.SM XA.XIR[4].XIC[9].icell.Ien Iout.t190 VGND.t1708 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2017 VGND.t520 XThC.Tn[6].t35 XA.XIR[10].XIC[6].icell.PDM VGND.t519 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2018 VPWR.t1241 XThR.Tn[12].t55 XA.XIR[13].XIC[4].icell.PUM VPWR.t1240 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2019 a_n1331_2891# data[5].t4 VGND.t320 VGND.t319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2020 VGND.t1378 Vbias.t180 XA.XIR[13].XIC[8].icell.SM VGND.t1377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2021 XA.XIR[12].XIC[9].icell.Ien XThR.Tn[12].t56 VPWR.t1243 VPWR.t1242 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2022 VPWR.t1446 VPWR.t1444 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1445 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2023 VGND.t1207 XThC.Tn[7].t27 XA.XIR[13].XIC[7].icell.PDM VGND.t1206 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2024 VPWR.t204 XThR.Tn[14].t55 XA.XIR[15].XIC[5].icell.PUM VPWR.t203 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2025 XThR.XTB7.B data[6].t1 VGND.t763 VGND.t762 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2026 XThR.Tn[2].t2 XThR.XTBN.Y.t89 a_n1049_7493# VPWR.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2027 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[9].t50 VGND.t524 VGND.t523 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2028 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[9].t51 VGND.t526 VGND.t525 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2029 XA.XIR[2].XIC[11].icell.Ien XThR.Tn[2].t50 VPWR.t790 VPWR.t789 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2030 XA.XIR[9].XIC[6].icell.SM XA.XIR[9].XIC[6].icell.Ien Iout.t211 VGND.t2089 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2031 VGND.t2549 XThC.Tn[12].t34 XA.XIR[1].XIC[12].icell.PDM VGND.t2548 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2032 VGND.t848 XThC.Tn[13].t35 XA.XIR[4].XIC[13].icell.PDM VGND.t847 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2033 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t2027 XA.XIR[4].XIC_dummy_left.icell.Ien VGND.t2579 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2034 XA.XIR[15].XIC[7].icell.PDM VPWR.t2028 XA.XIR[15].XIC[7].icell.Ien VGND.t2580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2035 VGND.t1380 Vbias.t181 XA.XIR[0].XIC[0].icell.SM VGND.t1379 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2036 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12].t57 XA.XIR[12].XIC[3].icell.Ien VGND.t2114 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2037 VPWR.t231 XThC.XTBN.Y.t90 XThC.Tn[8].t10 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2038 XThR.Tn[10].t5 XThR.XTB3.Y VPWR.t645 VPWR.t644 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2039 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7].t53 XA.XIR[7].XIC_15.icell.Ien VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2040 XA.XIR[11].XIC[4].icell.PUM XThC.Tn[4].t36 XA.XIR[11].XIC[4].icell.Ien VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2041 XThR.Tn[4].t9 XThR.XTBN.Y.t90 VGND.t381 VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2042 XA.XIR[15].XIC[12].icell.PUM XThC.Tn[12].t35 XA.XIR[15].XIC[12].icell.Ien VPWR.t1886 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2043 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1442 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1443 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2044 XA.XIR[2].XIC[2].icell.Ien XThR.Tn[2].t51 VPWR.t788 VPWR.t787 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2045 XA.XIR[11].XIC[13].icell.SM XA.XIR[11].XIC[13].icell.Ien Iout.t246 VGND.t2488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2046 VGND.t1921 XThR.XTB7.B XThR.XTB5.Y VGND.t1920 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2047 VGND.t1382 Vbias.t182 XA.XIR[12].XIC_15.icell.SM VGND.t1381 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2048 VGND.t1083 XThC.Tn[14].t34 XA.XIR[12].XIC[14].icell.PDM VGND.t1082 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2049 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[3].t60 XA.XIR[3].XIC[1].icell.Ien VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2050 XA.XIR[14].XIC[6].icell.Ien XThR.Tn[14].t56 VPWR.t206 VPWR.t205 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2051 VGND.t1052 XThC.Tn[8].t35 XA.XIR[12].XIC[8].icell.PDM VGND.t1051 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2052 VPWR.t1785 XThR.Tn[13].t54 XA.XIR[14].XIC[1].icell.PUM VPWR.t1784 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2053 XA.XIR[2].XIC[7].icell.PUM XThC.Tn[7].t28 XA.XIR[2].XIC[7].icell.Ien VPWR.t502 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2054 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[2].t52 XA.XIR[2].XIC[5].icell.Ien VGND.t1062 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2055 VPWR.t1245 XThR.Tn[12].t58 XA.XIR[13].XIC[0].icell.PUM VPWR.t1244 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2056 VPWR.t356 XThR.Tn[9].t52 XA.XIR[10].XIC[4].icell.PUM VPWR.t355 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2057 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6].t57 XA.XIR[6].XIC[13].icell.Ien VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2058 XA.XIR[1].XIC[3].icell.SM XA.XIR[1].XIC[3].icell.Ien Iout.t44 VGND.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2059 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14].t57 XA.XIR[14].XIC[9].icell.Ien VGND.t334 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2060 VPWR.t1144 XThR.Tn[11].t58 XA.XIR[12].XIC[14].icell.PUM VPWR.t1143 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2061 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t1 VGND.t1396 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2062 XThC.Tn[4].t4 XThC.XTBN.Y.t91 a_5155_9615# VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2063 XA.XIR[13].XIC[4].icell.Ien XThR.Tn[13].t55 VPWR.t1787 VPWR.t1786 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2064 VGND.t1384 Vbias.t183 XA.XIR[10].XIC[2].icell.SM VGND.t1383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2065 XA.XIR[4].XIC[4].icell.SM XA.XIR[4].XIC[4].icell.Ien Iout.t200 VGND.t1940 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2066 VGND.t1386 Vbias.t184 XA.XIR[9].XIC_15.icell.SM VGND.t1385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2067 XA.XIR[9].XIC[10].icell.SM XA.XIR[9].XIC[10].icell.Ien Iout.t37 VGND.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2068 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1439 VPWR.t1441 VPWR.t1440 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2069 VGND.t2194 XThC.Tn[10].t35 XA.XIR[1].XIC[10].icell.PDM VGND.t2193 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2070 VGND.t957 Vbias.t185 XA.XIR[13].XIC[3].icell.SM VGND.t956 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2071 XA.XIR[0].XIC[12].icell.PDM XThR.Tn[0].t59 XA.XIR[0].XIC[12].icell.Ien VGND.t1494 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2072 VPWR.t152 XThR.Tn[3].t61 XA.XIR[4].XIC[8].icell.PUM VPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2073 VGND.t382 XThR.XTBN.Y.t91 a_n997_1579# VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2074 VPWR.t703 XThR.Tn[10].t55 XA.XIR[11].XIC[12].icell.PUM VPWR.t702 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2075 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2029 VGND.t2582 VGND.t2581 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2076 XA.XIR[12].XIC[9].icell.PUM XThC.Tn[9].t35 XA.XIR[12].XIC[9].icell.Ien VPWR.t1303 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2077 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12].t59 XA.XIR[12].XIC[7].icell.Ien VGND.t2115 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2078 XA.XIR[15].XIC[10].icell.PUM XThC.Tn[10].t36 XA.XIR[15].XIC[10].icell.Ien VPWR.t1306 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2079 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[9].t53 VGND.t528 VGND.t527 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2080 XA.XIR[5].XIC[12].icell.SM XA.XIR[5].XIC[12].icell.Ien Iout.t230 VGND.t2386 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2081 XA.XIR[9].XIC[1].icell.SM XA.XIR[9].XIC[1].icell.Ien Iout.t165 VGND.t1388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2082 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t1 VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2083 XA.XIR[11].XIC[0].icell.PUM XThC.Tn[0].t32 XA.XIR[11].XIC[0].icell.Ien VPWR.t677 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2084 XA.XIR[8].XIC[13].icell.SM XA.XIR[8].XIC[13].icell.Ien Iout.t17 VGND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2085 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1437 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1438 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2086 XA.XIR[7].XIC[14].icell.SM XA.XIR[7].XIC[14].icell.Ien Iout.t21 VGND.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2087 XA.XIR[2].XIC[11].icell.PUM XThC.Tn[11].t33 XA.XIR[2].XIC[11].icell.Ien VPWR.t293 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2088 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[4].t60 VGND.t1957 VGND.t1956 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2089 XA.XIR[0].XIC[5].icell.PDM VGND.t1811 VGND.t1813 VGND.t1812 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2090 VPWR.t358 XThR.Tn[9].t54 XA.XIR[10].XIC[0].icell.PUM VPWR.t357 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2091 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[3].t62 VGND.t264 VGND.t263 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2092 XA.XIR[2].XIC[12].icell.SM XA.XIR[2].XIC[12].icell.Ien Iout.t149 VGND.t1223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2093 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[11].t59 VGND.t1969 VGND.t1968 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2094 VGND.t226 XThC.Tn[3].t36 XA.XIR[12].XIC[3].icell.PDM VGND.t225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2095 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14].t58 VPWR.t208 VPWR.t207 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2096 XThR.XTBN.Y.t2 XThR.XTBN.A VPWR.t190 VPWR.t189 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2097 VGND.t959 Vbias.t186 XA.XIR[15].XIC[11].icell.SM VGND.t958 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2098 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13].t56 VPWR.t1789 VPWR.t1788 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2099 VPWR.t1 XThR.Tn[7].t54 XA.XIR[8].XIC[9].icell.PUM VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2100 VGND.t1085 XThC.Tn[14].t35 XA.XIR[6].XIC[14].icell.PDM VGND.t1084 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2101 XA.XIR[0].XIC[10].icell.PDM XThR.Tn[0].t60 XA.XIR[0].XIC[10].icell.Ien VGND.t1495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2102 XA.XIR[2].XIC[2].icell.PUM XThC.Tn[2].t33 XA.XIR[2].XIC[2].icell.Ien VPWR.t1273 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2103 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[2].t53 XA.XIR[2].XIC[0].icell.Ien VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2104 VGND.t1054 XThC.Tn[8].t36 XA.XIR[6].XIC[8].icell.PDM VGND.t1053 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2105 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1434 VPWR.t1436 VPWR.t1435 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2106 VPWR.t705 XThR.Tn[10].t56 XA.XIR[11].XIC[10].icell.PUM VPWR.t704 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2107 XA.XIR[0].XIC_15.icell.PUM VPWR.t1432 XA.XIR[0].XIC_15.icell.Ien VPWR.t1433 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2108 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14].t59 XA.XIR[14].XIC[4].icell.Ien VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2109 XA.XIR[1].XIC[7].icell.Ien XThR.Tn[1].t54 VPWR.t142 VPWR.t141 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2110 VGND.t961 Vbias.t187 XA.XIR[2].XIC[6].icell.SM VGND.t960 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2111 VGND.t2679 XThC.Tn[1].t36 XA.XIR[7].XIC[1].icell.PDM VGND.t2678 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2112 VGND.t1236 XThC.Tn[5].t32 XA.XIR[2].XIC[5].icell.PDM VGND.t1235 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2113 VPWR.t242 XThR.XTBN.Y.t92 XThR.Tn[11].t9 VPWR.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2114 XA.XIR[4].XIC[8].icell.Ien XThR.Tn[4].t61 VPWR.t1124 VPWR.t1123 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2115 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[9].t55 VGND.t530 VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2116 VPWR.t160 data[1].t4 XThC.XTB7.A VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2117 VPWR.t154 XThR.Tn[3].t63 XA.XIR[4].XIC[3].icell.PUM VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2118 XA.XIR[11].XIC[12].icell.Ien XThR.Tn[11].t60 VPWR.t1146 VPWR.t1145 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2119 a_8739_9569# XThC.XTBN.Y.t92 VGND.t368 VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2120 VGND.t327 XThR.XTBN.A XThR.XTBN.Y.t0 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 XThC.Tn[6].t2 XThC.XTB7.Y VGND.t1303 VGND.t1302 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2122 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8].t59 XA.XIR[8].XIC[14].icell.Ien VGND.t1219 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2123 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8].t60 XA.XIR[8].XIC[8].icell.Ien VGND.t1220 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2124 XA.XIR[15].XIC[5].icell.PUM XThC.Tn[5].t33 XA.XIR[15].XIC[5].icell.Ien VPWR.t865 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2125 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[0].t61 VGND.t1497 VGND.t1496 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2126 XA.XIR[6].XIC[9].icell.PUM XThC.Tn[9].t36 XA.XIR[6].XIC[9].icell.Ien VPWR.t1262 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2127 XThR.Tn[12].t0 XThR.XTB5.Y a_n997_1803# VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2128 VGND.t2584 VPWR.t2030 XA.XIR[1].XIC_dummy_left.icell.PDM VGND.t2583 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2129 VGND.t963 Vbias.t188 XA.XIR[12].XIC[8].icell.SM VGND.t962 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2130 VGND.t430 XThC.Tn[11].t34 XA.XIR[3].XIC[11].icell.PDM VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2131 VGND.t684 XThC.Tn[7].t29 XA.XIR[12].XIC[7].icell.PDM VGND.t683 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2132 VGND.t965 Vbias.t189 XA.XIR[15].XIC[9].icell.SM VGND.t964 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2133 a_n997_3979# XThR.XTBN.Y.t93 VGND.t384 VGND.t383 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2134 XThC.XTB7.Y XThC.XTB7.B VGND.t1134 VGND.t1133 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2135 XA.XIR[0].XIC[0].icell.PDM VGND.t1808 VGND.t1810 VGND.t1809 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2136 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1429 VPWR.t1431 VPWR.t1430 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2137 VGND.t967 Vbias.t190 XA.XIR[6].XIC[7].icell.SM VGND.t966 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2138 XA.XIR[1].XIC[11].icell.Ien XThR.Tn[1].t55 VPWR.t144 VPWR.t143 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2139 VGND.t969 Vbias.t191 XA.XIR[2].XIC[10].icell.SM VGND.t968 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2140 XThC.Tn[8].t9 XThC.XTBN.Y.t93 VPWR.t233 VPWR.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2141 VGND.t2681 XThC.Tn[1].t37 XA.XIR[4].XIC[1].icell.PDM VGND.t2680 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2142 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[11].t61 VGND.t1971 VGND.t1970 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2143 VGND.t2148 XThC.Tn[2].t34 XA.XIR[3].XIC[2].icell.PDM VGND.t2147 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2144 VGND.t971 Vbias.t192 XA.XIR[9].XIC[8].icell.SM VGND.t970 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2145 XA.XIR[14].XIC[7].icell.PUM XThC.Tn[7].t30 XA.XIR[14].XIC[7].icell.Ien VPWR.t503 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2146 XA.XIR[8].XIC[9].icell.Ien XThR.Tn[8].t61 VPWR.t858 VPWR.t857 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2147 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t2031 VGND.t2586 VGND.t2585 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2148 VGND.t228 XThC.Tn[3].t37 XA.XIR[6].XIC[3].icell.PDM VGND.t227 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2149 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5].t55 XA.XIR[5].XIC[11].icell.Ien VGND.t2429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2150 XA.XIR[11].XIC[10].icell.Ien XThR.Tn[11].t62 VPWR.t1148 VPWR.t1147 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2151 a_n1049_6699# XThR.XTB4.Y VPWR.t466 VPWR.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2152 XA.XIR[13].XIC_15.icell.SM XA.XIR[13].XIC_15.icell.Ien Iout.t23 VGND.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2153 VPWR.t707 XThR.Tn[10].t57 XA.XIR[11].XIC[5].icell.PUM VPWR.t706 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2154 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9].t56 XA.XIR[9].XIC[11].icell.Ien VGND.t531 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2155 XA.XIR[10].XIC[4].icell.PUM XThC.Tn[4].t37 XA.XIR[10].XIC[4].icell.Ien VPWR.t76 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2156 XA.XIR[1].XIC[2].icell.Ien XThR.Tn[1].t56 VPWR.t146 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2157 VGND.t973 Vbias.t193 XA.XIR[2].XIC[1].icell.SM VGND.t972 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2158 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1427 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1428 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2159 XA.XIR[6].XIC[5].icell.SM XA.XIR[6].XIC[5].icell.Ien Iout.t186 VGND.t1579 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2160 VGND.t953 XThC.Tn[0].t33 XA.XIR[2].XIC[0].icell.PDM VGND.t952 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2161 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1425 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1426 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2162 XA.XIR[4].XIC[3].icell.Ien XThR.Tn[4].t62 VPWR.t1126 VPWR.t1125 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2163 VGND.t975 Vbias.t194 XA.XIR[0].XIC[14].icell.SM VGND.t974 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2164 VGND.t977 Vbias.t195 XA.XIR[14].XIC[5].icell.SM VGND.t976 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2165 VGND.t850 XThC.Tn[13].t36 XA.XIR[0].XIC[13].icell.PDM VGND.t849 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2166 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6].t58 XA.XIR[6].XIC[1].icell.Ien VGND.t671 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2167 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t2032 XA.XIR[0].XIC_dummy_left.icell.Ien VGND.t2587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2168 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[1].t57 XA.XIR[1].XIC[5].icell.Ien VGND.t252 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2169 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5].t56 XA.XIR[5].XIC[2].icell.Ien VGND.t2430 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2170 VGND.t2589 VPWR.t2033 XA.XIR[13].XIC_dummy_right.icell.PDM VGND.t2588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2171 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9].t57 XA.XIR[9].XIC[2].icell.Ien VGND.t532 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2172 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8].t62 XA.XIR[8].XIC[3].icell.Ien VGND.t1221 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2173 XA.XIR[3].XIC_15.icell.PDM XThR.Tn[3].t64 XA.XIR[3].XIC_15.icell.Ien VGND.t265 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2174 VGND.t1168 data[1].t5 XThC.XTB6.A VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2175 VPWR.t210 XThR.Tn[14].t60 XA.XIR[15].XIC[14].icell.PUM VPWR.t209 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2176 VPWR.t1424 VPWR.t1422 XA.XIR[14].XIC_15.icell.PUM VPWR.t1423 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2177 a_n997_2891# XThR.XTBN.Y.t94 VGND.t386 VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2178 VGND.t979 Vbias.t196 XA.XIR[12].XIC[3].icell.SM VGND.t978 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2179 VGND.t886 Vbias.t197 XA.XIR[3].XIC[7].icell.SM VGND.t885 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2180 VGND.t522 XThC.Tn[6].t36 XA.XIR[3].XIC[6].icell.PDM VGND.t521 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2181 XA.XIR[14].XIC[11].icell.PUM XThC.Tn[11].t35 XA.XIR[14].XIC[11].icell.Ien VPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2182 VPWR.t1817 XThR.Tn[5].t57 XA.XIR[6].XIC[4].icell.PUM VPWR.t1816 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2183 VPWR.t1421 VPWR.t1419 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1420 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2184 VGND.t888 Vbias.t198 XA.XIR[15].XIC[4].icell.SM VGND.t887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2185 VGND.t1807 VGND.t1805 XA.XIR[10].XIC_dummy_right.icell.SM VGND.t1806 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2186 VGND.t686 XThC.Tn[7].t31 XA.XIR[6].XIC[7].icell.PDM VGND.t685 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2187 VPWR.t1418 VPWR.t1416 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1417 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2188 VPWR.t1247 XThR.Tn[12].t60 XA.XIR[13].XIC[13].icell.PUM VPWR.t1246 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2189 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t2034 XA.XIR[15].XIC_dummy_right.icell.Ien VGND.t2590 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2190 XThR.Tn[11].t1 XThR.XTB4.Y a_n997_2667# VGND.t651 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2191 VGND.t890 Vbias.t199 XA.XIR[6].XIC[2].icell.SM VGND.t889 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2192 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[6].t59 VGND.t673 VGND.t672 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2193 VPWR.t409 XThC.XTB5.Y a_5155_9615# VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2194 XA.XIR[10].XIC[0].icell.PUM XThC.Tn[0].t34 XA.XIR[10].XIC[0].icell.Ien VPWR.t678 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2195 XA.XIR[3].XIC[5].icell.SM XA.XIR[3].XIC[5].icell.Ien Iout.t58 VGND.t498 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2196 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[2].t54 VGND.t1072 VGND.t1071 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2197 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[2].t55 VGND.t1070 VGND.t1069 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2198 VGND.t892 Vbias.t200 XA.XIR[9].XIC[3].icell.SM VGND.t891 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2199 XA.XIR[14].XIC[2].icell.PUM XThC.Tn[2].t35 XA.XIR[14].XIC[2].icell.Ien VPWR.t1274 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2200 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5].t58 XA.XIR[5].XIC[6].icell.Ien VGND.t2431 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2201 XA.XIR[11].XIC[5].icell.Ien XThR.Tn[11].t63 VPWR.t1150 VPWR.t1149 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2202 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[3].t65 VGND.t535 VGND.t534 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2203 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9].t58 XA.XIR[9].XIC[6].icell.Ien VGND.t533 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2204 VGND.t1238 XThC.Tn[5].t34 XA.XIR[14].XIC[5].icell.PDM VGND.t1237 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2205 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8].t63 XA.XIR[8].XIC[7].icell.Ien VGND.t1222 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2206 VGND.t435 XThR.XTBN.Y.t95 XThR.Tn[0].t9 VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2207 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[6].t60 VGND.t675 VGND.t674 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2208 XA.XIR[1].XIC[8].icell.PUM XThC.Tn[8].t37 XA.XIR[1].XIC[8].icell.Ien VPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2209 a_n1049_6405# XThR.XTB5.Y VPWR.t749 VPWR.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2210 XA.XIR[6].XIC[0].icell.SM XA.XIR[6].XIC[0].icell.Ien Iout.t176 VGND.t1492 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2211 XThR.Tn[8].t4 XThR.XTB1.Y VPWR.t1083 VPWR.t1082 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2212 XA.XIR[1].XIC[12].icell.SM XA.XIR[1].XIC[12].icell.Ien Iout.t189 VGND.t1603 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2213 XA.XIR[8].XIC[12].icell.PUM XThC.Tn[12].t36 XA.XIR[8].XIC[12].icell.Ien VPWR.t1887 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2214 VGND.t894 Vbias.t201 XA.XIR[14].XIC[0].icell.SM VGND.t893 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2215 XA.XIR[15].XIC[9].icell.PDM XThR.Tn[14].t61 VGND.t337 VGND.t336 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2216 XA.XIR[4].XIC[13].icell.SM XA.XIR[4].XIC[13].icell.Ien Iout.t13 VGND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2217 XA.XIR[5].XIC_15.icell.PDM VPWR.t2035 VGND.t2592 VGND.t2591 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2218 VGND.t896 Vbias.t202 XA.XIR[5].XIC_15.icell.SM VGND.t895 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2219 XA.XIR[11].XIC[13].icell.PUM XThC.Tn[13].t37 XA.XIR[11].XIC[13].icell.Ien VPWR.t627 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2220 VGND.t312 XThC.Tn[8].t38 XA.XIR[5].XIC[8].icell.PDM VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2221 VGND.t1087 XThC.Tn[14].t36 XA.XIR[5].XIC[14].icell.PDM VGND.t1086 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2222 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[1].t58 XA.XIR[1].XIC[0].icell.Ien VGND.t253 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2223 VGND.t898 Vbias.t203 XA.XIR[13].XIC[12].icell.SM VGND.t897 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2224 XThR.Tn[1].t1 XThR.XTB2.Y VGND.t1395 VGND.t1394 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2225 VGND.t1944 XThC.Tn[14].t37 XA.XIR[9].XIC[14].icell.PDM VGND.t1943 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2226 VGND.t314 XThC.Tn[8].t39 XA.XIR[9].XIC[8].icell.PDM VGND.t313 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2227 VPWR.t1819 XThR.Tn[5].t59 XA.XIR[6].XIC[0].icell.PUM VPWR.t1818 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2228 VGND.t369 XThC.XTBN.Y.t94 a_8739_9569# VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2229 XA.XIR[14].XIC_15.icell.Ien XThR.Tn[14].t62 VPWR.t212 VPWR.t211 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2230 VGND.t900 Vbias.t204 XA.XIR[1].XIC[6].icell.SM VGND.t899 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2231 VPWR.t1415 VPWR.t1413 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1414 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2232 XThC.Tn[1].t2 XThC.XTB2.Y VGND.t67 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2233 VGND.t1301 XThC.XTB7.Y XThC.Tn[6].t1 VGND.t1300 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2234 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t2036 XA.XIR[12].XIC_dummy_right.icell.Ien VGND.t2593 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2235 VPWR.t360 XThR.Tn[9].t59 XA.XIR[10].XIC[13].icell.PUM VPWR.t359 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2236 VPWR.t1412 VPWR.t1410 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1411 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2237 a_6243_9615# XThC.XTBN.Y.t95 XThC.Tn[6].t5 VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2238 VGND.t902 Vbias.t205 XA.XIR[3].XIC[2].icell.SM VGND.t901 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2239 VGND.t904 Vbias.t206 XA.XIR[11].XIC[11].icell.SM VGND.t903 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2240 XA.XIR[10].XIC[12].icell.Ien XThR.Tn[10].t58 VPWR.t709 VPWR.t708 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2241 XThR.Tn[2].t5 XThR.XTBN.Y.t96 a_n1049_7493# VPWR.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2242 VGND.t2595 VPWR.t2037 XA.XIR[7].XIC_15.icell.PDM VGND.t2594 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2243 XA.XIR[10].XIC[7].icell.SM XA.XIR[10].XIC[7].icell.Ien Iout.t250 VGND.t2505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2244 XA.XIR[13].XIC[13].icell.Ien XThR.Tn[13].t57 VPWR.t1791 VPWR.t1790 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2245 XA.XIR[13].XIC[8].icell.SM XA.XIR[13].XIC[8].icell.Ien Iout.t168 VGND.t1482 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2246 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[0].t62 VGND.t1499 VGND.t1498 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2247 XThR.Tn[13].t8 XThR.XTBN.Y.t97 VPWR.t297 VPWR.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2248 XA.XIR[5].XIC[9].icell.PUM XThC.Tn[9].t37 XA.XIR[5].XIC[9].icell.Ien VPWR.t1263 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2249 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[6].t61 VGND.t677 VGND.t676 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2250 XA.XIR[0].XIC[8].icell.Ien XThR.Tn[0].t63 VPWR.t962 VPWR.t961 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2251 XA.XIR[3].XIC[0].icell.SM XA.XIR[3].XIC[0].icell.Ien Iout.t66 VGND.t619 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2252 XA.XIR[9].XIC[9].icell.PUM XThC.Tn[9].t38 XA.XIR[9].XIC[9].icell.Ien VPWR.t1264 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2253 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[2].t56 VGND.t1068 VGND.t1067 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2254 XThR.Tn[10].t4 XThR.XTB3.Y VPWR.t643 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2255 XA.XIR[8].XIC[10].icell.PUM XThC.Tn[10].t37 XA.XIR[8].XIC[10].icell.Ien VPWR.t1307 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2256 XThR.Tn[4].t8 XThR.XTBN.Y.t98 VGND.t437 VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2257 VPWR.t1249 XThR.Tn[12].t61 XA.XIR[13].XIC[6].icell.PUM VPWR.t1248 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2258 VGND.t1804 VGND.t1802 XA.XIR[10].XIC_dummy_left.icell.SM VGND.t1803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2259 VGND.t208 XThR.XTB6.Y XThR.Tn[5].t0 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2260 VGND.t955 XThC.Tn[0].t35 XA.XIR[14].XIC[0].icell.PDM VGND.t954 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2261 XA.XIR[1].XIC[3].icell.PUM XThC.Tn[3].t38 XA.XIR[1].XIC[3].icell.Ien VPWR.t130 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2262 VGND.t906 Vbias.t207 XA.XIR[1].XIC[10].icell.SM VGND.t905 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2263 a_4861_9615# XThC.XTBN.Y.t96 XThC.Tn[3].t1 VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2264 XA.XIR[15].XIC[4].icell.PDM XThR.Tn[14].t63 VGND.t339 VGND.t338 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2265 XA.XIR[0].XIC[11].icell.SM XA.XIR[0].XIC[11].icell.Ien Iout.t49 VGND.t371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2266 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[13].t58 VGND.t2418 VGND.t2417 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2267 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2038 VGND.t2597 VGND.t2596 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2268 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t0 VGND.t1393 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2269 VGND.t230 XThC.Tn[3].t39 XA.XIR[5].XIC[3].icell.PDM VGND.t229 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2270 VGND.t908 Vbias.t208 XA.XIR[11].XIC[9].icell.SM VGND.t907 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2271 XA.XIR[10].XIC[10].icell.Ien XThR.Tn[10].t59 VPWR.t711 VPWR.t710 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2272 XA.XIR[12].XIC_15.icell.SM XA.XIR[12].XIC_15.icell.Ien Iout.t159 VGND.t1290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2273 VGND.t232 XThC.Tn[3].t40 XA.XIR[9].XIC[3].icell.PDM VGND.t231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2274 VGND.t1310 Vbias.t209 XA.XIR[8].XIC[11].icell.SM VGND.t1309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2275 XA.XIR[7].XIC[12].icell.Ien XThR.Tn[7].t55 VPWR.t3 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2276 VPWR.t1725 XThR.Tn[0].t64 XA.XIR[1].XIC[9].icell.PUM VPWR.t1724 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2277 VGND.t2599 VPWR.t2039 XA.XIR[4].XIC_15.icell.PDM VGND.t2598 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2278 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1407 VPWR.t1409 VPWR.t1408 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2279 VGND.t1312 Vbias.t210 XA.XIR[1].XIC[1].icell.SM VGND.t1311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2280 VPWR.t1128 XThR.Tn[4].t63 XA.XIR[5].XIC[9].icell.PUM VPWR.t1127 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2281 VGND.t2683 XThC.Tn[1].t38 XA.XIR[0].XIC[1].icell.PDM VGND.t2682 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2282 XA.XIR[11].XIC[6].icell.PUM XThC.Tn[6].t37 XA.XIR[11].XIC[6].icell.Ien VPWR.t353 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2283 XA.XIR[15].XIC[14].icell.PUM XThC.Tn[14].t38 XA.XIR[15].XIC[14].icell.Ien VPWR.t1109 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2284 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[2].t57 VGND.t1066 VGND.t1065 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2285 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14].t64 XA.XIR[14].XIC[13].icell.Ien VGND.t340 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2286 VGND.t2601 VPWR.t2040 XA.XIR[12].XIC_dummy_right.icell.PDM VGND.t2600 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2287 XA.XIR[10].XIC[2].icell.SM XA.XIR[10].XIC[2].icell.Ien Iout.t77 VGND.t723 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2288 VGND.t2126 XThC.Tn[9].t39 XA.XIR[11].XIC[9].icell.PDM VGND.t2125 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2289 VPWR.t641 XThR.XTB3.Y a_n1049_7493# VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2290 XA.XIR[13].XIC[3].icell.SM XA.XIR[13].XIC[3].icell.Ien Iout.t110 VGND.t1097 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2291 VPWR.t362 XThR.Tn[9].t60 XA.XIR[10].XIC[6].icell.PUM VPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2292 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6].t62 XA.XIR[6].XIC_15.icell.Ien VGND.t678 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2293 VPWR.t1779 XThR.Tn[11].t64 XA.XIR[12].XIC[8].icell.PUM VPWR.t1778 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2294 XA.XIR[0].XIC[3].icell.Ien XThR.Tn[0].t65 VPWR.t1727 VPWR.t1726 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2295 XA.XIR[8].XIC[5].icell.PUM XThC.Tn[5].t35 XA.XIR[8].XIC[5].icell.Ien VPWR.t866 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2296 XA.XIR[13].XIC[6].icell.Ien XThR.Tn[13].t59 VPWR.t1793 VPWR.t1792 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2297 XA.XIR[0].XIC[9].icell.SM XA.XIR[0].XIC[9].icell.Ien Iout.t209 VGND.t2085 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2298 VGND.t1314 Vbias.t211 XA.XIR[5].XIC[8].icell.SM VGND.t1313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2299 VGND.t688 XThC.Tn[7].t32 XA.XIR[5].XIC[7].icell.PDM VGND.t687 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2300 VPWR.t1251 XThR.Tn[12].t62 XA.XIR[13].XIC[1].icell.PUM VPWR.t1250 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2301 XThC.XTB2.Y XThC.XTB6.A a_3523_10575# VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2302 VPWR.t1406 VPWR.t1404 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1405 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2303 VGND.t690 XThC.Tn[7].t33 XA.XIR[9].XIC[7].icell.PDM VGND.t689 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2304 VGND.t1316 Vbias.t212 XA.XIR[8].XIC[9].icell.SM VGND.t1315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2305 XA.XIR[7].XIC[10].icell.Ien XThR.Tn[7].t56 VPWR.t5 VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2306 XThR.Tn[4].t1 XThR.XTB5.Y VGND.t1163 VGND.t209 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2307 VPWR.t298 XThR.XTBN.Y.t99 XThR.Tn[14].t8 VPWR.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2308 VPWR.t713 XThR.Tn[10].t60 XA.XIR[11].XIC[14].icell.PUM VPWR.t712 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2309 XThC.Tn[13].t5 XThC.XTB6.Y VPWR.t760 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2310 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13].t60 XA.XIR[13].XIC[9].icell.Ien VGND.t1597 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2311 VGND.t1174 XThC.XTB6.Y XThC.Tn[5].t0 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2312 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[13].t61 VGND.t1599 VGND.t1598 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2313 XA.XIR[5].XIC[6].icell.SM XA.XIR[5].XIC[6].icell.Ien Iout.t253 VGND.t2649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2314 VPWR.t300 XThR.XTBN.Y.t100 XThR.Tn[11].t8 VPWR.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2315 VGND.t1318 Vbias.t213 XA.XIR[11].XIC[4].icell.SM VGND.t1317 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2316 XA.XIR[10].XIC[5].icell.Ien XThR.Tn[10].t61 VPWR.t715 VPWR.t714 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2317 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[12].t63 VGND.t2117 VGND.t2116 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2318 VGND.t1801 VGND.t1799 XA.XIR[6].XIC_dummy_right.icell.SM VGND.t1800 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2319 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[11].t65 VGND.t2412 VGND.t2411 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2320 XA.XIR[15].XIC[11].icell.SM XA.XIR[15].XIC[11].icell.Ien Iout.t53 VGND.t414 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2321 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[2].t58 XA.XIR[2].XIC[11].icell.Ien VGND.t1064 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2322 XA.XIR[3].XIC[4].icell.PUM XThC.Tn[4].t38 XA.XIR[3].XIC[4].icell.Ien VPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2323 XThC.Tn[9].t0 XThC.XTB2.Y a_7875_9569# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2324 XA.XIR[4].XIC_15.icell.PDM VPWR.t2041 VGND.t2603 VGND.t2602 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2325 XA.XIR[11].XIC[1].icell.PUM XThC.Tn[1].t39 XA.XIR[11].XIC[1].icell.Ien VPWR.t1922 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2326 VGND.t115 XThC.XTB6.A XThC.XTB6.Y VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2327 VGND.t65 XThC.XTB2.Y XThC.Tn[1].t1 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 XA.XIR[10].XIC[13].icell.PUM XThC.Tn[13].t38 XA.XIR[10].XIC[13].icell.Ien VPWR.t1770 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2329 XA.XIR[2].XIC[6].icell.SM XA.XIR[2].XIC[6].icell.Ien Iout.t140 VGND.t1199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2330 VGND.t1320 Vbias.t214 XA.XIR[12].XIC[12].icell.SM VGND.t1319 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2331 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1402 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1403 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2332 XThC.Tn[6].t4 XThC.XTBN.Y.t97 a_6243_9615# VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2333 XA.XIR[6].XIC[14].icell.SM XA.XIR[6].XIC[14].icell.Ien Iout.t245 VGND.t2486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2334 VGND.t1322 Vbias.t215 XA.XIR[15].XIC[13].icell.SM VGND.t1321 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2335 VGND.t1324 Vbias.t216 XA.XIR[14].XIC[14].icell.SM VGND.t1323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2336 VGND.t2551 XThC.Tn[12].t37 XA.XIR[15].XIC[12].icell.PDM VGND.t2550 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2337 VGND.t85 XThC.Tn[4].t39 XA.XIR[11].XIC[4].icell.PDM VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2338 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[2].t59 XA.XIR[2].XIC[2].icell.Ien VGND.t1063 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2339 VPWR.t990 XThR.XTB7.Y a_n1049_5317# VPWR.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2340 VPWR.t364 XThR.Tn[9].t61 XA.XIR[10].XIC[1].icell.PUM VPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2341 VGND.t2605 VPWR.t2042 XA.XIR[6].XIC_dummy_right.icell.PDM VGND.t2604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2342 VPWR.t759 XThC.XTB6.Y XThC.Tn[13].t4 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2343 VPWR.t1781 XThR.Tn[11].t66 XA.XIR[12].XIC[3].icell.PUM VPWR.t1780 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2344 a_n997_3979# XThR.XTBN.Y.t101 VGND.t438 VGND.t378 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2345 XA.XIR[5].XIC[4].icell.Ien XThR.Tn[5].t60 VPWR.t1751 VPWR.t1750 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2346 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13].t62 VPWR.t1025 VPWR.t1024 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2347 XA.XIR[9].XIC[4].icell.Ien XThR.Tn[9].t62 VPWR.t366 VPWR.t365 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2348 XA.XIR[0].XIC[4].icell.SM XA.XIR[0].XIC[4].icell.Ien Iout.t184 VGND.t1568 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2349 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1399 VPWR.t1401 VPWR.t1400 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2350 VGND.t1326 Vbias.t217 XA.XIR[5].XIC[3].icell.SM VGND.t1325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2351 VGND.t1328 Vbias.t218 XA.XIR[9].XIC[12].icell.SM VGND.t1327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2352 XA.XIR[9].XIC[7].icell.SM XA.XIR[9].XIC[7].icell.Ien Iout.t117 VGND.t1123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2353 VGND.t650 XThR.XTB4.Y XThR.Tn[3].t0 VGND.t649 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2354 XA.XIR[5].XIC[10].icell.SM XA.XIR[5].XIC[10].icell.Ien Iout.t169 VGND.t1483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2355 a_7331_10587# data[0].t2 VPWR.t748 VPWR.t747 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2356 a_4067_9615# XThC.XTBN.Y.t98 XThC.Tn[2].t2 VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2357 VPWR.t786 XThR.Tn[2].t60 XA.XIR[3].XIC[12].icell.PUM VPWR.t785 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2358 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[12].t64 VGND.t2119 VGND.t2118 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2359 XA.XIR[12].XIC[8].icell.SM XA.XIR[12].XIC[8].icell.Ien Iout.t237 VGND.t2478 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2360 XA.XIR[11].XIC[14].icell.Ien XThR.Tn[11].t67 VPWR.t1783 VPWR.t1782 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2361 VGND.t1330 Vbias.t219 XA.XIR[8].XIC[4].icell.SM VGND.t1329 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2362 VGND.t1798 VGND.t1796 XA.XIR[3].XIC_dummy_right.icell.SM VGND.t1797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2363 XA.XIR[7].XIC[5].icell.Ien XThR.Tn[7].t57 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2364 VPWR.t488 XThR.Tn[6].t63 XA.XIR[7].XIC[12].icell.PUM VPWR.t487 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2365 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13].t63 XA.XIR[13].XIC[4].icell.Ien VGND.t1600 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2366 XA.XIR[15].XIC[9].icell.SM XA.XIR[15].XIC[9].icell.Ien Iout.t75 VGND.t719 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2367 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t2043 XA.XIR[8].XIC_dummy_right.icell.Ien VGND.t2606 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2368 VPWR.t1753 XThR.Tn[5].t61 XA.XIR[6].XIC[13].icell.PUM VPWR.t1752 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2369 a_n1049_6699# XThR.XTBN.Y.t102 XThR.Tn[3].t4 VPWR.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2370 XA.XIR[0].XIC[11].icell.PDM VGND.t1793 VGND.t1795 VGND.t1794 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2371 XA.XIR[3].XIC[0].icell.PUM XThC.Tn[0].t36 XA.XIR[3].XIC[0].icell.Ien VPWR.t1880 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2372 XA.XIR[1].XIC_15.icell.PDM VPWR.t2044 VGND.t2608 VGND.t2607 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2373 XA.XIR[5].XIC[1].icell.SM XA.XIR[5].XIC[1].icell.Ien Iout.t251 VGND.t2506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2374 XA.XIR[2].XIC[10].icell.SM XA.XIR[2].XIC[10].icell.Ien Iout.t226 VGND.t2268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2375 XThC.Tn[3].t0 XThC.XTBN.Y.t99 a_4861_9615# VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2376 XA.XIR[3].XIC[14].icell.SM XA.XIR[3].XIC[14].icell.Ien Iout.t2 VGND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2377 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1397 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1398 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2378 XThC.XTB5.A data[0].t3 VGND.t1161 VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2379 VGND.t2196 XThC.Tn[10].t38 XA.XIR[15].XIC[10].icell.PDM VGND.t2195 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2380 VPWR.t464 XThR.XTB4.Y XThR.Tn[11].t5 VPWR.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2381 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[2].t61 XA.XIR[2].XIC[6].icell.Ien VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2382 XA.XIR[0].XIC[2].icell.PDM VGND.t1790 VGND.t1792 VGND.t1791 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2383 XA.XIR[2].XIC[1].icell.SM XA.XIR[2].XIC[1].icell.Ien Iout.t144 VGND.t1211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2384 VGND.t432 XThC.Tn[11].t36 XA.XIR[2].XIC[11].icell.PDM VGND.t431 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2385 VGND.t440 XThR.XTBN.Y.t103 a_n997_715# VGND.t439 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2386 a_n997_2891# XThR.XTBN.Y.t104 VGND.t441 VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2387 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[7].t58 VGND.t4 VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2388 VGND.t1789 VGND.t1787 XA.XIR[6].XIC_dummy_left.icell.SM VGND.t1788 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2389 XA.XIR[5].XIC[0].icell.Ien XThR.Tn[5].t62 VPWR.t1755 VPWR.t1754 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2390 VPWR.t370 XThR.Tn[3].t66 XA.XIR[4].XIC[9].icell.PUM VPWR.t369 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2391 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9].t63 VPWR.t368 VPWR.t367 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2392 VPWR.t784 XThR.Tn[2].t62 XA.XIR[3].XIC[10].icell.PUM VPWR.t783 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2393 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1394 VPWR.t1396 VPWR.t1395 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2394 VPWR.t490 XThR.Tn[6].t64 XA.XIR[7].XIC[10].icell.PUM VPWR.t489 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2395 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14].t65 XA.XIR[14].XIC[1].icell.Ien VGND.t341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2396 XA.XIR[10].XIC[6].icell.PUM XThC.Tn[6].t38 XA.XIR[10].XIC[6].icell.Ien VPWR.t354 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2397 XThR.Tn[11].t0 XThR.XTB4.Y a_n997_2667# VGND.t648 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2398 VPWR.t1393 VPWR.t1391 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1392 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2399 VGND.t2150 XThC.Tn[2].t36 XA.XIR[2].XIC[2].icell.PDM VGND.t2149 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2400 XA.XIR[13].XIC[7].icell.PUM XThC.Tn[7].t34 XA.XIR[13].XIC[7].icell.Ien VPWR.t504 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2401 XA.XIR[9].XIC[2].icell.SM XA.XIR[9].XIC[2].icell.Ien Iout.t187 VGND.t1596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2402 VPWR.t50 XThC.XTB2.Y XThC.Tn[9].t4 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2403 XA.XIR[3].XIC[12].icell.Ien XThR.Tn[3].t67 VPWR.t372 VPWR.t371 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2404 a_n997_3979# XThR.XTB1.Y XThR.Tn[8].t1 VGND.t1396 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2405 VGND.t2610 VPWR.t2045 XA.XIR[0].XIC_15.icell.PDM VGND.t2609 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2406 VGND.t2128 XThC.Tn[9].t40 XA.XIR[10].XIC[9].icell.PDM VGND.t2127 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2407 XA.XIR[12].XIC[3].icell.SM XA.XIR[12].XIC[3].icell.Ien Iout.t154 VGND.t1274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2408 VPWR.t444 XThC.XTBN.Y.t100 XThC.Tn[8].t8 VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2409 XA.XIR[15].XIC[4].icell.SM XA.XIR[15].XIC[4].icell.Ien Iout.t15 VGND.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2410 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[4].t64 XA.XIR[4].XIC[8].icell.Ien VGND.t241 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2411 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[4].t65 XA.XIR[4].XIC[14].icell.Ien VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2412 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout VGND.t2371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2413 a_n1335_8331# XThR.XTB5.A XThR.XTB1.Y VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2414 VPWR.t180 XThR.Tn[14].t66 XA.XIR[15].XIC[8].icell.PUM VPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2415 XA.XIR[0].XIC[6].icell.PDM VGND.t1784 VGND.t1786 VGND.t1785 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2416 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11].t68 XA.XIR[11].XIC[12].icell.Ien VGND.t2413 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2417 a_n1049_6405# XThR.XTBN.Y.t105 XThR.Tn[4].t4 VPWR.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2418 XA.XIR[15].XIC[7].icell.Ien VPWR.t1388 VPWR.t1390 VPWR.t1389 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2419 XThR.Tn[7].t4 XThR.XTBN.Y.t106 VPWR.t303 VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2420 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2046 VGND.t2612 VGND.t2611 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2421 VPWR.t1757 XThR.Tn[5].t63 XA.XIR[6].XIC[6].icell.PUM VPWR.t1756 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2422 VGND.t1783 VGND.t1781 XA.XIR[3].XIC_dummy_left.icell.SM VGND.t1782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2423 VPWR.t1219 XThR.Tn[8].t64 XA.XIR[9].XIC[7].icell.PUM VPWR.t1218 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2424 XThC.Tn[9].t8 XThC.XTBN.Y.t101 VPWR.t445 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2425 XThR.Tn[1].t9 XThR.XTBN.Y.t107 VGND.t443 VGND.t442 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2426 VPWR.t1374 VPWR.t1372 XA.XIR[13].XIC_15.icell.PUM VPWR.t1373 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2427 VGND.t1332 Vbias.t220 XA.XIR[2].XIC[7].icell.SM VGND.t1331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2428 VGND.t479 XThC.Tn[6].t39 XA.XIR[2].XIC[6].icell.PDM VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2429 XA.XIR[13].XIC[11].icell.PUM XThC.Tn[11].t37 XA.XIR[13].XIC[11].icell.Ien VPWR.t295 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2430 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[11].t69 VGND.t2415 VGND.t2414 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2431 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[7].t59 VGND.t793 VGND.t792 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2432 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2047 VGND.t2614 VGND.t2613 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2433 XA.XIR[4].XIC[9].icell.Ien XThR.Tn[4].t66 VPWR.t138 VPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2434 XA.XIR[3].XIC[10].icell.Ien XThR.Tn[3].t68 VPWR.t374 VPWR.t373 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2435 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[10].t62 VGND.t1099 VGND.t1098 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2436 XA.XIR[14].XIC[11].icell.SM XA.XIR[14].XIC[11].icell.Ien Iout.t84 VGND.t770 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2437 XA.XIR[15].XIC[13].icell.PDM XThR.Tn[14].t67 VGND.t322 VGND.t321 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2438 VPWR.t446 XThC.XTBN.Y.t102 XThC.Tn[11].t3 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2439 VPWR.t782 XThR.Tn[2].t63 XA.XIR[3].XIC[5].icell.PUM VPWR.t781 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2440 VPWR.t119 XThR.XTB6.Y a_n1049_5611# VPWR.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2441 VGND.t2616 VPWR.t2048 XA.XIR[15].XIC_dummy_left.icell.PDM VGND.t2615 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2442 a_n997_2891# XThR.XTB3.Y XThR.Tn[10].t1 VGND.t657 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2443 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[1].t59 XA.XIR[1].XIC[11].icell.Ien VGND.t254 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2444 XA.XIR[13].XIC[12].icell.SM XA.XIR[13].XIC[12].icell.Ien Iout.t80 VGND.t748 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2445 VPWR.t492 XThR.Tn[6].t65 XA.XIR[7].XIC[5].icell.PUM VPWR.t491 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2446 XA.XIR[10].XIC[1].icell.PUM XThC.Tn[1].t40 XA.XIR[10].XIC[1].icell.Ien VPWR.t1923 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2447 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1386 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1387 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2448 XA.XIR[1].XIC[6].icell.SM XA.XIR[1].XIC[6].icell.Ien Iout.t131 VGND.t1173 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2449 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[1].t60 VGND.t2104 VGND.t2103 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2450 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[1].t61 VGND.t2106 VGND.t2105 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2451 XA.XIR[13].XIC[2].icell.PUM XThC.Tn[2].t37 XA.XIR[13].XIC[2].icell.Ien VPWR.t1275 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2452 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11].t70 XA.XIR[11].XIC[10].icell.Ien VGND.t2416 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2453 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[8].t65 VGND.t2095 VGND.t2094 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2454 XA.XIR[8].XIC[14].icell.PUM XThC.Tn[14].t39 XA.XIR[8].XIC[14].icell.Ien VPWR.t1110 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2455 VGND.t1714 Vbias.t221 XA.XIR[10].XIC[5].icell.SM VGND.t1713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2456 XA.XIR[15].XIC[11].icell.Ien VPWR.t1383 VPWR.t1385 VPWR.t1384 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2457 VGND.t87 XThC.Tn[4].t40 XA.XIR[10].XIC[4].icell.PDM VGND.t86 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2458 VGND.t2618 VPWR.t2049 XA.XIR[5].XIC_dummy_right.icell.PDM VGND.t2617 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2459 XA.XIR[11].XIC_15.icell.PUM VPWR.t1381 XA.XIR[11].XIC_15.icell.Ien VPWR.t1382 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2460 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[1].t62 XA.XIR[1].XIC[2].icell.Ien VGND.t2107 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2461 VGND.t1716 Vbias.t222 XA.XIR[13].XIC[6].icell.SM VGND.t1715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2462 XA.XIR[12].XIC[7].icell.Ien XThR.Tn[12].t65 VPWR.t1253 VPWR.t1252 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2463 VGND.t1240 XThC.Tn[5].t36 XA.XIR[13].XIC[5].icell.PDM VGND.t1239 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2464 VGND.t2620 VPWR.t2050 XA.XIR[9].XIC_dummy_right.icell.PDM VGND.t2619 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2465 XThC.Tn[2].t1 XThC.XTBN.Y.t103 a_4067_9615# VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2466 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[4].t67 XA.XIR[4].XIC[3].icell.Ien VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2467 VPWR.t1221 XThR.Tn[8].t66 XA.XIR[9].XIC[11].icell.PUM VPWR.t1220 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2468 VPWR.t182 XThR.Tn[14].t68 XA.XIR[15].XIC[3].icell.PUM VPWR.t181 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2469 XA.XIR[7].XIC[12].icell.PUM XThC.Tn[12].t38 XA.XIR[7].XIC[12].icell.Ien VPWR.t995 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2470 VGND.t1919 XThR.XTB7.B XThR.XTB4.Y VGND.t1918 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2471 VPWR.t1380 VPWR.t1378 XA.XIR[10].XIC_15.icell.PUM VPWR.t1379 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2472 VGND.t1718 Vbias.t223 XA.XIR[4].XIC_15.icell.SM VGND.t1717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2473 XA.XIR[15].XIC[2].icell.Ien VPWR.t1375 VPWR.t1377 VPWR.t1376 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2474 VGND.t1720 Vbias.t224 XA.XIR[11].XIC[13].icell.SM VGND.t1719 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2475 XA.XIR[10].XIC[14].icell.Ien XThR.Tn[10].t63 VPWR.t717 VPWR.t716 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2476 VGND.t1910 XThR.XTB1.Y XThR.Tn[0].t0 VGND.t1397 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2477 VPWR.t1229 XThR.Tn[1].t63 XA.XIR[2].XIC[4].icell.PUM VPWR.t1228 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2478 VPWR.t1759 XThR.Tn[5].t64 XA.XIR[6].XIC[1].icell.PUM VPWR.t1758 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2479 XA.XIR[13].XIC_15.icell.Ien XThR.Tn[13].t64 VPWR.t1027 VPWR.t1026 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2480 XA.XIR[14].XIC[9].icell.SM XA.XIR[14].XIC[9].icell.Ien Iout.t240 VGND.t2481 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2481 VPWR.t1223 XThR.Tn[8].t67 XA.XIR[9].XIC[2].icell.PUM VPWR.t1222 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2482 XA.XIR[15].XIC[5].icell.PDM VPWR.t2051 XA.XIR[15].XIC[5].icell.Ien VGND.t2621 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2483 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout VGND.t1484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2484 VGND.t434 XThC.Tn[11].t38 XA.XIR[14].XIC[11].icell.PDM VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2485 VGND.t1722 Vbias.t225 XA.XIR[2].XIC[2].icell.SM VGND.t1721 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2486 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1369 VPWR.t1371 VPWR.t1370 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2487 XA.XIR[1].XIC[10].icell.SM XA.XIR[1].XIC[10].icell.Ien Iout.t54 VGND.t467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2488 a_8739_9569# XThC.XTBN.Y.t104 VGND.t595 VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2489 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[8].t68 VGND.t2097 VGND.t2096 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2490 XThC.Tn[6].t0 XThC.XTB7.Y VGND.t1299 VGND.t1298 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2491 XA.XIR[3].XIC[5].icell.Ien XThR.Tn[3].t69 VPWR.t376 VPWR.t375 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2492 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[10].t64 VGND.t1101 VGND.t1100 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2493 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[5].t65 VGND.t2251 VGND.t2250 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2494 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[1].t64 XA.XIR[1].XIC[6].icell.Ien VGND.t2108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2495 VGND.t1724 Vbias.t226 XA.XIR[13].XIC[10].icell.SM VGND.t1723 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2496 VGND.t597 XThC.XTBN.Y.t105 XThC.Tn[7].t0 VGND.t596 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2497 XThC.Tn[12].t8 XThC.XTBN.Y.t106 VPWR.t447 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2498 XA.XIR[12].XIC[11].icell.Ien XThR.Tn[12].t66 VPWR.t943 VPWR.t942 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2499 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[4].t68 XA.XIR[4].XIC[7].icell.Ien VGND.t244 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2500 VGND.t2152 XThC.Tn[2].t38 XA.XIR[14].XIC[2].icell.PDM VGND.t2151 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2501 XThC.Tn[12].t0 XThC.XTB5.Y a_9827_9569# VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2502 XA.XIR[1].XIC[1].icell.SM XA.XIR[1].XIC[1].icell.Ien Iout.t30 VGND.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2503 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[1].t65 VGND.t2110 VGND.t2109 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2504 XA.XIR[7].XIC[10].icell.PUM XThC.Tn[10].t39 XA.XIR[7].XIC[10].icell.Ien VPWR.t1308 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2505 XA.XIR[4].XIC[12].icell.PUM XThC.Tn[12].t39 XA.XIR[4].XIC[12].icell.Ien VPWR.t996 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2506 a_8963_9569# XThC.XTB4.Y.t15 XThC.Tn[11].t9 VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2507 XA.XIR[0].XIC[13].icell.SM XA.XIR[0].XIC[13].icell.Ien Iout.t91 VGND.t876 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2508 XA.XIR[3].XIC[13].icell.PUM XThC.Tn[13].t39 XA.XIR[3].XIC[13].icell.Ien VPWR.t1771 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2509 VGND.t1726 Vbias.t227 XA.XIR[10].XIC[0].icell.SM VGND.t1725 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2510 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1367 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1368 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2511 VGND.t1728 Vbias.t228 XA.XIR[5].XIC[12].icell.SM VGND.t1727 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2512 VGND.t316 XThC.Tn[8].t40 XA.XIR[1].XIC[8].icell.PDM VGND.t315 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2513 VGND.t1946 XThC.Tn[14].t40 XA.XIR[1].XIC[14].icell.PDM VGND.t1945 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2514 XThR.Tn[13].t5 XThR.XTB6.Y VPWR.t117 VPWR.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2515 VGND.t1730 Vbias.t229 XA.XIR[13].XIC[1].icell.SM VGND.t1729 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2516 XA.XIR[12].XIC[2].icell.Ien XThR.Tn[12].t67 VPWR.t945 VPWR.t944 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2517 VGND.t2529 XThC.Tn[0].t37 XA.XIR[13].XIC[0].icell.PDM VGND.t2528 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2518 VGND.t1732 Vbias.t230 XA.XIR[8].XIC[13].icell.SM VGND.t1731 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2519 XA.XIR[7].XIC[14].icell.Ien XThR.Tn[7].t60 VPWR.t594 VPWR.t593 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2520 VGND.t1560 XThC.Tn[12].t40 XA.XIR[8].XIC[12].icell.PDM VGND.t1559 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2521 VPWR.t1231 XThR.Tn[1].t66 XA.XIR[2].XIC[0].icell.PUM VPWR.t1230 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2522 VGND.t2270 XThC.Tn[13].t40 XA.XIR[11].XIC[13].icell.PDM VGND.t2269 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2523 XA.XIR[12].XIC[7].icell.PUM XThC.Tn[7].t35 XA.XIR[12].XIC[7].icell.Ien VPWR.t317 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2524 VGND.t598 XThC.XTBN.Y.t107 a_7875_9569# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2525 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12].t68 XA.XIR[12].XIC[5].icell.Ien VGND.t1410 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2526 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2052 XA.XIR[11].XIC_dummy_left.icell.Ien VGND.t2622 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2527 XA.XIR[15].XIC[8].icell.PUM XThC.Tn[8].t41 XA.XIR[15].XIC[8].icell.Ien VPWR.t177 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2528 XA.XIR[2].XIC[4].icell.Ien XThR.Tn[2].t64 VPWR.t780 VPWR.t779 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2529 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14].t69 XA.XIR[14].XIC_15.icell.Ien VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2530 XA.XIR[11].XIC_15.icell.SM XA.XIR[11].XIC_15.icell.Ien Iout.t127 VGND.t1152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2531 VGND.t1734 Vbias.t231 XA.XIR[7].XIC[11].icell.SM VGND.t1733 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2532 XA.XIR[6].XIC[12].icell.Ien XThR.Tn[6].t66 VPWR.t494 VPWR.t493 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2533 XA.XIR[5].XIC[13].icell.Ien XThR.Tn[5].t66 VPWR.t1761 VPWR.t1760 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2534 XA.XIR[14].XIC[4].icell.SM XA.XIR[14].XIC[4].icell.Ien Iout.t238 VGND.t2479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2535 XA.XIR[9].XIC[13].icell.Ien XThR.Tn[9].t64 VPWR.t382 VPWR.t381 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2536 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[5].t67 VGND.t2253 VGND.t2252 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2537 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout VGND.t1445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2538 VPWR.t1054 VGND.t2700 XA.XIR[0].XIC[12].icell.PUM VPWR.t1053 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2539 XA.XIR[15].XIC[0].icell.PDM VPWR.t2053 XA.XIR[15].XIC[0].icell.Ien VGND.t2623 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2540 a_8963_9569# XThC.XTBN.Y.t108 VGND.t599 VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2541 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10].t65 XA.XIR[10].XIC[12].icell.Ien VGND.t1102 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2542 VGND.t481 XThC.Tn[6].t40 XA.XIR[14].XIC[6].icell.PDM VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2543 XA.XIR[1].XIC[9].icell.PUM XThC.Tn[9].t41 XA.XIR[1].XIC[9].icell.Ien VPWR.t1265 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2544 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[1].t67 VGND.t2092 VGND.t2091 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2545 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13].t65 XA.XIR[13].XIC[13].icell.Ien VGND.t1601 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2546 VPWR.t1366 VPWR.t1364 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1365 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2547 XA.XIR[4].XIC[10].icell.PUM XThC.Tn[10].t40 XA.XIR[4].XIC[10].icell.Ien VPWR.t1309 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2548 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[13].t66 VGND.t2553 VGND.t2552 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2549 XA.XIR[0].XIC[8].icell.PDM XThR.Tn[0].t66 XA.XIR[0].XIC[8].icell.Ien VGND.t2233 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2550 XA.XIR[0].XIC[14].icell.PDM XThR.Tn[0].t67 XA.XIR[0].XIC[14].icell.Ien VGND.t2234 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2551 VPWR.t596 XThR.Tn[7].t61 XA.XIR[8].XIC[7].icell.PUM VPWR.t595 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2552 VGND.t2198 XThC.Tn[10].t41 XA.XIR[8].XIC[10].icell.PDM VGND.t2197 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2553 XThC.Tn[11].t2 XThC.XTBN.Y.t109 VPWR.t1326 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2554 VPWR.t1913 XThR.Tn[10].t66 XA.XIR[11].XIC[8].icell.PUM VPWR.t1912 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2555 VGND.t1736 Vbias.t232 XA.XIR[1].XIC[7].icell.SM VGND.t1735 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2556 XThR.Tn[6].t5 XThR.XTBN.Y.t108 a_n1049_5317# VPWR.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2557 XA.XIR[7].XIC[5].icell.PUM XThC.Tn[5].t37 XA.XIR[7].XIC[5].icell.Ien VPWR.t999 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2558 VPWR.t156 XThC.XTB4.Y.t16 XThC.Tn[11].t0 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2559 XThR.XTB7.Y XThR.XTB7.B a_n1319_5317# VPWR.t1098 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2560 XA.XIR[12].XIC[11].icell.PUM XThC.Tn[11].t39 XA.XIR[12].XIC[11].icell.Ien VPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2561 VGND.t1743 Vbias.t233 XA.XIR[4].XIC[8].icell.SM VGND.t1742 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2562 XA.XIR[15].XIC[1].icell.PDM XThR.Tn[14].t70 VGND.t325 VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2563 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[13].t67 VGND.t2555 VGND.t2554 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2564 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[9].t65 VGND.t539 VGND.t538 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2565 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2054 VGND.t2625 VGND.t2624 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2566 VGND.t234 XThC.Tn[3].t41 XA.XIR[1].XIC[3].icell.PDM VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2567 VGND.t1745 Vbias.t234 XA.XIR[7].XIC[9].icell.SM VGND.t1744 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2568 XA.XIR[6].XIC[10].icell.Ien XThR.Tn[6].t67 VPWR.t496 VPWR.t495 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2569 XA.XIR[2].XIC[0].icell.Ien XThR.Tn[2].t65 VPWR.t778 VPWR.t777 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2570 XA.XIR[12].XIC_15.icell.PDM VPWR.t2055 VGND.t2627 VGND.t2626 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2571 XA.XIR[12].XIC[12].icell.SM XA.XIR[12].XIC[12].icell.Ien Iout.t163 VGND.t1296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2572 XA.XIR[8].XIC_15.icell.SM XA.XIR[8].XIC_15.icell.Ien Iout.t197 VGND.t1937 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2573 XA.XIR[15].XIC[13].icell.SM XA.XIR[15].XIC[13].icell.Ien Iout.t106 VGND.t1073 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2574 VPWR.t1052 VGND.t2701 XA.XIR[0].XIC[10].icell.PUM VPWR.t1051 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2575 VPWR.t631 XThC.XTB3.Y.t14 a_4067_9615# VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2576 XA.XIR[3].XIC[6].icell.PUM XThC.Tn[6].t41 XA.XIR[3].XIC[6].icell.Ien VPWR.t327 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2577 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12].t69 XA.XIR[12].XIC[0].icell.Ien VGND.t1411 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2578 XA.XIR[12].XIC[2].icell.PUM XThC.Tn[2].t39 XA.XIR[12].XIC[2].icell.Ien VPWR.t1276 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2579 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10].t67 XA.XIR[10].XIC[10].icell.Ien VGND.t2669 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2580 VGND.t351 XThR.XTBN.Y.t109 a_n997_1803# VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2581 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7].t62 XA.XIR[7].XIC[12].icell.Ien VGND.t794 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2582 XA.XIR[0].XIC[9].icell.Ien XThR.Tn[0].t68 VPWR.t1729 VPWR.t1728 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2583 XA.XIR[15].XIC[3].icell.PUM XThC.Tn[3].t42 XA.XIR[15].XIC[3].icell.Ien VPWR.t131 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2584 XA.XIR[6].XIC[7].icell.PUM XThC.Tn[7].t36 XA.XIR[6].XIC[7].icell.Ien VPWR.t318 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2585 XA.XIR[10].XIC_15.icell.PUM VPWR.t1362 XA.XIR[10].XIC_15.icell.Ien VPWR.t1363 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2586 a_3773_9615# XThC.XTB2.Y VPWR.t48 VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2587 VPWR.t1361 VPWR.t1359 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1360 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2588 VGND.t1747 Vbias.t235 XA.XIR[12].XIC[6].icell.SM VGND.t1746 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2589 VGND.t2130 XThC.Tn[9].t42 XA.XIR[3].XIC[9].icell.PDM VGND.t2129 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2590 VGND.t1570 XThC.Tn[5].t38 XA.XIR[12].XIC[5].icell.PDM VGND.t1569 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2591 VPWR.t598 XThR.Tn[7].t63 XA.XIR[8].XIC[11].icell.PUM VPWR.t597 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2592 XA.XIR[2].XIC[4].icell.PUM XThC.Tn[4].t41 XA.XIR[2].XIC[4].icell.Ien VPWR.t78 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2593 VPWR.t462 XThR.XTB4.Y XThR.Tn[11].t4 VPWR.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2594 a_n997_715# XThR.XTBN.Y.t110 VGND.t353 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2595 VGND.t1749 Vbias.t236 XA.XIR[6].XIC[5].icell.SM VGND.t1748 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2596 VPWR.t1081 XThR.XTB1.Y a_n1049_8581# VPWR.t1080 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2597 XA.XIR[4].XIC[5].icell.PUM XThC.Tn[5].t39 XA.XIR[4].XIC[5].icell.Ien VPWR.t1000 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2598 XA.XIR[5].XIC[6].icell.Ien XThR.Tn[5].t68 VPWR.t1763 VPWR.t1762 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2599 XThR.Tn[14].t5 XThR.XTB7.Y VPWR.t989 VPWR.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2600 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[13].t68 VGND.t2557 VGND.t2556 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2601 XA.XIR[9].XIC[6].icell.Ien XThR.Tn[9].t66 VPWR.t384 VPWR.t383 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2602 VGND.t1751 Vbias.t237 XA.XIR[9].XIC[6].icell.SM VGND.t1750 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2603 VGND.t2213 XThC.XTBN.Y.t110 XThC.Tn[3].t5 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2604 XA.XIR[8].XIC[7].icell.Ien XThR.Tn[8].t69 VPWR.t1225 VPWR.t1224 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2605 VGND.t469 XThC.Tn[7].t37 XA.XIR[1].XIC[7].icell.PDM VGND.t468 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2606 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2056 VGND.t2629 VGND.t2628 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2607 XA.XIR[0].XIC[3].icell.PDM XThR.Tn[0].t69 XA.XIR[0].XIC[3].icell.Ien VGND.t2235 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2608 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout VGND.t177 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2609 VPWR.t600 XThR.Tn[7].t64 XA.XIR[8].XIC[2].icell.PUM VPWR.t599 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2610 XThC.Tn[1].t0 XThC.XTB2.Y VGND.t64 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2611 VPWR.t776 XThR.Tn[2].t66 XA.XIR[3].XIC[14].icell.PUM VPWR.t775 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2612 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5].t69 XA.XIR[5].XIC[9].icell.Ien VGND.t1055 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2613 XA.XIR[11].XIC[8].icell.Ien XThR.Tn[11].t71 VPWR.t91 VPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2614 VPWR.t1199 XThC.XTBN.A XThC.XTBN.Y.t2 VPWR.t1198 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2615 VPWR.t1915 XThR.Tn[10].t68 XA.XIR[11].XIC[3].icell.PUM VPWR.t1914 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2616 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9].t67 XA.XIR[9].XIC[9].icell.Ien VGND.t540 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2617 VPWR.t498 XThR.Tn[6].t68 XA.XIR[7].XIC[14].icell.PUM VPWR.t497 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2618 VGND.t1753 Vbias.t238 XA.XIR[1].XIC[2].icell.SM VGND.t1752 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2619 VPWR.t1358 VPWR.t1356 XA.XIR[6].XIC_15.icell.PUM VPWR.t1357 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2620 VGND.t1755 Vbias.t239 XA.XIR[4].XIC[3].icell.SM VGND.t1754 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2621 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7].t65 XA.XIR[7].XIC[10].icell.Ien VGND.t795 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2622 XThR.Tn[2].t7 XThR.XTB3.Y VGND.t867 VGND.t655 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2623 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[9].t68 VGND.t542 VGND.t541 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2624 XA.XIR[6].XIC[11].icell.PUM XThC.Tn[11].t40 XA.XIR[6].XIC[11].icell.Ien VPWR.t281 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2625 XA.XIR[11].XIC[8].icell.SM XA.XIR[11].XIC[8].icell.Ien Iout.t74 VGND.t691 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2626 VGND.t1757 Vbias.t240 XA.XIR[7].XIC[4].icell.SM VGND.t1756 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2627 XA.XIR[6].XIC[5].icell.Ien XThR.Tn[6].t69 VPWR.t500 VPWR.t499 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2628 VGND.t1780 VGND.t1778 XA.XIR[2].XIC_dummy_right.icell.SM VGND.t1779 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2629 VGND.t1759 Vbias.t241 XA.XIR[12].XIC[10].icell.SM VGND.t1758 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2630 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[7].t66 VGND.t797 VGND.t796 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2631 a_n997_3979# XThR.XTB1.Y XThR.Tn[8].t0 VGND.t1393 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2632 XA.XIR[7].XIC[11].icell.SM XA.XIR[7].XIC[11].icell.Ien Iout.t218 VGND.t2168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2633 a_3299_10575# XThC.XTB7.B VGND.t1132 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2634 VGND.t2631 VPWR.t2057 XA.XIR[8].XIC_dummy_left.icell.PDM VGND.t2630 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2635 VGND.t355 XThR.XTBN.Y.t111 XThR.Tn[6].t8 VGND.t354 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2636 VPWR.t1050 VGND.t2702 XA.XIR[0].XIC[5].icell.PUM VPWR.t1049 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2637 XA.XIR[3].XIC[1].icell.PUM XThC.Tn[1].t41 XA.XIR[3].XIC[1].icell.Ien VPWR.t1924 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2638 XA.XIR[2].XIC[0].icell.PUM XThC.Tn[0].t38 XA.XIR[2].XIC[0].icell.Ien VPWR.t1881 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2639 VPWR.t93 XThR.Tn[11].t72 XA.XIR[12].XIC[9].icell.PUM VPWR.t92 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2640 XA.XIR[6].XIC[2].icell.PUM XThC.Tn[2].t40 XA.XIR[6].XIC[2].icell.Ien VPWR.t1277 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2641 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1353 VPWR.t1355 VPWR.t1354 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2642 VGND.t1761 Vbias.t242 XA.XIR[12].XIC[1].icell.SM VGND.t1760 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2643 VGND.t1763 Vbias.t243 XA.XIR[3].XIC[5].icell.SM VGND.t1762 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2644 VGND.t2531 XThC.Tn[0].t39 XA.XIR[12].XIC[0].icell.PDM VGND.t2530 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2645 VGND.t89 XThC.Tn[4].t42 XA.XIR[3].XIC[4].icell.PDM VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2646 VGND.t1765 Vbias.t244 XA.XIR[9].XIC[10].icell.SM VGND.t1764 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2647 XA.XIR[8].XIC[11].icell.Ien XThR.Tn[8].t70 VPWR.t1227 VPWR.t1226 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2648 VGND.t1419 XThC.Tn[1].t42 XA.XIR[11].XIC[1].icell.PDM VGND.t1418 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2649 VGND.t1524 Vbias.t245 XA.XIR[10].XIC[14].icell.SM VGND.t1523 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2650 XA.XIR[0].XIC[7].icell.PDM XThR.Tn[0].t70 XA.XIR[0].XIC[7].icell.Ien VGND.t2236 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2651 VGND.t1572 XThC.Tn[5].t40 XA.XIR[6].XIC[5].icell.PDM VGND.t1571 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2652 VPWR.t1327 XThC.XTBN.Y.t111 XThC.Tn[10].t7 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2653 VGND.t2272 XThC.Tn[13].t41 XA.XIR[10].XIC[13].icell.PDM VGND.t2271 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2654 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2058 XA.XIR[10].XIC_dummy_left.icell.Ien VGND.t2632 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2655 XA.XIR[0].XIC[12].icell.PUM XThC.Tn[12].t41 XA.XIR[0].XIC[12].icell.Ien VPWR.t997 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2656 VGND.t2214 XThC.XTBN.Y.t112 a_8963_9569# VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2657 XA.XIR[5].XIC[1].icell.Ien XThR.Tn[5].t70 VPWR.t696 VPWR.t695 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2658 VGND.t1526 Vbias.t246 XA.XIR[6].XIC[0].icell.SM VGND.t1525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2659 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[6].t70 VGND.t591 VGND.t590 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2660 VPWR.t550 XThC.XTB5.A a_5155_10571# VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2661 VPWR.t911 XThC.XTB7.Y XThC.Tn[14].t4 VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2662 XThR.Tn[1].t8 XThR.XTBN.Y.t112 VGND.t357 VGND.t356 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2663 XA.XIR[1].XIC[4].icell.Ien XThR.Tn[1].t68 VPWR.t1207 VPWR.t1206 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2664 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9].t69 VPWR.t386 VPWR.t385 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2665 VGND.t1528 Vbias.t247 XA.XIR[9].XIC[1].icell.SM VGND.t1527 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2666 XA.XIR[8].XIC[2].icell.Ien XThR.Tn[8].t71 VPWR.t725 VPWR.t724 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2667 XA.XIR[3].XIC[14].icell.Ien XThR.Tn[3].t70 VPWR.t378 VPWR.t377 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2668 XA.XIR[5].XIC[7].icell.SM XA.XIR[5].XIC[7].icell.Ien Iout.t64 VGND.t589 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2669 VPWR.t1854 XThC.XTB7.A XThC.XTB3.Y.t2 VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2670 XA.XIR[11].XIC[3].icell.Ien XThR.Tn[11].t73 VPWR.t95 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2671 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5].t71 XA.XIR[5].XIC[4].icell.Ien VGND.t1056 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2672 XA.XIR[8].XIC[8].icell.SM XA.XIR[8].XIC[8].icell.Ien Iout.t155 VGND.t1276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2673 XA.XIR[7].XIC[9].icell.SM XA.XIR[7].XIC[9].icell.Ien Iout.t134 VGND.t1180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2674 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13].t69 XA.XIR[13].XIC[1].icell.Ien VGND.t2558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2675 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9].t70 XA.XIR[9].XIC[4].icell.Ien VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2676 XThR.Tn[8].t8 XThR.XTBN.Y.t113 VPWR.t224 VPWR.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2677 VPWR.t1209 XThR.Tn[1].t69 XA.XIR[2].XIC[13].icell.PUM VPWR.t1208 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2678 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t2059 XA.XIR[4].XIC_dummy_right.icell.Ien VGND.t2633 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2679 XThR.Tn[5].t8 XThR.XTBN.Y.t114 a_n1049_5611# VPWR.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2680 a_n997_2891# XThR.XTB3.Y XThR.Tn[10].t0 VGND.t654 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2681 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8].t72 XA.XIR[8].XIC[5].icell.Ien VGND.t1107 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2682 XThR.XTB6.Y XThR.XTB7.B a_n1319_5611# VPWR.t1098 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2683 VPWR.t1352 VPWR.t1350 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1351 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2684 XA.XIR[2].XIC[7].icell.SM XA.XIR[2].XIC[7].icell.Ien Iout.t52 VGND.t397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2685 XA.XIR[11].XIC[3].icell.SM XA.XIR[11].XIC[3].icell.Ien Iout.t112 VGND.t1104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2686 a_n1049_7787# XThR.XTBN.Y.t115 XThR.Tn[1].t4 VPWR.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2687 a_3773_9615# XThC.XTBN.Y.t113 XThC.Tn[1].t5 VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2688 VPWR.t1097 XThR.XTB7.B XThR.XTB3.Y VPWR.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2689 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t2060 XA.XIR[7].XIC_dummy_left.icell.Ien VGND.t2634 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2690 XA.XIR[0].XIC[10].icell.PUM XThC.Tn[10].t42 XA.XIR[0].XIC[10].icell.Ien VPWR.t1310 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2691 a_4067_9615# XThC.XTB3.Y.t15 VPWR.t1311 VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2692 VGND.t1530 Vbias.t248 XA.XIR[3].XIC[0].icell.SM VGND.t1529 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2693 VPWR.t1312 XThC.XTB3.Y.t16 XThC.Tn[10].t5 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2694 VPWR.t1328 XThC.XTBN.Y.t114 XThC.Tn[14].t9 VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2695 XA.XIR[1].XIC[0].icell.Ien XThR.Tn[1].t70 VPWR.t1211 VPWR.t1210 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2696 VGND.t1777 VGND.t1775 XA.XIR[2].XIC_dummy_left.icell.SM VGND.t1776 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2697 XA.XIR[14].XIC[4].icell.PUM XThC.Tn[4].t43 XA.XIR[14].XIC[4].icell.Ien VPWR.t79 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2698 XA.XIR[15].XIC_15.icell.PDM VPWR.t2061 VGND.t2636 VGND.t2635 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2699 XA.XIR[10].XIC[5].icell.SM XA.XIR[10].XIC[5].icell.Ien Iout.t31 VGND.t202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2700 VGND.t2533 XThC.Tn[0].t40 XA.XIR[6].XIC[0].icell.PDM VGND.t2532 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2701 XA.XIR[14].XIC[13].icell.SM XA.XIR[14].XIC[13].icell.Ien Iout.t16 VGND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2702 VGND.t359 XThR.XTBN.Y.t116 XThR.Tn[0].t8 VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2703 XA.XIR[13].XIC[6].icell.SM XA.XIR[13].XIC[6].icell.Ien Iout.t68 VGND.t645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2704 VGND.t2201 XThC.XTB3.Y.t17 XThC.Tn[2].t9 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2705 XA.XIR[5].XIC[7].icell.PUM XThC.Tn[7].t38 XA.XIR[5].XIC[7].icell.Ien VPWR.t319 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2706 XThR.Tn[10].t8 XThR.XTBN.Y.t117 VPWR.t227 VPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2707 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[6].t71 VGND.t593 VGND.t592 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2708 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2062 VGND.t2638 VGND.t2637 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2709 XA.XIR[9].XIC[7].icell.PUM XThC.Tn[7].t39 XA.XIR[9].XIC[7].icell.Ien VPWR.t320 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2710 XA.XIR[5].XIC[2].icell.SM XA.XIR[5].XIC[2].icell.Ien Iout.t239 VGND.t2480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2711 XA.XIR[8].XIC[8].icell.PUM XThC.Tn[8].t42 XA.XIR[8].XIC[8].icell.Ien VPWR.t178 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2712 VGND.t1532 Vbias.t249 XA.XIR[0].XIC[11].icell.SM VGND.t1531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2713 VPWR.t758 XThC.XTB6.Y a_5949_9615# VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2714 XThR.Tn[1].t0 XThR.XTB2.Y VGND.t1392 VGND.t1391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2715 XA.XIR[4].XIC_15.icell.SM XA.XIR[4].XIC_15.icell.Ien Iout.t89 VGND.t865 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2716 VGND.t361 XThR.XTBN.Y.t118 a_n997_3755# VGND.t360 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2717 VPWR.t501 data[3].t1 XThC.XTBN.A VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2718 XA.XIR[8].XIC[3].icell.SM XA.XIR[8].XIC[3].icell.Ien Iout.t217 VGND.t2111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2719 a_2979_9615# XThC.XTB1.Y.t17 VPWR.t1118 VPWR.t1117 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2720 XThC.Tn[3].t4 XThC.XTBN.Y.t115 VGND.t2215 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2721 XA.XIR[2].XIC[13].icell.Ien XThR.Tn[2].t67 VPWR.t774 VPWR.t773 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2722 XA.XIR[7].XIC[4].icell.SM XA.XIR[7].XIC[4].icell.Ien Iout.t97 VGND.t882 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2723 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8].t73 XA.XIR[8].XIC[0].icell.Ien VGND.t1108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2724 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[3].t71 XA.XIR[3].XIC[12].icell.Ien VGND.t536 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2725 XA.XIR[7].XIC[14].icell.PUM XThC.Tn[14].t41 XA.XIR[7].XIC[14].icell.Ien VPWR.t1111 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2726 VPWR.t1889 XThR.Tn[13].t70 XA.XIR[14].XIC[12].icell.PUM VPWR.t1888 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2727 XA.XIR[2].XIC[2].icell.SM XA.XIR[2].XIC[2].icell.Ien Iout.t19 VGND.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2728 XA.XIR[10].XIC[8].icell.Ien XThR.Tn[10].t69 VPWR.t1917 VPWR.t1916 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2729 a_5949_10571# XThC.XTB7.B XThC.XTB6.Y VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2730 VPWR.t1213 XThR.Tn[1].t71 XA.XIR[2].XIC[6].icell.PUM VPWR.t1212 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2731 VPWR.t480 XThR.Tn[0].t71 XA.XIR[1].XIC[7].icell.PUM VPWR.t479 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2732 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[10].t70 VGND.t2671 VGND.t2670 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2733 XA.XIR[14].XIC[0].icell.PUM XThC.Tn[0].t41 XA.XIR[14].XIC[0].icell.Ien VPWR.t1882 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2734 XThR.Tn[13].t4 XThR.XTB6.Y VPWR.t115 VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2735 VPWR.t140 XThR.Tn[4].t69 XA.XIR[5].XIC[7].icell.PUM VPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2736 XA.XIR[13].XIC[10].icell.SM XA.XIR[13].XIC[10].icell.Ien Iout.t101 VGND.t938 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2737 a_n1049_7493# XThR.XTB3.Y VPWR.t639 VPWR.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2738 XA.XIR[0].XIC[5].icell.PUM XThC.Tn[5].t41 XA.XIR[0].XIC[5].icell.Ien VPWR.t1001 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2739 XA.XIR[5].XIC[11].icell.PUM XThC.Tn[11].t41 XA.XIR[5].XIC[11].icell.Ien VPWR.t282 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2740 XA.XIR[9].XIC[11].icell.PUM XThC.Tn[11].t42 XA.XIR[9].XIC[11].icell.Ien VPWR.t283 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2741 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[7].t67 VGND.t799 VGND.t798 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2742 VGND.t1774 VGND.t1772 XA.XIR[1].XIC_dummy_right.icell.SM VGND.t1773 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2743 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[2].t68 VGND.t62 VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2744 VGND.t1534 Vbias.t250 XA.XIR[0].XIC[9].icell.SM VGND.t1533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2745 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[10].t71 VGND.t2673 VGND.t2672 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2746 XA.XIR[10].XIC[0].icell.SM XA.XIR[10].XIC[0].icell.Ien Iout.t14 VGND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2747 VPWR.t1120 XThC.XTB1.Y.t18 XThC.Tn[8].t4 VPWR.t1119 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2748 VGND.t416 XThC.Tn[11].t43 XA.XIR[13].XIC[11].icell.PDM VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2749 XA.XIR[13].XIC[1].icell.SM XA.XIR[13].XIC[1].icell.Ien Iout.t99 VGND.t924 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2750 VGND.t1162 XThR.XTB5.Y XThR.Tn[4].t0 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2751 XThC.Tn[10].t8 XThC.XTBN.Y.t116 VPWR.t1329 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2752 VGND.t2217 XThC.XTBN.Y.t117 XThC.Tn[6].t8 VGND.t2216 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2753 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[3].t72 XA.XIR[3].XIC[10].icell.Ien VGND.t537 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2754 XA.XIR[5].XIC[2].icell.PUM XThC.Tn[2].t41 XA.XIR[5].XIC[2].icell.Ien VPWR.t1278 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2755 VPWR.t184 XThR.Tn[14].t71 XA.XIR[15].XIC[9].icell.PUM VPWR.t183 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2756 VPWR.t1891 XThR.Tn[13].t71 XA.XIR[14].XIC[10].icell.PUM VPWR.t1890 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2757 XA.XIR[9].XIC[2].icell.PUM XThC.Tn[2].t42 XA.XIR[9].XIC[2].icell.Ien VPWR.t951 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2758 XA.XIR[4].XIC[14].icell.PUM XThC.Tn[14].t42 XA.XIR[4].XIC[14].icell.Ien VPWR.t1112 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2759 XA.XIR[8].XIC[3].icell.PUM XThC.Tn[3].t43 XA.XIR[8].XIC[3].icell.Ien VPWR.t132 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2760 XA.XIR[3].XIC_15.icell.PUM VPWR.t1348 XA.XIR[3].XIC_15.icell.Ien VPWR.t1349 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2761 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[4].t70 VGND.t246 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2762 VGND.t1536 Vbias.t251 XA.XIR[5].XIC[6].icell.SM VGND.t1535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2763 VGND.t1421 XThC.Tn[1].t43 XA.XIR[10].XIC[1].icell.PDM VGND.t1420 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2764 VGND.t2640 VPWR.t2063 XA.XIR[1].XIC_dummy_right.icell.PDM VGND.t2639 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2765 VGND.t1574 XThC.Tn[5].t42 XA.XIR[5].XIC[5].icell.PDM VGND.t1573 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2766 VGND.t1444 XThC.Tn[2].t43 XA.XIR[13].XIC[2].icell.PDM VGND.t1443 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2767 VGND.t1576 XThC.Tn[5].t43 XA.XIR[9].XIC[5].icell.PDM VGND.t1575 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2768 VPWR.t482 XThR.Tn[0].t72 XA.XIR[1].XIC[11].icell.PUM VPWR.t481 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2769 XA.XIR[7].XIC[8].icell.Ien XThR.Tn[7].t68 VPWR.t602 VPWR.t601 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2770 VPWR.t158 XThC.XTB4.Y.t17 a_4861_9615# VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2771 VPWR.t1203 XThR.Tn[4].t71 XA.XIR[5].XIC[11].icell.PUM VPWR.t1202 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2772 XA.XIR[14].XIC[12].icell.Ien XThR.Tn[14].t72 VPWR.t186 VPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2773 XA.XIR[15].XIC[11].icell.PDM VPWR.t2064 XA.XIR[15].XIC[11].icell.Ien VGND.t2641 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2774 VGND.t2643 VPWR.t2065 XA.XIR[11].XIC_15.icell.PDM VGND.t2642 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2775 XA.XIR[2].XIC[13].icell.PUM XThC.Tn[13].t42 XA.XIR[2].XIC[13].icell.Ien VPWR.t1772 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2776 VGND.t1538 Vbias.t252 XA.XIR[4].XIC[12].icell.SM VGND.t1537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2777 XThR.Tn[6].t4 XThR.XTBN.Y.t119 a_n1049_5317# VPWR.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2778 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1346 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1347 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2779 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t0 VGND.t1297 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2780 XA.XIR[2].XIC[6].icell.Ien XThR.Tn[2].t69 VPWR.t772 VPWR.t771 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2781 XA.XIR[10].XIC[3].icell.Ien XThR.Tn[10].t72 VPWR.t1919 VPWR.t1918 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2782 VGND.t1540 Vbias.t253 XA.XIR[7].XIC[13].icell.SM VGND.t1539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2783 XA.XIR[6].XIC[14].icell.Ien XThR.Tn[6].t72 VPWR.t442 VPWR.t441 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2784 VGND.t2219 XThC.XTBN.Y.t118 a_10915_9569# VGND.t2218 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2785 VPWR.t1215 XThR.Tn[1].t72 XA.XIR[2].XIC[1].icell.PUM VPWR.t1214 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2786 XA.XIR[5].XIC_15.icell.Ien XThR.Tn[5].t72 VPWR.t698 VPWR.t697 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2787 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[10].t73 VGND.t2675 VGND.t2674 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2788 VGND.t1562 XThC.Tn[12].t42 XA.XIR[7].XIC[12].icell.PDM VGND.t1561 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2789 VGND.t1542 Vbias.t254 XA.XIR[6].XIC[14].icell.SM VGND.t1541 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2790 VPWR.t484 XThR.Tn[0].t73 XA.XIR[1].XIC[2].icell.PUM VPWR.t483 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2791 XA.XIR[9].XIC_15.icell.Ien XThR.Tn[9].t71 VPWR.t388 VPWR.t387 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2792 VPWR.t1205 XThR.Tn[4].t72 XA.XIR[5].XIC[2].icell.PUM VPWR.t1204 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2793 VPWR.t1048 VGND.t2703 XA.XIR[0].XIC[14].icell.PUM VPWR.t1047 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2794 XA.XIR[15].XIC[2].icell.PDM VPWR.t2066 XA.XIR[15].XIC[2].icell.Ien VGND.t2644 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2795 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[2].t70 XA.XIR[2].XIC[9].icell.Ien VGND.t682 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2796 XThC.Tn[1].t4 XThC.XTBN.Y.t119 a_3773_9615# VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2797 XA.XIR[1].XIC[7].icell.SM XA.XIR[1].XIC[7].icell.Ien Iout.t180 VGND.t1519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2798 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13].t72 XA.XIR[13].XIC_15.icell.Ien VGND.t664 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2799 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[2].t71 VGND.t681 VGND.t680 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2800 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[4].t73 VGND.t2087 VGND.t2086 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2801 VGND.t1544 Vbias.t255 XA.XIR[0].XIC[4].icell.SM VGND.t1543 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2802 XA.XIR[4].XIC[8].icell.SM XA.XIR[4].XIC[8].icell.Ien Iout.t102 VGND.t939 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2803 XThC.Tn[14].t8 XThC.XTBN.Y.t120 VPWR.t448 VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2804 VGND.t1546 Vbias.t256 XA.XIR[5].XIC[10].icell.SM VGND.t1545 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2805 VGND.t1040 Vbias.t257 XA.XIR[13].XIC[7].icell.SM VGND.t1039 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2806 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2067 XA.XIR[0].XIC_dummy_right.icell.Ien VGND.t2645 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2807 VGND.t483 XThC.Tn[6].t42 XA.XIR[13].XIC[6].icell.PDM VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2808 VGND.t363 XThR.XTBN.Y.t120 a_n997_715# VGND.t362 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2809 VPWR.t1345 VPWR.t1343 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1344 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2810 XA.XIR[14].XIC[10].icell.Ien XThR.Tn[14].t73 VPWR.t188 VPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2811 VPWR.t478 XThR.Tn[13].t73 XA.XIR[14].XIC[5].icell.PUM VPWR.t477 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2812 VPWR.t988 XThR.XTB7.Y XThR.Tn[14].t4 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2813 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12].t70 XA.XIR[12].XIC[11].icell.Ien VGND.t1412 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2814 VGND.t1771 VGND.t1769 XA.XIR[1].XIC_dummy_left.icell.SM VGND.t1770 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2815 VGND.t1042 Vbias.t258 XA.XIR[5].XIC[1].icell.SM VGND.t1041 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2816 XA.XIR[9].XIC[5].icell.SM XA.XIR[9].XIC[5].icell.Ien Iout.t39 VGND.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2817 XThR.XTB6.A data[5].t5 VGND.t769 VGND.t768 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2818 XThR.Tn[0].t4 XThR.XTBN.Y.t121 a_n1049_8581# VPWR.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2819 VGND.t2535 XThC.Tn[0].t42 XA.XIR[5].XIC[0].icell.PDM VGND.t2534 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2820 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[12].t71 VGND.t1414 VGND.t1413 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2821 a_5949_9615# XThC.XTB6.Y VPWR.t757 VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2822 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[12].t72 VGND.t1416 VGND.t1415 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2823 XA.XIR[12].XIC[6].icell.SM XA.XIR[12].XIC[6].icell.Ien Iout.t45 VGND.t266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2824 VGND.t2537 XThC.Tn[0].t43 XA.XIR[9].XIC[0].icell.PDM VGND.t2536 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2825 VGND.t2200 XThC.Tn[10].t43 XA.XIR[7].XIC[10].icell.PDM VGND.t2199 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2826 XA.XIR[7].XIC[3].icell.Ien XThR.Tn[7].t69 VPWR.t604 VPWR.t603 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2827 VGND.t601 XThC.XTBN.Y.t121 a_10051_9569# VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2828 VGND.t1044 Vbias.t259 XA.XIR[3].XIC[14].icell.SM VGND.t1043 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2829 VGND.t1564 XThC.Tn[12].t43 XA.XIR[4].XIC[12].icell.PDM VGND.t1563 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2830 VGND.t2274 XThC.Tn[13].t43 XA.XIR[3].XIC[13].icell.PDM VGND.t2273 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2831 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2068 XA.XIR[3].XIC_dummy_left.icell.Ien VGND.t2646 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2832 XA.XIR[15].XIC[6].icell.PDM VPWR.t2069 XA.XIR[15].XIC[6].icell.Ien VGND.t2647 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2833 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12].t73 XA.XIR[12].XIC[2].icell.Ien VGND.t1417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2834 XA.XIR[0].XIC[9].icell.PDM VGND.t1766 VGND.t1768 VGND.t1767 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2835 VPWR.t449 XThC.XTBN.Y.t122 XThC.Tn[11].t1 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2836 VGND.t603 XThC.XTBN.Y.t123 a_7651_9569# VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2837 XA.XIR[2].XIC[1].icell.Ien XThR.Tn[2].t72 VPWR.t770 VPWR.t769 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2838 Vbias.t4 bias[1].t0 VPWR.t694 VPWR.t693 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
X2839 XA.XIR[11].XIC[12].icell.SM XA.XIR[11].XIC[12].icell.Ien Iout.t22 VGND.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2840 XA.XIR[1].XIC[13].icell.Ien XThR.Tn[1].t73 VPWR.t1217 VPWR.t1216 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2841 XThR.Tn[2].t0 XThR.XTBN.Y.t122 VGND.t343 VGND.t342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2842 VPWR.t987 XThR.XTB7.Y a_n1049_5317# VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2843 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout VGND.t767 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2844 VGND.t1046 Vbias.t260 XA.XIR[15].XIC_15.icell.SM VGND.t1045 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2845 a_8739_9569# XThC.XTB3.Y.t18 XThC.Tn[10].t6 VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2846 XA.XIR[2].XIC[6].icell.PUM XThC.Tn[6].t43 XA.XIR[2].XIC[6].icell.Ien VPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2847 VGND.t1948 XThC.Tn[14].t43 XA.XIR[15].XIC[14].icell.PDM VGND.t1947 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2848 VGND.t318 XThC.Tn[8].t43 XA.XIR[15].XIC[8].icell.PDM VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2849 VPWR.t215 XThR.XTBN.Y.t123 XThR.Tn[12].t8 VPWR.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2850 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[2].t73 XA.XIR[2].XIC[4].icell.Ien VGND.t679 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2851 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6].t73 XA.XIR[6].XIC[12].icell.Ien VGND.t594 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2852 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5].t73 XA.XIR[5].XIC[13].icell.Ien VGND.t1057 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2853 XA.XIR[1].XIC[2].icell.SM XA.XIR[1].XIC[2].icell.Ien Iout.t63 VGND.t561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2854 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9].t72 XA.XIR[9].XIC[13].icell.Ien VGND.t544 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2855 VPWR.t1342 VPWR.t1340 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1341 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2856 VGND.t2132 XThC.Tn[9].t43 XA.XIR[2].XIC[9].icell.PDM VGND.t2131 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2857 XA.XIR[4].XIC[3].icell.SM XA.XIR[4].XIC[3].icell.Ien Iout.t151 VGND.t1242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2858 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[9].t73 VGND.t546 VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2859 VGND.t1048 Vbias.t261 XA.XIR[13].XIC[2].icell.SM VGND.t1047 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2860 VPWR.t380 XThR.Tn[3].t73 XA.XIR[4].XIC[7].icell.PUM VPWR.t379 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
R0 VGND.n3019 VGND.n3018 15660.6
R1 VGND.n196 VGND.n195 13477
R2 VGND.n3018 VGND.n7 11578
R3 VGND.n195 VGND.n7 10429.6
R4 VGND.n3012 VGND.n8 9309.26
R5 VGND.n200 VGND.n199 9223.7
R6 VGND.n198 VGND.n197 9223.7
R7 VGND.n197 VGND.n196 9223.7
R8 VGND.n2969 VGND.n200 9223.7
R9 VGND.n2969 VGND.n2968 7447.41
R10 VGND.n2249 VGND.n2248 7387.65
R11 VGND.n2250 VGND.n2249 7387.65
R12 VGND.n2285 VGND.n2284 7387.65
R13 VGND.n3017 VGND.n3016 7387.65
R14 VGND.n3016 VGND.n3015 7387.65
R15 VGND.n3015 VGND.n3014 7387.65
R16 VGND.n3014 VGND.n3013 7387.65
R17 VGND.n3013 VGND.n3012 7387.65
R18 VGND.n2351 VGND.n2285 6674.35
R19 VGND.n1386 VGND.t2248 6324.96
R20 VGND.n199 VGND.n198 5231.11
R21 VGND.n1336 VGND.t2364 5168.13
R22 VGND.n2967 VGND.n8 5074.71
R23 VGND.n3018 VGND.n3017 5063.19
R24 VGND.n1154 VGND.n806 4539.15
R25 VGND VGND.n8 4240.58
R26 VGND.t1770 VGND.t883 4212.19
R27 VGND.t1776 VGND.t2079 4212.19
R28 VGND.t1782 VGND.t1181 4212.19
R29 VGND.t1869 VGND.t556 4212.19
R30 VGND.t1875 VGND.t557 4212.19
R31 VGND.t1788 VGND.t660 4212.19
R32 VGND.t1830 VGND.t1077 4212.19
R33 VGND.t1488 VGND.t1881 4212.19
R34 VGND.t177 VGND.t1803 4212.19
R35 VGND.t1484 VGND.t1848 4212.19
R36 VGND.t466 VGND.t1887 4212.19
R37 VGND.t2487 VGND.t1899 4212.19
R38 VGND.t942 VGND.t1815 4212.19
R39 VGND.t1407 VGND.t1857 4212.19
R40 VGND.n2919 VGND.n222 4077.12
R41 VGND.n1340 VGND.n1338 3417.39
R42 VGND.n1340 VGND.n1339 3417.39
R43 VGND.n1388 VGND.n1387 3417.39
R44 VGND.n2180 VGND.n504 3417.39
R45 VGND.n503 VGND.n473 3417.39
R46 VGND.n2353 VGND.n2352 3417.39
R47 VGND.n2920 VGND.n2919 3331.79
R48 VGND.n2921 VGND.n2920 3331.79
R49 VGND.n2922 VGND.n2921 3331.79
R50 VGND.n2923 VGND.n2922 3331.79
R51 VGND.n2924 VGND.n2923 3331.79
R52 VGND.n2925 VGND.n2924 3331.79
R53 VGND.n2926 VGND.n2925 3331.79
R54 VGND.n2927 VGND.n2926 3331.79
R55 VGND.n2928 VGND.n2927 3331.79
R56 VGND.n2929 VGND.n2928 3331.79
R57 VGND.n2930 VGND.n2929 3331.79
R58 VGND.n2931 VGND.n2930 3331.79
R59 VGND.n2932 VGND.n2931 3331.79
R60 VGND.n2933 VGND.n2932 3331.79
R61 VGND.n2934 VGND.n2933 3331.79
R62 VGND.n1339 VGND.n806 3273.91
R63 VGND.n2181 VGND.n539 3265.22
R64 VGND.n2934 VGND.n201 2725.63
R65 VGND.n197 VGND.t451 2655.17
R66 VGND.n196 VGND.t391 2655.17
R67 VGND.n2353 VGND.n2285 2517.39
R68 VGND.t2075 VGND.n201 2334.15
R69 VGND.t2587 VGND.n2701 2307.69
R70 VGND.n359 VGND.t2324 2307.69
R71 VGND.n360 VGND.t2311 2307.69
R72 VGND.n370 VGND.t2646 2307.69
R73 VGND.n371 VGND.t2579 2307.69
R74 VGND.n381 VGND.t2298 2307.69
R75 VGND.n382 VGND.t1662 2307.69
R76 VGND.t2634 VGND.n327 2307.69
R77 VGND.n2705 VGND.t2360 2307.69
R78 VGND.n2728 VGND.t2299 2307.69
R79 VGND.n2738 VGND.t2632 2307.69
R80 VGND.t2622 VGND.n2737 2307.69
R81 VGND.n2731 VGND.t2351 2307.69
R82 VGND.n2776 VGND.t1701 2307.69
R83 VGND.t1678 VGND.n2775 2307.69
R84 VGND.n2943 VGND.t2348 2307.69
R85 VGND.t1821 VGND.n2703 2280.49
R86 VGND.n3020 VGND.n5 2229.43
R87 VGND.n3020 VGND.n6 2229.43
R88 VGND.n2348 VGND.n6 2229.43
R89 VGND.n2348 VGND.n5 2229.43
R90 VGND.n1338 VGND.n1337 2173.91
R91 VGND.n2704 VGND.t145 2132.93
R92 VGND.n2701 VGND.t1665 2123.08
R93 VGND.t2581 VGND.n359 2123.08
R94 VGND.n360 VGND.t2559 2123.08
R95 VGND.t1663 VGND.n370 2123.08
R96 VGND.n371 VGND.t1652 2123.08
R97 VGND.t2628 VGND.n381 2123.08
R98 VGND.n382 VGND.t2300 2123.08
R99 VGND.n2705 VGND.t2624 2123.08
R100 VGND.t2354 VGND.n2728 2123.08
R101 VGND.n2738 VGND.t2342 2123.08
R102 VGND.n2737 VGND.t1681 2123.08
R103 VGND.n2731 VGND.t2611 2123.08
R104 VGND.n2776 VGND.t2330 2123.08
R105 VGND.n2775 VGND.t1695 2123.08
R106 VGND.n2704 VGND.t1845 2079.27
R107 VGND.t883 VGND.t1821 2012.2
R108 VGND.t2079 VGND.t1770 2012.2
R109 VGND.t1181 VGND.t1776 2012.2
R110 VGND.t556 VGND.t1782 2012.2
R111 VGND.t557 VGND.t1869 2012.2
R112 VGND.t660 VGND.t1875 2012.2
R113 VGND.t1077 VGND.t1788 2012.2
R114 VGND.t145 VGND.t1830 2012.2
R115 VGND.t1845 VGND.t1488 2012.2
R116 VGND.t1881 VGND.t177 2012.2
R117 VGND.t1803 VGND.t1484 2012.2
R118 VGND.t1848 VGND.t466 2012.2
R119 VGND.t1887 VGND.t2487 2012.2
R120 VGND.t1899 VGND.t942 2012.2
R121 VGND.t1815 VGND.t1407 2012.2
R122 VGND.t1857 VGND.t2075 2012.2
R123 VGND.n199 VGND 1997.7
R124 VGND.n200 VGND 1997.7
R125 VGND VGND.n2969 1997.7
R126 VGND.n2968 VGND.n2944 1907.51
R127 VGND.n2284 VGND.n2251 1831.57
R128 VGND.n198 VGND.t354 1807.04
R129 VGND.n2970 VGND.t2100 1785.51
R130 VGND.n2352 VGND.n2351 1760.87
R131 VGND.n2702 VGND.t2312 1738.46
R132 VGND.n2250 VGND.n504 1691.3
R133 VGND.n2351 VGND.n2350 1656.52
R134 VGND.t1402 VGND.n66 1618.39
R135 VGND.n3011 VGND.t651 1618.39
R136 VGND.n2971 VGND.t212 1618.39
R137 VGND.n2702 VGND.n7 1604.17
R138 VGND.n2350 VGND.n328 1517.39
R139 VGND.n195 VGND.t401 1517.24
R140 VGND.n2248 VGND.n540 1513.49
R141 VGND.t2277 VGND.n2704 1507.69
R142 VGND.n2703 VGND.n2702 1441.28
R143 VGND.n1386 VGND.n540 1370.36
R144 VGND.t2312 VGND.t1667 1353.85
R145 VGND.t1667 VGND.t2587 1353.85
R146 VGND.t2583 VGND.t1665 1353.85
R147 VGND.t2324 VGND.t2583 1353.85
R148 VGND.t2316 VGND.t2581 1353.85
R149 VGND.t2311 VGND.t2316 1353.85
R150 VGND.t2559 VGND.t2296 1353.85
R151 VGND.t2296 VGND.t2646 1353.85
R152 VGND.t1660 VGND.t1663 1353.85
R153 VGND.t2579 VGND.t1660 1353.85
R154 VGND.t1652 VGND.t2561 1353.85
R155 VGND.t2561 VGND.t2298 1353.85
R156 VGND.t2358 VGND.t2628 1353.85
R157 VGND.t1662 VGND.t2358 1353.85
R158 VGND.t2300 VGND.t1656 1353.85
R159 VGND.t1656 VGND.t2634 1353.85
R160 VGND.t2630 VGND.t2277 1353.85
R161 VGND.t2360 VGND.t2630 1353.85
R162 VGND.t2624 VGND.t2563 1353.85
R163 VGND.t2563 VGND.t2299 1353.85
R164 VGND.t2279 VGND.t2354 1353.85
R165 VGND.t2632 VGND.t2279 1353.85
R166 VGND.t2342 VGND.t1697 1353.85
R167 VGND.t1697 VGND.t2622 1353.85
R168 VGND.t2356 VGND.t1681 1353.85
R169 VGND.t2351 VGND.t2356 1353.85
R170 VGND.t2611 VGND.t2344 1353.85
R171 VGND.t2344 VGND.t1701 1353.85
R172 VGND.t2330 VGND.t2328 1353.85
R173 VGND.t2328 VGND.t1678 1353.85
R174 VGND.t1695 VGND.t2615 1353.85
R175 VGND.t2615 VGND.t2348 1353.85
R176 VGND.n2944 VGND.n201 1301.35
R177 VGND.n2703 VGND.n328 1278.26
R178 VGND.t1767 VGND.n540 1270.28
R179 VGND.n1127 VGND.t600 1268.93
R180 VGND.n1127 VGND.t366 1268.93
R181 VGND.n502 VGND.t63 1253.59
R182 VGND.t551 VGND.n502 1253.59
R183 VGND.n2283 VGND.t1136 1253.59
R184 VGND.t364 VGND.n2283 1253.59
R185 VGND.n538 VGND.t114 1253.59
R186 VGND.t548 VGND.n538 1253.59
R187 VGND.n2247 VGND.t66 1253.59
R188 VGND.t602 VGND.n2247 1253.59
R189 VGND.n1385 VGND.t488 1253.59
R190 VGND.t330 VGND.n1385 1253.59
R191 VGND.n1337 VGND.n1336 1243.48
R192 VGND.n2251 VGND.t1812 1237.71
R193 VGND.n66 VGND.t238 1213.79
R194 VGND.n2967 VGND.n2966 1198.25
R195 VGND.n1155 VGND.n1154 1198.25
R196 VGND.n2943 VGND.n2942 1180.79
R197 VGND.n2936 VGND.n2935 1180.79
R198 VGND.n2534 VGND.n208 1180.79
R199 VGND.n2529 VGND.n209 1180.79
R200 VGND.n2817 VGND.n210 1180.79
R201 VGND.n1989 VGND.n211 1180.79
R202 VGND.n1996 VGND.n212 1180.79
R203 VGND.n2842 VGND.n213 1180.79
R204 VGND.n1829 VGND.n214 1180.79
R205 VGND.n1836 VGND.n215 1180.79
R206 VGND.n2867 VGND.n216 1180.79
R207 VGND.n1655 VGND.n217 1180.79
R208 VGND.n1650 VGND.n218 1180.79
R209 VGND.n2892 VGND.n219 1180.79
R210 VGND.n1607 VGND.n220 1180.79
R211 VGND.n2912 VGND.n221 1180.79
R212 VGND.n1282 VGND.n222 1180.79
R213 VGND.n2918 VGND.n2917 1180.79
R214 VGND.n1335 VGND.n1334 1180.46
R215 VGND.n929 VGND.n890 1180.46
R216 VGND.n934 VGND.n933 1180.46
R217 VGND.n939 VGND.n938 1180.46
R218 VGND.n944 VGND.n943 1180.46
R219 VGND.n949 VGND.n948 1180.46
R220 VGND.n954 VGND.n953 1180.46
R221 VGND.n959 VGND.n958 1180.46
R222 VGND.n964 VGND.n963 1180.46
R223 VGND.n969 VGND.n968 1180.46
R224 VGND.n974 VGND.n973 1180.46
R225 VGND.n979 VGND.n978 1180.46
R226 VGND.n984 VGND.n983 1180.46
R227 VGND.n989 VGND.n988 1180.46
R228 VGND.n991 VGND.n990 1180.46
R229 VGND.n1279 VGND.n1278 1180.46
R230 VGND.n1277 VGND.n1276 1180.46
R231 VGND.n1234 VGND.n1233 1180.46
R232 VGND.n1239 VGND.n1238 1180.46
R233 VGND.n1241 VGND.n1240 1180.46
R234 VGND.n1246 VGND.n1245 1180.46
R235 VGND.n1248 VGND.n1247 1180.46
R236 VGND.n1220 VGND.n1219 1180.46
R237 VGND.n1209 VGND.n1208 1180.46
R238 VGND.n1207 VGND.n1206 1180.46
R239 VGND.n1190 VGND.n1189 1180.46
R240 VGND.n1188 VGND.n1187 1180.46
R241 VGND.n1177 VGND.n1176 1180.46
R242 VGND.n1175 VGND.n1174 1180.46
R243 VGND.n1167 VGND.n1166 1180.46
R244 VGND.n2775 VGND.n2774 1180.46
R245 VGND.n2777 VGND.n2776 1180.46
R246 VGND.n2732 VGND.n2731 1180.46
R247 VGND.n2737 VGND.n2736 1180.46
R248 VGND.n2739 VGND.n2738 1180.46
R249 VGND.n2728 VGND.n2727 1180.46
R250 VGND.n2706 VGND.n2705 1180.46
R251 VGND.n388 VGND.n327 1180.46
R252 VGND.n383 VGND.n382 1180.46
R253 VGND.n381 VGND.n380 1180.46
R254 VGND.n372 VGND.n371 1180.46
R255 VGND.n370 VGND.n369 1180.46
R256 VGND.n361 VGND.n360 1180.46
R257 VGND.n359 VGND.n333 1180.46
R258 VGND.n2701 VGND.n2700 1180.46
R259 VGND.n2641 VGND.n2640 1180.46
R260 VGND.n2646 VGND.n2645 1180.46
R261 VGND.n2651 VGND.n2650 1180.46
R262 VGND.n2656 VGND.n2655 1180.46
R263 VGND.n2661 VGND.n2660 1180.46
R264 VGND.n2666 VGND.n2665 1180.46
R265 VGND.n2671 VGND.n2670 1180.46
R266 VGND.n2673 VGND.n2672 1180.46
R267 VGND.n2717 VGND.n2716 1180.46
R268 VGND.n2719 VGND.n2718 1180.46
R269 VGND.n2750 VGND.n2749 1180.46
R270 VGND.n2757 VGND.n2756 1180.46
R271 VGND.n2755 VGND.n2754 1180.46
R272 VGND.n2790 VGND.n2789 1180.46
R273 VGND.n2792 VGND.n2791 1180.46
R274 VGND.n2345 VGND.n2344 1180.46
R275 VGND.n2340 VGND.n2339 1180.46
R276 VGND.n2335 VGND.n2334 1180.46
R277 VGND.n2330 VGND.n2329 1180.46
R278 VGND.n2325 VGND.n2324 1180.46
R279 VGND.n2320 VGND.n2319 1180.46
R280 VGND.n2315 VGND.n2314 1180.46
R281 VGND.n2310 VGND.n2309 1180.46
R282 VGND.n2305 VGND.n2304 1180.46
R283 VGND.n2300 VGND.n2299 1180.46
R284 VGND.n2295 VGND.n2294 1180.46
R285 VGND.n2290 VGND.n2289 1180.46
R286 VGND.n2545 VGND.n2544 1180.46
R287 VGND.n2543 VGND.n2542 1180.46
R288 VGND.n2538 VGND.n2537 1180.46
R289 VGND.n2355 VGND.n2354 1180.46
R290 VGND.n2379 VGND.n2378 1180.46
R291 VGND.n2381 VGND.n2380 1180.46
R292 VGND.n2405 VGND.n2404 1180.46
R293 VGND.n2407 VGND.n2406 1180.46
R294 VGND.n2431 VGND.n2430 1180.46
R295 VGND.n2433 VGND.n2432 1180.46
R296 VGND.n2457 VGND.n2456 1180.46
R297 VGND.n2459 VGND.n2458 1180.46
R298 VGND.n2483 VGND.n2482 1180.46
R299 VGND.n2485 VGND.n2484 1180.46
R300 VGND.n2514 VGND.n2513 1180.46
R301 VGND.n2519 VGND.n2518 1180.46
R302 VGND.n2524 VGND.n2523 1180.46
R303 VGND.n2526 VGND.n2525 1180.46
R304 VGND.n2366 VGND.n2365 1180.46
R305 VGND.n2368 VGND.n2367 1180.46
R306 VGND.n2392 VGND.n2391 1180.46
R307 VGND.n2394 VGND.n2393 1180.46
R308 VGND.n2418 VGND.n2417 1180.46
R309 VGND.n2420 VGND.n2419 1180.46
R310 VGND.n2444 VGND.n2443 1180.46
R311 VGND.n2446 VGND.n2445 1180.46
R312 VGND.n2470 VGND.n2469 1180.46
R313 VGND.n2472 VGND.n2471 1180.46
R314 VGND.n2496 VGND.n2495 1180.46
R315 VGND.n2503 VGND.n2502 1180.46
R316 VGND.n2501 VGND.n2500 1180.46
R317 VGND.n2812 VGND.n2811 1180.46
R318 VGND.n2814 VGND.n2813 1180.46
R319 VGND.n1913 VGND.n1912 1180.46
R320 VGND.n1915 VGND.n1914 1180.46
R321 VGND.n1924 VGND.n1923 1180.46
R322 VGND.n1926 VGND.n1925 1180.46
R323 VGND.n1935 VGND.n1934 1180.46
R324 VGND.n1937 VGND.n1936 1180.46
R325 VGND.n1946 VGND.n1945 1180.46
R326 VGND.n1948 VGND.n1947 1180.46
R327 VGND.n1957 VGND.n1956 1180.46
R328 VGND.n1959 VGND.n1958 1180.46
R329 VGND.n1968 VGND.n1967 1180.46
R330 VGND.n1970 VGND.n1969 1180.46
R331 VGND.n1979 VGND.n1978 1180.46
R332 VGND.n1984 VGND.n1983 1180.46
R333 VGND.n1986 VGND.n1985 1180.46
R334 VGND.n599 VGND.n598 1180.46
R335 VGND.n2060 VGND.n2059 1180.46
R336 VGND.n2058 VGND.n2057 1180.46
R337 VGND.n2053 VGND.n2052 1180.46
R338 VGND.n2048 VGND.n2047 1180.46
R339 VGND.n2043 VGND.n2042 1180.46
R340 VGND.n2038 VGND.n2037 1180.46
R341 VGND.n2033 VGND.n2032 1180.46
R342 VGND.n2028 VGND.n2027 1180.46
R343 VGND.n2023 VGND.n2022 1180.46
R344 VGND.n2018 VGND.n2017 1180.46
R345 VGND.n2013 VGND.n2012 1180.46
R346 VGND.n2008 VGND.n2007 1180.46
R347 VGND.n2003 VGND.n2002 1180.46
R348 VGND.n602 VGND.n601 1180.46
R349 VGND.n2072 VGND.n2071 1180.46
R350 VGND.n2077 VGND.n2076 1180.46
R351 VGND.n2082 VGND.n2081 1180.46
R352 VGND.n2087 VGND.n2086 1180.46
R353 VGND.n2092 VGND.n2091 1180.46
R354 VGND.n2097 VGND.n2096 1180.46
R355 VGND.n2102 VGND.n2101 1180.46
R356 VGND.n2107 VGND.n2106 1180.46
R357 VGND.n2112 VGND.n2111 1180.46
R358 VGND.n2117 VGND.n2116 1180.46
R359 VGND.n2122 VGND.n2121 1180.46
R360 VGND.n2129 VGND.n2128 1180.46
R361 VGND.n2127 VGND.n2126 1180.46
R362 VGND.n2837 VGND.n2836 1180.46
R363 VGND.n2839 VGND.n2838 1180.46
R364 VGND.n2179 VGND.n2178 1180.46
R365 VGND.n1754 VGND.n550 1180.46
R366 VGND.n1764 VGND.n1763 1180.46
R367 VGND.n1766 VGND.n1765 1180.46
R368 VGND.n1775 VGND.n1774 1180.46
R369 VGND.n1777 VGND.n1776 1180.46
R370 VGND.n1786 VGND.n1785 1180.46
R371 VGND.n1788 VGND.n1787 1180.46
R372 VGND.n1797 VGND.n1796 1180.46
R373 VGND.n1799 VGND.n1798 1180.46
R374 VGND.n1808 VGND.n1807 1180.46
R375 VGND.n1810 VGND.n1809 1180.46
R376 VGND.n1819 VGND.n1818 1180.46
R377 VGND.n1824 VGND.n1823 1180.46
R378 VGND.n1826 VGND.n1825 1180.46
R379 VGND.n1681 VGND.n1680 1180.46
R380 VGND.n1683 VGND.n1682 1180.46
R381 VGND.n1692 VGND.n1691 1180.46
R382 VGND.n1697 VGND.n1696 1180.46
R383 VGND.n1702 VGND.n1701 1180.46
R384 VGND.n1707 VGND.n1706 1180.46
R385 VGND.n1712 VGND.n1711 1180.46
R386 VGND.n1717 VGND.n1716 1180.46
R387 VGND.n1722 VGND.n1721 1180.46
R388 VGND.n1727 VGND.n1726 1180.46
R389 VGND.n1732 VGND.n1731 1180.46
R390 VGND.n1850 VGND.n1849 1180.46
R391 VGND.n1848 VGND.n1847 1180.46
R392 VGND.n1843 VGND.n1842 1180.46
R393 VGND.n1735 VGND.n1734 1180.46
R394 VGND.n672 VGND.n671 1180.46
R395 VGND.n677 VGND.n676 1180.46
R396 VGND.n682 VGND.n681 1180.46
R397 VGND.n687 VGND.n686 1180.46
R398 VGND.n692 VGND.n691 1180.46
R399 VGND.n697 VGND.n696 1180.46
R400 VGND.n702 VGND.n701 1180.46
R401 VGND.n707 VGND.n706 1180.46
R402 VGND.n712 VGND.n711 1180.46
R403 VGND.n717 VGND.n716 1180.46
R404 VGND.n722 VGND.n721 1180.46
R405 VGND.n729 VGND.n728 1180.46
R406 VGND.n727 VGND.n726 1180.46
R407 VGND.n2862 VGND.n2861 1180.46
R408 VGND.n2864 VGND.n2863 1180.46
R409 VGND.n1355 VGND.n1354 1180.46
R410 VGND.n877 VGND.n876 1180.46
R411 VGND.n872 VGND.n871 1180.46
R412 VGND.n821 VGND.n808 1180.46
R413 VGND.n826 VGND.n825 1180.46
R414 VGND.n831 VGND.n830 1180.46
R415 VGND.n836 VGND.n835 1180.46
R416 VGND.n841 VGND.n840 1180.46
R417 VGND.n846 VGND.n845 1180.46
R418 VGND.n851 VGND.n850 1180.46
R419 VGND.n858 VGND.n857 1180.46
R420 VGND.n856 VGND.n855 1180.46
R421 VGND.n1666 VGND.n1665 1180.46
R422 VGND.n1664 VGND.n1663 1180.46
R423 VGND.n1659 VGND.n1658 1180.46
R424 VGND.n1393 VGND.n1392 1180.46
R425 VGND.n1398 VGND.n1397 1180.46
R426 VGND.n1400 VGND.n1399 1180.46
R427 VGND.n1493 VGND.n1492 1180.46
R428 VGND.n1495 VGND.n1494 1180.46
R429 VGND.n1519 VGND.n1518 1180.46
R430 VGND.n1521 VGND.n1520 1180.46
R431 VGND.n1545 VGND.n1544 1180.46
R432 VGND.n1550 VGND.n1549 1180.46
R433 VGND.n1557 VGND.n1556 1180.46
R434 VGND.n1555 VGND.n1554 1180.46
R435 VGND.n1635 VGND.n1634 1180.46
R436 VGND.n1640 VGND.n1639 1180.46
R437 VGND.n1645 VGND.n1644 1180.46
R438 VGND.n1647 VGND.n1646 1180.46
R439 VGND.n1413 VGND.n1412 1180.46
R440 VGND.n1415 VGND.n1414 1180.46
R441 VGND.n1480 VGND.n1479 1180.46
R442 VGND.n1482 VGND.n1481 1180.46
R443 VGND.n1506 VGND.n1505 1180.46
R444 VGND.n1508 VGND.n1507 1180.46
R445 VGND.n1532 VGND.n1531 1180.46
R446 VGND.n1534 VGND.n1533 1180.46
R447 VGND.n1569 VGND.n1568 1180.46
R448 VGND.n1586 VGND.n1585 1180.46
R449 VGND.n1584 VGND.n1583 1180.46
R450 VGND.n1579 VGND.n1578 1180.46
R451 VGND.n1574 VGND.n1573 1180.46
R452 VGND.n2887 VGND.n2886 1180.46
R453 VGND.n2889 VGND.n2888 1180.46
R454 VGND.n1342 VGND.n1341 1180.46
R455 VGND.n1426 VGND.n1425 1180.46
R456 VGND.n1431 VGND.n1430 1180.46
R457 VGND.n1436 VGND.n1435 1180.46
R458 VGND.n1441 VGND.n1440 1180.46
R459 VGND.n1446 VGND.n1445 1180.46
R460 VGND.n1451 VGND.n1450 1180.46
R461 VGND.n1456 VGND.n1455 1180.46
R462 VGND.n1463 VGND.n1462 1180.46
R463 VGND.n1461 VGND.n1460 1180.46
R464 VGND.n1598 VGND.n1597 1180.46
R465 VGND.n1603 VGND.n1602 1180.46
R466 VGND.n1618 VGND.n1617 1180.46
R467 VGND.n1616 VGND.n1615 1180.46
R468 VGND.n1611 VGND.n1610 1180.46
R469 VGND.n1034 VGND.n1033 1180.46
R470 VGND.n1039 VGND.n1038 1180.46
R471 VGND.n1099 VGND.n1098 1180.46
R472 VGND.n1097 VGND.n1096 1180.46
R473 VGND.n1092 VGND.n1091 1180.46
R474 VGND.n1087 VGND.n1086 1180.46
R475 VGND.n1082 VGND.n1081 1180.46
R476 VGND.n1077 VGND.n1076 1180.46
R477 VGND.n1072 VGND.n1071 1180.46
R478 VGND.n1050 VGND.n1041 1180.46
R479 VGND.n1055 VGND.n1054 1180.46
R480 VGND.n1060 VGND.n1059 1180.46
R481 VGND.n1062 VGND.n1061 1180.46
R482 VGND.n2907 VGND.n2906 1180.46
R483 VGND.n2909 VGND.n2908 1180.46
R484 VGND.t237 VGND.n3011 1180.08
R485 VGND.n1387 VGND.n1386 1169.57
R486 VGND.n3015 VGND.t57 1146.36
R487 VGND.n3017 VGND.t56 1112.64
R488 VGND.n3016 VGND.t1194 1112.64
R489 VGND.n2351 VGND.n2349 1070.21
R490 VGND.n2968 VGND 1055.35
R491 VGND.n2251 VGND.n2250 1052.29
R492 VGND.t484 VGND.n2181 1032.59
R493 VGND.t1270 VGND.n2641 988.926
R494 VGND.t1966 VGND.n2646 988.926
R495 VGND.t680 VGND.n2651 988.926
R496 VGND.t858 VGND.n2656 988.926
R497 VGND.t694 VGND.n2661 988.926
R498 VGND.t2048 VGND.n2666 988.926
R499 VGND.t668 VGND.n2671 988.926
R500 VGND.n2672 VGND.t421 988.926
R501 VGND.t1933 VGND.n2717 988.926
R502 VGND.n2718 VGND.t541 988.926
R503 VGND.t1100 VGND.n2750 988.926
R504 VGND.n2756 VGND.t1981 988.926
R505 VGND.n2755 VGND.t728 988.926
R506 VGND.t1598 VGND.n2790 988.926
R507 VGND.n2791 VGND.t1584 988.926
R508 VGND.n2345 VGND.t1498 988.926
R509 VGND.n2340 VGND.t1958 988.926
R510 VGND.n2335 VGND.t2495 988.926
R511 VGND.n2330 VGND.t534 988.926
R512 VGND.n2325 VGND.t1956 988.926
R513 VGND.n2320 VGND.t80 988.926
R514 VGND.n2315 VGND.t2123 988.926
R515 VGND.n2310 VGND.t798 988.926
R516 VGND.n2305 VGND.t780 988.926
R517 VGND.n2300 VGND.t585 988.926
R518 VGND.n2295 VGND.t2469 988.926
R519 VGND.n2290 VGND.t2414 988.926
R520 VGND.n2544 VGND.t2162 988.926
R521 VGND.n2543 VGND.t1260 988.926
R522 VGND.n2538 VGND.t324 988.926
R523 VGND.n2354 VGND.t2664 988.926
R524 VGND.t2654 VGND.n2379 988.926
R525 VGND.n2380 VGND.t1156 988.926
R526 VGND.t1737 VGND.n2405 988.926
R527 VGND.n2406 VGND.t700 988.926
R528 VGND.t1987 VGND.n2431 988.926
R529 VGND.n2432 VGND.t674 988.926
R530 VGND.t1121 VGND.n2457 988.926
R531 VGND.n2458 VGND.t708 988.926
R532 VGND.t784 VGND.n2483 988.926
R533 VGND.n2484 VGND.t2672 988.926
R534 VGND.t1974 VGND.n2514 988.926
R535 VGND.t734 VGND.n2519 988.926
R536 VGND.t2554 VGND.n2524 988.926
R537 VGND.n2525 VGND.t1591 988.926
R538 VGND.t1284 VGND.n2366 988.926
R539 VGND.n2367 VGND.t2109 988.926
R540 VGND.t1067 VGND.n2392 988.926
R541 VGND.n2393 VGND.t986 988.926
R542 VGND.t872 VGND.n2418 988.926
R543 VGND.n2419 VGND.t750 988.926
R544 VGND.t2243 VGND.n2444 988.926
R545 VGND.n2445 VGND.t1150 988.926
R546 VGND.t1112 VGND.n2470 988.926
R547 VGND.n2471 VGND.t527 988.926
R548 VGND.t1092 VGND.n2496 988.926
R549 VGND.n2502 VGND.t138 988.926
R550 VGND.n2501 VGND.t1502 988.926
R551 VGND.t13 VGND.n2812 988.926
R552 VGND.n2813 VGND.t1253 988.926
R553 VGND.t813 VGND.n1913 988.926
R554 VGND.n1914 VGND.t1185 988.926
R555 VGND.t2489 VGND.n1924 988.926
R556 VGND.n1925 VGND.t259 988.926
R557 VGND.t2069 VGND.n1935 988.926
R558 VGND.n1936 VGND.t76 988.926
R559 VGND.t592 VGND.n1946 988.926
R560 VGND.n1947 VGND.t792 988.926
R561 VGND.t157 VGND.n1957 988.926
R562 VGND.n1958 VGND.t580 988.926
R563 VGND.t2465 VGND.n1968 988.926
R564 VGND.n1969 VGND.t1970 988.926
R565 VGND.t2156 VGND.n1979 988.926
R566 VGND.t42 VGND.n1984 988.926
R567 VGND.n1985 VGND.t338 988.926
R568 VGND.t1268 VGND.n599 988.926
R569 VGND.n2059 VGND.t1964 988.926
R570 VGND.n2058 VGND.t61 988.926
R571 VGND.n2053 VGND.t856 988.926
R572 VGND.n2048 VGND.t692 988.926
R573 VGND.n2043 VGND.t2046 988.926
R574 VGND.n2038 VGND.t666 988.926
R575 VGND.n2033 VGND.t419 988.926
R576 VGND.n2028 VGND.t1931 988.926
R577 VGND.n2023 VGND.t538 988.926
R578 VGND.n2018 VGND.t1098 988.926
R579 VGND.n2013 VGND.t2419 988.926
R580 VGND.n2008 VGND.t726 988.926
R581 VGND.n2003 VGND.t2417 988.926
R582 VGND.n601 VGND.t1582 988.926
R583 VGND.t2666 VGND.n2072 988.926
R584 VGND.t2656 VGND.n2077 988.926
R585 VGND.t1154 VGND.n2082 988.926
R586 VGND.t1739 VGND.n2087 988.926
R587 VGND.t2210 VGND.n2092 988.926
R588 VGND.t1989 VGND.n2097 988.926
R589 VGND.t676 VGND.n2102 988.926
R590 VGND.t0 VGND.n2107 988.926
R591 VGND.t710 VGND.n2112 988.926
R592 VGND.t786 VGND.n2117 988.926
R593 VGND.t2674 VGND.n2122 988.926
R594 VGND.n2128 VGND.t1976 988.926
R595 VGND.n2127 VGND.t736 988.926
R596 VGND.t2556 VGND.n2837 988.926
R597 VGND.n2838 VGND.t332 988.926
R598 VGND.n2179 VGND.t1286 988.926
R599 VGND.t2091 VGND.n1754 988.926
R600 VGND.t1065 VGND.n1764 988.926
R601 VGND.n1765 VGND.t988 988.926
R602 VGND.t874 VGND.n1775 988.926
R603 VGND.n1776 VGND.t752 988.926
R604 VGND.t2245 VGND.n1786 988.926
R605 VGND.n1787 VGND.t1214 988.926
R606 VGND.t1114 VGND.n1797 988.926
R607 VGND.n1798 VGND.t529 988.926
R608 VGND.t1094 VGND.n1808 988.926
R609 VGND.n1809 VGND.t140 988.926
R610 VGND.t1504 VGND.n1819 988.926
R611 VGND.t33 VGND.n1824 988.926
R612 VGND.n1825 VGND.t1255 988.926
R613 VGND.t1279 VGND.n1681 988.926
R614 VGND.n1682 VGND.t2103 988.926
R615 VGND.t1071 VGND.n1692 988.926
R616 VGND.t982 VGND.n1697 988.926
R617 VGND.t169 VGND.n1702 988.926
R618 VGND.t2055 VGND.n1707 988.926
R619 VGND.t2239 VGND.n1712 988.926
R620 VGND.t1146 VGND.n1717 988.926
R621 VGND.t1227 VGND.n1722 988.926
R622 VGND.t525 VGND.n1727 988.926
R623 VGND.t1090 VGND.n1732 988.926
R624 VGND.n1849 VGND.t2425 988.926
R625 VGND.n1848 VGND.t1415 988.926
R626 VGND.n1843 VGND.t9 988.926
R627 VGND.n1734 VGND.t1251 988.926
R628 VGND.t811 VGND.n672 988.926
R629 VGND.t1183 VGND.n677 988.926
R630 VGND.t2491 VGND.n682 988.926
R631 VGND.t257 VGND.n687 988.926
R632 VGND.t2067 VGND.n692 988.926
R633 VGND.t74 VGND.n697 988.926
R634 VGND.t590 VGND.n702 988.926
R635 VGND.t3 VGND.n707 988.926
R636 VGND.t155 VGND.n712 988.926
R637 VGND.t790 VGND.n717 988.926
R638 VGND.t2463 VGND.n722 988.926
R639 VGND.n728 VGND.t1968 988.926
R640 VGND.n727 VGND.t2154 988.926
R641 VGND.t40 VGND.n2862 988.926
R642 VGND.n2863 VGND.t336 988.926
R643 VGND.n1355 VGND.t2166 988.926
R644 VGND.n877 VGND.t250 988.926
R645 VGND.n872 VGND.t1058 988.926
R646 VGND.t2228 VGND.n821 988.926
R647 VGND.t2086 VGND.n826 988.926
R648 VGND.t2252 VGND.n831 988.926
R649 VGND.t2513 VGND.n836 988.926
R650 VGND.t773 VGND.n841 988.926
R651 VGND.t2096 VGND.n846 988.926
R652 VGND.t505 VGND.n851 988.926
R653 VGND.n857 VGND.t344 988.926
R654 VGND.n856 VGND.t1337 988.926
R655 VGND.n1665 VGND.t2118 988.926
R656 VGND.n1664 VGND.t5 988.926
R657 VGND.n1659 VGND.t1243 988.926
R658 VGND.t2662 VGND.n1393 988.926
R659 VGND.t2652 VGND.n1398 988.926
R660 VGND.n1399 VGND.t1158 988.926
R661 VGND.t863 VGND.n1493 988.926
R662 VGND.n1494 VGND.t698 988.926
R663 VGND.t1985 VGND.n1519 988.926
R664 VGND.n1520 VGND.t672 988.926
R665 VGND.t1119 VGND.n1545 988.926
R666 VGND.t706 VGND.n1550 988.926
R667 VGND.n1556 VGND.t545 988.926
R668 VGND.n1555 VGND.t2670 988.926
R669 VGND.t1972 VGND.n1635 988.926
R670 VGND.t732 VGND.n1640 988.926
R671 VGND.t2552 VGND.n1645 988.926
R672 VGND.n1646 VGND.t1589 988.926
R673 VGND.t2164 VGND.n1413 988.926
R674 VGND.n1414 VGND.t704 988.926
R675 VGND.t1060 VGND.n1480 988.926
R676 VGND.n1481 VGND.t2226 988.926
R677 VGND.t245 VGND.n1506 988.926
R678 VGND.n1507 VGND.t2250 988.926
R679 VGND.t2511 VGND.n1532 988.926
R680 VGND.n1533 VGND.t771 988.926
R681 VGND.t2094 VGND.n1569 988.926
R682 VGND.n1585 VGND.t503 988.926
R683 VGND.n1584 VGND.t721 988.926
R684 VGND.n1579 VGND.t1335 988.926
R685 VGND.n1574 VGND.t2116 988.926
R686 VGND.t17 VGND.n2887 988.926
R687 VGND.n2888 VGND.t295 988.926
R688 VGND.n1341 VGND.t1496 988.926
R689 VGND.t1189 VGND.n1426 988.926
R690 VGND.t713 VGND.n1431 988.926
R691 VGND.t263 VGND.n1436 988.926
R692 VGND.t1954 VGND.n1441 988.926
R693 VGND.t78 VGND.n1446 988.926
R694 VGND.t2121 VGND.n1451 988.926
R695 VGND.t796 VGND.n1456 988.926
R696 VGND.n1462 VGND.t778 988.926
R697 VGND.n1461 VGND.t582 988.926
R698 VGND.t2467 VGND.n1598 988.926
R699 VGND.t2411 VGND.n1603 988.926
R700 VGND.n1617 VGND.t2160 988.926
R701 VGND.n1616 VGND.t1257 988.926
R702 VGND.n1611 VGND.t321 988.926
R703 VGND.t1281 VGND.n1034 988.926
R704 VGND.t2105 VGND.n1039 988.926
R705 VGND.n1098 VGND.t1069 988.926
R706 VGND.n1097 VGND.t984 988.926
R707 VGND.n1092 VGND.t171 988.926
R708 VGND.n1087 VGND.t2053 988.926
R709 VGND.n1082 VGND.t2237 988.926
R710 VGND.n1077 VGND.t1144 988.926
R711 VGND.n1072 VGND.t1225 988.926
R712 VGND.t523 VGND.n1050 988.926
R713 VGND.t1088 VGND.n1055 988.926
R714 VGND.t2423 VGND.n1060 988.926
R715 VGND.n1061 VGND.t1413 988.926
R716 VGND.t11 VGND.n2907 988.926
R717 VGND.n2908 VGND.t1249 988.926
R718 VGND.n1335 VGND.t2607 988.926
R719 VGND.t2336 VGND.n929 988.926
R720 VGND.t2314 VGND.n934 988.926
R721 VGND.t2602 VGND.n939 988.926
R722 VGND.t2591 VGND.n944 988.926
R723 VGND.t2572 VGND.n949 988.926
R724 VGND.t1675 VGND.n954 988.926
R725 VGND.t1654 VGND.n959 988.926
R726 VGND.t2568 VGND.n964 988.926
R727 VGND.t2302 VGND.n969 988.926
R728 VGND.t2289 VGND.n974 988.926
R729 VGND.t2626 VGND.n979 988.926
R730 VGND.t2362 VGND.n984 988.926
R731 VGND.t1704 VGND.n989 988.926
R732 VGND.n990 VGND.t2635 988.926
R733 VGND.n2248 VGND.n539 934.784
R734 VGND.n116 VGND 927.203
R735 VGND.n134 VGND 927.203
R736 VGND.n2182 VGND 918.774
R737 VGND.n194 VGND 910.346
R738 VGND.n165 VGND 910.346
R739 VGND.t1556 VGND.n2967 909.365
R740 VGND.n2285 VGND.n473 900
R741 VGND.n2641 VGND.t1208 852.769
R742 VGND.n2646 VGND.t52 852.769
R743 VGND.n2651 VGND.t1167 852.769
R744 VGND.n2656 VGND.t619 852.769
R745 VGND.n2661 VGND.t1172 852.769
R746 VGND.n2666 VGND.t2220 852.769
R747 VGND.n2671 VGND.t1492 852.769
R748 VGND.n2672 VGND.t495 852.769
R749 VGND.n2717 VGND.t1241 852.769
R750 VGND.n2718 VGND.t720 852.769
R751 VGND.n2750 VGND.t55 852.769
R752 VGND.n2756 VGND.t2660 852.769
R753 VGND.t560 VGND.n2755 852.769
R754 VGND.n2790 VGND.t204 852.769
R755 VGND.n2791 VGND.t1109 852.769
R756 VGND.n2935 VGND.t747 852.769
R757 VGND.t2482 VGND.n2345 852.769
R758 VGND.t176 VGND.n2340 852.769
R759 VGND.t1211 VGND.n2335 852.769
R760 VGND.t2099 VGND.n2330 852.769
R761 VGND.t1266 VGND.n2325 852.769
R762 VGND.t2506 VGND.n2320 852.769
R763 VGND.t470 VGND.n2315 852.769
R764 VGND.t1995 VGND.n2310 852.769
R765 VGND.t661 VGND.n2305 852.769
R766 VGND.t1388 VGND.n2300 852.769
R767 VGND.t618 VGND.n2295 852.769
R768 VGND.t2077 VGND.n2290 852.769
R769 VGND.n2544 VGND.t2093 852.769
R770 VGND.t924 VGND.n2543 852.769
R771 VGND.t1518 VGND.n2538 852.769
R772 VGND.t2225 VGND.n208 852.769
R773 VGND.n2354 VGND.t1389 852.769
R774 VGND.n2379 VGND.t561 852.769
R775 VGND.n2380 VGND.t127 852.769
R776 VGND.n2405 VGND.t1125 852.769
R777 VGND.n2406 VGND.t1942 852.769
R778 VGND.n2431 VGND.t2480 852.769
R779 VGND.n2432 VGND.t1291 852.769
R780 VGND.n2457 VGND.t2484 852.769
R781 VGND.n2458 VGND.t1909 852.769
R782 VGND.n2483 VGND.t1596 852.769
R783 VGND.n2484 VGND.t723 852.769
R784 VGND.n2514 VGND.t766 852.769
R785 VGND.n2519 VGND.t44 852.769
R786 VGND.n2524 VGND.t164 852.769
R787 VGND.n2525 VGND.t852 852.769
R788 VGND.t2438 VGND.n209 852.769
R789 VGND.n2366 VGND.t558 852.769
R790 VGND.n2367 VGND.t255 852.769
R791 VGND.n2392 VGND.t2648 852.769
R792 VGND.n2393 VGND.t879 852.769
R793 VGND.n2418 VGND.t1242 852.769
R794 VGND.n2419 VGND.t1126 852.769
R795 VGND.n2444 VGND.t940 852.769
R796 VGND.n2445 VGND.t162 852.769
R797 VGND.n2470 VGND.t2111 852.769
R798 VGND.n2471 VGND.t559 852.769
R799 VGND.n2496 VGND.t1213 852.769
R800 VGND.n2502 VGND.t1104 852.769
R801 VGND.t1274 VGND.n2501 852.769
R802 VGND.n2812 VGND.t1097 852.769
R803 VGND.n2813 VGND.t45 852.769
R804 VGND.t50 VGND.n210 852.769
R805 VGND.n1913 VGND.t1568 852.769
R806 VGND.n1914 VGND.t206 852.769
R807 VGND.n1924 VGND.t1941 852.769
R808 VGND.n1925 VGND.t1193 852.769
R809 VGND.n1935 VGND.t1940 852.769
R810 VGND.n1936 VGND.t2471 852.769
R811 VGND.n1946 VGND.t646 852.769
R812 VGND.n1947 VGND.t882 852.769
R813 VGND.n1957 VGND.t877 852.769
R814 VGND.n1958 VGND.t925 852.769
R815 VGND.n1968 VGND.t782 852.769
R816 VGND.n1969 VGND.t1076 852.769
R817 VGND.n1979 VGND.t1192 852.769
R818 VGND.n1984 VGND.t2223 852.769
R819 VGND.n1985 VGND.t2479 852.769
R820 VGND.t69 VGND.n211 852.769
R821 VGND.n599 VGND.t2222 852.769
R822 VGND.n2059 VGND.t881 852.769
R823 VGND.t236 VGND.n2058 852.769
R824 VGND.t498 VGND.n2053 852.769
R825 VGND.t783 VGND.n2048 852.769
R826 VGND.t1387 VGND.n2043 852.769
R827 VGND.t1579 VGND.n2038 852.769
R828 VGND.t268 VGND.n2033 852.769
R829 VGND.t1210 VGND.n2028 852.769
R830 VGND.t222 VGND.n2023 852.769
R831 VGND.t202 VGND.n2018 852.769
R832 VGND.t943 VGND.n2013 852.769
R833 VGND.t2483 VGND.n2008 852.769
R834 VGND.t765 VGND.n2003 852.769
R835 VGND.n601 VGND.t1565 852.769
R836 VGND.t880 VGND.n212 852.769
R837 VGND.n2072 VGND.t2221 852.769
R838 VGND.n2077 VGND.t1173 852.769
R839 VGND.n2082 VGND.t1199 852.769
R840 VGND.n2087 VGND.t154 852.769
R841 VGND.n2092 VGND.t1262 852.769
R842 VGND.n2097 VGND.t2649 852.769
R843 VGND.n2102 VGND.t496 852.769
R844 VGND.n2107 VGND.t878 852.769
R845 VGND.n2112 VGND.t647 852.769
R846 VGND.n2117 VGND.t2089 852.769
R847 VGND.n2122 VGND.t2387 852.769
R848 VGND.n2128 VGND.t1491 852.769
R849 VGND.t266 VGND.n2127 852.769
R850 VGND.n2837 VGND.t645 852.769
R851 VGND.n2838 VGND.t219 852.769
R852 VGND.t203 VGND.n213 852.769
R853 VGND.t372 VGND.n2179 852.769
R854 VGND.n1754 VGND.t1519 852.769
R855 VGND.n1764 VGND.t397 852.769
R856 VGND.n1765 VGND.t49 852.769
R857 VGND.n1775 VGND.t1489 852.769
R858 VGND.n1776 VGND.t589 852.769
R859 VGND.n1786 VGND.t1178 852.769
R860 VGND.n1787 VGND.t2076 852.769
R861 VGND.n1797 VGND.t1994 852.769
R862 VGND.n1798 VGND.t1123 852.769
R863 VGND.n1808 VGND.t2505 852.769
R864 VGND.n1809 VGND.t1129 852.769
R865 VGND.n1819 VGND.t205 852.769
R866 VGND.n1824 VGND.t1106 852.769
R867 VGND.n1825 VGND.t1128 852.769
R868 VGND.t20 VGND.n214 852.769
R869 VGND.n1681 VGND.t163 852.769
R870 VGND.n1682 VGND.t1216 852.769
R871 VGND.n1692 VGND.t2088 852.769
R872 VGND.n1697 VGND.t1197 852.769
R873 VGND.n1702 VGND.t939 852.769
R874 VGND.n1707 VGND.t1915 852.769
R875 VGND.n1712 VGND.t1487 852.769
R876 VGND.n1717 VGND.t2078 852.769
R877 VGND.n1722 VGND.t1276 852.769
R878 VGND.n1727 VGND.t499 852.769
R879 VGND.n1732 VGND.t2224 852.769
R880 VGND.n1849 VGND.t691 852.769
R881 VGND.t2478 VGND.n1848 852.769
R882 VGND.t1482 VGND.n1843 852.769
R883 VGND.n1734 VGND.t46 852.769
R884 VGND.t1074 VGND.n215 852.769
R885 VGND.n672 VGND.t2085 852.769
R886 VGND.n677 VGND.t941 852.769
R887 VGND.n682 VGND.t165 852.769
R888 VGND.n687 VGND.t1521 852.769
R889 VGND.n692 VGND.t1708 852.769
R890 VGND.n697 VGND.t866 852.769
R891 VGND.n702 VGND.t1166 852.769
R892 VGND.n707 VGND.t1180 852.769
R893 VGND.n712 VGND.t240 852.769
R894 VGND.n717 VGND.t1277 852.769
R895 VGND.n722 VGND.t2388 852.769
R896 VGND.n728 VGND.t373 852.769
R897 VGND.t1116 VGND.n727 852.769
R898 VGND.n2862 VGND.t1917 852.769
R899 VGND.n2863 VGND.t2481 852.769
R900 VGND.t719 VGND.n216 852.769
R901 VGND.t1288 VGND.n1355 852.769
R902 VGND.t467 VGND.n877 852.769
R903 VGND.t2268 VGND.n872 852.769
R904 VGND.n821 VGND.t267 852.769
R905 VGND.n826 VGND.t2372 852.769
R906 VGND.n831 VGND.t1483 852.769
R907 VGND.n836 VGND.t853 852.769
R908 VGND.n841 VGND.t1294 852.769
R909 VGND.n846 VGND.t2504 852.769
R910 VGND.n851 VGND.t220 852.769
R911 VGND.n857 VGND.t1289 852.769
R912 VGND.t662 VGND.n856 852.769
R913 VGND.n1665 VGND.t2232 852.769
R914 VGND.t938 VGND.n1664 852.769
R915 VGND.t1103 VGND.n1659 852.769
R916 VGND.t221 VGND.n217 852.769
R917 VGND.n1393 VGND.t371 852.769
R918 VGND.n1398 VGND.t663 852.769
R919 VGND.n1399 VGND.t1127 852.769
R920 VGND.n1493 VGND.t1105 852.769
R921 VGND.n1494 VGND.t1212 852.769
R922 VGND.n1519 VGND.t1939 852.769
R923 VGND.n1520 VGND.t2485 852.769
R924 VGND.n1545 VGND.t2168 852.769
R925 VGND.n1550 VGND.t2080 852.769
R926 VGND.n1556 VGND.t1711 852.769
R927 VGND.t2102 VGND.n1555 852.769
R928 VGND.n1635 VGND.t1075 852.769
R929 VGND.n1640 VGND.t174 852.769
R930 VGND.n1645 VGND.t2098 852.769
R931 VGND.n1646 VGND.t770 852.769
R932 VGND.t414 VGND.n218 852.769
R933 VGND.n1413 VGND.t644 852.769
R934 VGND.n1414 VGND.t1603 852.769
R935 VGND.n1480 VGND.t1223 852.769
R936 VGND.n1481 VGND.t53 852.769
R937 VGND.n1506 VGND.t2502 852.769
R938 VGND.n1507 VGND.t2386 852.769
R939 VGND.n1532 VGND.t2385 852.769
R940 VGND.n1533 VGND.t1124 852.769
R941 VGND.n1569 VGND.t249 852.769
R942 VGND.n1585 VGND.t1500 852.769
R943 VGND.t235 VGND.n1584 852.769
R944 VGND.t160 VGND.n1579 852.769
R945 VGND.t1296 VGND.n1574 852.769
R946 VGND.n2887 VGND.t748 852.769
R947 VGND.n2888 VGND.t1130 852.769
R948 VGND.t2437 VGND.n219 852.769
R949 VGND.n1341 VGND.t876 852.769
R950 VGND.n1426 VGND.t1493 852.769
R951 VGND.n1431 VGND.t2503 852.769
R952 VGND.n1436 VGND.t1938 852.769
R953 VGND.n1441 VGND.t54 852.769
R954 VGND.n1446 VGND.t761 852.769
R955 VGND.n1451 VGND.t175 852.769
R956 VGND.n1456 VGND.t2370 852.769
R957 VGND.n1462 VGND.t71 852.769
R958 VGND.t1916 VGND.n1461 852.769
R959 VGND.n1598 VGND.t1486 852.769
R960 VGND.n1603 VGND.t2488 852.769
R961 VGND.n1617 VGND.t19 852.769
R962 VGND.t1578 VGND.n1616 852.769
R963 VGND.t70 VGND.n1611 852.769
R964 VGND.t1073 VGND.n220 852.769
R965 VGND.n1034 VGND.t1179 852.769
R966 VGND.n1039 VGND.t1141 852.769
R967 VGND.n1098 VGND.t32 852.769
R968 VGND.t21 VGND.n1097 852.769
R969 VGND.t2661 VGND.n1092 852.769
R970 VGND.t48 VGND.n1087 852.769
R971 VGND.t2486 VGND.n1082 852.769
R972 VGND.t159 VGND.n1077 852.769
R973 VGND.t2090 VGND.n1072 852.769
R974 VGND.n1050 VGND.t1485 852.769
R975 VGND.n1055 VGND.t1602 852.769
R976 VGND.n1060 VGND.t1182 852.769
R977 VGND.n1061 VGND.t1198 852.769
R978 VGND.n2907 VGND.t47 852.769
R979 VGND.n2908 VGND.t1131 852.769
R980 VGND.t923 VGND.n221 852.769
R981 VGND.t370 VGND.n1335 852.769
R982 VGND.n929 VGND.t1520 852.769
R983 VGND.n934 VGND.t1293 852.769
R984 VGND.n939 VGND.t746 852.769
R985 VGND.n944 VGND.t865 852.769
R986 VGND.n949 VGND.t1914 852.769
R987 VGND.n954 VGND.t126 852.769
R988 VGND.n959 VGND.t2436 852.769
R989 VGND.n964 VGND.t1937 852.769
R990 VGND.n969 VGND.t1390 852.769
R991 VGND.n974 VGND.t1218 852.769
R992 VGND.n979 VGND.t1152 852.769
R993 VGND.n984 VGND.t1290 852.769
R994 VGND.n989 VGND.t161 852.769
R995 VGND.n990 VGND.t1209 852.769
R996 VGND.n2918 VGND.t1490 852.769
R997 VGND.n2249 VGND 851.341
R998 VGND.n2944 VGND.n2943 846.154
R999 VGND.n2350 VGND.t1809 809.773
R1000 VGND.n2352 VGND.t1884 809.773
R1001 VGND.t1791 VGND.n2353 809.773
R1002 VGND.n473 VGND.t1833 809.773
R1003 VGND.t1905 VGND.n503 809.773
R1004 VGND.t1785 VGND.n504 809.773
R1005 VGND.n2180 VGND.t1827 809.773
R1006 VGND.t1839 VGND.n539 809.773
R1007 VGND.n1387 VGND.t1863 809.773
R1008 VGND.t1794 VGND.n1388 809.773
R1009 VGND.n1339 VGND.t1866 809.773
R1010 VGND.t1896 VGND.n1340 809.773
R1011 VGND.n1338 VGND.t1836 809.773
R1012 VGND.n1336 VGND.t1690 809.773
R1013 VGND.t401 VGND.t356 708.047
R1014 VGND.t356 VGND.t358 708.047
R1015 VGND.t358 VGND.t442 708.047
R1016 VGND.t442 VGND.t1397 708.047
R1017 VGND.t1397 VGND.t1394 708.047
R1018 VGND.t1394 VGND.t1400 708.047
R1019 VGND.t1400 VGND.t1391 708.047
R1020 VGND.t1923 VGND.t56 708.047
R1021 VGND.t378 VGND.t410 708.047
R1022 VGND.t410 VGND.t383 708.047
R1023 VGND.t383 VGND.t360 708.047
R1024 VGND.t360 VGND.t1393 708.047
R1025 VGND.t1393 VGND.t1399 708.047
R1026 VGND.t1399 VGND.t1396 708.047
R1027 VGND.t1396 VGND.t1402 708.047
R1028 VGND.t451 VGND.t436 708.047
R1029 VGND.t436 VGND.t404 708.047
R1030 VGND.t404 VGND.t380 708.047
R1031 VGND.t380 VGND.t217 708.047
R1032 VGND.t217 VGND.t213 708.047
R1033 VGND.t213 VGND.t207 708.047
R1034 VGND.t207 VGND.t209 708.047
R1035 VGND.t1920 VGND.t57 708.047
R1036 VGND.t391 VGND.t458 708.047
R1037 VGND.t458 VGND.t374 708.047
R1038 VGND.t374 VGND.t342 708.047
R1039 VGND.t342 VGND.t658 708.047
R1040 VGND.t658 VGND.t655 708.047
R1041 VGND.t655 VGND.t649 708.047
R1042 VGND.t649 VGND.t652 708.047
R1043 VGND.t408 VGND.t387 708.047
R1044 VGND.t387 VGND.t385 708.047
R1045 VGND.t385 VGND.t376 708.047
R1046 VGND.t376 VGND.t654 708.047
R1047 VGND.t654 VGND.t648 708.047
R1048 VGND.t648 VGND.t657 708.047
R1049 VGND.t657 VGND.t651 708.047
R1050 VGND.t350 VGND.t398 708.047
R1051 VGND.t455 VGND.t350 708.047
R1052 VGND.t406 VGND.t455 708.047
R1053 VGND.t215 VGND.t406 708.047
R1054 VGND.t211 VGND.t215 708.047
R1055 VGND.t216 VGND.t211 708.047
R1056 VGND.t212 VGND.t216 708.047
R1057 VGND.n2971 VGND.n2970 708.047
R1058 VGND.t326 VGND.t1195 691.188
R1059 VGND.t2081 VGND.t2498 691.188
R1060 VGND.t2454 VGND.t412 657.471
R1061 VGND.t389 VGND.t1557 657.471
R1062 VGND.t453 VGND.t1553 657.471
R1063 VGND.t475 VGND.t1547 657.471
R1064 VGND.t1452 VGND.t1302 657.471
R1065 VGND.t2259 VGND.t1300 657.471
R1066 VGND.t596 VGND.t1298 657.471
R1067 VGND.t491 VGND.t1434 657.471
R1068 VGND.t412 VGND.t462 654.197
R1069 VGND.t1434 VGND.t1436 654.197
R1070 VGND VGND.n194 640.614
R1071 VGND VGND.n134 640.614
R1072 VGND VGND.n165 640.614
R1073 VGND.n2182 VGND 640.614
R1074 VGND.n116 VGND 632.184
R1075 VGND.t944 VGND.t1594 630.62
R1076 VGND.t253 VGND.t2518 630.62
R1077 VGND.t59 VGND.t952 630.62
R1078 VGND.t855 VGND.t950 630.62
R1079 VGND.t167 VGND.t2526 630.62
R1080 VGND.t2428 VGND.t2534 630.62
R1081 VGND.t2516 VGND.t2532 630.62
R1082 VGND.t1142 VGND.t2524 630.62
R1083 VGND.t2522 VGND.t1108 630.62
R1084 VGND.t508 VGND.t2536 630.62
R1085 VGND.t948 VGND.t2450 630.62
R1086 VGND.t2422 VGND.t946 630.62
R1087 VGND.t2530 VGND.t1411 630.62
R1088 VGND.t2528 VGND.t8 630.62
R1089 VGND.t1581 VGND.t954 630.62
R1090 VGND.t2520 VGND.t2623 630.62
R1091 VGND.t2682 VGND.t1273 630.62
R1092 VGND.t2063 VGND.t2651 630.62
R1093 VGND.t610 VGND.t1153 630.62
R1094 VGND.t1408 VGND.t262 630.62
R1095 VGND.t2680 VGND.t697 630.62
R1096 VGND.t2059 VGND.t2052 630.62
R1097 VGND.t2057 VGND.t671 630.62
R1098 VGND.t2678 VGND.t1118 630.62
R1099 VGND.t2676 VGND.t1936 630.62
R1100 VGND.t2061 VGND.t788 630.62
R1101 VGND.t1420 VGND.t349 630.62
R1102 VGND.t1418 VGND.t1978 630.62
R1103 VGND.t616 VGND.t731 630.62
R1104 VGND.t614 VGND.t2558 630.62
R1105 VGND.t612 VGND.t341 630.62
R1106 VGND.t2065 VGND.t2283 630.62
R1107 VGND.t1278 VGND.t2141 630.62
R1108 VGND.t1426 VGND.t2107 630.62
R1109 VGND.t1063 VGND.t2149 630.62
R1110 VGND.t2147 VGND.t861 630.62
R1111 VGND.t173 VGND.t2139 630.62
R1112 VGND.t1422 VGND.t2430 630.62
R1113 VGND.t2241 VGND.t2686 630.62
R1114 VGND.t2137 VGND.t1148 630.62
R1115 VGND.t1110 VGND.t1430 630.62
R1116 VGND.t1424 VGND.t532 630.62
R1117 VGND.t2452 VGND.t2145 630.62
R1118 VGND.t2143 VGND.t143 630.62
R1119 VGND.t1417 VGND.t2684 630.62
R1120 VGND.t36 VGND.t1443 630.62
R1121 VGND.t1587 VGND.t2151 630.62
R1122 VGND.t1428 VGND.t2644 630.62
R1123 VGND.t2443 VGND.t2235 630.62
R1124 VGND.t702 VGND.t233 630.62
R1125 VGND.t606 VGND.t715 630.62
R1126 VGND.t980 VGND.t604 630.62
R1127 VGND.t2441 VGND.t243 630.62
R1128 VGND.t1993 VGND.t229 630.62
R1129 VGND.t227 VGND.t2509 630.62
R1130 VGND.t82 VGND.t2439 630.62
R1131 VGND.t2135 VGND.t1221 630.62
R1132 VGND.t501 VGND.t231 630.62
R1133 VGND.t2447 VGND.t1951 630.62
R1134 VGND.t1333 VGND.t2445 630.62
R1135 VGND.t225 VGND.t2114 630.62
R1136 VGND.t223 VGND.t15 630.62
R1137 VGND.t1247 VGND.t608 630.62
R1138 VGND.t2133 VGND.t2578 630.62
R1139 VGND.t1267 VGND.t124 630.62
R1140 VGND.t1963 VGND.t936 630.62
R1141 VGND.t2474 VGND.t679 630.62
R1142 VGND.t256 VGND.t88 630.62
R1143 VGND.t122 VGND.t563 630.62
R1144 VGND.t1056 VGND.t932 630.62
R1145 VGND.t930 VGND.t665 630.62
R1146 VGND.t418 VGND.t120 630.62
R1147 VGND.t118 VGND.t1930 630.62
R1148 VGND.t543 VGND.t934 630.62
R1149 VGND.t86 VGND.t347 630.62
R1150 VGND.t1983 VGND.t84 630.62
R1151 VGND.t928 VGND.t725 630.62
R1152 VGND.t1600 VGND.t926 630.62
R1153 VGND.t335 VGND.t2476 630.62
R1154 VGND.t116 VGND.t1688 630.62
R1155 VGND.t1593 VGND.t2383 630.62
R1156 VGND.t252 VGND.t2373 630.62
R1157 VGND.t1235 VGND.t1062 630.62
R1158 VGND.t1233 VGND.t854 630.62
R1159 VGND.t2381 VGND.t166 630.62
R1160 VGND.t1573 VGND.t2427 630.62
R1161 VGND.t1571 VGND.t2515 630.62
R1162 VGND.t2379 VGND.t775 630.62
R1163 VGND.t2377 VGND.t1107 630.62
R1164 VGND.t1575 VGND.t507 630.62
R1165 VGND.t1231 VGND.t2449 630.62
R1166 VGND.t1229 VGND.t2421 630.62
R1167 VGND.t1569 VGND.t1410 630.62
R1168 VGND.t1239 VGND.t7 630.62
R1169 VGND.t1580 VGND.t1237 630.62
R1170 VGND.t2375 VGND.t2621 630.62
R1171 VGND.t1283 VGND.t515 630.62
R1172 VGND.t2108 VGND.t576 630.62
R1173 VGND.t60 VGND.t478 630.62
R1174 VGND.t862 VGND.t521 630.62
R1175 VGND.t871 VGND.t513 630.62
R1176 VGND.t2431 VGND.t572 630.62
R1177 VGND.t2242 VGND.t570 630.62
R1178 VGND.t1149 VGND.t511 630.62
R1179 VGND.t1111 VGND.t509 630.62
R1180 VGND.t533 VGND.t574 630.62
R1181 VGND.t2453 VGND.t519 630.62
R1182 VGND.t144 VGND.t517 630.62
R1183 VGND.t568 VGND.t1501 630.62
R1184 VGND.t482 VGND.t37 630.62
R1185 VGND.t1588 VGND.t480 630.62
R1186 VGND.t578 VGND.t2647 630.62
R1187 VGND.t755 VGND.t2236 630.62
R1188 VGND.t703 VGND.t468 630.62
R1189 VGND.t718 VGND.t1202 630.62
R1190 VGND.t981 VGND.t1200 630.62
R1191 VGND.t152 VGND.t244 630.62
R1192 VGND.t73 VGND.t687 630.62
R1193 VGND.t685 VGND.t2510 630.62
R1194 VGND.t83 VGND.t150 630.62
R1195 VGND.t148 VGND.t1222 630.62
R1196 VGND.t502 VGND.t689 630.62
R1197 VGND.t759 VGND.t1952 630.62
R1198 VGND.t1334 VGND.t757 630.62
R1199 VGND.t683 VGND.t2115 630.62
R1200 VGND.t16 VGND.t1206 630.62
R1201 VGND.t1248 VGND.t1204 630.62
R1202 VGND.t146 VGND.t2580 630.62
R1203 VGND.t2233 VGND.t742 630.62
R1204 VGND.t1961 VGND.t315 630.62
R1205 VGND.t2206 VGND.t717 630.62
R1206 VGND.t2231 VGND.t2204 630.62
R1207 VGND.t241 VGND.t740 630.62
R1208 VGND.t1991 VGND.t311 630.62
R1209 VGND.t2508 VGND.t1053 630.62
R1210 VGND.t248 VGND.t738 630.62
R1211 VGND.t1220 VGND.t2044 630.62
R1212 VGND.t500 VGND.t313 630.62
R1213 VGND.t1950 VGND.t2202 630.62
R1214 VGND.t1908 VGND.t744 630.62
R1215 VGND.t1051 VGND.t2113 630.62
R1216 VGND.t1049 VGND.t1265 630.62
R1217 VGND.t1245 VGND.t2208 630.62
R1218 VGND.t317 VGND.t2571 630.62
R1219 VGND.t1275 VGND.t2181 630.62
R1220 VGND.t1962 VGND.t2171 630.62
R1221 VGND.t682 VGND.t2131 630.62
R1222 VGND.t1741 VGND.t2129 630.62
R1223 VGND.t562 VGND.t2179 630.62
R1224 VGND.t1055 VGND.t30 630.62
R1225 VGND.t2247 VGND.t28 630.62
R1226 VGND.t417 VGND.t2177 630.62
R1227 VGND.t2659 VGND.t2175 630.62
R1228 VGND.t540 VGND.t2169 630.62
R1229 VGND.t346 VGND.t2127 630.62
R1230 VGND.t1980 VGND.t2125 630.62
R1231 VGND.t26 VGND.t724 630.62
R1232 VGND.t24 VGND.t1597 630.62
R1233 VGND.t334 VGND.t22 630.62
R1234 VGND.t2173 VGND.t1683 630.62
R1235 VGND.t299 VGND.t1495 630.62
R1236 VGND.t2193 VGND.t1188 630.62
R1237 VGND.t307 VGND.t2494 630.62
R1238 VGND.t537 VGND.t305 630.62
R1239 VGND.t1953 VGND.t297 630.62
R1240 VGND.t2051 VGND.t2189 630.62
R1241 VGND.t2120 VGND.t2187 630.62
R1242 VGND.t795 VGND.t2199 630.62
R1243 VGND.t777 VGND.t2197 630.62
R1244 VGND.t587 VGND.t2191 630.62
R1245 VGND.t2669 VGND.t303 630.62
R1246 VGND.t301 VGND.t2416 630.62
R1247 VGND.t2185 VGND.t2159 630.62
R1248 VGND.t2183 VGND.t1263 630.62
R1249 VGND.t309 VGND.t294 630.62
R1250 VGND.t2195 VGND.t2341 630.62
R1251 VGND.t1595 VGND.t423 630.62
R1252 VGND.t254 VGND.t913 630.62
R1253 VGND.t1064 VGND.t431 630.62
R1254 VGND.t429 VGND.t860 630.62
R1255 VGND.t168 VGND.t921 630.62
R1256 VGND.t909 VGND.t2429 630.62
R1257 VGND.t2517 VGND.t2434 630.62
R1258 VGND.t919 VGND.t1143 630.62
R1259 VGND.t1224 VGND.t917 630.62
R1260 VGND.t531 VGND.t911 630.62
R1261 VGND.t427 VGND.t2451 630.62
R1262 VGND.t425 VGND.t142 630.62
R1263 VGND.t1412 VGND.t2432 630.62
R1264 VGND.t35 VGND.t415 630.62
R1265 VGND.t1586 VGND.t433 630.62
R1266 VGND.t915 VGND.t2641 630.62
R1267 VGND.t2500 VGND.t1494 630.62
R1268 VGND.t1187 VGND.t2548 630.62
R1269 VGND.t807 VGND.t2497 630.62
R1270 VGND.t536 VGND.t805 630.62
R1271 VGND.t1563 VGND.t2071 630.62
R1272 VGND.t2050 VGND.t2544 630.62
R1273 VGND.t2542 VGND.t594 630.62
R1274 VGND.t794 VGND.t1561 630.62
R1275 VGND.t1559 VGND.t776 630.62
R1276 VGND.t584 VGND.t2546 630.62
R1277 VGND.t803 VGND.t1102 630.62
R1278 VGND.t801 VGND.t2413 630.62
R1279 VGND.t2540 VGND.t2158 630.62
R1280 VGND.t2538 VGND.t1259 630.62
R1281 VGND.t293 VGND.t809 630.62
R1282 VGND.t2550 VGND.t2338 630.62
R1283 VGND.t1272 VGND.t849 630.62
R1284 VGND.t839 VGND.t2650 630.62
R1285 VGND.t1160 VGND.t1566 630.62
R1286 VGND.t261 VGND.t2273 630.62
R1287 VGND.t696 VGND.t847 630.62
R1288 VGND.t1057 VGND.t1514 630.62
R1289 VGND.t670 VGND.t1512 630.62
R1290 VGND.t1117 VGND.t845 630.62
R1291 VGND.t1935 VGND.t843 630.62
R1292 VGND.t1516 VGND.t544 630.62
R1293 VGND.t2271 VGND.t348 630.62
R1294 VGND.t1984 VGND.t2269 630.62
R1295 VGND.t730 VGND.t1510 630.62
R1296 VGND.t1508 VGND.t1601 630.62
R1297 VGND.t1506 VGND.t340 630.62
R1298 VGND.t841 VGND.t1703 630.62
R1299 VGND.t2234 VGND.t134 630.62
R1300 VGND.t1960 VGND.t1945 630.62
R1301 VGND.t716 VGND.t448 630.62
R1302 VGND.t446 VGND.t2230 630.62
R1303 VGND.t132 VGND.t242 630.62
R1304 VGND.t1086 VGND.t1992 630.62
R1305 VGND.t1084 VGND.t2507 630.62
R1306 VGND.t130 VGND.t247 630.62
R1307 VGND.t128 VGND.t1219 630.62
R1308 VGND.t588 VGND.t1943 630.62
R1309 VGND.t1949 VGND.t444 630.62
R1310 VGND.t1907 VGND.t136 630.62
R1311 VGND.t2112 VGND.t1082 630.62
R1312 VGND.t1080 VGND.t1264 630.62
R1313 VGND.t1246 VGND.t1078 630.62
R1314 VGND.t1947 VGND.t2570 630.62
R1315 VGND.t2609 VGND.t2668 630.62
R1316 VGND.t2658 VGND.t2339 630.62
R1317 VGND.t2493 VGND.t1693 630.62
R1318 VGND.t265 VGND.t1671 630.62
R1319 VGND.t2212 VGND.t2598 630.62
R1320 VGND.t754 VGND.t2320 630.62
R1321 VGND.t678 VGND.t2309 630.62
R1322 VGND.t2 VGND.t2594 630.62
R1323 VGND.t712 VGND.t2576 630.62
R1324 VGND.t789 VGND.t2322 630.62
R1325 VGND.t1096 VGND.t1658 630.62
R1326 VGND.t1979 VGND.t2642 630.62
R1327 VGND.t2153 VGND.t2304 630.62
R1328 VGND.t664 VGND.t2291 630.62
R1329 VGND.t323 VGND.t1699 630.62
R1330 VGND.t2366 VGND.t2295 630.62
R1331 VGND.n2704 VGND.n327 615.385
R1332 VGND.n2349 VGND.t1456 602.708
R1333 VGND.n3019 VGND.t1456 602.708
R1334 VGND.n3011 VGND.n3010 599.125
R1335 VGND.n194 VGND.n193 599.125
R1336 VGND.n66 VGND.n65 599.125
R1337 VGND.n117 VGND.n116 599.125
R1338 VGND.n134 VGND.n133 599.125
R1339 VGND.n165 VGND.n164 599.125
R1340 VGND.n2210 VGND.n2182 599.125
R1341 VGND.n2972 VGND.n2971 599.125
R1342 VGND VGND.t319 581.61
R1343 VGND.t1391 VGND 573.181
R1344 VGND VGND.t1549 573.181
R1345 VGND.t209 VGND 573.181
R1346 VGND.t652 VGND 573.181
R1347 VGND.n3013 VGND 564.751
R1348 VGND.t328 VGND 564.751
R1349 VGND.n3014 VGND 564.751
R1350 VGND.n3012 VGND 556.322
R1351 VGND.t1169 VGND 539.465
R1352 VGND VGND.t1133 539.465
R1353 VGND.t600 VGND.n806 494.779
R1354 VGND.n1166 VGND.t2287 492.058
R1355 VGND.t2637 VGND.n1175 492.058
R1356 VGND.n1176 VGND.t2613 492.058
R1357 VGND.t2285 VGND.n1188 492.058
R1358 VGND.n1189 VGND.t1706 492.058
R1359 VGND.t1684 VGND.n1207 492.058
R1360 VGND.n1208 VGND.t2352 492.058
R1361 VGND.t2332 VGND.n1220 492.058
R1362 VGND.n1247 VGND.t1679 492.058
R1363 VGND.n1246 VGND.t2596 492.058
R1364 VGND.n1240 VGND.t2585 492.058
R1365 VGND.n1239 VGND.t2307 492.058
R1366 VGND.n1233 VGND.t1669 492.058
R1367 VGND.t2574 VGND.n1277 492.058
R1368 VGND.n1278 VGND.t2318 492.058
R1369 VGND.t393 VGND.t354 481.877
R1370 VGND.t462 VGND.t393 481.877
R1371 VGND.t1436 VGND.t2216 481.877
R1372 VGND.t2216 VGND.t484 481.877
R1373 VGND.t2248 VGND 452.382
R1374 VGND.n1166 VGND.t497 424.312
R1375 VGND.n1175 VGND.t38 424.312
R1376 VGND.n1176 VGND.t1712 424.312
R1377 VGND.n1188 VGND.t764 424.312
R1378 VGND.n1189 VGND.t39 424.312
R1379 VGND.n1207 VGND.t767 424.312
R1380 VGND.n1208 VGND.t1292 424.312
R1381 VGND.n1220 VGND.t1171 424.312
R1382 VGND.n1247 VGND.t1295 424.312
R1383 VGND.t1445 VGND.n1246 424.312
R1384 VGND.n1240 VGND.t2371 424.312
R1385 VGND.t800 VGND.n1239 424.312
R1386 VGND.n1233 VGND.t72 424.312
R1387 VGND.n1277 VGND.t51 424.312
R1388 VGND.n1278 VGND.t884 424.312
R1389 VGND.t1217 VGND.n222 424.312
R1390 VGND.t366 VGND 419.68
R1391 VGND.n2284 VGND.n503 413.043
R1392 VGND.t1809 VGND.t1379 408.469
R1393 VGND.t283 VGND.t1270 408.469
R1394 VGND.t2401 VGND.t1966 408.469
R1395 VGND.t1529 VGND.t680 408.469
R1396 VGND.t1027 VGND.t858 408.469
R1397 VGND.t2040 VGND.t694 408.469
R1398 VGND.t1525 VGND.t2048 408.469
R1399 VGND.t106 VGND.t668 408.469
R1400 VGND.t421 VGND.t2016 408.469
R1401 VGND.t1472 VGND.t1933 408.469
R1402 VGND.t541 VGND.t1725 408.469
R1403 VGND.t2004 VGND.t1100 408.469
R1404 VGND.t1981 VGND.t1464 408.469
R1405 VGND.t728 VGND.t620 408.469
R1406 VGND.t893 VGND.t1598 408.469
R1407 VGND.t1584 VGND.t1636 408.469
R1408 VGND.t1884 VGND.t1009 408.469
R1409 VGND.t1498 VGND.t1311 408.469
R1410 VGND.t1958 VGND.t972 408.469
R1411 VGND.t2495 VGND.t1363 408.469
R1412 VGND.t534 VGND.t285 408.469
R1413 VGND.t1956 VGND.t1041 408.469
R1414 VGND.t80 VGND.t110 408.469
R1415 VGND.t2123 VGND.t1029 408.469
R1416 VGND.t798 VGND.t2042 408.469
R1417 VGND.t780 VGND.t1527 408.469
R1418 VGND.t585 VGND.t1353 408.469
R1419 VGND.t2469 VGND.t2028 408.469
R1420 VGND.t2414 VGND.t1760 408.469
R1421 VGND.t2162 VGND.t1729 408.469
R1422 VGND.t1260 VGND.t1638 408.469
R1423 VGND.t324 VGND.t1466 408.469
R1424 VGND.t2014 VGND.t1791 408.469
R1425 VGND.t2664 VGND.t1752 408.469
R1426 VGND.t1721 VGND.t2654 408.469
R1427 VGND.t1156 VGND.t901 408.469
R1428 VGND.t642 VGND.t1737 408.469
R1429 VGND.t700 VGND.t821 408.469
R1430 VGND.t889 VGND.t1987 408.469
R1431 VGND.t674 VGND.t1628 408.469
R1432 VGND.t993 VGND.t1121 408.469
R1433 VGND.t708 VGND.t271 408.469
R1434 VGND.t1383 VGND.t784 408.469
R1435 VGND.t2672 VGND.t1035 408.469
R1436 VGND.t2405 VGND.t1974 408.469
R1437 VGND.t1047 VGND.t734 408.469
R1438 VGND.t1361 VGND.t2554 408.469
R1439 VGND.t1591 VGND.t1624 408.469
R1440 VGND.t1833 VGND.t2036 408.469
R1441 VGND.t98 VGND.t1284 408.469
R1442 VGND.t2109 VGND.t1347 408.469
R1443 VGND.t1644 VGND.t1067 408.469
R1444 VGND.t986 VGND.t1754 408.469
R1445 VGND.t1325 VGND.t872 408.469
R1446 VGND.t750 VGND.t1630 408.469
R1447 VGND.t1458 VGND.t2243 408.469
R1448 VGND.t1150 VGND.t823 408.469
R1449 VGND.t891 VGND.t1112 408.469
R1450 VGND.t527 VGND.t1013 408.469
R1451 VGND.t815 VGND.t1092 408.469
R1452 VGND.t138 VGND.t978 408.469
R1453 VGND.t1502 VGND.t956 408.469
R1454 VGND.t1626 VGND.t13 408.469
R1455 VGND.t1253 VGND.t2409 408.469
R1456 VGND.t1543 VGND.t1905 408.469
R1457 VGND.t1021 VGND.t813 408.469
R1458 VGND.t1185 VGND.t1612 408.469
R1459 VGND.t1476 VGND.t2489 408.469
R1460 VGND.t259 VGND.t100 408.469
R1461 VGND.t2010 VGND.t2069 408.469
R1462 VGND.t76 VGND.t1460 408.469
R1463 VGND.t1756 VGND.t592 408.469
R1464 VGND.t792 VGND.t1329 408.469
R1465 VGND.t1632 VGND.t157 408.469
R1466 VGND.t580 VGND.t837 408.469
R1467 VGND.t1317 VGND.t2465 408.469
R1468 VGND.t1970 VGND.t200 408.469
R1469 VGND.t178 VGND.t2156 408.469
R1470 VGND.t269 VGND.t42 408.469
R1471 VGND.t338 VGND.t887 408.469
R1472 VGND.t1369 VGND.t1812 408.469
R1473 VGND.t275 VGND.t1268 408.469
R1474 VGND.t1964 VGND.t2391 408.469
R1475 VGND.t61 VGND.t1762 408.469
R1476 VGND.t856 VGND.t1017 408.469
R1477 VGND.t692 VGND.t2020 408.469
R1478 VGND.t2046 VGND.t1748 408.469
R1479 VGND.t666 VGND.t94 408.469
R1480 VGND.t419 VGND.t1998 408.469
R1481 VGND.t1931 VGND.t638 408.469
R1482 VGND.t538 VGND.t1713 408.469
R1483 VGND.t1098 VGND.t1648 408.469
R1484 VGND.t2419 VGND.t634 408.469
R1485 VGND.t726 VGND.t831 408.469
R1486 VGND.t976 VGND.t2417 408.469
R1487 VGND.t1582 VGND.t194 408.469
R1488 VGND.t999 VGND.t1785 408.469
R1489 VGND.t899 VGND.t2666 408.469
R1490 VGND.t960 VGND.t2656 408.469
R1491 VGND.t104 VGND.t1154 408.469
R1492 VGND.t277 VGND.t1739 408.469
R1493 VGND.t1535 VGND.t2210 408.469
R1494 VGND.t96 VGND.t1989 408.469
R1495 VGND.t1019 VGND.t676 408.469
R1496 VGND.t2026 VGND.t0 408.469
R1497 VGND.t1750 VGND.t710 408.469
R1498 VGND.t1341 VGND.t786 408.469
R1499 VGND.t1478 VGND.t2674 408.469
R1500 VGND.t1976 VGND.t1746 408.469
R1501 VGND.t736 VGND.t1715 408.469
R1502 VGND.t196 VGND.t2556 408.469
R1503 VGND.t332 VGND.t636 408.469
R1504 VGND.t1827 VGND.t1996 408.469
R1505 VGND.t1735 VGND.t1286 408.469
R1506 VGND.t1331 VGND.t2091 408.469
R1507 VGND.t885 VGND.t1065 408.469
R1508 VGND.t988 VGND.t626 408.469
R1509 VGND.t289 VGND.t874 408.469
R1510 VGND.t752 VGND.t966 408.469
R1511 VGND.t188 VGND.t2245 408.469
R1512 VGND.t1214 VGND.t1033 408.469
R1513 VGND.t2399 VGND.t1114 408.469
R1514 VGND.t529 VGND.t1375 408.469
R1515 VGND.t1023 VGND.t1094 408.469
R1516 VGND.t140 VGND.t2393 408.469
R1517 VGND.t1039 VGND.t1504 408.469
R1518 VGND.t1349 VGND.t33 408.469
R1519 VGND.t1255 VGND.t1614 408.469
R1520 VGND.t1480 VGND.t1839 408.469
R1521 VGND.t90 VGND.t1279 408.469
R1522 VGND.t2103 VGND.t1339 408.469
R1523 VGND.t198 VGND.t1071 408.469
R1524 VGND.t1742 VGND.t982 408.469
R1525 VGND.t1313 VGND.t169 408.469
R1526 VGND.t190 VGND.t2055 408.469
R1527 VGND.t628 VGND.t2239 408.469
R1528 VGND.t291 VGND.t1146 408.469
R1529 VGND.t970 VGND.t1227 408.469
R1530 VGND.t1003 VGND.t525 408.469
R1531 VGND.t281 VGND.t1090 408.469
R1532 VGND.t2425 VGND.t962 408.469
R1533 VGND.t1415 VGND.t1377 408.469
R1534 VGND.t1616 VGND.t9 408.469
R1535 VGND.t1251 VGND.t2395 408.469
R1536 VGND.t1533 VGND.t1767 408.469
R1537 VGND.t1015 VGND.t811 408.469
R1538 VGND.t1610 VGND.t1183 408.469
R1539 VGND.t640 VGND.t2491 408.469
R1540 VGND.t92 VGND.t257 408.469
R1541 VGND.t1650 VGND.t2067 408.469
R1542 VGND.t630 VGND.t74 408.469
R1543 VGND.t1744 VGND.t590 408.469
R1544 VGND.t1315 VGND.t3 408.469
R1545 VGND.t192 VGND.t155 408.469
R1546 VGND.t829 VGND.t790 408.469
R1547 VGND.t907 VGND.t2463 408.469
R1548 VGND.t1968 VGND.t186 408.469
R1549 VGND.t2154 VGND.t1005 408.469
R1550 VGND.t2397 VGND.t40 408.469
R1551 VGND.t336 VGND.t964 408.469
R1552 VGND.t1863 VGND.t1007 408.469
R1553 VGND.t2166 VGND.t905 408.469
R1554 VGND.t250 VGND.t968 408.469
R1555 VGND.t112 VGND.t1058 408.469
R1556 VGND.t279 VGND.t2228 408.469
R1557 VGND.t1545 VGND.t2086 408.469
R1558 VGND.t102 VGND.t2252 408.469
R1559 VGND.t1025 VGND.t2513 408.469
R1560 VGND.t2038 VGND.t773 408.469
R1561 VGND.t1764 VGND.t2096 408.469
R1562 VGND.t1351 VGND.t505 408.469
R1563 VGND.t344 VGND.t2022 408.469
R1564 VGND.t1337 VGND.t1758 408.469
R1565 VGND.t2118 VGND.t1723 408.469
R1566 VGND.t5 VGND.t1634 408.469
R1567 VGND.t1243 VGND.t1462 408.469
R1568 VGND.t1531 VGND.t1794 408.469
R1569 VGND.t1620 VGND.t2662 408.469
R1570 VGND.t1606 VGND.t2652 408.469
R1571 VGND.t1158 VGND.t632 408.469
R1572 VGND.t1359 VGND.t863 408.469
R1573 VGND.t698 VGND.t1646 408.469
R1574 VGND.t624 VGND.t1985 408.469
R1575 VGND.t672 VGND.t1733 408.469
R1576 VGND.t1309 VGND.t1119 408.469
R1577 VGND.t184 VGND.t706 408.469
R1578 VGND.t545 VGND.t825 408.469
R1579 VGND.t2670 VGND.t903 408.469
R1580 VGND.t182 VGND.t1972 408.469
R1581 VGND.t995 VGND.t732 408.469
R1582 VGND.t2389 VGND.t2552 408.469
R1583 VGND.t1589 VGND.t958 408.469
R1584 VGND.t1866 VGND.t1622 408.469
R1585 VGND.t1367 VGND.t2164 408.469
R1586 VGND.t704 VGND.t108 408.469
R1587 VGND.t2018 VGND.t1060 408.469
R1588 VGND.t2226 VGND.t1537 408.469
R1589 VGND.t1727 VGND.t245 408.469
R1590 VGND.t2250 VGND.t2008 408.469
R1591 VGND.t2030 VGND.t2511 408.469
R1592 VGND.t771 VGND.t622 408.469
R1593 VGND.t1327 VGND.t2094 408.469
R1594 VGND.t503 VGND.t1640 408.469
R1595 VGND.t721 VGND.t833 408.469
R1596 VGND.t1335 VGND.t1319 408.469
R1597 VGND.t2116 VGND.t897 408.469
R1598 VGND.t1037 VGND.t17 408.469
R1599 VGND.t295 VGND.t817 408.469
R1600 VGND.t2403 VGND.t1896 408.469
R1601 VGND.t1496 VGND.t997 408.469
R1602 VGND.t1031 VGND.t1189 408.469
R1603 VGND.t1604 VGND.t713 408.469
R1604 VGND.t1371 VGND.t263 408.469
R1605 VGND.t1355 VGND.t1954 408.469
R1606 VGND.t2032 VGND.t78 408.469
R1607 VGND.t1539 VGND.t2121 408.469
R1608 VGND.t1731 VGND.t796 408.469
R1609 VGND.t778 VGND.t2012 408.469
R1610 VGND.t582 VGND.t1468 408.469
R1611 VGND.t1719 VGND.t2467 408.469
R1612 VGND.t2000 VGND.t2411 408.469
R1613 VGND.t2160 VGND.t1642 408.469
R1614 VGND.t1257 VGND.t819 408.469
R1615 VGND.t321 VGND.t1321 408.469
R1616 VGND.t974 VGND.t1836 408.469
R1617 VGND.t827 VGND.t1281 408.469
R1618 VGND.t287 VGND.t2105 408.469
R1619 VGND.t1069 VGND.t1043 408.469
R1620 VGND.t984 VGND.t1001 408.469
R1621 VGND.t171 VGND.t1618 408.469
R1622 VGND.t2053 VGND.t1541 408.469
R1623 VGND.t2237 VGND.t1373 408.469
R1624 VGND.t1144 VGND.t1357 408.469
R1625 VGND.t2034 VGND.t1225 408.469
R1626 VGND.t1523 VGND.t523 408.469
R1627 VGND.t1345 VGND.t1088 408.469
R1628 VGND.t2024 VGND.t2423 408.469
R1629 VGND.t1413 VGND.t1470 408.469
R1630 VGND.t1323 VGND.t11 408.469
R1631 VGND.t1249 VGND.t2002 408.469
R1632 VGND.t1690 VGND.t1474 408.469
R1633 VGND.t1343 VGND.t2607 408.469
R1634 VGND.t2006 VGND.t2336 408.469
R1635 VGND.t180 VGND.t2314 408.469
R1636 VGND.t1717 VGND.t2602 408.469
R1637 VGND.t895 VGND.t2591 408.469
R1638 VGND.t1011 VGND.t2572 408.469
R1639 VGND.t835 VGND.t1675 408.469
R1640 VGND.t273 VGND.t1654 408.469
R1641 VGND.t1385 VGND.t2568 408.469
R1642 VGND.t991 VGND.t2302 408.469
R1643 VGND.t2407 VGND.t2289 408.469
R1644 VGND.t1381 VGND.t2626 408.469
R1645 VGND.t1365 VGND.t2362 408.469
R1646 VGND.t1608 VGND.t1704 408.469
R1647 VGND.t2635 VGND.t1045 408.469
R1648 VGND.t464 VGND.t362 397.848
R1649 VGND.t362 VGND.t352 397.848
R1650 VGND.t352 VGND.t439 397.848
R1651 VGND.t439 VGND.t1551 397.848
R1652 VGND.t1551 VGND.t1552 397.848
R1653 VGND.t1552 VGND.t1555 397.848
R1654 VGND.t1555 VGND.t1556 397.848
R1655 VGND.t1918 VGND.t1194 396.17
R1656 VGND.t762 VGND.t237 396.17
R1657 VGND.n2935 VGND.n2934 394.137
R1658 VGND.n2933 VGND.n208 394.137
R1659 VGND.n2932 VGND.n209 394.137
R1660 VGND.n2931 VGND.n210 394.137
R1661 VGND.n2930 VGND.n211 394.137
R1662 VGND.n2929 VGND.n212 394.137
R1663 VGND.n2928 VGND.n213 394.137
R1664 VGND.n2927 VGND.n214 394.137
R1665 VGND.n2926 VGND.n215 394.137
R1666 VGND.n2925 VGND.n216 394.137
R1667 VGND.n2924 VGND.n217 394.137
R1668 VGND.n2923 VGND.n218 394.137
R1669 VGND.n2922 VGND.n219 394.137
R1670 VGND.n2921 VGND.n220 394.137
R1671 VGND.n2920 VGND.n221 394.137
R1672 VGND.n2919 VGND.n2918 394.137
R1673 VGND.n2285 VGND.t63 387.421
R1674 VGND.n2284 VGND.t1136 387.421
R1675 VGND.n2250 VGND.t114 387.421
R1676 VGND.n2248 VGND.t66 387.421
R1677 VGND.n1386 VGND.t488 387.421
R1678 VGND.t238 VGND.t768 362.452
R1679 VGND.t768 VGND.t1169 345.594
R1680 VGND VGND.t551 328.616
R1681 VGND VGND.t364 328.616
R1682 VGND VGND.t548 328.616
R1683 VGND VGND.t602 328.616
R1684 VGND VGND.t330 328.616
R1685 VGND.t2645 VGND.t2293 313.776
R1686 VGND.t2639 VGND.t2565 313.776
R1687 VGND.t2361 VGND.t2368 313.776
R1688 VGND.t2346 VGND.t1702 313.776
R1689 VGND.t2633 VGND.t2281 313.776
R1690 VGND.t2617 VGND.t2349 313.776
R1691 VGND.t2284 VGND.t2604 313.776
R1692 VGND.t2275 VGND.t1692 313.776
R1693 VGND.t2606 VGND.t1686 313.776
R1694 VGND.t2619 VGND.t2350 313.776
R1695 VGND.t1689 VGND.t2334 313.776
R1696 VGND.t2325 VGND.t1677 313.776
R1697 VGND.t2593 VGND.t2600 313.776
R1698 VGND.t2588 VGND.t2327 313.776
R1699 VGND.t2306 VGND.t2566 313.776
R1700 VGND.t1673 VGND.t2590 313.776
R1701 VGND.t1927 VGND.t1918 311.877
R1702 VGND.t319 VGND.t762 311.877
R1703 VGND VGND.t1923 303.449
R1704 VGND VGND.t1927 295.019
R1705 VGND.n101 VGND.t355 287.832
R1706 VGND VGND.t1305 286.591
R1707 VGND.n93 VGND.t476 282.327
R1708 VGND.n2184 VGND.t1453 282.327
R1709 VGND.n104 VGND.t2455 281.13
R1710 VGND.n2189 VGND.t492 281.13
R1711 VGND.n177 VGND.t435 280.978
R1712 VGND.n177 VGND.t402 280.978
R1713 VGND.n78 VGND.t2458 280.978
R1714 VGND.n78 VGND.t452 280.978
R1715 VGND.n146 VGND.t392 280.978
R1716 VGND.n146 VGND.t457 280.978
R1717 VGND.n482 VGND.t1432 280.978
R1718 VGND.n482 VGND.t1450 280.978
R1719 VGND.n2263 VGND.t493 280.978
R1720 VGND.n2263 VGND.t2215 280.978
R1721 VGND.n518 VGND.t2256 280.978
R1722 VGND.n518 VGND.t1447 280.978
R1723 VGND.n2194 VGND.t485 280.978
R1724 VGND.t2083 VGND 278.161
R1725 VGND.n2970 VGND 271.014
R1726 VGND.n3021 VGND.n4 259.389
R1727 VGND.n2347 VGND.n4 259.389
R1728 VGND.n3022 VGND.n3 252.988
R1729 VGND VGND.t378 252.875
R1730 VGND VGND.t1925 252.875
R1731 VGND VGND.t1920 252.875
R1732 VGND VGND.t408 252.875
R1733 VGND.t398 VGND 252.875
R1734 VGND.n887 VGND.t1475 241.393
R1735 VGND.n330 VGND.t1822 241.393
R1736 VGND.n396 VGND.t1380 241.393
R1737 VGND.n400 VGND.t1010 241.393
R1738 VGND.n469 VGND.t2015 241.393
R1739 VGND.n466 VGND.t2037 241.393
R1740 VGND.n625 VGND.t1544 241.393
R1741 VGND.n590 VGND.t1370 241.393
R1742 VGND.n587 VGND.t1000 241.393
R1743 VGND.n547 VGND.t1997 241.393
R1744 VGND.n628 VGND.t1481 241.393
R1745 VGND.n632 VGND.t1534 241.393
R1746 VGND.n879 VGND.t1008 241.393
R1747 VGND.n800 VGND.t1532 241.393
R1748 VGND.n797 VGND.t1623 241.393
R1749 VGND.n882 VGND.t2404 241.393
R1750 VGND.n1024 VGND.t975 241.393
R1751 VGND.n1014 VGND.t1825 241.393
R1752 VGND.n1333 VGND.t1344 241.284
R1753 VGND.n894 VGND.t2007 241.284
R1754 VGND.n932 VGND.t181 241.284
R1755 VGND.n937 VGND.t1718 241.284
R1756 VGND.n942 VGND.t896 241.284
R1757 VGND.n947 VGND.t1012 241.284
R1758 VGND.n952 VGND.t836 241.284
R1759 VGND.n957 VGND.t274 241.284
R1760 VGND.n962 VGND.t1386 241.284
R1761 VGND.n967 VGND.t992 241.284
R1762 VGND.n972 VGND.t2408 241.284
R1763 VGND.n977 VGND.t1382 241.284
R1764 VGND.n982 VGND.t1366 241.284
R1765 VGND.n987 VGND.t1609 241.284
R1766 VGND.n1280 VGND.t1861 241.284
R1767 VGND.n1275 VGND.t1819 241.284
R1768 VGND.n1232 VGND.t1903 241.284
R1769 VGND.n1237 VGND.t1894 241.284
R1770 VGND.n1225 VGND.t1855 241.284
R1771 VGND.n1244 VGND.t1807 241.284
R1772 VGND.n1001 VGND.t1891 241.284
R1773 VGND.n1218 VGND.t1852 241.284
R1774 VGND.n1210 VGND.t1843 241.284
R1775 VGND.n1205 VGND.t1801 241.284
R1776 VGND.n1009 VGND.t1879 241.284
R1777 VGND.n1186 VGND.t1873 241.284
R1778 VGND.n1178 VGND.t1798 241.284
R1779 VGND.n1173 VGND.t1780 241.284
R1780 VGND.n1168 VGND.t1774 241.284
R1781 VGND.n2773 VGND.t1858 241.284
R1782 VGND.n294 VGND.t1816 241.284
R1783 VGND.n2730 VGND.t1900 241.284
R1784 VGND.n2735 VGND.t1888 241.284
R1785 VGND.n312 VGND.t1849 241.284
R1786 VGND.n2726 VGND.t1804 241.284
R1787 VGND.n326 VGND.t1882 241.284
R1788 VGND.n387 VGND.t1846 241.284
R1789 VGND.n384 VGND.t1831 241.284
R1790 VGND.n379 VGND.t1789 241.284
R1791 VGND.n373 VGND.t1876 241.284
R1792 VGND.n368 VGND.t1870 241.284
R1793 VGND.n362 VGND.t1783 241.284
R1794 VGND.n355 VGND.t1777 241.284
R1795 VGND.n2699 VGND.t1771 241.284
R1796 VGND.n2639 VGND.t284 241.284
R1797 VGND.n2644 VGND.t2402 241.284
R1798 VGND.n2649 VGND.t1530 241.284
R1799 VGND.n2654 VGND.t1028 241.284
R1800 VGND.n2659 VGND.t2041 241.284
R1801 VGND.n2664 VGND.t1526 241.284
R1802 VGND.n2669 VGND.t107 241.284
R1803 VGND.n394 VGND.t2017 241.284
R1804 VGND.n2715 VGND.t1473 241.284
R1805 VGND.n320 VGND.t1726 241.284
R1806 VGND.n2748 VGND.t2005 241.284
R1807 VGND.n304 VGND.t1465 241.284
R1808 VGND.n2753 VGND.t621 241.284
R1809 VGND.n2788 VGND.t894 241.284
R1810 VGND.n287 VGND.t1637 241.284
R1811 VGND.n2343 VGND.t1312 241.284
R1812 VGND.n2338 VGND.t973 241.284
R1813 VGND.n2333 VGND.t1364 241.284
R1814 VGND.n2328 VGND.t286 241.284
R1815 VGND.n2323 VGND.t1042 241.284
R1816 VGND.n2318 VGND.t111 241.284
R1817 VGND.n2313 VGND.t1030 241.284
R1818 VGND.n2308 VGND.t2043 241.284
R1819 VGND.n2303 VGND.t1528 241.284
R1820 VGND.n2298 VGND.t1354 241.284
R1821 VGND.n2293 VGND.t2029 241.284
R1822 VGND.n2288 VGND.t1761 241.284
R1823 VGND.n415 VGND.t1730 241.284
R1824 VGND.n2541 VGND.t1639 241.284
R1825 VGND.n2536 VGND.t1467 241.284
R1826 VGND.n472 VGND.t1753 241.284
R1827 VGND.n2377 VGND.t1722 241.284
R1828 VGND.n460 VGND.t902 241.284
R1829 VGND.n2403 VGND.t643 241.284
R1830 VGND.n452 VGND.t822 241.284
R1831 VGND.n2429 VGND.t890 241.284
R1832 VGND.n444 VGND.t1629 241.284
R1833 VGND.n2455 VGND.t994 241.284
R1834 VGND.n436 VGND.t272 241.284
R1835 VGND.n2481 VGND.t1384 241.284
R1836 VGND.n428 VGND.t1036 241.284
R1837 VGND.n2512 VGND.t2406 241.284
R1838 VGND.n2517 VGND.t1048 241.284
R1839 VGND.n2522 VGND.t1362 241.284
R1840 VGND.n2527 VGND.t1625 241.284
R1841 VGND.n2364 VGND.t99 241.284
R1842 VGND.n464 VGND.t1348 241.284
R1843 VGND.n2390 VGND.t1645 241.284
R1844 VGND.n456 VGND.t1755 241.284
R1845 VGND.n2416 VGND.t1326 241.284
R1846 VGND.n448 VGND.t1631 241.284
R1847 VGND.n2442 VGND.t1459 241.284
R1848 VGND.n440 VGND.t824 241.284
R1849 VGND.n2468 VGND.t892 241.284
R1850 VGND.n432 VGND.t1014 241.284
R1851 VGND.n2494 VGND.t816 241.284
R1852 VGND.n424 VGND.t979 241.284
R1853 VGND.n2499 VGND.t957 241.284
R1854 VGND.n2810 VGND.t1627 241.284
R1855 VGND.n2815 VGND.t2410 241.284
R1856 VGND.n1911 VGND.t1022 241.284
R1857 VGND.n623 VGND.t1613 241.284
R1858 VGND.n1922 VGND.t1477 241.284
R1859 VGND.n620 VGND.t101 241.284
R1860 VGND.n1933 VGND.t2011 241.284
R1861 VGND.n617 VGND.t1461 241.284
R1862 VGND.n1944 VGND.t1757 241.284
R1863 VGND.n614 VGND.t1330 241.284
R1864 VGND.n1955 VGND.t1633 241.284
R1865 VGND.n611 VGND.t838 241.284
R1866 VGND.n1966 VGND.t1318 241.284
R1867 VGND.n608 VGND.t201 241.284
R1868 VGND.n1977 VGND.t179 241.284
R1869 VGND.n1982 VGND.t270 241.284
R1870 VGND.n1987 VGND.t888 241.284
R1871 VGND.n597 VGND.t276 241.284
R1872 VGND.n594 VGND.t2392 241.284
R1873 VGND.n2056 VGND.t1763 241.284
R1874 VGND.n2051 VGND.t1018 241.284
R1875 VGND.n2046 VGND.t2021 241.284
R1876 VGND.n2041 VGND.t1749 241.284
R1877 VGND.n2036 VGND.t95 241.284
R1878 VGND.n2031 VGND.t1999 241.284
R1879 VGND.n2026 VGND.t639 241.284
R1880 VGND.n2021 VGND.t1714 241.284
R1881 VGND.n2016 VGND.t1649 241.284
R1882 VGND.n2011 VGND.t635 241.284
R1883 VGND.n2006 VGND.t832 241.284
R1884 VGND.n2001 VGND.t977 241.284
R1885 VGND.n1994 VGND.t195 241.284
R1886 VGND.n2070 VGND.t900 241.284
R1887 VGND.n2075 VGND.t961 241.284
R1888 VGND.n2080 VGND.t105 241.284
R1889 VGND.n2085 VGND.t278 241.284
R1890 VGND.n2090 VGND.t1536 241.284
R1891 VGND.n2095 VGND.t97 241.284
R1892 VGND.n2100 VGND.t1020 241.284
R1893 VGND.n2105 VGND.t2027 241.284
R1894 VGND.n2110 VGND.t1751 241.284
R1895 VGND.n2115 VGND.t1342 241.284
R1896 VGND.n2120 VGND.t1479 241.284
R1897 VGND.n585 VGND.t1747 241.284
R1898 VGND.n2125 VGND.t1716 241.284
R1899 VGND.n2835 VGND.t197 241.284
R1900 VGND.n2840 VGND.t637 241.284
R1901 VGND.n2177 VGND.t1736 241.284
R1902 VGND.n1756 VGND.t1332 241.284
R1903 VGND.n1762 VGND.t886 241.284
R1904 VGND.n1753 VGND.t627 241.284
R1905 VGND.n1773 VGND.t290 241.284
R1906 VGND.n1750 VGND.t967 241.284
R1907 VGND.n1784 VGND.t189 241.284
R1908 VGND.n1747 VGND.t1034 241.284
R1909 VGND.n1795 VGND.t2400 241.284
R1910 VGND.n1744 VGND.t1376 241.284
R1911 VGND.n1806 VGND.t1024 241.284
R1912 VGND.n1741 VGND.t2394 241.284
R1913 VGND.n1817 VGND.t1040 241.284
R1914 VGND.n1822 VGND.t1350 241.284
R1915 VGND.n1827 VGND.t1615 241.284
R1916 VGND.n1679 VGND.t91 241.284
R1917 VGND.n1676 VGND.t1340 241.284
R1918 VGND.n1690 VGND.t199 241.284
R1919 VGND.n1695 VGND.t1743 241.284
R1920 VGND.n1700 VGND.t1314 241.284
R1921 VGND.n1705 VGND.t191 241.284
R1922 VGND.n1710 VGND.t629 241.284
R1923 VGND.n1715 VGND.t292 241.284
R1924 VGND.n1720 VGND.t971 241.284
R1925 VGND.n1725 VGND.t1004 241.284
R1926 VGND.n1730 VGND.t282 241.284
R1927 VGND.n1673 VGND.t963 241.284
R1928 VGND.n1846 VGND.t1378 241.284
R1929 VGND.n1841 VGND.t1617 241.284
R1930 VGND.n1834 VGND.t2396 241.284
R1931 VGND.n670 VGND.t1016 241.284
R1932 VGND.n675 VGND.t1611 241.284
R1933 VGND.n680 VGND.t641 241.284
R1934 VGND.n685 VGND.t93 241.284
R1935 VGND.n690 VGND.t1651 241.284
R1936 VGND.n695 VGND.t631 241.284
R1937 VGND.n700 VGND.t1745 241.284
R1938 VGND.n705 VGND.t1316 241.284
R1939 VGND.n710 VGND.t193 241.284
R1940 VGND.n715 VGND.t830 241.284
R1941 VGND.n720 VGND.t908 241.284
R1942 VGND.n667 VGND.t187 241.284
R1943 VGND.n725 VGND.t1006 241.284
R1944 VGND.n2860 VGND.t2398 241.284
R1945 VGND.n2865 VGND.t965 241.284
R1946 VGND.n1353 VGND.t906 241.284
R1947 VGND.n875 VGND.t969 241.284
R1948 VGND.n870 VGND.t113 241.284
R1949 VGND.n810 VGND.t280 241.284
R1950 VGND.n824 VGND.t1546 241.284
R1951 VGND.n829 VGND.t103 241.284
R1952 VGND.n834 VGND.t1026 241.284
R1953 VGND.n839 VGND.t2039 241.284
R1954 VGND.n844 VGND.t1765 241.284
R1955 VGND.n849 VGND.t1352 241.284
R1956 VGND.n820 VGND.t2023 241.284
R1957 VGND.n854 VGND.t1759 241.284
R1958 VGND.n735 VGND.t1724 241.284
R1959 VGND.n1662 VGND.t1635 241.284
R1960 VGND.n1657 VGND.t1463 241.284
R1961 VGND.n1391 VGND.t1621 241.284
R1962 VGND.n1396 VGND.t1607 241.284
R1963 VGND.n805 VGND.t633 241.284
R1964 VGND.n1491 VGND.t1360 241.284
R1965 VGND.n777 VGND.t1647 241.284
R1966 VGND.n1517 VGND.t625 241.284
R1967 VGND.n769 VGND.t1734 241.284
R1968 VGND.n1543 VGND.t1310 241.284
R1969 VGND.n1548 VGND.t185 241.284
R1970 VGND.n761 VGND.t826 241.284
R1971 VGND.n1553 VGND.t904 241.284
R1972 VGND.n1633 VGND.t183 241.284
R1973 VGND.n1638 VGND.t996 241.284
R1974 VGND.n1643 VGND.t2390 241.284
R1975 VGND.n1648 VGND.t959 241.284
R1976 VGND.n1411 VGND.t1368 241.284
R1977 VGND.n795 VGND.t109 241.284
R1978 VGND.n1478 VGND.t2019 241.284
R1979 VGND.n781 VGND.t1538 241.284
R1980 VGND.n1504 VGND.t1728 241.284
R1981 VGND.n773 VGND.t2009 241.284
R1982 VGND.n1530 VGND.t2031 241.284
R1983 VGND.n765 VGND.t623 241.284
R1984 VGND.n1567 VGND.t1328 241.284
R1985 VGND.n756 VGND.t1641 241.284
R1986 VGND.n1582 VGND.t834 241.284
R1987 VGND.n1577 VGND.t1320 241.284
R1988 VGND.n1572 VGND.t898 241.284
R1989 VGND.n2885 VGND.t1038 241.284
R1990 VGND.n2890 VGND.t818 241.284
R1991 VGND.n885 VGND.t998 241.284
R1992 VGND.n1424 VGND.t1032 241.284
R1993 VGND.n1429 VGND.t1605 241.284
R1994 VGND.n1434 VGND.t1372 241.284
R1995 VGND.n1439 VGND.t1356 241.284
R1996 VGND.n1444 VGND.t2033 241.284
R1997 VGND.n1449 VGND.t1540 241.284
R1998 VGND.n1454 VGND.t1732 241.284
R1999 VGND.n791 VGND.t2013 241.284
R2000 VGND.n1459 VGND.t1469 241.284
R2001 VGND.n1596 VGND.t1720 241.284
R2002 VGND.n1601 VGND.t2001 241.284
R2003 VGND.n750 VGND.t1643 241.284
R2004 VGND.n1614 VGND.t820 241.284
R2005 VGND.n1609 VGND.t1322 241.284
R2006 VGND.n1032 VGND.t828 241.284
R2007 VGND.n1037 VGND.t288 241.284
R2008 VGND.n1029 VGND.t1044 241.284
R2009 VGND.n1095 VGND.t1002 241.284
R2010 VGND.n1090 VGND.t1619 241.284
R2011 VGND.n1085 VGND.t1542 241.284
R2012 VGND.n1080 VGND.t1374 241.284
R2013 VGND.n1075 VGND.t1358 241.284
R2014 VGND.n1070 VGND.t2035 241.284
R2015 VGND.n1043 VGND.t1524 241.284
R2016 VGND.n1053 VGND.t1346 241.284
R2017 VGND.n1058 VGND.t2025 241.284
R2018 VGND.n1049 VGND.t1471 241.284
R2019 VGND.n2905 VGND.t1324 241.284
R2020 VGND.n2910 VGND.t2003 241.284
R2021 VGND.n928 VGND.t1046 241.284
R2022 VGND.t1379 VGND.t944 222.15
R2023 VGND.t1594 VGND.t1208 222.15
R2024 VGND.t2518 VGND.t283 222.15
R2025 VGND.t52 VGND.t253 222.15
R2026 VGND.t952 VGND.t2401 222.15
R2027 VGND.t1167 VGND.t59 222.15
R2028 VGND.t950 VGND.t1529 222.15
R2029 VGND.t619 VGND.t855 222.15
R2030 VGND.t2526 VGND.t1027 222.15
R2031 VGND.t1172 VGND.t167 222.15
R2032 VGND.t2534 VGND.t2040 222.15
R2033 VGND.t2220 VGND.t2428 222.15
R2034 VGND.t2532 VGND.t1525 222.15
R2035 VGND.t1492 VGND.t2516 222.15
R2036 VGND.t2524 VGND.t106 222.15
R2037 VGND.t495 VGND.t1142 222.15
R2038 VGND.t2016 VGND.t2522 222.15
R2039 VGND.t1108 VGND.t1241 222.15
R2040 VGND.t2536 VGND.t1472 222.15
R2041 VGND.t720 VGND.t508 222.15
R2042 VGND.t1725 VGND.t948 222.15
R2043 VGND.t2450 VGND.t55 222.15
R2044 VGND.t946 VGND.t2004 222.15
R2045 VGND.t2660 VGND.t2422 222.15
R2046 VGND.t1464 VGND.t2530 222.15
R2047 VGND.t1411 VGND.t560 222.15
R2048 VGND.t620 VGND.t2528 222.15
R2049 VGND.t8 VGND.t204 222.15
R2050 VGND.t954 VGND.t893 222.15
R2051 VGND.t1109 VGND.t1581 222.15
R2052 VGND.t1636 VGND.t2520 222.15
R2053 VGND.t2623 VGND.t747 222.15
R2054 VGND.t1009 VGND.t2682 222.15
R2055 VGND.t1273 VGND.t2482 222.15
R2056 VGND.t1311 VGND.t2063 222.15
R2057 VGND.t2651 VGND.t176 222.15
R2058 VGND.t972 VGND.t610 222.15
R2059 VGND.t1153 VGND.t1211 222.15
R2060 VGND.t1363 VGND.t1408 222.15
R2061 VGND.t262 VGND.t2099 222.15
R2062 VGND.t285 VGND.t2680 222.15
R2063 VGND.t697 VGND.t1266 222.15
R2064 VGND.t1041 VGND.t2059 222.15
R2065 VGND.t2052 VGND.t2506 222.15
R2066 VGND.t110 VGND.t2057 222.15
R2067 VGND.t671 VGND.t470 222.15
R2068 VGND.t1029 VGND.t2678 222.15
R2069 VGND.t1118 VGND.t1995 222.15
R2070 VGND.t2042 VGND.t2676 222.15
R2071 VGND.t1936 VGND.t661 222.15
R2072 VGND.t1527 VGND.t2061 222.15
R2073 VGND.t788 VGND.t1388 222.15
R2074 VGND.t1353 VGND.t1420 222.15
R2075 VGND.t349 VGND.t618 222.15
R2076 VGND.t2028 VGND.t1418 222.15
R2077 VGND.t1978 VGND.t2077 222.15
R2078 VGND.t1760 VGND.t616 222.15
R2079 VGND.t731 VGND.t2093 222.15
R2080 VGND.t1729 VGND.t614 222.15
R2081 VGND.t2558 VGND.t924 222.15
R2082 VGND.t1638 VGND.t612 222.15
R2083 VGND.t341 VGND.t1518 222.15
R2084 VGND.t1466 VGND.t2065 222.15
R2085 VGND.t2283 VGND.t2225 222.15
R2086 VGND.t2141 VGND.t2014 222.15
R2087 VGND.t1389 VGND.t1278 222.15
R2088 VGND.t1752 VGND.t1426 222.15
R2089 VGND.t2107 VGND.t561 222.15
R2090 VGND.t2149 VGND.t1721 222.15
R2091 VGND.t127 VGND.t1063 222.15
R2092 VGND.t901 VGND.t2147 222.15
R2093 VGND.t861 VGND.t1125 222.15
R2094 VGND.t2139 VGND.t642 222.15
R2095 VGND.t1942 VGND.t173 222.15
R2096 VGND.t821 VGND.t1422 222.15
R2097 VGND.t2430 VGND.t2480 222.15
R2098 VGND.t2686 VGND.t889 222.15
R2099 VGND.t1291 VGND.t2241 222.15
R2100 VGND.t1628 VGND.t2137 222.15
R2101 VGND.t1148 VGND.t2484 222.15
R2102 VGND.t1430 VGND.t993 222.15
R2103 VGND.t1909 VGND.t1110 222.15
R2104 VGND.t271 VGND.t1424 222.15
R2105 VGND.t532 VGND.t1596 222.15
R2106 VGND.t2145 VGND.t1383 222.15
R2107 VGND.t723 VGND.t2452 222.15
R2108 VGND.t1035 VGND.t2143 222.15
R2109 VGND.t143 VGND.t766 222.15
R2110 VGND.t2684 VGND.t2405 222.15
R2111 VGND.t44 VGND.t1417 222.15
R2112 VGND.t1443 VGND.t1047 222.15
R2113 VGND.t164 VGND.t36 222.15
R2114 VGND.t2151 VGND.t1361 222.15
R2115 VGND.t852 VGND.t1587 222.15
R2116 VGND.t1624 VGND.t1428 222.15
R2117 VGND.t2644 VGND.t2438 222.15
R2118 VGND.t2036 VGND.t2443 222.15
R2119 VGND.t2235 VGND.t558 222.15
R2120 VGND.t233 VGND.t98 222.15
R2121 VGND.t255 VGND.t702 222.15
R2122 VGND.t1347 VGND.t606 222.15
R2123 VGND.t715 VGND.t2648 222.15
R2124 VGND.t604 VGND.t1644 222.15
R2125 VGND.t879 VGND.t980 222.15
R2126 VGND.t1754 VGND.t2441 222.15
R2127 VGND.t243 VGND.t1242 222.15
R2128 VGND.t229 VGND.t1325 222.15
R2129 VGND.t1126 VGND.t1993 222.15
R2130 VGND.t1630 VGND.t227 222.15
R2131 VGND.t2509 VGND.t940 222.15
R2132 VGND.t2439 VGND.t1458 222.15
R2133 VGND.t162 VGND.t82 222.15
R2134 VGND.t823 VGND.t2135 222.15
R2135 VGND.t1221 VGND.t2111 222.15
R2136 VGND.t231 VGND.t891 222.15
R2137 VGND.t559 VGND.t501 222.15
R2138 VGND.t1013 VGND.t2447 222.15
R2139 VGND.t1951 VGND.t1213 222.15
R2140 VGND.t2445 VGND.t815 222.15
R2141 VGND.t1104 VGND.t1333 222.15
R2142 VGND.t978 VGND.t225 222.15
R2143 VGND.t2114 VGND.t1274 222.15
R2144 VGND.t956 VGND.t223 222.15
R2145 VGND.t15 VGND.t1097 222.15
R2146 VGND.t608 VGND.t1626 222.15
R2147 VGND.t45 VGND.t1247 222.15
R2148 VGND.t2409 VGND.t2133 222.15
R2149 VGND.t2578 VGND.t50 222.15
R2150 VGND.t124 VGND.t1543 222.15
R2151 VGND.t1568 VGND.t1267 222.15
R2152 VGND.t936 VGND.t1021 222.15
R2153 VGND.t206 VGND.t1963 222.15
R2154 VGND.t1612 VGND.t2474 222.15
R2155 VGND.t679 VGND.t1941 222.15
R2156 VGND.t88 VGND.t1476 222.15
R2157 VGND.t1193 VGND.t256 222.15
R2158 VGND.t100 VGND.t122 222.15
R2159 VGND.t563 VGND.t1940 222.15
R2160 VGND.t932 VGND.t2010 222.15
R2161 VGND.t2471 VGND.t1056 222.15
R2162 VGND.t1460 VGND.t930 222.15
R2163 VGND.t665 VGND.t646 222.15
R2164 VGND.t120 VGND.t1756 222.15
R2165 VGND.t882 VGND.t418 222.15
R2166 VGND.t1329 VGND.t118 222.15
R2167 VGND.t1930 VGND.t877 222.15
R2168 VGND.t934 VGND.t1632 222.15
R2169 VGND.t925 VGND.t543 222.15
R2170 VGND.t837 VGND.t86 222.15
R2171 VGND.t347 VGND.t782 222.15
R2172 VGND.t84 VGND.t1317 222.15
R2173 VGND.t1076 VGND.t1983 222.15
R2174 VGND.t200 VGND.t928 222.15
R2175 VGND.t725 VGND.t1192 222.15
R2176 VGND.t926 VGND.t178 222.15
R2177 VGND.t2223 VGND.t1600 222.15
R2178 VGND.t2476 VGND.t269 222.15
R2179 VGND.t2479 VGND.t335 222.15
R2180 VGND.t887 VGND.t116 222.15
R2181 VGND.t1688 VGND.t69 222.15
R2182 VGND.t2383 VGND.t1369 222.15
R2183 VGND.t2222 VGND.t1593 222.15
R2184 VGND.t2373 VGND.t275 222.15
R2185 VGND.t881 VGND.t252 222.15
R2186 VGND.t2391 VGND.t1235 222.15
R2187 VGND.t1062 VGND.t236 222.15
R2188 VGND.t1762 VGND.t1233 222.15
R2189 VGND.t854 VGND.t498 222.15
R2190 VGND.t1017 VGND.t2381 222.15
R2191 VGND.t166 VGND.t783 222.15
R2192 VGND.t2020 VGND.t1573 222.15
R2193 VGND.t2427 VGND.t1387 222.15
R2194 VGND.t1748 VGND.t1571 222.15
R2195 VGND.t2515 VGND.t1579 222.15
R2196 VGND.t94 VGND.t2379 222.15
R2197 VGND.t775 VGND.t268 222.15
R2198 VGND.t1998 VGND.t2377 222.15
R2199 VGND.t1107 VGND.t1210 222.15
R2200 VGND.t638 VGND.t1575 222.15
R2201 VGND.t507 VGND.t222 222.15
R2202 VGND.t1713 VGND.t1231 222.15
R2203 VGND.t2449 VGND.t202 222.15
R2204 VGND.t1648 VGND.t1229 222.15
R2205 VGND.t2421 VGND.t943 222.15
R2206 VGND.t634 VGND.t1569 222.15
R2207 VGND.t1410 VGND.t2483 222.15
R2208 VGND.t831 VGND.t1239 222.15
R2209 VGND.t7 VGND.t765 222.15
R2210 VGND.t1237 VGND.t976 222.15
R2211 VGND.t1565 VGND.t1580 222.15
R2212 VGND.t194 VGND.t2375 222.15
R2213 VGND.t2621 VGND.t880 222.15
R2214 VGND.t515 VGND.t999 222.15
R2215 VGND.t2221 VGND.t1283 222.15
R2216 VGND.t576 VGND.t899 222.15
R2217 VGND.t1173 VGND.t2108 222.15
R2218 VGND.t478 VGND.t960 222.15
R2219 VGND.t1199 VGND.t60 222.15
R2220 VGND.t521 VGND.t104 222.15
R2221 VGND.t154 VGND.t862 222.15
R2222 VGND.t513 VGND.t277 222.15
R2223 VGND.t1262 VGND.t871 222.15
R2224 VGND.t572 VGND.t1535 222.15
R2225 VGND.t2649 VGND.t2431 222.15
R2226 VGND.t570 VGND.t96 222.15
R2227 VGND.t496 VGND.t2242 222.15
R2228 VGND.t511 VGND.t1019 222.15
R2229 VGND.t878 VGND.t1149 222.15
R2230 VGND.t509 VGND.t2026 222.15
R2231 VGND.t647 VGND.t1111 222.15
R2232 VGND.t574 VGND.t1750 222.15
R2233 VGND.t2089 VGND.t533 222.15
R2234 VGND.t519 VGND.t1341 222.15
R2235 VGND.t2387 VGND.t2453 222.15
R2236 VGND.t517 VGND.t1478 222.15
R2237 VGND.t1491 VGND.t144 222.15
R2238 VGND.t1746 VGND.t568 222.15
R2239 VGND.t1501 VGND.t266 222.15
R2240 VGND.t1715 VGND.t482 222.15
R2241 VGND.t37 VGND.t645 222.15
R2242 VGND.t480 VGND.t196 222.15
R2243 VGND.t219 VGND.t1588 222.15
R2244 VGND.t636 VGND.t578 222.15
R2245 VGND.t2647 VGND.t203 222.15
R2246 VGND.t1996 VGND.t755 222.15
R2247 VGND.t2236 VGND.t372 222.15
R2248 VGND.t468 VGND.t1735 222.15
R2249 VGND.t1519 VGND.t703 222.15
R2250 VGND.t1202 VGND.t1331 222.15
R2251 VGND.t397 VGND.t718 222.15
R2252 VGND.t1200 VGND.t885 222.15
R2253 VGND.t49 VGND.t981 222.15
R2254 VGND.t626 VGND.t152 222.15
R2255 VGND.t244 VGND.t1489 222.15
R2256 VGND.t687 VGND.t289 222.15
R2257 VGND.t589 VGND.t73 222.15
R2258 VGND.t966 VGND.t685 222.15
R2259 VGND.t2510 VGND.t1178 222.15
R2260 VGND.t150 VGND.t188 222.15
R2261 VGND.t2076 VGND.t83 222.15
R2262 VGND.t1033 VGND.t148 222.15
R2263 VGND.t1222 VGND.t1994 222.15
R2264 VGND.t689 VGND.t2399 222.15
R2265 VGND.t1123 VGND.t502 222.15
R2266 VGND.t1375 VGND.t759 222.15
R2267 VGND.t1952 VGND.t2505 222.15
R2268 VGND.t757 VGND.t1023 222.15
R2269 VGND.t1129 VGND.t1334 222.15
R2270 VGND.t2393 VGND.t683 222.15
R2271 VGND.t2115 VGND.t205 222.15
R2272 VGND.t1206 VGND.t1039 222.15
R2273 VGND.t1106 VGND.t16 222.15
R2274 VGND.t1204 VGND.t1349 222.15
R2275 VGND.t1128 VGND.t1248 222.15
R2276 VGND.t1614 VGND.t146 222.15
R2277 VGND.t2580 VGND.t20 222.15
R2278 VGND.t742 VGND.t1480 222.15
R2279 VGND.t163 VGND.t2233 222.15
R2280 VGND.t315 VGND.t90 222.15
R2281 VGND.t1216 VGND.t1961 222.15
R2282 VGND.t1339 VGND.t2206 222.15
R2283 VGND.t717 VGND.t2088 222.15
R2284 VGND.t2204 VGND.t198 222.15
R2285 VGND.t1197 VGND.t2231 222.15
R2286 VGND.t740 VGND.t1742 222.15
R2287 VGND.t939 VGND.t241 222.15
R2288 VGND.t311 VGND.t1313 222.15
R2289 VGND.t1915 VGND.t1991 222.15
R2290 VGND.t1053 VGND.t190 222.15
R2291 VGND.t1487 VGND.t2508 222.15
R2292 VGND.t738 VGND.t628 222.15
R2293 VGND.t2078 VGND.t248 222.15
R2294 VGND.t2044 VGND.t291 222.15
R2295 VGND.t1276 VGND.t1220 222.15
R2296 VGND.t313 VGND.t970 222.15
R2297 VGND.t499 VGND.t500 222.15
R2298 VGND.t2202 VGND.t1003 222.15
R2299 VGND.t2224 VGND.t1950 222.15
R2300 VGND.t744 VGND.t281 222.15
R2301 VGND.t691 VGND.t1908 222.15
R2302 VGND.t962 VGND.t1051 222.15
R2303 VGND.t2113 VGND.t2478 222.15
R2304 VGND.t1377 VGND.t1049 222.15
R2305 VGND.t1265 VGND.t1482 222.15
R2306 VGND.t2208 VGND.t1616 222.15
R2307 VGND.t46 VGND.t1245 222.15
R2308 VGND.t2395 VGND.t317 222.15
R2309 VGND.t2571 VGND.t1074 222.15
R2310 VGND.t2181 VGND.t1533 222.15
R2311 VGND.t2085 VGND.t1275 222.15
R2312 VGND.t2171 VGND.t1015 222.15
R2313 VGND.t941 VGND.t1962 222.15
R2314 VGND.t2131 VGND.t1610 222.15
R2315 VGND.t165 VGND.t682 222.15
R2316 VGND.t2129 VGND.t640 222.15
R2317 VGND.t1521 VGND.t1741 222.15
R2318 VGND.t2179 VGND.t92 222.15
R2319 VGND.t1708 VGND.t562 222.15
R2320 VGND.t30 VGND.t1650 222.15
R2321 VGND.t866 VGND.t1055 222.15
R2322 VGND.t28 VGND.t630 222.15
R2323 VGND.t1166 VGND.t2247 222.15
R2324 VGND.t2177 VGND.t1744 222.15
R2325 VGND.t1180 VGND.t417 222.15
R2326 VGND.t2175 VGND.t1315 222.15
R2327 VGND.t240 VGND.t2659 222.15
R2328 VGND.t2169 VGND.t192 222.15
R2329 VGND.t1277 VGND.t540 222.15
R2330 VGND.t2127 VGND.t829 222.15
R2331 VGND.t2388 VGND.t346 222.15
R2332 VGND.t2125 VGND.t907 222.15
R2333 VGND.t373 VGND.t1980 222.15
R2334 VGND.t186 VGND.t26 222.15
R2335 VGND.t724 VGND.t1116 222.15
R2336 VGND.t1005 VGND.t24 222.15
R2337 VGND.t1597 VGND.t1917 222.15
R2338 VGND.t22 VGND.t2397 222.15
R2339 VGND.t2481 VGND.t334 222.15
R2340 VGND.t964 VGND.t2173 222.15
R2341 VGND.t1683 VGND.t719 222.15
R2342 VGND.t1007 VGND.t299 222.15
R2343 VGND.t1495 VGND.t1288 222.15
R2344 VGND.t905 VGND.t2193 222.15
R2345 VGND.t1188 VGND.t467 222.15
R2346 VGND.t968 VGND.t307 222.15
R2347 VGND.t2494 VGND.t2268 222.15
R2348 VGND.t305 VGND.t112 222.15
R2349 VGND.t267 VGND.t537 222.15
R2350 VGND.t297 VGND.t279 222.15
R2351 VGND.t2372 VGND.t1953 222.15
R2352 VGND.t2189 VGND.t1545 222.15
R2353 VGND.t1483 VGND.t2051 222.15
R2354 VGND.t2187 VGND.t102 222.15
R2355 VGND.t853 VGND.t2120 222.15
R2356 VGND.t2199 VGND.t1025 222.15
R2357 VGND.t1294 VGND.t795 222.15
R2358 VGND.t2197 VGND.t2038 222.15
R2359 VGND.t2504 VGND.t777 222.15
R2360 VGND.t2191 VGND.t1764 222.15
R2361 VGND.t220 VGND.t587 222.15
R2362 VGND.t303 VGND.t1351 222.15
R2363 VGND.t1289 VGND.t2669 222.15
R2364 VGND.t2022 VGND.t301 222.15
R2365 VGND.t2416 VGND.t662 222.15
R2366 VGND.t1758 VGND.t2185 222.15
R2367 VGND.t2159 VGND.t2232 222.15
R2368 VGND.t1723 VGND.t2183 222.15
R2369 VGND.t1263 VGND.t938 222.15
R2370 VGND.t1634 VGND.t309 222.15
R2371 VGND.t294 VGND.t1103 222.15
R2372 VGND.t1462 VGND.t2195 222.15
R2373 VGND.t2341 VGND.t221 222.15
R2374 VGND.t423 VGND.t1531 222.15
R2375 VGND.t371 VGND.t1595 222.15
R2376 VGND.t913 VGND.t1620 222.15
R2377 VGND.t663 VGND.t254 222.15
R2378 VGND.t431 VGND.t1606 222.15
R2379 VGND.t1127 VGND.t1064 222.15
R2380 VGND.t632 VGND.t429 222.15
R2381 VGND.t860 VGND.t1105 222.15
R2382 VGND.t921 VGND.t1359 222.15
R2383 VGND.t1212 VGND.t168 222.15
R2384 VGND.t1646 VGND.t909 222.15
R2385 VGND.t2429 VGND.t1939 222.15
R2386 VGND.t2434 VGND.t624 222.15
R2387 VGND.t2485 VGND.t2517 222.15
R2388 VGND.t1733 VGND.t919 222.15
R2389 VGND.t1143 VGND.t2168 222.15
R2390 VGND.t917 VGND.t1309 222.15
R2391 VGND.t2080 VGND.t1224 222.15
R2392 VGND.t911 VGND.t184 222.15
R2393 VGND.t1711 VGND.t531 222.15
R2394 VGND.t825 VGND.t427 222.15
R2395 VGND.t2451 VGND.t2102 222.15
R2396 VGND.t903 VGND.t425 222.15
R2397 VGND.t142 VGND.t1075 222.15
R2398 VGND.t2432 VGND.t182 222.15
R2399 VGND.t174 VGND.t1412 222.15
R2400 VGND.t415 VGND.t995 222.15
R2401 VGND.t2098 VGND.t35 222.15
R2402 VGND.t433 VGND.t2389 222.15
R2403 VGND.t770 VGND.t1586 222.15
R2404 VGND.t958 VGND.t915 222.15
R2405 VGND.t2641 VGND.t414 222.15
R2406 VGND.t1622 VGND.t2500 222.15
R2407 VGND.t1494 VGND.t644 222.15
R2408 VGND.t2548 VGND.t1367 222.15
R2409 VGND.t1603 VGND.t1187 222.15
R2410 VGND.t108 VGND.t807 222.15
R2411 VGND.t2497 VGND.t1223 222.15
R2412 VGND.t805 VGND.t2018 222.15
R2413 VGND.t53 VGND.t536 222.15
R2414 VGND.t1537 VGND.t1563 222.15
R2415 VGND.t2071 VGND.t2502 222.15
R2416 VGND.t2544 VGND.t1727 222.15
R2417 VGND.t2386 VGND.t2050 222.15
R2418 VGND.t2008 VGND.t2542 222.15
R2419 VGND.t594 VGND.t2385 222.15
R2420 VGND.t1561 VGND.t2030 222.15
R2421 VGND.t1124 VGND.t794 222.15
R2422 VGND.t622 VGND.t1559 222.15
R2423 VGND.t776 VGND.t249 222.15
R2424 VGND.t2546 VGND.t1327 222.15
R2425 VGND.t1500 VGND.t584 222.15
R2426 VGND.t1640 VGND.t803 222.15
R2427 VGND.t1102 VGND.t235 222.15
R2428 VGND.t833 VGND.t801 222.15
R2429 VGND.t2413 VGND.t160 222.15
R2430 VGND.t1319 VGND.t2540 222.15
R2431 VGND.t2158 VGND.t1296 222.15
R2432 VGND.t897 VGND.t2538 222.15
R2433 VGND.t1259 VGND.t748 222.15
R2434 VGND.t809 VGND.t1037 222.15
R2435 VGND.t1130 VGND.t293 222.15
R2436 VGND.t817 VGND.t2550 222.15
R2437 VGND.t2338 VGND.t2437 222.15
R2438 VGND.t849 VGND.t2403 222.15
R2439 VGND.t876 VGND.t1272 222.15
R2440 VGND.t997 VGND.t839 222.15
R2441 VGND.t2650 VGND.t1493 222.15
R2442 VGND.t1566 VGND.t1031 222.15
R2443 VGND.t2503 VGND.t1160 222.15
R2444 VGND.t2273 VGND.t1604 222.15
R2445 VGND.t1938 VGND.t261 222.15
R2446 VGND.t847 VGND.t1371 222.15
R2447 VGND.t54 VGND.t696 222.15
R2448 VGND.t1514 VGND.t1355 222.15
R2449 VGND.t761 VGND.t1057 222.15
R2450 VGND.t1512 VGND.t2032 222.15
R2451 VGND.t175 VGND.t670 222.15
R2452 VGND.t845 VGND.t1539 222.15
R2453 VGND.t2370 VGND.t1117 222.15
R2454 VGND.t843 VGND.t1731 222.15
R2455 VGND.t71 VGND.t1935 222.15
R2456 VGND.t2012 VGND.t1516 222.15
R2457 VGND.t544 VGND.t1916 222.15
R2458 VGND.t1468 VGND.t2271 222.15
R2459 VGND.t348 VGND.t1486 222.15
R2460 VGND.t2269 VGND.t1719 222.15
R2461 VGND.t2488 VGND.t1984 222.15
R2462 VGND.t1510 VGND.t2000 222.15
R2463 VGND.t19 VGND.t730 222.15
R2464 VGND.t1642 VGND.t1508 222.15
R2465 VGND.t1601 VGND.t1578 222.15
R2466 VGND.t819 VGND.t1506 222.15
R2467 VGND.t340 VGND.t70 222.15
R2468 VGND.t1321 VGND.t841 222.15
R2469 VGND.t1703 VGND.t1073 222.15
R2470 VGND.t134 VGND.t974 222.15
R2471 VGND.t1179 VGND.t2234 222.15
R2472 VGND.t1945 VGND.t827 222.15
R2473 VGND.t1141 VGND.t1960 222.15
R2474 VGND.t448 VGND.t287 222.15
R2475 VGND.t32 VGND.t716 222.15
R2476 VGND.t1043 VGND.t446 222.15
R2477 VGND.t2230 VGND.t21 222.15
R2478 VGND.t1001 VGND.t132 222.15
R2479 VGND.t242 VGND.t2661 222.15
R2480 VGND.t1618 VGND.t1086 222.15
R2481 VGND.t1992 VGND.t48 222.15
R2482 VGND.t1541 VGND.t1084 222.15
R2483 VGND.t2507 VGND.t2486 222.15
R2484 VGND.t1373 VGND.t130 222.15
R2485 VGND.t247 VGND.t159 222.15
R2486 VGND.t1357 VGND.t128 222.15
R2487 VGND.t1219 VGND.t2090 222.15
R2488 VGND.t1943 VGND.t2034 222.15
R2489 VGND.t1485 VGND.t588 222.15
R2490 VGND.t444 VGND.t1523 222.15
R2491 VGND.t1602 VGND.t1949 222.15
R2492 VGND.t136 VGND.t1345 222.15
R2493 VGND.t1182 VGND.t1907 222.15
R2494 VGND.t1082 VGND.t2024 222.15
R2495 VGND.t1198 VGND.t2112 222.15
R2496 VGND.t1470 VGND.t1080 222.15
R2497 VGND.t1264 VGND.t47 222.15
R2498 VGND.t1078 VGND.t1323 222.15
R2499 VGND.t1131 VGND.t1246 222.15
R2500 VGND.t2002 VGND.t1947 222.15
R2501 VGND.t2570 VGND.t923 222.15
R2502 VGND.t1474 VGND.t2609 222.15
R2503 VGND.t2668 VGND.t370 222.15
R2504 VGND.t2339 VGND.t1343 222.15
R2505 VGND.t1520 VGND.t2658 222.15
R2506 VGND.t1693 VGND.t2006 222.15
R2507 VGND.t1293 VGND.t2493 222.15
R2508 VGND.t1671 VGND.t180 222.15
R2509 VGND.t746 VGND.t265 222.15
R2510 VGND.t2598 VGND.t1717 222.15
R2511 VGND.t865 VGND.t2212 222.15
R2512 VGND.t2320 VGND.t895 222.15
R2513 VGND.t1914 VGND.t754 222.15
R2514 VGND.t2309 VGND.t1011 222.15
R2515 VGND.t126 VGND.t678 222.15
R2516 VGND.t2594 VGND.t835 222.15
R2517 VGND.t2436 VGND.t2 222.15
R2518 VGND.t2576 VGND.t273 222.15
R2519 VGND.t1937 VGND.t712 222.15
R2520 VGND.t2322 VGND.t1385 222.15
R2521 VGND.t1390 VGND.t789 222.15
R2522 VGND.t1658 VGND.t991 222.15
R2523 VGND.t1218 VGND.t1096 222.15
R2524 VGND.t2642 VGND.t2407 222.15
R2525 VGND.t1152 VGND.t1979 222.15
R2526 VGND.t2304 VGND.t1381 222.15
R2527 VGND.t1290 VGND.t2153 222.15
R2528 VGND.t2291 VGND.t1365 222.15
R2529 VGND.t161 VGND.t664 222.15
R2530 VGND.t1699 VGND.t1608 222.15
R2531 VGND.t1209 VGND.t323 222.15
R2532 VGND.t1045 VGND.t2366 222.15
R2533 VGND.t2295 VGND.t1490 222.15
R2534 VGND.n2346 VGND.n3 218.73
R2535 VGND.n489 VGND.n487 214.365
R2536 VGND.n489 VGND.n488 214.365
R2537 VGND.n479 VGND.n477 214.365
R2538 VGND.n479 VGND.n478 214.365
R2539 VGND.n497 VGND.n495 214.365
R2540 VGND.n497 VGND.n496 214.365
R2541 VGND.n2270 VGND.n2268 214.365
R2542 VGND.n2270 VGND.n2269 214.365
R2543 VGND.n2260 VGND.n2258 214.365
R2544 VGND.n2260 VGND.n2259 214.365
R2545 VGND.n2278 VGND.n2276 214.365
R2546 VGND.n2278 VGND.n2277 214.365
R2547 VGND.n525 VGND.n523 214.365
R2548 VGND.n525 VGND.n524 214.365
R2549 VGND.n515 VGND.n513 214.365
R2550 VGND.n515 VGND.n514 214.365
R2551 VGND.n533 VGND.n531 214.365
R2552 VGND.n533 VGND.n532 214.365
R2553 VGND.n2191 VGND.n2190 214.365
R2554 VGND.n1140 VGND.n1139 213.613
R2555 VGND.n1142 VGND.n1141 213.613
R2556 VGND.n1112 VGND.n1110 213.613
R2557 VGND.n1112 VGND.n1111 213.613
R2558 VGND.n1115 VGND.n1113 213.613
R2559 VGND.n1115 VGND.n1114 213.613
R2560 VGND.n2236 VGND.n2229 213.613
R2561 VGND.n2236 VGND.n2230 213.613
R2562 VGND.n2234 VGND.n2231 213.613
R2563 VGND.n2234 VGND.n2233 213.613
R2564 VGND.n1374 VGND.n1367 213.613
R2565 VGND.n1374 VGND.n1368 213.613
R2566 VGND.n1372 VGND.n1369 213.613
R2567 VGND.n1372 VGND.n1371 213.613
R2568 VGND.n1154 VGND.t1297 211.359
R2569 VGND.n179 VGND.n175 207.965
R2570 VGND.n179 VGND.n176 207.965
R2571 VGND.n173 VGND.n171 207.965
R2572 VGND.n173 VGND.n172 207.965
R2573 VGND.n186 VGND.n169 207.965
R2574 VGND.n186 VGND.n170 207.965
R2575 VGND.n98 VGND.n97 207.965
R2576 VGND.n110 VGND.n95 207.965
R2577 VGND.n102 VGND.n100 207.965
R2578 VGND.n80 VGND.n76 207.965
R2579 VGND.n80 VGND.n77 207.965
R2580 VGND.n74 VGND.n72 207.965
R2581 VGND.n74 VGND.n73 207.965
R2582 VGND.n87 VGND.n70 207.965
R2583 VGND.n87 VGND.n71 207.965
R2584 VGND.n148 VGND.n144 207.965
R2585 VGND.n148 VGND.n145 207.965
R2586 VGND.n142 VGND.n140 207.965
R2587 VGND.n142 VGND.n141 207.965
R2588 VGND.n155 VGND.n138 207.965
R2589 VGND.n155 VGND.n139 207.965
R2590 VGND.n2188 VGND.n2187 207.965
R2591 VGND.n2205 VGND.n2185 207.965
R2592 VGND.n2981 VGND.n2979 207.213
R2593 VGND.n2981 VGND.n2980 207.213
R2594 VGND.n2985 VGND.n2976 207.213
R2595 VGND.n2985 VGND.n2977 207.213
R2596 VGND.n18 VGND.n16 207.213
R2597 VGND.n18 VGND.n17 207.213
R2598 VGND.n22 VGND.n14 207.213
R2599 VGND.n22 VGND.n15 207.213
R2600 VGND.n2951 VGND.n2950 207.213
R2601 VGND.n2955 VGND.n2949 207.213
R2602 VGND.n44 VGND.n42 207.213
R2603 VGND.n44 VGND.n43 207.213
R2604 VGND.n48 VGND.n40 207.213
R2605 VGND.n48 VGND.n41 207.213
R2606 VGND.n109 VGND.n96 207.213
R2607 VGND.n2204 VGND.n2186 207.213
R2608 VGND.t1824 VGND.t2364 203.242
R2609 VGND.t2287 VGND.t1773 203.242
R2610 VGND.t1779 VGND.t2637 203.242
R2611 VGND.t2613 VGND.t1797 203.242
R2612 VGND.t1872 VGND.t2285 203.242
R2613 VGND.t1706 VGND.t1878 203.242
R2614 VGND.t1800 VGND.t1684 203.242
R2615 VGND.t2352 VGND.t1842 203.242
R2616 VGND.t1851 VGND.t2332 203.242
R2617 VGND.t1679 VGND.t1890 203.242
R2618 VGND.t1806 VGND.t2596 203.242
R2619 VGND.t2585 VGND.t1854 203.242
R2620 VGND.t1893 VGND.t2307 203.242
R2621 VGND.t1669 VGND.t1902 203.242
R2622 VGND.t1818 VGND.t2574 203.242
R2623 VGND.t2318 VGND.t1860 203.242
R2624 VGND VGND.n332 194.419
R2625 VGND VGND.n356 194.419
R2626 VGND VGND.n363 194.419
R2627 VGND VGND.n366 194.419
R2628 VGND VGND.n374 194.419
R2629 VGND VGND.n377 194.419
R2630 VGND VGND.n385 194.419
R2631 VGND VGND.n324 194.419
R2632 VGND VGND.n313 194.419
R2633 VGND VGND.n308 194.419
R2634 VGND VGND.n310 194.419
R2635 VGND VGND.n2729 194.419
R2636 VGND VGND.n292 194.419
R2637 VGND VGND.n295 194.419
R2638 VGND VGND.n202 194.419
R2639 VGND.n887 VGND.n886 194.391
R2640 VGND.n1332 VGND.n889 194.391
R2641 VGND.n895 VGND.n893 194.391
R2642 VGND.n931 VGND.n930 194.391
R2643 VGND.n936 VGND.n935 194.391
R2644 VGND.n941 VGND.n940 194.391
R2645 VGND.n946 VGND.n945 194.391
R2646 VGND.n951 VGND.n950 194.391
R2647 VGND.n956 VGND.n955 194.391
R2648 VGND.n961 VGND.n960 194.391
R2649 VGND.n966 VGND.n965 194.391
R2650 VGND.n971 VGND.n970 194.391
R2651 VGND.n976 VGND.n975 194.391
R2652 VGND.n981 VGND.n980 194.391
R2653 VGND.n986 VGND.n985 194.391
R2654 VGND.n1281 VGND.n996 194.391
R2655 VGND.n1274 VGND.n1273 194.391
R2656 VGND.n1231 VGND.n1230 194.391
R2657 VGND.n1236 VGND.n1229 194.391
R2658 VGND.n1227 VGND.n1226 194.391
R2659 VGND.n1243 VGND.n1224 194.391
R2660 VGND.n1222 VGND.n1221 194.391
R2661 VGND.n1217 VGND.n1216 194.391
R2662 VGND.n1211 VGND.n1002 194.391
R2663 VGND.n1204 VGND.n1203 194.391
R2664 VGND.n1008 VGND.n1007 194.391
R2665 VGND.n1185 VGND.n1184 194.391
R2666 VGND.n1179 VGND.n1010 194.391
R2667 VGND.n1172 VGND.n1171 194.391
R2668 VGND.n1169 VGND.n1012 194.391
R2669 VGND.n330 VGND.n329 194.391
R2670 VGND.n396 VGND.n395 194.391
R2671 VGND.n2638 VGND.n2637 194.391
R2672 VGND.n2643 VGND.n2642 194.391
R2673 VGND.n2648 VGND.n2647 194.391
R2674 VGND.n2653 VGND.n2652 194.391
R2675 VGND.n2658 VGND.n2657 194.391
R2676 VGND.n2663 VGND.n2662 194.391
R2677 VGND.n2668 VGND.n2667 194.391
R2678 VGND.n393 VGND.n392 194.391
R2679 VGND.n2714 VGND.n2713 194.391
R2680 VGND.n319 VGND.n318 194.391
R2681 VGND.n2747 VGND.n2746 194.391
R2682 VGND.n303 VGND.n302 194.391
R2683 VGND.n2752 VGND.n2751 194.391
R2684 VGND.n2787 VGND.n2786 194.391
R2685 VGND.n286 VGND.n285 194.391
R2686 VGND.n400 VGND.n399 194.391
R2687 VGND.n2342 VGND.n2341 194.391
R2688 VGND.n2337 VGND.n2336 194.391
R2689 VGND.n2332 VGND.n2331 194.391
R2690 VGND.n2327 VGND.n2326 194.391
R2691 VGND.n2322 VGND.n2321 194.391
R2692 VGND.n2317 VGND.n2316 194.391
R2693 VGND.n2312 VGND.n2311 194.391
R2694 VGND.n2307 VGND.n2306 194.391
R2695 VGND.n2302 VGND.n2301 194.391
R2696 VGND.n2297 VGND.n2296 194.391
R2697 VGND.n2292 VGND.n2291 194.391
R2698 VGND.n2287 VGND.n2286 194.391
R2699 VGND.n414 VGND.n413 194.391
R2700 VGND.n2540 VGND.n2539 194.391
R2701 VGND.n2535 VGND.n416 194.391
R2702 VGND.n469 VGND.n468 194.391
R2703 VGND.n471 VGND.n470 194.391
R2704 VGND.n2376 VGND.n2375 194.391
R2705 VGND.n459 VGND.n458 194.391
R2706 VGND.n2402 VGND.n2401 194.391
R2707 VGND.n451 VGND.n450 194.391
R2708 VGND.n2428 VGND.n2427 194.391
R2709 VGND.n443 VGND.n442 194.391
R2710 VGND.n2454 VGND.n2453 194.391
R2711 VGND.n435 VGND.n434 194.391
R2712 VGND.n2480 VGND.n2479 194.391
R2713 VGND.n427 VGND.n426 194.391
R2714 VGND.n2511 VGND.n2510 194.391
R2715 VGND.n2516 VGND.n2515 194.391
R2716 VGND.n2521 VGND.n2520 194.391
R2717 VGND.n2528 VGND.n418 194.391
R2718 VGND.n466 VGND.n465 194.391
R2719 VGND.n2363 VGND.n2362 194.391
R2720 VGND.n463 VGND.n462 194.391
R2721 VGND.n2389 VGND.n2388 194.391
R2722 VGND.n455 VGND.n454 194.391
R2723 VGND.n2415 VGND.n2414 194.391
R2724 VGND.n447 VGND.n446 194.391
R2725 VGND.n2441 VGND.n2440 194.391
R2726 VGND.n439 VGND.n438 194.391
R2727 VGND.n2467 VGND.n2466 194.391
R2728 VGND.n431 VGND.n430 194.391
R2729 VGND.n2493 VGND.n2492 194.391
R2730 VGND.n423 VGND.n422 194.391
R2731 VGND.n2498 VGND.n2497 194.391
R2732 VGND.n2809 VGND.n2808 194.391
R2733 VGND.n2816 VGND.n276 194.391
R2734 VGND.n625 VGND.n624 194.391
R2735 VGND.n1910 VGND.n1909 194.391
R2736 VGND.n622 VGND.n621 194.391
R2737 VGND.n1921 VGND.n1920 194.391
R2738 VGND.n619 VGND.n618 194.391
R2739 VGND.n1932 VGND.n1931 194.391
R2740 VGND.n616 VGND.n615 194.391
R2741 VGND.n1943 VGND.n1942 194.391
R2742 VGND.n613 VGND.n612 194.391
R2743 VGND.n1954 VGND.n1953 194.391
R2744 VGND.n610 VGND.n609 194.391
R2745 VGND.n1965 VGND.n1964 194.391
R2746 VGND.n607 VGND.n606 194.391
R2747 VGND.n1976 VGND.n1975 194.391
R2748 VGND.n1981 VGND.n1980 194.391
R2749 VGND.n1988 VGND.n605 194.391
R2750 VGND.n590 VGND.n589 194.391
R2751 VGND.n596 VGND.n595 194.391
R2752 VGND.n593 VGND.n592 194.391
R2753 VGND.n2055 VGND.n2054 194.391
R2754 VGND.n2050 VGND.n2049 194.391
R2755 VGND.n2045 VGND.n2044 194.391
R2756 VGND.n2040 VGND.n2039 194.391
R2757 VGND.n2035 VGND.n2034 194.391
R2758 VGND.n2030 VGND.n2029 194.391
R2759 VGND.n2025 VGND.n2024 194.391
R2760 VGND.n2020 VGND.n2019 194.391
R2761 VGND.n2015 VGND.n2014 194.391
R2762 VGND.n2010 VGND.n2009 194.391
R2763 VGND.n2005 VGND.n2004 194.391
R2764 VGND.n2000 VGND.n600 194.391
R2765 VGND.n1995 VGND.n1993 194.391
R2766 VGND.n587 VGND.n586 194.391
R2767 VGND.n2069 VGND.n2068 194.391
R2768 VGND.n2074 VGND.n2073 194.391
R2769 VGND.n2079 VGND.n2078 194.391
R2770 VGND.n2084 VGND.n2083 194.391
R2771 VGND.n2089 VGND.n2088 194.391
R2772 VGND.n2094 VGND.n2093 194.391
R2773 VGND.n2099 VGND.n2098 194.391
R2774 VGND.n2104 VGND.n2103 194.391
R2775 VGND.n2109 VGND.n2108 194.391
R2776 VGND.n2114 VGND.n2113 194.391
R2777 VGND.n2119 VGND.n2118 194.391
R2778 VGND.n584 VGND.n583 194.391
R2779 VGND.n2124 VGND.n2123 194.391
R2780 VGND.n2834 VGND.n2833 194.391
R2781 VGND.n2841 VGND.n264 194.391
R2782 VGND.n547 VGND.n546 194.391
R2783 VGND.n2176 VGND.n549 194.391
R2784 VGND.n1757 VGND.n1755 194.391
R2785 VGND.n1761 VGND.n1760 194.391
R2786 VGND.n1752 VGND.n1751 194.391
R2787 VGND.n1772 VGND.n1771 194.391
R2788 VGND.n1749 VGND.n1748 194.391
R2789 VGND.n1783 VGND.n1782 194.391
R2790 VGND.n1746 VGND.n1745 194.391
R2791 VGND.n1794 VGND.n1793 194.391
R2792 VGND.n1743 VGND.n1742 194.391
R2793 VGND.n1805 VGND.n1804 194.391
R2794 VGND.n1740 VGND.n1739 194.391
R2795 VGND.n1816 VGND.n1815 194.391
R2796 VGND.n1821 VGND.n1820 194.391
R2797 VGND.n1828 VGND.n1738 194.391
R2798 VGND.n628 VGND.n627 194.391
R2799 VGND.n1678 VGND.n1677 194.391
R2800 VGND.n1675 VGND.n1674 194.391
R2801 VGND.n1689 VGND.n1688 194.391
R2802 VGND.n1694 VGND.n1693 194.391
R2803 VGND.n1699 VGND.n1698 194.391
R2804 VGND.n1704 VGND.n1703 194.391
R2805 VGND.n1709 VGND.n1708 194.391
R2806 VGND.n1714 VGND.n1713 194.391
R2807 VGND.n1719 VGND.n1718 194.391
R2808 VGND.n1724 VGND.n1723 194.391
R2809 VGND.n1729 VGND.n1728 194.391
R2810 VGND.n1672 VGND.n1671 194.391
R2811 VGND.n1845 VGND.n1844 194.391
R2812 VGND.n1840 VGND.n1733 194.391
R2813 VGND.n1835 VGND.n1833 194.391
R2814 VGND.n632 VGND.n631 194.391
R2815 VGND.n669 VGND.n668 194.391
R2816 VGND.n674 VGND.n673 194.391
R2817 VGND.n679 VGND.n678 194.391
R2818 VGND.n684 VGND.n683 194.391
R2819 VGND.n689 VGND.n688 194.391
R2820 VGND.n694 VGND.n693 194.391
R2821 VGND.n699 VGND.n698 194.391
R2822 VGND.n704 VGND.n703 194.391
R2823 VGND.n709 VGND.n708 194.391
R2824 VGND.n714 VGND.n713 194.391
R2825 VGND.n719 VGND.n718 194.391
R2826 VGND.n666 VGND.n665 194.391
R2827 VGND.n724 VGND.n723 194.391
R2828 VGND.n2859 VGND.n2858 194.391
R2829 VGND.n2866 VGND.n252 194.391
R2830 VGND.n879 VGND.n878 194.391
R2831 VGND.n1352 VGND.n1351 194.391
R2832 VGND.n874 VGND.n873 194.391
R2833 VGND.n869 VGND.n807 194.391
R2834 VGND.n811 VGND.n809 194.391
R2835 VGND.n823 VGND.n822 194.391
R2836 VGND.n828 VGND.n827 194.391
R2837 VGND.n833 VGND.n832 194.391
R2838 VGND.n838 VGND.n837 194.391
R2839 VGND.n843 VGND.n842 194.391
R2840 VGND.n848 VGND.n847 194.391
R2841 VGND.n819 VGND.n818 194.391
R2842 VGND.n853 VGND.n852 194.391
R2843 VGND.n734 VGND.n733 194.391
R2844 VGND.n1661 VGND.n1660 194.391
R2845 VGND.n1656 VGND.n736 194.391
R2846 VGND.n800 VGND.n799 194.391
R2847 VGND.n1390 VGND.n1389 194.391
R2848 VGND.n1395 VGND.n1394 194.391
R2849 VGND.n804 VGND.n803 194.391
R2850 VGND.n1490 VGND.n1489 194.391
R2851 VGND.n776 VGND.n775 194.391
R2852 VGND.n1516 VGND.n1515 194.391
R2853 VGND.n768 VGND.n767 194.391
R2854 VGND.n1542 VGND.n1541 194.391
R2855 VGND.n1547 VGND.n1546 194.391
R2856 VGND.n760 VGND.n759 194.391
R2857 VGND.n1552 VGND.n1551 194.391
R2858 VGND.n1632 VGND.n1631 194.391
R2859 VGND.n1637 VGND.n1636 194.391
R2860 VGND.n1642 VGND.n1641 194.391
R2861 VGND.n1649 VGND.n739 194.391
R2862 VGND.n797 VGND.n796 194.391
R2863 VGND.n1410 VGND.n1409 194.391
R2864 VGND.n794 VGND.n793 194.391
R2865 VGND.n1477 VGND.n1476 194.391
R2866 VGND.n780 VGND.n779 194.391
R2867 VGND.n1503 VGND.n1502 194.391
R2868 VGND.n772 VGND.n771 194.391
R2869 VGND.n1529 VGND.n1528 194.391
R2870 VGND.n764 VGND.n763 194.391
R2871 VGND.n1566 VGND.n1565 194.391
R2872 VGND.n755 VGND.n754 194.391
R2873 VGND.n1581 VGND.n1580 194.391
R2874 VGND.n1576 VGND.n1575 194.391
R2875 VGND.n1571 VGND.n1570 194.391
R2876 VGND.n2884 VGND.n2883 194.391
R2877 VGND.n2891 VGND.n239 194.391
R2878 VGND.n882 VGND.n881 194.391
R2879 VGND.n884 VGND.n883 194.391
R2880 VGND.n1423 VGND.n1422 194.391
R2881 VGND.n1428 VGND.n1427 194.391
R2882 VGND.n1433 VGND.n1432 194.391
R2883 VGND.n1438 VGND.n1437 194.391
R2884 VGND.n1443 VGND.n1442 194.391
R2885 VGND.n1448 VGND.n1447 194.391
R2886 VGND.n1453 VGND.n1452 194.391
R2887 VGND.n790 VGND.n789 194.391
R2888 VGND.n1458 VGND.n1457 194.391
R2889 VGND.n1595 VGND.n1594 194.391
R2890 VGND.n1600 VGND.n1599 194.391
R2891 VGND.n749 VGND.n748 194.391
R2892 VGND.n1613 VGND.n1612 194.391
R2893 VGND.n1608 VGND.n1604 194.391
R2894 VGND.n1024 VGND.n1023 194.391
R2895 VGND.n1031 VGND.n1030 194.391
R2896 VGND.n1036 VGND.n1035 194.391
R2897 VGND.n1028 VGND.n1027 194.391
R2898 VGND.n1094 VGND.n1093 194.391
R2899 VGND.n1089 VGND.n1088 194.391
R2900 VGND.n1084 VGND.n1083 194.391
R2901 VGND.n1079 VGND.n1078 194.391
R2902 VGND.n1074 VGND.n1073 194.391
R2903 VGND.n1069 VGND.n1040 194.391
R2904 VGND.n1044 VGND.n1042 194.391
R2905 VGND.n1052 VGND.n1051 194.391
R2906 VGND.n1057 VGND.n1056 194.391
R2907 VGND.n1048 VGND.n1047 194.391
R2908 VGND.n2904 VGND.n2903 194.391
R2909 VGND.n2911 VGND.n227 194.391
R2910 VGND.n1014 VGND.n1013 194.391
R2911 VGND.n927 VGND.n926 194.391
R2912 VGND.n2606 VGND.n2605 161.308
R2913 VGND.n2603 VGND.n2602 161.308
R2914 VGND.n2600 VGND.n2599 161.308
R2915 VGND.n2597 VGND.n2596 161.308
R2916 VGND.n2594 VGND.n2593 161.308
R2917 VGND.n2591 VGND.n2590 161.308
R2918 VGND.n2588 VGND.n2587 161.308
R2919 VGND.n2585 VGND.n2584 161.308
R2920 VGND.n2582 VGND.n2581 161.308
R2921 VGND.n2579 VGND.n2578 161.308
R2922 VGND.n2576 VGND.n2575 161.308
R2923 VGND.n2573 VGND.n2572 161.308
R2924 VGND.n2570 VGND.n2569 161.308
R2925 VGND.n2567 VGND.n2566 161.308
R2926 VGND.n2564 VGND.n2563 161.308
R2927 VGND.n2605 VGND.t2696 159.978
R2928 VGND.n2602 VGND.t2699 159.978
R2929 VGND.n2599 VGND.t2694 159.978
R2930 VGND.n2596 VGND.t2689 159.978
R2931 VGND.n2593 VGND.t2695 159.978
R2932 VGND.n2590 VGND.t2702 159.978
R2933 VGND.n2587 VGND.t2698 159.978
R2934 VGND.n2584 VGND.t2692 159.978
R2935 VGND.n2581 VGND.t2688 159.978
R2936 VGND.n2578 VGND.t2690 159.978
R2937 VGND.n2575 VGND.t2701 159.978
R2938 VGND.n2572 VGND.t2693 159.978
R2939 VGND.n2569 VGND.t2700 159.978
R2940 VGND.n2566 VGND.t2697 159.978
R2941 VGND.n2563 VGND.t2703 159.978
R2942 VGND.n123 VGND.t329 159.315
R2943 VGND.n2216 VGND.t2084 159.315
R2944 VGND.n1132 VGND.t2249 158.361
R2945 VGND.n2999 VGND.t2101 158.361
R2946 VGND.n121 VGND.t327 157.291
R2947 VGND.n544 VGND.t2082 157.291
R2948 VGND.n68 VGND.t1921 156.915
R2949 VGND.n506 VGND.t1140 156.915
R2950 VGND.n68 VGND.t1922 156.915
R2951 VGND.n506 VGND.t1138 156.915
R2952 VGND.n36 VGND.t239 154.131
R2953 VGND.n123 VGND.t1196 154.131
R2954 VGND.n128 VGND.t58 154.131
R2955 VGND.n128 VGND.t1191 154.131
R2956 VGND.n508 VGND.t749 154.131
R2957 VGND.n508 VGND.t115 154.131
R2958 VGND.n2216 VGND.t2499 154.131
R2959 VGND.n541 VGND.t1161 154.131
R2960 VGND.n3005 VGND.t763 153.631
R2961 VGND.n60 VGND.t769 153.631
R2962 VGND.n160 VGND.t1919 153.631
R2963 VGND.n2255 VGND.t1137 153.631
R2964 VGND.n2222 VGND.t1168 153.631
R2965 VGND.n1360 VGND.t1577 153.631
R2966 VGND.n59 VGND.t1170 152.757
R2967 VGND.n2221 VGND.t990 152.757
R2968 VGND.n92 VGND.t1926 152.381
R2969 VGND.n2211 VGND.t1134 152.381
R2970 VGND.n2181 VGND.n2180 152.174
R2971 VGND.n167 VGND.t1929 150.922
R2972 VGND.n167 VGND.t1924 150.922
R2973 VGND.n475 VGND.t1139 150.922
R2974 VGND.n475 VGND.t1132 150.922
R2975 VGND.n166 VGND.t1392 150.922
R2976 VGND.n67 VGND.t210 150.922
R2977 VGND.n135 VGND.t653 150.922
R2978 VGND.n474 VGND.t68 150.922
R2979 VGND.n2253 VGND.t2472 150.922
R2980 VGND.n505 VGND.t1174 150.922
R2981 VGND.n166 VGND.t1912 150.922
R2982 VGND.n67 VGND.t1163 150.922
R2983 VGND.n135 VGND.t870 150.922
R2984 VGND.n474 VGND.t1522 150.922
R2985 VGND.n2253 VGND.t2201 150.922
R2986 VGND.n505 VGND.t564 150.922
R2987 VGND.n3004 VGND.t320 147.411
R2988 VGND.n159 VGND.t1928 147.411
R2989 VGND.n2254 VGND.t1135 147.411
R2990 VGND.n1359 VGND.t331 147.411
R2991 VGND.n115 VGND.t1550 146.964
R2992 VGND.n545 VGND.t1306 146.964
R2993 VGND.n2605 VGND.t1808 143.911
R2994 VGND.n2602 VGND.t1883 143.911
R2995 VGND.n2599 VGND.t1790 143.911
R2996 VGND.n2596 VGND.t1832 143.911
R2997 VGND.n2593 VGND.t1904 143.911
R2998 VGND.n2590 VGND.t1811 143.911
R2999 VGND.n2587 VGND.t1784 143.911
R3000 VGND.n2584 VGND.t1826 143.911
R3001 VGND.n2581 VGND.t1838 143.911
R3002 VGND.n2578 VGND.t1766 143.911
R3003 VGND.n2575 VGND.t1862 143.911
R3004 VGND.n2572 VGND.t1793 143.911
R3005 VGND.n2569 VGND.t1865 143.911
R3006 VGND.n2566 VGND.t1895 143.911
R3007 VGND.n2563 VGND.t1835 143.911
R3008 VGND.n1388 VGND.n806 143.478
R3009 VGND VGND.t464 142.089
R3010 VGND.n1021 VGND.t1823 119.309
R3011 VGND.n994 VGND.t1859 119.309
R3012 VGND.n2630 VGND.t1820 119.309
R3013 VGND.n204 VGND.t1856 119.309
R3014 VGND.n334 VGND.t1769 119.309
R3015 VGND.n2626 VGND.t1775 119.309
R3016 VGND.n2623 VGND.t1781 119.309
R3017 VGND.n2620 VGND.t1868 119.309
R3018 VGND.n2617 VGND.t1874 119.309
R3019 VGND.n2614 VGND.t1787 119.309
R3020 VGND.n2611 VGND.t1829 119.309
R3021 VGND.n322 VGND.t1844 119.309
R3022 VGND.n315 VGND.t1880 119.309
R3023 VGND.n306 VGND.t1802 119.309
R3024 VGND.n299 VGND.t1847 119.309
R3025 VGND.n2765 VGND.t1886 119.309
R3026 VGND.n290 VGND.t1898 119.309
R3027 VGND.n297 VGND.t1814 119.309
R3028 VGND.n1018 VGND.t1772 119.309
R3029 VGND.n1015 VGND.t1778 119.309
R3030 VGND.n1180 VGND.t1796 119.309
R3031 VGND.n1006 VGND.t1871 119.309
R3032 VGND.n1004 VGND.t1877 119.309
R3033 VGND.n1195 VGND.t1799 119.309
R3034 VGND.n1212 VGND.t1841 119.309
R3035 VGND.n1000 VGND.t1850 119.309
R3036 VGND.n1253 VGND.t1889 119.309
R3037 VGND.n1256 VGND.t1805 119.309
R3038 VGND.n1259 VGND.t1853 119.309
R3039 VGND.n1262 VGND.t1892 119.309
R3040 VGND.n998 VGND.t1901 119.309
R3041 VGND.n1265 VGND.t1817 119.309
R3042 VGND.n5 VGND.n3 117.001
R3043 VGND.t1456 VGND.n5 117.001
R3044 VGND.n6 VGND.n4 117.001
R3045 VGND.n328 VGND.n6 117.001
R3046 VGND.t2293 VGND.t1824 110.535
R3047 VGND.t497 VGND.t2645 110.535
R3048 VGND.t1773 VGND.t2639 110.535
R3049 VGND.t2565 VGND.t38 110.535
R3050 VGND.t2368 VGND.t1779 110.535
R3051 VGND.t1712 VGND.t2361 110.535
R3052 VGND.t1797 VGND.t2346 110.535
R3053 VGND.t1702 VGND.t764 110.535
R3054 VGND.t2281 VGND.t1872 110.535
R3055 VGND.t39 VGND.t2633 110.535
R3056 VGND.t1878 VGND.t2617 110.535
R3057 VGND.t2349 VGND.t767 110.535
R3058 VGND.t2604 VGND.t1800 110.535
R3059 VGND.t1292 VGND.t2284 110.535
R3060 VGND.t1842 VGND.t2275 110.535
R3061 VGND.t1692 VGND.t1171 110.535
R3062 VGND.t1686 VGND.t1851 110.535
R3063 VGND.t1295 VGND.t2606 110.535
R3064 VGND.t1890 VGND.t2619 110.535
R3065 VGND.t2350 VGND.t1445 110.535
R3066 VGND.t2334 VGND.t1806 110.535
R3067 VGND.t2371 VGND.t1689 110.535
R3068 VGND.t1854 VGND.t2325 110.535
R3069 VGND.t1677 VGND.t800 110.535
R3070 VGND.t2600 VGND.t1893 110.535
R3071 VGND.t72 VGND.t2593 110.535
R3072 VGND.t1902 VGND.t2588 110.535
R3073 VGND.t2327 VGND.t51 110.535
R3074 VGND.t2566 VGND.t1818 110.535
R3075 VGND.t884 VGND.t2306 110.535
R3076 VGND.t1860 VGND.t1673 110.535
R3077 VGND.t2590 VGND.t1217 110.535
R3078 VGND.t1297 VGND.t1307 92.4699
R3079 VGND.t1307 VGND.t1304 92.4699
R3080 VGND.t1304 VGND.t1308 92.4699
R3081 VGND.t1308 VGND.t1454 92.4699
R3082 VGND.t1454 VGND.t2261 92.4699
R3083 VGND.t2261 VGND.t1439 92.4699
R3084 VGND.t1439 VGND.t2218 92.4699
R3085 VGND VGND.n806 80.9529
R3086 VGND VGND.n806 75.1009
R3087 VGND.n1337 VGND 74.8566
R3088 VGND.t2218 VGND 70.4533
R3089 VGND.n2285 VGND 58.8055
R3090 VGND.n2284 VGND 58.8055
R3091 VGND.n2250 VGND 58.8055
R3092 VGND.n2248 VGND 58.8055
R3093 VGND.n1386 VGND 58.8055
R3094 VGND.n2348 VGND.n2347 53.1823
R3095 VGND.n2349 VGND.n2348 53.1823
R3096 VGND.n3021 VGND.n3020 53.1823
R3097 VGND.n3020 VGND.n3019 53.1823
R3098 VGND.t1557 VGND.t2454 50.5752
R3099 VGND.t1553 VGND.t389 50.5752
R3100 VGND.t1547 VGND.t453 50.5752
R3101 VGND.t1549 VGND.t475 50.5752
R3102 VGND.t1305 VGND.t1452 50.5752
R3103 VGND.t1302 VGND.t2259 50.5752
R3104 VGND.t1300 VGND.t596 50.5752
R3105 VGND.t1298 VGND.t491 50.5752
R3106 VGND VGND.n2981 43.2063
R3107 VGND VGND.n18 43.2063
R3108 VGND VGND.n2951 43.2063
R3109 VGND VGND.n44 43.2063
R3110 VGND.n2347 VGND.n2346 40.6593
R3111 VGND.n886 VGND.t1691 34.8005
R3112 VGND.n886 VGND.t2610 34.8005
R3113 VGND.n889 VGND.t2608 34.8005
R3114 VGND.n889 VGND.t2340 34.8005
R3115 VGND.n893 VGND.t2337 34.8005
R3116 VGND.n893 VGND.t1694 34.8005
R3117 VGND.n930 VGND.t2315 34.8005
R3118 VGND.n930 VGND.t1672 34.8005
R3119 VGND.n935 VGND.t2603 34.8005
R3120 VGND.n935 VGND.t2599 34.8005
R3121 VGND.n940 VGND.t2592 34.8005
R3122 VGND.n940 VGND.t2321 34.8005
R3123 VGND.n945 VGND.t2573 34.8005
R3124 VGND.n945 VGND.t2310 34.8005
R3125 VGND.n950 VGND.t1676 34.8005
R3126 VGND.n950 VGND.t2595 34.8005
R3127 VGND.n955 VGND.t1655 34.8005
R3128 VGND.n955 VGND.t2577 34.8005
R3129 VGND.n960 VGND.t2569 34.8005
R3130 VGND.n960 VGND.t2323 34.8005
R3131 VGND.n965 VGND.t2303 34.8005
R3132 VGND.n965 VGND.t1659 34.8005
R3133 VGND.n970 VGND.t2290 34.8005
R3134 VGND.n970 VGND.t2643 34.8005
R3135 VGND.n975 VGND.t2627 34.8005
R3136 VGND.n975 VGND.t2305 34.8005
R3137 VGND.n980 VGND.t2363 34.8005
R3138 VGND.n980 VGND.t2292 34.8005
R3139 VGND.n985 VGND.t1705 34.8005
R3140 VGND.n985 VGND.t1700 34.8005
R3141 VGND.n996 VGND.t2319 34.8005
R3142 VGND.n996 VGND.t1674 34.8005
R3143 VGND.n1273 VGND.t2575 34.8005
R3144 VGND.n1273 VGND.t2567 34.8005
R3145 VGND.n1230 VGND.t1670 34.8005
R3146 VGND.n1230 VGND.t2589 34.8005
R3147 VGND.n1229 VGND.t2308 34.8005
R3148 VGND.n1229 VGND.t2601 34.8005
R3149 VGND.n1226 VGND.t2586 34.8005
R3150 VGND.n1226 VGND.t2326 34.8005
R3151 VGND.n1224 VGND.t2597 34.8005
R3152 VGND.n1224 VGND.t2335 34.8005
R3153 VGND.n1221 VGND.t1680 34.8005
R3154 VGND.n1221 VGND.t2620 34.8005
R3155 VGND.n1216 VGND.t2333 34.8005
R3156 VGND.n1216 VGND.t1687 34.8005
R3157 VGND.n1002 VGND.t2353 34.8005
R3158 VGND.n1002 VGND.t2276 34.8005
R3159 VGND.n1203 VGND.t1685 34.8005
R3160 VGND.n1203 VGND.t2605 34.8005
R3161 VGND.n1007 VGND.t1707 34.8005
R3162 VGND.n1007 VGND.t2618 34.8005
R3163 VGND.n1184 VGND.t2286 34.8005
R3164 VGND.n1184 VGND.t2282 34.8005
R3165 VGND.n1010 VGND.t2614 34.8005
R3166 VGND.n1010 VGND.t2347 34.8005
R3167 VGND.n1171 VGND.t2638 34.8005
R3168 VGND.n1171 VGND.t2369 34.8005
R3169 VGND.n1012 VGND.t2288 34.8005
R3170 VGND.n1012 VGND.t2640 34.8005
R3171 VGND.n329 VGND.t2313 34.8005
R3172 VGND.n329 VGND.t1668 34.8005
R3173 VGND.n332 VGND.t1666 34.8005
R3174 VGND.n332 VGND.t2584 34.8005
R3175 VGND.n356 VGND.t2582 34.8005
R3176 VGND.n356 VGND.t2317 34.8005
R3177 VGND.n363 VGND.t2560 34.8005
R3178 VGND.n363 VGND.t2297 34.8005
R3179 VGND.n366 VGND.t1664 34.8005
R3180 VGND.n366 VGND.t1661 34.8005
R3181 VGND.n374 VGND.t1653 34.8005
R3182 VGND.n374 VGND.t2562 34.8005
R3183 VGND.n377 VGND.t2629 34.8005
R3184 VGND.n377 VGND.t2359 34.8005
R3185 VGND.n385 VGND.t2301 34.8005
R3186 VGND.n385 VGND.t1657 34.8005
R3187 VGND.n324 VGND.t2278 34.8005
R3188 VGND.n324 VGND.t2631 34.8005
R3189 VGND.n313 VGND.t2625 34.8005
R3190 VGND.n313 VGND.t2564 34.8005
R3191 VGND.n308 VGND.t2355 34.8005
R3192 VGND.n308 VGND.t2280 34.8005
R3193 VGND.n310 VGND.t2343 34.8005
R3194 VGND.n310 VGND.t1698 34.8005
R3195 VGND.n2729 VGND.t1682 34.8005
R3196 VGND.n2729 VGND.t2357 34.8005
R3197 VGND.n292 VGND.t2612 34.8005
R3198 VGND.n292 VGND.t2345 34.8005
R3199 VGND.n295 VGND.t2331 34.8005
R3200 VGND.n295 VGND.t2329 34.8005
R3201 VGND.n202 VGND.t1696 34.8005
R3202 VGND.n202 VGND.t2616 34.8005
R3203 VGND.n395 VGND.t1810 34.8005
R3204 VGND.n395 VGND.t945 34.8005
R3205 VGND.n2637 VGND.t1271 34.8005
R3206 VGND.n2637 VGND.t2519 34.8005
R3207 VGND.n2642 VGND.t1967 34.8005
R3208 VGND.n2642 VGND.t953 34.8005
R3209 VGND.n2647 VGND.t681 34.8005
R3210 VGND.n2647 VGND.t951 34.8005
R3211 VGND.n2652 VGND.t859 34.8005
R3212 VGND.n2652 VGND.t2527 34.8005
R3213 VGND.n2657 VGND.t695 34.8005
R3214 VGND.n2657 VGND.t2535 34.8005
R3215 VGND.n2662 VGND.t2049 34.8005
R3216 VGND.n2662 VGND.t2533 34.8005
R3217 VGND.n2667 VGND.t669 34.8005
R3218 VGND.n2667 VGND.t2525 34.8005
R3219 VGND.n392 VGND.t422 34.8005
R3220 VGND.n392 VGND.t2523 34.8005
R3221 VGND.n2713 VGND.t1934 34.8005
R3222 VGND.n2713 VGND.t2537 34.8005
R3223 VGND.n318 VGND.t542 34.8005
R3224 VGND.n318 VGND.t949 34.8005
R3225 VGND.n2746 VGND.t1101 34.8005
R3226 VGND.n2746 VGND.t947 34.8005
R3227 VGND.n302 VGND.t1982 34.8005
R3228 VGND.n302 VGND.t2531 34.8005
R3229 VGND.n2751 VGND.t729 34.8005
R3230 VGND.n2751 VGND.t2529 34.8005
R3231 VGND.n2786 VGND.t1599 34.8005
R3232 VGND.n2786 VGND.t955 34.8005
R3233 VGND.n285 VGND.t1585 34.8005
R3234 VGND.n285 VGND.t2521 34.8005
R3235 VGND.n399 VGND.t1885 34.8005
R3236 VGND.n399 VGND.t2683 34.8005
R3237 VGND.n2341 VGND.t1499 34.8005
R3238 VGND.n2341 VGND.t2064 34.8005
R3239 VGND.n2336 VGND.t1959 34.8005
R3240 VGND.n2336 VGND.t611 34.8005
R3241 VGND.n2331 VGND.t2496 34.8005
R3242 VGND.n2331 VGND.t1409 34.8005
R3243 VGND.n2326 VGND.t535 34.8005
R3244 VGND.n2326 VGND.t2681 34.8005
R3245 VGND.n2321 VGND.t1957 34.8005
R3246 VGND.n2321 VGND.t2060 34.8005
R3247 VGND.n2316 VGND.t81 34.8005
R3248 VGND.n2316 VGND.t2058 34.8005
R3249 VGND.n2311 VGND.t2124 34.8005
R3250 VGND.n2311 VGND.t2679 34.8005
R3251 VGND.n2306 VGND.t799 34.8005
R3252 VGND.n2306 VGND.t2677 34.8005
R3253 VGND.n2301 VGND.t781 34.8005
R3254 VGND.n2301 VGND.t2062 34.8005
R3255 VGND.n2296 VGND.t586 34.8005
R3256 VGND.n2296 VGND.t1421 34.8005
R3257 VGND.n2291 VGND.t2470 34.8005
R3258 VGND.n2291 VGND.t1419 34.8005
R3259 VGND.n2286 VGND.t2415 34.8005
R3260 VGND.n2286 VGND.t617 34.8005
R3261 VGND.n413 VGND.t2163 34.8005
R3262 VGND.n413 VGND.t615 34.8005
R3263 VGND.n2539 VGND.t1261 34.8005
R3264 VGND.n2539 VGND.t613 34.8005
R3265 VGND.n416 VGND.t325 34.8005
R3266 VGND.n416 VGND.t2066 34.8005
R3267 VGND.n468 VGND.t1792 34.8005
R3268 VGND.n468 VGND.t2142 34.8005
R3269 VGND.n470 VGND.t2665 34.8005
R3270 VGND.n470 VGND.t1427 34.8005
R3271 VGND.n2375 VGND.t2655 34.8005
R3272 VGND.n2375 VGND.t2150 34.8005
R3273 VGND.n458 VGND.t1157 34.8005
R3274 VGND.n458 VGND.t2148 34.8005
R3275 VGND.n2401 VGND.t1738 34.8005
R3276 VGND.n2401 VGND.t2140 34.8005
R3277 VGND.n450 VGND.t701 34.8005
R3278 VGND.n450 VGND.t1423 34.8005
R3279 VGND.n2427 VGND.t1988 34.8005
R3280 VGND.n2427 VGND.t2687 34.8005
R3281 VGND.n442 VGND.t675 34.8005
R3282 VGND.n442 VGND.t2138 34.8005
R3283 VGND.n2453 VGND.t1122 34.8005
R3284 VGND.n2453 VGND.t1431 34.8005
R3285 VGND.n434 VGND.t709 34.8005
R3286 VGND.n434 VGND.t1425 34.8005
R3287 VGND.n2479 VGND.t785 34.8005
R3288 VGND.n2479 VGND.t2146 34.8005
R3289 VGND.n426 VGND.t2673 34.8005
R3290 VGND.n426 VGND.t2144 34.8005
R3291 VGND.n2510 VGND.t1975 34.8005
R3292 VGND.n2510 VGND.t2685 34.8005
R3293 VGND.n2515 VGND.t735 34.8005
R3294 VGND.n2515 VGND.t1444 34.8005
R3295 VGND.n2520 VGND.t2555 34.8005
R3296 VGND.n2520 VGND.t2152 34.8005
R3297 VGND.n418 VGND.t1592 34.8005
R3298 VGND.n418 VGND.t1429 34.8005
R3299 VGND.n465 VGND.t1834 34.8005
R3300 VGND.n465 VGND.t2444 34.8005
R3301 VGND.n2362 VGND.t1285 34.8005
R3302 VGND.n2362 VGND.t234 34.8005
R3303 VGND.n462 VGND.t2110 34.8005
R3304 VGND.n462 VGND.t607 34.8005
R3305 VGND.n2388 VGND.t1068 34.8005
R3306 VGND.n2388 VGND.t605 34.8005
R3307 VGND.n454 VGND.t987 34.8005
R3308 VGND.n454 VGND.t2442 34.8005
R3309 VGND.n2414 VGND.t873 34.8005
R3310 VGND.n2414 VGND.t230 34.8005
R3311 VGND.n446 VGND.t751 34.8005
R3312 VGND.n446 VGND.t228 34.8005
R3313 VGND.n2440 VGND.t2244 34.8005
R3314 VGND.n2440 VGND.t2440 34.8005
R3315 VGND.n438 VGND.t1151 34.8005
R3316 VGND.n438 VGND.t2136 34.8005
R3317 VGND.n2466 VGND.t1113 34.8005
R3318 VGND.n2466 VGND.t232 34.8005
R3319 VGND.n430 VGND.t528 34.8005
R3320 VGND.n430 VGND.t2448 34.8005
R3321 VGND.n2492 VGND.t1093 34.8005
R3322 VGND.n2492 VGND.t2446 34.8005
R3323 VGND.n422 VGND.t139 34.8005
R3324 VGND.n422 VGND.t226 34.8005
R3325 VGND.n2497 VGND.t1503 34.8005
R3326 VGND.n2497 VGND.t224 34.8005
R3327 VGND.n2808 VGND.t14 34.8005
R3328 VGND.n2808 VGND.t609 34.8005
R3329 VGND.n276 VGND.t1254 34.8005
R3330 VGND.n276 VGND.t2134 34.8005
R3331 VGND.n624 VGND.t1906 34.8005
R3332 VGND.n624 VGND.t125 34.8005
R3333 VGND.n1909 VGND.t814 34.8005
R3334 VGND.n1909 VGND.t937 34.8005
R3335 VGND.n621 VGND.t1186 34.8005
R3336 VGND.n621 VGND.t2475 34.8005
R3337 VGND.n1920 VGND.t2490 34.8005
R3338 VGND.n1920 VGND.t89 34.8005
R3339 VGND.n618 VGND.t260 34.8005
R3340 VGND.n618 VGND.t123 34.8005
R3341 VGND.n1931 VGND.t2070 34.8005
R3342 VGND.n1931 VGND.t933 34.8005
R3343 VGND.n615 VGND.t77 34.8005
R3344 VGND.n615 VGND.t931 34.8005
R3345 VGND.n1942 VGND.t593 34.8005
R3346 VGND.n1942 VGND.t121 34.8005
R3347 VGND.n612 VGND.t793 34.8005
R3348 VGND.n612 VGND.t119 34.8005
R3349 VGND.n1953 VGND.t158 34.8005
R3350 VGND.n1953 VGND.t935 34.8005
R3351 VGND.n609 VGND.t581 34.8005
R3352 VGND.n609 VGND.t87 34.8005
R3353 VGND.n1964 VGND.t2466 34.8005
R3354 VGND.n1964 VGND.t85 34.8005
R3355 VGND.n606 VGND.t1971 34.8005
R3356 VGND.n606 VGND.t929 34.8005
R3357 VGND.n1975 VGND.t2157 34.8005
R3358 VGND.n1975 VGND.t927 34.8005
R3359 VGND.n1980 VGND.t43 34.8005
R3360 VGND.n1980 VGND.t2477 34.8005
R3361 VGND.n605 VGND.t339 34.8005
R3362 VGND.n605 VGND.t117 34.8005
R3363 VGND.n589 VGND.t1813 34.8005
R3364 VGND.n589 VGND.t2384 34.8005
R3365 VGND.n595 VGND.t1269 34.8005
R3366 VGND.n595 VGND.t2374 34.8005
R3367 VGND.n592 VGND.t1965 34.8005
R3368 VGND.n592 VGND.t1236 34.8005
R3369 VGND.n2054 VGND.t62 34.8005
R3370 VGND.n2054 VGND.t1234 34.8005
R3371 VGND.n2049 VGND.t857 34.8005
R3372 VGND.n2049 VGND.t2382 34.8005
R3373 VGND.n2044 VGND.t693 34.8005
R3374 VGND.n2044 VGND.t1574 34.8005
R3375 VGND.n2039 VGND.t2047 34.8005
R3376 VGND.n2039 VGND.t1572 34.8005
R3377 VGND.n2034 VGND.t667 34.8005
R3378 VGND.n2034 VGND.t2380 34.8005
R3379 VGND.n2029 VGND.t420 34.8005
R3380 VGND.n2029 VGND.t2378 34.8005
R3381 VGND.n2024 VGND.t1932 34.8005
R3382 VGND.n2024 VGND.t1576 34.8005
R3383 VGND.n2019 VGND.t539 34.8005
R3384 VGND.n2019 VGND.t1232 34.8005
R3385 VGND.n2014 VGND.t1099 34.8005
R3386 VGND.n2014 VGND.t1230 34.8005
R3387 VGND.n2009 VGND.t2420 34.8005
R3388 VGND.n2009 VGND.t1570 34.8005
R3389 VGND.n2004 VGND.t727 34.8005
R3390 VGND.n2004 VGND.t1240 34.8005
R3391 VGND.n600 VGND.t2418 34.8005
R3392 VGND.n600 VGND.t1238 34.8005
R3393 VGND.n1993 VGND.t1583 34.8005
R3394 VGND.n1993 VGND.t2376 34.8005
R3395 VGND.n586 VGND.t1786 34.8005
R3396 VGND.n586 VGND.t516 34.8005
R3397 VGND.n2068 VGND.t2667 34.8005
R3398 VGND.n2068 VGND.t577 34.8005
R3399 VGND.n2073 VGND.t2657 34.8005
R3400 VGND.n2073 VGND.t479 34.8005
R3401 VGND.n2078 VGND.t1155 34.8005
R3402 VGND.n2078 VGND.t522 34.8005
R3403 VGND.n2083 VGND.t1740 34.8005
R3404 VGND.n2083 VGND.t514 34.8005
R3405 VGND.n2088 VGND.t2211 34.8005
R3406 VGND.n2088 VGND.t573 34.8005
R3407 VGND.n2093 VGND.t1990 34.8005
R3408 VGND.n2093 VGND.t571 34.8005
R3409 VGND.n2098 VGND.t677 34.8005
R3410 VGND.n2098 VGND.t512 34.8005
R3411 VGND.n2103 VGND.t1 34.8005
R3412 VGND.n2103 VGND.t510 34.8005
R3413 VGND.n2108 VGND.t711 34.8005
R3414 VGND.n2108 VGND.t575 34.8005
R3415 VGND.n2113 VGND.t787 34.8005
R3416 VGND.n2113 VGND.t520 34.8005
R3417 VGND.n2118 VGND.t2675 34.8005
R3418 VGND.n2118 VGND.t518 34.8005
R3419 VGND.n583 VGND.t1977 34.8005
R3420 VGND.n583 VGND.t569 34.8005
R3421 VGND.n2123 VGND.t737 34.8005
R3422 VGND.n2123 VGND.t483 34.8005
R3423 VGND.n2833 VGND.t2557 34.8005
R3424 VGND.n2833 VGND.t481 34.8005
R3425 VGND.n264 VGND.t333 34.8005
R3426 VGND.n264 VGND.t579 34.8005
R3427 VGND.n546 VGND.t1828 34.8005
R3428 VGND.n546 VGND.t756 34.8005
R3429 VGND.n549 VGND.t1287 34.8005
R3430 VGND.n549 VGND.t469 34.8005
R3431 VGND.n1755 VGND.t2092 34.8005
R3432 VGND.n1755 VGND.t1203 34.8005
R3433 VGND.n1760 VGND.t1066 34.8005
R3434 VGND.n1760 VGND.t1201 34.8005
R3435 VGND.n1751 VGND.t989 34.8005
R3436 VGND.n1751 VGND.t153 34.8005
R3437 VGND.n1771 VGND.t875 34.8005
R3438 VGND.n1771 VGND.t688 34.8005
R3439 VGND.n1748 VGND.t753 34.8005
R3440 VGND.n1748 VGND.t686 34.8005
R3441 VGND.n1782 VGND.t2246 34.8005
R3442 VGND.n1782 VGND.t151 34.8005
R3443 VGND.n1745 VGND.t1215 34.8005
R3444 VGND.n1745 VGND.t149 34.8005
R3445 VGND.n1793 VGND.t1115 34.8005
R3446 VGND.n1793 VGND.t690 34.8005
R3447 VGND.n1742 VGND.t530 34.8005
R3448 VGND.n1742 VGND.t760 34.8005
R3449 VGND.n1804 VGND.t1095 34.8005
R3450 VGND.n1804 VGND.t758 34.8005
R3451 VGND.n1739 VGND.t141 34.8005
R3452 VGND.n1739 VGND.t684 34.8005
R3453 VGND.n1815 VGND.t1505 34.8005
R3454 VGND.n1815 VGND.t1207 34.8005
R3455 VGND.n1820 VGND.t34 34.8005
R3456 VGND.n1820 VGND.t1205 34.8005
R3457 VGND.n1738 VGND.t1256 34.8005
R3458 VGND.n1738 VGND.t147 34.8005
R3459 VGND.n627 VGND.t1840 34.8005
R3460 VGND.n627 VGND.t743 34.8005
R3461 VGND.n1677 VGND.t1280 34.8005
R3462 VGND.n1677 VGND.t316 34.8005
R3463 VGND.n1674 VGND.t2104 34.8005
R3464 VGND.n1674 VGND.t2207 34.8005
R3465 VGND.n1688 VGND.t1072 34.8005
R3466 VGND.n1688 VGND.t2205 34.8005
R3467 VGND.n1693 VGND.t983 34.8005
R3468 VGND.n1693 VGND.t741 34.8005
R3469 VGND.n1698 VGND.t170 34.8005
R3470 VGND.n1698 VGND.t312 34.8005
R3471 VGND.n1703 VGND.t2056 34.8005
R3472 VGND.n1703 VGND.t1054 34.8005
R3473 VGND.n1708 VGND.t2240 34.8005
R3474 VGND.n1708 VGND.t739 34.8005
R3475 VGND.n1713 VGND.t1147 34.8005
R3476 VGND.n1713 VGND.t2045 34.8005
R3477 VGND.n1718 VGND.t1228 34.8005
R3478 VGND.n1718 VGND.t314 34.8005
R3479 VGND.n1723 VGND.t526 34.8005
R3480 VGND.n1723 VGND.t2203 34.8005
R3481 VGND.n1728 VGND.t1091 34.8005
R3482 VGND.n1728 VGND.t745 34.8005
R3483 VGND.n1671 VGND.t2426 34.8005
R3484 VGND.n1671 VGND.t1052 34.8005
R3485 VGND.n1844 VGND.t1416 34.8005
R3486 VGND.n1844 VGND.t1050 34.8005
R3487 VGND.n1733 VGND.t10 34.8005
R3488 VGND.n1733 VGND.t2209 34.8005
R3489 VGND.n1833 VGND.t1252 34.8005
R3490 VGND.n1833 VGND.t318 34.8005
R3491 VGND.n631 VGND.t1768 34.8005
R3492 VGND.n631 VGND.t2182 34.8005
R3493 VGND.n668 VGND.t812 34.8005
R3494 VGND.n668 VGND.t2172 34.8005
R3495 VGND.n673 VGND.t1184 34.8005
R3496 VGND.n673 VGND.t2132 34.8005
R3497 VGND.n678 VGND.t2492 34.8005
R3498 VGND.n678 VGND.t2130 34.8005
R3499 VGND.n683 VGND.t258 34.8005
R3500 VGND.n683 VGND.t2180 34.8005
R3501 VGND.n688 VGND.t2068 34.8005
R3502 VGND.n688 VGND.t31 34.8005
R3503 VGND.n693 VGND.t75 34.8005
R3504 VGND.n693 VGND.t29 34.8005
R3505 VGND.n698 VGND.t591 34.8005
R3506 VGND.n698 VGND.t2178 34.8005
R3507 VGND.n703 VGND.t4 34.8005
R3508 VGND.n703 VGND.t2176 34.8005
R3509 VGND.n708 VGND.t156 34.8005
R3510 VGND.n708 VGND.t2170 34.8005
R3511 VGND.n713 VGND.t791 34.8005
R3512 VGND.n713 VGND.t2128 34.8005
R3513 VGND.n718 VGND.t2464 34.8005
R3514 VGND.n718 VGND.t2126 34.8005
R3515 VGND.n665 VGND.t1969 34.8005
R3516 VGND.n665 VGND.t27 34.8005
R3517 VGND.n723 VGND.t2155 34.8005
R3518 VGND.n723 VGND.t25 34.8005
R3519 VGND.n2858 VGND.t41 34.8005
R3520 VGND.n2858 VGND.t23 34.8005
R3521 VGND.n252 VGND.t337 34.8005
R3522 VGND.n252 VGND.t2174 34.8005
R3523 VGND.n878 VGND.t1864 34.8005
R3524 VGND.n878 VGND.t300 34.8005
R3525 VGND.n1351 VGND.t2167 34.8005
R3526 VGND.n1351 VGND.t2194 34.8005
R3527 VGND.n873 VGND.t251 34.8005
R3528 VGND.n873 VGND.t308 34.8005
R3529 VGND.n807 VGND.t1059 34.8005
R3530 VGND.n807 VGND.t306 34.8005
R3531 VGND.n809 VGND.t2229 34.8005
R3532 VGND.n809 VGND.t298 34.8005
R3533 VGND.n822 VGND.t2087 34.8005
R3534 VGND.n822 VGND.t2190 34.8005
R3535 VGND.n827 VGND.t2253 34.8005
R3536 VGND.n827 VGND.t2188 34.8005
R3537 VGND.n832 VGND.t2514 34.8005
R3538 VGND.n832 VGND.t2200 34.8005
R3539 VGND.n837 VGND.t774 34.8005
R3540 VGND.n837 VGND.t2198 34.8005
R3541 VGND.n842 VGND.t2097 34.8005
R3542 VGND.n842 VGND.t2192 34.8005
R3543 VGND.n847 VGND.t506 34.8005
R3544 VGND.n847 VGND.t304 34.8005
R3545 VGND.n818 VGND.t345 34.8005
R3546 VGND.n818 VGND.t302 34.8005
R3547 VGND.n852 VGND.t1338 34.8005
R3548 VGND.n852 VGND.t2186 34.8005
R3549 VGND.n733 VGND.t2119 34.8005
R3550 VGND.n733 VGND.t2184 34.8005
R3551 VGND.n1660 VGND.t6 34.8005
R3552 VGND.n1660 VGND.t310 34.8005
R3553 VGND.n736 VGND.t1244 34.8005
R3554 VGND.n736 VGND.t2196 34.8005
R3555 VGND.n799 VGND.t1795 34.8005
R3556 VGND.n799 VGND.t424 34.8005
R3557 VGND.n1389 VGND.t2663 34.8005
R3558 VGND.n1389 VGND.t914 34.8005
R3559 VGND.n1394 VGND.t2653 34.8005
R3560 VGND.n1394 VGND.t432 34.8005
R3561 VGND.n803 VGND.t1159 34.8005
R3562 VGND.n803 VGND.t430 34.8005
R3563 VGND.n1489 VGND.t864 34.8005
R3564 VGND.n1489 VGND.t922 34.8005
R3565 VGND.n775 VGND.t699 34.8005
R3566 VGND.n775 VGND.t910 34.8005
R3567 VGND.n1515 VGND.t1986 34.8005
R3568 VGND.n1515 VGND.t2435 34.8005
R3569 VGND.n767 VGND.t673 34.8005
R3570 VGND.n767 VGND.t920 34.8005
R3571 VGND.n1541 VGND.t1120 34.8005
R3572 VGND.n1541 VGND.t918 34.8005
R3573 VGND.n1546 VGND.t707 34.8005
R3574 VGND.n1546 VGND.t912 34.8005
R3575 VGND.n759 VGND.t546 34.8005
R3576 VGND.n759 VGND.t428 34.8005
R3577 VGND.n1551 VGND.t2671 34.8005
R3578 VGND.n1551 VGND.t426 34.8005
R3579 VGND.n1631 VGND.t1973 34.8005
R3580 VGND.n1631 VGND.t2433 34.8005
R3581 VGND.n1636 VGND.t733 34.8005
R3582 VGND.n1636 VGND.t416 34.8005
R3583 VGND.n1641 VGND.t2553 34.8005
R3584 VGND.n1641 VGND.t434 34.8005
R3585 VGND.n739 VGND.t1590 34.8005
R3586 VGND.n739 VGND.t916 34.8005
R3587 VGND.n796 VGND.t1867 34.8005
R3588 VGND.n796 VGND.t2501 34.8005
R3589 VGND.n1409 VGND.t2165 34.8005
R3590 VGND.n1409 VGND.t2549 34.8005
R3591 VGND.n793 VGND.t705 34.8005
R3592 VGND.n793 VGND.t808 34.8005
R3593 VGND.n1476 VGND.t1061 34.8005
R3594 VGND.n1476 VGND.t806 34.8005
R3595 VGND.n779 VGND.t2227 34.8005
R3596 VGND.n779 VGND.t1564 34.8005
R3597 VGND.n1502 VGND.t246 34.8005
R3598 VGND.n1502 VGND.t2545 34.8005
R3599 VGND.n771 VGND.t2251 34.8005
R3600 VGND.n771 VGND.t2543 34.8005
R3601 VGND.n1528 VGND.t2512 34.8005
R3602 VGND.n1528 VGND.t1562 34.8005
R3603 VGND.n763 VGND.t772 34.8005
R3604 VGND.n763 VGND.t1560 34.8005
R3605 VGND.n1565 VGND.t2095 34.8005
R3606 VGND.n1565 VGND.t2547 34.8005
R3607 VGND.n754 VGND.t504 34.8005
R3608 VGND.n754 VGND.t804 34.8005
R3609 VGND.n1580 VGND.t722 34.8005
R3610 VGND.n1580 VGND.t802 34.8005
R3611 VGND.n1575 VGND.t1336 34.8005
R3612 VGND.n1575 VGND.t2541 34.8005
R3613 VGND.n1570 VGND.t2117 34.8005
R3614 VGND.n1570 VGND.t2539 34.8005
R3615 VGND.n2883 VGND.t18 34.8005
R3616 VGND.n2883 VGND.t810 34.8005
R3617 VGND.n239 VGND.t296 34.8005
R3618 VGND.n239 VGND.t2551 34.8005
R3619 VGND.n881 VGND.t1897 34.8005
R3620 VGND.n881 VGND.t850 34.8005
R3621 VGND.n883 VGND.t1497 34.8005
R3622 VGND.n883 VGND.t840 34.8005
R3623 VGND.n1422 VGND.t1190 34.8005
R3624 VGND.n1422 VGND.t1567 34.8005
R3625 VGND.n1427 VGND.t714 34.8005
R3626 VGND.n1427 VGND.t2274 34.8005
R3627 VGND.n1432 VGND.t264 34.8005
R3628 VGND.n1432 VGND.t848 34.8005
R3629 VGND.n1437 VGND.t1955 34.8005
R3630 VGND.n1437 VGND.t1515 34.8005
R3631 VGND.n1442 VGND.t79 34.8005
R3632 VGND.n1442 VGND.t1513 34.8005
R3633 VGND.n1447 VGND.t2122 34.8005
R3634 VGND.n1447 VGND.t846 34.8005
R3635 VGND.n1452 VGND.t797 34.8005
R3636 VGND.n1452 VGND.t844 34.8005
R3637 VGND.n789 VGND.t779 34.8005
R3638 VGND.n789 VGND.t1517 34.8005
R3639 VGND.n1457 VGND.t583 34.8005
R3640 VGND.n1457 VGND.t2272 34.8005
R3641 VGND.n1594 VGND.t2468 34.8005
R3642 VGND.n1594 VGND.t2270 34.8005
R3643 VGND.n1599 VGND.t2412 34.8005
R3644 VGND.n1599 VGND.t1511 34.8005
R3645 VGND.n748 VGND.t2161 34.8005
R3646 VGND.n748 VGND.t1509 34.8005
R3647 VGND.n1612 VGND.t1258 34.8005
R3648 VGND.n1612 VGND.t1507 34.8005
R3649 VGND.n1604 VGND.t322 34.8005
R3650 VGND.n1604 VGND.t842 34.8005
R3651 VGND.n1023 VGND.t1837 34.8005
R3652 VGND.n1023 VGND.t135 34.8005
R3653 VGND.n1030 VGND.t1282 34.8005
R3654 VGND.n1030 VGND.t1946 34.8005
R3655 VGND.n1035 VGND.t2106 34.8005
R3656 VGND.n1035 VGND.t449 34.8005
R3657 VGND.n1027 VGND.t1070 34.8005
R3658 VGND.n1027 VGND.t447 34.8005
R3659 VGND.n1093 VGND.t985 34.8005
R3660 VGND.n1093 VGND.t133 34.8005
R3661 VGND.n1088 VGND.t172 34.8005
R3662 VGND.n1088 VGND.t1087 34.8005
R3663 VGND.n1083 VGND.t2054 34.8005
R3664 VGND.n1083 VGND.t1085 34.8005
R3665 VGND.n1078 VGND.t2238 34.8005
R3666 VGND.n1078 VGND.t131 34.8005
R3667 VGND.n1073 VGND.t1145 34.8005
R3668 VGND.n1073 VGND.t129 34.8005
R3669 VGND.n1040 VGND.t1226 34.8005
R3670 VGND.n1040 VGND.t1944 34.8005
R3671 VGND.n1042 VGND.t524 34.8005
R3672 VGND.n1042 VGND.t445 34.8005
R3673 VGND.n1051 VGND.t1089 34.8005
R3674 VGND.n1051 VGND.t137 34.8005
R3675 VGND.n1056 VGND.t2424 34.8005
R3676 VGND.n1056 VGND.t1083 34.8005
R3677 VGND.n1047 VGND.t1414 34.8005
R3678 VGND.n1047 VGND.t1081 34.8005
R3679 VGND.n2903 VGND.t12 34.8005
R3680 VGND.n2903 VGND.t1079 34.8005
R3681 VGND.n227 VGND.t1250 34.8005
R3682 VGND.n227 VGND.t1948 34.8005
R3683 VGND.n1013 VGND.t2365 34.8005
R3684 VGND.n1013 VGND.t2294 34.8005
R3685 VGND.n926 VGND.t2636 34.8005
R3686 VGND.n926 VGND.t2367 34.8005
R3687 VGND.n105 VGND.n103 34.6358
R3688 VGND.n2984 VGND.n2978 34.6358
R3689 VGND.n2987 VGND.n2986 34.6358
R3690 VGND.n2987 VGND.n2974 34.6358
R3691 VGND.n2991 VGND.n2974 34.6358
R3692 VGND.n2992 VGND.n2991 34.6358
R3693 VGND.n2993 VGND.n2992 34.6358
R3694 VGND.n21 VGND.n20 34.6358
R3695 VGND.n23 VGND.n12 34.6358
R3696 VGND.n27 VGND.n12 34.6358
R3697 VGND.n28 VGND.n27 34.6358
R3698 VGND.n29 VGND.n28 34.6358
R3699 VGND.n29 VGND.n9 34.6358
R3700 VGND.n3006 VGND.n10 34.6358
R3701 VGND.n181 VGND.n180 34.6358
R3702 VGND.n185 VGND.n184 34.6358
R3703 VGND.n2954 VGND.n2953 34.6358
R3704 VGND.n2956 VGND.n2947 34.6358
R3705 VGND.n2960 VGND.n2947 34.6358
R3706 VGND.n2961 VGND.n2960 34.6358
R3707 VGND.n2962 VGND.n2961 34.6358
R3708 VGND.n2962 VGND.n2945 34.6358
R3709 VGND.n47 VGND.n46 34.6358
R3710 VGND.n49 VGND.n38 34.6358
R3711 VGND.n53 VGND.n38 34.6358
R3712 VGND.n54 VGND.n53 34.6358
R3713 VGND.n55 VGND.n54 34.6358
R3714 VGND.n55 VGND.n35 34.6358
R3715 VGND.n109 VGND.n108 34.6358
R3716 VGND.n82 VGND.n81 34.6358
R3717 VGND.n86 VGND.n85 34.6358
R3718 VGND.n150 VGND.n149 34.6358
R3719 VGND.n154 VGND.n153 34.6358
R3720 VGND.n1153 VGND.n1135 34.6358
R3721 VGND.n1149 VGND.n1135 34.6358
R3722 VGND.n1149 VGND.n1148 34.6358
R3723 VGND.n1148 VGND.n1147 34.6358
R3724 VGND.n1147 VGND.n1137 34.6358
R3725 VGND.n1131 VGND.n1105 34.6358
R3726 VGND.n1126 VGND.n1106 34.6358
R3727 VGND.n1122 VGND.n1106 34.6358
R3728 VGND.n1122 VGND.n1121 34.6358
R3729 VGND.n1121 VGND.n1120 34.6358
R3730 VGND.n1120 VGND.n1108 34.6358
R3731 VGND.n486 VGND.n481 34.6358
R3732 VGND.n491 VGND.n490 34.6358
R3733 VGND.n2267 VGND.n2262 34.6358
R3734 VGND.n2272 VGND.n2271 34.6358
R3735 VGND.n522 VGND.n517 34.6358
R3736 VGND.n527 VGND.n526 34.6358
R3737 VGND.n2196 VGND.n2195 34.6358
R3738 VGND.n2204 VGND.n2203 34.6358
R3739 VGND.n2200 VGND.n2199 34.6358
R3740 VGND.n2243 VGND.n542 34.6358
R3741 VGND.n2243 VGND.n2242 34.6358
R3742 VGND.n2242 VGND.n2241 34.6358
R3743 VGND.n2241 VGND.n2227 34.6358
R3744 VGND.n2237 VGND.n2227 34.6358
R3745 VGND.n1361 VGND.n1356 34.6358
R3746 VGND.n1381 VGND.n1357 34.6358
R3747 VGND.n1381 VGND.n1380 34.6358
R3748 VGND.n1380 VGND.n1379 34.6358
R3749 VGND.n1379 VGND.n1365 34.6358
R3750 VGND.n1375 VGND.n1365 34.6358
R3751 VGND.n2998 VGND.n2997 34.6358
R3752 VGND.n2 VGND.t1457 34.4422
R3753 VGND.n122 VGND.n121 33.1299
R3754 VGND.n2215 VGND.n544 33.1299
R3755 VGND.n111 VGND.n93 32.377
R3756 VGND.n187 VGND.n186 32.377
R3757 VGND.n111 VGND.n110 32.377
R3758 VGND.n88 VGND.n87 32.377
R3759 VGND.n156 VGND.n155 32.377
R3760 VGND.n2206 VGND.n2205 32.377
R3761 VGND.n2206 VGND.n2184 32.0005
R3762 VGND.n497 VGND.n494 30.4946
R3763 VGND.n2278 VGND.n2275 30.4946
R3764 VGND.n533 VGND.n530 30.4946
R3765 VGND.n190 VGND.n167 29.8709
R3766 VGND.n1143 VGND.n1142 28.9887
R3767 VGND.n1116 VGND.n1115 28.9887
R3768 VGND.n2235 VGND.n2234 28.9887
R3769 VGND.n1373 VGND.n1372 28.9887
R3770 VGND.n2985 VGND.n2984 27.8593
R3771 VGND.n22 VGND.n21 27.8593
R3772 VGND.n2955 VGND.n2954 27.8593
R3773 VGND.n48 VGND.n47 27.8593
R3774 VGND.n2256 VGND.n2255 27.0003
R3775 VGND.n161 VGND.n160 26.8591
R3776 VGND.n184 VGND.n173 26.3534
R3777 VGND.n108 VGND.n98 26.3534
R3778 VGND.n85 VGND.n74 26.3534
R3779 VGND.n153 VGND.n142 26.3534
R3780 VGND.n2203 VGND.n2188 26.3534
R3781 VGND.n129 VGND.n68 25.977
R3782 VGND.n498 VGND.n497 25.977
R3783 VGND.n2279 VGND.n2278 25.977
R3784 VGND.n534 VGND.n533 25.977
R3785 VGND.n509 VGND.n506 25.977
R3786 VGND.n2980 VGND.t2456 24.9236
R3787 VGND.n2980 VGND.t382 24.9236
R3788 VGND.n2979 VGND.t399 24.9236
R3789 VGND.n2979 VGND.t351 24.9236
R3790 VGND.n2977 VGND.t456 24.9236
R3791 VGND.n2977 VGND.t407 24.9236
R3792 VGND.n2976 VGND.t2459 24.9236
R3793 VGND.n2976 VGND.t471 24.9236
R3794 VGND.n17 VGND.t409 24.9236
R3795 VGND.n17 VGND.t450 24.9236
R3796 VGND.n16 VGND.t441 24.9236
R3797 VGND.n16 VGND.t388 24.9236
R3798 VGND.n15 VGND.t400 24.9236
R3799 VGND.n15 VGND.t377 24.9236
R3800 VGND.n14 VGND.t386 24.9236
R3801 VGND.n14 VGND.t461 24.9236
R3802 VGND.n176 VGND.t357 24.9236
R3803 VGND.n176 VGND.t395 24.9236
R3804 VGND.n175 VGND.t403 24.9236
R3805 VGND.n175 VGND.t359 24.9236
R3806 VGND.n172 VGND.t443 24.9236
R3807 VGND.n172 VGND.t1398 24.9236
R3808 VGND.n171 VGND.t2461 24.9236
R3809 VGND.n171 VGND.t1910 24.9236
R3810 VGND.n170 VGND.t1395 24.9236
R3811 VGND.n170 VGND.t1401 24.9236
R3812 VGND.n169 VGND.t1913 24.9236
R3813 VGND.n169 VGND.t1911 24.9236
R3814 VGND.n2950 VGND.t465 24.9236
R3815 VGND.n2950 VGND.t363 24.9236
R3816 VGND.n2949 VGND.t353 24.9236
R3817 VGND.n2949 VGND.t440 24.9236
R3818 VGND.n43 VGND.t379 24.9236
R3819 VGND.n43 VGND.t2462 24.9236
R3820 VGND.n42 VGND.t438 24.9236
R3821 VGND.n42 VGND.t411 24.9236
R3822 VGND.n41 VGND.t474 24.9236
R3823 VGND.n41 VGND.t361 24.9236
R3824 VGND.n40 VGND.t384 24.9236
R3825 VGND.n40 VGND.t460 24.9236
R3826 VGND.n96 VGND.t390 24.9236
R3827 VGND.n96 VGND.t454 24.9236
R3828 VGND.n97 VGND.t413 24.9236
R3829 VGND.n97 VGND.t1558 24.9236
R3830 VGND.n95 VGND.t1554 24.9236
R3831 VGND.n95 VGND.t1548 24.9236
R3832 VGND.n100 VGND.t394 24.9236
R3833 VGND.n100 VGND.t463 24.9236
R3834 VGND.n77 VGND.t473 24.9236
R3835 VGND.n77 VGND.t2457 24.9236
R3836 VGND.n76 VGND.t437 24.9236
R3837 VGND.n76 VGND.t405 24.9236
R3838 VGND.n73 VGND.t396 24.9236
R3839 VGND.n73 VGND.t218 24.9236
R3840 VGND.n72 VGND.t381 24.9236
R3841 VGND.n72 VGND.t1165 24.9236
R3842 VGND.n71 VGND.t214 24.9236
R3843 VGND.n71 VGND.t208 24.9236
R3844 VGND.n70 VGND.t1164 24.9236
R3845 VGND.n70 VGND.t1162 24.9236
R3846 VGND.n145 VGND.t477 24.9236
R3847 VGND.n145 VGND.t2460 24.9236
R3848 VGND.n144 VGND.t459 24.9236
R3849 VGND.n144 VGND.t375 24.9236
R3850 VGND.n141 VGND.t472 24.9236
R3851 VGND.n141 VGND.t659 24.9236
R3852 VGND.n140 VGND.t343 24.9236
R3853 VGND.n140 VGND.t868 24.9236
R3854 VGND.n139 VGND.t656 24.9236
R3855 VGND.n139 VGND.t650 24.9236
R3856 VGND.n138 VGND.t867 24.9236
R3857 VGND.n138 VGND.t869 24.9236
R3858 VGND.n1139 VGND.t1455 24.9236
R3859 VGND.n1139 VGND.t2262 24.9236
R3860 VGND.n1141 VGND.t1440 24.9236
R3861 VGND.n1141 VGND.t2219 24.9236
R3862 VGND.n1111 VGND.t555 24.9236
R3863 VGND.n1111 VGND.t1403 24.9236
R3864 VGND.n1110 VGND.t2254 24.9236
R3865 VGND.n1110 VGND.t2264 24.9236
R3866 VGND.n1114 VGND.t1404 24.9236
R3867 VGND.n1114 VGND.t367 24.9236
R3868 VGND.n1113 VGND.t1441 24.9236
R3869 VGND.n1113 VGND.t601 24.9236
R3870 VGND.n488 VGND.t553 24.9236
R3871 VGND.n488 VGND.t2257 24.9236
R3872 VGND.n487 VGND.t547 24.9236
R3873 VGND.n487 VGND.t1448 24.9236
R3874 VGND.n478 VGND.t2074 24.9236
R3875 VGND.n478 VGND.t552 24.9236
R3876 VGND.n477 VGND.t64 24.9236
R3877 VGND.n477 VGND.t494 24.9236
R3878 VGND.n496 VGND.t2072 24.9236
R3879 VGND.n496 VGND.t2073 24.9236
R3880 VGND.n495 VGND.t67 24.9236
R3881 VGND.n495 VGND.t65 24.9236
R3882 VGND.n2269 VGND.t365 24.9236
R3883 VGND.n2269 VGND.t487 24.9236
R3884 VGND.n2268 VGND.t1433 24.9236
R3885 VGND.n2268 VGND.t2213 24.9236
R3886 VGND.n2259 VGND.t851 24.9236
R3887 VGND.n2259 VGND.t1438 24.9236
R3888 VGND.n2258 VGND.t1710 24.9236
R3889 VGND.n2258 VGND.t2258 24.9236
R3890 VGND.n2277 VGND.t2266 24.9236
R3891 VGND.n2277 VGND.t2267 24.9236
R3892 VGND.n2276 VGND.t2473 24.9236
R3893 VGND.n2276 VGND.t1709 24.9236
R3894 VGND.n524 VGND.t550 24.9236
R3895 VGND.n524 VGND.t1451 24.9236
R3896 VGND.n523 VGND.t490 24.9236
R3897 VGND.n523 VGND.t1406 24.9236
R3898 VGND.n514 VGND.t565 24.9236
R3899 VGND.n514 VGND.t549 24.9236
R3900 VGND.n513 VGND.t1175 24.9236
R3901 VGND.n513 VGND.t486 24.9236
R3902 VGND.n532 VGND.t567 24.9236
R3903 VGND.n532 VGND.t566 24.9236
R3904 VGND.n531 VGND.t1177 24.9236
R3905 VGND.n531 VGND.t1176 24.9236
R3906 VGND.n2186 VGND.t2260 24.9236
R3907 VGND.n2186 VGND.t597 24.9236
R3908 VGND.n2187 VGND.t1299 24.9236
R3909 VGND.n2187 VGND.t1435 24.9236
R3910 VGND.n2185 VGND.t1303 24.9236
R3911 VGND.n2185 VGND.t1301 24.9236
R3912 VGND.n2190 VGND.t1437 24.9236
R3913 VGND.n2190 VGND.t2217 24.9236
R3914 VGND.n2230 VGND.t2255 24.9236
R3915 VGND.n2230 VGND.t2265 24.9236
R3916 VGND.n2229 VGND.t1446 24.9236
R3917 VGND.n2229 VGND.t1449 24.9236
R3918 VGND.n2233 VGND.t1442 24.9236
R3919 VGND.n2233 VGND.t603 24.9236
R3920 VGND.n2231 VGND.t2263 24.9236
R3921 VGND.n2231 VGND.t598 24.9236
R3922 VGND.n1368 VGND.t368 24.9236
R3923 VGND.n1368 VGND.t369 24.9236
R3924 VGND.n1367 VGND.t599 24.9236
R3925 VGND.n1367 VGND.t2214 24.9236
R3926 VGND.n1371 VGND.t595 24.9236
R3927 VGND.n1371 VGND.t554 24.9236
R3928 VGND.n1369 VGND.t489 24.9236
R3929 VGND.n1369 VGND.t1405 24.9236
R3930 VGND.n187 VGND.n166 24.4711
R3931 VGND.n61 VGND.n36 24.4711
R3932 VGND.n123 VGND.n122 24.4711
R3933 VGND.n88 VGND.n67 24.4711
R3934 VGND.n129 VGND.n128 24.4711
R3935 VGND.n156 VGND.n135 24.4711
R3936 VGND.n498 VGND.n474 24.4711
R3937 VGND.n2279 VGND.n2253 24.4711
R3938 VGND.n534 VGND.n505 24.4711
R3939 VGND.n509 VGND.n508 24.4711
R3940 VGND.n2216 VGND.n2215 24.4711
R3941 VGND.n2223 VGND.n541 24.4711
R3942 VGND.n164 VGND.n136 23.7181
R3943 VGND.n2993 VGND.n2972 23.7181
R3944 VGND.n3010 VGND.n9 23.7181
R3945 VGND.n3010 VGND.n10 23.7181
R3946 VGND.n2966 VGND.n2945 23.7181
R3947 VGND.n65 VGND.n35 23.7181
R3948 VGND.n1155 VGND.n1153 23.7181
R3949 VGND.n1127 VGND.n1105 23.7181
R3950 VGND.n1127 VGND.n1126 23.7181
R3951 VGND.n2283 VGND.n2252 23.7181
R3952 VGND.n2210 VGND.n545 23.7181
R3953 VGND.n2247 VGND.n542 23.7181
R3954 VGND.n1385 VGND.n1356 23.7181
R3955 VGND.n1385 VGND.n1357 23.7181
R3956 VGND.n2997 VGND.n2972 23.7181
R3957 VGND.n117 VGND.n115 23.3417
R3958 VGND.n117 VGND.n92 23.3417
R3959 VGND.n2211 VGND.n2210 23.3417
R3960 VGND.n1143 VGND.n1140 21.4593
R3961 VGND.n1116 VGND.n1112 21.4593
R3962 VGND.n2236 VGND.n2235 21.4593
R3963 VGND.n1374 VGND.n1373 21.4593
R3964 VGND.n179 VGND.n178 21.0905
R3965 VGND.n102 VGND.n101 21.0905
R3966 VGND.n80 VGND.n79 21.0905
R3967 VGND.n148 VGND.n147 21.0905
R3968 VGND.n180 VGND.n179 20.3299
R3969 VGND.n103 VGND.n102 20.3299
R3970 VGND.n81 VGND.n80 20.3299
R3971 VGND.n149 VGND.n148 20.3299
R3972 VGND.n494 VGND.n479 19.9534
R3973 VGND.n2275 VGND.n2260 19.9534
R3974 VGND.n530 VGND.n515 19.9534
R3975 VGND.n3006 VGND.n3005 19.2005
R3976 VGND.n61 VGND.n60 19.2005
R3977 VGND.n2223 VGND.n2222 19.2005
R3978 VGND.n1361 VGND.n1360 19.2005
R3979 VGND.t1925 VGND.t326 16.8587
R3980 VGND.t1195 VGND.t328 16.8587
R3981 VGND.t2498 VGND.t2083 16.8587
R3982 VGND.t1133 VGND.t2081 16.8587
R3983 VGND.n1133 VGND.n1132 16.077
R3984 VGND.n3000 VGND.n2999 16.077
R3985 VGND.n60 VGND.n59 15.4358
R3986 VGND.n2222 VGND.n2221 15.4358
R3987 VGND.n3005 VGND.n3004 14.6829
R3988 VGND.n160 VGND.n159 14.6829
R3989 VGND.n2255 VGND.n2254 14.6829
R3990 VGND.n1360 VGND.n1359 14.6829
R3991 VGND.n483 VGND.n482 14.5711
R3992 VGND.n2264 VGND.n2263 14.5711
R3993 VGND.n519 VGND.n518 14.5711
R3994 VGND.n2194 VGND.n2193 14.5711
R3995 VGND.n133 VGND.n68 14.3064
R3996 VGND.n538 VGND.n506 14.3064
R3997 VGND.n490 VGND.n489 13.9299
R3998 VGND.n2271 VGND.n2270 13.9299
R3999 VGND.n526 VGND.n525 13.9299
R4000 VGND.n2199 VGND.n2191 13.9299
R4001 VGND.n65 VGND.n36 13.5534
R4002 VGND.n2247 VGND.n541 13.5534
R4003 VGND.n193 VGND.n166 13.177
R4004 VGND.n133 VGND.n67 13.177
R4005 VGND.n164 VGND.n135 13.177
R4006 VGND.n502 VGND.n474 13.177
R4007 VGND.n2283 VGND.n2253 13.177
R4008 VGND.n538 VGND.n505 13.177
R4009 VGND.n193 VGND.n167 12.8005
R4010 VGND.n502 VGND.n475 12.8005
R4011 VGND.n3023 VGND.t2691 12.5645
R4012 VGND.n1132 VGND.n1131 10.5417
R4013 VGND.n2999 VGND.n2998 10.5417
R4014 VGND.n3004 VGND.n3003 10.0534
R4015 VGND.n1359 VGND.n1358 10.0534
R4016 VGND.n20 VGND.n19 9.3005
R4017 VGND.n21 VGND.n13 9.3005
R4018 VGND.n24 VGND.n23 9.3005
R4019 VGND.n25 VGND.n12 9.3005
R4020 VGND.n27 VGND.n26 9.3005
R4021 VGND.n28 VGND.n11 9.3005
R4022 VGND.n30 VGND.n29 9.3005
R4023 VGND.n31 VGND.n9 9.3005
R4024 VGND.n3008 VGND.n10 9.3005
R4025 VGND.n3007 VGND.n3006 9.3005
R4026 VGND.n3010 VGND.n3009 9.3005
R4027 VGND.n191 VGND.n167 9.3005
R4028 VGND.n180 VGND.n174 9.3005
R4029 VGND.n182 VGND.n181 9.3005
R4030 VGND.n184 VGND.n183 9.3005
R4031 VGND.n185 VGND.n168 9.3005
R4032 VGND.n188 VGND.n187 9.3005
R4033 VGND.n189 VGND.n166 9.3005
R4034 VGND.n193 VGND.n192 9.3005
R4035 VGND.n2953 VGND.n2952 9.3005
R4036 VGND.n2954 VGND.n2948 9.3005
R4037 VGND.n2957 VGND.n2956 9.3005
R4038 VGND.n2958 VGND.n2947 9.3005
R4039 VGND.n2960 VGND.n2959 9.3005
R4040 VGND.n2961 VGND.n2946 9.3005
R4041 VGND.n2963 VGND.n2962 9.3005
R4042 VGND.n2964 VGND.n2945 9.3005
R4043 VGND.n2966 VGND.n2965 9.3005
R4044 VGND.n59 VGND.n58 9.3005
R4045 VGND.n46 VGND.n45 9.3005
R4046 VGND.n47 VGND.n39 9.3005
R4047 VGND.n50 VGND.n49 9.3005
R4048 VGND.n51 VGND.n38 9.3005
R4049 VGND.n53 VGND.n52 9.3005
R4050 VGND.n54 VGND.n37 9.3005
R4051 VGND.n56 VGND.n55 9.3005
R4052 VGND.n57 VGND.n35 9.3005
R4053 VGND.n63 VGND.n36 9.3005
R4054 VGND.n62 VGND.n61 9.3005
R4055 VGND.n65 VGND.n64 9.3005
R4056 VGND.n124 VGND.n123 9.3005
R4057 VGND.n103 VGND.n99 9.3005
R4058 VGND.n106 VGND.n105 9.3005
R4059 VGND.n108 VGND.n107 9.3005
R4060 VGND.n109 VGND.n94 9.3005
R4061 VGND.n112 VGND.n111 9.3005
R4062 VGND.n114 VGND.n113 9.3005
R4063 VGND.n120 VGND.n119 9.3005
R4064 VGND.n122 VGND.n91 9.3005
R4065 VGND.n118 VGND.n117 9.3005
R4066 VGND.n128 VGND.n127 9.3005
R4067 VGND.n81 VGND.n75 9.3005
R4068 VGND.n83 VGND.n82 9.3005
R4069 VGND.n85 VGND.n84 9.3005
R4070 VGND.n86 VGND.n69 9.3005
R4071 VGND.n89 VGND.n88 9.3005
R4072 VGND.n90 VGND.n67 9.3005
R4073 VGND.n131 VGND.n68 9.3005
R4074 VGND.n130 VGND.n129 9.3005
R4075 VGND.n133 VGND.n132 9.3005
R4076 VGND.n162 VGND.n136 9.3005
R4077 VGND.n149 VGND.n143 9.3005
R4078 VGND.n151 VGND.n150 9.3005
R4079 VGND.n153 VGND.n152 9.3005
R4080 VGND.n154 VGND.n137 9.3005
R4081 VGND.n157 VGND.n156 9.3005
R4082 VGND.n158 VGND.n135 9.3005
R4083 VGND.n164 VGND.n163 9.3005
R4084 VGND.n1144 VGND.n1143 9.3005
R4085 VGND.n1145 VGND.n1137 9.3005
R4086 VGND.n1147 VGND.n1146 9.3005
R4087 VGND.n1148 VGND.n1136 9.3005
R4088 VGND.n1150 VGND.n1149 9.3005
R4089 VGND.n1151 VGND.n1135 9.3005
R4090 VGND.n1153 VGND.n1152 9.3005
R4091 VGND.n1156 VGND.n1155 9.3005
R4092 VGND.n1117 VGND.n1116 9.3005
R4093 VGND.n1118 VGND.n1108 9.3005
R4094 VGND.n1120 VGND.n1119 9.3005
R4095 VGND.n1121 VGND.n1107 9.3005
R4096 VGND.n1123 VGND.n1122 9.3005
R4097 VGND.n1124 VGND.n1106 9.3005
R4098 VGND.n1126 VGND.n1125 9.3005
R4099 VGND.n1129 VGND.n1105 9.3005
R4100 VGND.n1131 VGND.n1130 9.3005
R4101 VGND.n1128 VGND.n1127 9.3005
R4102 VGND.n500 VGND.n474 9.3005
R4103 VGND.n484 VGND.n481 9.3005
R4104 VGND.n486 VGND.n485 9.3005
R4105 VGND.n490 VGND.n480 9.3005
R4106 VGND.n492 VGND.n491 9.3005
R4107 VGND.n494 VGND.n493 9.3005
R4108 VGND.n497 VGND.n476 9.3005
R4109 VGND.n499 VGND.n498 9.3005
R4110 VGND.n502 VGND.n501 9.3005
R4111 VGND.n2281 VGND.n2253 9.3005
R4112 VGND.n2265 VGND.n2262 9.3005
R4113 VGND.n2267 VGND.n2266 9.3005
R4114 VGND.n2271 VGND.n2261 9.3005
R4115 VGND.n2273 VGND.n2272 9.3005
R4116 VGND.n2275 VGND.n2274 9.3005
R4117 VGND.n2278 VGND.n2257 9.3005
R4118 VGND.n2280 VGND.n2279 9.3005
R4119 VGND.n2256 VGND.n2252 9.3005
R4120 VGND.n2283 VGND.n2282 9.3005
R4121 VGND.n508 VGND.n507 9.3005
R4122 VGND.n511 VGND.n506 9.3005
R4123 VGND.n536 VGND.n505 9.3005
R4124 VGND.n520 VGND.n517 9.3005
R4125 VGND.n522 VGND.n521 9.3005
R4126 VGND.n526 VGND.n516 9.3005
R4127 VGND.n528 VGND.n527 9.3005
R4128 VGND.n530 VGND.n529 9.3005
R4129 VGND.n533 VGND.n512 9.3005
R4130 VGND.n535 VGND.n534 9.3005
R4131 VGND.n510 VGND.n509 9.3005
R4132 VGND.n538 VGND.n537 9.3005
R4133 VGND.n2217 VGND.n2216 9.3005
R4134 VGND.n2208 VGND.n545 9.3005
R4135 VGND.n2195 VGND.n2192 9.3005
R4136 VGND.n2197 VGND.n2196 9.3005
R4137 VGND.n2199 VGND.n2198 9.3005
R4138 VGND.n2201 VGND.n2200 9.3005
R4139 VGND.n2203 VGND.n2202 9.3005
R4140 VGND.n2204 VGND.n2183 9.3005
R4141 VGND.n2207 VGND.n2206 9.3005
R4142 VGND.n2213 VGND.n2212 9.3005
R4143 VGND.n2215 VGND.n2214 9.3005
R4144 VGND.n2210 VGND.n2209 9.3005
R4145 VGND.n2235 VGND.n2228 9.3005
R4146 VGND.n2238 VGND.n2237 9.3005
R4147 VGND.n2239 VGND.n2227 9.3005
R4148 VGND.n2241 VGND.n2240 9.3005
R4149 VGND.n2242 VGND.n2226 9.3005
R4150 VGND.n2244 VGND.n2243 9.3005
R4151 VGND.n2245 VGND.n542 9.3005
R4152 VGND.n2225 VGND.n541 9.3005
R4153 VGND.n2224 VGND.n2223 9.3005
R4154 VGND.n2221 VGND.n2220 9.3005
R4155 VGND.n2247 VGND.n2246 9.3005
R4156 VGND.n1373 VGND.n1366 9.3005
R4157 VGND.n1376 VGND.n1375 9.3005
R4158 VGND.n1377 VGND.n1365 9.3005
R4159 VGND.n1379 VGND.n1378 9.3005
R4160 VGND.n1380 VGND.n1364 9.3005
R4161 VGND.n1382 VGND.n1381 9.3005
R4162 VGND.n1383 VGND.n1357 9.3005
R4163 VGND.n1363 VGND.n1356 9.3005
R4164 VGND.n1362 VGND.n1361 9.3005
R4165 VGND.n1385 VGND.n1384 9.3005
R4166 VGND.n2982 VGND.n2978 9.3005
R4167 VGND.n2984 VGND.n2983 9.3005
R4168 VGND.n2986 VGND.n2975 9.3005
R4169 VGND.n2988 VGND.n2987 9.3005
R4170 VGND.n2989 VGND.n2974 9.3005
R4171 VGND.n2991 VGND.n2990 9.3005
R4172 VGND.n2992 VGND.n2973 9.3005
R4173 VGND.n2994 VGND.n2993 9.3005
R4174 VGND.n2995 VGND.n2972 9.3005
R4175 VGND.n2997 VGND.n2996 9.3005
R4176 VGND.n2998 VGND.n34 9.3005
R4177 VGND.n181 VGND.n173 8.28285
R4178 VGND.n82 VGND.n74 8.28285
R4179 VGND.n150 VGND.n142 8.28285
R4180 VGND.n2636 VGND.n2635 7.9105
R4181 VGND.n2693 VGND.n337 7.9105
R4182 VGND.n2692 VGND.n338 7.9105
R4183 VGND.n2687 VGND.n343 7.9105
R4184 VGND.n2686 VGND.n344 7.9105
R4185 VGND.n2681 VGND.n349 7.9105
R4186 VGND.n2680 VGND.n350 7.9105
R4187 VGND.n2675 VGND.n2674 7.9105
R4188 VGND.n2712 VGND.n2711 7.9105
R4189 VGND.n2721 VGND.n2720 7.9105
R4190 VGND.n2745 VGND.n2744 7.9105
R4191 VGND.n2759 VGND.n2758 7.9105
R4192 VGND.n2783 VGND.n288 7.9105
R4193 VGND.n2785 VGND.n2784 7.9105
R4194 VGND.n2794 VGND.n2793 7.9105
R4195 VGND.n2937 VGND.n2936 7.9105
R4196 VGND.n2559 VGND.n401 7.9105
R4197 VGND.n2558 VGND.n402 7.9105
R4198 VGND.n2557 VGND.n403 7.9105
R4199 VGND.n2556 VGND.n404 7.9105
R4200 VGND.n2555 VGND.n405 7.9105
R4201 VGND.n2554 VGND.n406 7.9105
R4202 VGND.n2553 VGND.n407 7.9105
R4203 VGND.n2552 VGND.n408 7.9105
R4204 VGND.n2551 VGND.n409 7.9105
R4205 VGND.n2550 VGND.n410 7.9105
R4206 VGND.n2549 VGND.n411 7.9105
R4207 VGND.n2548 VGND.n412 7.9105
R4208 VGND.n2547 VGND.n2546 7.9105
R4209 VGND.n2798 VGND.n282 7.9105
R4210 VGND.n2797 VGND.n283 7.9105
R4211 VGND.n2534 VGND.n2533 7.9105
R4212 VGND.n2357 VGND.n2356 7.9105
R4213 VGND.n2374 VGND.n2373 7.9105
R4214 VGND.n2383 VGND.n2382 7.9105
R4215 VGND.n2400 VGND.n2399 7.9105
R4216 VGND.n2409 VGND.n2408 7.9105
R4217 VGND.n2426 VGND.n2425 7.9105
R4218 VGND.n2435 VGND.n2434 7.9105
R4219 VGND.n2452 VGND.n2451 7.9105
R4220 VGND.n2461 VGND.n2460 7.9105
R4221 VGND.n2478 VGND.n2477 7.9105
R4222 VGND.n2487 VGND.n2486 7.9105
R4223 VGND.n2509 VGND.n2508 7.9105
R4224 VGND.n2802 VGND.n279 7.9105
R4225 VGND.n2801 VGND.n280 7.9105
R4226 VGND.n420 VGND.n419 7.9105
R4227 VGND.n2530 VGND.n2529 7.9105
R4228 VGND.n2361 VGND.n2360 7.9105
R4229 VGND.n2370 VGND.n2369 7.9105
R4230 VGND.n2387 VGND.n2386 7.9105
R4231 VGND.n2396 VGND.n2395 7.9105
R4232 VGND.n2413 VGND.n2412 7.9105
R4233 VGND.n2422 VGND.n2421 7.9105
R4234 VGND.n2439 VGND.n2438 7.9105
R4235 VGND.n2448 VGND.n2447 7.9105
R4236 VGND.n2465 VGND.n2464 7.9105
R4237 VGND.n2474 VGND.n2473 7.9105
R4238 VGND.n2491 VGND.n2490 7.9105
R4239 VGND.n2505 VGND.n2504 7.9105
R4240 VGND.n2805 VGND.n277 7.9105
R4241 VGND.n2807 VGND.n2806 7.9105
R4242 VGND.n2819 VGND.n273 7.9105
R4243 VGND.n2818 VGND.n2817 7.9105
R4244 VGND.n1908 VGND.n1907 7.9105
R4245 VGND.n1917 VGND.n1916 7.9105
R4246 VGND.n1919 VGND.n1918 7.9105
R4247 VGND.n1928 VGND.n1927 7.9105
R4248 VGND.n1930 VGND.n1929 7.9105
R4249 VGND.n1939 VGND.n1938 7.9105
R4250 VGND.n1941 VGND.n1940 7.9105
R4251 VGND.n1950 VGND.n1949 7.9105
R4252 VGND.n1952 VGND.n1951 7.9105
R4253 VGND.n1961 VGND.n1960 7.9105
R4254 VGND.n1963 VGND.n1962 7.9105
R4255 VGND.n1972 VGND.n1971 7.9105
R4256 VGND.n1974 VGND.n1973 7.9105
R4257 VGND.n2823 VGND.n270 7.9105
R4258 VGND.n2822 VGND.n271 7.9105
R4259 VGND.n1990 VGND.n1989 7.9105
R4260 VGND.n2063 VGND.n591 7.9105
R4261 VGND.n2062 VGND.n2061 7.9105
R4262 VGND.n2167 VGND.n556 7.9105
R4263 VGND.n2166 VGND.n557 7.9105
R4264 VGND.n2159 VGND.n562 7.9105
R4265 VGND.n2158 VGND.n563 7.9105
R4266 VGND.n2151 VGND.n568 7.9105
R4267 VGND.n2150 VGND.n569 7.9105
R4268 VGND.n2143 VGND.n574 7.9105
R4269 VGND.n2142 VGND.n575 7.9105
R4270 VGND.n2135 VGND.n580 7.9105
R4271 VGND.n2134 VGND.n581 7.9105
R4272 VGND.n2827 VGND.n267 7.9105
R4273 VGND.n2826 VGND.n268 7.9105
R4274 VGND.n1999 VGND.n1998 7.9105
R4275 VGND.n1997 VGND.n1996 7.9105
R4276 VGND.n2067 VGND.n2066 7.9105
R4277 VGND.n2171 VGND.n553 7.9105
R4278 VGND.n2170 VGND.n554 7.9105
R4279 VGND.n2163 VGND.n559 7.9105
R4280 VGND.n2162 VGND.n560 7.9105
R4281 VGND.n2155 VGND.n565 7.9105
R4282 VGND.n2154 VGND.n566 7.9105
R4283 VGND.n2147 VGND.n571 7.9105
R4284 VGND.n2146 VGND.n572 7.9105
R4285 VGND.n2139 VGND.n577 7.9105
R4286 VGND.n2138 VGND.n578 7.9105
R4287 VGND.n2131 VGND.n2130 7.9105
R4288 VGND.n2830 VGND.n265 7.9105
R4289 VGND.n2832 VGND.n2831 7.9105
R4290 VGND.n2844 VGND.n261 7.9105
R4291 VGND.n2843 VGND.n2842 7.9105
R4292 VGND.n1901 VGND.n548 7.9105
R4293 VGND.n2175 VGND.n2174 7.9105
R4294 VGND.n1759 VGND.n1758 7.9105
R4295 VGND.n1768 VGND.n1767 7.9105
R4296 VGND.n1770 VGND.n1769 7.9105
R4297 VGND.n1779 VGND.n1778 7.9105
R4298 VGND.n1781 VGND.n1780 7.9105
R4299 VGND.n1790 VGND.n1789 7.9105
R4300 VGND.n1792 VGND.n1791 7.9105
R4301 VGND.n1801 VGND.n1800 7.9105
R4302 VGND.n1803 VGND.n1802 7.9105
R4303 VGND.n1812 VGND.n1811 7.9105
R4304 VGND.n1814 VGND.n1813 7.9105
R4305 VGND.n2848 VGND.n258 7.9105
R4306 VGND.n2847 VGND.n259 7.9105
R4307 VGND.n1830 VGND.n1829 7.9105
R4308 VGND.n1899 VGND.n629 7.9105
R4309 VGND.n1685 VGND.n1684 7.9105
R4310 VGND.n1687 VGND.n1686 7.9105
R4311 VGND.n1884 VGND.n643 7.9105
R4312 VGND.n1883 VGND.n644 7.9105
R4313 VGND.n1876 VGND.n649 7.9105
R4314 VGND.n1875 VGND.n650 7.9105
R4315 VGND.n1868 VGND.n655 7.9105
R4316 VGND.n1867 VGND.n656 7.9105
R4317 VGND.n1860 VGND.n661 7.9105
R4318 VGND.n1859 VGND.n662 7.9105
R4319 VGND.n1852 VGND.n1851 7.9105
R4320 VGND.n2852 VGND.n255 7.9105
R4321 VGND.n2851 VGND.n256 7.9105
R4322 VGND.n1839 VGND.n1838 7.9105
R4323 VGND.n1837 VGND.n1836 7.9105
R4324 VGND.n1896 VGND.n633 7.9105
R4325 VGND.n1895 VGND.n634 7.9105
R4326 VGND.n1888 VGND.n640 7.9105
R4327 VGND.n1887 VGND.n641 7.9105
R4328 VGND.n1880 VGND.n646 7.9105
R4329 VGND.n1879 VGND.n647 7.9105
R4330 VGND.n1872 VGND.n652 7.9105
R4331 VGND.n1871 VGND.n653 7.9105
R4332 VGND.n1864 VGND.n658 7.9105
R4333 VGND.n1863 VGND.n659 7.9105
R4334 VGND.n1856 VGND.n664 7.9105
R4335 VGND.n1855 VGND.n730 7.9105
R4336 VGND.n2855 VGND.n253 7.9105
R4337 VGND.n2857 VGND.n2856 7.9105
R4338 VGND.n2869 VGND.n249 7.9105
R4339 VGND.n2868 VGND.n2867 7.9105
R4340 VGND.n1350 VGND.n1349 7.9105
R4341 VGND.n1892 VGND.n636 7.9105
R4342 VGND.n1891 VGND.n637 7.9105
R4343 VGND.n868 VGND.n867 7.9105
R4344 VGND.n866 VGND.n812 7.9105
R4345 VGND.n865 VGND.n813 7.9105
R4346 VGND.n864 VGND.n814 7.9105
R4347 VGND.n863 VGND.n815 7.9105
R4348 VGND.n862 VGND.n816 7.9105
R4349 VGND.n861 VGND.n817 7.9105
R4350 VGND.n860 VGND.n859 7.9105
R4351 VGND.n1669 VGND.n732 7.9105
R4352 VGND.n1668 VGND.n1667 7.9105
R4353 VGND.n2873 VGND.n246 7.9105
R4354 VGND.n2872 VGND.n247 7.9105
R4355 VGND.n1655 VGND.n1654 7.9105
R4356 VGND.n1404 VGND.n801 7.9105
R4357 VGND.n1403 VGND.n802 7.9105
R4358 VGND.n1402 VGND.n1401 7.9105
R4359 VGND.n1488 VGND.n1487 7.9105
R4360 VGND.n1497 VGND.n1496 7.9105
R4361 VGND.n1514 VGND.n1513 7.9105
R4362 VGND.n1523 VGND.n1522 7.9105
R4363 VGND.n1540 VGND.n1539 7.9105
R4364 VGND.n1560 VGND.n758 7.9105
R4365 VGND.n1559 VGND.n1558 7.9105
R4366 VGND.n1628 VGND.n742 7.9105
R4367 VGND.n1630 VGND.n1629 7.9105
R4368 VGND.n2877 VGND.n243 7.9105
R4369 VGND.n2876 VGND.n244 7.9105
R4370 VGND.n741 VGND.n740 7.9105
R4371 VGND.n1651 VGND.n1650 7.9105
R4372 VGND.n1408 VGND.n1407 7.9105
R4373 VGND.n1417 VGND.n1416 7.9105
R4374 VGND.n1475 VGND.n1474 7.9105
R4375 VGND.n1484 VGND.n1483 7.9105
R4376 VGND.n1501 VGND.n1500 7.9105
R4377 VGND.n1510 VGND.n1509 7.9105
R4378 VGND.n1527 VGND.n1526 7.9105
R4379 VGND.n1536 VGND.n1535 7.9105
R4380 VGND.n1564 VGND.n1563 7.9105
R4381 VGND.n1588 VGND.n1587 7.9105
R4382 VGND.n1625 VGND.n744 7.9105
R4383 VGND.n1624 VGND.n745 7.9105
R4384 VGND.n2880 VGND.n240 7.9105
R4385 VGND.n2882 VGND.n2881 7.9105
R4386 VGND.n2894 VGND.n236 7.9105
R4387 VGND.n2893 VGND.n2892 7.9105
R4388 VGND.n1344 VGND.n1343 7.9105
R4389 VGND.n1421 VGND.n1420 7.9105
R4390 VGND.n1471 VGND.n783 7.9105
R4391 VGND.n1470 VGND.n784 7.9105
R4392 VGND.n1469 VGND.n785 7.9105
R4393 VGND.n1468 VGND.n786 7.9105
R4394 VGND.n1467 VGND.n787 7.9105
R4395 VGND.n1466 VGND.n788 7.9105
R4396 VGND.n1465 VGND.n1464 7.9105
R4397 VGND.n1591 VGND.n751 7.9105
R4398 VGND.n1593 VGND.n1592 7.9105
R4399 VGND.n1621 VGND.n747 7.9105
R4400 VGND.n1620 VGND.n1619 7.9105
R4401 VGND.n2898 VGND.n231 7.9105
R4402 VGND.n2897 VGND.n232 7.9105
R4403 VGND.n1607 VGND.n1606 7.9105
R4404 VGND.n1103 VGND.n1025 7.9105
R4405 VGND.n1102 VGND.n1026 7.9105
R4406 VGND.n1101 VGND.n1100 7.9105
R4407 VGND.n1321 VGND.n899 7.9105
R4408 VGND.n1320 VGND.n900 7.9105
R4409 VGND.n1313 VGND.n905 7.9105
R4410 VGND.n1312 VGND.n906 7.9105
R4411 VGND.n1305 VGND.n911 7.9105
R4412 VGND.n1304 VGND.n912 7.9105
R4413 VGND.n1068 VGND.n1067 7.9105
R4414 VGND.n1066 VGND.n1045 7.9105
R4415 VGND.n1065 VGND.n1046 7.9105
R4416 VGND.n1064 VGND.n1063 7.9105
R4417 VGND.n2902 VGND.n2901 7.9105
R4418 VGND.n233 VGND.n228 7.9105
R4419 VGND.n2913 VGND.n2912 7.9105
R4420 VGND.n1161 VGND.n888 7.9105
R4421 VGND.n1331 VGND.n1330 7.9105
R4422 VGND.n1325 VGND.n896 7.9105
R4423 VGND.n1324 VGND.n897 7.9105
R4424 VGND.n1317 VGND.n902 7.9105
R4425 VGND.n1316 VGND.n903 7.9105
R4426 VGND.n1309 VGND.n908 7.9105
R4427 VGND.n1308 VGND.n909 7.9105
R4428 VGND.n1301 VGND.n914 7.9105
R4429 VGND.n1300 VGND.n915 7.9105
R4430 VGND.n1295 VGND.n919 7.9105
R4431 VGND.n1294 VGND.n920 7.9105
R4432 VGND.n1289 VGND.n924 7.9105
R4433 VGND.n1288 VGND.n925 7.9105
R4434 VGND.n1287 VGND.n992 7.9105
R4435 VGND.n2917 VGND.n2916 7.9105
R4436 VGND.n489 VGND.n486 7.90638
R4437 VGND.n482 VGND.n481 7.90638
R4438 VGND.n2270 VGND.n2267 7.90638
R4439 VGND.n2263 VGND.n2262 7.90638
R4440 VGND.n525 VGND.n522 7.90638
R4441 VGND.n518 VGND.n517 7.90638
R4442 VGND.n2196 VGND.n2191 7.90638
R4443 VGND.n2195 VGND.n2194 7.90638
R4444 VGND.n1142 VGND.n1138 7.4049
R4445 VGND.n1115 VGND.n1109 7.4049
R4446 VGND.n2234 VGND.n2232 7.4049
R4447 VGND.n1372 VGND.n1370 7.4049
R4448 VGND VGND.n475 7.12482
R4449 VGND.n178 VGND.n177 6.85473
R4450 VGND.n79 VGND.n78 6.85473
R4451 VGND.n147 VGND.n146 6.85473
R4452 VGND.n2986 VGND.n2985 6.77697
R4453 VGND.n23 VGND.n22 6.77697
R4454 VGND.n2956 VGND.n2955 6.77697
R4455 VGND.n49 VGND.n48 6.77697
R4456 VGND.n3022 VGND.n3021 6.4005
R4457 VGND.n104 VGND.n98 5.27109
R4458 VGND.n2189 VGND.n2188 5.27109
R4459 VGND.n2565 VGND.n2564 4.5005
R4460 VGND.n2568 VGND.n2567 4.5005
R4461 VGND.n2571 VGND.n2570 4.5005
R4462 VGND.n2574 VGND.n2573 4.5005
R4463 VGND.n2577 VGND.n2576 4.5005
R4464 VGND.n2580 VGND.n2579 4.5005
R4465 VGND.n2583 VGND.n2582 4.5005
R4466 VGND.n2586 VGND.n2585 4.5005
R4467 VGND.n2589 VGND.n2588 4.5005
R4468 VGND.n2592 VGND.n2591 4.5005
R4469 VGND.n2595 VGND.n2594 4.5005
R4470 VGND.n2598 VGND.n2597 4.5005
R4471 VGND.n2601 VGND.n2600 4.5005
R4472 VGND.n2604 VGND.n2603 4.5005
R4473 VGND.n2607 VGND.n2606 4.5005
R4474 VGND.n335 VGND.n334 4.5005
R4475 VGND.n2627 VGND.n2626 4.5005
R4476 VGND.n2624 VGND.n2623 4.5005
R4477 VGND.n2621 VGND.n2620 4.5005
R4478 VGND.n2618 VGND.n2617 4.5005
R4479 VGND.n2615 VGND.n2614 4.5005
R4480 VGND.n2612 VGND.n2611 4.5005
R4481 VGND.n323 VGND.n322 4.5005
R4482 VGND.n316 VGND.n315 4.5005
R4483 VGND.n307 VGND.n306 4.5005
R4484 VGND.n2763 VGND.n299 4.5005
R4485 VGND.n2766 VGND.n2765 4.5005
R4486 VGND.n291 VGND.n290 4.5005
R4487 VGND.n2770 VGND.n297 4.5005
R4488 VGND.n205 VGND.n204 4.5005
R4489 VGND.n2631 VGND.n2630 4.5005
R4490 VGND.n2632 VGND.n331 4.5005
R4491 VGND.n2697 VGND.n2696 4.5005
R4492 VGND.n358 VGND.n340 4.5005
R4493 VGND.n365 VGND.n341 4.5005
R4494 VGND.n354 VGND.n346 4.5005
R4495 VGND.n376 VGND.n347 4.5005
R4496 VGND.n353 VGND.n352 4.5005
R4497 VGND.n390 VGND.n389 4.5005
R4498 VGND.n2708 VGND.n2707 4.5005
R4499 VGND.n2725 VGND.n2724 4.5005
R4500 VGND.n2741 VGND.n2740 4.5005
R4501 VGND.n2762 VGND.n300 4.5005
R4502 VGND.n2733 VGND.n289 4.5005
R4503 VGND.n2779 VGND.n2778 4.5005
R4504 VGND.n2772 VGND.n2771 4.5005
R4505 VGND.n2942 VGND.n2941 4.5005
R4506 VGND.n1019 VGND.n1018 4.5005
R4507 VGND.n1016 VGND.n1015 4.5005
R4508 VGND.n1181 VGND.n1180 4.5005
R4509 VGND.n1193 VGND.n1006 4.5005
R4510 VGND.n1200 VGND.n1004 4.5005
R4511 VGND.n1197 VGND.n1195 4.5005
R4512 VGND.n1213 VGND.n1212 4.5005
R4513 VGND.n1251 VGND.n1000 4.5005
R4514 VGND.n1254 VGND.n1253 4.5005
R4515 VGND.n1257 VGND.n1256 4.5005
R4516 VGND.n1260 VGND.n1259 4.5005
R4517 VGND.n1263 VGND.n1262 4.5005
R4518 VGND.n1269 VGND.n998 4.5005
R4519 VGND.n1266 VGND.n1265 4.5005
R4520 VGND.n995 VGND.n994 4.5005
R4521 VGND.n1022 VGND.n1021 4.5005
R4522 VGND.n1165 VGND.n1164 4.5005
R4523 VGND.n1170 VGND.n891 4.5005
R4524 VGND.n1011 VGND.n892 4.5005
R4525 VGND.n1183 VGND.n1182 4.5005
R4526 VGND.n1192 VGND.n1191 4.5005
R4527 VGND.n1202 VGND.n1201 4.5005
R4528 VGND.n1196 VGND.n1003 4.5005
R4529 VGND.n1215 VGND.n1214 4.5005
R4530 VGND.n1250 VGND.n1249 4.5005
R4531 VGND.n1223 VGND.n916 4.5005
R4532 VGND.n1242 VGND.n917 4.5005
R4533 VGND.n1228 VGND.n921 4.5005
R4534 VGND.n1235 VGND.n922 4.5005
R4535 VGND.n1272 VGND.n1271 4.5005
R4536 VGND.n997 VGND.n993 4.5005
R4537 VGND.n1283 VGND.n1282 4.5005
R4538 VGND.n1157 VGND.n1156 4.41365
R4539 VGND VGND.n33 4.35375
R4540 VGND.n1134 VGND.n1133 4.05427
R4541 VGND.n507 VGND.n0 4.05427
R4542 VGND.n2218 VGND.n2217 4.05427
R4543 VGND.n2220 VGND.n2219 4.05427
R4544 VGND.n1358 VGND.n543 4.05427
R4545 VGND VGND.n3002 3.99438
R4546 VGND VGND.n32 3.99438
R4547 VGND.n125 VGND 3.99438
R4548 VGND VGND.n126 3.99438
R4549 VGND.n3001 VGND 3.99437
R4550 VGND.n1284 VGND.n223 3.77268
R4551 VGND.n2940 VGND.n206 3.77268
R4552 VGND.n1163 VGND.n1162 3.77268
R4553 VGND.n2634 VGND.n2633 3.77268
R4554 VGND.n1327 VGND.n1326 3.77268
R4555 VGND.n2691 VGND.n2690 3.77268
R4556 VGND.n1323 VGND.n898 3.77268
R4557 VGND.n2689 VGND.n2688 3.77268
R4558 VGND.n1318 VGND.n901 3.77268
R4559 VGND.n2685 VGND.n2684 3.77268
R4560 VGND.n1315 VGND.n904 3.77268
R4561 VGND.n2683 VGND.n2682 3.77268
R4562 VGND.n1310 VGND.n907 3.77268
R4563 VGND.n2679 VGND.n2678 3.77268
R4564 VGND.n1307 VGND.n910 3.77268
R4565 VGND.n2677 VGND.n2676 3.77268
R4566 VGND.n1302 VGND.n913 3.77268
R4567 VGND.n2710 VGND.n2709 3.77268
R4568 VGND.n1299 VGND.n1298 3.77268
R4569 VGND.n2723 VGND.n2722 3.77268
R4570 VGND.n1297 VGND.n1296 3.77268
R4571 VGND.n2743 VGND.n2742 3.77268
R4572 VGND.n1293 VGND.n1292 3.77268
R4573 VGND.n2761 VGND.n2760 3.77268
R4574 VGND.n1291 VGND.n1290 3.77268
R4575 VGND.n2782 VGND.n2781 3.77268
R4576 VGND.n1270 VGND.n229 3.77268
R4577 VGND.n2780 VGND.n281 3.77268
R4578 VGND.n1286 VGND.n1285 3.77268
R4579 VGND.n2795 VGND.n284 3.77268
R4580 VGND.n1329 VGND.n1328 3.77268
R4581 VGND.n2695 VGND.n2694 3.77268
R4582 VGND.n2769 VGND.n205 3.75914
R4583 VGND.n2631 VGND.n2629 3.75914
R4584 VGND.n1267 VGND.n995 3.75914
R4585 VGND.n1022 VGND.n1020 3.75914
R4586 VGND.n2771 VGND.n284 3.4105
R4587 VGND.n2780 VGND.n2779 3.4105
R4588 VGND.n2781 VGND.n289 3.4105
R4589 VGND.n2762 VGND.n2761 3.4105
R4590 VGND.n2742 VGND.n2741 3.4105
R4591 VGND.n2724 VGND.n2723 3.4105
R4592 VGND.n2709 VGND.n2708 3.4105
R4593 VGND.n2677 VGND.n390 3.4105
R4594 VGND.n2678 VGND.n352 3.4105
R4595 VGND.n2683 VGND.n347 3.4105
R4596 VGND.n2684 VGND.n346 3.4105
R4597 VGND.n2689 VGND.n341 3.4105
R4598 VGND.n2690 VGND.n340 3.4105
R4599 VGND.n2696 VGND.n2695 3.4105
R4600 VGND.n2941 VGND.n2940 3.4105
R4601 VGND.n2770 VGND.n2769 3.4105
R4602 VGND.n2768 VGND.n291 3.4105
R4603 VGND.n2767 VGND.n2766 3.4105
R4604 VGND.n2764 VGND.n2763 3.4105
R4605 VGND.n307 VGND.n298 3.4105
R4606 VGND.n2609 VGND.n316 3.4105
R4607 VGND.n2610 VGND.n323 3.4105
R4608 VGND.n2613 VGND.n2612 3.4105
R4609 VGND.n2616 VGND.n2615 3.4105
R4610 VGND.n2619 VGND.n2618 3.4105
R4611 VGND.n2622 VGND.n2621 3.4105
R4612 VGND.n2625 VGND.n2624 3.4105
R4613 VGND.n2628 VGND.n2627 3.4105
R4614 VGND.n2629 VGND.n335 3.4105
R4615 VGND.n2633 VGND.n2632 3.4105
R4616 VGND.n2937 VGND.n206 3.4105
R4617 VGND.n2635 VGND.n2634 3.4105
R4618 VGND.n2559 VGND.n397 3.4105
R4619 VGND.n2533 VGND.n2532 3.4105
R4620 VGND.n2557 VGND.n339 3.4105
R4621 VGND.n2692 VGND.n2691 3.4105
R4622 VGND.n2384 VGND.n2383 3.4105
R4623 VGND.n2358 VGND.n2357 3.4105
R4624 VGND.n2531 VGND.n2530 3.4105
R4625 VGND.n2399 VGND.n2398 3.4105
R4626 VGND.n2556 VGND.n342 3.4105
R4627 VGND.n2688 VGND.n2687 3.4105
R4628 VGND.n2397 VGND.n2396 3.4105
R4629 VGND.n2386 VGND.n2385 3.4105
R4630 VGND.n2360 VGND.n2359 3.4105
R4631 VGND.n2818 VGND.n274 3.4105
R4632 VGND.n2412 VGND.n2411 3.4105
R4633 VGND.n2410 VGND.n2409 3.4105
R4634 VGND.n2555 VGND.n345 3.4105
R4635 VGND.n2686 VGND.n2685 3.4105
R4636 VGND.n1929 VGND.n449 3.4105
R4637 VGND.n1928 VGND.n453 3.4105
R4638 VGND.n1918 VGND.n457 3.4105
R4639 VGND.n1907 VGND.n467 3.4105
R4640 VGND.n1990 VGND.n604 3.4105
R4641 VGND.n1939 VGND.n445 3.4105
R4642 VGND.n2423 VGND.n2422 3.4105
R4643 VGND.n2425 VGND.n2424 3.4105
R4644 VGND.n2554 VGND.n348 3.4105
R4645 VGND.n2682 VGND.n2681 3.4105
R4646 VGND.n2158 VGND.n2157 3.4105
R4647 VGND.n2160 VGND.n2159 3.4105
R4648 VGND.n2166 VGND.n2165 3.4105
R4649 VGND.n2168 VGND.n2167 3.4105
R4650 VGND.n2064 VGND.n2063 3.4105
R4651 VGND.n1997 VGND.n603 3.4105
R4652 VGND.n2152 VGND.n2151 3.4105
R4653 VGND.n1940 VGND.n441 3.4105
R4654 VGND.n2438 VGND.n2437 3.4105
R4655 VGND.n2436 VGND.n2435 3.4105
R4656 VGND.n2553 VGND.n351 3.4105
R4657 VGND.n2680 VGND.n2679 3.4105
R4658 VGND.n2154 VGND.n2153 3.4105
R4659 VGND.n2156 VGND.n2155 3.4105
R4660 VGND.n2162 VGND.n2161 3.4105
R4661 VGND.n2164 VGND.n2163 3.4105
R4662 VGND.n2170 VGND.n2169 3.4105
R4663 VGND.n2066 VGND.n2065 3.4105
R4664 VGND.n2843 VGND.n262 3.4105
R4665 VGND.n2148 VGND.n2147 3.4105
R4666 VGND.n2150 VGND.n2149 3.4105
R4667 VGND.n1950 VGND.n437 3.4105
R4668 VGND.n2449 VGND.n2448 3.4105
R4669 VGND.n2451 VGND.n2450 3.4105
R4670 VGND.n2552 VGND.n391 3.4105
R4671 VGND.n2676 VGND.n2675 3.4105
R4672 VGND.n1790 VGND.n570 3.4105
R4673 VGND.n1780 VGND.n567 3.4105
R4674 VGND.n1779 VGND.n564 3.4105
R4675 VGND.n1769 VGND.n561 3.4105
R4676 VGND.n1768 VGND.n558 3.4105
R4677 VGND.n1758 VGND.n555 3.4105
R4678 VGND.n1901 VGND.n588 3.4105
R4679 VGND.n1830 VGND.n1737 3.4105
R4680 VGND.n1791 VGND.n573 3.4105
R4681 VGND.n2146 VGND.n2145 3.4105
R4682 VGND.n2144 VGND.n2143 3.4105
R4683 VGND.n1951 VGND.n433 3.4105
R4684 VGND.n2464 VGND.n2463 3.4105
R4685 VGND.n2462 VGND.n2461 3.4105
R4686 VGND.n2551 VGND.n321 3.4105
R4687 VGND.n2711 VGND.n2710 3.4105
R4688 VGND.n1867 VGND.n1866 3.4105
R4689 VGND.n1869 VGND.n1868 3.4105
R4690 VGND.n1875 VGND.n1874 3.4105
R4691 VGND.n1877 VGND.n1876 3.4105
R4692 VGND.n1883 VGND.n1882 3.4105
R4693 VGND.n1885 VGND.n1884 3.4105
R4694 VGND.n1686 VGND.n639 3.4105
R4695 VGND.n1899 VGND.n1898 3.4105
R4696 VGND.n1837 VGND.n1736 3.4105
R4697 VGND.n1861 VGND.n1860 3.4105
R4698 VGND.n1801 VGND.n576 3.4105
R4699 VGND.n2140 VGND.n2139 3.4105
R4700 VGND.n2142 VGND.n2141 3.4105
R4701 VGND.n1961 VGND.n429 3.4105
R4702 VGND.n2475 VGND.n2474 3.4105
R4703 VGND.n2477 VGND.n2476 3.4105
R4704 VGND.n2550 VGND.n317 3.4105
R4705 VGND.n2722 VGND.n2721 3.4105
R4706 VGND.n1863 VGND.n1862 3.4105
R4707 VGND.n1865 VGND.n1864 3.4105
R4708 VGND.n1871 VGND.n1870 3.4105
R4709 VGND.n1873 VGND.n1872 3.4105
R4710 VGND.n1879 VGND.n1878 3.4105
R4711 VGND.n1881 VGND.n1880 3.4105
R4712 VGND.n1887 VGND.n1886 3.4105
R4713 VGND.n1889 VGND.n1888 3.4105
R4714 VGND.n1897 VGND.n1896 3.4105
R4715 VGND.n2868 VGND.n250 3.4105
R4716 VGND.n1857 VGND.n1856 3.4105
R4717 VGND.n1859 VGND.n1858 3.4105
R4718 VGND.n1802 VGND.n579 3.4105
R4719 VGND.n2138 VGND.n2137 3.4105
R4720 VGND.n2136 VGND.n2135 3.4105
R4721 VGND.n1962 VGND.n425 3.4105
R4722 VGND.n2490 VGND.n2489 3.4105
R4723 VGND.n2488 VGND.n2487 3.4105
R4724 VGND.n2549 VGND.n305 3.4105
R4725 VGND.n2744 VGND.n2743 3.4105
R4726 VGND.n860 VGND.n663 3.4105
R4727 VGND.n861 VGND.n660 3.4105
R4728 VGND.n862 VGND.n657 3.4105
R4729 VGND.n863 VGND.n654 3.4105
R4730 VGND.n864 VGND.n651 3.4105
R4731 VGND.n865 VGND.n648 3.4105
R4732 VGND.n866 VGND.n645 3.4105
R4733 VGND.n867 VGND.n642 3.4105
R4734 VGND.n1891 VGND.n1890 3.4105
R4735 VGND.n1349 VGND.n630 3.4105
R4736 VGND.n1654 VGND.n737 3.4105
R4737 VGND.n1670 VGND.n1669 3.4105
R4738 VGND.n1855 VGND.n1854 3.4105
R4739 VGND.n1853 VGND.n1852 3.4105
R4740 VGND.n1812 VGND.n582 3.4105
R4741 VGND.n2132 VGND.n2131 3.4105
R4742 VGND.n2134 VGND.n2133 3.4105
R4743 VGND.n1972 VGND.n421 3.4105
R4744 VGND.n2506 VGND.n2505 3.4105
R4745 VGND.n2508 VGND.n2507 3.4105
R4746 VGND.n2548 VGND.n301 3.4105
R4747 VGND.n2760 VGND.n2759 3.4105
R4748 VGND.n1629 VGND.n731 3.4105
R4749 VGND.n1628 VGND.n1627 3.4105
R4750 VGND.n1559 VGND.n753 3.4105
R4751 VGND.n1561 VGND.n1560 3.4105
R4752 VGND.n1539 VGND.n1538 3.4105
R4753 VGND.n1524 VGND.n1523 3.4105
R4754 VGND.n1513 VGND.n1512 3.4105
R4755 VGND.n1498 VGND.n1497 3.4105
R4756 VGND.n1487 VGND.n1486 3.4105
R4757 VGND.n1402 VGND.n638 3.4105
R4758 VGND.n1405 VGND.n1404 3.4105
R4759 VGND.n1651 VGND.n738 3.4105
R4760 VGND.n2878 VGND.n2877 3.4105
R4761 VGND.n1668 VGND.n242 3.4105
R4762 VGND.n2855 VGND.n2854 3.4105
R4763 VGND.n2853 VGND.n2852 3.4105
R4764 VGND.n1813 VGND.n254 3.4105
R4765 VGND.n2830 VGND.n2829 3.4105
R4766 VGND.n2828 VGND.n2827 3.4105
R4767 VGND.n1973 VGND.n266 3.4105
R4768 VGND.n2805 VGND.n2804 3.4105
R4769 VGND.n2803 VGND.n2802 3.4105
R4770 VGND.n2547 VGND.n278 3.4105
R4771 VGND.n2783 VGND.n2782 3.4105
R4772 VGND.n2880 VGND.n2879 3.4105
R4773 VGND.n1624 VGND.n1623 3.4105
R4774 VGND.n1626 VGND.n1625 3.4105
R4775 VGND.n1589 VGND.n1588 3.4105
R4776 VGND.n1563 VGND.n1562 3.4105
R4777 VGND.n1537 VGND.n1536 3.4105
R4778 VGND.n1526 VGND.n1525 3.4105
R4779 VGND.n1511 VGND.n1510 3.4105
R4780 VGND.n1500 VGND.n1499 3.4105
R4781 VGND.n1485 VGND.n1484 3.4105
R4782 VGND.n1474 VGND.n1473 3.4105
R4783 VGND.n1407 VGND.n1406 3.4105
R4784 VGND.n2893 VGND.n237 3.4105
R4785 VGND.n2881 VGND.n230 3.4105
R4786 VGND.n2876 VGND.n2875 3.4105
R4787 VGND.n2874 VGND.n2873 3.4105
R4788 VGND.n2856 VGND.n245 3.4105
R4789 VGND.n2851 VGND.n2850 3.4105
R4790 VGND.n2849 VGND.n2848 3.4105
R4791 VGND.n2831 VGND.n257 3.4105
R4792 VGND.n2826 VGND.n2825 3.4105
R4793 VGND.n2824 VGND.n2823 3.4105
R4794 VGND.n2806 VGND.n269 3.4105
R4795 VGND.n2801 VGND.n2800 3.4105
R4796 VGND.n2799 VGND.n2798 3.4105
R4797 VGND.n2784 VGND.n281 3.4105
R4798 VGND.n2899 VGND.n2898 3.4105
R4799 VGND.n1620 VGND.n241 3.4105
R4800 VGND.n1622 VGND.n1621 3.4105
R4801 VGND.n1592 VGND.n743 3.4105
R4802 VGND.n1591 VGND.n1590 3.4105
R4803 VGND.n1465 VGND.n757 3.4105
R4804 VGND.n1466 VGND.n762 3.4105
R4805 VGND.n1467 VGND.n766 3.4105
R4806 VGND.n1468 VGND.n770 3.4105
R4807 VGND.n1469 VGND.n774 3.4105
R4808 VGND.n1470 VGND.n778 3.4105
R4809 VGND.n1472 VGND.n1471 3.4105
R4810 VGND.n1344 VGND.n798 3.4105
R4811 VGND.n1606 VGND.n1605 3.4105
R4812 VGND.n2897 VGND.n2896 3.4105
R4813 VGND.n2895 VGND.n2894 3.4105
R4814 VGND.n740 VGND.n235 3.4105
R4815 VGND.n2872 VGND.n2871 3.4105
R4816 VGND.n2870 VGND.n2869 3.4105
R4817 VGND.n1838 VGND.n248 3.4105
R4818 VGND.n2847 VGND.n2846 3.4105
R4819 VGND.n2845 VGND.n2844 3.4105
R4820 VGND.n1998 VGND.n260 3.4105
R4821 VGND.n2822 VGND.n2821 3.4105
R4822 VGND.n2820 VGND.n2819 3.4105
R4823 VGND.n419 VGND.n272 3.4105
R4824 VGND.n2797 VGND.n2796 3.4105
R4825 VGND.n2795 VGND.n2794 3.4105
R4826 VGND.n234 VGND.n233 3.4105
R4827 VGND.n2901 VGND.n2900 3.4105
R4828 VGND.n1064 VGND.n923 3.4105
R4829 VGND.n1065 VGND.n746 3.4105
R4830 VGND.n1066 VGND.n918 3.4105
R4831 VGND.n1067 VGND.n752 3.4105
R4832 VGND.n1304 VGND.n1303 3.4105
R4833 VGND.n1306 VGND.n1305 3.4105
R4834 VGND.n1312 VGND.n1311 3.4105
R4835 VGND.n1314 VGND.n1313 3.4105
R4836 VGND.n1320 VGND.n1319 3.4105
R4837 VGND.n1322 VGND.n1321 3.4105
R4838 VGND.n1101 VGND.n782 3.4105
R4839 VGND.n1104 VGND.n1103 3.4105
R4840 VGND.n2913 VGND.n226 3.4105
R4841 VGND.n1102 VGND.n792 3.4105
R4842 VGND.n1420 VGND.n1419 3.4105
R4843 VGND.n1418 VGND.n1417 3.4105
R4844 VGND.n1403 VGND.n635 3.4105
R4845 VGND.n1893 VGND.n1892 3.4105
R4846 VGND.n1895 VGND.n1894 3.4105
R4847 VGND.n1685 VGND.n551 3.4105
R4848 VGND.n2174 VGND.n2173 3.4105
R4849 VGND.n2172 VGND.n2171 3.4105
R4850 VGND.n2062 VGND.n552 3.4105
R4851 VGND.n1917 VGND.n461 3.4105
R4852 VGND.n2371 VGND.n2370 3.4105
R4853 VGND.n2373 VGND.n2372 3.4105
R4854 VGND.n2558 VGND.n336 3.4105
R4855 VGND.n2694 VGND.n2693 3.4105
R4856 VGND.n1285 VGND.n993 3.4105
R4857 VGND.n1271 VGND.n1270 3.4105
R4858 VGND.n1291 VGND.n922 3.4105
R4859 VGND.n1292 VGND.n921 3.4105
R4860 VGND.n1297 VGND.n917 3.4105
R4861 VGND.n1298 VGND.n916 3.4105
R4862 VGND.n1250 VGND.n913 3.4105
R4863 VGND.n1214 VGND.n910 3.4105
R4864 VGND.n1196 VGND.n907 3.4105
R4865 VGND.n1201 VGND.n904 3.4105
R4866 VGND.n1192 VGND.n901 3.4105
R4867 VGND.n1182 VGND.n898 3.4105
R4868 VGND.n1327 VGND.n892 3.4105
R4869 VGND.n1328 VGND.n891 3.4105
R4870 VGND.n1284 VGND.n1283 3.4105
R4871 VGND.n1267 VGND.n1266 3.4105
R4872 VGND.n1269 VGND.n1268 3.4105
R4873 VGND.n1264 VGND.n1263 3.4105
R4874 VGND.n1261 VGND.n1260 3.4105
R4875 VGND.n1258 VGND.n1257 3.4105
R4876 VGND.n1255 VGND.n1254 3.4105
R4877 VGND.n1252 VGND.n1251 3.4105
R4878 VGND.n1213 VGND.n999 3.4105
R4879 VGND.n1198 VGND.n1197 3.4105
R4880 VGND.n1200 VGND.n1199 3.4105
R4881 VGND.n1194 VGND.n1193 3.4105
R4882 VGND.n1181 VGND.n1005 3.4105
R4883 VGND.n1017 VGND.n1016 3.4105
R4884 VGND.n1020 VGND.n1019 3.4105
R4885 VGND.n1164 VGND.n1163 3.4105
R4886 VGND.n1287 VGND.n1286 3.4105
R4887 VGND.n1288 VGND.n229 3.4105
R4888 VGND.n1290 VGND.n1289 3.4105
R4889 VGND.n1294 VGND.n1293 3.4105
R4890 VGND.n1296 VGND.n1295 3.4105
R4891 VGND.n1300 VGND.n1299 3.4105
R4892 VGND.n1302 VGND.n1301 3.4105
R4893 VGND.n1308 VGND.n1307 3.4105
R4894 VGND.n1310 VGND.n1309 3.4105
R4895 VGND.n1316 VGND.n1315 3.4105
R4896 VGND.n1318 VGND.n1317 3.4105
R4897 VGND.n1324 VGND.n1323 3.4105
R4898 VGND.n1326 VGND.n1325 3.4105
R4899 VGND.n1330 VGND.n1329 3.4105
R4900 VGND.n1162 VGND.n1161 3.4105
R4901 VGND.n2916 VGND.n223 3.4105
R4902 VGND.n105 VGND.n104 3.01226
R4903 VGND.n2200 VGND.n2189 3.01226
R4904 VGND.n2184 VGND.n545 2.63579
R4905 VGND.n2565 VGND 2.52282
R4906 VGND.n2568 VGND 2.52282
R4907 VGND.n2571 VGND 2.52282
R4908 VGND.n2574 VGND 2.52282
R4909 VGND.n2577 VGND 2.52282
R4910 VGND.n2580 VGND 2.52282
R4911 VGND.n2583 VGND 2.52282
R4912 VGND.n2586 VGND 2.52282
R4913 VGND.n2589 VGND 2.52282
R4914 VGND.n2592 VGND 2.52282
R4915 VGND.n2595 VGND 2.52282
R4916 VGND.n2598 VGND 2.52282
R4917 VGND.n2601 VGND 2.52282
R4918 VGND.n2604 VGND 2.52282
R4919 VGND.n2607 VGND 2.52282
R4920 VGND.n186 VGND.n185 2.25932
R4921 VGND.n114 VGND.n93 2.25932
R4922 VGND.n110 VGND.n109 2.25932
R4923 VGND.n87 VGND.n86 2.25932
R4924 VGND.n155 VGND.n154 2.25932
R4925 VGND.n2205 VGND.n2204 2.25932
R4926 VGND.n491 VGND.n479 1.88285
R4927 VGND.n2272 VGND.n2260 1.88285
R4928 VGND.n527 VGND.n515 1.88285
R4929 VGND.n2608 VGND 1.79514
R4930 VGND.n1158 VGND.n224 1.76378
R4931 VGND.n2608 VGND 1.57193
R4932 VGND.n2940 VGND.n2939 1.54254
R4933 VGND.n2938 VGND.n2937 1.54254
R4934 VGND.n2533 VGND.n207 1.54254
R4935 VGND.n2530 VGND.n417 1.54254
R4936 VGND.n2818 VGND.n275 1.54254
R4937 VGND.n1991 VGND.n1990 1.54254
R4938 VGND.n1997 VGND.n1992 1.54254
R4939 VGND.n2843 VGND.n263 1.54254
R4940 VGND.n1831 VGND.n1830 1.54254
R4941 VGND.n1837 VGND.n1832 1.54254
R4942 VGND.n2868 VGND.n251 1.54254
R4943 VGND.n1654 VGND.n1653 1.54254
R4944 VGND.n1652 VGND.n1651 1.54254
R4945 VGND.n2893 VGND.n238 1.54254
R4946 VGND.n1606 VGND.n225 1.54254
R4947 VGND.n2914 VGND.n2913 1.54254
R4948 VGND.n1284 VGND.n224 1.54254
R4949 VGND.n2916 VGND.n2915 1.54254
R4950 VGND.n121 VGND.n120 1.50638
R4951 VGND.n2212 VGND.n544 1.50638
R4952 VGND VGND.n2562 1.3946
R4953 VGND.n2561 VGND 1.3946
R4954 VGND.n2560 VGND 1.3946
R4955 VGND VGND.n398 1.3946
R4956 VGND.n1905 VGND 1.3946
R4957 VGND VGND.n1906 1.3946
R4958 VGND.n1904 VGND 1.3946
R4959 VGND.n1903 VGND 1.3946
R4960 VGND.n1902 VGND 1.3946
R4961 VGND.n1900 VGND 1.3946
R4962 VGND VGND.n626 1.3946
R4963 VGND VGND.n1348 1.3946
R4964 VGND.n1347 VGND 1.3946
R4965 VGND.n1346 VGND 1.3946
R4966 VGND.n1345 VGND 1.3946
R4967 VGND VGND.n880 1.3946
R4968 VGND.n1159 VGND 1.3946
R4969 VGND VGND.n1160 1.3946
R4970 VGND.n1158 VGND.n1157 1.04899
R4971 VGND.n2696 VGND.n335 1.00149
R4972 VGND.n2627 VGND.n340 1.00149
R4973 VGND.n2624 VGND.n341 1.00149
R4974 VGND.n2621 VGND.n346 1.00149
R4975 VGND.n2618 VGND.n347 1.00149
R4976 VGND.n2615 VGND.n352 1.00149
R4977 VGND.n2612 VGND.n390 1.00149
R4978 VGND.n2708 VGND.n323 1.00149
R4979 VGND.n2724 VGND.n316 1.00149
R4980 VGND.n2741 VGND.n307 1.00149
R4981 VGND.n2763 VGND.n2762 1.00149
R4982 VGND.n2766 VGND.n289 1.00149
R4983 VGND.n2779 VGND.n291 1.00149
R4984 VGND.n2771 VGND.n2770 1.00149
R4985 VGND.n2941 VGND.n205 1.00149
R4986 VGND.n1019 VGND.n891 1.00149
R4987 VGND.n1016 VGND.n892 1.00149
R4988 VGND.n1182 VGND.n1181 1.00149
R4989 VGND.n1193 VGND.n1192 1.00149
R4990 VGND.n1201 VGND.n1200 1.00149
R4991 VGND.n1197 VGND.n1196 1.00149
R4992 VGND.n1214 VGND.n1213 1.00149
R4993 VGND.n1251 VGND.n1250 1.00149
R4994 VGND.n1254 VGND.n916 1.00149
R4995 VGND.n1257 VGND.n917 1.00149
R4996 VGND.n1260 VGND.n921 1.00149
R4997 VGND.n1263 VGND.n922 1.00149
R4998 VGND.n1271 VGND.n1269 1.00149
R4999 VGND.n1266 VGND.n993 1.00149
R5000 VGND.n1283 VGND.n995 1.00149
R5001 VGND.n1164 VGND.n1022 1.00149
R5002 VGND.n2632 VGND.n2631 0.973133
R5003 VGND.n2346 VGND.n2 0.9305
R5004 VGND.n178 VGND.n174 0.929432
R5005 VGND.n101 VGND.n99 0.929432
R5006 VGND.n79 VGND.n75 0.929432
R5007 VGND.n147 VGND.n143 0.929432
R5008 VGND.n126 VGND.n1 0.916608
R5009 VGND VGND.n2565 0.839786
R5010 VGND VGND.n2568 0.839786
R5011 VGND VGND.n2571 0.839786
R5012 VGND VGND.n2574 0.839786
R5013 VGND VGND.n2577 0.839786
R5014 VGND VGND.n2580 0.839786
R5015 VGND VGND.n2583 0.839786
R5016 VGND VGND.n2586 0.839786
R5017 VGND VGND.n2589 0.839786
R5018 VGND VGND.n2592 0.839786
R5019 VGND VGND.n2595 0.839786
R5020 VGND VGND.n2598 0.839786
R5021 VGND VGND.n2601 0.839786
R5022 VGND VGND.n2604 0.839786
R5023 VGND VGND.n2607 0.839786
R5024 VGND.n3023 VGND.n3022 0.7755
R5025 VGND.n3024 VGND.n3023 0.774207
R5026 VGND.n2981 VGND.n2978 0.753441
R5027 VGND.n20 VGND.n18 0.753441
R5028 VGND.n2953 VGND.n2951 0.753441
R5029 VGND.n46 VGND.n44 0.753441
R5030 VGND.n159 VGND.n136 0.753441
R5031 VGND.n2254 VGND.n2252 0.753441
R5032 VGND.n3025 VGND 0.706681
R5033 VGND VGND.n0 0.542567
R5034 VGND.n3025 VGND.n1 0.507317
R5035 VGND.n2939 VGND.n33 0.404308
R5036 VGND.n115 VGND.n114 0.376971
R5037 VGND.n120 VGND.n92 0.376971
R5038 VGND.n1140 VGND.n1137 0.376971
R5039 VGND.n1112 VGND.n1108 0.376971
R5040 VGND.n2212 VGND.n2211 0.376971
R5041 VGND.n2237 VGND.n2236 0.376971
R5042 VGND.n1375 VGND.n1374 0.376971
R5043 VGND VGND.n3025 0.37415
R5044 VGND.n226 VGND.n223 0.362676
R5045 VGND.n1605 VGND.n226 0.362676
R5046 VGND.n1605 VGND.n237 0.362676
R5047 VGND.n738 VGND.n237 0.362676
R5048 VGND.n738 VGND.n737 0.362676
R5049 VGND.n737 VGND.n250 0.362676
R5050 VGND.n1736 VGND.n250 0.362676
R5051 VGND.n1737 VGND.n1736 0.362676
R5052 VGND.n1737 VGND.n262 0.362676
R5053 VGND.n603 VGND.n262 0.362676
R5054 VGND.n604 VGND.n603 0.362676
R5055 VGND.n604 VGND.n274 0.362676
R5056 VGND.n2531 VGND.n274 0.362676
R5057 VGND.n2532 VGND.n2531 0.362676
R5058 VGND.n2532 VGND.n206 0.362676
R5059 VGND.n1162 VGND.n1104 0.362676
R5060 VGND.n1104 VGND.n798 0.362676
R5061 VGND.n1406 VGND.n798 0.362676
R5062 VGND.n1406 VGND.n1405 0.362676
R5063 VGND.n1405 VGND.n630 0.362676
R5064 VGND.n1897 VGND.n630 0.362676
R5065 VGND.n1898 VGND.n1897 0.362676
R5066 VGND.n1898 VGND.n588 0.362676
R5067 VGND.n2065 VGND.n588 0.362676
R5068 VGND.n2065 VGND.n2064 0.362676
R5069 VGND.n2064 VGND.n467 0.362676
R5070 VGND.n2359 VGND.n467 0.362676
R5071 VGND.n2359 VGND.n2358 0.362676
R5072 VGND.n2358 VGND.n397 0.362676
R5073 VGND.n2634 VGND.n397 0.362676
R5074 VGND.n1326 VGND.n782 0.362676
R5075 VGND.n1472 VGND.n782 0.362676
R5076 VGND.n1473 VGND.n1472 0.362676
R5077 VGND.n1473 VGND.n638 0.362676
R5078 VGND.n1890 VGND.n638 0.362676
R5079 VGND.n1890 VGND.n1889 0.362676
R5080 VGND.n1889 VGND.n639 0.362676
R5081 VGND.n639 VGND.n555 0.362676
R5082 VGND.n2169 VGND.n555 0.362676
R5083 VGND.n2169 VGND.n2168 0.362676
R5084 VGND.n2168 VGND.n457 0.362676
R5085 VGND.n2385 VGND.n457 0.362676
R5086 VGND.n2385 VGND.n2384 0.362676
R5087 VGND.n2384 VGND.n339 0.362676
R5088 VGND.n2691 VGND.n339 0.362676
R5089 VGND.n1323 VGND.n1322 0.362676
R5090 VGND.n1322 VGND.n778 0.362676
R5091 VGND.n1485 VGND.n778 0.362676
R5092 VGND.n1486 VGND.n1485 0.362676
R5093 VGND.n1486 VGND.n642 0.362676
R5094 VGND.n1886 VGND.n642 0.362676
R5095 VGND.n1886 VGND.n1885 0.362676
R5096 VGND.n1885 VGND.n558 0.362676
R5097 VGND.n2164 VGND.n558 0.362676
R5098 VGND.n2165 VGND.n2164 0.362676
R5099 VGND.n2165 VGND.n453 0.362676
R5100 VGND.n2397 VGND.n453 0.362676
R5101 VGND.n2398 VGND.n2397 0.362676
R5102 VGND.n2398 VGND.n342 0.362676
R5103 VGND.n2688 VGND.n342 0.362676
R5104 VGND.n1319 VGND.n1318 0.362676
R5105 VGND.n1319 VGND.n774 0.362676
R5106 VGND.n1499 VGND.n774 0.362676
R5107 VGND.n1499 VGND.n1498 0.362676
R5108 VGND.n1498 VGND.n645 0.362676
R5109 VGND.n1881 VGND.n645 0.362676
R5110 VGND.n1882 VGND.n1881 0.362676
R5111 VGND.n1882 VGND.n561 0.362676
R5112 VGND.n2161 VGND.n561 0.362676
R5113 VGND.n2161 VGND.n2160 0.362676
R5114 VGND.n2160 VGND.n449 0.362676
R5115 VGND.n2411 VGND.n449 0.362676
R5116 VGND.n2411 VGND.n2410 0.362676
R5117 VGND.n2410 VGND.n345 0.362676
R5118 VGND.n2685 VGND.n345 0.362676
R5119 VGND.n1315 VGND.n1314 0.362676
R5120 VGND.n1314 VGND.n770 0.362676
R5121 VGND.n1511 VGND.n770 0.362676
R5122 VGND.n1512 VGND.n1511 0.362676
R5123 VGND.n1512 VGND.n648 0.362676
R5124 VGND.n1878 VGND.n648 0.362676
R5125 VGND.n1878 VGND.n1877 0.362676
R5126 VGND.n1877 VGND.n564 0.362676
R5127 VGND.n2156 VGND.n564 0.362676
R5128 VGND.n2157 VGND.n2156 0.362676
R5129 VGND.n2157 VGND.n445 0.362676
R5130 VGND.n2423 VGND.n445 0.362676
R5131 VGND.n2424 VGND.n2423 0.362676
R5132 VGND.n2424 VGND.n348 0.362676
R5133 VGND.n2682 VGND.n348 0.362676
R5134 VGND.n1311 VGND.n1310 0.362676
R5135 VGND.n1311 VGND.n766 0.362676
R5136 VGND.n1525 VGND.n766 0.362676
R5137 VGND.n1525 VGND.n1524 0.362676
R5138 VGND.n1524 VGND.n651 0.362676
R5139 VGND.n1873 VGND.n651 0.362676
R5140 VGND.n1874 VGND.n1873 0.362676
R5141 VGND.n1874 VGND.n567 0.362676
R5142 VGND.n2153 VGND.n567 0.362676
R5143 VGND.n2153 VGND.n2152 0.362676
R5144 VGND.n2152 VGND.n441 0.362676
R5145 VGND.n2437 VGND.n441 0.362676
R5146 VGND.n2437 VGND.n2436 0.362676
R5147 VGND.n2436 VGND.n351 0.362676
R5148 VGND.n2679 VGND.n351 0.362676
R5149 VGND.n1307 VGND.n1306 0.362676
R5150 VGND.n1306 VGND.n762 0.362676
R5151 VGND.n1537 VGND.n762 0.362676
R5152 VGND.n1538 VGND.n1537 0.362676
R5153 VGND.n1538 VGND.n654 0.362676
R5154 VGND.n1870 VGND.n654 0.362676
R5155 VGND.n1870 VGND.n1869 0.362676
R5156 VGND.n1869 VGND.n570 0.362676
R5157 VGND.n2148 VGND.n570 0.362676
R5158 VGND.n2149 VGND.n2148 0.362676
R5159 VGND.n2149 VGND.n437 0.362676
R5160 VGND.n2449 VGND.n437 0.362676
R5161 VGND.n2450 VGND.n2449 0.362676
R5162 VGND.n2450 VGND.n391 0.362676
R5163 VGND.n2676 VGND.n391 0.362676
R5164 VGND.n1303 VGND.n1302 0.362676
R5165 VGND.n1303 VGND.n757 0.362676
R5166 VGND.n1562 VGND.n757 0.362676
R5167 VGND.n1562 VGND.n1561 0.362676
R5168 VGND.n1561 VGND.n657 0.362676
R5169 VGND.n1865 VGND.n657 0.362676
R5170 VGND.n1866 VGND.n1865 0.362676
R5171 VGND.n1866 VGND.n573 0.362676
R5172 VGND.n2145 VGND.n573 0.362676
R5173 VGND.n2145 VGND.n2144 0.362676
R5174 VGND.n2144 VGND.n433 0.362676
R5175 VGND.n2463 VGND.n433 0.362676
R5176 VGND.n2463 VGND.n2462 0.362676
R5177 VGND.n2462 VGND.n321 0.362676
R5178 VGND.n2710 VGND.n321 0.362676
R5179 VGND.n1299 VGND.n752 0.362676
R5180 VGND.n1590 VGND.n752 0.362676
R5181 VGND.n1590 VGND.n1589 0.362676
R5182 VGND.n1589 VGND.n753 0.362676
R5183 VGND.n753 VGND.n660 0.362676
R5184 VGND.n1862 VGND.n660 0.362676
R5185 VGND.n1862 VGND.n1861 0.362676
R5186 VGND.n1861 VGND.n576 0.362676
R5187 VGND.n2140 VGND.n576 0.362676
R5188 VGND.n2141 VGND.n2140 0.362676
R5189 VGND.n2141 VGND.n429 0.362676
R5190 VGND.n2475 VGND.n429 0.362676
R5191 VGND.n2476 VGND.n2475 0.362676
R5192 VGND.n2476 VGND.n317 0.362676
R5193 VGND.n2722 VGND.n317 0.362676
R5194 VGND.n1296 VGND.n918 0.362676
R5195 VGND.n918 VGND.n743 0.362676
R5196 VGND.n1626 VGND.n743 0.362676
R5197 VGND.n1627 VGND.n1626 0.362676
R5198 VGND.n1627 VGND.n663 0.362676
R5199 VGND.n1857 VGND.n663 0.362676
R5200 VGND.n1858 VGND.n1857 0.362676
R5201 VGND.n1858 VGND.n579 0.362676
R5202 VGND.n2137 VGND.n579 0.362676
R5203 VGND.n2137 VGND.n2136 0.362676
R5204 VGND.n2136 VGND.n425 0.362676
R5205 VGND.n2489 VGND.n425 0.362676
R5206 VGND.n2489 VGND.n2488 0.362676
R5207 VGND.n2488 VGND.n305 0.362676
R5208 VGND.n2743 VGND.n305 0.362676
R5209 VGND.n1293 VGND.n746 0.362676
R5210 VGND.n1622 VGND.n746 0.362676
R5211 VGND.n1623 VGND.n1622 0.362676
R5212 VGND.n1623 VGND.n731 0.362676
R5213 VGND.n1670 VGND.n731 0.362676
R5214 VGND.n1854 VGND.n1670 0.362676
R5215 VGND.n1854 VGND.n1853 0.362676
R5216 VGND.n1853 VGND.n582 0.362676
R5217 VGND.n2132 VGND.n582 0.362676
R5218 VGND.n2133 VGND.n2132 0.362676
R5219 VGND.n2133 VGND.n421 0.362676
R5220 VGND.n2506 VGND.n421 0.362676
R5221 VGND.n2507 VGND.n2506 0.362676
R5222 VGND.n2507 VGND.n301 0.362676
R5223 VGND.n2760 VGND.n301 0.362676
R5224 VGND.n1290 VGND.n923 0.362676
R5225 VGND.n923 VGND.n241 0.362676
R5226 VGND.n2879 VGND.n241 0.362676
R5227 VGND.n2879 VGND.n2878 0.362676
R5228 VGND.n2878 VGND.n242 0.362676
R5229 VGND.n2854 VGND.n242 0.362676
R5230 VGND.n2854 VGND.n2853 0.362676
R5231 VGND.n2853 VGND.n254 0.362676
R5232 VGND.n2829 VGND.n254 0.362676
R5233 VGND.n2829 VGND.n2828 0.362676
R5234 VGND.n2828 VGND.n266 0.362676
R5235 VGND.n2804 VGND.n266 0.362676
R5236 VGND.n2804 VGND.n2803 0.362676
R5237 VGND.n2803 VGND.n278 0.362676
R5238 VGND.n2782 VGND.n278 0.362676
R5239 VGND.n2900 VGND.n229 0.362676
R5240 VGND.n2900 VGND.n2899 0.362676
R5241 VGND.n2899 VGND.n230 0.362676
R5242 VGND.n2875 VGND.n230 0.362676
R5243 VGND.n2875 VGND.n2874 0.362676
R5244 VGND.n2874 VGND.n245 0.362676
R5245 VGND.n2850 VGND.n245 0.362676
R5246 VGND.n2850 VGND.n2849 0.362676
R5247 VGND.n2849 VGND.n257 0.362676
R5248 VGND.n2825 VGND.n257 0.362676
R5249 VGND.n2825 VGND.n2824 0.362676
R5250 VGND.n2824 VGND.n269 0.362676
R5251 VGND.n2800 VGND.n269 0.362676
R5252 VGND.n2800 VGND.n2799 0.362676
R5253 VGND.n2799 VGND.n281 0.362676
R5254 VGND.n1286 VGND.n234 0.362676
R5255 VGND.n2896 VGND.n234 0.362676
R5256 VGND.n2896 VGND.n2895 0.362676
R5257 VGND.n2895 VGND.n235 0.362676
R5258 VGND.n2871 VGND.n235 0.362676
R5259 VGND.n2871 VGND.n2870 0.362676
R5260 VGND.n2870 VGND.n248 0.362676
R5261 VGND.n2846 VGND.n248 0.362676
R5262 VGND.n2846 VGND.n2845 0.362676
R5263 VGND.n2845 VGND.n260 0.362676
R5264 VGND.n2821 VGND.n260 0.362676
R5265 VGND.n2821 VGND.n2820 0.362676
R5266 VGND.n2820 VGND.n272 0.362676
R5267 VGND.n2796 VGND.n272 0.362676
R5268 VGND.n2796 VGND.n2795 0.362676
R5269 VGND.n1329 VGND.n792 0.362676
R5270 VGND.n1419 VGND.n792 0.362676
R5271 VGND.n1419 VGND.n1418 0.362676
R5272 VGND.n1418 VGND.n635 0.362676
R5273 VGND.n1893 VGND.n635 0.362676
R5274 VGND.n1894 VGND.n1893 0.362676
R5275 VGND.n1894 VGND.n551 0.362676
R5276 VGND.n2173 VGND.n551 0.362676
R5277 VGND.n2173 VGND.n2172 0.362676
R5278 VGND.n2172 VGND.n552 0.362676
R5279 VGND.n552 VGND.n461 0.362676
R5280 VGND.n2371 VGND.n461 0.362676
R5281 VGND.n2372 VGND.n2371 0.362676
R5282 VGND.n2372 VGND.n336 0.362676
R5283 VGND.n2694 VGND.n336 0.362676
R5284 VGND.n2769 VGND.n2768 0.349144
R5285 VGND.n2768 VGND.n2767 0.349144
R5286 VGND.n2767 VGND.n2764 0.349144
R5287 VGND.n2764 VGND.n298 0.349144
R5288 VGND.n2609 VGND.n298 0.349144
R5289 VGND.n2610 VGND.n2609 0.349144
R5290 VGND.n2613 VGND.n2610 0.349144
R5291 VGND.n2616 VGND.n2613 0.349144
R5292 VGND.n2619 VGND.n2616 0.349144
R5293 VGND.n2622 VGND.n2619 0.349144
R5294 VGND.n2625 VGND.n2622 0.349144
R5295 VGND.n2628 VGND.n2625 0.349144
R5296 VGND.n2629 VGND.n2628 0.349144
R5297 VGND.n1268 VGND.n1267 0.349144
R5298 VGND.n1268 VGND.n1264 0.349144
R5299 VGND.n1264 VGND.n1261 0.349144
R5300 VGND.n1261 VGND.n1258 0.349144
R5301 VGND.n1258 VGND.n1255 0.349144
R5302 VGND.n1255 VGND.n1252 0.349144
R5303 VGND.n1252 VGND.n999 0.349144
R5304 VGND.n1198 VGND.n999 0.349144
R5305 VGND.n1199 VGND.n1198 0.349144
R5306 VGND.n1199 VGND.n1194 0.349144
R5307 VGND.n1194 VGND.n1005 0.349144
R5308 VGND.n1017 VGND.n1005 0.349144
R5309 VGND.n1020 VGND.n1017 0.349144
R5310 VGND.n2700 VGND.n331 0.327628
R5311 VGND.n2697 VGND.n333 0.327628
R5312 VGND.n361 VGND.n358 0.327628
R5313 VGND.n369 VGND.n365 0.327628
R5314 VGND.n372 VGND.n354 0.327628
R5315 VGND.n380 VGND.n376 0.327628
R5316 VGND.n383 VGND.n353 0.327628
R5317 VGND.n389 VGND.n388 0.327628
R5318 VGND.n2707 VGND.n2706 0.327628
R5319 VGND.n2727 VGND.n2725 0.327628
R5320 VGND.n2740 VGND.n2739 0.327628
R5321 VGND.n2736 VGND.n300 0.327628
R5322 VGND.n2733 VGND.n2732 0.327628
R5323 VGND.n2778 VGND.n2777 0.327628
R5324 VGND.n2774 VGND.n2772 0.327628
R5325 VGND.n2793 VGND.n2792 0.327628
R5326 VGND.n2789 VGND.n2785 0.327628
R5327 VGND.n2754 VGND.n288 0.327628
R5328 VGND.n2758 VGND.n2757 0.327628
R5329 VGND.n2749 VGND.n2745 0.327628
R5330 VGND.n2720 VGND.n2719 0.327628
R5331 VGND.n2716 VGND.n2712 0.327628
R5332 VGND.n2674 VGND.n2673 0.327628
R5333 VGND.n2670 VGND.n350 0.327628
R5334 VGND.n2665 VGND.n349 0.327628
R5335 VGND.n2660 VGND.n344 0.327628
R5336 VGND.n2655 VGND.n343 0.327628
R5337 VGND.n2650 VGND.n338 0.327628
R5338 VGND.n2645 VGND.n337 0.327628
R5339 VGND.n2640 VGND.n2636 0.327628
R5340 VGND.n2537 VGND.n283 0.327628
R5341 VGND.n2542 VGND.n282 0.327628
R5342 VGND.n2546 VGND.n2545 0.327628
R5343 VGND.n2289 VGND.n412 0.327628
R5344 VGND.n2294 VGND.n411 0.327628
R5345 VGND.n2299 VGND.n410 0.327628
R5346 VGND.n2304 VGND.n409 0.327628
R5347 VGND.n2309 VGND.n408 0.327628
R5348 VGND.n2314 VGND.n407 0.327628
R5349 VGND.n2319 VGND.n406 0.327628
R5350 VGND.n2324 VGND.n405 0.327628
R5351 VGND.n2329 VGND.n404 0.327628
R5352 VGND.n2334 VGND.n403 0.327628
R5353 VGND.n2339 VGND.n402 0.327628
R5354 VGND.n2344 VGND.n401 0.327628
R5355 VGND.n2526 VGND.n420 0.327628
R5356 VGND.n2523 VGND.n280 0.327628
R5357 VGND.n2518 VGND.n279 0.327628
R5358 VGND.n2513 VGND.n2509 0.327628
R5359 VGND.n2486 VGND.n2485 0.327628
R5360 VGND.n2482 VGND.n2478 0.327628
R5361 VGND.n2460 VGND.n2459 0.327628
R5362 VGND.n2456 VGND.n2452 0.327628
R5363 VGND.n2434 VGND.n2433 0.327628
R5364 VGND.n2430 VGND.n2426 0.327628
R5365 VGND.n2408 VGND.n2407 0.327628
R5366 VGND.n2404 VGND.n2400 0.327628
R5367 VGND.n2382 VGND.n2381 0.327628
R5368 VGND.n2378 VGND.n2374 0.327628
R5369 VGND.n2356 VGND.n2355 0.327628
R5370 VGND.n2814 VGND.n273 0.327628
R5371 VGND.n2811 VGND.n2807 0.327628
R5372 VGND.n2500 VGND.n277 0.327628
R5373 VGND.n2504 VGND.n2503 0.327628
R5374 VGND.n2495 VGND.n2491 0.327628
R5375 VGND.n2473 VGND.n2472 0.327628
R5376 VGND.n2469 VGND.n2465 0.327628
R5377 VGND.n2447 VGND.n2446 0.327628
R5378 VGND.n2443 VGND.n2439 0.327628
R5379 VGND.n2421 VGND.n2420 0.327628
R5380 VGND.n2417 VGND.n2413 0.327628
R5381 VGND.n2395 VGND.n2394 0.327628
R5382 VGND.n2391 VGND.n2387 0.327628
R5383 VGND.n2369 VGND.n2368 0.327628
R5384 VGND.n2365 VGND.n2361 0.327628
R5385 VGND.n1986 VGND.n271 0.327628
R5386 VGND.n1983 VGND.n270 0.327628
R5387 VGND.n1978 VGND.n1974 0.327628
R5388 VGND.n1971 VGND.n1970 0.327628
R5389 VGND.n1967 VGND.n1963 0.327628
R5390 VGND.n1960 VGND.n1959 0.327628
R5391 VGND.n1956 VGND.n1952 0.327628
R5392 VGND.n1949 VGND.n1948 0.327628
R5393 VGND.n1945 VGND.n1941 0.327628
R5394 VGND.n1938 VGND.n1937 0.327628
R5395 VGND.n1934 VGND.n1930 0.327628
R5396 VGND.n1927 VGND.n1926 0.327628
R5397 VGND.n1923 VGND.n1919 0.327628
R5398 VGND.n1916 VGND.n1915 0.327628
R5399 VGND.n1912 VGND.n1908 0.327628
R5400 VGND.n1999 VGND.n602 0.327628
R5401 VGND.n2002 VGND.n268 0.327628
R5402 VGND.n2007 VGND.n267 0.327628
R5403 VGND.n2012 VGND.n581 0.327628
R5404 VGND.n2017 VGND.n580 0.327628
R5405 VGND.n2022 VGND.n575 0.327628
R5406 VGND.n2027 VGND.n574 0.327628
R5407 VGND.n2032 VGND.n569 0.327628
R5408 VGND.n2037 VGND.n568 0.327628
R5409 VGND.n2042 VGND.n563 0.327628
R5410 VGND.n2047 VGND.n562 0.327628
R5411 VGND.n2052 VGND.n557 0.327628
R5412 VGND.n2057 VGND.n556 0.327628
R5413 VGND.n2061 VGND.n2060 0.327628
R5414 VGND.n598 VGND.n591 0.327628
R5415 VGND.n2839 VGND.n261 0.327628
R5416 VGND.n2836 VGND.n2832 0.327628
R5417 VGND.n2126 VGND.n265 0.327628
R5418 VGND.n2130 VGND.n2129 0.327628
R5419 VGND.n2121 VGND.n578 0.327628
R5420 VGND.n2116 VGND.n577 0.327628
R5421 VGND.n2111 VGND.n572 0.327628
R5422 VGND.n2106 VGND.n571 0.327628
R5423 VGND.n2101 VGND.n566 0.327628
R5424 VGND.n2096 VGND.n565 0.327628
R5425 VGND.n2091 VGND.n560 0.327628
R5426 VGND.n2086 VGND.n559 0.327628
R5427 VGND.n2081 VGND.n554 0.327628
R5428 VGND.n2076 VGND.n553 0.327628
R5429 VGND.n2071 VGND.n2067 0.327628
R5430 VGND.n1826 VGND.n259 0.327628
R5431 VGND.n1823 VGND.n258 0.327628
R5432 VGND.n1818 VGND.n1814 0.327628
R5433 VGND.n1811 VGND.n1810 0.327628
R5434 VGND.n1807 VGND.n1803 0.327628
R5435 VGND.n1800 VGND.n1799 0.327628
R5436 VGND.n1796 VGND.n1792 0.327628
R5437 VGND.n1789 VGND.n1788 0.327628
R5438 VGND.n1785 VGND.n1781 0.327628
R5439 VGND.n1778 VGND.n1777 0.327628
R5440 VGND.n1774 VGND.n1770 0.327628
R5441 VGND.n1767 VGND.n1766 0.327628
R5442 VGND.n1763 VGND.n1759 0.327628
R5443 VGND.n2175 VGND.n550 0.327628
R5444 VGND.n2178 VGND.n548 0.327628
R5445 VGND.n1839 VGND.n1735 0.327628
R5446 VGND.n1842 VGND.n256 0.327628
R5447 VGND.n1847 VGND.n255 0.327628
R5448 VGND.n1851 VGND.n1850 0.327628
R5449 VGND.n1731 VGND.n662 0.327628
R5450 VGND.n1726 VGND.n661 0.327628
R5451 VGND.n1721 VGND.n656 0.327628
R5452 VGND.n1716 VGND.n655 0.327628
R5453 VGND.n1711 VGND.n650 0.327628
R5454 VGND.n1706 VGND.n649 0.327628
R5455 VGND.n1701 VGND.n644 0.327628
R5456 VGND.n1696 VGND.n643 0.327628
R5457 VGND.n1691 VGND.n1687 0.327628
R5458 VGND.n1684 VGND.n1683 0.327628
R5459 VGND.n1680 VGND.n629 0.327628
R5460 VGND.n2864 VGND.n249 0.327628
R5461 VGND.n2861 VGND.n2857 0.327628
R5462 VGND.n726 VGND.n253 0.327628
R5463 VGND.n730 VGND.n729 0.327628
R5464 VGND.n721 VGND.n664 0.327628
R5465 VGND.n716 VGND.n659 0.327628
R5466 VGND.n711 VGND.n658 0.327628
R5467 VGND.n706 VGND.n653 0.327628
R5468 VGND.n701 VGND.n652 0.327628
R5469 VGND.n696 VGND.n647 0.327628
R5470 VGND.n691 VGND.n646 0.327628
R5471 VGND.n686 VGND.n641 0.327628
R5472 VGND.n681 VGND.n640 0.327628
R5473 VGND.n676 VGND.n634 0.327628
R5474 VGND.n671 VGND.n633 0.327628
R5475 VGND.n1658 VGND.n247 0.327628
R5476 VGND.n1663 VGND.n246 0.327628
R5477 VGND.n1667 VGND.n1666 0.327628
R5478 VGND.n855 VGND.n732 0.327628
R5479 VGND.n859 VGND.n858 0.327628
R5480 VGND.n850 VGND.n817 0.327628
R5481 VGND.n845 VGND.n816 0.327628
R5482 VGND.n840 VGND.n815 0.327628
R5483 VGND.n835 VGND.n814 0.327628
R5484 VGND.n830 VGND.n813 0.327628
R5485 VGND.n825 VGND.n812 0.327628
R5486 VGND.n868 VGND.n808 0.327628
R5487 VGND.n871 VGND.n637 0.327628
R5488 VGND.n876 VGND.n636 0.327628
R5489 VGND.n1354 VGND.n1350 0.327628
R5490 VGND.n1647 VGND.n741 0.327628
R5491 VGND.n1644 VGND.n244 0.327628
R5492 VGND.n1639 VGND.n243 0.327628
R5493 VGND.n1634 VGND.n1630 0.327628
R5494 VGND.n1554 VGND.n742 0.327628
R5495 VGND.n1558 VGND.n1557 0.327628
R5496 VGND.n1549 VGND.n758 0.327628
R5497 VGND.n1544 VGND.n1540 0.327628
R5498 VGND.n1522 VGND.n1521 0.327628
R5499 VGND.n1518 VGND.n1514 0.327628
R5500 VGND.n1496 VGND.n1495 0.327628
R5501 VGND.n1492 VGND.n1488 0.327628
R5502 VGND.n1401 VGND.n1400 0.327628
R5503 VGND.n1397 VGND.n802 0.327628
R5504 VGND.n1392 VGND.n801 0.327628
R5505 VGND.n2889 VGND.n236 0.327628
R5506 VGND.n2886 VGND.n2882 0.327628
R5507 VGND.n1573 VGND.n240 0.327628
R5508 VGND.n1578 VGND.n745 0.327628
R5509 VGND.n1583 VGND.n744 0.327628
R5510 VGND.n1587 VGND.n1586 0.327628
R5511 VGND.n1568 VGND.n1564 0.327628
R5512 VGND.n1535 VGND.n1534 0.327628
R5513 VGND.n1531 VGND.n1527 0.327628
R5514 VGND.n1509 VGND.n1508 0.327628
R5515 VGND.n1505 VGND.n1501 0.327628
R5516 VGND.n1483 VGND.n1482 0.327628
R5517 VGND.n1479 VGND.n1475 0.327628
R5518 VGND.n1416 VGND.n1415 0.327628
R5519 VGND.n1412 VGND.n1408 0.327628
R5520 VGND.n1610 VGND.n232 0.327628
R5521 VGND.n1615 VGND.n231 0.327628
R5522 VGND.n1619 VGND.n1618 0.327628
R5523 VGND.n1602 VGND.n747 0.327628
R5524 VGND.n1597 VGND.n1593 0.327628
R5525 VGND.n1460 VGND.n751 0.327628
R5526 VGND.n1464 VGND.n1463 0.327628
R5527 VGND.n1455 VGND.n788 0.327628
R5528 VGND.n1450 VGND.n787 0.327628
R5529 VGND.n1445 VGND.n786 0.327628
R5530 VGND.n1440 VGND.n785 0.327628
R5531 VGND.n1435 VGND.n784 0.327628
R5532 VGND.n1430 VGND.n783 0.327628
R5533 VGND.n1425 VGND.n1421 0.327628
R5534 VGND.n1343 VGND.n1342 0.327628
R5535 VGND.n2909 VGND.n228 0.327628
R5536 VGND.n2906 VGND.n2902 0.327628
R5537 VGND.n1063 VGND.n1062 0.327628
R5538 VGND.n1059 VGND.n1046 0.327628
R5539 VGND.n1054 VGND.n1045 0.327628
R5540 VGND.n1068 VGND.n1041 0.327628
R5541 VGND.n1071 VGND.n912 0.327628
R5542 VGND.n1076 VGND.n911 0.327628
R5543 VGND.n1081 VGND.n906 0.327628
R5544 VGND.n1086 VGND.n905 0.327628
R5545 VGND.n1091 VGND.n900 0.327628
R5546 VGND.n1096 VGND.n899 0.327628
R5547 VGND.n1100 VGND.n1099 0.327628
R5548 VGND.n1038 VGND.n1026 0.327628
R5549 VGND.n1033 VGND.n1025 0.327628
R5550 VGND.n1167 VGND.n1165 0.327628
R5551 VGND.n1174 VGND.n1170 0.327628
R5552 VGND.n1177 VGND.n1011 0.327628
R5553 VGND.n1187 VGND.n1183 0.327628
R5554 VGND.n1191 VGND.n1190 0.327628
R5555 VGND.n1206 VGND.n1202 0.327628
R5556 VGND.n1209 VGND.n1003 0.327628
R5557 VGND.n1219 VGND.n1215 0.327628
R5558 VGND.n1249 VGND.n1248 0.327628
R5559 VGND.n1245 VGND.n1223 0.327628
R5560 VGND.n1242 VGND.n1241 0.327628
R5561 VGND.n1238 VGND.n1228 0.327628
R5562 VGND.n1235 VGND.n1234 0.327628
R5563 VGND.n1276 VGND.n1272 0.327628
R5564 VGND.n1279 VGND.n997 0.327628
R5565 VGND.n992 VGND.n991 0.327628
R5566 VGND.n988 VGND.n925 0.327628
R5567 VGND.n983 VGND.n924 0.327628
R5568 VGND.n978 VGND.n920 0.327628
R5569 VGND.n973 VGND.n919 0.327628
R5570 VGND.n968 VGND.n915 0.327628
R5571 VGND.n963 VGND.n914 0.327628
R5572 VGND.n958 VGND.n909 0.327628
R5573 VGND.n953 VGND.n908 0.327628
R5574 VGND.n948 VGND.n903 0.327628
R5575 VGND.n943 VGND.n902 0.327628
R5576 VGND.n938 VGND.n897 0.327628
R5577 VGND.n933 VGND.n896 0.327628
R5578 VGND.n1331 VGND.n890 0.327628
R5579 VGND.n1334 VGND.n888 0.327628
R5580 VGND.n126 VGND.n125 0.213567
R5581 VGND.n125 VGND.n32 0.213567
R5582 VGND.n3002 VGND.n32 0.213567
R5583 VGND.n3002 VGND.n3001 0.213567
R5584 VGND.n1157 VGND.n1134 0.213567
R5585 VGND.n1134 VGND.n543 0.213567
R5586 VGND.n2219 VGND.n543 0.213567
R5587 VGND.n2219 VGND.n2218 0.213567
R5588 VGND.n2218 VGND.n0 0.213567
R5589 VGND.n3001 VGND.n33 0.2073
R5590 VGND.n3024 VGND.n2 0.18968
R5591 VGND.n1159 VGND.n1158 0.175967
R5592 VGND.n2633 VGND 0.169807
R5593 VGND.n2695 VGND 0.169807
R5594 VGND.n2690 VGND 0.169807
R5595 VGND.n2689 VGND 0.169807
R5596 VGND.n2684 VGND 0.169807
R5597 VGND.n2683 VGND 0.169807
R5598 VGND.n2678 VGND 0.169807
R5599 VGND.n2677 VGND 0.169807
R5600 VGND.n2709 VGND 0.169807
R5601 VGND.n2723 VGND 0.169807
R5602 VGND.n2742 VGND 0.169807
R5603 VGND.n2761 VGND 0.169807
R5604 VGND.n2781 VGND 0.169807
R5605 VGND.n2780 VGND 0.169807
R5606 VGND.n284 VGND 0.169807
R5607 VGND.n2635 VGND 0.169807
R5608 VGND.n2693 VGND 0.169807
R5609 VGND.n2692 VGND 0.169807
R5610 VGND.n2687 VGND 0.169807
R5611 VGND.n2686 VGND 0.169807
R5612 VGND.n2681 VGND 0.169807
R5613 VGND.n2680 VGND 0.169807
R5614 VGND.n2675 VGND 0.169807
R5615 VGND.n2711 VGND 0.169807
R5616 VGND.n2721 VGND 0.169807
R5617 VGND.n2744 VGND 0.169807
R5618 VGND.n2759 VGND 0.169807
R5619 VGND VGND.n2783 0.169807
R5620 VGND.n2784 VGND 0.169807
R5621 VGND.n2794 VGND 0.169807
R5622 VGND.n2559 VGND 0.169807
R5623 VGND.n2558 VGND 0.169807
R5624 VGND.n2557 VGND 0.169807
R5625 VGND.n2556 VGND 0.169807
R5626 VGND.n2555 VGND 0.169807
R5627 VGND.n2554 VGND 0.169807
R5628 VGND.n2553 VGND 0.169807
R5629 VGND.n2552 VGND 0.169807
R5630 VGND.n2551 VGND 0.169807
R5631 VGND.n2550 VGND 0.169807
R5632 VGND.n2549 VGND 0.169807
R5633 VGND.n2548 VGND 0.169807
R5634 VGND.n2547 VGND 0.169807
R5635 VGND.n2798 VGND 0.169807
R5636 VGND.n2797 VGND 0.169807
R5637 VGND.n2357 VGND 0.169807
R5638 VGND.n2373 VGND 0.169807
R5639 VGND.n2383 VGND 0.169807
R5640 VGND.n2399 VGND 0.169807
R5641 VGND.n2409 VGND 0.169807
R5642 VGND.n2425 VGND 0.169807
R5643 VGND.n2435 VGND 0.169807
R5644 VGND.n2451 VGND 0.169807
R5645 VGND.n2461 VGND 0.169807
R5646 VGND.n2477 VGND 0.169807
R5647 VGND.n2487 VGND 0.169807
R5648 VGND.n2508 VGND 0.169807
R5649 VGND.n2802 VGND 0.169807
R5650 VGND.n2801 VGND 0.169807
R5651 VGND.n419 VGND 0.169807
R5652 VGND.n2360 VGND 0.169807
R5653 VGND.n2370 VGND 0.169807
R5654 VGND.n2386 VGND 0.169807
R5655 VGND.n2396 VGND 0.169807
R5656 VGND.n2412 VGND 0.169807
R5657 VGND.n2422 VGND 0.169807
R5658 VGND.n2438 VGND 0.169807
R5659 VGND.n2448 VGND 0.169807
R5660 VGND.n2464 VGND 0.169807
R5661 VGND.n2474 VGND 0.169807
R5662 VGND.n2490 VGND 0.169807
R5663 VGND.n2505 VGND 0.169807
R5664 VGND VGND.n2805 0.169807
R5665 VGND.n2806 VGND 0.169807
R5666 VGND.n2819 VGND 0.169807
R5667 VGND.n1907 VGND 0.169807
R5668 VGND VGND.n1917 0.169807
R5669 VGND.n1918 VGND 0.169807
R5670 VGND VGND.n1928 0.169807
R5671 VGND.n1929 VGND 0.169807
R5672 VGND VGND.n1939 0.169807
R5673 VGND.n1940 VGND 0.169807
R5674 VGND VGND.n1950 0.169807
R5675 VGND.n1951 VGND 0.169807
R5676 VGND VGND.n1961 0.169807
R5677 VGND.n1962 VGND 0.169807
R5678 VGND VGND.n1972 0.169807
R5679 VGND.n1973 VGND 0.169807
R5680 VGND.n2823 VGND 0.169807
R5681 VGND.n2822 VGND 0.169807
R5682 VGND.n2063 VGND 0.169807
R5683 VGND.n2062 VGND 0.169807
R5684 VGND.n2167 VGND 0.169807
R5685 VGND.n2166 VGND 0.169807
R5686 VGND.n2159 VGND 0.169807
R5687 VGND.n2158 VGND 0.169807
R5688 VGND.n2151 VGND 0.169807
R5689 VGND.n2150 VGND 0.169807
R5690 VGND.n2143 VGND 0.169807
R5691 VGND.n2142 VGND 0.169807
R5692 VGND.n2135 VGND 0.169807
R5693 VGND.n2134 VGND 0.169807
R5694 VGND.n2827 VGND 0.169807
R5695 VGND.n2826 VGND 0.169807
R5696 VGND.n1998 VGND 0.169807
R5697 VGND.n2066 VGND 0.169807
R5698 VGND.n2171 VGND 0.169807
R5699 VGND.n2170 VGND 0.169807
R5700 VGND.n2163 VGND 0.169807
R5701 VGND.n2162 VGND 0.169807
R5702 VGND.n2155 VGND 0.169807
R5703 VGND.n2154 VGND 0.169807
R5704 VGND.n2147 VGND 0.169807
R5705 VGND.n2146 VGND 0.169807
R5706 VGND.n2139 VGND 0.169807
R5707 VGND.n2138 VGND 0.169807
R5708 VGND.n2131 VGND 0.169807
R5709 VGND VGND.n2830 0.169807
R5710 VGND.n2831 VGND 0.169807
R5711 VGND.n2844 VGND 0.169807
R5712 VGND.n1901 VGND 0.169807
R5713 VGND.n2174 VGND 0.169807
R5714 VGND.n1758 VGND 0.169807
R5715 VGND VGND.n1768 0.169807
R5716 VGND.n1769 VGND 0.169807
R5717 VGND VGND.n1779 0.169807
R5718 VGND.n1780 VGND 0.169807
R5719 VGND VGND.n1790 0.169807
R5720 VGND.n1791 VGND 0.169807
R5721 VGND VGND.n1801 0.169807
R5722 VGND.n1802 VGND 0.169807
R5723 VGND VGND.n1812 0.169807
R5724 VGND.n1813 VGND 0.169807
R5725 VGND.n2848 VGND 0.169807
R5726 VGND.n2847 VGND 0.169807
R5727 VGND.n1899 VGND 0.169807
R5728 VGND VGND.n1685 0.169807
R5729 VGND.n1686 VGND 0.169807
R5730 VGND.n1884 VGND 0.169807
R5731 VGND.n1883 VGND 0.169807
R5732 VGND.n1876 VGND 0.169807
R5733 VGND.n1875 VGND 0.169807
R5734 VGND.n1868 VGND 0.169807
R5735 VGND.n1867 VGND 0.169807
R5736 VGND.n1860 VGND 0.169807
R5737 VGND.n1859 VGND 0.169807
R5738 VGND.n1852 VGND 0.169807
R5739 VGND.n2852 VGND 0.169807
R5740 VGND.n2851 VGND 0.169807
R5741 VGND.n1838 VGND 0.169807
R5742 VGND.n1896 VGND 0.169807
R5743 VGND.n1895 VGND 0.169807
R5744 VGND.n1888 VGND 0.169807
R5745 VGND.n1887 VGND 0.169807
R5746 VGND.n1880 VGND 0.169807
R5747 VGND.n1879 VGND 0.169807
R5748 VGND.n1872 VGND 0.169807
R5749 VGND.n1871 VGND 0.169807
R5750 VGND.n1864 VGND 0.169807
R5751 VGND.n1863 VGND 0.169807
R5752 VGND.n1856 VGND 0.169807
R5753 VGND.n1855 VGND 0.169807
R5754 VGND VGND.n2855 0.169807
R5755 VGND.n2856 VGND 0.169807
R5756 VGND.n2869 VGND 0.169807
R5757 VGND.n1349 VGND 0.169807
R5758 VGND.n1892 VGND 0.169807
R5759 VGND.n1891 VGND 0.169807
R5760 VGND.n867 VGND 0.169807
R5761 VGND.n866 VGND 0.169807
R5762 VGND.n865 VGND 0.169807
R5763 VGND.n864 VGND 0.169807
R5764 VGND.n863 VGND 0.169807
R5765 VGND.n862 VGND 0.169807
R5766 VGND.n861 VGND 0.169807
R5767 VGND.n860 VGND 0.169807
R5768 VGND.n1669 VGND 0.169807
R5769 VGND.n1668 VGND 0.169807
R5770 VGND.n2873 VGND 0.169807
R5771 VGND.n2872 VGND 0.169807
R5772 VGND.n1404 VGND 0.169807
R5773 VGND.n1403 VGND 0.169807
R5774 VGND.n1402 VGND 0.169807
R5775 VGND.n1487 VGND 0.169807
R5776 VGND.n1497 VGND 0.169807
R5777 VGND.n1513 VGND 0.169807
R5778 VGND.n1523 VGND 0.169807
R5779 VGND.n1539 VGND 0.169807
R5780 VGND.n1560 VGND 0.169807
R5781 VGND.n1559 VGND 0.169807
R5782 VGND VGND.n1628 0.169807
R5783 VGND.n1629 VGND 0.169807
R5784 VGND.n2877 VGND 0.169807
R5785 VGND.n2876 VGND 0.169807
R5786 VGND.n740 VGND 0.169807
R5787 VGND.n1407 VGND 0.169807
R5788 VGND.n1417 VGND 0.169807
R5789 VGND.n1474 VGND 0.169807
R5790 VGND.n1484 VGND 0.169807
R5791 VGND.n1500 VGND 0.169807
R5792 VGND.n1510 VGND 0.169807
R5793 VGND.n1526 VGND 0.169807
R5794 VGND.n1536 VGND 0.169807
R5795 VGND.n1563 VGND 0.169807
R5796 VGND.n1588 VGND 0.169807
R5797 VGND.n1625 VGND 0.169807
R5798 VGND.n1624 VGND 0.169807
R5799 VGND VGND.n2880 0.169807
R5800 VGND.n2881 VGND 0.169807
R5801 VGND.n2894 VGND 0.169807
R5802 VGND.n1344 VGND 0.169807
R5803 VGND.n1420 VGND 0.169807
R5804 VGND.n1471 VGND 0.169807
R5805 VGND.n1470 VGND 0.169807
R5806 VGND.n1469 VGND 0.169807
R5807 VGND.n1468 VGND 0.169807
R5808 VGND.n1467 VGND 0.169807
R5809 VGND.n1466 VGND 0.169807
R5810 VGND.n1465 VGND 0.169807
R5811 VGND VGND.n1591 0.169807
R5812 VGND.n1592 VGND 0.169807
R5813 VGND.n1621 VGND 0.169807
R5814 VGND.n1620 VGND 0.169807
R5815 VGND.n2898 VGND 0.169807
R5816 VGND.n2897 VGND 0.169807
R5817 VGND.n1103 VGND 0.169807
R5818 VGND.n1102 VGND 0.169807
R5819 VGND.n1101 VGND 0.169807
R5820 VGND.n1321 VGND 0.169807
R5821 VGND.n1320 VGND 0.169807
R5822 VGND.n1313 VGND 0.169807
R5823 VGND.n1312 VGND 0.169807
R5824 VGND.n1305 VGND 0.169807
R5825 VGND.n1304 VGND 0.169807
R5826 VGND.n1067 VGND 0.169807
R5827 VGND.n1066 VGND 0.169807
R5828 VGND.n1065 VGND 0.169807
R5829 VGND.n1064 VGND 0.169807
R5830 VGND.n2901 VGND 0.169807
R5831 VGND.n233 VGND 0.169807
R5832 VGND.n1163 VGND 0.169807
R5833 VGND.n1328 VGND 0.169807
R5834 VGND.n1327 VGND 0.169807
R5835 VGND VGND.n898 0.169807
R5836 VGND VGND.n901 0.169807
R5837 VGND VGND.n904 0.169807
R5838 VGND VGND.n907 0.169807
R5839 VGND VGND.n910 0.169807
R5840 VGND VGND.n913 0.169807
R5841 VGND.n1298 VGND 0.169807
R5842 VGND.n1297 VGND 0.169807
R5843 VGND.n1292 VGND 0.169807
R5844 VGND.n1291 VGND 0.169807
R5845 VGND.n1270 VGND 0.169807
R5846 VGND.n1285 VGND 0.169807
R5847 VGND.n1161 VGND 0.169807
R5848 VGND.n1330 VGND 0.169807
R5849 VGND.n1325 VGND 0.169807
R5850 VGND.n1324 VGND 0.169807
R5851 VGND.n1317 VGND 0.169807
R5852 VGND.n1316 VGND 0.169807
R5853 VGND.n1309 VGND 0.169807
R5854 VGND.n1308 VGND 0.169807
R5855 VGND.n1301 VGND 0.169807
R5856 VGND.n1300 VGND 0.169807
R5857 VGND.n1295 VGND 0.169807
R5858 VGND.n1294 VGND 0.169807
R5859 VGND.n1289 VGND 0.169807
R5860 VGND.n1288 VGND 0.169807
R5861 VGND.n1287 VGND 0.169807
R5862 VGND.n190 VGND 0.159538
R5863 VGND.n161 VGND 0.159538
R5864 VGND.n2915 VGND.n224 0.154425
R5865 VGND.n2915 VGND.n2914 0.154425
R5866 VGND.n2914 VGND.n225 0.154425
R5867 VGND.n238 VGND.n225 0.154425
R5868 VGND.n1652 VGND.n238 0.154425
R5869 VGND.n1653 VGND.n1652 0.154425
R5870 VGND.n1653 VGND.n251 0.154425
R5871 VGND.n1832 VGND.n251 0.154425
R5872 VGND.n1832 VGND.n1831 0.154425
R5873 VGND.n1831 VGND.n263 0.154425
R5874 VGND.n1992 VGND.n263 0.154425
R5875 VGND.n1992 VGND.n1991 0.154425
R5876 VGND.n1991 VGND.n275 0.154425
R5877 VGND.n417 VGND.n275 0.154425
R5878 VGND.n417 VGND.n207 0.154425
R5879 VGND.n2938 VGND.n207 0.154425
R5880 VGND.n2939 VGND.n2938 0.154425
R5881 VGND.n1160 VGND.n1159 0.154425
R5882 VGND.n1160 VGND.n880 0.154425
R5883 VGND.n1345 VGND.n880 0.154425
R5884 VGND.n1346 VGND.n1345 0.154425
R5885 VGND.n1347 VGND.n1346 0.154425
R5886 VGND.n1348 VGND.n1347 0.154425
R5887 VGND.n1348 VGND.n626 0.154425
R5888 VGND.n1900 VGND.n626 0.154425
R5889 VGND.n1902 VGND.n1900 0.154425
R5890 VGND.n1903 VGND.n1902 0.154425
R5891 VGND.n1904 VGND.n1903 0.154425
R5892 VGND.n1906 VGND.n1904 0.154425
R5893 VGND.n1906 VGND.n1905 0.154425
R5894 VGND.n1905 VGND.n398 0.154425
R5895 VGND.n2560 VGND.n398 0.154425
R5896 VGND.n2561 VGND.n2560 0.154425
R5897 VGND.n2562 VGND.n2561 0.154425
R5898 VGND.n1144 VGND.n1138 0.144904
R5899 VGND.n1117 VGND.n1109 0.144904
R5900 VGND.n2232 VGND.n2228 0.144904
R5901 VGND.n1370 VGND.n1366 0.144904
R5902 VGND.n2632 VGND.n2608 0.138284
R5903 VGND.n2700 VGND.n2699 0.13638
R5904 VGND.n355 VGND.n333 0.13638
R5905 VGND.n362 VGND.n361 0.13638
R5906 VGND.n369 VGND.n368 0.13638
R5907 VGND.n373 VGND.n372 0.13638
R5908 VGND.n380 VGND.n379 0.13638
R5909 VGND.n384 VGND.n383 0.13638
R5910 VGND.n388 VGND.n387 0.13638
R5911 VGND.n2706 VGND.n326 0.13638
R5912 VGND.n2727 VGND.n2726 0.13638
R5913 VGND.n2739 VGND.n312 0.13638
R5914 VGND.n2736 VGND.n2735 0.13638
R5915 VGND.n2732 VGND.n2730 0.13638
R5916 VGND.n2777 VGND.n294 0.13638
R5917 VGND.n2774 VGND.n2773 0.13638
R5918 VGND.n2792 VGND.n287 0.13638
R5919 VGND.n2789 VGND.n2788 0.13638
R5920 VGND.n2754 VGND.n2753 0.13638
R5921 VGND.n2757 VGND.n304 0.13638
R5922 VGND.n2749 VGND.n2748 0.13638
R5923 VGND.n2719 VGND.n320 0.13638
R5924 VGND.n2716 VGND.n2715 0.13638
R5925 VGND.n2673 VGND.n394 0.13638
R5926 VGND.n2670 VGND.n2669 0.13638
R5927 VGND.n2665 VGND.n2664 0.13638
R5928 VGND.n2660 VGND.n2659 0.13638
R5929 VGND.n2655 VGND.n2654 0.13638
R5930 VGND.n2650 VGND.n2649 0.13638
R5931 VGND.n2645 VGND.n2644 0.13638
R5932 VGND.n2640 VGND.n2639 0.13638
R5933 VGND.n2537 VGND.n2536 0.13638
R5934 VGND.n2542 VGND.n2541 0.13638
R5935 VGND.n2545 VGND.n415 0.13638
R5936 VGND.n2289 VGND.n2288 0.13638
R5937 VGND.n2294 VGND.n2293 0.13638
R5938 VGND.n2299 VGND.n2298 0.13638
R5939 VGND.n2304 VGND.n2303 0.13638
R5940 VGND.n2309 VGND.n2308 0.13638
R5941 VGND.n2314 VGND.n2313 0.13638
R5942 VGND.n2319 VGND.n2318 0.13638
R5943 VGND.n2324 VGND.n2323 0.13638
R5944 VGND.n2329 VGND.n2328 0.13638
R5945 VGND.n2334 VGND.n2333 0.13638
R5946 VGND.n2339 VGND.n2338 0.13638
R5947 VGND.n2344 VGND.n2343 0.13638
R5948 VGND.n2527 VGND.n2526 0.13638
R5949 VGND.n2523 VGND.n2522 0.13638
R5950 VGND.n2518 VGND.n2517 0.13638
R5951 VGND.n2513 VGND.n2512 0.13638
R5952 VGND.n2485 VGND.n428 0.13638
R5953 VGND.n2482 VGND.n2481 0.13638
R5954 VGND.n2459 VGND.n436 0.13638
R5955 VGND.n2456 VGND.n2455 0.13638
R5956 VGND.n2433 VGND.n444 0.13638
R5957 VGND.n2430 VGND.n2429 0.13638
R5958 VGND.n2407 VGND.n452 0.13638
R5959 VGND.n2404 VGND.n2403 0.13638
R5960 VGND.n2381 VGND.n460 0.13638
R5961 VGND.n2378 VGND.n2377 0.13638
R5962 VGND.n2355 VGND.n472 0.13638
R5963 VGND.n2815 VGND.n2814 0.13638
R5964 VGND.n2811 VGND.n2810 0.13638
R5965 VGND.n2500 VGND.n2499 0.13638
R5966 VGND.n2503 VGND.n424 0.13638
R5967 VGND.n2495 VGND.n2494 0.13638
R5968 VGND.n2472 VGND.n432 0.13638
R5969 VGND.n2469 VGND.n2468 0.13638
R5970 VGND.n2446 VGND.n440 0.13638
R5971 VGND.n2443 VGND.n2442 0.13638
R5972 VGND.n2420 VGND.n448 0.13638
R5973 VGND.n2417 VGND.n2416 0.13638
R5974 VGND.n2394 VGND.n456 0.13638
R5975 VGND.n2391 VGND.n2390 0.13638
R5976 VGND.n2368 VGND.n464 0.13638
R5977 VGND.n2365 VGND.n2364 0.13638
R5978 VGND.n1987 VGND.n1986 0.13638
R5979 VGND.n1983 VGND.n1982 0.13638
R5980 VGND.n1978 VGND.n1977 0.13638
R5981 VGND.n1970 VGND.n608 0.13638
R5982 VGND.n1967 VGND.n1966 0.13638
R5983 VGND.n1959 VGND.n611 0.13638
R5984 VGND.n1956 VGND.n1955 0.13638
R5985 VGND.n1948 VGND.n614 0.13638
R5986 VGND.n1945 VGND.n1944 0.13638
R5987 VGND.n1937 VGND.n617 0.13638
R5988 VGND.n1934 VGND.n1933 0.13638
R5989 VGND.n1926 VGND.n620 0.13638
R5990 VGND.n1923 VGND.n1922 0.13638
R5991 VGND.n1915 VGND.n623 0.13638
R5992 VGND.n1912 VGND.n1911 0.13638
R5993 VGND.n1994 VGND.n602 0.13638
R5994 VGND.n2002 VGND.n2001 0.13638
R5995 VGND.n2007 VGND.n2006 0.13638
R5996 VGND.n2012 VGND.n2011 0.13638
R5997 VGND.n2017 VGND.n2016 0.13638
R5998 VGND.n2022 VGND.n2021 0.13638
R5999 VGND.n2027 VGND.n2026 0.13638
R6000 VGND.n2032 VGND.n2031 0.13638
R6001 VGND.n2037 VGND.n2036 0.13638
R6002 VGND.n2042 VGND.n2041 0.13638
R6003 VGND.n2047 VGND.n2046 0.13638
R6004 VGND.n2052 VGND.n2051 0.13638
R6005 VGND.n2057 VGND.n2056 0.13638
R6006 VGND.n2060 VGND.n594 0.13638
R6007 VGND.n598 VGND.n597 0.13638
R6008 VGND.n2840 VGND.n2839 0.13638
R6009 VGND.n2836 VGND.n2835 0.13638
R6010 VGND.n2126 VGND.n2125 0.13638
R6011 VGND.n2129 VGND.n585 0.13638
R6012 VGND.n2121 VGND.n2120 0.13638
R6013 VGND.n2116 VGND.n2115 0.13638
R6014 VGND.n2111 VGND.n2110 0.13638
R6015 VGND.n2106 VGND.n2105 0.13638
R6016 VGND.n2101 VGND.n2100 0.13638
R6017 VGND.n2096 VGND.n2095 0.13638
R6018 VGND.n2091 VGND.n2090 0.13638
R6019 VGND.n2086 VGND.n2085 0.13638
R6020 VGND.n2081 VGND.n2080 0.13638
R6021 VGND.n2076 VGND.n2075 0.13638
R6022 VGND.n2071 VGND.n2070 0.13638
R6023 VGND.n1827 VGND.n1826 0.13638
R6024 VGND.n1823 VGND.n1822 0.13638
R6025 VGND.n1818 VGND.n1817 0.13638
R6026 VGND.n1810 VGND.n1741 0.13638
R6027 VGND.n1807 VGND.n1806 0.13638
R6028 VGND.n1799 VGND.n1744 0.13638
R6029 VGND.n1796 VGND.n1795 0.13638
R6030 VGND.n1788 VGND.n1747 0.13638
R6031 VGND.n1785 VGND.n1784 0.13638
R6032 VGND.n1777 VGND.n1750 0.13638
R6033 VGND.n1774 VGND.n1773 0.13638
R6034 VGND.n1766 VGND.n1753 0.13638
R6035 VGND.n1763 VGND.n1762 0.13638
R6036 VGND.n1756 VGND.n550 0.13638
R6037 VGND.n2178 VGND.n2177 0.13638
R6038 VGND.n1834 VGND.n1735 0.13638
R6039 VGND.n1842 VGND.n1841 0.13638
R6040 VGND.n1847 VGND.n1846 0.13638
R6041 VGND.n1850 VGND.n1673 0.13638
R6042 VGND.n1731 VGND.n1730 0.13638
R6043 VGND.n1726 VGND.n1725 0.13638
R6044 VGND.n1721 VGND.n1720 0.13638
R6045 VGND.n1716 VGND.n1715 0.13638
R6046 VGND.n1711 VGND.n1710 0.13638
R6047 VGND.n1706 VGND.n1705 0.13638
R6048 VGND.n1701 VGND.n1700 0.13638
R6049 VGND.n1696 VGND.n1695 0.13638
R6050 VGND.n1691 VGND.n1690 0.13638
R6051 VGND.n1683 VGND.n1676 0.13638
R6052 VGND.n1680 VGND.n1679 0.13638
R6053 VGND.n2865 VGND.n2864 0.13638
R6054 VGND.n2861 VGND.n2860 0.13638
R6055 VGND.n726 VGND.n725 0.13638
R6056 VGND.n729 VGND.n667 0.13638
R6057 VGND.n721 VGND.n720 0.13638
R6058 VGND.n716 VGND.n715 0.13638
R6059 VGND.n711 VGND.n710 0.13638
R6060 VGND.n706 VGND.n705 0.13638
R6061 VGND.n701 VGND.n700 0.13638
R6062 VGND.n696 VGND.n695 0.13638
R6063 VGND.n691 VGND.n690 0.13638
R6064 VGND.n686 VGND.n685 0.13638
R6065 VGND.n681 VGND.n680 0.13638
R6066 VGND.n676 VGND.n675 0.13638
R6067 VGND.n671 VGND.n670 0.13638
R6068 VGND.n1658 VGND.n1657 0.13638
R6069 VGND.n1663 VGND.n1662 0.13638
R6070 VGND.n1666 VGND.n735 0.13638
R6071 VGND.n855 VGND.n854 0.13638
R6072 VGND.n858 VGND.n820 0.13638
R6073 VGND.n850 VGND.n849 0.13638
R6074 VGND.n845 VGND.n844 0.13638
R6075 VGND.n840 VGND.n839 0.13638
R6076 VGND.n835 VGND.n834 0.13638
R6077 VGND.n830 VGND.n829 0.13638
R6078 VGND.n825 VGND.n824 0.13638
R6079 VGND.n810 VGND.n808 0.13638
R6080 VGND.n871 VGND.n870 0.13638
R6081 VGND.n876 VGND.n875 0.13638
R6082 VGND.n1354 VGND.n1353 0.13638
R6083 VGND.n1648 VGND.n1647 0.13638
R6084 VGND.n1644 VGND.n1643 0.13638
R6085 VGND.n1639 VGND.n1638 0.13638
R6086 VGND.n1634 VGND.n1633 0.13638
R6087 VGND.n1554 VGND.n1553 0.13638
R6088 VGND.n1557 VGND.n761 0.13638
R6089 VGND.n1549 VGND.n1548 0.13638
R6090 VGND.n1544 VGND.n1543 0.13638
R6091 VGND.n1521 VGND.n769 0.13638
R6092 VGND.n1518 VGND.n1517 0.13638
R6093 VGND.n1495 VGND.n777 0.13638
R6094 VGND.n1492 VGND.n1491 0.13638
R6095 VGND.n1400 VGND.n805 0.13638
R6096 VGND.n1397 VGND.n1396 0.13638
R6097 VGND.n1392 VGND.n1391 0.13638
R6098 VGND.n2890 VGND.n2889 0.13638
R6099 VGND.n2886 VGND.n2885 0.13638
R6100 VGND.n1573 VGND.n1572 0.13638
R6101 VGND.n1578 VGND.n1577 0.13638
R6102 VGND.n1583 VGND.n1582 0.13638
R6103 VGND.n1586 VGND.n756 0.13638
R6104 VGND.n1568 VGND.n1567 0.13638
R6105 VGND.n1534 VGND.n765 0.13638
R6106 VGND.n1531 VGND.n1530 0.13638
R6107 VGND.n1508 VGND.n773 0.13638
R6108 VGND.n1505 VGND.n1504 0.13638
R6109 VGND.n1482 VGND.n781 0.13638
R6110 VGND.n1479 VGND.n1478 0.13638
R6111 VGND.n1415 VGND.n795 0.13638
R6112 VGND.n1412 VGND.n1411 0.13638
R6113 VGND.n1610 VGND.n1609 0.13638
R6114 VGND.n1615 VGND.n1614 0.13638
R6115 VGND.n1618 VGND.n750 0.13638
R6116 VGND.n1602 VGND.n1601 0.13638
R6117 VGND.n1597 VGND.n1596 0.13638
R6118 VGND.n1460 VGND.n1459 0.13638
R6119 VGND.n1463 VGND.n791 0.13638
R6120 VGND.n1455 VGND.n1454 0.13638
R6121 VGND.n1450 VGND.n1449 0.13638
R6122 VGND.n1445 VGND.n1444 0.13638
R6123 VGND.n1440 VGND.n1439 0.13638
R6124 VGND.n1435 VGND.n1434 0.13638
R6125 VGND.n1430 VGND.n1429 0.13638
R6126 VGND.n1425 VGND.n1424 0.13638
R6127 VGND.n1342 VGND.n885 0.13638
R6128 VGND.n2910 VGND.n2909 0.13638
R6129 VGND.n2906 VGND.n2905 0.13638
R6130 VGND.n1062 VGND.n1049 0.13638
R6131 VGND.n1059 VGND.n1058 0.13638
R6132 VGND.n1054 VGND.n1053 0.13638
R6133 VGND.n1043 VGND.n1041 0.13638
R6134 VGND.n1071 VGND.n1070 0.13638
R6135 VGND.n1076 VGND.n1075 0.13638
R6136 VGND.n1081 VGND.n1080 0.13638
R6137 VGND.n1086 VGND.n1085 0.13638
R6138 VGND.n1091 VGND.n1090 0.13638
R6139 VGND.n1096 VGND.n1095 0.13638
R6140 VGND.n1099 VGND.n1029 0.13638
R6141 VGND.n1038 VGND.n1037 0.13638
R6142 VGND.n1033 VGND.n1032 0.13638
R6143 VGND.n1168 VGND.n1167 0.13638
R6144 VGND.n1174 VGND.n1173 0.13638
R6145 VGND.n1178 VGND.n1177 0.13638
R6146 VGND.n1187 VGND.n1186 0.13638
R6147 VGND.n1190 VGND.n1009 0.13638
R6148 VGND.n1206 VGND.n1205 0.13638
R6149 VGND.n1210 VGND.n1209 0.13638
R6150 VGND.n1219 VGND.n1218 0.13638
R6151 VGND.n1248 VGND.n1001 0.13638
R6152 VGND.n1245 VGND.n1244 0.13638
R6153 VGND.n1241 VGND.n1225 0.13638
R6154 VGND.n1238 VGND.n1237 0.13638
R6155 VGND.n1234 VGND.n1232 0.13638
R6156 VGND.n1276 VGND.n1275 0.13638
R6157 VGND.n1280 VGND.n1279 0.13638
R6158 VGND.n991 VGND.n928 0.13638
R6159 VGND.n988 VGND.n987 0.13638
R6160 VGND.n983 VGND.n982 0.13638
R6161 VGND.n978 VGND.n977 0.13638
R6162 VGND.n973 VGND.n972 0.13638
R6163 VGND.n968 VGND.n967 0.13638
R6164 VGND.n963 VGND.n962 0.13638
R6165 VGND.n958 VGND.n957 0.13638
R6166 VGND.n953 VGND.n952 0.13638
R6167 VGND.n948 VGND.n947 0.13638
R6168 VGND.n943 VGND.n942 0.13638
R6169 VGND.n938 VGND.n937 0.13638
R6170 VGND.n933 VGND.n932 0.13638
R6171 VGND.n894 VGND.n890 0.13638
R6172 VGND.n1334 VGND.n1333 0.13638
R6173 VGND VGND.n190 0.120838
R6174 VGND.n19 VGND.n13 0.120292
R6175 VGND.n24 VGND.n13 0.120292
R6176 VGND.n25 VGND.n24 0.120292
R6177 VGND.n26 VGND.n25 0.120292
R6178 VGND.n26 VGND.n11 0.120292
R6179 VGND.n30 VGND.n11 0.120292
R6180 VGND.n31 VGND.n30 0.120292
R6181 VGND.n3008 VGND.n3007 0.120292
R6182 VGND.n3007 VGND.n3003 0.120292
R6183 VGND.n182 VGND.n174 0.120292
R6184 VGND.n183 VGND.n182 0.120292
R6185 VGND.n183 VGND.n168 0.120292
R6186 VGND.n188 VGND.n168 0.120292
R6187 VGND.n189 VGND.n188 0.120292
R6188 VGND.n2952 VGND.n2948 0.120292
R6189 VGND.n2957 VGND.n2948 0.120292
R6190 VGND.n2958 VGND.n2957 0.120292
R6191 VGND.n2959 VGND.n2958 0.120292
R6192 VGND.n2959 VGND.n2946 0.120292
R6193 VGND.n2963 VGND.n2946 0.120292
R6194 VGND.n2964 VGND.n2963 0.120292
R6195 VGND.n45 VGND.n39 0.120292
R6196 VGND.n50 VGND.n39 0.120292
R6197 VGND.n51 VGND.n50 0.120292
R6198 VGND.n52 VGND.n51 0.120292
R6199 VGND.n52 VGND.n37 0.120292
R6200 VGND.n56 VGND.n37 0.120292
R6201 VGND.n57 VGND.n56 0.120292
R6202 VGND.n63 VGND.n62 0.120292
R6203 VGND.n62 VGND.n58 0.120292
R6204 VGND.n106 VGND.n99 0.120292
R6205 VGND.n107 VGND.n106 0.120292
R6206 VGND.n107 VGND.n94 0.120292
R6207 VGND.n112 VGND.n94 0.120292
R6208 VGND.n113 VGND.n112 0.120292
R6209 VGND.n124 VGND.n91 0.120292
R6210 VGND.n83 VGND.n75 0.120292
R6211 VGND.n84 VGND.n83 0.120292
R6212 VGND.n84 VGND.n69 0.120292
R6213 VGND.n89 VGND.n69 0.120292
R6214 VGND.n90 VGND.n89 0.120292
R6215 VGND.n130 VGND.n127 0.120292
R6216 VGND.n151 VGND.n143 0.120292
R6217 VGND.n152 VGND.n151 0.120292
R6218 VGND.n152 VGND.n137 0.120292
R6219 VGND.n157 VGND.n137 0.120292
R6220 VGND.n158 VGND.n157 0.120292
R6221 VGND.n1152 VGND.n1151 0.120292
R6222 VGND.n1151 VGND.n1150 0.120292
R6223 VGND.n1150 VGND.n1136 0.120292
R6224 VGND.n1146 VGND.n1136 0.120292
R6225 VGND.n1146 VGND.n1145 0.120292
R6226 VGND.n1145 VGND.n1144 0.120292
R6227 VGND.n1130 VGND.n1129 0.120292
R6228 VGND.n1125 VGND.n1124 0.120292
R6229 VGND.n1124 VGND.n1123 0.120292
R6230 VGND.n1123 VGND.n1107 0.120292
R6231 VGND.n1119 VGND.n1107 0.120292
R6232 VGND.n1119 VGND.n1118 0.120292
R6233 VGND.n1118 VGND.n1117 0.120292
R6234 VGND.n499 VGND.n476 0.120292
R6235 VGND.n493 VGND.n476 0.120292
R6236 VGND.n493 VGND.n492 0.120292
R6237 VGND.n492 VGND.n480 0.120292
R6238 VGND.n485 VGND.n480 0.120292
R6239 VGND.n485 VGND.n484 0.120292
R6240 VGND.n484 VGND.n483 0.120292
R6241 VGND.n2280 VGND.n2257 0.120292
R6242 VGND.n2274 VGND.n2257 0.120292
R6243 VGND.n2274 VGND.n2273 0.120292
R6244 VGND.n2273 VGND.n2261 0.120292
R6245 VGND.n2266 VGND.n2261 0.120292
R6246 VGND.n2266 VGND.n2265 0.120292
R6247 VGND.n2265 VGND.n2264 0.120292
R6248 VGND.n510 VGND.n507 0.120292
R6249 VGND.n511 VGND.n510 0.120292
R6250 VGND.n535 VGND.n512 0.120292
R6251 VGND.n529 VGND.n512 0.120292
R6252 VGND.n529 VGND.n528 0.120292
R6253 VGND.n528 VGND.n516 0.120292
R6254 VGND.n521 VGND.n516 0.120292
R6255 VGND.n521 VGND.n520 0.120292
R6256 VGND.n520 VGND.n519 0.120292
R6257 VGND.n2214 VGND.n2213 0.120292
R6258 VGND.n2207 VGND.n2183 0.120292
R6259 VGND.n2202 VGND.n2183 0.120292
R6260 VGND.n2202 VGND.n2201 0.120292
R6261 VGND.n2198 VGND.n2197 0.120292
R6262 VGND.n2197 VGND.n2192 0.120292
R6263 VGND.n2193 VGND.n2192 0.120292
R6264 VGND.n2225 VGND.n2224 0.120292
R6265 VGND.n2245 VGND.n2244 0.120292
R6266 VGND.n2244 VGND.n2226 0.120292
R6267 VGND.n2240 VGND.n2226 0.120292
R6268 VGND.n2240 VGND.n2239 0.120292
R6269 VGND.n2239 VGND.n2238 0.120292
R6270 VGND.n2238 VGND.n2228 0.120292
R6271 VGND.n1363 VGND.n1362 0.120292
R6272 VGND.n1383 VGND.n1382 0.120292
R6273 VGND.n1382 VGND.n1364 0.120292
R6274 VGND.n1378 VGND.n1364 0.120292
R6275 VGND.n1378 VGND.n1377 0.120292
R6276 VGND.n1377 VGND.n1376 0.120292
R6277 VGND.n1376 VGND.n1366 0.120292
R6278 VGND.n2983 VGND.n2982 0.120292
R6279 VGND.n2983 VGND.n2975 0.120292
R6280 VGND.n2988 VGND.n2975 0.120292
R6281 VGND.n2989 VGND.n2988 0.120292
R6282 VGND.n2990 VGND.n2989 0.120292
R6283 VGND.n2990 VGND.n2973 0.120292
R6284 VGND.n2994 VGND.n2973 0.120292
R6285 VGND.n2996 VGND.n34 0.120292
R6286 VGND.n3000 VGND.n34 0.120292
R6287 VGND VGND.n161 0.119536
R6288 VGND.n1138 VGND 0.117202
R6289 VGND.n1109 VGND 0.117202
R6290 VGND.n2232 VGND 0.117202
R6291 VGND.n1370 VGND 0.117202
R6292 VGND.n287 VGND.n286 0.110872
R6293 VGND.n2788 VGND.n2787 0.110872
R6294 VGND.n2753 VGND.n2752 0.110872
R6295 VGND.n304 VGND.n303 0.110872
R6296 VGND.n2748 VGND.n2747 0.110872
R6297 VGND.n320 VGND.n319 0.110872
R6298 VGND.n2715 VGND.n2714 0.110872
R6299 VGND.n394 VGND.n393 0.110872
R6300 VGND.n2669 VGND.n2668 0.110872
R6301 VGND.n2664 VGND.n2663 0.110872
R6302 VGND.n2659 VGND.n2658 0.110872
R6303 VGND.n2654 VGND.n2653 0.110872
R6304 VGND.n2649 VGND.n2648 0.110872
R6305 VGND.n2644 VGND.n2643 0.110872
R6306 VGND.n2639 VGND.n2638 0.110872
R6307 VGND.n2536 VGND.n2535 0.110872
R6308 VGND.n2541 VGND.n2540 0.110872
R6309 VGND.n415 VGND.n414 0.110872
R6310 VGND.n2288 VGND.n2287 0.110872
R6311 VGND.n2293 VGND.n2292 0.110872
R6312 VGND.n2298 VGND.n2297 0.110872
R6313 VGND.n2303 VGND.n2302 0.110872
R6314 VGND.n2308 VGND.n2307 0.110872
R6315 VGND.n2313 VGND.n2312 0.110872
R6316 VGND.n2318 VGND.n2317 0.110872
R6317 VGND.n2323 VGND.n2322 0.110872
R6318 VGND.n2328 VGND.n2327 0.110872
R6319 VGND.n2333 VGND.n2332 0.110872
R6320 VGND.n2338 VGND.n2337 0.110872
R6321 VGND.n2343 VGND.n2342 0.110872
R6322 VGND.n2528 VGND.n2527 0.110872
R6323 VGND.n2522 VGND.n2521 0.110872
R6324 VGND.n2517 VGND.n2516 0.110872
R6325 VGND.n2512 VGND.n2511 0.110872
R6326 VGND.n428 VGND.n427 0.110872
R6327 VGND.n2481 VGND.n2480 0.110872
R6328 VGND.n436 VGND.n435 0.110872
R6329 VGND.n2455 VGND.n2454 0.110872
R6330 VGND.n444 VGND.n443 0.110872
R6331 VGND.n2429 VGND.n2428 0.110872
R6332 VGND.n452 VGND.n451 0.110872
R6333 VGND.n2403 VGND.n2402 0.110872
R6334 VGND.n460 VGND.n459 0.110872
R6335 VGND.n2377 VGND.n2376 0.110872
R6336 VGND.n472 VGND.n471 0.110872
R6337 VGND.n2816 VGND.n2815 0.110872
R6338 VGND.n2810 VGND.n2809 0.110872
R6339 VGND.n2499 VGND.n2498 0.110872
R6340 VGND.n424 VGND.n423 0.110872
R6341 VGND.n2494 VGND.n2493 0.110872
R6342 VGND.n432 VGND.n431 0.110872
R6343 VGND.n2468 VGND.n2467 0.110872
R6344 VGND.n440 VGND.n439 0.110872
R6345 VGND.n2442 VGND.n2441 0.110872
R6346 VGND.n448 VGND.n447 0.110872
R6347 VGND.n2416 VGND.n2415 0.110872
R6348 VGND.n456 VGND.n455 0.110872
R6349 VGND.n2390 VGND.n2389 0.110872
R6350 VGND.n464 VGND.n463 0.110872
R6351 VGND.n2364 VGND.n2363 0.110872
R6352 VGND.n1988 VGND.n1987 0.110872
R6353 VGND.n1982 VGND.n1981 0.110872
R6354 VGND.n1977 VGND.n1976 0.110872
R6355 VGND.n608 VGND.n607 0.110872
R6356 VGND.n1966 VGND.n1965 0.110872
R6357 VGND.n611 VGND.n610 0.110872
R6358 VGND.n1955 VGND.n1954 0.110872
R6359 VGND.n614 VGND.n613 0.110872
R6360 VGND.n1944 VGND.n1943 0.110872
R6361 VGND.n617 VGND.n616 0.110872
R6362 VGND.n1933 VGND.n1932 0.110872
R6363 VGND.n620 VGND.n619 0.110872
R6364 VGND.n1922 VGND.n1921 0.110872
R6365 VGND.n623 VGND.n622 0.110872
R6366 VGND.n1911 VGND.n1910 0.110872
R6367 VGND.n1995 VGND.n1994 0.110872
R6368 VGND.n2001 VGND.n2000 0.110872
R6369 VGND.n2006 VGND.n2005 0.110872
R6370 VGND.n2011 VGND.n2010 0.110872
R6371 VGND.n2016 VGND.n2015 0.110872
R6372 VGND.n2021 VGND.n2020 0.110872
R6373 VGND.n2026 VGND.n2025 0.110872
R6374 VGND.n2031 VGND.n2030 0.110872
R6375 VGND.n2036 VGND.n2035 0.110872
R6376 VGND.n2041 VGND.n2040 0.110872
R6377 VGND.n2046 VGND.n2045 0.110872
R6378 VGND.n2051 VGND.n2050 0.110872
R6379 VGND.n2056 VGND.n2055 0.110872
R6380 VGND.n594 VGND.n593 0.110872
R6381 VGND.n597 VGND.n596 0.110872
R6382 VGND.n2841 VGND.n2840 0.110872
R6383 VGND.n2835 VGND.n2834 0.110872
R6384 VGND.n2125 VGND.n2124 0.110872
R6385 VGND.n585 VGND.n584 0.110872
R6386 VGND.n2120 VGND.n2119 0.110872
R6387 VGND.n2115 VGND.n2114 0.110872
R6388 VGND.n2110 VGND.n2109 0.110872
R6389 VGND.n2105 VGND.n2104 0.110872
R6390 VGND.n2100 VGND.n2099 0.110872
R6391 VGND.n2095 VGND.n2094 0.110872
R6392 VGND.n2090 VGND.n2089 0.110872
R6393 VGND.n2085 VGND.n2084 0.110872
R6394 VGND.n2080 VGND.n2079 0.110872
R6395 VGND.n2075 VGND.n2074 0.110872
R6396 VGND.n2070 VGND.n2069 0.110872
R6397 VGND.n1828 VGND.n1827 0.110872
R6398 VGND.n1822 VGND.n1821 0.110872
R6399 VGND.n1817 VGND.n1816 0.110872
R6400 VGND.n1741 VGND.n1740 0.110872
R6401 VGND.n1806 VGND.n1805 0.110872
R6402 VGND.n1744 VGND.n1743 0.110872
R6403 VGND.n1795 VGND.n1794 0.110872
R6404 VGND.n1747 VGND.n1746 0.110872
R6405 VGND.n1784 VGND.n1783 0.110872
R6406 VGND.n1750 VGND.n1749 0.110872
R6407 VGND.n1773 VGND.n1772 0.110872
R6408 VGND.n1753 VGND.n1752 0.110872
R6409 VGND.n1762 VGND.n1761 0.110872
R6410 VGND.n1757 VGND.n1756 0.110872
R6411 VGND.n2177 VGND.n2176 0.110872
R6412 VGND.n1835 VGND.n1834 0.110872
R6413 VGND.n1841 VGND.n1840 0.110872
R6414 VGND.n1846 VGND.n1845 0.110872
R6415 VGND.n1673 VGND.n1672 0.110872
R6416 VGND.n1730 VGND.n1729 0.110872
R6417 VGND.n1725 VGND.n1724 0.110872
R6418 VGND.n1720 VGND.n1719 0.110872
R6419 VGND.n1715 VGND.n1714 0.110872
R6420 VGND.n1710 VGND.n1709 0.110872
R6421 VGND.n1705 VGND.n1704 0.110872
R6422 VGND.n1700 VGND.n1699 0.110872
R6423 VGND.n1695 VGND.n1694 0.110872
R6424 VGND.n1690 VGND.n1689 0.110872
R6425 VGND.n1676 VGND.n1675 0.110872
R6426 VGND.n1679 VGND.n1678 0.110872
R6427 VGND.n2866 VGND.n2865 0.110872
R6428 VGND.n2860 VGND.n2859 0.110872
R6429 VGND.n725 VGND.n724 0.110872
R6430 VGND.n667 VGND.n666 0.110872
R6431 VGND.n720 VGND.n719 0.110872
R6432 VGND.n715 VGND.n714 0.110872
R6433 VGND.n710 VGND.n709 0.110872
R6434 VGND.n705 VGND.n704 0.110872
R6435 VGND.n700 VGND.n699 0.110872
R6436 VGND.n695 VGND.n694 0.110872
R6437 VGND.n690 VGND.n689 0.110872
R6438 VGND.n685 VGND.n684 0.110872
R6439 VGND.n680 VGND.n679 0.110872
R6440 VGND.n675 VGND.n674 0.110872
R6441 VGND.n670 VGND.n669 0.110872
R6442 VGND.n1657 VGND.n1656 0.110872
R6443 VGND.n1662 VGND.n1661 0.110872
R6444 VGND.n735 VGND.n734 0.110872
R6445 VGND.n854 VGND.n853 0.110872
R6446 VGND.n820 VGND.n819 0.110872
R6447 VGND.n849 VGND.n848 0.110872
R6448 VGND.n844 VGND.n843 0.110872
R6449 VGND.n839 VGND.n838 0.110872
R6450 VGND.n834 VGND.n833 0.110872
R6451 VGND.n829 VGND.n828 0.110872
R6452 VGND.n824 VGND.n823 0.110872
R6453 VGND.n811 VGND.n810 0.110872
R6454 VGND.n870 VGND.n869 0.110872
R6455 VGND.n875 VGND.n874 0.110872
R6456 VGND.n1353 VGND.n1352 0.110872
R6457 VGND.n1649 VGND.n1648 0.110872
R6458 VGND.n1643 VGND.n1642 0.110872
R6459 VGND.n1638 VGND.n1637 0.110872
R6460 VGND.n1633 VGND.n1632 0.110872
R6461 VGND.n1553 VGND.n1552 0.110872
R6462 VGND.n761 VGND.n760 0.110872
R6463 VGND.n1548 VGND.n1547 0.110872
R6464 VGND.n1543 VGND.n1542 0.110872
R6465 VGND.n769 VGND.n768 0.110872
R6466 VGND.n1517 VGND.n1516 0.110872
R6467 VGND.n777 VGND.n776 0.110872
R6468 VGND.n1491 VGND.n1490 0.110872
R6469 VGND.n805 VGND.n804 0.110872
R6470 VGND.n1396 VGND.n1395 0.110872
R6471 VGND.n1391 VGND.n1390 0.110872
R6472 VGND.n2891 VGND.n2890 0.110872
R6473 VGND.n2885 VGND.n2884 0.110872
R6474 VGND.n1572 VGND.n1571 0.110872
R6475 VGND.n1577 VGND.n1576 0.110872
R6476 VGND.n1582 VGND.n1581 0.110872
R6477 VGND.n756 VGND.n755 0.110872
R6478 VGND.n1567 VGND.n1566 0.110872
R6479 VGND.n765 VGND.n764 0.110872
R6480 VGND.n1530 VGND.n1529 0.110872
R6481 VGND.n773 VGND.n772 0.110872
R6482 VGND.n1504 VGND.n1503 0.110872
R6483 VGND.n781 VGND.n780 0.110872
R6484 VGND.n1478 VGND.n1477 0.110872
R6485 VGND.n795 VGND.n794 0.110872
R6486 VGND.n1411 VGND.n1410 0.110872
R6487 VGND.n1609 VGND.n1608 0.110872
R6488 VGND.n1614 VGND.n1613 0.110872
R6489 VGND.n750 VGND.n749 0.110872
R6490 VGND.n1601 VGND.n1600 0.110872
R6491 VGND.n1596 VGND.n1595 0.110872
R6492 VGND.n1459 VGND.n1458 0.110872
R6493 VGND.n791 VGND.n790 0.110872
R6494 VGND.n1454 VGND.n1453 0.110872
R6495 VGND.n1449 VGND.n1448 0.110872
R6496 VGND.n1444 VGND.n1443 0.110872
R6497 VGND.n1439 VGND.n1438 0.110872
R6498 VGND.n1434 VGND.n1433 0.110872
R6499 VGND.n1429 VGND.n1428 0.110872
R6500 VGND.n1424 VGND.n1423 0.110872
R6501 VGND.n885 VGND.n884 0.110872
R6502 VGND.n2911 VGND.n2910 0.110872
R6503 VGND.n2905 VGND.n2904 0.110872
R6504 VGND.n1049 VGND.n1048 0.110872
R6505 VGND.n1058 VGND.n1057 0.110872
R6506 VGND.n1053 VGND.n1052 0.110872
R6507 VGND.n1044 VGND.n1043 0.110872
R6508 VGND.n1070 VGND.n1069 0.110872
R6509 VGND.n1075 VGND.n1074 0.110872
R6510 VGND.n1080 VGND.n1079 0.110872
R6511 VGND.n1085 VGND.n1084 0.110872
R6512 VGND.n1090 VGND.n1089 0.110872
R6513 VGND.n1095 VGND.n1094 0.110872
R6514 VGND.n1029 VGND.n1028 0.110872
R6515 VGND.n1037 VGND.n1036 0.110872
R6516 VGND.n1032 VGND.n1031 0.110872
R6517 VGND.n1169 VGND.n1168 0.110872
R6518 VGND.n1173 VGND.n1172 0.110872
R6519 VGND.n1179 VGND.n1178 0.110872
R6520 VGND.n1186 VGND.n1185 0.110872
R6521 VGND.n1009 VGND.n1008 0.110872
R6522 VGND.n1205 VGND.n1204 0.110872
R6523 VGND.n1211 VGND.n1210 0.110872
R6524 VGND.n1218 VGND.n1217 0.110872
R6525 VGND.n1222 VGND.n1001 0.110872
R6526 VGND.n1244 VGND.n1243 0.110872
R6527 VGND.n1227 VGND.n1225 0.110872
R6528 VGND.n1237 VGND.n1236 0.110872
R6529 VGND.n1232 VGND.n1231 0.110872
R6530 VGND.n1275 VGND.n1274 0.110872
R6531 VGND.n1281 VGND.n1280 0.110872
R6532 VGND.n928 VGND.n927 0.110872
R6533 VGND.n987 VGND.n986 0.110872
R6534 VGND.n982 VGND.n981 0.110872
R6535 VGND.n977 VGND.n976 0.110872
R6536 VGND.n972 VGND.n971 0.110872
R6537 VGND.n967 VGND.n966 0.110872
R6538 VGND.n962 VGND.n961 0.110872
R6539 VGND.n957 VGND.n956 0.110872
R6540 VGND.n952 VGND.n951 0.110872
R6541 VGND.n947 VGND.n946 0.110872
R6542 VGND.n942 VGND.n941 0.110872
R6543 VGND.n937 VGND.n936 0.110872
R6544 VGND.n932 VGND.n931 0.110872
R6545 VGND.n895 VGND.n894 0.110872
R6546 VGND.n1333 VGND.n1332 0.110872
R6547 VGND.n1130 VGND 0.0981562
R6548 VGND.n2214 VGND 0.0981562
R6549 VGND.n1362 VGND 0.0981562
R6550 VGND.n19 VGND 0.0968542
R6551 VGND.n2952 VGND 0.0968542
R6552 VGND.n45 VGND 0.0968542
R6553 VGND VGND.n91 0.0968542
R6554 VGND VGND.n130 0.0968542
R6555 VGND VGND.n499 0.0968542
R6556 VGND VGND.n2280 0.0968542
R6557 VGND VGND.n535 0.0968542
R6558 VGND VGND.n2207 0.0968542
R6559 VGND.n2224 VGND 0.0968542
R6560 VGND.n2982 VGND 0.0968542
R6561 VGND.n2562 VGND 0.088625
R6562 VGND.n2633 VGND 0.0790114
R6563 VGND.n2695 VGND 0.0790114
R6564 VGND.n2690 VGND 0.0790114
R6565 VGND VGND.n2689 0.0790114
R6566 VGND.n2684 VGND 0.0790114
R6567 VGND VGND.n2683 0.0790114
R6568 VGND.n2678 VGND 0.0790114
R6569 VGND VGND.n2677 0.0790114
R6570 VGND.n2709 VGND 0.0790114
R6571 VGND.n2723 VGND 0.0790114
R6572 VGND.n2742 VGND 0.0790114
R6573 VGND.n2761 VGND 0.0790114
R6574 VGND.n2781 VGND 0.0790114
R6575 VGND VGND.n2780 0.0790114
R6576 VGND VGND.n284 0.0790114
R6577 VGND.n2940 VGND 0.0790114
R6578 VGND.n2635 VGND 0.0790114
R6579 VGND.n2693 VGND 0.0790114
R6580 VGND VGND.n2692 0.0790114
R6581 VGND.n2687 VGND 0.0790114
R6582 VGND VGND.n2686 0.0790114
R6583 VGND.n2681 VGND 0.0790114
R6584 VGND VGND.n2680 0.0790114
R6585 VGND.n2675 VGND 0.0790114
R6586 VGND.n2711 VGND 0.0790114
R6587 VGND.n2721 VGND 0.0790114
R6588 VGND.n2744 VGND 0.0790114
R6589 VGND.n2759 VGND 0.0790114
R6590 VGND.n2783 VGND 0.0790114
R6591 VGND.n2784 VGND 0.0790114
R6592 VGND.n2794 VGND 0.0790114
R6593 VGND.n2937 VGND 0.0790114
R6594 VGND VGND.n2559 0.0790114
R6595 VGND VGND.n2558 0.0790114
R6596 VGND VGND.n2557 0.0790114
R6597 VGND VGND.n2556 0.0790114
R6598 VGND VGND.n2555 0.0790114
R6599 VGND VGND.n2554 0.0790114
R6600 VGND VGND.n2553 0.0790114
R6601 VGND VGND.n2552 0.0790114
R6602 VGND VGND.n2551 0.0790114
R6603 VGND VGND.n2550 0.0790114
R6604 VGND VGND.n2549 0.0790114
R6605 VGND VGND.n2548 0.0790114
R6606 VGND VGND.n2547 0.0790114
R6607 VGND.n2798 VGND 0.0790114
R6608 VGND VGND.n2797 0.0790114
R6609 VGND.n2533 VGND 0.0790114
R6610 VGND.n2357 VGND 0.0790114
R6611 VGND.n2373 VGND 0.0790114
R6612 VGND.n2383 VGND 0.0790114
R6613 VGND.n2399 VGND 0.0790114
R6614 VGND.n2409 VGND 0.0790114
R6615 VGND.n2425 VGND 0.0790114
R6616 VGND.n2435 VGND 0.0790114
R6617 VGND.n2451 VGND 0.0790114
R6618 VGND.n2461 VGND 0.0790114
R6619 VGND.n2477 VGND 0.0790114
R6620 VGND.n2487 VGND 0.0790114
R6621 VGND.n2508 VGND 0.0790114
R6622 VGND.n2802 VGND 0.0790114
R6623 VGND VGND.n2801 0.0790114
R6624 VGND.n419 VGND 0.0790114
R6625 VGND.n2530 VGND 0.0790114
R6626 VGND.n2360 VGND 0.0790114
R6627 VGND.n2370 VGND 0.0790114
R6628 VGND.n2386 VGND 0.0790114
R6629 VGND.n2396 VGND 0.0790114
R6630 VGND.n2412 VGND 0.0790114
R6631 VGND.n2422 VGND 0.0790114
R6632 VGND.n2438 VGND 0.0790114
R6633 VGND.n2448 VGND 0.0790114
R6634 VGND.n2464 VGND 0.0790114
R6635 VGND.n2474 VGND 0.0790114
R6636 VGND.n2490 VGND 0.0790114
R6637 VGND.n2505 VGND 0.0790114
R6638 VGND.n2805 VGND 0.0790114
R6639 VGND.n2806 VGND 0.0790114
R6640 VGND.n2819 VGND 0.0790114
R6641 VGND VGND.n2818 0.0790114
R6642 VGND.n1907 VGND 0.0790114
R6643 VGND.n1917 VGND 0.0790114
R6644 VGND.n1918 VGND 0.0790114
R6645 VGND.n1928 VGND 0.0790114
R6646 VGND.n1929 VGND 0.0790114
R6647 VGND.n1939 VGND 0.0790114
R6648 VGND.n1940 VGND 0.0790114
R6649 VGND.n1950 VGND 0.0790114
R6650 VGND.n1951 VGND 0.0790114
R6651 VGND.n1961 VGND 0.0790114
R6652 VGND.n1962 VGND 0.0790114
R6653 VGND.n1972 VGND 0.0790114
R6654 VGND.n1973 VGND 0.0790114
R6655 VGND.n2823 VGND 0.0790114
R6656 VGND VGND.n2822 0.0790114
R6657 VGND.n1990 VGND 0.0790114
R6658 VGND.n2063 VGND 0.0790114
R6659 VGND VGND.n2062 0.0790114
R6660 VGND.n2167 VGND 0.0790114
R6661 VGND VGND.n2166 0.0790114
R6662 VGND.n2159 VGND 0.0790114
R6663 VGND VGND.n2158 0.0790114
R6664 VGND.n2151 VGND 0.0790114
R6665 VGND VGND.n2150 0.0790114
R6666 VGND.n2143 VGND 0.0790114
R6667 VGND VGND.n2142 0.0790114
R6668 VGND.n2135 VGND 0.0790114
R6669 VGND VGND.n2134 0.0790114
R6670 VGND.n2827 VGND 0.0790114
R6671 VGND VGND.n2826 0.0790114
R6672 VGND.n1998 VGND 0.0790114
R6673 VGND VGND.n1997 0.0790114
R6674 VGND.n2066 VGND 0.0790114
R6675 VGND.n2171 VGND 0.0790114
R6676 VGND VGND.n2170 0.0790114
R6677 VGND.n2163 VGND 0.0790114
R6678 VGND VGND.n2162 0.0790114
R6679 VGND.n2155 VGND 0.0790114
R6680 VGND VGND.n2154 0.0790114
R6681 VGND.n2147 VGND 0.0790114
R6682 VGND VGND.n2146 0.0790114
R6683 VGND.n2139 VGND 0.0790114
R6684 VGND VGND.n2138 0.0790114
R6685 VGND.n2131 VGND 0.0790114
R6686 VGND.n2830 VGND 0.0790114
R6687 VGND.n2831 VGND 0.0790114
R6688 VGND.n2844 VGND 0.0790114
R6689 VGND VGND.n2843 0.0790114
R6690 VGND VGND.n1901 0.0790114
R6691 VGND.n2174 VGND 0.0790114
R6692 VGND.n1758 VGND 0.0790114
R6693 VGND.n1768 VGND 0.0790114
R6694 VGND.n1769 VGND 0.0790114
R6695 VGND.n1779 VGND 0.0790114
R6696 VGND.n1780 VGND 0.0790114
R6697 VGND.n1790 VGND 0.0790114
R6698 VGND.n1791 VGND 0.0790114
R6699 VGND.n1801 VGND 0.0790114
R6700 VGND.n1802 VGND 0.0790114
R6701 VGND.n1812 VGND 0.0790114
R6702 VGND.n1813 VGND 0.0790114
R6703 VGND.n2848 VGND 0.0790114
R6704 VGND VGND.n2847 0.0790114
R6705 VGND.n1830 VGND 0.0790114
R6706 VGND VGND.n1899 0.0790114
R6707 VGND.n1685 VGND 0.0790114
R6708 VGND.n1686 VGND 0.0790114
R6709 VGND.n1884 VGND 0.0790114
R6710 VGND VGND.n1883 0.0790114
R6711 VGND.n1876 VGND 0.0790114
R6712 VGND VGND.n1875 0.0790114
R6713 VGND.n1868 VGND 0.0790114
R6714 VGND VGND.n1867 0.0790114
R6715 VGND.n1860 VGND 0.0790114
R6716 VGND VGND.n1859 0.0790114
R6717 VGND.n1852 VGND 0.0790114
R6718 VGND.n2852 VGND 0.0790114
R6719 VGND VGND.n2851 0.0790114
R6720 VGND.n1838 VGND 0.0790114
R6721 VGND VGND.n1837 0.0790114
R6722 VGND.n1896 VGND 0.0790114
R6723 VGND VGND.n1895 0.0790114
R6724 VGND.n1888 VGND 0.0790114
R6725 VGND VGND.n1887 0.0790114
R6726 VGND.n1880 VGND 0.0790114
R6727 VGND VGND.n1879 0.0790114
R6728 VGND.n1872 VGND 0.0790114
R6729 VGND VGND.n1871 0.0790114
R6730 VGND.n1864 VGND 0.0790114
R6731 VGND VGND.n1863 0.0790114
R6732 VGND.n1856 VGND 0.0790114
R6733 VGND VGND.n1855 0.0790114
R6734 VGND.n2855 VGND 0.0790114
R6735 VGND.n2856 VGND 0.0790114
R6736 VGND.n2869 VGND 0.0790114
R6737 VGND VGND.n2868 0.0790114
R6738 VGND.n1349 VGND 0.0790114
R6739 VGND.n1892 VGND 0.0790114
R6740 VGND VGND.n1891 0.0790114
R6741 VGND.n867 VGND 0.0790114
R6742 VGND VGND.n866 0.0790114
R6743 VGND VGND.n865 0.0790114
R6744 VGND VGND.n864 0.0790114
R6745 VGND VGND.n863 0.0790114
R6746 VGND VGND.n862 0.0790114
R6747 VGND VGND.n861 0.0790114
R6748 VGND VGND.n860 0.0790114
R6749 VGND.n1669 VGND 0.0790114
R6750 VGND VGND.n1668 0.0790114
R6751 VGND.n2873 VGND 0.0790114
R6752 VGND VGND.n2872 0.0790114
R6753 VGND.n1654 VGND 0.0790114
R6754 VGND.n1404 VGND 0.0790114
R6755 VGND VGND.n1403 0.0790114
R6756 VGND VGND.n1402 0.0790114
R6757 VGND.n1487 VGND 0.0790114
R6758 VGND.n1497 VGND 0.0790114
R6759 VGND.n1513 VGND 0.0790114
R6760 VGND.n1523 VGND 0.0790114
R6761 VGND.n1539 VGND 0.0790114
R6762 VGND.n1560 VGND 0.0790114
R6763 VGND VGND.n1559 0.0790114
R6764 VGND.n1628 VGND 0.0790114
R6765 VGND.n1629 VGND 0.0790114
R6766 VGND.n2877 VGND 0.0790114
R6767 VGND VGND.n2876 0.0790114
R6768 VGND.n740 VGND 0.0790114
R6769 VGND.n1651 VGND 0.0790114
R6770 VGND.n1407 VGND 0.0790114
R6771 VGND.n1417 VGND 0.0790114
R6772 VGND.n1474 VGND 0.0790114
R6773 VGND.n1484 VGND 0.0790114
R6774 VGND.n1500 VGND 0.0790114
R6775 VGND.n1510 VGND 0.0790114
R6776 VGND.n1526 VGND 0.0790114
R6777 VGND.n1536 VGND 0.0790114
R6778 VGND.n1563 VGND 0.0790114
R6779 VGND.n1588 VGND 0.0790114
R6780 VGND.n1625 VGND 0.0790114
R6781 VGND VGND.n1624 0.0790114
R6782 VGND.n2880 VGND 0.0790114
R6783 VGND.n2881 VGND 0.0790114
R6784 VGND.n2894 VGND 0.0790114
R6785 VGND VGND.n2893 0.0790114
R6786 VGND VGND.n1344 0.0790114
R6787 VGND.n1420 VGND 0.0790114
R6788 VGND.n1471 VGND 0.0790114
R6789 VGND VGND.n1470 0.0790114
R6790 VGND VGND.n1469 0.0790114
R6791 VGND VGND.n1468 0.0790114
R6792 VGND VGND.n1467 0.0790114
R6793 VGND VGND.n1466 0.0790114
R6794 VGND VGND.n1465 0.0790114
R6795 VGND.n1591 VGND 0.0790114
R6796 VGND.n1592 VGND 0.0790114
R6797 VGND.n1621 VGND 0.0790114
R6798 VGND VGND.n1620 0.0790114
R6799 VGND.n2898 VGND 0.0790114
R6800 VGND VGND.n2897 0.0790114
R6801 VGND.n1606 VGND 0.0790114
R6802 VGND.n1103 VGND 0.0790114
R6803 VGND VGND.n1102 0.0790114
R6804 VGND VGND.n1101 0.0790114
R6805 VGND.n1321 VGND 0.0790114
R6806 VGND VGND.n1320 0.0790114
R6807 VGND.n1313 VGND 0.0790114
R6808 VGND VGND.n1312 0.0790114
R6809 VGND.n1305 VGND 0.0790114
R6810 VGND VGND.n1304 0.0790114
R6811 VGND.n1067 VGND 0.0790114
R6812 VGND VGND.n1066 0.0790114
R6813 VGND VGND.n1065 0.0790114
R6814 VGND VGND.n1064 0.0790114
R6815 VGND.n2901 VGND 0.0790114
R6816 VGND.n233 VGND 0.0790114
R6817 VGND.n2913 VGND 0.0790114
R6818 VGND.n1163 VGND 0.0790114
R6819 VGND.n1328 VGND 0.0790114
R6820 VGND VGND.n1327 0.0790114
R6821 VGND.n898 VGND 0.0790114
R6822 VGND.n901 VGND 0.0790114
R6823 VGND.n904 VGND 0.0790114
R6824 VGND.n907 VGND 0.0790114
R6825 VGND.n910 VGND 0.0790114
R6826 VGND.n913 VGND 0.0790114
R6827 VGND.n1298 VGND 0.0790114
R6828 VGND VGND.n1297 0.0790114
R6829 VGND.n1292 VGND 0.0790114
R6830 VGND VGND.n1291 0.0790114
R6831 VGND.n1270 VGND 0.0790114
R6832 VGND.n1285 VGND 0.0790114
R6833 VGND VGND.n1284 0.0790114
R6834 VGND.n1161 VGND 0.0790114
R6835 VGND.n1330 VGND 0.0790114
R6836 VGND.n1325 VGND 0.0790114
R6837 VGND VGND.n1324 0.0790114
R6838 VGND.n1317 VGND 0.0790114
R6839 VGND VGND.n1316 0.0790114
R6840 VGND.n1309 VGND 0.0790114
R6841 VGND VGND.n1308 0.0790114
R6842 VGND.n1301 VGND 0.0790114
R6843 VGND VGND.n1300 0.0790114
R6844 VGND.n1295 VGND 0.0790114
R6845 VGND VGND.n1294 0.0790114
R6846 VGND.n1289 VGND 0.0790114
R6847 VGND VGND.n1288 0.0790114
R6848 VGND VGND.n1287 0.0790114
R6849 VGND.n2916 VGND 0.0790114
R6850 VGND.n2699 VGND.n2698 0.0656596
R6851 VGND.n357 VGND.n355 0.0656596
R6852 VGND.n364 VGND.n362 0.0656596
R6853 VGND.n368 VGND.n367 0.0656596
R6854 VGND.n375 VGND.n373 0.0656596
R6855 VGND.n379 VGND.n378 0.0656596
R6856 VGND.n386 VGND.n384 0.0656596
R6857 VGND.n387 VGND.n325 0.0656596
R6858 VGND.n326 VGND.n314 0.0656596
R6859 VGND.n2726 VGND.n309 0.0656596
R6860 VGND.n312 VGND.n311 0.0656596
R6861 VGND.n2735 VGND.n2734 0.0656596
R6862 VGND.n2730 VGND.n293 0.0656596
R6863 VGND.n296 VGND.n294 0.0656596
R6864 VGND.n2773 VGND.n203 0.0656596
R6865 VGND.n2606 VGND 0.063
R6866 VGND.n2603 VGND 0.063
R6867 VGND.n2600 VGND 0.063
R6868 VGND.n2597 VGND 0.063
R6869 VGND.n2594 VGND 0.063
R6870 VGND.n2591 VGND 0.063
R6871 VGND.n2588 VGND 0.063
R6872 VGND.n2585 VGND 0.063
R6873 VGND.n2582 VGND 0.063
R6874 VGND.n2579 VGND 0.063
R6875 VGND.n2576 VGND 0.063
R6876 VGND.n2573 VGND 0.063
R6877 VGND.n2570 VGND 0.063
R6878 VGND.n2567 VGND 0.063
R6879 VGND.n2564 VGND 0.063
R6880 VGND VGND.n31 0.0603958
R6881 VGND.n3009 VGND 0.0603958
R6882 VGND VGND.n3008 0.0603958
R6883 VGND.n192 VGND 0.0603958
R6884 VGND VGND.n191 0.0603958
R6885 VGND VGND.n2964 0.0603958
R6886 VGND.n2965 VGND 0.0603958
R6887 VGND VGND.n57 0.0603958
R6888 VGND.n64 VGND 0.0603958
R6889 VGND VGND.n63 0.0603958
R6890 VGND.n118 VGND 0.0603958
R6891 VGND.n119 VGND 0.0603958
R6892 VGND.n132 VGND 0.0603958
R6893 VGND VGND.n131 0.0603958
R6894 VGND.n127 VGND 0.0603958
R6895 VGND.n163 VGND 0.0603958
R6896 VGND VGND.n162 0.0603958
R6897 VGND.n1152 VGND 0.0603958
R6898 VGND.n1129 VGND 0.0603958
R6899 VGND VGND.n1128 0.0603958
R6900 VGND.n1125 VGND 0.0603958
R6901 VGND.n501 VGND 0.0603958
R6902 VGND VGND.n500 0.0603958
R6903 VGND.n483 VGND 0.0603958
R6904 VGND.n2282 VGND 0.0603958
R6905 VGND VGND.n2281 0.0603958
R6906 VGND.n2264 VGND 0.0603958
R6907 VGND.n537 VGND 0.0603958
R6908 VGND VGND.n536 0.0603958
R6909 VGND.n519 VGND 0.0603958
R6910 VGND.n2209 VGND 0.0603958
R6911 VGND VGND.n2208 0.0603958
R6912 VGND.n2201 VGND 0.0603958
R6913 VGND.n2198 VGND 0.0603958
R6914 VGND.n2193 VGND 0.0603958
R6915 VGND VGND.n2225 0.0603958
R6916 VGND.n2246 VGND 0.0603958
R6917 VGND VGND.n2245 0.0603958
R6918 VGND VGND.n1363 0.0603958
R6919 VGND.n1384 VGND 0.0603958
R6920 VGND VGND.n1383 0.0603958
R6921 VGND VGND.n2994 0.0603958
R6922 VGND.n2995 VGND 0.0603958
R6923 VGND.n2996 VGND 0.0603958
R6924 VGND.n2698 VGND 0.0574853
R6925 VGND.n357 VGND 0.0574853
R6926 VGND.n364 VGND 0.0574853
R6927 VGND.n367 VGND 0.0574853
R6928 VGND.n375 VGND 0.0574853
R6929 VGND.n378 VGND 0.0574853
R6930 VGND.n386 VGND 0.0574853
R6931 VGND.n325 VGND 0.0574853
R6932 VGND.n314 VGND 0.0574853
R6933 VGND.n309 VGND 0.0574853
R6934 VGND.n311 VGND 0.0574853
R6935 VGND.n2734 VGND 0.0574853
R6936 VGND.n293 VGND 0.0574853
R6937 VGND.n296 VGND 0.0574853
R6938 VGND.n203 VGND 0.0574853
R6939 VGND.n1021 VGND 0.0489375
R6940 VGND.n994 VGND 0.0489375
R6941 VGND.n2630 VGND 0.0489375
R6942 VGND.n204 VGND 0.0489375
R6943 VGND.n334 VGND 0.0489375
R6944 VGND.n2626 VGND 0.0489375
R6945 VGND.n2623 VGND 0.0489375
R6946 VGND.n2620 VGND 0.0489375
R6947 VGND.n2617 VGND 0.0489375
R6948 VGND.n2614 VGND 0.0489375
R6949 VGND.n2611 VGND 0.0489375
R6950 VGND.n322 VGND 0.0489375
R6951 VGND.n315 VGND 0.0489375
R6952 VGND.n306 VGND 0.0489375
R6953 VGND.n299 VGND 0.0489375
R6954 VGND.n2765 VGND 0.0489375
R6955 VGND.n290 VGND 0.0489375
R6956 VGND.n297 VGND 0.0489375
R6957 VGND.n1018 VGND 0.0489375
R6958 VGND.n1015 VGND 0.0489375
R6959 VGND.n1180 VGND 0.0489375
R6960 VGND.n1006 VGND 0.0489375
R6961 VGND.n1004 VGND 0.0489375
R6962 VGND.n1195 VGND 0.0489375
R6963 VGND.n1212 VGND 0.0489375
R6964 VGND.n1000 VGND 0.0489375
R6965 VGND.n1253 VGND 0.0489375
R6966 VGND.n1256 VGND 0.0489375
R6967 VGND.n1259 VGND 0.0489375
R6968 VGND.n1262 VGND 0.0489375
R6969 VGND.n998 VGND 0.0489375
R6970 VGND.n1265 VGND 0.0489375
R6971 VGND VGND.n330 0.037734
R6972 VGND.n286 VGND 0.037734
R6973 VGND.n2787 VGND 0.037734
R6974 VGND.n2752 VGND 0.037734
R6975 VGND.n303 VGND 0.037734
R6976 VGND.n2747 VGND 0.037734
R6977 VGND.n319 VGND 0.037734
R6978 VGND.n2714 VGND 0.037734
R6979 VGND.n393 VGND 0.037734
R6980 VGND.n2668 VGND 0.037734
R6981 VGND.n2663 VGND 0.037734
R6982 VGND.n2658 VGND 0.037734
R6983 VGND.n2653 VGND 0.037734
R6984 VGND.n2648 VGND 0.037734
R6985 VGND.n2643 VGND 0.037734
R6986 VGND.n2638 VGND 0.037734
R6987 VGND VGND.n396 0.037734
R6988 VGND.n2535 VGND 0.037734
R6989 VGND.n2540 VGND 0.037734
R6990 VGND.n414 VGND 0.037734
R6991 VGND.n2287 VGND 0.037734
R6992 VGND.n2292 VGND 0.037734
R6993 VGND.n2297 VGND 0.037734
R6994 VGND.n2302 VGND 0.037734
R6995 VGND.n2307 VGND 0.037734
R6996 VGND.n2312 VGND 0.037734
R6997 VGND.n2317 VGND 0.037734
R6998 VGND.n2322 VGND 0.037734
R6999 VGND.n2327 VGND 0.037734
R7000 VGND.n2332 VGND 0.037734
R7001 VGND.n2337 VGND 0.037734
R7002 VGND.n2342 VGND 0.037734
R7003 VGND VGND.n400 0.037734
R7004 VGND VGND.n2528 0.037734
R7005 VGND.n2521 VGND 0.037734
R7006 VGND.n2516 VGND 0.037734
R7007 VGND.n2511 VGND 0.037734
R7008 VGND.n427 VGND 0.037734
R7009 VGND.n2480 VGND 0.037734
R7010 VGND.n435 VGND 0.037734
R7011 VGND.n2454 VGND 0.037734
R7012 VGND.n443 VGND 0.037734
R7013 VGND.n2428 VGND 0.037734
R7014 VGND.n451 VGND 0.037734
R7015 VGND.n2402 VGND 0.037734
R7016 VGND.n459 VGND 0.037734
R7017 VGND.n2376 VGND 0.037734
R7018 VGND.n471 VGND 0.037734
R7019 VGND VGND.n469 0.037734
R7020 VGND VGND.n2816 0.037734
R7021 VGND.n2809 VGND 0.037734
R7022 VGND.n2498 VGND 0.037734
R7023 VGND.n423 VGND 0.037734
R7024 VGND.n2493 VGND 0.037734
R7025 VGND.n431 VGND 0.037734
R7026 VGND.n2467 VGND 0.037734
R7027 VGND.n439 VGND 0.037734
R7028 VGND.n2441 VGND 0.037734
R7029 VGND.n447 VGND 0.037734
R7030 VGND.n2415 VGND 0.037734
R7031 VGND.n455 VGND 0.037734
R7032 VGND.n2389 VGND 0.037734
R7033 VGND.n463 VGND 0.037734
R7034 VGND.n2363 VGND 0.037734
R7035 VGND VGND.n466 0.037734
R7036 VGND VGND.n1988 0.037734
R7037 VGND.n1981 VGND 0.037734
R7038 VGND.n1976 VGND 0.037734
R7039 VGND.n607 VGND 0.037734
R7040 VGND.n1965 VGND 0.037734
R7041 VGND.n610 VGND 0.037734
R7042 VGND.n1954 VGND 0.037734
R7043 VGND.n613 VGND 0.037734
R7044 VGND.n1943 VGND 0.037734
R7045 VGND.n616 VGND 0.037734
R7046 VGND.n1932 VGND 0.037734
R7047 VGND.n619 VGND 0.037734
R7048 VGND.n1921 VGND 0.037734
R7049 VGND.n622 VGND 0.037734
R7050 VGND.n1910 VGND 0.037734
R7051 VGND VGND.n625 0.037734
R7052 VGND VGND.n1995 0.037734
R7053 VGND.n2000 VGND 0.037734
R7054 VGND.n2005 VGND 0.037734
R7055 VGND.n2010 VGND 0.037734
R7056 VGND.n2015 VGND 0.037734
R7057 VGND.n2020 VGND 0.037734
R7058 VGND.n2025 VGND 0.037734
R7059 VGND.n2030 VGND 0.037734
R7060 VGND.n2035 VGND 0.037734
R7061 VGND.n2040 VGND 0.037734
R7062 VGND.n2045 VGND 0.037734
R7063 VGND.n2050 VGND 0.037734
R7064 VGND.n2055 VGND 0.037734
R7065 VGND.n593 VGND 0.037734
R7066 VGND.n596 VGND 0.037734
R7067 VGND VGND.n590 0.037734
R7068 VGND VGND.n2841 0.037734
R7069 VGND.n2834 VGND 0.037734
R7070 VGND.n2124 VGND 0.037734
R7071 VGND.n584 VGND 0.037734
R7072 VGND.n2119 VGND 0.037734
R7073 VGND.n2114 VGND 0.037734
R7074 VGND.n2109 VGND 0.037734
R7075 VGND.n2104 VGND 0.037734
R7076 VGND.n2099 VGND 0.037734
R7077 VGND.n2094 VGND 0.037734
R7078 VGND.n2089 VGND 0.037734
R7079 VGND.n2084 VGND 0.037734
R7080 VGND.n2079 VGND 0.037734
R7081 VGND.n2074 VGND 0.037734
R7082 VGND.n2069 VGND 0.037734
R7083 VGND VGND.n587 0.037734
R7084 VGND VGND.n1828 0.037734
R7085 VGND.n1821 VGND 0.037734
R7086 VGND.n1816 VGND 0.037734
R7087 VGND.n1740 VGND 0.037734
R7088 VGND.n1805 VGND 0.037734
R7089 VGND.n1743 VGND 0.037734
R7090 VGND.n1794 VGND 0.037734
R7091 VGND.n1746 VGND 0.037734
R7092 VGND.n1783 VGND 0.037734
R7093 VGND.n1749 VGND 0.037734
R7094 VGND.n1772 VGND 0.037734
R7095 VGND.n1752 VGND 0.037734
R7096 VGND.n1761 VGND 0.037734
R7097 VGND VGND.n1757 0.037734
R7098 VGND.n2176 VGND 0.037734
R7099 VGND VGND.n547 0.037734
R7100 VGND VGND.n1835 0.037734
R7101 VGND.n1840 VGND 0.037734
R7102 VGND.n1845 VGND 0.037734
R7103 VGND.n1672 VGND 0.037734
R7104 VGND.n1729 VGND 0.037734
R7105 VGND.n1724 VGND 0.037734
R7106 VGND.n1719 VGND 0.037734
R7107 VGND.n1714 VGND 0.037734
R7108 VGND.n1709 VGND 0.037734
R7109 VGND.n1704 VGND 0.037734
R7110 VGND.n1699 VGND 0.037734
R7111 VGND.n1694 VGND 0.037734
R7112 VGND.n1689 VGND 0.037734
R7113 VGND.n1675 VGND 0.037734
R7114 VGND.n1678 VGND 0.037734
R7115 VGND VGND.n628 0.037734
R7116 VGND VGND.n2866 0.037734
R7117 VGND.n2859 VGND 0.037734
R7118 VGND.n724 VGND 0.037734
R7119 VGND.n666 VGND 0.037734
R7120 VGND.n719 VGND 0.037734
R7121 VGND.n714 VGND 0.037734
R7122 VGND.n709 VGND 0.037734
R7123 VGND.n704 VGND 0.037734
R7124 VGND.n699 VGND 0.037734
R7125 VGND.n694 VGND 0.037734
R7126 VGND.n689 VGND 0.037734
R7127 VGND.n684 VGND 0.037734
R7128 VGND.n679 VGND 0.037734
R7129 VGND.n674 VGND 0.037734
R7130 VGND.n669 VGND 0.037734
R7131 VGND VGND.n632 0.037734
R7132 VGND.n1656 VGND 0.037734
R7133 VGND.n1661 VGND 0.037734
R7134 VGND.n734 VGND 0.037734
R7135 VGND.n853 VGND 0.037734
R7136 VGND.n819 VGND 0.037734
R7137 VGND.n848 VGND 0.037734
R7138 VGND.n843 VGND 0.037734
R7139 VGND.n838 VGND 0.037734
R7140 VGND.n833 VGND 0.037734
R7141 VGND.n828 VGND 0.037734
R7142 VGND.n823 VGND 0.037734
R7143 VGND VGND.n811 0.037734
R7144 VGND.n869 VGND 0.037734
R7145 VGND.n874 VGND 0.037734
R7146 VGND.n1352 VGND 0.037734
R7147 VGND VGND.n879 0.037734
R7148 VGND VGND.n1649 0.037734
R7149 VGND.n1642 VGND 0.037734
R7150 VGND.n1637 VGND 0.037734
R7151 VGND.n1632 VGND 0.037734
R7152 VGND.n1552 VGND 0.037734
R7153 VGND.n760 VGND 0.037734
R7154 VGND.n1547 VGND 0.037734
R7155 VGND.n1542 VGND 0.037734
R7156 VGND.n768 VGND 0.037734
R7157 VGND.n1516 VGND 0.037734
R7158 VGND.n776 VGND 0.037734
R7159 VGND.n1490 VGND 0.037734
R7160 VGND.n804 VGND 0.037734
R7161 VGND.n1395 VGND 0.037734
R7162 VGND.n1390 VGND 0.037734
R7163 VGND VGND.n800 0.037734
R7164 VGND VGND.n2891 0.037734
R7165 VGND.n2884 VGND 0.037734
R7166 VGND.n1571 VGND 0.037734
R7167 VGND.n1576 VGND 0.037734
R7168 VGND.n1581 VGND 0.037734
R7169 VGND.n755 VGND 0.037734
R7170 VGND.n1566 VGND 0.037734
R7171 VGND.n764 VGND 0.037734
R7172 VGND.n1529 VGND 0.037734
R7173 VGND.n772 VGND 0.037734
R7174 VGND.n1503 VGND 0.037734
R7175 VGND.n780 VGND 0.037734
R7176 VGND.n1477 VGND 0.037734
R7177 VGND.n794 VGND 0.037734
R7178 VGND.n1410 VGND 0.037734
R7179 VGND VGND.n797 0.037734
R7180 VGND.n1608 VGND 0.037734
R7181 VGND.n1613 VGND 0.037734
R7182 VGND.n749 VGND 0.037734
R7183 VGND.n1600 VGND 0.037734
R7184 VGND.n1595 VGND 0.037734
R7185 VGND.n1458 VGND 0.037734
R7186 VGND.n790 VGND 0.037734
R7187 VGND.n1453 VGND 0.037734
R7188 VGND.n1448 VGND 0.037734
R7189 VGND.n1443 VGND 0.037734
R7190 VGND.n1438 VGND 0.037734
R7191 VGND.n1433 VGND 0.037734
R7192 VGND.n1428 VGND 0.037734
R7193 VGND.n1423 VGND 0.037734
R7194 VGND.n884 VGND 0.037734
R7195 VGND VGND.n882 0.037734
R7196 VGND VGND.n2911 0.037734
R7197 VGND.n2904 VGND 0.037734
R7198 VGND.n1048 VGND 0.037734
R7199 VGND.n1057 VGND 0.037734
R7200 VGND.n1052 VGND 0.037734
R7201 VGND VGND.n1044 0.037734
R7202 VGND.n1069 VGND 0.037734
R7203 VGND.n1074 VGND 0.037734
R7204 VGND.n1079 VGND 0.037734
R7205 VGND.n1084 VGND 0.037734
R7206 VGND.n1089 VGND 0.037734
R7207 VGND.n1094 VGND 0.037734
R7208 VGND.n1028 VGND 0.037734
R7209 VGND.n1036 VGND 0.037734
R7210 VGND.n1031 VGND 0.037734
R7211 VGND VGND.n1024 0.037734
R7212 VGND VGND.n1014 0.037734
R7213 VGND VGND.n1169 0.037734
R7214 VGND.n1172 VGND 0.037734
R7215 VGND VGND.n1179 0.037734
R7216 VGND.n1185 VGND 0.037734
R7217 VGND.n1008 VGND 0.037734
R7218 VGND.n1204 VGND 0.037734
R7219 VGND VGND.n1211 0.037734
R7220 VGND.n1217 VGND 0.037734
R7221 VGND VGND.n1222 0.037734
R7222 VGND.n1243 VGND 0.037734
R7223 VGND VGND.n1227 0.037734
R7224 VGND.n1236 VGND 0.037734
R7225 VGND.n1231 VGND 0.037734
R7226 VGND.n1274 VGND 0.037734
R7227 VGND VGND.n1281 0.037734
R7228 VGND.n927 VGND 0.037734
R7229 VGND.n986 VGND 0.037734
R7230 VGND.n981 VGND 0.037734
R7231 VGND.n976 VGND 0.037734
R7232 VGND.n971 VGND 0.037734
R7233 VGND.n966 VGND 0.037734
R7234 VGND.n961 VGND 0.037734
R7235 VGND.n956 VGND 0.037734
R7236 VGND.n951 VGND 0.037734
R7237 VGND.n946 VGND 0.037734
R7238 VGND.n941 VGND 0.037734
R7239 VGND.n936 VGND 0.037734
R7240 VGND.n931 VGND 0.037734
R7241 VGND VGND.n895 0.037734
R7242 VGND.n1332 VGND 0.037734
R7243 VGND VGND.n887 0.037734
R7244 VGND.n1156 VGND 0.0343542
R7245 VGND.n1128 VGND 0.0343542
R7246 VGND.n501 VGND 0.0343542
R7247 VGND.n2282 VGND 0.0343542
R7248 VGND.n537 VGND 0.0343542
R7249 VGND.n2209 VGND 0.0343542
R7250 VGND.n2246 VGND 0.0343542
R7251 VGND.n1384 VGND 0.0343542
R7252 VGND.n3009 VGND 0.0330521
R7253 VGND.n192 VGND 0.0330521
R7254 VGND.n2965 VGND 0.0330521
R7255 VGND.n64 VGND 0.0330521
R7256 VGND VGND.n118 0.0330521
R7257 VGND.n132 VGND 0.0330521
R7258 VGND.n163 VGND 0.0330521
R7259 VGND VGND.n2995 0.0330521
R7260 VGND.n33 VGND 0.024
R7261 VGND.n1 VGND 0.024
R7262 VGND.n119 VGND 0.0239375
R7263 VGND.n131 VGND 0.0239375
R7264 VGND.n500 VGND 0.0239375
R7265 VGND.n2281 VGND 0.0239375
R7266 VGND.n536 VGND 0.0239375
R7267 VGND.n3003 VGND 0.0226354
R7268 VGND VGND.n124 0.0226354
R7269 VGND.n1133 VGND 0.0226354
R7270 VGND VGND.n2256 0.0226354
R7271 VGND.n2217 VGND 0.0226354
R7272 VGND.n2208 VGND 0.0226354
R7273 VGND.n2220 VGND 0.0226354
R7274 VGND VGND.n3000 0.0226354
R7275 VGND VGND.n189 0.0213333
R7276 VGND.n191 VGND 0.0213333
R7277 VGND.n58 VGND 0.0213333
R7278 VGND.n113 VGND 0.0213333
R7279 VGND VGND.n90 0.0213333
R7280 VGND VGND.n158 0.0213333
R7281 VGND.n162 VGND 0.0213333
R7282 VGND VGND.n511 0.0213333
R7283 VGND.n2213 VGND 0.0213333
R7284 VGND.n1358 VGND 0.0213333
R7285 VGND VGND.n3024 0.0193356
R7286 VGND.n33 VGND 0.0161667
R7287 VGND.n331 VGND 0.00980851
R7288 VGND.n2936 VGND 0.00980851
R7289 VGND.n2793 VGND 0.00980851
R7290 VGND.n2785 VGND 0.00980851
R7291 VGND VGND.n288 0.00980851
R7292 VGND.n2758 VGND 0.00980851
R7293 VGND.n2745 VGND 0.00980851
R7294 VGND.n2720 VGND 0.00980851
R7295 VGND.n2712 VGND 0.00980851
R7296 VGND.n2674 VGND 0.00980851
R7297 VGND VGND.n350 0.00980851
R7298 VGND VGND.n349 0.00980851
R7299 VGND VGND.n344 0.00980851
R7300 VGND VGND.n343 0.00980851
R7301 VGND VGND.n338 0.00980851
R7302 VGND VGND.n337 0.00980851
R7303 VGND.n2636 VGND 0.00980851
R7304 VGND VGND.n2534 0.00980851
R7305 VGND VGND.n283 0.00980851
R7306 VGND VGND.n282 0.00980851
R7307 VGND.n2546 VGND 0.00980851
R7308 VGND VGND.n412 0.00980851
R7309 VGND VGND.n411 0.00980851
R7310 VGND VGND.n410 0.00980851
R7311 VGND VGND.n409 0.00980851
R7312 VGND VGND.n408 0.00980851
R7313 VGND VGND.n407 0.00980851
R7314 VGND VGND.n406 0.00980851
R7315 VGND VGND.n405 0.00980851
R7316 VGND VGND.n404 0.00980851
R7317 VGND VGND.n403 0.00980851
R7318 VGND VGND.n402 0.00980851
R7319 VGND.n401 VGND 0.00980851
R7320 VGND.n2529 VGND 0.00980851
R7321 VGND VGND.n420 0.00980851
R7322 VGND VGND.n280 0.00980851
R7323 VGND VGND.n279 0.00980851
R7324 VGND.n2509 VGND 0.00980851
R7325 VGND.n2486 VGND 0.00980851
R7326 VGND.n2478 VGND 0.00980851
R7327 VGND.n2460 VGND 0.00980851
R7328 VGND.n2452 VGND 0.00980851
R7329 VGND.n2434 VGND 0.00980851
R7330 VGND.n2426 VGND 0.00980851
R7331 VGND.n2408 VGND 0.00980851
R7332 VGND.n2400 VGND 0.00980851
R7333 VGND.n2382 VGND 0.00980851
R7334 VGND.n2374 VGND 0.00980851
R7335 VGND.n2356 VGND 0.00980851
R7336 VGND.n2817 VGND 0.00980851
R7337 VGND VGND.n273 0.00980851
R7338 VGND.n2807 VGND 0.00980851
R7339 VGND VGND.n277 0.00980851
R7340 VGND.n2504 VGND 0.00980851
R7341 VGND.n2491 VGND 0.00980851
R7342 VGND.n2473 VGND 0.00980851
R7343 VGND.n2465 VGND 0.00980851
R7344 VGND.n2447 VGND 0.00980851
R7345 VGND.n2439 VGND 0.00980851
R7346 VGND.n2421 VGND 0.00980851
R7347 VGND.n2413 VGND 0.00980851
R7348 VGND.n2395 VGND 0.00980851
R7349 VGND.n2387 VGND 0.00980851
R7350 VGND.n2369 VGND 0.00980851
R7351 VGND.n2361 VGND 0.00980851
R7352 VGND.n1989 VGND 0.00980851
R7353 VGND VGND.n271 0.00980851
R7354 VGND VGND.n270 0.00980851
R7355 VGND.n1974 VGND 0.00980851
R7356 VGND.n1971 VGND 0.00980851
R7357 VGND.n1963 VGND 0.00980851
R7358 VGND.n1960 VGND 0.00980851
R7359 VGND.n1952 VGND 0.00980851
R7360 VGND.n1949 VGND 0.00980851
R7361 VGND.n1941 VGND 0.00980851
R7362 VGND.n1938 VGND 0.00980851
R7363 VGND.n1930 VGND 0.00980851
R7364 VGND.n1927 VGND 0.00980851
R7365 VGND.n1919 VGND 0.00980851
R7366 VGND.n1916 VGND 0.00980851
R7367 VGND.n1908 VGND 0.00980851
R7368 VGND.n1996 VGND 0.00980851
R7369 VGND VGND.n1999 0.00980851
R7370 VGND VGND.n268 0.00980851
R7371 VGND VGND.n267 0.00980851
R7372 VGND VGND.n581 0.00980851
R7373 VGND VGND.n580 0.00980851
R7374 VGND VGND.n575 0.00980851
R7375 VGND VGND.n574 0.00980851
R7376 VGND VGND.n569 0.00980851
R7377 VGND VGND.n568 0.00980851
R7378 VGND VGND.n563 0.00980851
R7379 VGND VGND.n562 0.00980851
R7380 VGND VGND.n557 0.00980851
R7381 VGND VGND.n556 0.00980851
R7382 VGND.n2061 VGND 0.00980851
R7383 VGND.n591 VGND 0.00980851
R7384 VGND.n2842 VGND 0.00980851
R7385 VGND VGND.n261 0.00980851
R7386 VGND.n2832 VGND 0.00980851
R7387 VGND VGND.n265 0.00980851
R7388 VGND.n2130 VGND 0.00980851
R7389 VGND VGND.n578 0.00980851
R7390 VGND VGND.n577 0.00980851
R7391 VGND VGND.n572 0.00980851
R7392 VGND VGND.n571 0.00980851
R7393 VGND VGND.n566 0.00980851
R7394 VGND VGND.n565 0.00980851
R7395 VGND VGND.n560 0.00980851
R7396 VGND VGND.n559 0.00980851
R7397 VGND VGND.n554 0.00980851
R7398 VGND VGND.n553 0.00980851
R7399 VGND.n2067 VGND 0.00980851
R7400 VGND.n1829 VGND 0.00980851
R7401 VGND VGND.n259 0.00980851
R7402 VGND VGND.n258 0.00980851
R7403 VGND.n1814 VGND 0.00980851
R7404 VGND.n1811 VGND 0.00980851
R7405 VGND.n1803 VGND 0.00980851
R7406 VGND.n1800 VGND 0.00980851
R7407 VGND.n1792 VGND 0.00980851
R7408 VGND.n1789 VGND 0.00980851
R7409 VGND.n1781 VGND 0.00980851
R7410 VGND.n1778 VGND 0.00980851
R7411 VGND.n1770 VGND 0.00980851
R7412 VGND.n1767 VGND 0.00980851
R7413 VGND.n1759 VGND 0.00980851
R7414 VGND VGND.n2175 0.00980851
R7415 VGND.n548 VGND 0.00980851
R7416 VGND.n1836 VGND 0.00980851
R7417 VGND VGND.n1839 0.00980851
R7418 VGND VGND.n256 0.00980851
R7419 VGND VGND.n255 0.00980851
R7420 VGND.n1851 VGND 0.00980851
R7421 VGND VGND.n662 0.00980851
R7422 VGND VGND.n661 0.00980851
R7423 VGND VGND.n656 0.00980851
R7424 VGND VGND.n655 0.00980851
R7425 VGND VGND.n650 0.00980851
R7426 VGND VGND.n649 0.00980851
R7427 VGND VGND.n644 0.00980851
R7428 VGND VGND.n643 0.00980851
R7429 VGND.n1687 VGND 0.00980851
R7430 VGND.n1684 VGND 0.00980851
R7431 VGND.n629 VGND 0.00980851
R7432 VGND.n2867 VGND 0.00980851
R7433 VGND VGND.n249 0.00980851
R7434 VGND.n2857 VGND 0.00980851
R7435 VGND VGND.n253 0.00980851
R7436 VGND.n730 VGND 0.00980851
R7437 VGND VGND.n664 0.00980851
R7438 VGND VGND.n659 0.00980851
R7439 VGND VGND.n658 0.00980851
R7440 VGND VGND.n653 0.00980851
R7441 VGND VGND.n652 0.00980851
R7442 VGND VGND.n647 0.00980851
R7443 VGND VGND.n646 0.00980851
R7444 VGND VGND.n641 0.00980851
R7445 VGND VGND.n640 0.00980851
R7446 VGND VGND.n634 0.00980851
R7447 VGND.n633 VGND 0.00980851
R7448 VGND VGND.n1655 0.00980851
R7449 VGND VGND.n247 0.00980851
R7450 VGND VGND.n246 0.00980851
R7451 VGND.n1667 VGND 0.00980851
R7452 VGND VGND.n732 0.00980851
R7453 VGND.n859 VGND 0.00980851
R7454 VGND VGND.n817 0.00980851
R7455 VGND VGND.n816 0.00980851
R7456 VGND VGND.n815 0.00980851
R7457 VGND VGND.n814 0.00980851
R7458 VGND VGND.n813 0.00980851
R7459 VGND.n812 VGND 0.00980851
R7460 VGND VGND.n868 0.00980851
R7461 VGND VGND.n637 0.00980851
R7462 VGND VGND.n636 0.00980851
R7463 VGND.n1350 VGND 0.00980851
R7464 VGND.n1650 VGND 0.00980851
R7465 VGND VGND.n741 0.00980851
R7466 VGND VGND.n244 0.00980851
R7467 VGND VGND.n243 0.00980851
R7468 VGND.n1630 VGND 0.00980851
R7469 VGND VGND.n742 0.00980851
R7470 VGND.n1558 VGND 0.00980851
R7471 VGND VGND.n758 0.00980851
R7472 VGND.n1540 VGND 0.00980851
R7473 VGND.n1522 VGND 0.00980851
R7474 VGND.n1514 VGND 0.00980851
R7475 VGND.n1496 VGND 0.00980851
R7476 VGND.n1488 VGND 0.00980851
R7477 VGND.n1401 VGND 0.00980851
R7478 VGND VGND.n802 0.00980851
R7479 VGND.n801 VGND 0.00980851
R7480 VGND.n2892 VGND 0.00980851
R7481 VGND VGND.n236 0.00980851
R7482 VGND.n2882 VGND 0.00980851
R7483 VGND VGND.n240 0.00980851
R7484 VGND VGND.n745 0.00980851
R7485 VGND VGND.n744 0.00980851
R7486 VGND.n1587 VGND 0.00980851
R7487 VGND.n1564 VGND 0.00980851
R7488 VGND.n1535 VGND 0.00980851
R7489 VGND.n1527 VGND 0.00980851
R7490 VGND.n1509 VGND 0.00980851
R7491 VGND.n1501 VGND 0.00980851
R7492 VGND.n1483 VGND 0.00980851
R7493 VGND.n1475 VGND 0.00980851
R7494 VGND.n1416 VGND 0.00980851
R7495 VGND.n1408 VGND 0.00980851
R7496 VGND VGND.n1607 0.00980851
R7497 VGND VGND.n232 0.00980851
R7498 VGND VGND.n231 0.00980851
R7499 VGND.n1619 VGND 0.00980851
R7500 VGND VGND.n747 0.00980851
R7501 VGND.n1593 VGND 0.00980851
R7502 VGND VGND.n751 0.00980851
R7503 VGND.n1464 VGND 0.00980851
R7504 VGND VGND.n788 0.00980851
R7505 VGND VGND.n787 0.00980851
R7506 VGND VGND.n786 0.00980851
R7507 VGND VGND.n785 0.00980851
R7508 VGND VGND.n784 0.00980851
R7509 VGND VGND.n783 0.00980851
R7510 VGND.n1421 VGND 0.00980851
R7511 VGND.n1343 VGND 0.00980851
R7512 VGND.n2912 VGND 0.00980851
R7513 VGND VGND.n228 0.00980851
R7514 VGND.n2902 VGND 0.00980851
R7515 VGND.n1063 VGND 0.00980851
R7516 VGND VGND.n1046 0.00980851
R7517 VGND.n1045 VGND 0.00980851
R7518 VGND VGND.n1068 0.00980851
R7519 VGND VGND.n912 0.00980851
R7520 VGND VGND.n911 0.00980851
R7521 VGND VGND.n906 0.00980851
R7522 VGND VGND.n905 0.00980851
R7523 VGND VGND.n900 0.00980851
R7524 VGND VGND.n899 0.00980851
R7525 VGND.n1100 VGND 0.00980851
R7526 VGND VGND.n1026 0.00980851
R7527 VGND.n1025 VGND 0.00980851
R7528 VGND.n1165 VGND 0.00980851
R7529 VGND.n1170 VGND 0.00980851
R7530 VGND VGND.n1011 0.00980851
R7531 VGND.n1183 VGND 0.00980851
R7532 VGND.n1191 VGND 0.00980851
R7533 VGND.n1202 VGND 0.00980851
R7534 VGND VGND.n1003 0.00980851
R7535 VGND.n1215 VGND 0.00980851
R7536 VGND.n1249 VGND 0.00980851
R7537 VGND.n1223 VGND 0.00980851
R7538 VGND VGND.n1242 0.00980851
R7539 VGND.n1228 VGND 0.00980851
R7540 VGND VGND.n1235 0.00980851
R7541 VGND.n1272 VGND 0.00980851
R7542 VGND VGND.n997 0.00980851
R7543 VGND.n1282 VGND 0.00980851
R7544 VGND.n2917 VGND 0.00980851
R7545 VGND.n992 VGND 0.00980851
R7546 VGND VGND.n925 0.00980851
R7547 VGND VGND.n924 0.00980851
R7548 VGND VGND.n920 0.00980851
R7549 VGND VGND.n919 0.00980851
R7550 VGND VGND.n915 0.00980851
R7551 VGND VGND.n914 0.00980851
R7552 VGND VGND.n909 0.00980851
R7553 VGND VGND.n908 0.00980851
R7554 VGND VGND.n903 0.00980851
R7555 VGND VGND.n902 0.00980851
R7556 VGND VGND.n897 0.00980851
R7557 VGND.n896 VGND 0.00980851
R7558 VGND VGND.n1331 0.00980851
R7559 VGND.n888 VGND 0.00980851
R7560 VGND.n2698 VGND.n2697 0.00182979
R7561 VGND.n358 VGND.n357 0.00182979
R7562 VGND.n365 VGND.n364 0.00182979
R7563 VGND.n367 VGND.n354 0.00182979
R7564 VGND.n376 VGND.n375 0.00182979
R7565 VGND.n378 VGND.n353 0.00182979
R7566 VGND.n389 VGND.n386 0.00182979
R7567 VGND.n2707 VGND.n325 0.00182979
R7568 VGND.n2725 VGND.n314 0.00182979
R7569 VGND.n2740 VGND.n309 0.00182979
R7570 VGND.n311 VGND.n300 0.00182979
R7571 VGND.n2734 VGND.n2733 0.00182979
R7572 VGND.n2778 VGND.n293 0.00182979
R7573 VGND.n2772 VGND.n296 0.00182979
R7574 VGND.n2942 VGND.n203 0.00182979
R7575 XThR.Tn[2].n2 XThR.Tn[2].n1 332.332
R7576 XThR.Tn[2].n2 XThR.Tn[2].n0 296.493
R7577 XThR.Tn[2] XThR.Tn[2].n82 161.363
R7578 XThR.Tn[2] XThR.Tn[2].n77 161.363
R7579 XThR.Tn[2] XThR.Tn[2].n72 161.363
R7580 XThR.Tn[2] XThR.Tn[2].n67 161.363
R7581 XThR.Tn[2] XThR.Tn[2].n62 161.363
R7582 XThR.Tn[2] XThR.Tn[2].n57 161.363
R7583 XThR.Tn[2] XThR.Tn[2].n52 161.363
R7584 XThR.Tn[2] XThR.Tn[2].n47 161.363
R7585 XThR.Tn[2] XThR.Tn[2].n42 161.363
R7586 XThR.Tn[2] XThR.Tn[2].n37 161.363
R7587 XThR.Tn[2] XThR.Tn[2].n32 161.363
R7588 XThR.Tn[2] XThR.Tn[2].n27 161.363
R7589 XThR.Tn[2] XThR.Tn[2].n22 161.363
R7590 XThR.Tn[2] XThR.Tn[2].n17 161.363
R7591 XThR.Tn[2] XThR.Tn[2].n12 161.363
R7592 XThR.Tn[2] XThR.Tn[2].n10 161.363
R7593 XThR.Tn[2].n84 XThR.Tn[2].n83 161.3
R7594 XThR.Tn[2].n79 XThR.Tn[2].n78 161.3
R7595 XThR.Tn[2].n74 XThR.Tn[2].n73 161.3
R7596 XThR.Tn[2].n69 XThR.Tn[2].n68 161.3
R7597 XThR.Tn[2].n64 XThR.Tn[2].n63 161.3
R7598 XThR.Tn[2].n59 XThR.Tn[2].n58 161.3
R7599 XThR.Tn[2].n54 XThR.Tn[2].n53 161.3
R7600 XThR.Tn[2].n49 XThR.Tn[2].n48 161.3
R7601 XThR.Tn[2].n44 XThR.Tn[2].n43 161.3
R7602 XThR.Tn[2].n39 XThR.Tn[2].n38 161.3
R7603 XThR.Tn[2].n34 XThR.Tn[2].n33 161.3
R7604 XThR.Tn[2].n29 XThR.Tn[2].n28 161.3
R7605 XThR.Tn[2].n24 XThR.Tn[2].n23 161.3
R7606 XThR.Tn[2].n19 XThR.Tn[2].n18 161.3
R7607 XThR.Tn[2].n14 XThR.Tn[2].n13 161.3
R7608 XThR.Tn[2].n82 XThR.Tn[2].t65 161.106
R7609 XThR.Tn[2].n77 XThR.Tn[2].t72 161.106
R7610 XThR.Tn[2].n72 XThR.Tn[2].t51 161.106
R7611 XThR.Tn[2].n67 XThR.Tn[2].t36 161.106
R7612 XThR.Tn[2].n62 XThR.Tn[2].t64 161.106
R7613 XThR.Tn[2].n57 XThR.Tn[2].t26 161.106
R7614 XThR.Tn[2].n52 XThR.Tn[2].t69 161.106
R7615 XThR.Tn[2].n47 XThR.Tn[2].t49 161.106
R7616 XThR.Tn[2].n42 XThR.Tn[2].t35 161.106
R7617 XThR.Tn[2].n37 XThR.Tn[2].t41 161.106
R7618 XThR.Tn[2].n32 XThR.Tn[2].t25 161.106
R7619 XThR.Tn[2].n27 XThR.Tn[2].t50 161.106
R7620 XThR.Tn[2].n22 XThR.Tn[2].t23 161.106
R7621 XThR.Tn[2].n17 XThR.Tn[2].t67 161.106
R7622 XThR.Tn[2].n12 XThR.Tn[2].t31 161.106
R7623 XThR.Tn[2].n10 XThR.Tn[2].t14 161.106
R7624 XThR.Tn[2].n83 XThR.Tn[2].t38 159.978
R7625 XThR.Tn[2].n78 XThR.Tn[2].t46 159.978
R7626 XThR.Tn[2].n73 XThR.Tn[2].t29 159.978
R7627 XThR.Tn[2].n68 XThR.Tn[2].t13 159.978
R7628 XThR.Tn[2].n63 XThR.Tn[2].t37 159.978
R7629 XThR.Tn[2].n58 XThR.Tn[2].t63 159.978
R7630 XThR.Tn[2].n53 XThR.Tn[2].t45 159.978
R7631 XThR.Tn[2].n48 XThR.Tn[2].t27 159.978
R7632 XThR.Tn[2].n43 XThR.Tn[2].t12 159.978
R7633 XThR.Tn[2].n38 XThR.Tn[2].t20 159.978
R7634 XThR.Tn[2].n33 XThR.Tn[2].t62 159.978
R7635 XThR.Tn[2].n28 XThR.Tn[2].t28 159.978
R7636 XThR.Tn[2].n23 XThR.Tn[2].t60 159.978
R7637 XThR.Tn[2].n18 XThR.Tn[2].t43 159.978
R7638 XThR.Tn[2].n13 XThR.Tn[2].t66 159.978
R7639 XThR.Tn[2].n82 XThR.Tn[2].t53 145.038
R7640 XThR.Tn[2].n77 XThR.Tn[2].t19 145.038
R7641 XThR.Tn[2].n72 XThR.Tn[2].t59 145.038
R7642 XThR.Tn[2].n67 XThR.Tn[2].t42 145.038
R7643 XThR.Tn[2].n62 XThR.Tn[2].t73 145.038
R7644 XThR.Tn[2].n57 XThR.Tn[2].t52 145.038
R7645 XThR.Tn[2].n52 XThR.Tn[2].t61 145.038
R7646 XThR.Tn[2].n47 XThR.Tn[2].t44 145.038
R7647 XThR.Tn[2].n42 XThR.Tn[2].t39 145.038
R7648 XThR.Tn[2].n37 XThR.Tn[2].t70 145.038
R7649 XThR.Tn[2].n32 XThR.Tn[2].t34 145.038
R7650 XThR.Tn[2].n27 XThR.Tn[2].t58 145.038
R7651 XThR.Tn[2].n22 XThR.Tn[2].t32 145.038
R7652 XThR.Tn[2].n17 XThR.Tn[2].t15 145.038
R7653 XThR.Tn[2].n12 XThR.Tn[2].t40 145.038
R7654 XThR.Tn[2].n10 XThR.Tn[2].t21 145.038
R7655 XThR.Tn[2].n83 XThR.Tn[2].t71 143.911
R7656 XThR.Tn[2].n78 XThR.Tn[2].t33 143.911
R7657 XThR.Tn[2].n73 XThR.Tn[2].t17 143.911
R7658 XThR.Tn[2].n68 XThR.Tn[2].t56 143.911
R7659 XThR.Tn[2].n63 XThR.Tn[2].t24 143.911
R7660 XThR.Tn[2].n58 XThR.Tn[2].t68 143.911
R7661 XThR.Tn[2].n53 XThR.Tn[2].t18 143.911
R7662 XThR.Tn[2].n48 XThR.Tn[2].t57 143.911
R7663 XThR.Tn[2].n43 XThR.Tn[2].t54 143.911
R7664 XThR.Tn[2].n38 XThR.Tn[2].t22 143.911
R7665 XThR.Tn[2].n33 XThR.Tn[2].t48 143.911
R7666 XThR.Tn[2].n28 XThR.Tn[2].t16 143.911
R7667 XThR.Tn[2].n23 XThR.Tn[2].t47 143.911
R7668 XThR.Tn[2].n18 XThR.Tn[2].t30 143.911
R7669 XThR.Tn[2].n13 XThR.Tn[2].t55 143.911
R7670 XThR.Tn[2].n6 XThR.Tn[2].n4 135.249
R7671 XThR.Tn[2].n9 XThR.Tn[2].n3 98.982
R7672 XThR.Tn[2].n6 XThR.Tn[2].n5 98.982
R7673 XThR.Tn[2].n8 XThR.Tn[2].n7 98.982
R7674 XThR.Tn[2].n8 XThR.Tn[2].n6 36.2672
R7675 XThR.Tn[2].n9 XThR.Tn[2].n8 36.2672
R7676 XThR.Tn[2].n88 XThR.Tn[2].n9 32.6405
R7677 XThR.Tn[2].n1 XThR.Tn[2].t4 26.5955
R7678 XThR.Tn[2].n1 XThR.Tn[2].t2 26.5955
R7679 XThR.Tn[2].n0 XThR.Tn[2].t11 26.5955
R7680 XThR.Tn[2].n0 XThR.Tn[2].t5 26.5955
R7681 XThR.Tn[2].n3 XThR.Tn[2].t3 24.9236
R7682 XThR.Tn[2].n3 XThR.Tn[2].t6 24.9236
R7683 XThR.Tn[2].n4 XThR.Tn[2].t9 24.9236
R7684 XThR.Tn[2].n4 XThR.Tn[2].t10 24.9236
R7685 XThR.Tn[2].n5 XThR.Tn[2].t8 24.9236
R7686 XThR.Tn[2].n5 XThR.Tn[2].t7 24.9236
R7687 XThR.Tn[2].n7 XThR.Tn[2].t1 24.9236
R7688 XThR.Tn[2].n7 XThR.Tn[2].t0 24.9236
R7689 XThR.Tn[2] XThR.Tn[2].n2 23.3605
R7690 XThR.Tn[2] XThR.Tn[2].n88 6.7205
R7691 XThR.Tn[2].n88 XThR.Tn[2] 6.30883
R7692 XThR.Tn[2] XThR.Tn[2].n11 5.34038
R7693 XThR.Tn[2].n16 XThR.Tn[2].n15 4.5005
R7694 XThR.Tn[2].n21 XThR.Tn[2].n20 4.5005
R7695 XThR.Tn[2].n26 XThR.Tn[2].n25 4.5005
R7696 XThR.Tn[2].n31 XThR.Tn[2].n30 4.5005
R7697 XThR.Tn[2].n36 XThR.Tn[2].n35 4.5005
R7698 XThR.Tn[2].n41 XThR.Tn[2].n40 4.5005
R7699 XThR.Tn[2].n46 XThR.Tn[2].n45 4.5005
R7700 XThR.Tn[2].n51 XThR.Tn[2].n50 4.5005
R7701 XThR.Tn[2].n56 XThR.Tn[2].n55 4.5005
R7702 XThR.Tn[2].n61 XThR.Tn[2].n60 4.5005
R7703 XThR.Tn[2].n66 XThR.Tn[2].n65 4.5005
R7704 XThR.Tn[2].n71 XThR.Tn[2].n70 4.5005
R7705 XThR.Tn[2].n76 XThR.Tn[2].n75 4.5005
R7706 XThR.Tn[2].n81 XThR.Tn[2].n80 4.5005
R7707 XThR.Tn[2].n86 XThR.Tn[2].n85 4.5005
R7708 XThR.Tn[2].n87 XThR.Tn[2] 3.70586
R7709 XThR.Tn[2].n16 XThR.Tn[2] 2.52282
R7710 XThR.Tn[2].n21 XThR.Tn[2] 2.52282
R7711 XThR.Tn[2].n26 XThR.Tn[2] 2.52282
R7712 XThR.Tn[2].n31 XThR.Tn[2] 2.52282
R7713 XThR.Tn[2].n36 XThR.Tn[2] 2.52282
R7714 XThR.Tn[2].n41 XThR.Tn[2] 2.52282
R7715 XThR.Tn[2].n46 XThR.Tn[2] 2.52282
R7716 XThR.Tn[2].n51 XThR.Tn[2] 2.52282
R7717 XThR.Tn[2].n56 XThR.Tn[2] 2.52282
R7718 XThR.Tn[2].n61 XThR.Tn[2] 2.52282
R7719 XThR.Tn[2].n66 XThR.Tn[2] 2.52282
R7720 XThR.Tn[2].n71 XThR.Tn[2] 2.52282
R7721 XThR.Tn[2].n76 XThR.Tn[2] 2.52282
R7722 XThR.Tn[2].n81 XThR.Tn[2] 2.52282
R7723 XThR.Tn[2].n86 XThR.Tn[2] 2.52282
R7724 XThR.Tn[2].n84 XThR.Tn[2] 1.08677
R7725 XThR.Tn[2].n79 XThR.Tn[2] 1.08677
R7726 XThR.Tn[2].n74 XThR.Tn[2] 1.08677
R7727 XThR.Tn[2].n69 XThR.Tn[2] 1.08677
R7728 XThR.Tn[2].n64 XThR.Tn[2] 1.08677
R7729 XThR.Tn[2].n59 XThR.Tn[2] 1.08677
R7730 XThR.Tn[2].n54 XThR.Tn[2] 1.08677
R7731 XThR.Tn[2].n49 XThR.Tn[2] 1.08677
R7732 XThR.Tn[2].n44 XThR.Tn[2] 1.08677
R7733 XThR.Tn[2].n39 XThR.Tn[2] 1.08677
R7734 XThR.Tn[2].n34 XThR.Tn[2] 1.08677
R7735 XThR.Tn[2].n29 XThR.Tn[2] 1.08677
R7736 XThR.Tn[2].n24 XThR.Tn[2] 1.08677
R7737 XThR.Tn[2].n19 XThR.Tn[2] 1.08677
R7738 XThR.Tn[2].n14 XThR.Tn[2] 1.08677
R7739 XThR.Tn[2] XThR.Tn[2].n16 0.839786
R7740 XThR.Tn[2] XThR.Tn[2].n21 0.839786
R7741 XThR.Tn[2] XThR.Tn[2].n26 0.839786
R7742 XThR.Tn[2] XThR.Tn[2].n31 0.839786
R7743 XThR.Tn[2] XThR.Tn[2].n36 0.839786
R7744 XThR.Tn[2] XThR.Tn[2].n41 0.839786
R7745 XThR.Tn[2] XThR.Tn[2].n46 0.839786
R7746 XThR.Tn[2] XThR.Tn[2].n51 0.839786
R7747 XThR.Tn[2] XThR.Tn[2].n56 0.839786
R7748 XThR.Tn[2] XThR.Tn[2].n61 0.839786
R7749 XThR.Tn[2] XThR.Tn[2].n66 0.839786
R7750 XThR.Tn[2] XThR.Tn[2].n71 0.839786
R7751 XThR.Tn[2] XThR.Tn[2].n76 0.839786
R7752 XThR.Tn[2] XThR.Tn[2].n81 0.839786
R7753 XThR.Tn[2] XThR.Tn[2].n86 0.839786
R7754 XThR.Tn[2].n11 XThR.Tn[2] 0.499542
R7755 XThR.Tn[2].n85 XThR.Tn[2] 0.063
R7756 XThR.Tn[2].n80 XThR.Tn[2] 0.063
R7757 XThR.Tn[2].n75 XThR.Tn[2] 0.063
R7758 XThR.Tn[2].n70 XThR.Tn[2] 0.063
R7759 XThR.Tn[2].n65 XThR.Tn[2] 0.063
R7760 XThR.Tn[2].n60 XThR.Tn[2] 0.063
R7761 XThR.Tn[2].n55 XThR.Tn[2] 0.063
R7762 XThR.Tn[2].n50 XThR.Tn[2] 0.063
R7763 XThR.Tn[2].n45 XThR.Tn[2] 0.063
R7764 XThR.Tn[2].n40 XThR.Tn[2] 0.063
R7765 XThR.Tn[2].n35 XThR.Tn[2] 0.063
R7766 XThR.Tn[2].n30 XThR.Tn[2] 0.063
R7767 XThR.Tn[2].n25 XThR.Tn[2] 0.063
R7768 XThR.Tn[2].n20 XThR.Tn[2] 0.063
R7769 XThR.Tn[2].n15 XThR.Tn[2] 0.063
R7770 XThR.Tn[2].n87 XThR.Tn[2] 0.0540714
R7771 XThR.Tn[2] XThR.Tn[2].n87 0.038
R7772 XThR.Tn[2].n11 XThR.Tn[2] 0.0143889
R7773 XThR.Tn[2].n85 XThR.Tn[2].n84 0.00771154
R7774 XThR.Tn[2].n80 XThR.Tn[2].n79 0.00771154
R7775 XThR.Tn[2].n75 XThR.Tn[2].n74 0.00771154
R7776 XThR.Tn[2].n70 XThR.Tn[2].n69 0.00771154
R7777 XThR.Tn[2].n65 XThR.Tn[2].n64 0.00771154
R7778 XThR.Tn[2].n60 XThR.Tn[2].n59 0.00771154
R7779 XThR.Tn[2].n55 XThR.Tn[2].n54 0.00771154
R7780 XThR.Tn[2].n50 XThR.Tn[2].n49 0.00771154
R7781 XThR.Tn[2].n45 XThR.Tn[2].n44 0.00771154
R7782 XThR.Tn[2].n40 XThR.Tn[2].n39 0.00771154
R7783 XThR.Tn[2].n35 XThR.Tn[2].n34 0.00771154
R7784 XThR.Tn[2].n30 XThR.Tn[2].n29 0.00771154
R7785 XThR.Tn[2].n25 XThR.Tn[2].n24 0.00771154
R7786 XThR.Tn[2].n20 XThR.Tn[2].n19 0.00771154
R7787 XThR.Tn[2].n15 XThR.Tn[2].n14 0.00771154
R7788 VPWR.n2837 VPWR.n2823 2618.82
R7789 VPWR.n2835 VPWR.n2829 2618.82
R7790 VPWR.n2853 VPWR.n2823 1916.47
R7791 VPWR.n2828 VPWR.n2827 1916.47
R7792 VPWR.n2827 VPWR.n2821 1916.47
R7793 VPWR.n2829 VPWR.n2822 1916.47
R7794 VPWR.n2852 VPWR.n2824 1912.94
R7795 VPWR.n2849 VPWR.n2843 1560
R7796 VPWR.n2850 VPWR.n2824 1408.24
R7797 VPWR.n2853 VPWR.n2852 1210.59
R7798 VPWR.n2851 VPWR.n2821 1210.59
R7799 VPWR.n2380 VPWR.t1488 1005.7
R7800 VPWR.t1706 VPWR.n485 1005.7
R7801 VPWR.t1555 VPWR.n2210 1005.7
R7802 VPWR.n639 VPWR.t1663 1005.7
R7803 VPWR.n2184 VPWR.t1389 1005.7
R7804 VPWR.t1496 VPWR.n677 1005.7
R7805 VPWR.t1456 VPWR.n2014 1005.7
R7806 VPWR.n831 VPWR.t1561 1005.7
R7807 VPWR.n1988 VPWR.t1384 1005.7
R7808 VPWR.t1568 VPWR.n869 1005.7
R7809 VPWR.n447 VPWR.t1376 1005.7
R7810 VPWR.t1676 VPWR.n1818 1005.7
R7811 VPWR.t1658 VPWR.n2406 1005.7
R7812 VPWR.n1023 VPWR.t1528 1005.7
R7813 VPWR.t1698 VPWR.n293 1005.7
R7814 VPWR.n1792 VPWR.t1639 1005.7
R7815 VPWR.n2591 VPWR.t1590 1005.7
R7816 VPWR.n1062 VPWR.t1474 1005.7
R7817 VPWR.t957 VPWR.n2309 983.14
R7818 VPWR.n2310 VPWR.t1129 983.14
R7819 VPWR.t827 VPWR.n2319 983.14
R7820 VPWR.n2320 VPWR.t153 983.14
R7821 VPWR.t1121 VPWR.n2329 983.14
R7822 VPWR.n2330 VPWR.t1176 983.14
R7823 VPWR.t1256 VPWR.n2339 983.14
R7824 VPWR.n2340 VPWR.t736 983.14
R7825 VPWR.t579 VPWR.n2349 983.14
R7826 VPWR.n2350 VPWR.t431 983.14
R7827 VPWR.t1914 VPWR.n2359 983.14
R7828 VPWR.n2360 VPWR.t1780 983.14
R7829 VPWR.t545 VPWR.n2369 983.14
R7830 VPWR.n2370 VPWR.t883 983.14
R7831 VPWR.t181 VPWR.n2379 983.14
R7832 VPWR.n542 VPWR.t1020 983.14
R7833 VPWR.n541 VPWR.t1228 983.14
R7834 VPWR.n537 VPWR.t803 983.14
R7835 VPWR.n533 VPWR.t679 983.14
R7836 VPWR.n529 VPWR.t112 983.14
R7837 VPWR.n525 VPWR.t1816 983.14
R7838 VPWR.n521 VPWR.t1730 983.14
R7839 VPWR.n517 VPWR.t65 983.14
R7840 VPWR.n513 VPWR.t726 983.14
R7841 VPWR.n509 VPWR.t355 983.14
R7842 VPWR.n505 VPWR.t1828 983.14
R7843 VPWR.n501 VPWR.t96 983.14
R7844 VPWR.n497 VPWR.t1240 983.14
R7845 VPWR.n493 VPWR.t16 983.14
R7846 VPWR.n489 VPWR.t877 983.14
R7847 VPWR.n2281 VPWR.t1910 983.14
R7848 VPWR.n2280 VPWR.t259 983.14
R7849 VPWR.n2271 VPWR.t781 983.14
R7850 VPWR.n2270 VPWR.t1041 983.14
R7851 VPWR.n2261 VPWR.t1320 983.14
R7852 VPWR.n2260 VPWR.t557 983.14
R7853 VPWR.n2251 VPWR.t491 983.14
R7854 VPWR.n2250 VPWR.t849 983.14
R7855 VPWR.n2241 VPWR.t519 983.14
R7856 VPWR.n2240 VPWR.t587 983.14
R7857 VPWR.n2231 VPWR.t706 983.14
R7858 VPWR.n2230 VPWR.t1141 983.14
R7859 VPWR.n2221 VPWR.t971 983.14
R7860 VPWR.n2220 VPWR.t477 983.14
R7861 VPWR.n2211 VPWR.t203 983.14
R7862 VPWR.t897 VPWR.n582 983.14
R7863 VPWR.t1212 VPWR.n586 983.14
R7864 VPWR.t795 VPWR.n590 983.14
R7865 VPWR.t685 VPWR.n594 983.14
R7866 VPWR.t399 VPWR.n598 983.14
R7867 VPWR.t1756 VPWR.n602 983.14
R7868 VPWR.t1740 VPWR.n606 983.14
R7869 VPWR.t73 VPWR.n610 983.14
R7870 VPWR.t1898 VPWR.n614 983.14
R7871 VPWR.t361 VPWR.n618 983.14
R7872 VPWR.t529 VPWR.n622 983.14
R7873 VPWR.t1796 VPWR.n626 983.14
R7874 VPWR.t1248 VPWR.n630 983.14
R7875 VPWR.t33 VPWR.n634 983.14
R7876 VPWR.t1004 VPWR.n638 983.14
R7877 VPWR.t479 VPWR.n2113 983.14
R7878 VPWR.n2114 VPWR.t509 983.14
R7879 VPWR.t817 VPWR.n2123 983.14
R7880 VPWR.n2124 VPWR.t379 983.14
R7881 VPWR.t139 VPWR.n2133 983.14
R7882 VPWR.n2134 VPWR.t57 983.14
R7883 VPWR.t1861 VPWR.n2143 983.14
R7884 VPWR.n2144 VPWR.t595 983.14
R7885 VPWR.t1218 VPWR.n2153 983.14
R7886 VPWR.n2154 VPWR.t336 983.14
R7887 VPWR.t1837 VPWR.n2163 983.14
R7888 VPWR.n2164 VPWR.t919 983.14
R7889 VPWR.t1289 VPWR.n2173 983.14
R7890 VPWR.n2174 VPWR.t22 983.14
R7891 VPWR.t165 VPWR.n2183 983.14
R7892 VPWR.n734 VPWR.t620 983.14
R7893 VPWR.n733 VPWR.t767 983.14
R7894 VPWR.n729 VPWR.t829 983.14
R7895 VPWR.n725 VPWR.t151 983.14
R7896 VPWR.n721 VPWR.t1190 983.14
R7897 VPWR.n717 VPWR.t1174 983.14
R7898 VPWR.n713 VPWR.t1254 983.14
R7899 VPWR.n709 VPWR.t734 983.14
R7900 VPWR.n705 VPWR.t577 983.14
R7901 VPWR.n701 VPWR.t429 983.14
R7902 VPWR.n697 VPWR.t1912 983.14
R7903 VPWR.n693 VPWR.t1778 983.14
R7904 VPWR.n689 VPWR.t543 983.14
R7905 VPWR.n685 VPWR.t881 983.14
R7906 VPWR.n681 VPWR.t179 983.14
R7907 VPWR.n2085 VPWR.t1724 983.14
R7908 VPWR.n2084 VPWR.t1135 983.14
R7909 VPWR.n2075 VPWR.t823 983.14
R7910 VPWR.n2074 VPWR.t369 983.14
R7911 VPWR.n2065 VPWR.t1127 983.14
R7912 VPWR.n2064 VPWR.t1163 983.14
R7913 VPWR.n2055 VPWR.t1857 983.14
R7914 VPWR.n2054 VPWR.t0 983.14
R7915 VPWR.n2045 VPWR.t855 983.14
R7916 VPWR.n2044 VPWR.t437 983.14
R7917 VPWR.n2035 VPWR.t1113 983.14
R7918 VPWR.n2034 VPWR.t92 983.14
R7919 VPWR.n2025 VPWR.t1279 983.14
R7920 VPWR.n2024 VPWR.t889 983.14
R7921 VPWR.n2015 VPWR.t183 983.14
R7922 VPWR.t1908 VPWR.n774 983.14
R7923 VPWR.t257 VPWR.n778 983.14
R7924 VPWR.t783 VPWR.n782 983.14
R7925 VPWR.t1037 VPWR.n786 983.14
R7926 VPWR.t1318 VPWR.n790 983.14
R7927 VPWR.t555 VPWR.n794 983.14
R7928 VPWR.t489 VPWR.n798 983.14
R7929 VPWR.t845 VPWR.n802 983.14
R7930 VPWR.t517 VPWR.n806 983.14
R7931 VPWR.t585 VPWR.n810 983.14
R7932 VPWR.t704 VPWR.n814 983.14
R7933 VPWR.t1153 VPWR.n818 983.14
R7934 VPWR.t967 VPWR.n822 983.14
R7935 VPWR.t1890 VPWR.n826 983.14
R7936 VPWR.t199 VPWR.n830 983.14
R7937 VPWR.t481 VPWR.n1917 983.14
R7938 VPWR.n1918 VPWR.t511 983.14
R7939 VPWR.t815 VPWR.n1927 983.14
R7940 VPWR.n1928 VPWR.t1330 983.14
R7941 VPWR.t1202 VPWR.n1937 983.14
R7942 VPWR.n1938 VPWR.t59 983.14
R7943 VPWR.t1863 VPWR.n1947 983.14
R7944 VPWR.n1948 VPWR.t597 983.14
R7945 VPWR.t1220 VPWR.n1957 983.14
R7946 VPWR.n1958 VPWR.t338 983.14
R7947 VPWR.t1839 VPWR.n1967 983.14
R7948 VPWR.n1968 VPWR.t921 983.14
R7949 VPWR.t1291 VPWR.n1977 983.14
R7950 VPWR.n1978 VPWR.t24 983.14
R7951 VPWR.t867 VPWR.n1987 983.14
R7952 VPWR.n926 VPWR.t1906 983.14
R7953 VPWR.n925 VPWR.t255 983.14
R7954 VPWR.n921 VPWR.t785 983.14
R7955 VPWR.n917 VPWR.t1035 983.14
R7956 VPWR.n913 VPWR.t1316 983.14
R7957 VPWR.n909 VPWR.t553 983.14
R7958 VPWR.n905 VPWR.t487 983.14
R7959 VPWR.n901 VPWR.t841 983.14
R7960 VPWR.n897 VPWR.t515 983.14
R7961 VPWR.n893 VPWR.t583 983.14
R7962 VPWR.n889 VPWR.t702 983.14
R7963 VPWR.n885 VPWR.t1151 983.14
R7964 VPWR.n881 VPWR.t963 983.14
R7965 VPWR.n877 VPWR.t1888 983.14
R7966 VPWR.n873 VPWR.t197 983.14
R7967 VPWR.t483 VPWR.n390 983.14
R7968 VPWR.t513 VPWR.n394 983.14
R7969 VPWR.t813 VPWR.n398 983.14
R7970 VPWR.t1334 VPWR.n402 983.14
R7971 VPWR.t1204 VPWR.n406 983.14
R7972 VPWR.t61 VPWR.n410 983.14
R7973 VPWR.t1865 VPWR.n414 983.14
R7974 VPWR.t599 VPWR.n418 983.14
R7975 VPWR.t1222 VPWR.n422 983.14
R7976 VPWR.t340 VPWR.n426 983.14
R7977 VPWR.t1841 VPWR.n430 983.14
R7978 VPWR.t923 VPWR.n434 983.14
R7979 VPWR.t1293 VPWR.n438 983.14
R7980 VPWR.t8 VPWR.n442 983.14
R7981 VPWR.t871 VPWR.n446 983.14
R7982 VPWR.n1889 VPWR.t909 983.14
R7983 VPWR.n1888 VPWR.t1208 983.14
R7984 VPWR.n1879 VPWR.t797 983.14
R7985 VPWR.n1878 VPWR.t683 983.14
R7986 VPWR.n1869 VPWR.t658 983.14
R7987 VPWR.n1868 VPWR.t1752 983.14
R7988 VPWR.n1859 VPWR.t1736 983.14
R7989 VPWR.n1858 VPWR.t71 983.14
R7990 VPWR.n1849 VPWR.t1894 983.14
R7991 VPWR.n1848 VPWR.t359 983.14
R7992 VPWR.n1839 VPWR.t525 983.14
R7993 VPWR.n1838 VPWR.t1794 983.14
R7994 VPWR.n1829 VPWR.t1246 983.14
R7995 VPWR.n1828 VPWR.t31 983.14
R7996 VPWR.n1819 VPWR.t1002 983.14
R7997 VPWR.n2477 VPWR.t899 983.14
R7998 VPWR.n2476 VPWR.t1214 983.14
R7999 VPWR.n2467 VPWR.t793 983.14
R8000 VPWR.n2466 VPWR.t632 983.14
R8001 VPWR.n2457 VPWR.t401 983.14
R8002 VPWR.n2456 VPWR.t1758 983.14
R8003 VPWR.n2447 VPWR.t1742 983.14
R8004 VPWR.n2446 VPWR.t569 983.14
R8005 VPWR.n2437 VPWR.t1900 983.14
R8006 VPWR.n2436 VPWR.t363 983.14
R8007 VPWR.n2427 VPWR.t531 983.14
R8008 VPWR.n2426 VPWR.t1798 983.14
R8009 VPWR.n2417 VPWR.t1250 983.14
R8010 VPWR.n2416 VPWR.t1784 983.14
R8011 VPWR.n2407 VPWR.t1008 983.14
R8012 VPWR.t612 VPWR.n966 983.14
R8013 VPWR.t265 VPWR.n970 983.14
R8014 VPWR.t775 VPWR.n974 983.14
R8015 VPWR.t147 VPWR.n978 983.14
R8016 VPWR.t1184 VPWR.n982 983.14
R8017 VPWR.t563 VPWR.n986 983.14
R8018 VPWR.t497 VPWR.n990 983.14
R8019 VPWR.t284 VPWR.n994 983.14
R8020 VPWR.t106 VPWR.n998 983.14
R8021 VPWR.t589 VPWR.n1002 983.14
R8022 VPWR.t712 VPWR.n1006 983.14
R8023 VPWR.t1143 VPWR.n1010 983.14
R8024 VPWR.t535 VPWR.n1014 983.14
R8025 VPWR.t35 VPWR.n1018 983.14
R8026 VPWR.t209 VPWR.n1022 983.14
R8027 VPWR.n350 VPWR.t1022 983.14
R8028 VPWR.n349 VPWR.t1230 983.14
R8029 VPWR.n345 VPWR.t801 983.14
R8030 VPWR.n341 VPWR.t681 983.14
R8031 VPWR.n337 VPWR.t654 983.14
R8032 VPWR.n333 VPWR.t1818 983.14
R8033 VPWR.n329 VPWR.t1732 983.14
R8034 VPWR.n325 VPWR.t69 983.14
R8035 VPWR.n321 VPWR.t728 983.14
R8036 VPWR.n317 VPWR.t357 983.14
R8037 VPWR.n313 VPWR.t521 983.14
R8038 VPWR.n309 VPWR.t98 983.14
R8039 VPWR.n305 VPWR.t1244 983.14
R8040 VPWR.n301 VPWR.t18 983.14
R8041 VPWR.n297 VPWR.t879 983.14
R8042 VPWR.t1609 VPWR.n1468 983.14
R8043 VPWR.t1711 VPWR.n1475 983.14
R8044 VPWR.t1482 VPWR.n1481 983.14
R8045 VPWR.t1584 VPWR.n1492 983.14
R8046 VPWR.n1493 VPWR.t1606 983.14
R8047 VPWR.t1357 VPWR.n1506 983.14
R8048 VPWR.n1507 VPWR.t1479 983.14
R8049 VPWR.t1620 VPWR.n1520 983.14
R8050 VPWR.n1521 VPWR.t1636 983.14
R8051 VPWR.n1536 VPWR.t1379 983.14
R8052 VPWR.n1535 VPWR.t1509 983.14
R8053 VPWR.n1761 VPWR.t1550 983.14
R8054 VPWR.n1760 VPWR.t1373 983.14
R8055 VPWR.n1749 VPWR.t1423 983.14
R8056 VPWR.t1531 VPWR.n1791 983.14
R8057 VPWR.t1537 VPWR.n2506 983.14
R8058 VPWR.n2507 VPWR.t1649 983.14
R8059 VPWR.t1414 VPWR.n2518 983.14
R8060 VPWR.n2519 VPWR.t1525 983.14
R8061 VPWR.t1534 VPWR.n2530 983.14
R8062 VPWR.n2531 VPWR.t1690 983.14
R8063 VPWR.t1411 VPWR.n2542 983.14
R8064 VPWR.n2543 VPWR.t1571 983.14
R8065 VPWR.t1587 VPWR.n2554 983.14
R8066 VPWR.n2555 VPWR.t1717 983.14
R8067 VPWR.t1461 VPWR.n2566 983.14
R8068 VPWR.n2567 VPWR.t1491 983.14
R8069 VPWR.t1341 VPWR.n2578 983.14
R8070 VPWR.n2579 VPWR.t1360 983.14
R8071 VPWR.t1485 VPWR.n2590 983.14
R8072 VPWR.n1594 VPWR.t1420 983.14
R8073 VPWR.n1593 VPWR.t1522 983.14
R8074 VPWR.t1687 VPWR.n1182 983.14
R8075 VPWR.t1405 VPWR.n1185 983.14
R8076 VPWR.n1220 VPWR.t1417 983.14
R8077 VPWR.n1219 VPWR.t1576 983.14
R8078 VPWR.n1216 VPWR.t1684 983.14
R8079 VPWR.n1213 VPWR.t1445 983.14
R8080 VPWR.n1205 VPWR.t1471 983.14
R8081 VPWR.n1202 VPWR.t1598 983.14
R8082 VPWR.n1199 VPWR.t1344 983.14
R8083 VPWR.n1191 VPWR.t1365 983.14
R8084 VPWR.n1188 VPWR.t1603 983.14
R8085 VPWR.n1740 VPWR.t1631 983.14
R8086 VPWR.n1739 VPWR.t1351 983.14
R8087 VPWR.n1308 VPWR.t331 877.144
R8088 VPWR.n2723 VPWR.t249 877.144
R8089 VPWR.n2843 VPWR.n2822 857.648
R8090 VPWR.n1122 VPWR.t1653 738.074
R8091 VPWR.n99 VPWR.t1393 738.074
R8092 VPWR.n290 VPWR.t1062 738.074
R8093 VPWR.n68 VPWR.t1462 738.074
R8094 VPWR.n346 VPWR.t1023 738.074
R8095 VPWR.n98 VPWR.t1538 738.074
R8096 VPWR.n963 VPWR.t1048 738.074
R8097 VPWR.n356 VPWR.t1056 738.074
R8098 VPWR.n357 VPWR.t900 738.074
R8099 VPWR.n318 VPWR.t70 738.074
R8100 VPWR.n75 VPWR.t1572 738.074
R8101 VPWR.n971 VPWR.t266 738.074
R8102 VPWR.n369 VPWR.t1743 738.074
R8103 VPWR.n322 VPWR.t1733 738.074
R8104 VPWR.n80 VPWR.t1412 738.074
R8105 VPWR.n932 VPWR.t1060 738.074
R8106 VPWR.n933 VPWR.t910 738.074
R8107 VPWR.n936 VPWR.t1209 738.074
R8108 VPWR.n387 VPWR.t1066 738.074
R8109 VPWR.n391 VPWR.t484 738.074
R8110 VPWR.n395 VPWR.t514 738.074
R8111 VPWR.n365 VPWR.t402 738.074
R8112 VPWR.n330 VPWR.t655 738.074
R8113 VPWR.n86 VPWR.t1535 738.074
R8114 VPWR.n937 VPWR.t798 738.074
R8115 VPWR.n403 VPWR.t1335 738.074
R8116 VPWR.n364 VPWR.t633 738.074
R8117 VPWR.n334 VPWR.t682 738.074
R8118 VPWR.n87 VPWR.t1526 738.074
R8119 VPWR.n481 VPWR.t1075 738.074
R8120 VPWR.n480 VPWR.t958 738.074
R8121 VPWR.n477 VPWR.t1130 738.074
R8122 VPWR.n476 VPWR.t828 738.074
R8123 VPWR.n472 VPWR.t1122 738.074
R8124 VPWR.n469 VPWR.t1177 738.074
R8125 VPWR.n468 VPWR.t1257 738.074
R8126 VPWR.n465 VPWR.t737 738.074
R8127 VPWR.n464 VPWR.t580 738.074
R8128 VPWR.n461 VPWR.t432 738.074
R8129 VPWR.n460 VPWR.t1915 738.074
R8130 VPWR.n457 VPWR.t1781 738.074
R8131 VPWR.n456 VPWR.t546 738.074
R8132 VPWR.n453 VPWR.t884 738.074
R8133 VPWR.n452 VPWR.t182 738.074
R8134 VPWR.n473 VPWR.t154 738.074
R8135 VPWR.n482 VPWR.t1064 738.074
R8136 VPWR.n538 VPWR.t1021 738.074
R8137 VPWR.n534 VPWR.t1229 738.074
R8138 VPWR.n530 VPWR.t804 738.074
R8139 VPWR.n522 VPWR.t113 738.074
R8140 VPWR.n518 VPWR.t1817 738.074
R8141 VPWR.n514 VPWR.t1731 738.074
R8142 VPWR.n510 VPWR.t66 738.074
R8143 VPWR.n506 VPWR.t727 738.074
R8144 VPWR.n502 VPWR.t356 738.074
R8145 VPWR.n498 VPWR.t1829 738.074
R8146 VPWR.n494 VPWR.t97 738.074
R8147 VPWR.n490 VPWR.t1241 738.074
R8148 VPWR.n486 VPWR.t17 738.074
R8149 VPWR.n483 VPWR.t878 738.074
R8150 VPWR.n526 VPWR.t680 738.074
R8151 VPWR.n548 VPWR.t1050 738.074
R8152 VPWR.n549 VPWR.t1911 738.074
R8153 VPWR.n552 VPWR.t260 738.074
R8154 VPWR.n553 VPWR.t782 738.074
R8155 VPWR.n557 VPWR.t1321 738.074
R8156 VPWR.n560 VPWR.t558 738.074
R8157 VPWR.n561 VPWR.t492 738.074
R8158 VPWR.n564 VPWR.t850 738.074
R8159 VPWR.n565 VPWR.t520 738.074
R8160 VPWR.n568 VPWR.t588 738.074
R8161 VPWR.n569 VPWR.t707 738.074
R8162 VPWR.n572 VPWR.t1142 738.074
R8163 VPWR.n573 VPWR.t972 738.074
R8164 VPWR.n576 VPWR.t478 738.074
R8165 VPWR.n577 VPWR.t204 738.074
R8166 VPWR.n556 VPWR.t1042 738.074
R8167 VPWR.n579 VPWR.t1058 738.074
R8168 VPWR.n583 VPWR.t898 738.074
R8169 VPWR.n587 VPWR.t1213 738.074
R8170 VPWR.n591 VPWR.t796 738.074
R8171 VPWR.n599 VPWR.t400 738.074
R8172 VPWR.n603 VPWR.t1757 738.074
R8173 VPWR.n607 VPWR.t1741 738.074
R8174 VPWR.n611 VPWR.t74 738.074
R8175 VPWR.n615 VPWR.t1899 738.074
R8176 VPWR.n619 VPWR.t362 738.074
R8177 VPWR.n623 VPWR.t530 738.074
R8178 VPWR.n627 VPWR.t1797 738.074
R8179 VPWR.n631 VPWR.t1249 738.074
R8180 VPWR.n635 VPWR.t34 738.074
R8181 VPWR.n578 VPWR.t1005 738.074
R8182 VPWR.n595 VPWR.t686 738.074
R8183 VPWR.n673 VPWR.t1070 738.074
R8184 VPWR.n672 VPWR.t480 738.074
R8185 VPWR.n669 VPWR.t510 738.074
R8186 VPWR.n668 VPWR.t818 738.074
R8187 VPWR.n664 VPWR.t140 738.074
R8188 VPWR.n661 VPWR.t58 738.074
R8189 VPWR.n660 VPWR.t1862 738.074
R8190 VPWR.n657 VPWR.t596 738.074
R8191 VPWR.n656 VPWR.t1219 738.074
R8192 VPWR.n653 VPWR.t337 738.074
R8193 VPWR.n652 VPWR.t1838 738.074
R8194 VPWR.n649 VPWR.t920 738.074
R8195 VPWR.n648 VPWR.t1290 738.074
R8196 VPWR.n645 VPWR.t23 738.074
R8197 VPWR.n644 VPWR.t166 738.074
R8198 VPWR.n665 VPWR.t380 738.074
R8199 VPWR.n674 VPWR.t1077 738.074
R8200 VPWR.n730 VPWR.t621 738.074
R8201 VPWR.n726 VPWR.t768 738.074
R8202 VPWR.n722 VPWR.t830 738.074
R8203 VPWR.n714 VPWR.t1191 738.074
R8204 VPWR.n710 VPWR.t1175 738.074
R8205 VPWR.n706 VPWR.t1255 738.074
R8206 VPWR.n702 VPWR.t735 738.074
R8207 VPWR.n698 VPWR.t578 738.074
R8208 VPWR.n694 VPWR.t430 738.074
R8209 VPWR.n690 VPWR.t1913 738.074
R8210 VPWR.n686 VPWR.t1779 738.074
R8211 VPWR.n682 VPWR.t544 738.074
R8212 VPWR.n678 VPWR.t882 738.074
R8213 VPWR.n675 VPWR.t180 738.074
R8214 VPWR.n718 VPWR.t152 738.074
R8215 VPWR.n740 VPWR.t1073 738.074
R8216 VPWR.n741 VPWR.t1725 738.074
R8217 VPWR.n744 VPWR.t1136 738.074
R8218 VPWR.n745 VPWR.t824 738.074
R8219 VPWR.n749 VPWR.t1128 738.074
R8220 VPWR.n752 VPWR.t1164 738.074
R8221 VPWR.n753 VPWR.t1858 738.074
R8222 VPWR.n756 VPWR.t1 738.074
R8223 VPWR.n757 VPWR.t856 738.074
R8224 VPWR.n760 VPWR.t438 738.074
R8225 VPWR.n761 VPWR.t1114 738.074
R8226 VPWR.n764 VPWR.t93 738.074
R8227 VPWR.n765 VPWR.t1280 738.074
R8228 VPWR.n768 VPWR.t890 738.074
R8229 VPWR.n769 VPWR.t184 738.074
R8230 VPWR.n748 VPWR.t370 738.074
R8231 VPWR.n771 VPWR.t1052 738.074
R8232 VPWR.n775 VPWR.t1909 738.074
R8233 VPWR.n779 VPWR.t258 738.074
R8234 VPWR.n783 VPWR.t784 738.074
R8235 VPWR.n791 VPWR.t1319 738.074
R8236 VPWR.n795 VPWR.t556 738.074
R8237 VPWR.n799 VPWR.t490 738.074
R8238 VPWR.n803 VPWR.t846 738.074
R8239 VPWR.n807 VPWR.t518 738.074
R8240 VPWR.n811 VPWR.t586 738.074
R8241 VPWR.n815 VPWR.t705 738.074
R8242 VPWR.n819 VPWR.t1154 738.074
R8243 VPWR.n823 VPWR.t968 738.074
R8244 VPWR.n827 VPWR.t1891 738.074
R8245 VPWR.n770 VPWR.t200 738.074
R8246 VPWR.n787 VPWR.t1038 738.074
R8247 VPWR.n865 VPWR.t1068 738.074
R8248 VPWR.n864 VPWR.t482 738.074
R8249 VPWR.n861 VPWR.t512 738.074
R8250 VPWR.n860 VPWR.t816 738.074
R8251 VPWR.n856 VPWR.t1203 738.074
R8252 VPWR.n853 VPWR.t60 738.074
R8253 VPWR.n852 VPWR.t1864 738.074
R8254 VPWR.n849 VPWR.t598 738.074
R8255 VPWR.n848 VPWR.t1221 738.074
R8256 VPWR.n845 VPWR.t339 738.074
R8257 VPWR.n844 VPWR.t1840 738.074
R8258 VPWR.n841 VPWR.t922 738.074
R8259 VPWR.n840 VPWR.t1292 738.074
R8260 VPWR.n837 VPWR.t25 738.074
R8261 VPWR.n836 VPWR.t868 738.074
R8262 VPWR.n857 VPWR.t1331 738.074
R8263 VPWR.n866 VPWR.t1054 738.074
R8264 VPWR.n922 VPWR.t1907 738.074
R8265 VPWR.n918 VPWR.t256 738.074
R8266 VPWR.n914 VPWR.t786 738.074
R8267 VPWR.n906 VPWR.t1317 738.074
R8268 VPWR.n902 VPWR.t554 738.074
R8269 VPWR.n898 VPWR.t488 738.074
R8270 VPWR.n894 VPWR.t842 738.074
R8271 VPWR.n890 VPWR.t516 738.074
R8272 VPWR.n886 VPWR.t584 738.074
R8273 VPWR.n882 VPWR.t703 738.074
R8274 VPWR.n878 VPWR.t1152 738.074
R8275 VPWR.n874 VPWR.t964 738.074
R8276 VPWR.n870 VPWR.t1889 738.074
R8277 VPWR.n867 VPWR.t198 738.074
R8278 VPWR.n910 VPWR.t1036 738.074
R8279 VPWR.n940 VPWR.t684 738.074
R8280 VPWR.n979 VPWR.t148 738.074
R8281 VPWR.n1179 VPWR.t1406 738.074
R8282 VPWR.n399 VPWR.t814 738.074
R8283 VPWR.n361 VPWR.t794 738.074
R8284 VPWR.n338 VPWR.t802 738.074
R8285 VPWR.n92 VPWR.t1415 738.074
R8286 VPWR.n975 VPWR.t776 738.074
R8287 VPWR.n1183 VPWR.t1688 738.074
R8288 VPWR.n941 VPWR.t659 738.074
R8289 VPWR.n983 VPWR.t1185 738.074
R8290 VPWR.n1217 VPWR.t1418 738.074
R8291 VPWR.n407 VPWR.t1205 738.074
R8292 VPWR.n415 VPWR.t1866 738.074
R8293 VPWR.n419 VPWR.t600 738.074
R8294 VPWR.n423 VPWR.t1223 738.074
R8295 VPWR.n427 VPWR.t341 738.074
R8296 VPWR.n431 VPWR.t1842 738.074
R8297 VPWR.n435 VPWR.t924 738.074
R8298 VPWR.n439 VPWR.t1294 738.074
R8299 VPWR.n443 VPWR.t9 738.074
R8300 VPWR.n386 VPWR.t872 738.074
R8301 VPWR.n411 VPWR.t62 738.074
R8302 VPWR.n368 VPWR.t1759 738.074
R8303 VPWR.n326 VPWR.t1819 738.074
R8304 VPWR.n81 VPWR.t1691 738.074
R8305 VPWR.n987 VPWR.t564 738.074
R8306 VPWR.n1214 VPWR.t1577 738.074
R8307 VPWR.n944 VPWR.t1753 738.074
R8308 VPWR.n948 VPWR.t72 738.074
R8309 VPWR.n949 VPWR.t1895 738.074
R8310 VPWR.n952 VPWR.t360 738.074
R8311 VPWR.n953 VPWR.t526 738.074
R8312 VPWR.n956 VPWR.t1795 738.074
R8313 VPWR.n957 VPWR.t1247 738.074
R8314 VPWR.n960 VPWR.t32 738.074
R8315 VPWR.n961 VPWR.t1003 738.074
R8316 VPWR.n945 VPWR.t1737 738.074
R8317 VPWR.n991 VPWR.t498 738.074
R8318 VPWR.n1206 VPWR.t1685 738.074
R8319 VPWR.n360 VPWR.t1215 738.074
R8320 VPWR.n342 VPWR.t1231 738.074
R8321 VPWR.n93 VPWR.t1650 738.074
R8322 VPWR.n1180 VPWR.t1523 738.074
R8323 VPWR.n995 VPWR.t285 738.074
R8324 VPWR.n1203 VPWR.t1446 738.074
R8325 VPWR.n372 VPWR.t570 738.074
R8326 VPWR.n376 VPWR.t364 738.074
R8327 VPWR.n377 VPWR.t532 738.074
R8328 VPWR.n380 VPWR.t1799 738.074
R8329 VPWR.n381 VPWR.t1251 738.074
R8330 VPWR.n384 VPWR.t1785 738.074
R8331 VPWR.n385 VPWR.t1009 738.074
R8332 VPWR.n373 VPWR.t1901 738.074
R8333 VPWR.n314 VPWR.t729 738.074
R8334 VPWR.n74 VPWR.t1588 738.074
R8335 VPWR.n1200 VPWR.t1472 738.074
R8336 VPWR.n999 VPWR.t107 738.074
R8337 VPWR.n1003 VPWR.t590 738.074
R8338 VPWR.n1007 VPWR.t713 738.074
R8339 VPWR.n1011 VPWR.t1144 738.074
R8340 VPWR.n1015 VPWR.t536 738.074
R8341 VPWR.n1019 VPWR.t36 738.074
R8342 VPWR.n962 VPWR.t210 738.074
R8343 VPWR.n967 VPWR.t613 738.074
R8344 VPWR.n1123 VPWR.t1421 738.074
R8345 VPWR.n310 VPWR.t358 738.074
R8346 VPWR.n69 VPWR.t1718 738.074
R8347 VPWR.n1192 VPWR.t1599 738.074
R8348 VPWR.n1189 VPWR.t1345 738.074
R8349 VPWR.n306 VPWR.t522 738.074
R8350 VPWR.n302 VPWR.t99 738.074
R8351 VPWR.n294 VPWR.t19 738.074
R8352 VPWR.n291 VPWR.t880 738.074
R8353 VPWR.n298 VPWR.t1245 738.074
R8354 VPWR.n1058 VPWR.t1604 738.074
R8355 VPWR.n1186 VPWR.t1366 738.074
R8356 VPWR.n63 VPWR.t1492 738.074
R8357 VPWR.n62 VPWR.t1342 738.074
R8358 VPWR.n57 VPWR.t1361 738.074
R8359 VPWR.n56 VPWR.t1486 738.074
R8360 VPWR.n1059 VPWR.t1632 738.074
R8361 VPWR.n1061 VPWR.t1352 738.074
R8362 VPWR.n2856 VPWR.n2821 702.354
R8363 VPWR.n2856 VPWR.n2822 702.354
R8364 VPWR.n2854 VPWR.n2853 702.354
R8365 VPWR.n2854 VPWR.n2821 702.354
R8366 VPWR.n2837 VPWR.n2828 702.354
R8367 VPWR.n2850 VPWR.n2849 702.354
R8368 VPWR.n2835 VPWR.n2828 702.354
R8369 VPWR.n2815 VPWR.t194 651.634
R8370 VPWR.n2831 VPWR.t1071 651.505
R8371 VPWR.n2825 VPWR.t669 651.505
R8372 VPWR.n2862 VPWR.t694 651.431
R8373 VPWR.n1061 VPWR.t1475 646.071
R8374 VPWR.n1122 VPWR.t1371 646.071
R8375 VPWR.n1059 VPWR.t1624 646.071
R8376 VPWR.n56 VPWR.t1591 646.071
R8377 VPWR.n62 VPWR.t1715 646.071
R8378 VPWR.n99 VPWR.t1500 646.071
R8379 VPWR.n1053 VPWR.t542 646.071
R8380 VPWR.n1231 VPWR.t896 646.071
R8381 VPWR.n298 VPWR.t1789 646.071
R8382 VPWR.n290 VPWR.t904 646.071
R8383 VPWR.n306 VPWR.t1803 646.071
R8384 VPWR.n68 VPWR.t1454 646.071
R8385 VPWR.n1153 VPWR.t221 646.071
R8386 VPWR.n346 VPWR.t1211 646.071
R8387 VPWR.n98 VPWR.t1629 646.071
R8388 VPWR.n967 VPWR.t766 646.071
R8389 VPWR.n963 VPWR.t960 646.071
R8390 VPWR.n999 VPWR.t434 646.071
R8391 VPWR.n373 VPWR.t386 646.071
R8392 VPWR.n356 VPWR.t894 646.071
R8393 VPWR.n357 VPWR.t1140 646.071
R8394 VPWR.n372 VPWR.t1106 646.071
R8395 VPWR.n318 VPWR.t1897 646.071
R8396 VPWR.n75 VPWR.t1559 646.071
R8397 VPWR.n971 VPWR.t812 646.071
R8398 VPWR.n369 VPWR.t289 646.071
R8399 VPWR.n322 VPWR.t848 646.071
R8400 VPWR.n80 VPWR.t1431 646.071
R8401 VPWR.n945 VPWR.t852 646.071
R8402 VPWR.n932 VPWR.t906 646.071
R8403 VPWR.n933 VPWR.t1217 646.071
R8404 VPWR.n936 VPWR.t774 646.071
R8405 VPWR.n944 VPWR.t1745 646.071
R8406 VPWR.n411 VPWR.t1872 646.071
R8407 VPWR.n387 VPWR.t1019 646.071
R8408 VPWR.n391 VPWR.t146 646.071
R8409 VPWR.n395 VPWR.t788 646.071
R8410 VPWR.n407 VPWR.t1815 646.071
R8411 VPWR.n365 VPWR.t696 646.071
R8412 VPWR.n330 VPWR.t1755 646.071
R8413 VPWR.n86 VPWR.t1672 646.071
R8414 VPWR.n937 VPWR.t1040 646.071
R8415 VPWR.n403 VPWR.t723 646.071
R8416 VPWR.n364 VPWR.t408 646.071
R8417 VPWR.n334 VPWR.t661 646.071
R8418 VPWR.n87 VPWR.t1517 646.071
R8419 VPWR.n473 VPWR.t1126 646.071
R8420 VPWR.n481 VPWR.t1727 646.071
R8421 VPWR.n480 VPWR.t1134 646.071
R8422 VPWR.n477 VPWR.t806 646.071
R8423 VPWR.n476 VPWR.t1337 646.071
R8424 VPWR.n472 VPWR.t1162 646.071
R8425 VPWR.n469 VPWR.t1261 646.071
R8426 VPWR.n468 VPWR.t604 646.071
R8427 VPWR.n465 VPWR.t854 646.071
R8428 VPWR.n464 VPWR.t440 646.071
R8429 VPWR.n461 VPWR.t1919 646.071
R8430 VPWR.n460 VPWR.t95 646.071
R8431 VPWR.n457 VPWR.t1239 646.071
R8432 VPWR.n456 VPWR.t892 646.071
R8433 VPWR.n453 VPWR.t874 646.071
R8434 VPWR.n452 VPWR.t1489 646.071
R8435 VPWR.n526 VPWR.t657 646.071
R8436 VPWR.n482 VPWR.t902 646.071
R8437 VPWR.n538 VPWR.t1207 646.071
R8438 VPWR.n534 VPWR.t780 646.071
R8439 VPWR.n530 VPWR.t1032 646.071
R8440 VPWR.n522 VPWR.t1751 646.071
R8441 VPWR.n518 VPWR.t1735 646.071
R8442 VPWR.n514 VPWR.t844 646.071
R8443 VPWR.n510 VPWR.t731 646.071
R8444 VPWR.n506 VPWR.t366 646.071
R8445 VPWR.n502 VPWR.t524 646.071
R8446 VPWR.n498 VPWR.t1801 646.071
R8447 VPWR.n494 VPWR.t966 646.071
R8448 VPWR.n490 VPWR.t1787 646.071
R8449 VPWR.n486 VPWR.t1015 646.071
R8450 VPWR.n483 VPWR.t1707 646.071
R8451 VPWR.n556 VPWR.t1187 646.071
R8452 VPWR.n548 VPWR.t619 646.071
R8453 VPWR.n549 VPWR.t268 646.071
R8454 VPWR.n552 VPWR.t820 646.071
R8455 VPWR.n553 VPWR.t376 646.071
R8456 VPWR.n557 VPWR.t1171 646.071
R8457 VPWR.n560 VPWR.t500 646.071
R8458 VPWR.n561 VPWR.t7 646.071
R8459 VPWR.n564 VPWR.t109 646.071
R8460 VPWR.n565 VPWR.t428 646.071
R8461 VPWR.n568 VPWR.t715 646.071
R8462 VPWR.n569 VPWR.t1150 646.071
R8463 VPWR.n572 VPWR.t1286 646.071
R8464 VPWR.n573 VPWR.t42 646.071
R8465 VPWR.n576 VPWR.t162 646.071
R8466 VPWR.n577 VPWR.t1556 646.071
R8467 VPWR.n595 VPWR.t406 646.071
R8468 VPWR.n579 VPWR.t908 646.071
R8469 VPWR.n583 VPWR.t1138 646.071
R8470 VPWR.n587 VPWR.t772 646.071
R8471 VPWR.n591 VPWR.t1044 646.071
R8472 VPWR.n599 VPWR.t1763 646.071
R8473 VPWR.n603 VPWR.t1747 646.071
R8474 VPWR.n607 VPWR.t287 646.071
R8475 VPWR.n611 VPWR.t1905 646.071
R8476 VPWR.n615 VPWR.t384 646.071
R8477 VPWR.n619 VPWR.t217 646.071
R8478 VPWR.n623 VPWR.t1156 646.071
R8479 VPWR.n627 VPWR.t538 646.071
R8480 VPWR.n631 VPWR.t1793 646.071
R8481 VPWR.n635 VPWR.t206 646.071
R8482 VPWR.n578 VPWR.t1664 646.071
R8483 VPWR.n665 VPWR.t719 646.071
R8484 VPWR.n673 VPWR.t1296 646.071
R8485 VPWR.n672 VPWR.t142 646.071
R8486 VPWR.n669 VPWR.t792 646.071
R8487 VPWR.n668 VPWR.t688 646.071
R8488 VPWR.n664 VPWR.t64 646.071
R8489 VPWR.n661 VPWR.t1868 646.071
R8490 VPWR.n660 VPWR.t572 646.071
R8491 VPWR.n657 VPWR.t1225 646.071
R8492 VPWR.n656 VPWR.t343 646.071
R8493 VPWR.n653 VPWR.t1844 646.071
R8494 VPWR.n652 VPWR.t1807 646.071
R8495 VPWR.n649 VPWR.t1253 646.071
R8496 VPWR.n648 VPWR.t11 646.071
R8497 VPWR.n645 VPWR.t1007 646.071
R8498 VPWR.n644 VPWR.t1390 646.071
R8499 VPWR.n718 VPWR.t1124 646.071
R8500 VPWR.n674 VPWR.t962 646.071
R8501 VPWR.n730 VPWR.t1132 646.071
R8502 VPWR.n726 VPWR.t810 646.071
R8503 VPWR.n722 VPWR.t1333 646.071
R8504 VPWR.n714 VPWR.t1179 646.071
R8505 VPWR.n710 VPWR.t1259 646.071
R8506 VPWR.n706 VPWR.t602 646.071
R8507 VPWR.n702 VPWR.t582 646.071
R8508 VPWR.n698 VPWR.t436 646.071
R8509 VPWR.n694 VPWR.t1917 646.071
R8510 VPWR.n690 VPWR.t91 646.071
R8511 VPWR.n686 VPWR.t1237 646.071
R8512 VPWR.n682 VPWR.t888 646.071
R8513 VPWR.n678 VPWR.t870 646.071
R8514 VPWR.n675 VPWR.t1497 646.071
R8515 VPWR.n748 VPWR.t138 646.071
R8516 VPWR.n740 VPWR.t1729 646.071
R8517 VPWR.n741 VPWR.t508 646.071
R8518 VPWR.n744 VPWR.t800 646.071
R8519 VPWR.n745 VPWR.t1339 646.071
R8520 VPWR.n749 VPWR.t1166 646.071
R8521 VPWR.n752 VPWR.t1860 646.071
R8522 VPWR.n753 VPWR.t68 646.071
R8523 VPWR.n756 VPWR.t858 646.071
R8524 VPWR.n757 VPWR.t335 646.071
R8525 VPWR.n760 VPWR.t1116 646.071
R8526 VPWR.n761 VPWR.t1079 646.071
R8527 VPWR.n764 VPWR.t1243 646.071
R8528 VPWR.n765 VPWR.t21 646.071
R8529 VPWR.n768 VPWR.t876 646.071
R8530 VPWR.n769 VPWR.t1457 646.071
R8531 VPWR.n787 VPWR.t1325 646.071
R8532 VPWR.n771 VPWR.t617 646.071
R8533 VPWR.n775 VPWR.t264 646.071
R8534 VPWR.n779 VPWR.t808 646.071
R8535 VPWR.n783 VPWR.t374 646.071
R8536 VPWR.n791 VPWR.t562 646.071
R8537 VPWR.n795 VPWR.t496 646.071
R8538 VPWR.n799 VPWR.t5 646.071
R8539 VPWR.n803 VPWR.t105 646.071
R8540 VPWR.n807 VPWR.t426 646.071
R8541 VPWR.n811 VPWR.t711 646.071
R8542 VPWR.n815 VPWR.t1148 646.071
R8543 VPWR.n819 VPWR.t1284 646.071
R8544 VPWR.n823 VPWR.t40 646.071
R8545 VPWR.n827 VPWR.t188 646.071
R8546 VPWR.n770 VPWR.t1562 646.071
R8547 VPWR.n857 VPWR.t721 646.071
R8548 VPWR.n865 VPWR.t1017 646.071
R8549 VPWR.n864 VPWR.t144 646.071
R8550 VPWR.n861 VPWR.t790 646.071
R8551 VPWR.n860 VPWR.t635 646.071
R8552 VPWR.n856 VPWR.t1813 646.071
R8553 VPWR.n853 VPWR.t1870 646.071
R8554 VPWR.n852 VPWR.t574 646.071
R8555 VPWR.n849 VPWR.t1227 646.071
R8556 VPWR.n848 VPWR.t345 646.071
R8557 VPWR.n845 VPWR.t1825 646.071
R8558 VPWR.n844 VPWR.t1809 646.071
R8559 VPWR.n841 VPWR.t943 646.071
R8560 VPWR.n840 VPWR.t13 646.071
R8561 VPWR.n837 VPWR.t1011 646.071
R8562 VPWR.n836 VPWR.t1385 646.071
R8563 VPWR.n910 VPWR.t1323 646.071
R8564 VPWR.n866 VPWR.t615 646.071
R8565 VPWR.n922 VPWR.t262 646.071
R8566 VPWR.n918 VPWR.t822 646.071
R8567 VPWR.n914 VPWR.t372 646.071
R8568 VPWR.n906 VPWR.t560 646.071
R8569 VPWR.n902 VPWR.t494 646.071
R8570 VPWR.n898 VPWR.t3 646.071
R8571 VPWR.n894 VPWR.t103 646.071
R8572 VPWR.n890 VPWR.t592 646.071
R8573 VPWR.n886 VPWR.t709 646.071
R8574 VPWR.n882 VPWR.t1146 646.071
R8575 VPWR.n878 VPWR.t1282 646.071
R8576 VPWR.n874 VPWR.t38 646.071
R8577 VPWR.n870 VPWR.t186 646.071
R8578 VPWR.n867 VPWR.t1569 646.071
R8579 VPWR.n940 VPWR.t404 646.071
R8580 VPWR.n979 VPWR.t1189 646.071
R8581 VPWR.n1227 VPWR.t506 646.071
R8582 VPWR.n1179 VPWR.t1401 646.071
R8583 VPWR.n399 VPWR.t637 646.071
R8584 VPWR.n361 VPWR.t1046 646.071
R8585 VPWR.n338 VPWR.t1034 646.071
R8586 VPWR.n92 VPWR.t1409 646.071
R8587 VPWR.n975 VPWR.t378 646.071
R8588 VPWR.n1485 VPWR.t150 646.071
R8589 VPWR.n1183 VPWR.t1680 646.071
R8590 VPWR.n941 VPWR.t1761 646.071
R8591 VPWR.n983 VPWR.t1173 646.071
R8592 VPWR.n1173 VPWR.t698 646.071
R8593 VPWR.n1217 VPWR.t1548 646.071
R8594 VPWR.n415 VPWR.t576 646.071
R8595 VPWR.n419 VPWR.t725 646.071
R8596 VPWR.n423 VPWR.t347 646.071
R8597 VPWR.n427 VPWR.t1827 646.071
R8598 VPWR.n431 VPWR.t1811 646.071
R8599 VPWR.n435 VPWR.t945 646.071
R8600 VPWR.n439 VPWR.t15 646.071
R8601 VPWR.n443 VPWR.t1013 646.071
R8602 VPWR.n386 VPWR.t1377 646.071
R8603 VPWR.n368 VPWR.t1749 646.071
R8604 VPWR.n326 VPWR.t1739 646.071
R8605 VPWR.n81 VPWR.t1396 646.071
R8606 VPWR.n987 VPWR.t442 646.071
R8607 VPWR.n1169 VPWR.t486 646.071
R8608 VPWR.n1214 VPWR.t1656 646.071
R8609 VPWR.n948 VPWR.t1903 646.071
R8610 VPWR.n949 VPWR.t382 646.071
R8611 VPWR.n952 VPWR.t534 646.071
R8612 VPWR.n953 VPWR.t1805 646.071
R8613 VPWR.n956 VPWR.t974 646.071
R8614 VPWR.n957 VPWR.t1791 646.071
R8615 VPWR.n960 VPWR.t202 646.071
R8616 VPWR.n961 VPWR.t1677 646.071
R8617 VPWR.n991 VPWR.t594 646.071
R8618 VPWR.n1163 VPWR.t733 646.071
R8619 VPWR.n1206 VPWR.t1696 646.071
R8620 VPWR.n360 VPWR.t770 646.071
R8621 VPWR.n342 VPWR.t778 646.071
R8622 VPWR.n93 VPWR.t1647 646.071
R8623 VPWR.n1479 VPWR.t826 646.071
R8624 VPWR.n1180 VPWR.t1520 646.071
R8625 VPWR.n995 VPWR.t111 646.071
R8626 VPWR.n1159 VPWR.t1108 646.071
R8627 VPWR.n1203 VPWR.t1441 646.071
R8628 VPWR.n376 VPWR.t219 646.071
R8629 VPWR.n377 VPWR.t1158 646.071
R8630 VPWR.n380 VPWR.t540 646.071
R8631 VPWR.n381 VPWR.t1025 646.071
R8632 VPWR.n384 VPWR.t208 646.071
R8633 VPWR.n385 VPWR.t1659 646.071
R8634 VPWR.n314 VPWR.t368 646.071
R8635 VPWR.n74 VPWR.t1669 646.071
R8636 VPWR.n1149 VPWR.t388 646.071
R8637 VPWR.n1200 VPWR.t1545 646.071
R8638 VPWR.n1003 VPWR.t717 646.071
R8639 VPWR.n1007 VPWR.t1783 646.071
R8640 VPWR.n1011 VPWR.t1288 646.071
R8641 VPWR.n1015 VPWR.t886 646.071
R8642 VPWR.n1019 VPWR.t164 646.071
R8643 VPWR.n962 VPWR.t1529 646.071
R8644 VPWR.n1472 VPWR.t1893 646.071
R8645 VPWR.n1123 VPWR.t1507 646.071
R8646 VPWR.n310 VPWR.t528 646.071
R8647 VPWR.n69 VPWR.t1436 646.071
R8648 VPWR.n1192 VPWR.t1704 646.071
R8649 VPWR.n1049 VPWR.t1160 646.071
R8650 VPWR.n1189 VPWR.t1723 646.071
R8651 VPWR.n302 VPWR.t970 646.071
R8652 VPWR.n294 VPWR.t196 646.071
R8653 VPWR.n291 VPWR.t1699 646.071
R8654 VPWR.n1058 VPWR.t1596 646.071
R8655 VPWR.n1748 VPWR.t1027 646.071
R8656 VPWR.n1036 VPWR.t212 646.071
R8657 VPWR.n1032 VPWR.t1640 646.071
R8658 VPWR.n1186 VPWR.t1467 646.071
R8659 VPWR.n63 VPWR.t1582 646.071
R8660 VPWR.n57 VPWR.t1355 646.071
R8661 VPWR.n1230 VPWR.t1449 642.13
R8662 VPWR.n1152 VPWR.t1380 642.13
R8663 VPWR.n1226 VPWR.t1585 642.13
R8664 VPWR.n1484 VPWR.t1483 642.13
R8665 VPWR.n1172 VPWR.t1607 642.13
R8666 VPWR.n1168 VPWR.t1358 642.13
R8667 VPWR.n1162 VPWR.t1480 642.13
R8668 VPWR.n1478 VPWR.t1712 642.13
R8669 VPWR.n1158 VPWR.t1621 642.13
R8670 VPWR.n1148 VPWR.t1637 642.13
R8671 VPWR.n1471 VPWR.t1610 642.13
R8672 VPWR.n1048 VPWR.t1510 642.13
R8673 VPWR.n1747 VPWR.t1374 642.13
R8674 VPWR.n1035 VPWR.t1424 642.13
R8675 VPWR.n1031 VPWR.t1532 642.13
R8676 VPWR.n1052 VPWR.t1551 642.13
R8677 VPWR.n2309 VPWR.t1726 629.652
R8678 VPWR.n2310 VPWR.t1133 629.652
R8679 VPWR.n2319 VPWR.t805 629.652
R8680 VPWR.n2320 VPWR.t1336 629.652
R8681 VPWR.n2329 VPWR.t1125 629.652
R8682 VPWR.n2330 VPWR.t1161 629.652
R8683 VPWR.n2339 VPWR.t1260 629.652
R8684 VPWR.n2340 VPWR.t603 629.652
R8685 VPWR.n2349 VPWR.t853 629.652
R8686 VPWR.n2350 VPWR.t439 629.652
R8687 VPWR.n2359 VPWR.t1918 629.652
R8688 VPWR.n2360 VPWR.t94 629.652
R8689 VPWR.n2369 VPWR.t1238 629.652
R8690 VPWR.n2370 VPWR.t891 629.652
R8691 VPWR.n2379 VPWR.t873 629.652
R8692 VPWR.n542 VPWR.t901 629.652
R8693 VPWR.t1206 VPWR.n541 629.652
R8694 VPWR.t779 VPWR.n537 629.652
R8695 VPWR.t1031 VPWR.n533 629.652
R8696 VPWR.t656 VPWR.n529 629.652
R8697 VPWR.t1750 VPWR.n525 629.652
R8698 VPWR.t1734 VPWR.n521 629.652
R8699 VPWR.t843 VPWR.n517 629.652
R8700 VPWR.t730 VPWR.n513 629.652
R8701 VPWR.t365 VPWR.n509 629.652
R8702 VPWR.t523 VPWR.n505 629.652
R8703 VPWR.t1800 VPWR.n501 629.652
R8704 VPWR.t965 VPWR.n497 629.652
R8705 VPWR.t1786 VPWR.n493 629.652
R8706 VPWR.t1014 VPWR.n489 629.652
R8707 VPWR.n2281 VPWR.t618 629.652
R8708 VPWR.t267 VPWR.n2280 629.652
R8709 VPWR.n2271 VPWR.t819 629.652
R8710 VPWR.t375 VPWR.n2270 629.652
R8711 VPWR.n2261 VPWR.t1186 629.652
R8712 VPWR.t1170 VPWR.n2260 629.652
R8713 VPWR.n2251 VPWR.t499 629.652
R8714 VPWR.t6 VPWR.n2250 629.652
R8715 VPWR.n2241 VPWR.t108 629.652
R8716 VPWR.t427 VPWR.n2240 629.652
R8717 VPWR.n2231 VPWR.t714 629.652
R8718 VPWR.t1149 VPWR.n2230 629.652
R8719 VPWR.n2221 VPWR.t1285 629.652
R8720 VPWR.t41 VPWR.n2220 629.652
R8721 VPWR.n2211 VPWR.t161 629.652
R8722 VPWR.n582 VPWR.t907 629.652
R8723 VPWR.n586 VPWR.t1137 629.652
R8724 VPWR.n590 VPWR.t771 629.652
R8725 VPWR.n594 VPWR.t1043 629.652
R8726 VPWR.n598 VPWR.t405 629.652
R8727 VPWR.n602 VPWR.t1762 629.652
R8728 VPWR.n606 VPWR.t1746 629.652
R8729 VPWR.n610 VPWR.t286 629.652
R8730 VPWR.n614 VPWR.t1904 629.652
R8731 VPWR.n618 VPWR.t383 629.652
R8732 VPWR.n622 VPWR.t216 629.652
R8733 VPWR.n626 VPWR.t1155 629.652
R8734 VPWR.n630 VPWR.t537 629.652
R8735 VPWR.n634 VPWR.t1792 629.652
R8736 VPWR.n638 VPWR.t205 629.652
R8737 VPWR.n2113 VPWR.t1295 629.652
R8738 VPWR.n2114 VPWR.t141 629.652
R8739 VPWR.n2123 VPWR.t791 629.652
R8740 VPWR.n2124 VPWR.t687 629.652
R8741 VPWR.n2133 VPWR.t718 629.652
R8742 VPWR.n2134 VPWR.t63 629.652
R8743 VPWR.n2143 VPWR.t1867 629.652
R8744 VPWR.n2144 VPWR.t571 629.652
R8745 VPWR.n2153 VPWR.t1224 629.652
R8746 VPWR.n2154 VPWR.t342 629.652
R8747 VPWR.n2163 VPWR.t1843 629.652
R8748 VPWR.n2164 VPWR.t1806 629.652
R8749 VPWR.n2173 VPWR.t1252 629.652
R8750 VPWR.n2174 VPWR.t10 629.652
R8751 VPWR.n2183 VPWR.t1006 629.652
R8752 VPWR.n734 VPWR.t961 629.652
R8753 VPWR.t1131 VPWR.n733 629.652
R8754 VPWR.t809 VPWR.n729 629.652
R8755 VPWR.t1332 VPWR.n725 629.652
R8756 VPWR.t1123 VPWR.n721 629.652
R8757 VPWR.t1178 VPWR.n717 629.652
R8758 VPWR.t1258 VPWR.n713 629.652
R8759 VPWR.t601 VPWR.n709 629.652
R8760 VPWR.t581 VPWR.n705 629.652
R8761 VPWR.t435 VPWR.n701 629.652
R8762 VPWR.t1916 VPWR.n697 629.652
R8763 VPWR.t90 VPWR.n693 629.652
R8764 VPWR.t1236 VPWR.n689 629.652
R8765 VPWR.t887 VPWR.n685 629.652
R8766 VPWR.t869 VPWR.n681 629.652
R8767 VPWR.n2085 VPWR.t1728 629.652
R8768 VPWR.t507 VPWR.n2084 629.652
R8769 VPWR.n2075 VPWR.t799 629.652
R8770 VPWR.t1338 VPWR.n2074 629.652
R8771 VPWR.n2065 VPWR.t137 629.652
R8772 VPWR.t1165 VPWR.n2064 629.652
R8773 VPWR.n2055 VPWR.t1859 629.652
R8774 VPWR.t67 VPWR.n2054 629.652
R8775 VPWR.n2045 VPWR.t857 629.652
R8776 VPWR.t334 VPWR.n2044 629.652
R8777 VPWR.n2035 VPWR.t1115 629.652
R8778 VPWR.t1078 VPWR.n2034 629.652
R8779 VPWR.n2025 VPWR.t1242 629.652
R8780 VPWR.t20 VPWR.n2024 629.652
R8781 VPWR.n2015 VPWR.t875 629.652
R8782 VPWR.n774 VPWR.t616 629.652
R8783 VPWR.n778 VPWR.t263 629.652
R8784 VPWR.n782 VPWR.t807 629.652
R8785 VPWR.n786 VPWR.t373 629.652
R8786 VPWR.n790 VPWR.t1324 629.652
R8787 VPWR.n794 VPWR.t561 629.652
R8788 VPWR.n798 VPWR.t495 629.652
R8789 VPWR.n802 VPWR.t4 629.652
R8790 VPWR.n806 VPWR.t104 629.652
R8791 VPWR.n810 VPWR.t425 629.652
R8792 VPWR.n814 VPWR.t710 629.652
R8793 VPWR.n818 VPWR.t1147 629.652
R8794 VPWR.n822 VPWR.t1283 629.652
R8795 VPWR.n826 VPWR.t39 629.652
R8796 VPWR.n830 VPWR.t187 629.652
R8797 VPWR.n1917 VPWR.t1016 629.652
R8798 VPWR.n1918 VPWR.t143 629.652
R8799 VPWR.n1927 VPWR.t789 629.652
R8800 VPWR.n1928 VPWR.t634 629.652
R8801 VPWR.n1937 VPWR.t720 629.652
R8802 VPWR.n1938 VPWR.t1812 629.652
R8803 VPWR.n1947 VPWR.t1869 629.652
R8804 VPWR.n1948 VPWR.t573 629.652
R8805 VPWR.n1957 VPWR.t1226 629.652
R8806 VPWR.n1958 VPWR.t344 629.652
R8807 VPWR.n1967 VPWR.t1824 629.652
R8808 VPWR.n1968 VPWR.t1808 629.652
R8809 VPWR.n1977 VPWR.t942 629.652
R8810 VPWR.n1978 VPWR.t12 629.652
R8811 VPWR.n1987 VPWR.t1010 629.652
R8812 VPWR.n926 VPWR.t614 629.652
R8813 VPWR.t261 VPWR.n925 629.652
R8814 VPWR.t821 VPWR.n921 629.652
R8815 VPWR.t371 VPWR.n917 629.652
R8816 VPWR.t1322 VPWR.n913 629.652
R8817 VPWR.t559 VPWR.n909 629.652
R8818 VPWR.t493 VPWR.n905 629.652
R8819 VPWR.t2 VPWR.n901 629.652
R8820 VPWR.t102 VPWR.n897 629.652
R8821 VPWR.t591 VPWR.n893 629.652
R8822 VPWR.t708 VPWR.n889 629.652
R8823 VPWR.t1145 VPWR.n885 629.652
R8824 VPWR.t1281 VPWR.n881 629.652
R8825 VPWR.t37 VPWR.n877 629.652
R8826 VPWR.t185 VPWR.n873 629.652
R8827 VPWR.n390 VPWR.t1018 629.652
R8828 VPWR.n394 VPWR.t145 629.652
R8829 VPWR.n398 VPWR.t787 629.652
R8830 VPWR.n402 VPWR.t636 629.652
R8831 VPWR.n406 VPWR.t722 629.652
R8832 VPWR.n410 VPWR.t1814 629.652
R8833 VPWR.n414 VPWR.t1871 629.652
R8834 VPWR.n418 VPWR.t575 629.652
R8835 VPWR.n422 VPWR.t724 629.652
R8836 VPWR.n426 VPWR.t346 629.652
R8837 VPWR.n430 VPWR.t1826 629.652
R8838 VPWR.n434 VPWR.t1810 629.652
R8839 VPWR.n438 VPWR.t944 629.652
R8840 VPWR.n442 VPWR.t14 629.652
R8841 VPWR.n446 VPWR.t1012 629.652
R8842 VPWR.n1889 VPWR.t905 629.652
R8843 VPWR.t1216 VPWR.n1888 629.652
R8844 VPWR.n1879 VPWR.t773 629.652
R8845 VPWR.t1039 VPWR.n1878 629.652
R8846 VPWR.n1869 VPWR.t403 629.652
R8847 VPWR.t1760 VPWR.n1868 629.652
R8848 VPWR.n1859 VPWR.t1744 629.652
R8849 VPWR.t851 VPWR.n1858 629.652
R8850 VPWR.n1849 VPWR.t1902 629.652
R8851 VPWR.t381 VPWR.n1848 629.652
R8852 VPWR.n1839 VPWR.t533 629.652
R8853 VPWR.t1804 VPWR.n1838 629.652
R8854 VPWR.n1829 VPWR.t973 629.652
R8855 VPWR.t1790 VPWR.n1828 629.652
R8856 VPWR.n1819 VPWR.t201 629.652
R8857 VPWR.n2477 VPWR.t893 629.652
R8858 VPWR.t1139 VPWR.n2476 629.652
R8859 VPWR.n2467 VPWR.t769 629.652
R8860 VPWR.t1045 VPWR.n2466 629.652
R8861 VPWR.n2457 VPWR.t407 629.652
R8862 VPWR.t695 VPWR.n2456 629.652
R8863 VPWR.n2447 VPWR.t1748 629.652
R8864 VPWR.t288 VPWR.n2446 629.652
R8865 VPWR.n2437 VPWR.t1105 629.652
R8866 VPWR.t385 VPWR.n2436 629.652
R8867 VPWR.n2427 VPWR.t218 629.652
R8868 VPWR.t1157 VPWR.n2426 629.652
R8869 VPWR.n2417 VPWR.t539 629.652
R8870 VPWR.t1024 VPWR.n2416 629.652
R8871 VPWR.n2407 VPWR.t207 629.652
R8872 VPWR.n966 VPWR.t959 629.652
R8873 VPWR.n970 VPWR.t765 629.652
R8874 VPWR.n974 VPWR.t811 629.652
R8875 VPWR.n978 VPWR.t377 629.652
R8876 VPWR.n982 VPWR.t1188 629.652
R8877 VPWR.n986 VPWR.t1172 629.652
R8878 VPWR.n990 VPWR.t441 629.652
R8879 VPWR.n994 VPWR.t593 629.652
R8880 VPWR.n998 VPWR.t110 629.652
R8881 VPWR.n1002 VPWR.t433 629.652
R8882 VPWR.n1006 VPWR.t716 629.652
R8883 VPWR.n1010 VPWR.t1782 629.652
R8884 VPWR.n1014 VPWR.t1287 629.652
R8885 VPWR.n1018 VPWR.t885 629.652
R8886 VPWR.n1022 VPWR.t163 629.652
R8887 VPWR.n350 VPWR.t903 629.652
R8888 VPWR.t1210 VPWR.n349 629.652
R8889 VPWR.t777 VPWR.n345 629.652
R8890 VPWR.t1033 VPWR.n341 629.652
R8891 VPWR.t660 VPWR.n337 629.652
R8892 VPWR.t1754 VPWR.n333 629.652
R8893 VPWR.t1738 VPWR.n329 629.652
R8894 VPWR.t847 VPWR.n325 629.652
R8895 VPWR.t1896 VPWR.n321 629.652
R8896 VPWR.t367 VPWR.n317 629.652
R8897 VPWR.t527 VPWR.n313 629.652
R8898 VPWR.t1802 VPWR.n309 629.652
R8899 VPWR.t969 VPWR.n305 629.652
R8900 VPWR.t1788 VPWR.n301 629.652
R8901 VPWR.t195 VPWR.n297 629.652
R8902 VPWR.n1468 VPWR.t895 629.652
R8903 VPWR.n1475 VPWR.t1892 629.652
R8904 VPWR.n1481 VPWR.t825 629.652
R8905 VPWR.n1492 VPWR.t149 629.652
R8906 VPWR.n1493 VPWR.t505 629.652
R8907 VPWR.n1506 VPWR.t697 629.652
R8908 VPWR.n1507 VPWR.t485 629.652
R8909 VPWR.n1520 VPWR.t732 629.652
R8910 VPWR.n1521 VPWR.t1107 629.652
R8911 VPWR.n1536 VPWR.t387 629.652
R8912 VPWR.t220 VPWR.n1535 629.652
R8913 VPWR.n1761 VPWR.t1159 629.652
R8914 VPWR.t541 VPWR.n1760 629.652
R8915 VPWR.n1749 VPWR.t1026 629.652
R8916 VPWR.n1791 VPWR.t211 629.652
R8917 VPWR.n2506 VPWR.t1499 629.652
R8918 VPWR.n2507 VPWR.t1628 629.652
R8919 VPWR.n2518 VPWR.t1646 629.652
R8920 VPWR.n2519 VPWR.t1408 629.652
R8921 VPWR.n2530 VPWR.t1516 629.652
R8922 VPWR.n2531 VPWR.t1671 629.652
R8923 VPWR.n2542 VPWR.t1395 629.652
R8924 VPWR.n2543 VPWR.t1430 629.652
R8925 VPWR.n2554 VPWR.t1558 629.652
R8926 VPWR.n2555 VPWR.t1668 629.652
R8927 VPWR.n2566 VPWR.t1435 629.652
R8928 VPWR.n2567 VPWR.t1453 629.652
R8929 VPWR.n2578 VPWR.t1581 629.652
R8930 VPWR.n2579 VPWR.t1714 629.652
R8931 VPWR.n2590 VPWR.t1354 629.652
R8932 VPWR.n1594 VPWR.t1370 629.652
R8933 VPWR.t1506 VPWR.n1593 629.652
R8934 VPWR.n1182 VPWR.t1519 629.652
R8935 VPWR.n1185 VPWR.t1679 629.652
R8936 VPWR.n1220 VPWR.t1400 629.652
R8937 VPWR.t1547 VPWR.n1219 629.652
R8938 VPWR.t1655 VPWR.n1216 629.652
R8939 VPWR.t1695 VPWR.n1213 629.652
R8940 VPWR.t1440 VPWR.n1205 629.652
R8941 VPWR.t1544 VPWR.n1202 629.652
R8942 VPWR.t1703 VPWR.n1199 629.652
R8943 VPWR.t1722 VPWR.n1191 629.652
R8944 VPWR.t1466 VPWR.n1188 629.652
R8945 VPWR.n1740 VPWR.t1595 629.652
R8946 VPWR.t1623 VPWR.n1739 629.652
R8947 VPWR.n2836 VPWR.t668 531.804
R8948 VPWR.n2855 VPWR.t668 531.804
R8949 VPWR.n2851 VPWR.n2850 504.707
R8950 VPWR.t1726 VPWR.t1268 486.048
R8951 VPWR.t1133 VPWR.t130 486.048
R8952 VPWR.t1823 VPWR.t805 486.048
R8953 VPWR.t1336 VPWR.t1822 486.048
R8954 VPWR.t1267 VPWR.t1125 486.048
R8955 VPWR.t1161 VPWR.t454 486.048
R8956 VPWR.t453 VPWR.t1260 486.048
R8957 VPWR.t603 VPWR.t1266 486.048
R8958 VPWR.t132 VPWR.t853 486.048
R8959 VPWR.t439 VPWR.t455 486.048
R8960 VPWR.t1821 VPWR.t1918 486.048
R8961 VPWR.t94 VPWR.t1820 486.048
R8962 VPWR.t452 VPWR.t1238 486.048
R8963 VPWR.t891 VPWR.t451 486.048
R8964 VPWR.t450 VPWR.t873 486.048
R8965 VPWR.t1488 VPWR.t131 486.048
R8966 VPWR.t901 VPWR.t86 486.048
R8967 VPWR.t671 VPWR.t1206 486.048
R8968 VPWR.t78 VPWR.t779 486.048
R8969 VPWR.t77 VPWR.t1031 486.048
R8970 VPWR.t85 VPWR.t656 486.048
R8971 VPWR.t1851 VPWR.t1750 486.048
R8972 VPWR.t1850 VPWR.t1734 486.048
R8973 VPWR.t84 VPWR.t843 486.048
R8974 VPWR.t83 VPWR.t730 486.048
R8975 VPWR.t670 VPWR.t365 486.048
R8976 VPWR.t76 VPWR.t523 486.048
R8977 VPWR.t75 VPWR.t1800 486.048
R8978 VPWR.t1849 VPWR.t965 486.048
R8979 VPWR.t1848 VPWR.t1786 486.048
R8980 VPWR.t79 VPWR.t1014 486.048
R8981 VPWR.t672 VPWR.t1706 486.048
R8982 VPWR.t618 VPWR.t1001 486.048
R8983 VPWR.t864 VPWR.t267 486.048
R8984 VPWR.t819 VPWR.t1776 486.048
R8985 VPWR.t1775 VPWR.t375 486.048
R8986 VPWR.t1186 VPWR.t1000 486.048
R8987 VPWR.t862 VPWR.t1170 486.048
R8988 VPWR.t499 VPWR.t861 486.048
R8989 VPWR.t999 VPWR.t6 486.048
R8990 VPWR.t108 VPWR.t866 486.048
R8991 VPWR.t863 VPWR.t427 486.048
R8992 VPWR.t714 VPWR.t1774 486.048
R8993 VPWR.t1773 VPWR.t1149 486.048
R8994 VPWR.t1285 VPWR.t860 486.048
R8995 VPWR.t859 VPWR.t41 486.048
R8996 VPWR.t161 VPWR.t1777 486.048
R8997 VPWR.t865 VPWR.t1555 486.048
R8998 VPWR.t907 VPWR.t352 486.048
R8999 VPWR.t1137 VPWR.t424 486.048
R9000 VPWR.t771 VPWR.t328 486.048
R9001 VPWR.t1043 VPWR.t327 486.048
R9002 VPWR.t405 VPWR.t351 486.048
R9003 VPWR.t1762 VPWR.t422 486.048
R9004 VPWR.t1746 VPWR.t421 486.048
R9005 VPWR.t286 VPWR.t350 486.048
R9006 VPWR.t1904 VPWR.t349 486.048
R9007 VPWR.t383 VPWR.t423 486.048
R9008 VPWR.t216 VPWR.t354 486.048
R9009 VPWR.t1155 VPWR.t353 486.048
R9010 VPWR.t537 VPWR.t420 486.048
R9011 VPWR.t1792 VPWR.t419 486.048
R9012 VPWR.t205 VPWR.t418 486.048
R9013 VPWR.t1663 VPWR.t348 486.048
R9014 VPWR.t1295 VPWR.t568 486.048
R9015 VPWR.t141 VPWR.t100 486.048
R9016 VPWR.t502 VPWR.t791 486.048
R9017 VPWR.t687 VPWR.t839 486.048
R9018 VPWR.t567 VPWR.t718 486.048
R9019 VPWR.t63 VPWR.t319 486.048
R9020 VPWR.t318 VPWR.t1867 486.048
R9021 VPWR.t571 VPWR.t566 486.048
R9022 VPWR.t565 VPWR.t1224 486.048
R9023 VPWR.t342 VPWR.t320 486.048
R9024 VPWR.t838 VPWR.t1843 486.048
R9025 VPWR.t1806 VPWR.t837 486.048
R9026 VPWR.t317 VPWR.t1252 486.048
R9027 VPWR.t10 VPWR.t504 486.048
R9028 VPWR.t503 VPWR.t1006 486.048
R9029 VPWR.t1389 VPWR.t101 486.048
R9030 VPWR.t961 VPWR.t1169 486.048
R9031 VPWR.t176 VPWR.t1131 486.048
R9032 VPWR.t1313 VPWR.t809 486.048
R9033 VPWR.t549 VPWR.t1332 486.048
R9034 VPWR.t1168 VPWR.t1123 486.048
R9035 VPWR.t691 VPWR.t1178 486.048
R9036 VPWR.t690 VPWR.t1258 486.048
R9037 VPWR.t1167 VPWR.t601 486.048
R9038 VPWR.t178 VPWR.t581 486.048
R9039 VPWR.t692 VPWR.t435 486.048
R9040 VPWR.t548 VPWR.t1916 486.048
R9041 VPWR.t547 VPWR.t90 486.048
R9042 VPWR.t689 VPWR.t1236 486.048
R9043 VPWR.t1315 VPWR.t887 486.048
R9044 VPWR.t1314 VPWR.t869 486.048
R9045 VPWR.t177 VPWR.t1496 486.048
R9046 VPWR.t1728 VPWR.t30 486.048
R9047 VPWR.t1265 VPWR.t507 486.048
R9048 VPWR.t799 VPWR.t1300 486.048
R9049 VPWR.t1299 VPWR.t1338 486.048
R9050 VPWR.t137 VPWR.t29 486.048
R9051 VPWR.t1263 VPWR.t1165 486.048
R9052 VPWR.t1859 VPWR.t1262 486.048
R9053 VPWR.t28 VPWR.t67 486.048
R9054 VPWR.t857 VPWR.t27 486.048
R9055 VPWR.t1264 VPWR.t334 486.048
R9056 VPWR.t1115 VPWR.t1298 486.048
R9057 VPWR.t1297 VPWR.t1078 486.048
R9058 VPWR.t1242 VPWR.t1303 486.048
R9059 VPWR.t1302 VPWR.t20 486.048
R9060 VPWR.t875 VPWR.t1301 486.048
R9061 VPWR.t26 VPWR.t1456 486.048
R9062 VPWR.t616 VPWR.t1310 486.048
R9063 VPWR.t263 VPWR.t1305 486.048
R9064 VPWR.t807 VPWR.t170 486.048
R9065 VPWR.t373 VPWR.t169 486.048
R9066 VPWR.t1324 VPWR.t1309 486.048
R9067 VPWR.t561 VPWR.t175 486.048
R9068 VPWR.t495 VPWR.t174 486.048
R9069 VPWR.t4 VPWR.t1308 486.048
R9070 VPWR.t104 VPWR.t1307 486.048
R9071 VPWR.t425 VPWR.t1304 486.048
R9072 VPWR.t710 VPWR.t168 486.048
R9073 VPWR.t1147 VPWR.t167 486.048
R9074 VPWR.t1283 VPWR.t173 486.048
R9075 VPWR.t39 VPWR.t172 486.048
R9076 VPWR.t187 VPWR.t171 486.048
R9077 VPWR.t1561 VPWR.t1306 486.048
R9078 VPWR.t1016 VPWR.t667 486.048
R9079 VPWR.t143 VPWR.t662 486.048
R9080 VPWR.t293 VPWR.t789 486.048
R9081 VPWR.t634 VPWR.t292 486.048
R9082 VPWR.t666 VPWR.t720 486.048
R9083 VPWR.t1812 VPWR.t282 486.048
R9084 VPWR.t281 VPWR.t1869 486.048
R9085 VPWR.t573 VPWR.t665 486.048
R9086 VPWR.t664 VPWR.t1226 486.048
R9087 VPWR.t344 VPWR.t283 486.048
R9088 VPWR.t291 VPWR.t1824 486.048
R9089 VPWR.t1808 VPWR.t290 486.048
R9090 VPWR.t296 VPWR.t942 486.048
R9091 VPWR.t12 VPWR.t295 486.048
R9092 VPWR.t294 VPWR.t1010 486.048
R9093 VPWR.t1384 VPWR.t663 486.048
R9094 VPWR.t614 VPWR.t997 486.048
R9095 VPWR.t1885 VPWR.t261 486.048
R9096 VPWR.t607 VPWR.t821 486.048
R9097 VPWR.t606 VPWR.t371 486.048
R9098 VPWR.t996 VPWR.t1322 486.048
R9099 VPWR.t1883 VPWR.t559 486.048
R9100 VPWR.t611 VPWR.t493 486.048
R9101 VPWR.t995 VPWR.t2 486.048
R9102 VPWR.t1887 VPWR.t102 486.048
R9103 VPWR.t1884 VPWR.t591 486.048
R9104 VPWR.t605 VPWR.t708 486.048
R9105 VPWR.t1856 VPWR.t1145 486.048
R9106 VPWR.t610 VPWR.t1281 486.048
R9107 VPWR.t609 VPWR.t37 486.048
R9108 VPWR.t608 VPWR.t185 486.048
R9109 VPWR.t1886 VPWR.t1568 486.048
R9110 VPWR.t1018 VPWR.t1269 486.048
R9111 VPWR.t145 VPWR.t1925 486.048
R9112 VPWR.t787 VPWR.t1273 486.048
R9113 VPWR.t636 VPWR.t1272 486.048
R9114 VPWR.t722 VPWR.t949 486.048
R9115 VPWR.t1814 VPWR.t1278 486.048
R9116 VPWR.t1871 VPWR.t1277 486.048
R9117 VPWR.t575 VPWR.t948 486.048
R9118 VPWR.t724 VPWR.t947 486.048
R9119 VPWR.t346 VPWR.t951 486.048
R9120 VPWR.t1826 VPWR.t1271 486.048
R9121 VPWR.t1810 VPWR.t1270 486.048
R9122 VPWR.t944 VPWR.t1276 486.048
R9123 VPWR.t14 VPWR.t1275 486.048
R9124 VPWR.t1012 VPWR.t1274 486.048
R9125 VPWR.t1376 VPWR.t946 486.048
R9126 VPWR.t905 VPWR.t626 486.048
R9127 VPWR.t980 VPWR.t1216 486.048
R9128 VPWR.t773 VPWR.t1772 486.048
R9129 VPWR.t1771 VPWR.t1039 486.048
R9130 VPWR.t403 VPWR.t625 486.048
R9131 VPWR.t978 VPWR.t1760 486.048
R9132 VPWR.t1744 VPWR.t977 486.048
R9133 VPWR.t624 VPWR.t851 486.048
R9134 VPWR.t1902 VPWR.t623 486.048
R9135 VPWR.t979 VPWR.t381 486.048
R9136 VPWR.t533 VPWR.t1770 486.048
R9137 VPWR.t627 VPWR.t1804 486.048
R9138 VPWR.t973 VPWR.t976 486.048
R9139 VPWR.t975 VPWR.t1790 486.048
R9140 VPWR.t201 VPWR.t998 486.048
R9141 VPWR.t622 VPWR.t1676 486.048
R9142 VPWR.t893 VPWR.t1921 486.048
R9143 VPWR.t1180 VPWR.t1139 486.048
R9144 VPWR.t769 VPWR.t940 486.048
R9145 VPWR.t1924 VPWR.t1045 486.048
R9146 VPWR.t407 VPWR.t1920 486.048
R9147 VPWR.t459 VPWR.t695 486.048
R9148 VPWR.t1748 VPWR.t458 486.048
R9149 VPWR.t1183 VPWR.t288 486.048
R9150 VPWR.t1105 VPWR.t1182 486.048
R9151 VPWR.t460 VPWR.t385 486.048
R9152 VPWR.t218 VPWR.t1923 486.048
R9153 VPWR.t1922 VPWR.t1157 486.048
R9154 VPWR.t539 VPWR.t457 486.048
R9155 VPWR.t456 VPWR.t1024 486.048
R9156 VPWR.t207 VPWR.t941 486.048
R9157 VPWR.t1181 VPWR.t1658 486.048
R9158 VPWR.t959 VPWR.t1836 486.048
R9159 VPWR.t765 VPWR.t701 486.048
R9160 VPWR.t811 VPWR.t304 486.048
R9161 VPWR.t377 VPWR.t89 486.048
R9162 VPWR.t1188 VPWR.t1112 486.048
R9163 VPWR.t1172 VPWR.t699 486.048
R9164 VPWR.t441 VPWR.t308 486.048
R9165 VPWR.t593 VPWR.t1111 486.048
R9166 VPWR.t110 VPWR.t1110 486.048
R9167 VPWR.t433 VPWR.t700 486.048
R9168 VPWR.t716 VPWR.t88 486.048
R9169 VPWR.t1782 VPWR.t87 486.048
R9170 VPWR.t1287 VPWR.t307 486.048
R9171 VPWR.t885 VPWR.t306 486.048
R9172 VPWR.t163 VPWR.t305 486.048
R9173 VPWR.t1528 VPWR.t1109 486.048
R9174 VPWR.t903 VPWR.t676 486.048
R9175 VPWR.t1878 VPWR.t1210 486.048
R9176 VPWR.t1881 VPWR.t777 486.048
R9177 VPWR.t1880 VPWR.t1033 486.048
R9178 VPWR.t675 VPWR.t660 486.048
R9179 VPWR.t1876 VPWR.t1754 486.048
R9180 VPWR.t1875 VPWR.t1738 486.048
R9181 VPWR.t674 VPWR.t847 486.048
R9182 VPWR.t673 VPWR.t1896 486.048
R9183 VPWR.t1877 VPWR.t367 486.048
R9184 VPWR.t678 VPWR.t527 486.048
R9185 VPWR.t677 VPWR.t1802 486.048
R9186 VPWR.t1874 VPWR.t969 486.048
R9187 VPWR.t1873 VPWR.t1788 486.048
R9188 VPWR.t1882 VPWR.t195 486.048
R9189 VPWR.t1879 VPWR.t1698 486.048
R9190 VPWR.t895 VPWR.t1433 486.048
R9191 VPWR.t1892 VPWR.t1564 486.048
R9192 VPWR.t825 VPWR.t1693 486.048
R9193 VPWR.t149 VPWR.t1349 486.048
R9194 VPWR.t505 VPWR.t1459 486.048
R9195 VPWR.t1614 VPWR.t697 486.048
R9196 VPWR.t485 VPWR.t1616 486.048
R9197 VPWR.t1464 VPWR.t732 486.048
R9198 VPWR.t1107 VPWR.t1494 486.048
R9199 VPWR.t1612 VPWR.t387 486.048
R9200 VPWR.t1363 VPWR.t220 486.048
R9201 VPWR.t1382 VPWR.t1159 486.048
R9202 VPWR.t1626 VPWR.t541 486.048
R9203 VPWR.t1026 VPWR.t1644 486.048
R9204 VPWR.t1682 VPWR.t211 486.048
R9205 VPWR.t1639 VPWR.t1514 486.048
R9206 VPWR.t1499 VPWR.t1368 486.048
R9207 VPWR.t1628 VPWR.t1504 486.048
R9208 VPWR.t1634 VPWR.t1646 486.048
R9209 VPWR.t1408 VPWR.t1674 486.048
R9210 VPWR.t1398 VPWR.t1516 486.048
R9211 VPWR.t1671 VPWR.t1542 486.048
R9212 VPWR.t1566 VPWR.t1395 486.048
R9213 VPWR.t1430 VPWR.t1403 486.048
R9214 VPWR.t1438 VPWR.t1558 486.048
R9215 VPWR.t1668 VPWR.t1540 486.048
R9216 VPWR.t1701 VPWR.t1435 486.048
R9217 VPWR.t1453 VPWR.t1720 486.048
R9218 VPWR.t1574 VPWR.t1581 486.048
R9219 VPWR.t1714 VPWR.t1593 486.048
R9220 VPWR.t1618 VPWR.t1354 486.048
R9221 VPWR.t1590 VPWR.t1469 486.048
R9222 VPWR.t1370 VPWR.t1642 486.048
R9223 VPWR.t1387 VPWR.t1506 486.048
R9224 VPWR.t1519 VPWR.t1512 486.048
R9225 VPWR.t1679 VPWR.t1553 486.048
R9226 VPWR.t1400 VPWR.t1661 486.048
R9227 VPWR.t1428 VPWR.t1547 486.048
R9228 VPWR.t1443 VPWR.t1655 486.048
R9229 VPWR.t1666 VPWR.t1695 486.048
R9230 VPWR.t1709 VPWR.t1440 486.048
R9231 VPWR.t1426 VPWR.t1544 486.048
R9232 VPWR.t1579 VPWR.t1703 486.048
R9233 VPWR.t1601 VPWR.t1722 486.048
R9234 VPWR.t1451 VPWR.t1466 486.048
R9235 VPWR.t1477 VPWR.t1595 486.048
R9236 VPWR.t1502 VPWR.t1623 486.048
R9237 VPWR.t1474 VPWR.t1347 486.048
R9238 VPWR.t1268 VPWR.t1074 463.954
R9239 VPWR.t130 VPWR.t957 463.954
R9240 VPWR.t1129 VPWR.t1823 463.954
R9241 VPWR.t1822 VPWR.t827 463.954
R9242 VPWR.t153 VPWR.t1267 463.954
R9243 VPWR.t454 VPWR.t1121 463.954
R9244 VPWR.t1176 VPWR.t453 463.954
R9245 VPWR.t1266 VPWR.t1256 463.954
R9246 VPWR.t736 VPWR.t132 463.954
R9247 VPWR.t455 VPWR.t579 463.954
R9248 VPWR.t431 VPWR.t1821 463.954
R9249 VPWR.t1820 VPWR.t1914 463.954
R9250 VPWR.t1780 VPWR.t452 463.954
R9251 VPWR.t451 VPWR.t545 463.954
R9252 VPWR.t883 VPWR.t450 463.954
R9253 VPWR.t131 VPWR.t181 463.954
R9254 VPWR.t86 VPWR.t1063 463.954
R9255 VPWR.t1020 VPWR.t671 463.954
R9256 VPWR.t1228 VPWR.t78 463.954
R9257 VPWR.t803 VPWR.t77 463.954
R9258 VPWR.t679 VPWR.t85 463.954
R9259 VPWR.t112 VPWR.t1851 463.954
R9260 VPWR.t1816 VPWR.t1850 463.954
R9261 VPWR.t1730 VPWR.t84 463.954
R9262 VPWR.t65 VPWR.t83 463.954
R9263 VPWR.t726 VPWR.t670 463.954
R9264 VPWR.t355 VPWR.t76 463.954
R9265 VPWR.t1828 VPWR.t75 463.954
R9266 VPWR.t96 VPWR.t1849 463.954
R9267 VPWR.t1240 VPWR.t1848 463.954
R9268 VPWR.t16 VPWR.t79 463.954
R9269 VPWR.t877 VPWR.t672 463.954
R9270 VPWR.t1001 VPWR.t1049 463.954
R9271 VPWR.t1910 VPWR.t864 463.954
R9272 VPWR.t1776 VPWR.t259 463.954
R9273 VPWR.t781 VPWR.t1775 463.954
R9274 VPWR.t1000 VPWR.t1041 463.954
R9275 VPWR.t1320 VPWR.t862 463.954
R9276 VPWR.t861 VPWR.t557 463.954
R9277 VPWR.t491 VPWR.t999 463.954
R9278 VPWR.t866 VPWR.t849 463.954
R9279 VPWR.t519 VPWR.t863 463.954
R9280 VPWR.t1774 VPWR.t587 463.954
R9281 VPWR.t706 VPWR.t1773 463.954
R9282 VPWR.t860 VPWR.t1141 463.954
R9283 VPWR.t971 VPWR.t859 463.954
R9284 VPWR.t1777 VPWR.t477 463.954
R9285 VPWR.t203 VPWR.t865 463.954
R9286 VPWR.t352 VPWR.t1057 463.954
R9287 VPWR.t424 VPWR.t897 463.954
R9288 VPWR.t328 VPWR.t1212 463.954
R9289 VPWR.t327 VPWR.t795 463.954
R9290 VPWR.t351 VPWR.t685 463.954
R9291 VPWR.t422 VPWR.t399 463.954
R9292 VPWR.t421 VPWR.t1756 463.954
R9293 VPWR.t350 VPWR.t1740 463.954
R9294 VPWR.t349 VPWR.t73 463.954
R9295 VPWR.t423 VPWR.t1898 463.954
R9296 VPWR.t354 VPWR.t361 463.954
R9297 VPWR.t353 VPWR.t529 463.954
R9298 VPWR.t420 VPWR.t1796 463.954
R9299 VPWR.t419 VPWR.t1248 463.954
R9300 VPWR.t418 VPWR.t33 463.954
R9301 VPWR.t348 VPWR.t1004 463.954
R9302 VPWR.t568 VPWR.t1069 463.954
R9303 VPWR.t100 VPWR.t479 463.954
R9304 VPWR.t509 VPWR.t502 463.954
R9305 VPWR.t839 VPWR.t817 463.954
R9306 VPWR.t379 VPWR.t567 463.954
R9307 VPWR.t319 VPWR.t139 463.954
R9308 VPWR.t57 VPWR.t318 463.954
R9309 VPWR.t566 VPWR.t1861 463.954
R9310 VPWR.t595 VPWR.t565 463.954
R9311 VPWR.t320 VPWR.t1218 463.954
R9312 VPWR.t336 VPWR.t838 463.954
R9313 VPWR.t837 VPWR.t1837 463.954
R9314 VPWR.t919 VPWR.t317 463.954
R9315 VPWR.t504 VPWR.t1289 463.954
R9316 VPWR.t22 VPWR.t503 463.954
R9317 VPWR.t101 VPWR.t165 463.954
R9318 VPWR.t1169 VPWR.t1076 463.954
R9319 VPWR.t620 VPWR.t176 463.954
R9320 VPWR.t767 VPWR.t1313 463.954
R9321 VPWR.t829 VPWR.t549 463.954
R9322 VPWR.t151 VPWR.t1168 463.954
R9323 VPWR.t1190 VPWR.t691 463.954
R9324 VPWR.t1174 VPWR.t690 463.954
R9325 VPWR.t1254 VPWR.t1167 463.954
R9326 VPWR.t734 VPWR.t178 463.954
R9327 VPWR.t577 VPWR.t692 463.954
R9328 VPWR.t429 VPWR.t548 463.954
R9329 VPWR.t1912 VPWR.t547 463.954
R9330 VPWR.t1778 VPWR.t689 463.954
R9331 VPWR.t543 VPWR.t1315 463.954
R9332 VPWR.t881 VPWR.t1314 463.954
R9333 VPWR.t179 VPWR.t177 463.954
R9334 VPWR.t30 VPWR.t1072 463.954
R9335 VPWR.t1724 VPWR.t1265 463.954
R9336 VPWR.t1300 VPWR.t1135 463.954
R9337 VPWR.t823 VPWR.t1299 463.954
R9338 VPWR.t29 VPWR.t369 463.954
R9339 VPWR.t1127 VPWR.t1263 463.954
R9340 VPWR.t1262 VPWR.t1163 463.954
R9341 VPWR.t1857 VPWR.t28 463.954
R9342 VPWR.t27 VPWR.t0 463.954
R9343 VPWR.t855 VPWR.t1264 463.954
R9344 VPWR.t1298 VPWR.t437 463.954
R9345 VPWR.t1113 VPWR.t1297 463.954
R9346 VPWR.t1303 VPWR.t92 463.954
R9347 VPWR.t1279 VPWR.t1302 463.954
R9348 VPWR.t1301 VPWR.t889 463.954
R9349 VPWR.t183 VPWR.t26 463.954
R9350 VPWR.t1310 VPWR.t1051 463.954
R9351 VPWR.t1305 VPWR.t1908 463.954
R9352 VPWR.t170 VPWR.t257 463.954
R9353 VPWR.t169 VPWR.t783 463.954
R9354 VPWR.t1309 VPWR.t1037 463.954
R9355 VPWR.t175 VPWR.t1318 463.954
R9356 VPWR.t174 VPWR.t555 463.954
R9357 VPWR.t1308 VPWR.t489 463.954
R9358 VPWR.t1307 VPWR.t845 463.954
R9359 VPWR.t1304 VPWR.t517 463.954
R9360 VPWR.t168 VPWR.t585 463.954
R9361 VPWR.t167 VPWR.t704 463.954
R9362 VPWR.t173 VPWR.t1153 463.954
R9363 VPWR.t172 VPWR.t967 463.954
R9364 VPWR.t171 VPWR.t1890 463.954
R9365 VPWR.t1306 VPWR.t199 463.954
R9366 VPWR.t667 VPWR.t1067 463.954
R9367 VPWR.t662 VPWR.t481 463.954
R9368 VPWR.t511 VPWR.t293 463.954
R9369 VPWR.t292 VPWR.t815 463.954
R9370 VPWR.t1330 VPWR.t666 463.954
R9371 VPWR.t282 VPWR.t1202 463.954
R9372 VPWR.t59 VPWR.t281 463.954
R9373 VPWR.t665 VPWR.t1863 463.954
R9374 VPWR.t597 VPWR.t664 463.954
R9375 VPWR.t283 VPWR.t1220 463.954
R9376 VPWR.t338 VPWR.t291 463.954
R9377 VPWR.t290 VPWR.t1839 463.954
R9378 VPWR.t921 VPWR.t296 463.954
R9379 VPWR.t295 VPWR.t1291 463.954
R9380 VPWR.t24 VPWR.t294 463.954
R9381 VPWR.t663 VPWR.t867 463.954
R9382 VPWR.t997 VPWR.t1053 463.954
R9383 VPWR.t1906 VPWR.t1885 463.954
R9384 VPWR.t255 VPWR.t607 463.954
R9385 VPWR.t785 VPWR.t606 463.954
R9386 VPWR.t1035 VPWR.t996 463.954
R9387 VPWR.t1316 VPWR.t1883 463.954
R9388 VPWR.t553 VPWR.t611 463.954
R9389 VPWR.t487 VPWR.t995 463.954
R9390 VPWR.t841 VPWR.t1887 463.954
R9391 VPWR.t515 VPWR.t1884 463.954
R9392 VPWR.t583 VPWR.t605 463.954
R9393 VPWR.t702 VPWR.t1856 463.954
R9394 VPWR.t1151 VPWR.t610 463.954
R9395 VPWR.t963 VPWR.t609 463.954
R9396 VPWR.t1888 VPWR.t608 463.954
R9397 VPWR.t197 VPWR.t1886 463.954
R9398 VPWR.t1269 VPWR.t1065 463.954
R9399 VPWR.t1925 VPWR.t483 463.954
R9400 VPWR.t1273 VPWR.t513 463.954
R9401 VPWR.t1272 VPWR.t813 463.954
R9402 VPWR.t949 VPWR.t1334 463.954
R9403 VPWR.t1278 VPWR.t1204 463.954
R9404 VPWR.t1277 VPWR.t61 463.954
R9405 VPWR.t948 VPWR.t1865 463.954
R9406 VPWR.t947 VPWR.t599 463.954
R9407 VPWR.t951 VPWR.t1222 463.954
R9408 VPWR.t1271 VPWR.t340 463.954
R9409 VPWR.t1270 VPWR.t1841 463.954
R9410 VPWR.t1276 VPWR.t923 463.954
R9411 VPWR.t1275 VPWR.t1293 463.954
R9412 VPWR.t1274 VPWR.t8 463.954
R9413 VPWR.t946 VPWR.t871 463.954
R9414 VPWR.t626 VPWR.t1059 463.954
R9415 VPWR.t909 VPWR.t980 463.954
R9416 VPWR.t1772 VPWR.t1208 463.954
R9417 VPWR.t797 VPWR.t1771 463.954
R9418 VPWR.t625 VPWR.t683 463.954
R9419 VPWR.t658 VPWR.t978 463.954
R9420 VPWR.t977 VPWR.t1752 463.954
R9421 VPWR.t1736 VPWR.t624 463.954
R9422 VPWR.t623 VPWR.t71 463.954
R9423 VPWR.t1894 VPWR.t979 463.954
R9424 VPWR.t1770 VPWR.t359 463.954
R9425 VPWR.t525 VPWR.t627 463.954
R9426 VPWR.t976 VPWR.t1794 463.954
R9427 VPWR.t1246 VPWR.t975 463.954
R9428 VPWR.t998 VPWR.t31 463.954
R9429 VPWR.t1002 VPWR.t622 463.954
R9430 VPWR.t1921 VPWR.t1055 463.954
R9431 VPWR.t899 VPWR.t1180 463.954
R9432 VPWR.t940 VPWR.t1214 463.954
R9433 VPWR.t793 VPWR.t1924 463.954
R9434 VPWR.t1920 VPWR.t632 463.954
R9435 VPWR.t401 VPWR.t459 463.954
R9436 VPWR.t458 VPWR.t1758 463.954
R9437 VPWR.t1742 VPWR.t1183 463.954
R9438 VPWR.t1182 VPWR.t569 463.954
R9439 VPWR.t1900 VPWR.t460 463.954
R9440 VPWR.t1923 VPWR.t363 463.954
R9441 VPWR.t531 VPWR.t1922 463.954
R9442 VPWR.t457 VPWR.t1798 463.954
R9443 VPWR.t1250 VPWR.t456 463.954
R9444 VPWR.t941 VPWR.t1784 463.954
R9445 VPWR.t1008 VPWR.t1181 463.954
R9446 VPWR.t1836 VPWR.t1047 463.954
R9447 VPWR.t701 VPWR.t612 463.954
R9448 VPWR.t304 VPWR.t265 463.954
R9449 VPWR.t89 VPWR.t775 463.954
R9450 VPWR.t1112 VPWR.t147 463.954
R9451 VPWR.t699 VPWR.t1184 463.954
R9452 VPWR.t308 VPWR.t563 463.954
R9453 VPWR.t1111 VPWR.t497 463.954
R9454 VPWR.t1110 VPWR.t284 463.954
R9455 VPWR.t700 VPWR.t106 463.954
R9456 VPWR.t88 VPWR.t589 463.954
R9457 VPWR.t87 VPWR.t712 463.954
R9458 VPWR.t307 VPWR.t1143 463.954
R9459 VPWR.t306 VPWR.t535 463.954
R9460 VPWR.t305 VPWR.t35 463.954
R9461 VPWR.t1109 VPWR.t209 463.954
R9462 VPWR.t676 VPWR.t1061 463.954
R9463 VPWR.t1022 VPWR.t1878 463.954
R9464 VPWR.t1230 VPWR.t1881 463.954
R9465 VPWR.t801 VPWR.t1880 463.954
R9466 VPWR.t681 VPWR.t675 463.954
R9467 VPWR.t654 VPWR.t1876 463.954
R9468 VPWR.t1818 VPWR.t1875 463.954
R9469 VPWR.t1732 VPWR.t674 463.954
R9470 VPWR.t69 VPWR.t673 463.954
R9471 VPWR.t728 VPWR.t1877 463.954
R9472 VPWR.t357 VPWR.t678 463.954
R9473 VPWR.t521 VPWR.t677 463.954
R9474 VPWR.t98 VPWR.t1874 463.954
R9475 VPWR.t1244 VPWR.t1873 463.954
R9476 VPWR.t18 VPWR.t1882 463.954
R9477 VPWR.t879 VPWR.t1879 463.954
R9478 VPWR.t1433 VPWR.t1448 463.954
R9479 VPWR.t1564 VPWR.t1609 463.954
R9480 VPWR.t1693 VPWR.t1711 463.954
R9481 VPWR.t1349 VPWR.t1482 463.954
R9482 VPWR.t1459 VPWR.t1584 463.954
R9483 VPWR.t1606 VPWR.t1614 463.954
R9484 VPWR.t1616 VPWR.t1357 463.954
R9485 VPWR.t1479 VPWR.t1464 463.954
R9486 VPWR.t1494 VPWR.t1620 463.954
R9487 VPWR.t1636 VPWR.t1612 463.954
R9488 VPWR.t1379 VPWR.t1363 463.954
R9489 VPWR.t1509 VPWR.t1382 463.954
R9490 VPWR.t1550 VPWR.t1626 463.954
R9491 VPWR.t1644 VPWR.t1373 463.954
R9492 VPWR.t1423 VPWR.t1682 463.954
R9493 VPWR.t1514 VPWR.t1531 463.954
R9494 VPWR.t1368 VPWR.t1392 463.954
R9495 VPWR.t1504 VPWR.t1537 463.954
R9496 VPWR.t1649 VPWR.t1634 463.954
R9497 VPWR.t1674 VPWR.t1414 463.954
R9498 VPWR.t1525 VPWR.t1398 463.954
R9499 VPWR.t1542 VPWR.t1534 463.954
R9500 VPWR.t1690 VPWR.t1566 463.954
R9501 VPWR.t1403 VPWR.t1411 463.954
R9502 VPWR.t1571 VPWR.t1438 463.954
R9503 VPWR.t1540 VPWR.t1587 463.954
R9504 VPWR.t1717 VPWR.t1701 463.954
R9505 VPWR.t1720 VPWR.t1461 463.954
R9506 VPWR.t1491 VPWR.t1574 463.954
R9507 VPWR.t1593 VPWR.t1341 463.954
R9508 VPWR.t1360 VPWR.t1618 463.954
R9509 VPWR.t1469 VPWR.t1485 463.954
R9510 VPWR.t1642 VPWR.t1652 463.954
R9511 VPWR.t1420 VPWR.t1387 463.954
R9512 VPWR.t1512 VPWR.t1522 463.954
R9513 VPWR.t1553 VPWR.t1687 463.954
R9514 VPWR.t1661 VPWR.t1405 463.954
R9515 VPWR.t1417 VPWR.t1428 463.954
R9516 VPWR.t1576 VPWR.t1443 463.954
R9517 VPWR.t1684 VPWR.t1666 463.954
R9518 VPWR.t1445 VPWR.t1709 463.954
R9519 VPWR.t1471 VPWR.t1426 463.954
R9520 VPWR.t1598 VPWR.t1579 463.954
R9521 VPWR.t1344 VPWR.t1601 463.954
R9522 VPWR.t1365 VPWR.t1451 463.954
R9523 VPWR.t1603 VPWR.t1477 463.954
R9524 VPWR.t1631 VPWR.t1502 463.954
R9525 VPWR.t1347 VPWR.t1351 463.954
R9526 VPWR.n2626 VPWR.t116 428.822
R9527 VPWR.n1595 VPWR.n1594 376.045
R9528 VPWR.n2506 VPWR.n2505 376.045
R9529 VPWR.n1468 VPWR.n1467 376.045
R9530 VPWR.n351 VPWR.n350 376.045
R9531 VPWR.n2568 VPWR.n2567 376.045
R9532 VPWR.n1535 VPWR.n1534 376.045
R9533 VPWR.n349 VPWR.n348 376.045
R9534 VPWR.n2508 VPWR.n2507 376.045
R9535 VPWR.n966 VPWR.n965 376.045
R9536 VPWR.n2478 VPWR.n2477 376.045
R9537 VPWR.n2476 VPWR.n2475 376.045
R9538 VPWR.n321 VPWR.n320 376.045
R9539 VPWR.n2554 VPWR.n2553 376.045
R9540 VPWR.n974 VPWR.n973 376.045
R9541 VPWR.n2446 VPWR.n2445 376.045
R9542 VPWR.n325 VPWR.n324 376.045
R9543 VPWR.n2544 VPWR.n2543 376.045
R9544 VPWR.n1890 VPWR.n1889 376.045
R9545 VPWR.n1888 VPWR.n1887 376.045
R9546 VPWR.n1880 VPWR.n1879 376.045
R9547 VPWR.n390 VPWR.n389 376.045
R9548 VPWR.n394 VPWR.n393 376.045
R9549 VPWR.n398 VPWR.n397 376.045
R9550 VPWR.n2456 VPWR.n2455 376.045
R9551 VPWR.n333 VPWR.n332 376.045
R9552 VPWR.n2532 VPWR.n2531 376.045
R9553 VPWR.n1878 VPWR.n1877 376.045
R9554 VPWR.n406 VPWR.n405 376.045
R9555 VPWR.n2458 VPWR.n2457 376.045
R9556 VPWR.n337 VPWR.n336 376.045
R9557 VPWR.n2530 VPWR.n2529 376.045
R9558 VPWR.n2309 VPWR.n2308 376.045
R9559 VPWR.n2311 VPWR.n2310 376.045
R9560 VPWR.n2319 VPWR.n2318 376.045
R9561 VPWR.n2321 VPWR.n2320 376.045
R9562 VPWR.n2331 VPWR.n2330 376.045
R9563 VPWR.n2339 VPWR.n2338 376.045
R9564 VPWR.n2341 VPWR.n2340 376.045
R9565 VPWR.n2349 VPWR.n2348 376.045
R9566 VPWR.n2351 VPWR.n2350 376.045
R9567 VPWR.n2359 VPWR.n2358 376.045
R9568 VPWR.n2361 VPWR.n2360 376.045
R9569 VPWR.n2369 VPWR.n2368 376.045
R9570 VPWR.n2371 VPWR.n2370 376.045
R9571 VPWR.n2379 VPWR.n2378 376.045
R9572 VPWR.n2329 VPWR.n2328 376.045
R9573 VPWR.n543 VPWR.n542 376.045
R9574 VPWR.n541 VPWR.n540 376.045
R9575 VPWR.n537 VPWR.n536 376.045
R9576 VPWR.n533 VPWR.n532 376.045
R9577 VPWR.n525 VPWR.n524 376.045
R9578 VPWR.n521 VPWR.n520 376.045
R9579 VPWR.n517 VPWR.n516 376.045
R9580 VPWR.n513 VPWR.n512 376.045
R9581 VPWR.n509 VPWR.n508 376.045
R9582 VPWR.n505 VPWR.n504 376.045
R9583 VPWR.n501 VPWR.n500 376.045
R9584 VPWR.n497 VPWR.n496 376.045
R9585 VPWR.n493 VPWR.n492 376.045
R9586 VPWR.n489 VPWR.n488 376.045
R9587 VPWR.n529 VPWR.n528 376.045
R9588 VPWR.n2282 VPWR.n2281 376.045
R9589 VPWR.n2280 VPWR.n2279 376.045
R9590 VPWR.n2272 VPWR.n2271 376.045
R9591 VPWR.n2270 VPWR.n2269 376.045
R9592 VPWR.n2260 VPWR.n2259 376.045
R9593 VPWR.n2252 VPWR.n2251 376.045
R9594 VPWR.n2250 VPWR.n2249 376.045
R9595 VPWR.n2242 VPWR.n2241 376.045
R9596 VPWR.n2240 VPWR.n2239 376.045
R9597 VPWR.n2232 VPWR.n2231 376.045
R9598 VPWR.n2230 VPWR.n2229 376.045
R9599 VPWR.n2222 VPWR.n2221 376.045
R9600 VPWR.n2220 VPWR.n2219 376.045
R9601 VPWR.n2212 VPWR.n2211 376.045
R9602 VPWR.n2262 VPWR.n2261 376.045
R9603 VPWR.n582 VPWR.n581 376.045
R9604 VPWR.n586 VPWR.n585 376.045
R9605 VPWR.n590 VPWR.n589 376.045
R9606 VPWR.n594 VPWR.n593 376.045
R9607 VPWR.n602 VPWR.n601 376.045
R9608 VPWR.n606 VPWR.n605 376.045
R9609 VPWR.n610 VPWR.n609 376.045
R9610 VPWR.n614 VPWR.n613 376.045
R9611 VPWR.n618 VPWR.n617 376.045
R9612 VPWR.n622 VPWR.n621 376.045
R9613 VPWR.n626 VPWR.n625 376.045
R9614 VPWR.n630 VPWR.n629 376.045
R9615 VPWR.n634 VPWR.n633 376.045
R9616 VPWR.n638 VPWR.n637 376.045
R9617 VPWR.n598 VPWR.n597 376.045
R9618 VPWR.n2113 VPWR.n2112 376.045
R9619 VPWR.n2115 VPWR.n2114 376.045
R9620 VPWR.n2123 VPWR.n2122 376.045
R9621 VPWR.n2125 VPWR.n2124 376.045
R9622 VPWR.n2135 VPWR.n2134 376.045
R9623 VPWR.n2143 VPWR.n2142 376.045
R9624 VPWR.n2145 VPWR.n2144 376.045
R9625 VPWR.n2153 VPWR.n2152 376.045
R9626 VPWR.n2155 VPWR.n2154 376.045
R9627 VPWR.n2163 VPWR.n2162 376.045
R9628 VPWR.n2165 VPWR.n2164 376.045
R9629 VPWR.n2173 VPWR.n2172 376.045
R9630 VPWR.n2175 VPWR.n2174 376.045
R9631 VPWR.n2183 VPWR.n2182 376.045
R9632 VPWR.n2133 VPWR.n2132 376.045
R9633 VPWR.n735 VPWR.n734 376.045
R9634 VPWR.n733 VPWR.n732 376.045
R9635 VPWR.n729 VPWR.n728 376.045
R9636 VPWR.n725 VPWR.n724 376.045
R9637 VPWR.n717 VPWR.n716 376.045
R9638 VPWR.n713 VPWR.n712 376.045
R9639 VPWR.n709 VPWR.n708 376.045
R9640 VPWR.n705 VPWR.n704 376.045
R9641 VPWR.n701 VPWR.n700 376.045
R9642 VPWR.n697 VPWR.n696 376.045
R9643 VPWR.n693 VPWR.n692 376.045
R9644 VPWR.n689 VPWR.n688 376.045
R9645 VPWR.n685 VPWR.n684 376.045
R9646 VPWR.n681 VPWR.n680 376.045
R9647 VPWR.n721 VPWR.n720 376.045
R9648 VPWR.n2086 VPWR.n2085 376.045
R9649 VPWR.n2084 VPWR.n2083 376.045
R9650 VPWR.n2076 VPWR.n2075 376.045
R9651 VPWR.n2074 VPWR.n2073 376.045
R9652 VPWR.n2064 VPWR.n2063 376.045
R9653 VPWR.n2056 VPWR.n2055 376.045
R9654 VPWR.n2054 VPWR.n2053 376.045
R9655 VPWR.n2046 VPWR.n2045 376.045
R9656 VPWR.n2044 VPWR.n2043 376.045
R9657 VPWR.n2036 VPWR.n2035 376.045
R9658 VPWR.n2034 VPWR.n2033 376.045
R9659 VPWR.n2026 VPWR.n2025 376.045
R9660 VPWR.n2024 VPWR.n2023 376.045
R9661 VPWR.n2016 VPWR.n2015 376.045
R9662 VPWR.n2066 VPWR.n2065 376.045
R9663 VPWR.n774 VPWR.n773 376.045
R9664 VPWR.n778 VPWR.n777 376.045
R9665 VPWR.n782 VPWR.n781 376.045
R9666 VPWR.n786 VPWR.n785 376.045
R9667 VPWR.n794 VPWR.n793 376.045
R9668 VPWR.n798 VPWR.n797 376.045
R9669 VPWR.n802 VPWR.n801 376.045
R9670 VPWR.n806 VPWR.n805 376.045
R9671 VPWR.n810 VPWR.n809 376.045
R9672 VPWR.n814 VPWR.n813 376.045
R9673 VPWR.n818 VPWR.n817 376.045
R9674 VPWR.n822 VPWR.n821 376.045
R9675 VPWR.n826 VPWR.n825 376.045
R9676 VPWR.n830 VPWR.n829 376.045
R9677 VPWR.n790 VPWR.n789 376.045
R9678 VPWR.n1917 VPWR.n1916 376.045
R9679 VPWR.n1919 VPWR.n1918 376.045
R9680 VPWR.n1927 VPWR.n1926 376.045
R9681 VPWR.n1929 VPWR.n1928 376.045
R9682 VPWR.n1939 VPWR.n1938 376.045
R9683 VPWR.n1947 VPWR.n1946 376.045
R9684 VPWR.n1949 VPWR.n1948 376.045
R9685 VPWR.n1957 VPWR.n1956 376.045
R9686 VPWR.n1959 VPWR.n1958 376.045
R9687 VPWR.n1967 VPWR.n1966 376.045
R9688 VPWR.n1969 VPWR.n1968 376.045
R9689 VPWR.n1977 VPWR.n1976 376.045
R9690 VPWR.n1979 VPWR.n1978 376.045
R9691 VPWR.n1987 VPWR.n1986 376.045
R9692 VPWR.n1937 VPWR.n1936 376.045
R9693 VPWR.n927 VPWR.n926 376.045
R9694 VPWR.n925 VPWR.n924 376.045
R9695 VPWR.n921 VPWR.n920 376.045
R9696 VPWR.n917 VPWR.n916 376.045
R9697 VPWR.n909 VPWR.n908 376.045
R9698 VPWR.n905 VPWR.n904 376.045
R9699 VPWR.n901 VPWR.n900 376.045
R9700 VPWR.n897 VPWR.n896 376.045
R9701 VPWR.n893 VPWR.n892 376.045
R9702 VPWR.n889 VPWR.n888 376.045
R9703 VPWR.n885 VPWR.n884 376.045
R9704 VPWR.n881 VPWR.n880 376.045
R9705 VPWR.n877 VPWR.n876 376.045
R9706 VPWR.n873 VPWR.n872 376.045
R9707 VPWR.n913 VPWR.n912 376.045
R9708 VPWR.n1870 VPWR.n1869 376.045
R9709 VPWR.n982 VPWR.n981 376.045
R9710 VPWR.n1494 VPWR.n1493 376.045
R9711 VPWR.n1221 VPWR.n1220 376.045
R9712 VPWR.n402 VPWR.n401 376.045
R9713 VPWR.n2466 VPWR.n2465 376.045
R9714 VPWR.n341 VPWR.n340 376.045
R9715 VPWR.n2520 VPWR.n2519 376.045
R9716 VPWR.n978 VPWR.n977 376.045
R9717 VPWR.n1492 VPWR.n1491 376.045
R9718 VPWR.n1185 VPWR.n1184 376.045
R9719 VPWR.n1868 VPWR.n1867 376.045
R9720 VPWR.n986 VPWR.n985 376.045
R9721 VPWR.n1506 VPWR.n1505 376.045
R9722 VPWR.n1219 VPWR.n1218 376.045
R9723 VPWR.n410 VPWR.n409 376.045
R9724 VPWR.n418 VPWR.n417 376.045
R9725 VPWR.n422 VPWR.n421 376.045
R9726 VPWR.n426 VPWR.n425 376.045
R9727 VPWR.n430 VPWR.n429 376.045
R9728 VPWR.n434 VPWR.n433 376.045
R9729 VPWR.n438 VPWR.n437 376.045
R9730 VPWR.n442 VPWR.n441 376.045
R9731 VPWR.n446 VPWR.n445 376.045
R9732 VPWR.n414 VPWR.n413 376.045
R9733 VPWR.n2448 VPWR.n2447 376.045
R9734 VPWR.n329 VPWR.n328 376.045
R9735 VPWR.n2542 VPWR.n2541 376.045
R9736 VPWR.n990 VPWR.n989 376.045
R9737 VPWR.n1508 VPWR.n1507 376.045
R9738 VPWR.n1216 VPWR.n1215 376.045
R9739 VPWR.n1860 VPWR.n1859 376.045
R9740 VPWR.n1850 VPWR.n1849 376.045
R9741 VPWR.n1848 VPWR.n1847 376.045
R9742 VPWR.n1840 VPWR.n1839 376.045
R9743 VPWR.n1838 VPWR.n1837 376.045
R9744 VPWR.n1830 VPWR.n1829 376.045
R9745 VPWR.n1828 VPWR.n1827 376.045
R9746 VPWR.n1820 VPWR.n1819 376.045
R9747 VPWR.n1858 VPWR.n1857 376.045
R9748 VPWR.n994 VPWR.n993 376.045
R9749 VPWR.n1520 VPWR.n1519 376.045
R9750 VPWR.n1213 VPWR.n1212 376.045
R9751 VPWR.n2468 VPWR.n2467 376.045
R9752 VPWR.n345 VPWR.n344 376.045
R9753 VPWR.n2518 VPWR.n2517 376.045
R9754 VPWR.n1481 VPWR.n1480 376.045
R9755 VPWR.n1182 VPWR.n1181 376.045
R9756 VPWR.n998 VPWR.n997 376.045
R9757 VPWR.n1522 VPWR.n1521 376.045
R9758 VPWR.n1205 VPWR.n1204 376.045
R9759 VPWR.n2438 VPWR.n2437 376.045
R9760 VPWR.n2428 VPWR.n2427 376.045
R9761 VPWR.n2426 VPWR.n2425 376.045
R9762 VPWR.n2418 VPWR.n2417 376.045
R9763 VPWR.n2416 VPWR.n2415 376.045
R9764 VPWR.n2408 VPWR.n2407 376.045
R9765 VPWR.n2436 VPWR.n2435 376.045
R9766 VPWR.n317 VPWR.n316 376.045
R9767 VPWR.n2556 VPWR.n2555 376.045
R9768 VPWR.n1537 VPWR.n1536 376.045
R9769 VPWR.n1202 VPWR.n1201 376.045
R9770 VPWR.n1002 VPWR.n1001 376.045
R9771 VPWR.n1006 VPWR.n1005 376.045
R9772 VPWR.n1010 VPWR.n1009 376.045
R9773 VPWR.n1014 VPWR.n1013 376.045
R9774 VPWR.n1018 VPWR.n1017 376.045
R9775 VPWR.n1022 VPWR.n1021 376.045
R9776 VPWR.n970 VPWR.n969 376.045
R9777 VPWR.n1475 VPWR.n1474 376.045
R9778 VPWR.n1593 VPWR.n1592 376.045
R9779 VPWR.n313 VPWR.n312 376.045
R9780 VPWR.n2566 VPWR.n2565 376.045
R9781 VPWR.n1199 VPWR.n1198 376.045
R9782 VPWR.n1762 VPWR.n1761 376.045
R9783 VPWR.n1191 VPWR.n1190 376.045
R9784 VPWR.n309 VPWR.n308 376.045
R9785 VPWR.n305 VPWR.n304 376.045
R9786 VPWR.n297 VPWR.n296 376.045
R9787 VPWR.n301 VPWR.n300 376.045
R9788 VPWR.n1741 VPWR.n1740 376.045
R9789 VPWR.n1750 VPWR.n1749 376.045
R9790 VPWR.n1791 VPWR.n1790 376.045
R9791 VPWR.n1760 VPWR.n1759 376.045
R9792 VPWR.n1188 VPWR.n1187 376.045
R9793 VPWR.n2578 VPWR.n2577 376.045
R9794 VPWR.n2580 VPWR.n2579 376.045
R9795 VPWR.n2590 VPWR.n2589 376.045
R9796 VPWR.n1739 VPWR.n1738 376.045
R9797 VPWR.n1339 VPWR.t1312 342.841
R9798 VPWR.n1378 VPWR.t411 342.841
R9799 VPWR.n1415 VPWR.t917 342.841
R9800 VPWR.n2693 VPWR.t645 342.841
R9801 VPWR.n2656 VPWR.t752 342.841
R9802 VPWR.n2599 VPWR.t989 342.841
R9803 VPWR.n1339 VPWR.t55 342.839
R9804 VPWR.n1378 VPWR.t156 342.839
R9805 VPWR.n1415 VPWR.t759 342.839
R9806 VPWR.n2693 VPWR.t928 342.839
R9807 VPWR.n2656 VPWR.t474 342.839
R9808 VPWR.n2599 VPWR.t117 342.839
R9809 VPWR.n2842 VPWR.n2824 339.212
R9810 VPWR.n1306 VPWR.t1120 338.488
R9811 VPWR.n2729 VPWR.t1085 338.488
R9812 VPWR.n1315 VPWR.n1314 327.377
R9813 VPWR.n1308 VPWR.n1307 327.377
R9814 VPWR.n1322 VPWR.n1321 327.377
R9815 VPWR.n1352 VPWR.n1350 327.377
R9816 VPWR.n1345 VPWR.n1343 327.377
R9817 VPWR.n1360 VPWR.n1358 327.377
R9818 VPWR.n1391 VPWR.n1389 327.377
R9819 VPWR.n1384 VPWR.n1382 327.377
R9820 VPWR.n1399 VPWR.n1397 327.377
R9821 VPWR.n1428 VPWR.n1426 327.377
R9822 VPWR.n1421 VPWR.n1419 327.377
R9823 VPWR.n1436 VPWR.n1434 327.377
R9824 VPWR.n1324 VPWR.n1323 327.375
R9825 VPWR.n1352 VPWR.n1351 327.375
R9826 VPWR.n1345 VPWR.n1344 327.375
R9827 VPWR.n1360 VPWR.n1359 327.375
R9828 VPWR.n1391 VPWR.n1390 327.375
R9829 VPWR.n1384 VPWR.n1383 327.375
R9830 VPWR.n1399 VPWR.n1398 327.375
R9831 VPWR.n1428 VPWR.n1427 327.375
R9832 VPWR.n1421 VPWR.n1420 327.375
R9833 VPWR.n1436 VPWR.n1435 327.375
R9834 VPWR.n1 VPWR 325.546
R9835 VPWR.n2667 VPWR.t644 322.262
R9836 VPWR.n2630 VPWR.t473 322.262
R9837 VPWR.n2805 VPWR.n2804 321.642
R9838 VPWR.n2722 VPWR.n2712 320.976
R9839 VPWR.n2716 VPWR.n2715 320.976
R9840 VPWR.n2710 VPWR.n2709 320.976
R9841 VPWR.n2680 VPWR.n2679 320.976
R9842 VPWR.n2686 VPWR.n2675 320.976
R9843 VPWR.n2672 VPWR.n2671 320.976
R9844 VPWR.n2643 VPWR.n2642 320.976
R9845 VPWR.n2649 VPWR.n2638 320.976
R9846 VPWR.n2635 VPWR.n2634 320.976
R9847 VPWR.n2610 VPWR.n2606 320.976
R9848 VPWR.n2614 VPWR.n2613 320.976
R9849 VPWR.n2620 VPWR.n2602 320.976
R9850 VPWR.n2727 VPWR.n2708 320.976
R9851 VPWR.n2680 VPWR.n2678 320.976
R9852 VPWR.n2686 VPWR.n2674 320.976
R9853 VPWR.n2672 VPWR.n2670 320.976
R9854 VPWR.n2643 VPWR.n2641 320.976
R9855 VPWR.n2649 VPWR.n2637 320.976
R9856 VPWR.n2635 VPWR.n2633 320.976
R9857 VPWR.n2610 VPWR.n2605 320.976
R9858 VPWR.n2614 VPWR.n2612 320.976
R9859 VPWR.n2620 VPWR.n2601 320.976
R9860 VPWR.n2801 VPWR 319.627
R9861 VPWR.n6 VPWR.n5 316.245
R9862 VPWR.n1241 VPWR.n1239 316.245
R9863 VPWR.n1264 VPWR.n1262 316.245
R9864 VPWR.n1288 VPWR.n1286 316.245
R9865 VPWR.n2784 VPWR.n2783 316.245
R9866 VPWR.n2764 VPWR.n2763 316.245
R9867 VPWR.n2745 VPWR.n2744 316.245
R9868 VPWR.n1241 VPWR.n1240 316.245
R9869 VPWR.n1264 VPWR.n1263 316.245
R9870 VPWR.n1288 VPWR.n1287 316.245
R9871 VPWR.n2784 VPWR.n2782 316.245
R9872 VPWR.n2764 VPWR.n2762 316.245
R9873 VPWR.n2745 VPWR.n2743 316.245
R9874 VPWR.n2630 VPWR.t738 313.87
R9875 VPWR.n10 VPWR.n4 310.502
R9876 VPWR.n1246 VPWR.n1238 310.502
R9877 VPWR.n1269 VPWR.n1261 310.502
R9878 VPWR.n1293 VPWR.n1285 310.502
R9879 VPWR.n2803 VPWR.n2802 310.502
R9880 VPWR.n2788 VPWR.n2787 310.502
R9881 VPWR.n2768 VPWR.n2767 310.502
R9882 VPWR.n2749 VPWR.n2748 310.502
R9883 VPWR.n1246 VPWR.n1245 310.5
R9884 VPWR.n1269 VPWR.n1268 310.5
R9885 VPWR.n1293 VPWR.n1292 310.5
R9886 VPWR.n2788 VPWR.n2786 310.5
R9887 VPWR.n2768 VPWR.n2766 310.5
R9888 VPWR.n2749 VPWR.n2747 310.5
R9889 VPWR.n2834 VPWR.n2833 279.341
R9890 VPWR.n2839 VPWR.n2838 279.341
R9891 VPWR.n1412 VPWR.t501 255.905
R9892 VPWR.n2663 VPWR.t739 255.905
R9893 VPWR.n1275 VPWR.t744 255.904
R9894 VPWR.n1412 VPWR.t269 255.904
R9895 VPWR.n2774 VPWR.t1101 255.904
R9896 VPWR.n2663 VPWR.t840 255.904
R9897 VPWR.n1303 VPWR.t1201 254.019
R9898 VPWR.n2735 VPWR.t192 254.019
R9899 VPWR.n1335 VPWR.t1199 252.948
R9900 VPWR.n2737 VPWR.t190 252.948
R9901 VPWR.n1373 VPWR.t745 250.722
R9902 VPWR.n2700 VPWR.t1853 250.722
R9903 VPWR.n1310 VPWR.t394 249.901
R9904 VPWR.n1346 VPWR.t939 249.901
R9905 VPWR.n1385 VPWR.t447 249.901
R9906 VPWR.n1422 VPWR.t953 249.901
R9907 VPWR.n2714 VPWR.t273 249.901
R9908 VPWR.n2677 VPWR.t277 249.901
R9909 VPWR.n2640 VPWR.t315 249.901
R9910 VPWR.n2607 VPWR.t298 249.901
R9911 VPWR.n1346 VPWR.t445 249.901
R9912 VPWR.n1385 VPWR.t936 249.901
R9913 VPWR.n1422 VPWR.t950 249.901
R9914 VPWR.n2677 VPWR.t316 249.901
R9915 VPWR.n2640 VPWR.t300 249.901
R9916 VPWR.n2607 VPWR.t252 249.901
R9917 VPWR.n1253 VPWR.t1854 249.363
R9918 VPWR.n1338 VPWR.t746 249.363
R9919 VPWR.n2811 VPWR.t832 249.363
R9920 VPWR.n2795 VPWR.t835 249.363
R9921 VPWR.n2698 VPWR.t136 249.363
R9922 VPWR.n17 VPWR.t552 249.362
R9923 VPWR.n1253 VPWR.t80 249.362
R9924 VPWR.n2795 VPWR.t46 249.362
R9925 VPWR.t740 VPWR.t551 248.599
R9926 VPWR.t1117 VPWR.t981 248.599
R9927 VPWR.t981 VPWR.t985 248.599
R9928 VPWR.t985 VPWR.t1194 248.599
R9929 VPWR.t1194 VPWR.t329 248.599
R9930 VPWR.t329 VPWR.t332 248.599
R9931 VPWR.t332 VPWR.t938 248.599
R9932 VPWR.t938 VPWR.t955 248.599
R9933 VPWR.t232 VPWR.t443 248.599
R9934 VPWR.t443 VPWR.t393 248.599
R9935 VPWR.t313 VPWR.t247 248.599
R9936 VPWR.t326 VPWR.t313 248.599
R9937 VPWR.t213 VPWR.t326 248.599
R9938 VPWR.t1086 VPWR.t213 248.599
R9939 VPWR.t1080 VPWR.t1086 248.599
R9940 VPWR.t1092 VPWR.t1080 248.599
R9941 VPWR.t1094 VPWR.t1092 248.599
R9942 VPWR.t1102 VPWR.t831 248.599
R9943 VPWR.t223 VPWR.t272 248.599
R9944 VPWR.t1833 VPWR.t223 248.599
R9945 VPWR.n15 VPWR.t741 247.394
R9946 VPWR.n1251 VPWR.t743 247.394
R9947 VPWR.n2809 VPWR.t1103 247.394
R9948 VPWR.n2793 VPWR.t1097 247.394
R9949 VPWR.n1251 VPWR.t742 247.394
R9950 VPWR.n2793 VPWR.t1099 247.394
R9951 VPWR.n1304 VPWR.t397 244.737
R9952 VPWR.n2730 VPWR.t312 244.737
R9953 VPWR.n1374 VPWR.t160 243.886
R9954 VPWR.n2701 VPWR.t1234 243.886
R9955 VPWR.n1277 VPWR.t550 243.512
R9956 VPWR.n1300 VPWR.t1855 243.512
R9957 VPWR.n1303 VPWR.t748 243.512
R9958 VPWR.n2776 VPWR.t834 243.512
R9959 VPWR.n2756 VPWR.t836 243.512
R9960 VPWR.n2735 VPWR.t134 243.512
R9961 VPWR.n1300 VPWR.t82 243.512
R9962 VPWR.n2756 VPWR.t44 243.512
R9963 VPWR.n1329 VPWR.t1200 238.339
R9964 VPWR.n2705 VPWR.t191 238.339
R9965 VPWR.n2855 VPWR.t193 237.99
R9966 VPWR.n2667 VPWR.t135 234.982
R9967 VPWR.t230 VPWR.t232 228.101
R9968 VPWR.t322 VPWR.t1833 228.101
R9969 VPWR.n2801 VPWR 224.923
R9970 VPWR.n1 VPWR 219.004
R9971 VPWR.n1444 VPWR.n1443 214.613
R9972 VPWR.n1444 VPWR.n1442 214.613
R9973 VPWR.n1236 VPWR.n1235 214.326
R9974 VPWR.n1259 VPWR.n1258 214.326
R9975 VPWR.n1283 VPWR.n1282 214.326
R9976 VPWR.n1368 VPWR.n1367 214.326
R9977 VPWR.n1407 VPWR.n1406 214.326
R9978 VPWR.n1236 VPWR.n1234 214.326
R9979 VPWR.n1259 VPWR.n1257 214.326
R9980 VPWR.n1283 VPWR.n1281 214.326
R9981 VPWR.n1368 VPWR.n1366 214.326
R9982 VPWR.n1407 VPWR.n1405 214.326
R9983 VPWR.n2 VPWR.n1 213.119
R9984 VPWR.n2808 VPWR.n2801 213.119
R9985 VPWR VPWR.t740 207.166
R9986 VPWR.n2840 VPWR.n2839 204.424
R9987 VPWR.n2830 VPWR.n2817 204.424
R9988 VPWR.n2833 VPWR.n2820 204.424
R9989 VPWR.n2844 VPWR.n2841 204.048
R9990 VPWR VPWR.t1094 201.246
R9991 VPWR.t393 VPWR 189.409
R9992 VPWR.n2741 VPWR 184.63
R9993 VPWR.n1329 VPWR 182.952
R9994 VPWR.n2760 VPWR 182.952
R9995 VPWR.n2780 VPWR 181.273
R9996 VPWR.t738 VPWR 177.916
R9997 VPWR.n2848 VPWR.n2847 166.4
R9998 VPWR.n1770 VPWR.n1768 161.365
R9999 VPWR.n1041 VPWR.n1039 161.365
R10000 VPWR.n1545 VPWR.n1543 161.365
R10001 VPWR.n1550 VPWR.n1548 161.365
R10002 VPWR.n1555 VPWR.n1553 161.365
R10003 VPWR.n1560 VPWR.n1558 161.365
R10004 VPWR.n1565 VPWR.n1563 161.365
R10005 VPWR.n1570 VPWR.n1568 161.365
R10006 VPWR.n1575 VPWR.n1573 161.365
R10007 VPWR.n1580 VPWR.n1578 161.365
R10008 VPWR.n1135 VPWR.n1133 161.365
R10009 VPWR.n1460 VPWR.n1458 161.365
R10010 VPWR.n1455 VPWR.n1453 161.365
R10011 VPWR.n1775 VPWR.n1773 161.365
R10012 VPWR.n1783 VPWR.n1781 161.365
R10013 VPWR.n1779 VPWR.n1777 161.365
R10014 VPWR VPWR.n53 161.363
R10015 VPWR VPWR.n51 161.363
R10016 VPWR VPWR.n49 161.363
R10017 VPWR VPWR.n47 161.363
R10018 VPWR VPWR.n45 161.363
R10019 VPWR VPWR.n43 161.363
R10020 VPWR VPWR.n41 161.363
R10021 VPWR VPWR.n39 161.363
R10022 VPWR VPWR.n37 161.363
R10023 VPWR VPWR.n35 161.363
R10024 VPWR VPWR.n33 161.363
R10025 VPWR VPWR.n31 161.363
R10026 VPWR VPWR.n29 161.363
R10027 VPWR VPWR.n27 161.363
R10028 VPWR VPWR.n25 161.363
R10029 VPWR VPWR.n23 161.363
R10030 VPWR.n1115 VPWR.n1114 161.303
R10031 VPWR.n107 VPWR.n106 161.303
R10032 VPWR.n1120 VPWR.n1119 161.3
R10033 VPWR.n1599 VPWR.n1598 161.3
R10034 VPWR.n1602 VPWR.n1601 161.3
R10035 VPWR.n1111 VPWR.n1110 161.3
R10036 VPWR.n1126 VPWR.n1125 161.3
R10037 VPWR.n1107 VPWR.n1106 161.3
R10038 VPWR.n1612 VPWR.n1611 161.3
R10039 VPWR.n1615 VPWR.n1614 161.3
R10040 VPWR.n1618 VPWR.n1617 161.3
R10041 VPWR.n1623 VPWR.n1622 161.3
R10042 VPWR.n1626 VPWR.n1625 161.3
R10043 VPWR.n1629 VPWR.n1628 161.3
R10044 VPWR.n1101 VPWR.n1100 161.3
R10045 VPWR.n1177 VPWR.n1176 161.3
R10046 VPWR.n1097 VPWR.n1096 161.3
R10047 VPWR.n1639 VPWR.n1638 161.3
R10048 VPWR.n1642 VPWR.n1641 161.3
R10049 VPWR.n1645 VPWR.n1644 161.3
R10050 VPWR.n1650 VPWR.n1649 161.3
R10051 VPWR.n1653 VPWR.n1652 161.3
R10052 VPWR.n1656 VPWR.n1655 161.3
R10053 VPWR.n1091 VPWR.n1090 161.3
R10054 VPWR.n1209 VPWR.n1208 161.3
R10055 VPWR.n1087 VPWR.n1086 161.3
R10056 VPWR.n1666 VPWR.n1665 161.3
R10057 VPWR.n1669 VPWR.n1668 161.3
R10058 VPWR.n1672 VPWR.n1671 161.3
R10059 VPWR.n1677 VPWR.n1676 161.3
R10060 VPWR.n1680 VPWR.n1679 161.3
R10061 VPWR.n1683 VPWR.n1682 161.3
R10062 VPWR.n1081 VPWR.n1080 161.3
R10063 VPWR.n1195 VPWR.n1194 161.3
R10064 VPWR.n1077 VPWR.n1076 161.3
R10065 VPWR.n1693 VPWR.n1692 161.3
R10066 VPWR.n1696 VPWR.n1695 161.3
R10067 VPWR.n1699 VPWR.n1698 161.3
R10068 VPWR.n1704 VPWR.n1703 161.3
R10069 VPWR.n1707 VPWR.n1706 161.3
R10070 VPWR.n1710 VPWR.n1709 161.3
R10071 VPWR.n1070 VPWR.n1069 161.3
R10072 VPWR.n1719 VPWR.n1718 161.3
R10073 VPWR.n1722 VPWR.n1721 161.3
R10074 VPWR.n1717 VPWR.n1716 161.3
R10075 VPWR.n1734 VPWR.n1733 161.3
R10076 VPWR.n1117 VPWR.n1116 161.3
R10077 VPWR.n1731 VPWR.n1730 161.3
R10078 VPWR.n1065 VPWR.n1064 161.3
R10079 VPWR.n126 VPWR.n125 161.3
R10080 VPWR.n117 VPWR.n116 161.3
R10081 VPWR.n120 VPWR.n119 161.3
R10082 VPWR.n115 VPWR.n114 161.3
R10083 VPWR.n138 VPWR.n137 161.3
R10084 VPWR.n128 VPWR.n127 161.3
R10085 VPWR.n109 VPWR.n108 161.3
R10086 VPWR.n105 VPWR.n104 161.3
R10087 VPWR.n288 VPWR.n287 161.3
R10088 VPWR.n285 VPWR.n284 161.3
R10089 VPWR.n101 VPWR.n100 161.3
R10090 VPWR.n272 VPWR.n271 161.3
R10091 VPWR.n275 VPWR.n274 161.3
R10092 VPWR.n270 VPWR.n269 161.3
R10093 VPWR.n260 VPWR.n259 161.3
R10094 VPWR.n263 VPWR.n262 161.3
R10095 VPWR.n258 VPWR.n257 161.3
R10096 VPWR.n248 VPWR.n247 161.3
R10097 VPWR.n251 VPWR.n250 161.3
R10098 VPWR.n246 VPWR.n245 161.3
R10099 VPWR.n236 VPWR.n235 161.3
R10100 VPWR.n239 VPWR.n238 161.3
R10101 VPWR.n234 VPWR.n233 161.3
R10102 VPWR.n224 VPWR.n223 161.3
R10103 VPWR.n227 VPWR.n226 161.3
R10104 VPWR.n222 VPWR.n221 161.3
R10105 VPWR.n212 VPWR.n211 161.3
R10106 VPWR.n215 VPWR.n214 161.3
R10107 VPWR.n210 VPWR.n209 161.3
R10108 VPWR.n200 VPWR.n199 161.3
R10109 VPWR.n203 VPWR.n202 161.3
R10110 VPWR.n198 VPWR.n197 161.3
R10111 VPWR.n188 VPWR.n187 161.3
R10112 VPWR.n191 VPWR.n190 161.3
R10113 VPWR.n186 VPWR.n185 161.3
R10114 VPWR.n176 VPWR.n175 161.3
R10115 VPWR.n179 VPWR.n178 161.3
R10116 VPWR.n174 VPWR.n173 161.3
R10117 VPWR.n164 VPWR.n163 161.3
R10118 VPWR.n167 VPWR.n166 161.3
R10119 VPWR.n162 VPWR.n161 161.3
R10120 VPWR.n152 VPWR.n151 161.3
R10121 VPWR.n155 VPWR.n154 161.3
R10122 VPWR.n150 VPWR.n149 161.3
R10123 VPWR.n140 VPWR.n139 161.3
R10124 VPWR.n143 VPWR.n142 161.3
R10125 VPWR.n131 VPWR.n130 161.3
R10126 VPWR.n1601 VPWR.t1386 161.202
R10127 VPWR.n1106 VPWR.t1511 161.202
R10128 VPWR.n1617 VPWR.t1552 161.202
R10129 VPWR.n1628 VPWR.t1660 161.202
R10130 VPWR.n1096 VPWR.t1427 161.202
R10131 VPWR.n1644 VPWR.t1442 161.202
R10132 VPWR.n1655 VPWR.t1665 161.202
R10133 VPWR.n1086 VPWR.t1708 161.202
R10134 VPWR.n1671 VPWR.t1425 161.202
R10135 VPWR.n1682 VPWR.t1578 161.202
R10136 VPWR.n1076 VPWR.t1600 161.202
R10137 VPWR.n1698 VPWR.t1450 161.202
R10138 VPWR.n1709 VPWR.t1476 161.202
R10139 VPWR.n1721 VPWR.t1501 161.202
R10140 VPWR.n1116 VPWR.t1641 161.202
R10141 VPWR.n1730 VPWR.t1346 161.202
R10142 VPWR.n119 VPWR.t1468 161.202
R10143 VPWR.n108 VPWR.t1367 161.202
R10144 VPWR.n284 VPWR.t1503 161.202
R10145 VPWR.n274 VPWR.t1633 161.202
R10146 VPWR.n262 VPWR.t1673 161.202
R10147 VPWR.n250 VPWR.t1397 161.202
R10148 VPWR.n238 VPWR.t1541 161.202
R10149 VPWR.n226 VPWR.t1565 161.202
R10150 VPWR.n214 VPWR.t1402 161.202
R10151 VPWR.n202 VPWR.t1437 161.202
R10152 VPWR.n190 VPWR.t1539 161.202
R10153 VPWR.n178 VPWR.t1700 161.202
R10154 VPWR.n166 VPWR.t1719 161.202
R10155 VPWR.n154 VPWR.t1573 161.202
R10156 VPWR.n1768 VPWR.t1625 161.202
R10157 VPWR.n1039 VPWR.t1381 161.202
R10158 VPWR.n1543 VPWR.t1362 161.202
R10159 VPWR.n1548 VPWR.t1611 161.202
R10160 VPWR.n1553 VPWR.t1493 161.202
R10161 VPWR.n1558 VPWR.t1463 161.202
R10162 VPWR.n1563 VPWR.t1615 161.202
R10163 VPWR.n1568 VPWR.t1613 161.202
R10164 VPWR.n1573 VPWR.t1458 161.202
R10165 VPWR.n1578 VPWR.t1348 161.202
R10166 VPWR.n1133 VPWR.t1692 161.202
R10167 VPWR.n1458 VPWR.t1563 161.202
R10168 VPWR.n1453 VPWR.t1432 161.202
R10169 VPWR.n1773 VPWR.t1643 161.202
R10170 VPWR.n1781 VPWR.t1681 161.202
R10171 VPWR.n1777 VPWR.t1513 161.202
R10172 VPWR.n142 VPWR.t1592 161.202
R10173 VPWR.n130 VPWR.t1617 161.202
R10174 VPWR.n1119 VPWR.t1369 161.106
R10175 VPWR.n1110 VPWR.t1505 161.106
R10176 VPWR.n1611 VPWR.t1518 161.106
R10177 VPWR.n1622 VPWR.t1678 161.106
R10178 VPWR.n1100 VPWR.t1399 161.106
R10179 VPWR.n1638 VPWR.t1546 161.106
R10180 VPWR.n1649 VPWR.t1654 161.106
R10181 VPWR.n1090 VPWR.t1694 161.106
R10182 VPWR.n1665 VPWR.t1439 161.106
R10183 VPWR.n1676 VPWR.t1543 161.106
R10184 VPWR.n1080 VPWR.t1702 161.106
R10185 VPWR.n1692 VPWR.t1721 161.106
R10186 VPWR.n1703 VPWR.t1465 161.106
R10187 VPWR.n1069 VPWR.t1594 161.106
R10188 VPWR.n1716 VPWR.t1622 161.106
R10189 VPWR.n1064 VPWR.t1473 161.106
R10190 VPWR.n125 VPWR.t1353 161.106
R10191 VPWR.n114 VPWR.t1589 161.106
R10192 VPWR.n137 VPWR.t1713 161.106
R10193 VPWR.n104 VPWR.t1498 161.106
R10194 VPWR.n100 VPWR.t1627 161.106
R10195 VPWR.n269 VPWR.t1645 161.106
R10196 VPWR.n257 VPWR.t1407 161.106
R10197 VPWR.n245 VPWR.t1515 161.106
R10198 VPWR.n233 VPWR.t1670 161.106
R10199 VPWR.n221 VPWR.t1394 161.106
R10200 VPWR.n209 VPWR.t1429 161.106
R10201 VPWR.n197 VPWR.t1557 161.106
R10202 VPWR.n185 VPWR.t1667 161.106
R10203 VPWR.n173 VPWR.t1434 161.106
R10204 VPWR.n161 VPWR.t1452 161.106
R10205 VPWR.n149 VPWR.t1580 161.106
R10206 VPWR.n53 VPWR.t1697 161.106
R10207 VPWR.n51 VPWR.t1657 161.106
R10208 VPWR.n49 VPWR.t1375 161.106
R10209 VPWR.n47 VPWR.t1487 161.106
R10210 VPWR.n45 VPWR.t1705 161.106
R10211 VPWR.n43 VPWR.t1554 161.106
R10212 VPWR.n41 VPWR.t1662 161.106
R10213 VPWR.n39 VPWR.t1388 161.106
R10214 VPWR.n37 VPWR.t1495 161.106
R10215 VPWR.n35 VPWR.t1455 161.106
R10216 VPWR.n33 VPWR.t1560 161.106
R10217 VPWR.n31 VPWR.t1383 161.106
R10218 VPWR.n29 VPWR.t1567 161.106
R10219 VPWR.n27 VPWR.t1675 161.106
R10220 VPWR.n25 VPWR.t1527 161.106
R10221 VPWR.n23 VPWR.t1638 161.106
R10222 VPWR.n1598 VPWR.t1419 159.978
R10223 VPWR.n1125 VPWR.t1521 159.978
R10224 VPWR.n1614 VPWR.t1686 159.978
R10225 VPWR.n1625 VPWR.t1404 159.978
R10226 VPWR.n1176 VPWR.t1416 159.978
R10227 VPWR.n1641 VPWR.t1575 159.978
R10228 VPWR.n1652 VPWR.t1683 159.978
R10229 VPWR.n1208 VPWR.t1444 159.978
R10230 VPWR.n1668 VPWR.t1470 159.978
R10231 VPWR.n1679 VPWR.t1597 159.978
R10232 VPWR.n1194 VPWR.t1343 159.978
R10233 VPWR.n1695 VPWR.t1364 159.978
R10234 VPWR.n1706 VPWR.t1602 159.978
R10235 VPWR.n1718 VPWR.t1630 159.978
R10236 VPWR.n1733 VPWR.t1350 159.978
R10237 VPWR.n1114 VPWR.t1651 159.978
R10238 VPWR.n116 VPWR.t1484 159.978
R10239 VPWR.n127 VPWR.t1359 159.978
R10240 VPWR.n106 VPWR.t1391 159.978
R10241 VPWR.n287 VPWR.t1536 159.978
R10242 VPWR.n271 VPWR.t1648 159.978
R10243 VPWR.n259 VPWR.t1413 159.978
R10244 VPWR.n247 VPWR.t1524 159.978
R10245 VPWR.n235 VPWR.t1533 159.978
R10246 VPWR.n223 VPWR.t1689 159.978
R10247 VPWR.n211 VPWR.t1410 159.978
R10248 VPWR.n199 VPWR.t1570 159.978
R10249 VPWR.n187 VPWR.t1586 159.978
R10250 VPWR.n175 VPWR.t1716 159.978
R10251 VPWR.n163 VPWR.t1460 159.978
R10252 VPWR.n151 VPWR.t1490 159.978
R10253 VPWR.n1228 VPWR.t1447 159.978
R10254 VPWR.n1150 VPWR.t1378 159.978
R10255 VPWR.n1224 VPWR.t1583 159.978
R10256 VPWR.n1482 VPWR.t1481 159.978
R10257 VPWR.n1170 VPWR.t1605 159.978
R10258 VPWR.n1166 VPWR.t1356 159.978
R10259 VPWR.n1160 VPWR.t1478 159.978
R10260 VPWR.n1476 VPWR.t1710 159.978
R10261 VPWR.n1156 VPWR.t1619 159.978
R10262 VPWR.n1146 VPWR.t1635 159.978
R10263 VPWR.n1469 VPWR.t1608 159.978
R10264 VPWR.n1046 VPWR.t1508 159.978
R10265 VPWR.n1745 VPWR.t1372 159.978
R10266 VPWR.n1033 VPWR.t1422 159.978
R10267 VPWR.n1029 VPWR.t1530 159.978
R10268 VPWR.n1050 VPWR.t1549 159.978
R10269 VPWR.n139 VPWR.t1340 159.978
R10270 VPWR.n1229 VPWR.n1228 152
R10271 VPWR.n1151 VPWR.n1150 152
R10272 VPWR.n1225 VPWR.n1224 152
R10273 VPWR.n1483 VPWR.n1482 152
R10274 VPWR.n1171 VPWR.n1170 152
R10275 VPWR.n1167 VPWR.n1166 152
R10276 VPWR.n1161 VPWR.n1160 152
R10277 VPWR.n1477 VPWR.n1476 152
R10278 VPWR.n1157 VPWR.n1156 152
R10279 VPWR.n1147 VPWR.n1146 152
R10280 VPWR.n1470 VPWR.n1469 152
R10281 VPWR.n1047 VPWR.n1046 152
R10282 VPWR.n1746 VPWR.n1745 152
R10283 VPWR.n1034 VPWR.n1033 152
R10284 VPWR.n1030 VPWR.n1029 152
R10285 VPWR.n1051 VPWR.n1050 152
R10286 VPWR.n2845 VPWR.n2844 150.213
R10287 VPWR.n1601 VPWR.t2063 145.137
R10288 VPWR.n1106 VPWR.t2014 145.137
R10289 VPWR.n1617 VPWR.t2000 145.137
R10290 VPWR.n1628 VPWR.t1962 145.137
R10291 VPWR.n1096 VPWR.t2049 145.137
R10292 VPWR.n1644 VPWR.t2042 145.137
R10293 VPWR.n1655 VPWR.t1959 145.137
R10294 VPWR.n1086 VPWR.t1945 145.137
R10295 VPWR.n1671 VPWR.t2050 145.137
R10296 VPWR.n1682 VPWR.t1993 145.137
R10297 VPWR.n1076 VPWR.t1988 145.137
R10298 VPWR.n1698 VPWR.t2040 145.137
R10299 VPWR.n1709 VPWR.t2033 145.137
R10300 VPWR.n1721 VPWR.t2019 145.137
R10301 VPWR.n1116 VPWR.t1969 145.137
R10302 VPWR.n1730 VPWR.t1937 145.137
R10303 VPWR.n119 VPWR.t2048 145.137
R10304 VPWR.n108 VPWR.t1934 145.137
R10305 VPWR.n284 VPWR.t2030 145.137
R10306 VPWR.n274 VPWR.t1983 145.137
R10307 VPWR.n262 VPWR.t1971 145.137
R10308 VPWR.n250 VPWR.t1930 145.137
R10309 VPWR.n238 VPWR.t2016 145.137
R10310 VPWR.n226 VPWR.t2008 145.137
R10311 VPWR.n214 VPWR.t1928 145.137
R10312 VPWR.n202 VPWR.t2057 145.137
R10313 VPWR.n190 VPWR.t2017 145.137
R10314 VPWR.n178 VPWR.t1961 145.137
R10315 VPWR.n166 VPWR.t1952 145.137
R10316 VPWR.n154 VPWR.t2007 145.137
R10317 VPWR.n1768 VPWR.t1976 145.137
R10318 VPWR.n1039 VPWR.t2065 145.137
R10319 VPWR.n1543 VPWR.t1929 145.137
R10320 VPWR.n1548 VPWR.t1986 145.137
R10321 VPWR.n1553 VPWR.t2025 145.137
R10322 VPWR.n1558 VPWR.t2037 145.137
R10323 VPWR.n1563 VPWR.t1979 145.137
R10324 VPWR.n1568 VPWR.t1985 145.137
R10325 VPWR.n1573 VPWR.t2039 145.137
R10326 VPWR.n1578 VPWR.t1936 145.137
R10327 VPWR.n1133 VPWR.t1950 145.137
R10328 VPWR.n1458 VPWR.t1996 145.137
R10329 VPWR.n1453 VPWR.t2045 145.137
R10330 VPWR.n1773 VPWR.t1968 145.137
R10331 VPWR.n1781 VPWR.t1953 145.137
R10332 VPWR.n1777 VPWR.t2013 145.137
R10333 VPWR.n142 VPWR.t1999 145.137
R10334 VPWR.n130 VPWR.t1990 145.137
R10335 VPWR.n1119 VPWR.t2067 145.038
R10336 VPWR.n1110 VPWR.t2018 145.038
R10337 VPWR.n1611 VPWR.t2010 145.038
R10338 VPWR.n1622 VPWR.t1955 145.038
R10339 VPWR.n1100 VPWR.t2059 145.038
R10340 VPWR.n1638 VPWR.t2002 145.038
R10341 VPWR.n1649 VPWR.t1964 145.038
R10342 VPWR.n1090 VPWR.t1949 145.038
R10343 VPWR.n1665 VPWR.t2043 145.038
R10344 VPWR.n1676 VPWR.t2003 145.038
R10345 VPWR.n1080 VPWR.t1947 145.038
R10346 VPWR.n1692 VPWR.t1939 145.038
R10347 VPWR.n1703 VPWR.t2036 145.038
R10348 VPWR.n1069 VPWR.t1989 145.038
R10349 VPWR.n1716 VPWR.t1977 145.038
R10350 VPWR.n1064 VPWR.t2034 145.038
R10351 VPWR.n125 VPWR.t1940 145.038
R10352 VPWR.n114 VPWR.t2001 145.038
R10353 VPWR.n137 VPWR.t1954 145.038
R10354 VPWR.n104 VPWR.t2032 145.038
R10355 VPWR.n100 VPWR.t1987 145.038
R10356 VPWR.n269 VPWR.t1980 145.038
R10357 VPWR.n257 VPWR.t2068 145.038
R10358 VPWR.n245 VPWR.t2027 145.038
R10359 VPWR.n233 VPWR.t1972 145.038
R10360 VPWR.n221 VPWR.t1931 145.038
R10361 VPWR.n209 VPWR.t2060 145.038
R10362 VPWR.n197 VPWR.t2009 145.038
R10363 VPWR.n185 VPWR.t1973 145.038
R10364 VPWR.n173 VPWR.t2058 145.038
R10365 VPWR.n161 VPWR.t2052 145.038
R10366 VPWR.n149 VPWR.t2004 145.038
R10367 VPWR.n53 VPWR.t2053 145.038
R10368 VPWR.n51 VPWR.t1963 145.038
R10369 VPWR.n49 VPWR.t2066 145.038
R10370 VPWR.n47 VPWR.t2026 145.038
R10371 VPWR.n45 VPWR.t1946 145.038
R10372 VPWR.n43 VPWR.t2051 145.038
R10373 VPWR.n41 VPWR.t2069 145.038
R10374 VPWR.n39 VPWR.t2028 145.038
R10375 VPWR.n37 VPWR.t2022 145.038
R10376 VPWR.n35 VPWR.t1943 145.038
R10377 VPWR.n33 VPWR.t1997 145.038
R10378 VPWR.n31 VPWR.t2064 145.038
R10379 VPWR.n29 VPWR.t1995 145.038
R10380 VPWR.n27 VPWR.t1956 145.038
R10381 VPWR.n25 VPWR.t2021 145.038
R10382 VPWR.n23 VPWR.t1970 145.038
R10383 VPWR.n1598 VPWR.t1966 143.911
R10384 VPWR.n1125 VPWR.t2062 143.911
R10385 VPWR.n1614 VPWR.t2047 143.911
R10386 VPWR.n1625 VPWR.t1965 143.911
R10387 VPWR.n1176 VPWR.t1958 143.911
R10388 VPWR.n1641 VPWR.t1944 143.911
R10389 VPWR.n1652 VPWR.t2005 143.911
R10390 VPWR.n1208 VPWR.t1992 143.911
R10391 VPWR.n1668 VPWR.t1941 143.911
R10392 VPWR.n1679 VPWR.t2038 143.911
R10393 VPWR.n1194 VPWR.t2031 143.911
R10394 VPWR.n1695 VPWR.t1978 143.911
R10395 VPWR.n1706 VPWR.t1935 143.911
R10396 VPWR.n1718 VPWR.t2024 143.911
R10397 VPWR.n1733 VPWR.t1984 143.911
R10398 VPWR.n1114 VPWR.t2012 143.911
R10399 VPWR.n116 VPWR.t1951 143.911
R10400 VPWR.n127 VPWR.t1991 143.911
R10401 VPWR.n106 VPWR.t1981 143.911
R10402 VPWR.n287 VPWR.t1933 143.911
R10403 VPWR.n271 VPWR.t2029 143.911
R10404 VPWR.n259 VPWR.t2015 143.911
R10405 VPWR.n247 VPWR.t1932 143.911
R10406 VPWR.n235 VPWR.t1926 143.911
R10407 VPWR.n223 VPWR.t2056 143.911
R10408 VPWR.n211 VPWR.t1974 143.911
R10409 VPWR.n199 VPWR.t1960 143.911
R10410 VPWR.n187 VPWR.t2054 143.911
R10411 VPWR.n175 VPWR.t2006 143.911
R10412 VPWR.n163 VPWR.t1998 143.911
R10413 VPWR.n151 VPWR.t1942 143.911
R10414 VPWR.n1228 VPWR.t1948 143.911
R10415 VPWR.n1150 VPWR.t1975 143.911
R10416 VPWR.n1224 VPWR.t2041 143.911
R10417 VPWR.n1482 VPWR.t1982 143.911
R10418 VPWR.n1170 VPWR.t2035 143.911
R10419 VPWR.n1166 VPWR.t2023 143.911
R10420 VPWR.n1160 VPWR.t1938 143.911
R10421 VPWR.n1476 VPWR.t1994 143.911
R10422 VPWR.n1156 VPWR.t1927 143.911
R10423 VPWR.n1146 VPWR.t2020 143.911
R10424 VPWR.n1469 VPWR.t2044 143.911
R10425 VPWR.n1046 VPWR.t1967 143.911
R10426 VPWR.n1745 VPWR.t2011 143.911
R10427 VPWR.n1033 VPWR.t1957 143.911
R10428 VPWR.n1029 VPWR.t2061 143.911
R10429 VPWR.n1050 VPWR.t2055 143.911
R10430 VPWR.n139 VPWR.t2046 143.911
R10431 VPWR.t1192 VPWR.t230 140.989
R10432 VPWR.t250 VPWR.t225 140.989
R10433 VPWR.t278 VPWR.t250 140.989
R10434 VPWR.t241 VPWR.t278 140.989
R10435 VPWR.t652 VPWR.t241 140.989
R10436 VPWR.t646 VPWR.t652 140.989
R10437 VPWR.t638 VPWR.t646 140.989
R10438 VPWR.t640 VPWR.t638 140.989
R10439 VPWR.t1096 VPWR.t45 140.989
R10440 VPWR.t1832 VPWR.t237 140.989
R10441 VPWR.t301 VPWR.t1832 140.989
R10442 VPWR.t1831 VPWR.t301 140.989
R10443 VPWR.t465 VPWR.t1831 140.989
R10444 VPWR.t475 VPWR.t465 140.989
R10445 VPWR.t467 VPWR.t475 140.989
R10446 VPWR.t469 VPWR.t467 140.989
R10447 VPWR.t228 VPWR.t279 140.989
R10448 VPWR.t321 VPWR.t228 140.989
R10449 VPWR.t222 VPWR.t321 140.989
R10450 VPWR.t124 VPWR.t222 140.989
R10451 VPWR.t118 VPWR.t124 140.989
R10452 VPWR.t126 VPWR.t118 140.989
R10453 VPWR.t128 VPWR.t126 140.989
R10454 VPWR.t1088 VPWR.t322 140.989
R10455 VPWR.t226 VPWR.t276 140.989
R10456 VPWR.t309 VPWR.t226 140.989
R10457 VPWR.t274 VPWR.t309 140.989
R10458 VPWR.t648 VPWR.t274 140.989
R10459 VPWR.t642 VPWR.t648 140.989
R10460 VPWR.t650 VPWR.t642 140.989
R10461 VPWR.t644 VPWR.t650 140.989
R10462 VPWR.t235 VPWR.t299 140.989
R10463 VPWR.t214 VPWR.t235 140.989
R10464 VPWR.t270 VPWR.t214 140.989
R10465 VPWR.t461 VPWR.t270 140.989
R10466 VPWR.t471 VPWR.t461 140.989
R10467 VPWR.t463 VPWR.t471 140.989
R10468 VPWR.t473 VPWR.t463 140.989
R10469 VPWR.t239 VPWR.t251 140.989
R10470 VPWR.t245 VPWR.t239 140.989
R10471 VPWR.t253 VPWR.t245 140.989
R10472 VPWR.t120 VPWR.t253 140.989
R10473 VPWR.t114 VPWR.t120 140.989
R10474 VPWR.t122 VPWR.t114 140.989
R10475 VPWR.t116 VPWR.t122 140.989
R10476 VPWR VPWR.n1442 133.312
R10477 VPWR.n2841 VPWR.n2840 129.13
R10478 VPWR.n2858 VPWR.n2819 129.13
R10479 VPWR.n2780 VPWR 127.562
R10480 VPWR.n2760 VPWR 127.562
R10481 VPWR.n2741 VPWR 127.562
R10482 VPWR VPWR.t311 125.883
R10483 VPWR.n2705 VPWR 125.883
R10484 VPWR.t1098 VPWR.t43 120.849
R10485 VPWR.t747 VPWR.t1198 117.492
R10486 VPWR.t133 VPWR.t189 117.492
R10487 VPWR.t1233 VPWR 115.814
R10488 VPWR VPWR.t640 114.135
R10489 VPWR VPWR.t469 114.135
R10490 VPWR VPWR.t128 114.135
R10491 VPWR.n2859 VPWR.n2817 111.059
R10492 VPWR.t1235 VPWR 107.421
R10493 VPWR.n1330 VPWR.n1329 106.561
R10494 VPWR.n2781 VPWR.n2780 106.561
R10495 VPWR.n2761 VPWR.n2760 106.561
R10496 VPWR.n2742 VPWR.n2741 106.561
R10497 VPWR.n2706 VPWR.n2705 106.561
R10498 VPWR.n2668 VPWR.n2667 106.561
R10499 VPWR.n2631 VPWR.n2630 106.561
R10500 VPWR VPWR.t1102 106.543
R10501 VPWR VPWR.n1234 104.8
R10502 VPWR VPWR.n1257 104.8
R10503 VPWR VPWR.n1281 104.8
R10504 VPWR VPWR.n1366 104.8
R10505 VPWR VPWR.n1405 104.8
R10506 VPWR.n1443 VPWR 100.883
R10507 VPWR VPWR.t1117 100.624
R10508 VPWR.t693 VPWR.t193 97.9386
R10509 VPWR.n2859 VPWR.n2858 93.3652
R10510 VPWR.n1231 VPWR.n1230 91.8492
R10511 VPWR.n1153 VPWR.n1152 91.8492
R10512 VPWR.n1227 VPWR.n1226 91.8492
R10513 VPWR.n1485 VPWR.n1484 91.8492
R10514 VPWR.n1173 VPWR.n1172 91.8492
R10515 VPWR.n1169 VPWR.n1168 91.8492
R10516 VPWR.n1163 VPWR.n1162 91.8492
R10517 VPWR.n1479 VPWR.n1478 91.8492
R10518 VPWR.n1159 VPWR.n1158 91.8492
R10519 VPWR.n1149 VPWR.n1148 91.8492
R10520 VPWR.n1472 VPWR.n1471 91.8492
R10521 VPWR.n1049 VPWR.n1048 91.8492
R10522 VPWR.n1748 VPWR.n1747 91.8492
R10523 VPWR.n1036 VPWR.n1035 91.8492
R10524 VPWR.n1032 VPWR.n1031 91.8492
R10525 VPWR.n1053 VPWR.n1052 91.8492
R10526 VPWR.n2847 VPWR.n2820 91.4829
R10527 VPWR.t693 VPWR.n2842 90.0872
R10528 VPWR.t272 VPWR 88.7855
R10529 VPWR.n1235 VPWR 79.407
R10530 VPWR.n1258 VPWR 79.407
R10531 VPWR.n1282 VPWR 79.407
R10532 VPWR.n1367 VPWR 79.407
R10533 VPWR.n1406 VPWR 79.407
R10534 VPWR.t135 VPWR.t1852 78.8874
R10535 VPWR.n2840 VPWR.n2818 74.9181
R10536 VPWR.n2858 VPWR.n2818 74.9181
R10537 VPWR.n2858 VPWR.n2857 74.9181
R10538 VPWR.n2857 VPWR.n2820 74.9181
R10539 VPWR.t396 VPWR.t1119 70.4952
R10540 VPWR.t1119 VPWR.t933 70.4952
R10541 VPWR.t933 VPWR.t983 70.4952
R10542 VPWR.t983 VPWR.t1766 70.4952
R10543 VPWR.t1766 VPWR.t1196 70.4952
R10544 VPWR.t1196 VPWR.t330 70.4952
R10545 VPWR.t330 VPWR.t1192 70.4952
R10546 VPWR.t248 VPWR.t1088 70.4952
R10547 VPWR.t1082 VPWR.t248 70.4952
R10548 VPWR.t302 VPWR.t1082 70.4952
R10549 VPWR.t1090 VPWR.t302 70.4952
R10550 VPWR.t243 VPWR.t1090 70.4952
R10551 VPWR.t1084 VPWR.t243 70.4952
R10552 VPWR.t311 VPWR.t1084 70.4952
R10553 VPWR VPWR.t396 68.8168
R10554 VPWR.t1104 VPWR.t1100 68.8168
R10555 VPWR.t1852 VPWR.t1233 62.103
R10556 VPWR VPWR.t1096 60.4245
R10557 VPWR.n2849 VPWR.n2842 59.762
R10558 VPWR.n2845 VPWR.n2819 53.8358
R10559 VPWR.t1100 VPWR.t833 52.0323
R10560 VPWR.t1232 VPWR 50.3539
R10561 VPWR VPWR.t1104 50.3539
R10562 VPWR VPWR.t1098 50.3539
R10563 VPWR.t276 VPWR 50.3539
R10564 VPWR.t299 VPWR 50.3539
R10565 VPWR.t251 VPWR 50.3539
R10566 VPWR.n2854 VPWR.n2818 46.2505
R10567 VPWR.n2855 VPWR.n2854 46.2505
R10568 VPWR.n2835 VPWR.n2834 46.2505
R10569 VPWR.n2836 VPWR.n2835 46.2505
R10570 VPWR.n2838 VPWR.n2837 46.2505
R10571 VPWR.n2837 VPWR.n2836 46.2505
R10572 VPWR.n2844 VPWR.n2824 46.2505
R10573 VPWR.n2857 VPWR.n2856 46.2505
R10574 VPWR.n2856 VPWR.n2855 46.2505
R10575 VPWR.n2849 VPWR.n2848 46.2505
R10576 VPWR.n2846 VPWR.n2845 45.9299
R10577 VPWR.n2832 VPWR.n2830 44.8005
R10578 VPWR.n2830 VPWR.n2826 44.8005
R10579 VPWR.n2847 VPWR.n2843 37.0005
R10580 VPWR.n2843 VPWR.t193 37.0005
R10581 VPWR.n1230 VPWR.n1229 34.7473
R10582 VPWR.n1152 VPWR.n1151 34.7473
R10583 VPWR.n1226 VPWR.n1225 34.7473
R10584 VPWR.n1484 VPWR.n1483 34.7473
R10585 VPWR.n1172 VPWR.n1171 34.7473
R10586 VPWR.n1168 VPWR.n1167 34.7473
R10587 VPWR.n1162 VPWR.n1161 34.7473
R10588 VPWR.n1478 VPWR.n1477 34.7473
R10589 VPWR.n1158 VPWR.n1157 34.7473
R10590 VPWR.n1148 VPWR.n1147 34.7473
R10591 VPWR.n1471 VPWR.n1470 34.7473
R10592 VPWR.n1048 VPWR.n1047 34.7473
R10593 VPWR.n1747 VPWR.n1746 34.7473
R10594 VPWR.n1035 VPWR.n1034 34.7473
R10595 VPWR.n1031 VPWR.n1030 34.7473
R10596 VPWR.n1052 VPWR.n1051 34.7473
R10597 VPWR.n1299 VPWR.n1298 34.6358
R10598 VPWR.n1357 VPWR.n1341 34.6358
R10599 VPWR.n1362 VPWR.n1361 34.6358
R10600 VPWR.n1396 VPWR.n1380 34.6358
R10601 VPWR.n1401 VPWR.n1400 34.6358
R10602 VPWR.n1411 VPWR.n1377 34.6358
R10603 VPWR.n1433 VPWR.n1417 34.6358
R10604 VPWR.n1438 VPWR.n1437 34.6358
R10605 VPWR.n2755 VPWR.n2754 34.6358
R10606 VPWR.n2721 VPWR.n2713 34.6358
R10607 VPWR.n2728 VPWR.n2727 34.6358
R10608 VPWR.n2685 VPWR.n2676 34.6358
R10609 VPWR.n2688 VPWR.n2687 34.6358
R10610 VPWR.n2692 VPWR.n2691 34.6358
R10611 VPWR.n2648 VPWR.n2639 34.6358
R10612 VPWR.n2651 VPWR.n2650 34.6358
R10613 VPWR.n2655 VPWR.n2654 34.6358
R10614 VPWR.n2662 VPWR.n2661 34.6358
R10615 VPWR.n2615 VPWR.n2611 34.6358
R10616 VPWR.n2619 VPWR.n2603 34.6358
R10617 VPWR.n2622 VPWR.n2621 34.6358
R10618 VPWR.n1316 VPWR.n1315 32.0005
R10619 VPWR.n1353 VPWR.n1352 32.0005
R10620 VPWR.n1392 VPWR.n1391 32.0005
R10621 VPWR.n1429 VPWR.n1428 32.0005
R10622 VPWR.n2717 VPWR.n2716 30.8711
R10623 VPWR.n2681 VPWR.n2680 30.8711
R10624 VPWR.n2644 VPWR.n2643 30.8711
R10625 VPWR.n2610 VPWR.n2609 30.8711
R10626 VPWR.n2834 VPWR.n2832 30.1181
R10627 VPWR.n2838 VPWR.n2826 30.1181
R10628 VPWR.n2848 VPWR.n2846 28.9887
R10629 VPWR.n1325 VPWR.n1324 28.2358
R10630 VPWR.n5 VPWR.t986 26.5955
R10631 VPWR.n5 VPWR.t1195 26.5955
R10632 VPWR.n4 VPWR.t1118 26.5955
R10633 VPWR.n4 VPWR.t982 26.5955
R10634 VPWR.n1240 VPWR.t53 26.5955
R10635 VPWR.n1240 VPWR.t52 26.5955
R10636 VPWR.n1239 VPWR.t1311 26.5955
R10637 VPWR.n1239 VPWR.t1768 26.5955
R10638 VPWR.n1245 VPWR.t48 26.5955
R10639 VPWR.n1245 VPWR.t54 26.5955
R10640 VPWR.n1238 VPWR.t628 26.5955
R10641 VPWR.n1238 VPWR.t631 26.5955
R10642 VPWR.n1263 VPWR.t1845 26.5955
R10643 VPWR.n1263 VPWR.t1846 26.5955
R10644 VPWR.n1262 VPWR.t412 26.5955
R10645 VPWR.n1262 VPWR.t409 26.5955
R10646 VPWR.n1268 VPWR.t1030 26.5955
R10647 VPWR.n1268 VPWR.t158 26.5955
R10648 VPWR.n1261 VPWR.t415 26.5955
R10649 VPWR.n1261 VPWR.t413 26.5955
R10650 VPWR.n1287 VPWR.t757 26.5955
R10651 VPWR.n1287 VPWR.t764 26.5955
R10652 VPWR.n1286 VPWR.t915 26.5955
R10653 VPWR.n1286 VPWR.t914 26.5955
R10654 VPWR.n1292 VPWR.t761 26.5955
R10655 VPWR.n1292 VPWR.t758 26.5955
R10656 VPWR.n1285 VPWR.t918 26.5955
R10657 VPWR.n1285 VPWR.t916 26.5955
R10658 VPWR.n1314 VPWR.t233 26.5955
R10659 VPWR.n1314 VPWR.t444 26.5955
R10660 VPWR.n1307 VPWR.t1193 26.5955
R10661 VPWR.n1307 VPWR.t231 26.5955
R10662 VPWR.n1321 VPWR.t984 26.5955
R10663 VPWR.n1321 VPWR.t1197 26.5955
R10664 VPWR.n1323 VPWR.t934 26.5955
R10665 VPWR.n1323 VPWR.t1767 26.5955
R10666 VPWR.n1351 VPWR.t954 26.5955
R10667 VPWR.n1351 VPWR.t1764 26.5955
R10668 VPWR.n1350 VPWR.t1329 26.5955
R10669 VPWR.n1350 VPWR.t333 26.5955
R10670 VPWR.n1344 VPWR.t56 26.5955
R10671 VPWR.n1344 VPWR.t937 26.5955
R10672 VPWR.n1343 VPWR.t629 26.5955
R10673 VPWR.n1343 VPWR.t1327 26.5955
R10674 VPWR.n1359 VPWR.t51 26.5955
R10675 VPWR.n1359 VPWR.t50 26.5955
R10676 VPWR.n1358 VPWR.t1769 26.5955
R10677 VPWR.n1358 VPWR.t630 26.5955
R10678 VPWR.n1390 VPWR.t1326 26.5955
R10679 VPWR.n1390 VPWR.t449 26.5955
R10680 VPWR.n1389 VPWR.t956 26.5955
R10681 VPWR.n1389 VPWR.t1765 26.5955
R10682 VPWR.n1383 VPWR.t1028 26.5955
R10683 VPWR.n1383 VPWR.t446 26.5955
R10684 VPWR.n1382 VPWR.t416 26.5955
R10685 VPWR.n1382 VPWR.t952 26.5955
R10686 VPWR.n1398 VPWR.t1847 26.5955
R10687 VPWR.n1398 VPWR.t1029 26.5955
R10688 VPWR.n1397 VPWR.t417 26.5955
R10689 VPWR.n1397 VPWR.t414 26.5955
R10690 VPWR.n1427 VPWR.t395 26.5955
R10691 VPWR.n1427 VPWR.t935 26.5955
R10692 VPWR.n1426 VPWR.t448 26.5955
R10693 VPWR.n1426 VPWR.t390 26.5955
R10694 VPWR.n1420 VPWR.t760 26.5955
R10695 VPWR.n1420 VPWR.t392 26.5955
R10696 VPWR.n1419 VPWR.t912 26.5955
R10697 VPWR.n1419 VPWR.t1328 26.5955
R10698 VPWR.n1435 VPWR.t763 26.5955
R10699 VPWR.n1435 VPWR.t762 26.5955
R10700 VPWR.n1434 VPWR.t913 26.5955
R10701 VPWR.n1434 VPWR.t911 26.5955
R10702 VPWR.n2802 VPWR.t1093 26.5955
R10703 VPWR.n2802 VPWR.t1095 26.5955
R10704 VPWR.n2804 VPWR.t1087 26.5955
R10705 VPWR.n2804 VPWR.t1081 26.5955
R10706 VPWR.n2782 VPWR.t932 26.5955
R10707 VPWR.n2782 VPWR.t929 26.5955
R10708 VPWR.n2783 VPWR.t653 26.5955
R10709 VPWR.n2783 VPWR.t647 26.5955
R10710 VPWR.n2786 VPWR.t925 26.5955
R10711 VPWR.n2786 VPWR.t926 26.5955
R10712 VPWR.n2787 VPWR.t639 26.5955
R10713 VPWR.n2787 VPWR.t641 26.5955
R10714 VPWR.n2762 VPWR.t466 26.5955
R10715 VPWR.n2762 VPWR.t476 26.5955
R10716 VPWR.n2763 VPWR.t749 26.5955
R10717 VPWR.n2763 VPWR.t755 26.5955
R10718 VPWR.n2766 VPWR.t468 26.5955
R10719 VPWR.n2766 VPWR.t470 26.5955
R10720 VPWR.n2767 VPWR.t751 26.5955
R10721 VPWR.n2767 VPWR.t753 26.5955
R10722 VPWR.n2743 VPWR.t125 26.5955
R10723 VPWR.n2743 VPWR.t119 26.5955
R10724 VPWR.n2744 VPWR.t991 26.5955
R10725 VPWR.n2744 VPWR.t990 26.5955
R10726 VPWR.n2747 VPWR.t127 26.5955
R10727 VPWR.n2747 VPWR.t129 26.5955
R10728 VPWR.n2748 VPWR.t993 26.5955
R10729 VPWR.n2748 VPWR.t987 26.5955
R10730 VPWR.n2708 VPWR.t303 26.5955
R10731 VPWR.n2708 VPWR.t244 26.5955
R10732 VPWR.n2712 VPWR.t323 26.5955
R10733 VPWR.n2712 VPWR.t1089 26.5955
R10734 VPWR.n2715 VPWR.t224 26.5955
R10735 VPWR.n2715 VPWR.t1834 26.5955
R10736 VPWR.n2709 VPWR.t1083 26.5955
R10737 VPWR.n2709 VPWR.t1091 26.5955
R10738 VPWR.n2679 VPWR.t227 26.5955
R10739 VPWR.n2679 VPWR.t1835 26.5955
R10740 VPWR.n2678 VPWR.t238 26.5955
R10741 VPWR.n2678 VPWR.t310 26.5955
R10742 VPWR.n2675 VPWR.t324 26.5955
R10743 VPWR.n2675 VPWR.t649 26.5955
R10744 VPWR.n2674 VPWR.t275 26.5955
R10745 VPWR.n2674 VPWR.t930 26.5955
R10746 VPWR.n2671 VPWR.t643 26.5955
R10747 VPWR.n2671 VPWR.t651 26.5955
R10748 VPWR.n2670 VPWR.t927 26.5955
R10749 VPWR.n2670 VPWR.t931 26.5955
R10750 VPWR.n2642 VPWR.t236 26.5955
R10751 VPWR.n2642 VPWR.t215 26.5955
R10752 VPWR.n2641 VPWR.t280 26.5955
R10753 VPWR.n2641 VPWR.t242 26.5955
R10754 VPWR.n2638 VPWR.t271 26.5955
R10755 VPWR.n2638 VPWR.t754 26.5955
R10756 VPWR.n2637 VPWR.t314 26.5955
R10757 VPWR.n2637 VPWR.t462 26.5955
R10758 VPWR.n2634 VPWR.t750 26.5955
R10759 VPWR.n2634 VPWR.t756 26.5955
R10760 VPWR.n2633 VPWR.t472 26.5955
R10761 VPWR.n2633 VPWR.t464 26.5955
R10762 VPWR.n2606 VPWR.t240 26.5955
R10763 VPWR.n2606 VPWR.t325 26.5955
R10764 VPWR.n2605 VPWR.t1830 26.5955
R10765 VPWR.n2605 VPWR.t246 26.5955
R10766 VPWR.n2613 VPWR.t254 26.5955
R10767 VPWR.n2613 VPWR.t992 26.5955
R10768 VPWR.n2612 VPWR.t297 26.5955
R10769 VPWR.n2612 VPWR.t121 26.5955
R10770 VPWR.n2602 VPWR.t994 26.5955
R10771 VPWR.n2602 VPWR.t988 26.5955
R10772 VPWR.n2601 VPWR.t115 26.5955
R10773 VPWR.n2601 VPWR.t123 26.5955
R10774 VPWR.n17 VPWR.n16 25.977
R10775 VPWR.n1253 VPWR.n1252 25.977
R10776 VPWR.n1313 VPWR.n1310 25.977
R10777 VPWR.n1349 VPWR.n1346 25.977
R10778 VPWR.n1372 VPWR.n1338 25.977
R10779 VPWR.n1388 VPWR.n1385 25.977
R10780 VPWR.n1425 VPWR.n1422 25.977
R10781 VPWR.n2811 VPWR.n2810 25.977
R10782 VPWR.n2795 VPWR.n2794 25.977
R10783 VPWR.n2717 VPWR.n2714 25.977
R10784 VPWR.n2681 VPWR.n2677 25.977
R10785 VPWR.n2699 VPWR.n2698 25.977
R10786 VPWR.n2644 VPWR.n2640 25.977
R10787 VPWR.n2609 VPWR.n2607 25.977
R10788 VPWR.n1335 VPWR.n1334 25.224
R10789 VPWR.n2737 VPWR.n2736 25.224
R10790 VPWR.n2722 VPWR.n2721 24.8476
R10791 VPWR.n2686 VPWR.n2685 24.8476
R10792 VPWR.n2649 VPWR.n2648 24.8476
R10793 VPWR.n2615 VPWR.n2614 24.8476
R10794 VPWR.n16 VPWR.n15 24.4711
R10795 VPWR.n1252 VPWR.n1251 24.4711
R10796 VPWR.n1315 VPWR.n1313 24.4711
R10797 VPWR.n1352 VPWR.n1349 24.4711
R10798 VPWR.n1391 VPWR.n1388 24.4711
R10799 VPWR.n1428 VPWR.n1425 24.4711
R10800 VPWR.n2810 VPWR.n2809 24.4711
R10801 VPWR.n2794 VPWR.n2793 24.4711
R10802 VPWR.n11 VPWR.n2 23.7181
R10803 VPWR.n1247 VPWR.n1236 23.7181
R10804 VPWR.n1270 VPWR.n1259 23.7181
R10805 VPWR.n1274 VPWR.n1259 23.7181
R10806 VPWR.n1294 VPWR.n1283 23.7181
R10807 VPWR.n1298 VPWR.n1283 23.7181
R10808 VPWR.n1330 VPWR.n1328 23.7181
R10809 VPWR.n1368 VPWR.n1365 23.7181
R10810 VPWR.n1407 VPWR.n1404 23.7181
R10811 VPWR.n1407 VPWR.n1377 23.7181
R10812 VPWR.n1444 VPWR.n1441 23.7181
R10813 VPWR.n2808 VPWR.n2807 23.7181
R10814 VPWR.n2789 VPWR.n2781 23.7181
R10815 VPWR.n2769 VPWR.n2761 23.7181
R10816 VPWR.n2773 VPWR.n2761 23.7181
R10817 VPWR.n2750 VPWR.n2742 23.7181
R10818 VPWR.n2754 VPWR.n2742 23.7181
R10819 VPWR.n2731 VPWR.n2706 23.7181
R10820 VPWR.n2694 VPWR.n2668 23.7181
R10821 VPWR.n2657 VPWR.n2631 23.7181
R10822 VPWR.n2661 VPWR.n2631 23.7181
R10823 VPWR.n2626 VPWR.n2625 23.7181
R10824 VPWR.t1200 VPWR.t747 23.4987
R10825 VPWR.t191 VPWR.t133 23.4987
R10826 VPWR.n2852 VPWR.n2841 23.1255
R10827 VPWR.n2852 VPWR.t693 23.1255
R10828 VPWR.n2851 VPWR.n2819 23.1255
R10829 VPWR.t693 VPWR.n2851 23.1255
R10830 VPWR.n11 VPWR.n10 22.9652
R10831 VPWR.n1247 VPWR.n1246 22.9652
R10832 VPWR.n1270 VPWR.n1269 22.9652
R10833 VPWR.n1294 VPWR.n1293 22.9652
R10834 VPWR.n2807 VPWR.n2803 22.9652
R10835 VPWR.n2789 VPWR.n2788 22.9652
R10836 VPWR.n2769 VPWR.n2768 22.9652
R10837 VPWR.n2750 VPWR.n2749 22.9652
R10838 VPWR.n1320 VPWR.n1308 22.2123
R10839 VPWR.n2724 VPWR.n2723 22.2123
R10840 VPWR.n10 VPWR.n3 21.4593
R10841 VPWR.n1246 VPWR.n1237 21.4593
R10842 VPWR.n1269 VPWR.n1260 21.4593
R10843 VPWR.n1293 VPWR.n1284 21.4593
R10844 VPWR.n1442 VPWR.t389 20.5957
R10845 VPWR.n1443 VPWR.t391 20.5957
R10846 VPWR.n1277 VPWR.n1276 19.9534
R10847 VPWR.n1300 VPWR.n1299 19.9534
R10848 VPWR.n1334 VPWR.n1303 19.9534
R10849 VPWR.n2776 VPWR.n2775 19.9534
R10850 VPWR.n2756 VPWR.n2755 19.9534
R10851 VPWR.n2736 VPWR.n2735 19.9534
R10852 VPWR.n2724 VPWR.n2710 18.824
R10853 VPWR.n2688 VPWR.n2672 18.824
R10854 VPWR.n2651 VPWR.n2635 18.824
R10855 VPWR.n2620 VPWR.n2619 18.824
R10856 VPWR.n1316 VPWR.n1308 18.4476
R10857 VPWR.n1353 VPWR.n1345 18.4476
R10858 VPWR.n1373 VPWR.n1372 18.4476
R10859 VPWR.n1392 VPWR.n1384 18.4476
R10860 VPWR.n1429 VPWR.n1421 18.4476
R10861 VPWR.n2700 VPWR.n2699 18.4476
R10862 VPWR.n1413 VPWR.n1412 17.5829
R10863 VPWR.n2664 VPWR.n2663 17.5829
R10864 VPWR.n6 VPWR.n3 16.9417
R10865 VPWR.n1241 VPWR.n1237 16.9417
R10866 VPWR.n1264 VPWR.n1260 16.9417
R10867 VPWR.n1288 VPWR.n1284 16.9417
R10868 VPWR.n2730 VPWR.n2729 16.5652
R10869 VPWR.n1306 VPWR.n1304 16.1887
R10870 VPWR.n1374 VPWR.n1373 16.1887
R10871 VPWR.n2701 VPWR.n2700 16.1887
R10872 VPWR.n1235 VPWR.t47 16.0935
R10873 VPWR.n1258 VPWR.t157 16.0935
R10874 VPWR.n1282 VPWR.t81 16.0935
R10875 VPWR.n1367 VPWR.t49 16.0935
R10876 VPWR.n1406 VPWR.t155 16.0935
R10877 VPWR.n1234 VPWR.t398 16.0935
R10878 VPWR.n1257 VPWR.t229 16.0935
R10879 VPWR.n1281 VPWR.t234 16.0935
R10880 VPWR.n1366 VPWR.t159 16.0935
R10881 VPWR.n1405 VPWR.t410 16.0935
R10882 VPWR.n1325 VPWR.n1306 15.8123
R10883 VPWR.n2727 VPWR.n2710 15.8123
R10884 VPWR.n2729 VPWR.n2728 15.8123
R10885 VPWR.n2691 VPWR.n2672 15.8123
R10886 VPWR.n2654 VPWR.n2635 15.8123
R10887 VPWR.n2621 VPWR.n2620 15.8123
R10888 VPWR.n1330 VPWR.n1303 13.5534
R10889 VPWR.n2735 VPWR.n2706 13.5534
R10890 VPWR.n2839 VPWR.n2823 13.2148
R10891 VPWR.n2823 VPWR.t668 13.2148
R10892 VPWR.n2827 VPWR.n2817 13.2148
R10893 VPWR.n2827 VPWR.t668 13.2148
R10894 VPWR.n2833 VPWR.n2829 13.2148
R10895 VPWR.n2829 VPWR.t668 13.2148
R10896 VPWR.n15 VPWR.n2 12.8005
R10897 VPWR.n1251 VPWR.n1236 12.8005
R10898 VPWR.n1368 VPWR.n1338 12.8005
R10899 VPWR.n2809 VPWR.n2808 12.8005
R10900 VPWR.n2793 VPWR.n2781 12.8005
R10901 VPWR.n2698 VPWR.n2668 12.8005
R10902 VPWR.n1322 VPWR.n1320 12.424
R10903 VPWR.n1360 VPWR.n1357 12.424
R10904 VPWR.n1399 VPWR.n1396 12.424
R10905 VPWR.n1436 VPWR.n1433 12.424
R10906 VPWR.n1276 VPWR.n1275 10.5417
R10907 VPWR.n1412 VPWR.n1411 10.5417
R10908 VPWR.n2775 VPWR.n2774 10.5417
R10909 VPWR.n2663 VPWR.n2662 10.5417
R10910 VPWR.n2687 VPWR.n2686 9.78874
R10911 VPWR.n2650 VPWR.n2649 9.78874
R10912 VPWR.n2614 VPWR.n2603 9.78874
R10913 VPWR.n1361 VPWR.n1360 9.41227
R10914 VPWR.n1365 VPWR.n1339 9.41227
R10915 VPWR.n1400 VPWR.n1399 9.41227
R10916 VPWR.n1404 VPWR.n1378 9.41227
R10917 VPWR.n1437 VPWR.n1436 9.41227
R10918 VPWR.n1441 VPWR.n1415 9.41227
R10919 VPWR.n2694 VPWR.n2693 9.41227
R10920 VPWR.n2657 VPWR.n2656 9.41227
R10921 VPWR.n2625 VPWR.n2599 9.41227
R10922 VPWR.n1229 VPWR 9.37021
R10923 VPWR.n1151 VPWR 9.37021
R10924 VPWR.n1225 VPWR 9.37021
R10925 VPWR.n1483 VPWR 9.37021
R10926 VPWR.n1171 VPWR 9.37021
R10927 VPWR.n1167 VPWR 9.37021
R10928 VPWR.n1161 VPWR 9.37021
R10929 VPWR.n1477 VPWR 9.37021
R10930 VPWR.n1157 VPWR 9.37021
R10931 VPWR.n1147 VPWR 9.37021
R10932 VPWR.n1470 VPWR 9.37021
R10933 VPWR.n1047 VPWR 9.37021
R10934 VPWR.n1746 VPWR 9.37021
R10935 VPWR.n1034 VPWR 9.37021
R10936 VPWR.n1030 VPWR 9.37021
R10937 VPWR.n1051 VPWR 9.37021
R10938 VPWR.n1467 VPWR.n1466 9.33404
R10939 VPWR.n352 VPWR.n351 9.33404
R10940 VPWR.n1534 VPWR.n1533 9.33404
R10941 VPWR.n348 VPWR.n347 9.33404
R10942 VPWR.n965 VPWR.n964 9.33404
R10943 VPWR.n2479 VPWR.n2478 9.33404
R10944 VPWR.n2475 VPWR.n2474 9.33404
R10945 VPWR.n320 VPWR.n319 9.33404
R10946 VPWR.n973 VPWR.n972 9.33404
R10947 VPWR.n2445 VPWR.n2444 9.33404
R10948 VPWR.n324 VPWR.n323 9.33404
R10949 VPWR.n1891 VPWR.n1890 9.33404
R10950 VPWR.n1887 VPWR.n1886 9.33404
R10951 VPWR.n1881 VPWR.n1880 9.33404
R10952 VPWR.n389 VPWR.n388 9.33404
R10953 VPWR.n393 VPWR.n392 9.33404
R10954 VPWR.n397 VPWR.n396 9.33404
R10955 VPWR.n2455 VPWR.n2454 9.33404
R10956 VPWR.n332 VPWR.n331 9.33404
R10957 VPWR.n1877 VPWR.n1876 9.33404
R10958 VPWR.n405 VPWR.n404 9.33404
R10959 VPWR.n2459 VPWR.n2458 9.33404
R10960 VPWR.n336 VPWR.n335 9.33404
R10961 VPWR.n2308 VPWR.n2307 9.33404
R10962 VPWR.n2312 VPWR.n2311 9.33404
R10963 VPWR.n2318 VPWR.n2317 9.33404
R10964 VPWR.n2322 VPWR.n2321 9.33404
R10965 VPWR.n2332 VPWR.n2331 9.33404
R10966 VPWR.n2338 VPWR.n2337 9.33404
R10967 VPWR.n2342 VPWR.n2341 9.33404
R10968 VPWR.n2348 VPWR.n2347 9.33404
R10969 VPWR.n2352 VPWR.n2351 9.33404
R10970 VPWR.n2358 VPWR.n2357 9.33404
R10971 VPWR.n2362 VPWR.n2361 9.33404
R10972 VPWR.n2368 VPWR.n2367 9.33404
R10973 VPWR.n2372 VPWR.n2371 9.33404
R10974 VPWR.n2378 VPWR.n2377 9.33404
R10975 VPWR.n2381 VPWR.n2380 9.33404
R10976 VPWR.n2328 VPWR.n2327 9.33404
R10977 VPWR.n544 VPWR.n543 9.33404
R10978 VPWR.n540 VPWR.n539 9.33404
R10979 VPWR.n536 VPWR.n535 9.33404
R10980 VPWR.n532 VPWR.n531 9.33404
R10981 VPWR.n524 VPWR.n523 9.33404
R10982 VPWR.n520 VPWR.n519 9.33404
R10983 VPWR.n516 VPWR.n515 9.33404
R10984 VPWR.n512 VPWR.n511 9.33404
R10985 VPWR.n508 VPWR.n507 9.33404
R10986 VPWR.n504 VPWR.n503 9.33404
R10987 VPWR.n500 VPWR.n499 9.33404
R10988 VPWR.n496 VPWR.n495 9.33404
R10989 VPWR.n492 VPWR.n491 9.33404
R10990 VPWR.n488 VPWR.n487 9.33404
R10991 VPWR.n485 VPWR.n484 9.33404
R10992 VPWR.n528 VPWR.n527 9.33404
R10993 VPWR.n2283 VPWR.n2282 9.33404
R10994 VPWR.n2279 VPWR.n2278 9.33404
R10995 VPWR.n2273 VPWR.n2272 9.33404
R10996 VPWR.n2269 VPWR.n2268 9.33404
R10997 VPWR.n2259 VPWR.n2258 9.33404
R10998 VPWR.n2253 VPWR.n2252 9.33404
R10999 VPWR.n2249 VPWR.n2248 9.33404
R11000 VPWR.n2243 VPWR.n2242 9.33404
R11001 VPWR.n2239 VPWR.n2238 9.33404
R11002 VPWR.n2233 VPWR.n2232 9.33404
R11003 VPWR.n2229 VPWR.n2228 9.33404
R11004 VPWR.n2223 VPWR.n2222 9.33404
R11005 VPWR.n2219 VPWR.n2218 9.33404
R11006 VPWR.n2213 VPWR.n2212 9.33404
R11007 VPWR.n2210 VPWR.n2209 9.33404
R11008 VPWR.n2263 VPWR.n2262 9.33404
R11009 VPWR.n581 VPWR.n580 9.33404
R11010 VPWR.n585 VPWR.n584 9.33404
R11011 VPWR.n589 VPWR.n588 9.33404
R11012 VPWR.n593 VPWR.n592 9.33404
R11013 VPWR.n601 VPWR.n600 9.33404
R11014 VPWR.n605 VPWR.n604 9.33404
R11015 VPWR.n609 VPWR.n608 9.33404
R11016 VPWR.n613 VPWR.n612 9.33404
R11017 VPWR.n617 VPWR.n616 9.33404
R11018 VPWR.n621 VPWR.n620 9.33404
R11019 VPWR.n625 VPWR.n624 9.33404
R11020 VPWR.n629 VPWR.n628 9.33404
R11021 VPWR.n633 VPWR.n632 9.33404
R11022 VPWR.n637 VPWR.n636 9.33404
R11023 VPWR.n640 VPWR.n639 9.33404
R11024 VPWR.n597 VPWR.n596 9.33404
R11025 VPWR.n2112 VPWR.n2111 9.33404
R11026 VPWR.n2116 VPWR.n2115 9.33404
R11027 VPWR.n2122 VPWR.n2121 9.33404
R11028 VPWR.n2126 VPWR.n2125 9.33404
R11029 VPWR.n2136 VPWR.n2135 9.33404
R11030 VPWR.n2142 VPWR.n2141 9.33404
R11031 VPWR.n2146 VPWR.n2145 9.33404
R11032 VPWR.n2152 VPWR.n2151 9.33404
R11033 VPWR.n2156 VPWR.n2155 9.33404
R11034 VPWR.n2162 VPWR.n2161 9.33404
R11035 VPWR.n2166 VPWR.n2165 9.33404
R11036 VPWR.n2172 VPWR.n2171 9.33404
R11037 VPWR.n2176 VPWR.n2175 9.33404
R11038 VPWR.n2182 VPWR.n2181 9.33404
R11039 VPWR.n2185 VPWR.n2184 9.33404
R11040 VPWR.n2132 VPWR.n2131 9.33404
R11041 VPWR.n736 VPWR.n735 9.33404
R11042 VPWR.n732 VPWR.n731 9.33404
R11043 VPWR.n728 VPWR.n727 9.33404
R11044 VPWR.n724 VPWR.n723 9.33404
R11045 VPWR.n716 VPWR.n715 9.33404
R11046 VPWR.n712 VPWR.n711 9.33404
R11047 VPWR.n708 VPWR.n707 9.33404
R11048 VPWR.n704 VPWR.n703 9.33404
R11049 VPWR.n700 VPWR.n699 9.33404
R11050 VPWR.n696 VPWR.n695 9.33404
R11051 VPWR.n692 VPWR.n691 9.33404
R11052 VPWR.n688 VPWR.n687 9.33404
R11053 VPWR.n684 VPWR.n683 9.33404
R11054 VPWR.n680 VPWR.n679 9.33404
R11055 VPWR.n677 VPWR.n676 9.33404
R11056 VPWR.n720 VPWR.n719 9.33404
R11057 VPWR.n2087 VPWR.n2086 9.33404
R11058 VPWR.n2083 VPWR.n2082 9.33404
R11059 VPWR.n2077 VPWR.n2076 9.33404
R11060 VPWR.n2073 VPWR.n2072 9.33404
R11061 VPWR.n2063 VPWR.n2062 9.33404
R11062 VPWR.n2057 VPWR.n2056 9.33404
R11063 VPWR.n2053 VPWR.n2052 9.33404
R11064 VPWR.n2047 VPWR.n2046 9.33404
R11065 VPWR.n2043 VPWR.n2042 9.33404
R11066 VPWR.n2037 VPWR.n2036 9.33404
R11067 VPWR.n2033 VPWR.n2032 9.33404
R11068 VPWR.n2027 VPWR.n2026 9.33404
R11069 VPWR.n2023 VPWR.n2022 9.33404
R11070 VPWR.n2017 VPWR.n2016 9.33404
R11071 VPWR.n2014 VPWR.n2013 9.33404
R11072 VPWR.n2067 VPWR.n2066 9.33404
R11073 VPWR.n773 VPWR.n772 9.33404
R11074 VPWR.n777 VPWR.n776 9.33404
R11075 VPWR.n781 VPWR.n780 9.33404
R11076 VPWR.n785 VPWR.n784 9.33404
R11077 VPWR.n793 VPWR.n792 9.33404
R11078 VPWR.n797 VPWR.n796 9.33404
R11079 VPWR.n801 VPWR.n800 9.33404
R11080 VPWR.n805 VPWR.n804 9.33404
R11081 VPWR.n809 VPWR.n808 9.33404
R11082 VPWR.n813 VPWR.n812 9.33404
R11083 VPWR.n817 VPWR.n816 9.33404
R11084 VPWR.n821 VPWR.n820 9.33404
R11085 VPWR.n825 VPWR.n824 9.33404
R11086 VPWR.n829 VPWR.n828 9.33404
R11087 VPWR.n832 VPWR.n831 9.33404
R11088 VPWR.n789 VPWR.n788 9.33404
R11089 VPWR.n1916 VPWR.n1915 9.33404
R11090 VPWR.n1920 VPWR.n1919 9.33404
R11091 VPWR.n1926 VPWR.n1925 9.33404
R11092 VPWR.n1930 VPWR.n1929 9.33404
R11093 VPWR.n1940 VPWR.n1939 9.33404
R11094 VPWR.n1946 VPWR.n1945 9.33404
R11095 VPWR.n1950 VPWR.n1949 9.33404
R11096 VPWR.n1956 VPWR.n1955 9.33404
R11097 VPWR.n1960 VPWR.n1959 9.33404
R11098 VPWR.n1966 VPWR.n1965 9.33404
R11099 VPWR.n1970 VPWR.n1969 9.33404
R11100 VPWR.n1976 VPWR.n1975 9.33404
R11101 VPWR.n1980 VPWR.n1979 9.33404
R11102 VPWR.n1986 VPWR.n1985 9.33404
R11103 VPWR.n1989 VPWR.n1988 9.33404
R11104 VPWR.n1936 VPWR.n1935 9.33404
R11105 VPWR.n928 VPWR.n927 9.33404
R11106 VPWR.n924 VPWR.n923 9.33404
R11107 VPWR.n920 VPWR.n919 9.33404
R11108 VPWR.n916 VPWR.n915 9.33404
R11109 VPWR.n908 VPWR.n907 9.33404
R11110 VPWR.n904 VPWR.n903 9.33404
R11111 VPWR.n900 VPWR.n899 9.33404
R11112 VPWR.n896 VPWR.n895 9.33404
R11113 VPWR.n892 VPWR.n891 9.33404
R11114 VPWR.n888 VPWR.n887 9.33404
R11115 VPWR.n884 VPWR.n883 9.33404
R11116 VPWR.n880 VPWR.n879 9.33404
R11117 VPWR.n876 VPWR.n875 9.33404
R11118 VPWR.n872 VPWR.n871 9.33404
R11119 VPWR.n869 VPWR.n868 9.33404
R11120 VPWR.n912 VPWR.n911 9.33404
R11121 VPWR.n1871 VPWR.n1870 9.33404
R11122 VPWR.n981 VPWR.n980 9.33404
R11123 VPWR.n1495 VPWR.n1494 9.33404
R11124 VPWR.n401 VPWR.n400 9.33404
R11125 VPWR.n2465 VPWR.n2464 9.33404
R11126 VPWR.n340 VPWR.n339 9.33404
R11127 VPWR.n977 VPWR.n976 9.33404
R11128 VPWR.n1491 VPWR.n1490 9.33404
R11129 VPWR.n1867 VPWR.n1866 9.33404
R11130 VPWR.n985 VPWR.n984 9.33404
R11131 VPWR.n1505 VPWR.n1504 9.33404
R11132 VPWR.n409 VPWR.n408 9.33404
R11133 VPWR.n417 VPWR.n416 9.33404
R11134 VPWR.n421 VPWR.n420 9.33404
R11135 VPWR.n425 VPWR.n424 9.33404
R11136 VPWR.n429 VPWR.n428 9.33404
R11137 VPWR.n433 VPWR.n432 9.33404
R11138 VPWR.n437 VPWR.n436 9.33404
R11139 VPWR.n441 VPWR.n440 9.33404
R11140 VPWR.n445 VPWR.n444 9.33404
R11141 VPWR.n448 VPWR.n447 9.33404
R11142 VPWR.n413 VPWR.n412 9.33404
R11143 VPWR.n2449 VPWR.n2448 9.33404
R11144 VPWR.n328 VPWR.n327 9.33404
R11145 VPWR.n989 VPWR.n988 9.33404
R11146 VPWR.n1509 VPWR.n1508 9.33404
R11147 VPWR.n1861 VPWR.n1860 9.33404
R11148 VPWR.n1851 VPWR.n1850 9.33404
R11149 VPWR.n1847 VPWR.n1846 9.33404
R11150 VPWR.n1841 VPWR.n1840 9.33404
R11151 VPWR.n1837 VPWR.n1836 9.33404
R11152 VPWR.n1831 VPWR.n1830 9.33404
R11153 VPWR.n1827 VPWR.n1826 9.33404
R11154 VPWR.n1821 VPWR.n1820 9.33404
R11155 VPWR.n1818 VPWR.n1817 9.33404
R11156 VPWR.n1857 VPWR.n1856 9.33404
R11157 VPWR.n993 VPWR.n992 9.33404
R11158 VPWR.n1519 VPWR.n1518 9.33404
R11159 VPWR.n2469 VPWR.n2468 9.33404
R11160 VPWR.n344 VPWR.n343 9.33404
R11161 VPWR.n1480 VPWR.n1130 9.33404
R11162 VPWR.n997 VPWR.n996 9.33404
R11163 VPWR.n1523 VPWR.n1522 9.33404
R11164 VPWR.n2439 VPWR.n2438 9.33404
R11165 VPWR.n2429 VPWR.n2428 9.33404
R11166 VPWR.n2425 VPWR.n2424 9.33404
R11167 VPWR.n2419 VPWR.n2418 9.33404
R11168 VPWR.n2415 VPWR.n2414 9.33404
R11169 VPWR.n2409 VPWR.n2408 9.33404
R11170 VPWR.n2406 VPWR.n2405 9.33404
R11171 VPWR.n2435 VPWR.n2434 9.33404
R11172 VPWR.n316 VPWR.n315 9.33404
R11173 VPWR.n1538 VPWR.n1537 9.33404
R11174 VPWR.n1001 VPWR.n1000 9.33404
R11175 VPWR.n1005 VPWR.n1004 9.33404
R11176 VPWR.n1009 VPWR.n1008 9.33404
R11177 VPWR.n1013 VPWR.n1012 9.33404
R11178 VPWR.n1017 VPWR.n1016 9.33404
R11179 VPWR.n1021 VPWR.n1020 9.33404
R11180 VPWR.n1024 VPWR.n1023 9.33404
R11181 VPWR.n969 VPWR.n968 9.33404
R11182 VPWR.n1474 VPWR.n1473 9.33404
R11183 VPWR.n312 VPWR.n311 9.33404
R11184 VPWR.n1763 VPWR.n1762 9.33404
R11185 VPWR.n308 VPWR.n307 9.33404
R11186 VPWR.n304 VPWR.n303 9.33404
R11187 VPWR.n296 VPWR.n295 9.33404
R11188 VPWR.n293 VPWR.n292 9.33404
R11189 VPWR.n300 VPWR.n299 9.33404
R11190 VPWR.n1751 VPWR.n1750 9.33404
R11191 VPWR.n1790 VPWR.n1789 9.33404
R11192 VPWR.n1793 VPWR.n1792 9.33404
R11193 VPWR.n1759 VPWR.n1758 9.33404
R11194 VPWR.n2714 VPWR 9.32394
R11195 VPWR.n2677 VPWR 9.32394
R11196 VPWR.n2640 VPWR 9.32394
R11197 VPWR VPWR.n2607 9.32394
R11198 VPWR.n18 VPWR.n17 9.3005
R11199 VPWR.n15 VPWR.n14 9.3005
R11200 VPWR.n13 VPWR.n2 9.3005
R11201 VPWR.n10 VPWR.n9 9.3005
R11202 VPWR.n8 VPWR.n3 9.3005
R11203 VPWR.n12 VPWR.n11 9.3005
R11204 VPWR.n16 VPWR.n0 9.3005
R11205 VPWR.n1254 VPWR.n1253 9.3005
R11206 VPWR.n1251 VPWR.n1250 9.3005
R11207 VPWR.n1249 VPWR.n1236 9.3005
R11208 VPWR.n1246 VPWR.n1244 9.3005
R11209 VPWR.n1243 VPWR.n1237 9.3005
R11210 VPWR.n1248 VPWR.n1247 9.3005
R11211 VPWR.n1252 VPWR.n1233 9.3005
R11212 VPWR.n1278 VPWR.n1277 9.3005
R11213 VPWR.n1272 VPWR.n1259 9.3005
R11214 VPWR.n1269 VPWR.n1267 9.3005
R11215 VPWR.n1266 VPWR.n1260 9.3005
R11216 VPWR.n1271 VPWR.n1270 9.3005
R11217 VPWR.n1274 VPWR.n1273 9.3005
R11218 VPWR.n1276 VPWR.n1256 9.3005
R11219 VPWR.n1301 VPWR.n1300 9.3005
R11220 VPWR.n1296 VPWR.n1283 9.3005
R11221 VPWR.n1293 VPWR.n1291 9.3005
R11222 VPWR.n1290 VPWR.n1284 9.3005
R11223 VPWR.n1295 VPWR.n1294 9.3005
R11224 VPWR.n1298 VPWR.n1297 9.3005
R11225 VPWR.n1299 VPWR.n1280 9.3005
R11226 VPWR.n1332 VPWR.n1303 9.3005
R11227 VPWR.n1331 VPWR.n1330 9.3005
R11228 VPWR.n1311 VPWR.n1310 9.3005
R11229 VPWR.n1313 VPWR.n1312 9.3005
R11230 VPWR.n1315 VPWR.n1309 9.3005
R11231 VPWR.n1317 VPWR.n1316 9.3005
R11232 VPWR.n1318 VPWR.n1308 9.3005
R11233 VPWR.n1320 VPWR.n1319 9.3005
R11234 VPWR.n1324 VPWR.n1305 9.3005
R11235 VPWR.n1326 VPWR.n1325 9.3005
R11236 VPWR.n1328 VPWR.n1327 9.3005
R11237 VPWR.n1334 VPWR.n1333 9.3005
R11238 VPWR.n1336 VPWR.n1335 9.3005
R11239 VPWR.n1375 VPWR.n1374 9.3005
R11240 VPWR.n1370 VPWR.n1338 9.3005
R11241 VPWR.n1369 VPWR.n1368 9.3005
R11242 VPWR.n1347 VPWR.n1346 9.3005
R11243 VPWR.n1349 VPWR.n1348 9.3005
R11244 VPWR.n1352 VPWR.n1342 9.3005
R11245 VPWR.n1354 VPWR.n1353 9.3005
R11246 VPWR.n1355 VPWR.n1341 9.3005
R11247 VPWR.n1357 VPWR.n1356 9.3005
R11248 VPWR.n1361 VPWR.n1340 9.3005
R11249 VPWR.n1363 VPWR.n1362 9.3005
R11250 VPWR.n1365 VPWR.n1364 9.3005
R11251 VPWR.n1372 VPWR.n1371 9.3005
R11252 VPWR.n1408 VPWR.n1407 9.3005
R11253 VPWR.n1386 VPWR.n1385 9.3005
R11254 VPWR.n1388 VPWR.n1387 9.3005
R11255 VPWR.n1391 VPWR.n1381 9.3005
R11256 VPWR.n1393 VPWR.n1392 9.3005
R11257 VPWR.n1394 VPWR.n1380 9.3005
R11258 VPWR.n1396 VPWR.n1395 9.3005
R11259 VPWR.n1400 VPWR.n1379 9.3005
R11260 VPWR.n1402 VPWR.n1401 9.3005
R11261 VPWR.n1404 VPWR.n1403 9.3005
R11262 VPWR.n1409 VPWR.n1377 9.3005
R11263 VPWR.n1411 VPWR.n1410 9.3005
R11264 VPWR.n1445 VPWR.n1444 9.3005
R11265 VPWR.n1423 VPWR.n1422 9.3005
R11266 VPWR.n1425 VPWR.n1424 9.3005
R11267 VPWR.n1428 VPWR.n1418 9.3005
R11268 VPWR.n1430 VPWR.n1429 9.3005
R11269 VPWR.n1431 VPWR.n1417 9.3005
R11270 VPWR.n1433 VPWR.n1432 9.3005
R11271 VPWR.n1437 VPWR.n1416 9.3005
R11272 VPWR.n1439 VPWR.n1438 9.3005
R11273 VPWR.n1441 VPWR.n1440 9.3005
R11274 VPWR.n2807 VPWR.n2806 9.3005
R11275 VPWR.n2808 VPWR.n2800 9.3005
R11276 VPWR.n2809 VPWR.n2799 9.3005
R11277 VPWR.n2810 VPWR.n2798 9.3005
R11278 VPWR.n2812 VPWR.n2811 9.3005
R11279 VPWR.n2796 VPWR.n2795 9.3005
R11280 VPWR.n2790 VPWR.n2789 9.3005
R11281 VPWR.n2791 VPWR.n2781 9.3005
R11282 VPWR.n2793 VPWR.n2792 9.3005
R11283 VPWR.n2794 VPWR.n2779 9.3005
R11284 VPWR.n2777 VPWR.n2776 9.3005
R11285 VPWR.n2775 VPWR.n2759 9.3005
R11286 VPWR.n2770 VPWR.n2769 9.3005
R11287 VPWR.n2771 VPWR.n2761 9.3005
R11288 VPWR.n2773 VPWR.n2772 9.3005
R11289 VPWR.n2757 VPWR.n2756 9.3005
R11290 VPWR.n2751 VPWR.n2750 9.3005
R11291 VPWR.n2752 VPWR.n2742 9.3005
R11292 VPWR.n2754 VPWR.n2753 9.3005
R11293 VPWR.n2755 VPWR.n2740 9.3005
R11294 VPWR.n2738 VPWR.n2737 9.3005
R11295 VPWR.n2718 VPWR.n2717 9.3005
R11296 VPWR.n2719 VPWR.n2713 9.3005
R11297 VPWR.n2721 VPWR.n2720 9.3005
R11298 VPWR.n2723 VPWR.n2711 9.3005
R11299 VPWR.n2725 VPWR.n2724 9.3005
R11300 VPWR.n2727 VPWR.n2726 9.3005
R11301 VPWR.n2728 VPWR.n2707 9.3005
R11302 VPWR.n2732 VPWR.n2731 9.3005
R11303 VPWR.n2733 VPWR.n2706 9.3005
R11304 VPWR.n2735 VPWR.n2734 9.3005
R11305 VPWR.n2736 VPWR.n2704 9.3005
R11306 VPWR.n2702 VPWR.n2701 9.3005
R11307 VPWR.n2682 VPWR.n2681 9.3005
R11308 VPWR.n2683 VPWR.n2676 9.3005
R11309 VPWR.n2685 VPWR.n2684 9.3005
R11310 VPWR.n2687 VPWR.n2673 9.3005
R11311 VPWR.n2689 VPWR.n2688 9.3005
R11312 VPWR.n2691 VPWR.n2690 9.3005
R11313 VPWR.n2692 VPWR.n2669 9.3005
R11314 VPWR.n2695 VPWR.n2694 9.3005
R11315 VPWR.n2696 VPWR.n2668 9.3005
R11316 VPWR.n2698 VPWR.n2697 9.3005
R11317 VPWR.n2699 VPWR.n2666 9.3005
R11318 VPWR.n2645 VPWR.n2644 9.3005
R11319 VPWR.n2646 VPWR.n2639 9.3005
R11320 VPWR.n2648 VPWR.n2647 9.3005
R11321 VPWR.n2650 VPWR.n2636 9.3005
R11322 VPWR.n2652 VPWR.n2651 9.3005
R11323 VPWR.n2654 VPWR.n2653 9.3005
R11324 VPWR.n2655 VPWR.n2632 9.3005
R11325 VPWR.n2658 VPWR.n2657 9.3005
R11326 VPWR.n2659 VPWR.n2631 9.3005
R11327 VPWR.n2661 VPWR.n2660 9.3005
R11328 VPWR.n2662 VPWR.n2629 9.3005
R11329 VPWR.n2627 VPWR.n2626 9.3005
R11330 VPWR.n2609 VPWR.n2608 9.3005
R11331 VPWR.n2611 VPWR.n2604 9.3005
R11332 VPWR.n2616 VPWR.n2615 9.3005
R11333 VPWR.n2617 VPWR.n2603 9.3005
R11334 VPWR.n2619 VPWR.n2618 9.3005
R11335 VPWR.n2621 VPWR.n2600 9.3005
R11336 VPWR.n2623 VPWR.n2622 9.3005
R11337 VPWR.n2625 VPWR.n2624 9.3005
R11338 VPWR.n2505 VPWR.n2504 9.3005
R11339 VPWR.n2569 VPWR.n2568 9.3005
R11340 VPWR.n2509 VPWR.n2508 9.3005
R11341 VPWR.n2553 VPWR.n2552 9.3005
R11342 VPWR.n2545 VPWR.n2544 9.3005
R11343 VPWR.n2533 VPWR.n2532 9.3005
R11344 VPWR.n2529 VPWR.n2528 9.3005
R11345 VPWR.n1222 VPWR.n1221 9.3005
R11346 VPWR.n2521 VPWR.n2520 9.3005
R11347 VPWR.n1184 VPWR.n1102 9.3005
R11348 VPWR.n1218 VPWR.n1094 9.3005
R11349 VPWR.n2541 VPWR.n2540 9.3005
R11350 VPWR.n1215 VPWR.n1092 9.3005
R11351 VPWR.n1212 VPWR.n1211 9.3005
R11352 VPWR.n2517 VPWR.n2516 9.3005
R11353 VPWR.n1181 VPWR.n1104 9.3005
R11354 VPWR.n1204 VPWR.n1084 9.3005
R11355 VPWR.n2557 VPWR.n2556 9.3005
R11356 VPWR.n1201 VPWR.n1082 9.3005
R11357 VPWR.n1592 VPWR.n1591 9.3005
R11358 VPWR.n2565 VPWR.n2564 9.3005
R11359 VPWR.n1198 VPWR.n1197 9.3005
R11360 VPWR.n1190 VPWR.n1074 9.3005
R11361 VPWR.n1742 VPWR.n1741 9.3005
R11362 VPWR.n1187 VPWR.n1071 9.3005
R11363 VPWR.n2577 VPWR.n2576 9.3005
R11364 VPWR.n2581 VPWR.n2580 9.3005
R11365 VPWR.n2592 VPWR.n2591 9.3005
R11366 VPWR.n2589 VPWR.n2588 9.3005
R11367 VPWR.n1738 VPWR.n1737 9.3005
R11368 VPWR.n1063 VPWR.n1062 9.3005
R11369 VPWR.n1596 VPWR.n1595 9.3005
R11370 VPWR.n1275 VPWR.n1274 8.28285
R11371 VPWR.n2774 VPWR.n2773 8.28285
R11372 VPWR.n1607 VPWR.n1109 8.25914
R11373 VPWR.n1728 VPWR.n1727 8.25914
R11374 VPWR.n281 VPWR.n113 8.25914
R11375 VPWR.n136 VPWR.n124 8.25914
R11376 VPWR.n1780 VPWR.n1779 7.91351
R11377 VPWR.n1771 VPWR.n1770 7.9105
R11378 VPWR.n1042 VPWR.n1041 7.9105
R11379 VPWR.n1546 VPWR.n1545 7.9105
R11380 VPWR.n1551 VPWR.n1550 7.9105
R11381 VPWR.n1556 VPWR.n1555 7.9105
R11382 VPWR.n1561 VPWR.n1560 7.9105
R11383 VPWR.n1566 VPWR.n1565 7.9105
R11384 VPWR.n1571 VPWR.n1570 7.9105
R11385 VPWR.n1576 VPWR.n1575 7.9105
R11386 VPWR.n1581 VPWR.n1580 7.9105
R11387 VPWR.n1136 VPWR.n1135 7.9105
R11388 VPWR.n1461 VPWR.n1460 7.9105
R11389 VPWR.n1456 VPWR.n1455 7.9105
R11390 VPWR.n1776 VPWR.n1775 7.9105
R11391 VPWR.n1784 VPWR.n1783 7.9105
R11392 VPWR.n282 VPWR.n281 7.9105
R11393 VPWR.n280 VPWR.n279 7.9105
R11394 VPWR.n268 VPWR.n267 7.9105
R11395 VPWR.n256 VPWR.n255 7.9105
R11396 VPWR.n244 VPWR.n243 7.9105
R11397 VPWR.n232 VPWR.n231 7.9105
R11398 VPWR.n220 VPWR.n219 7.9105
R11399 VPWR.n208 VPWR.n207 7.9105
R11400 VPWR.n196 VPWR.n195 7.9105
R11401 VPWR.n184 VPWR.n183 7.9105
R11402 VPWR.n172 VPWR.n171 7.9105
R11403 VPWR.n160 VPWR.n159 7.9105
R11404 VPWR.n148 VPWR.n147 7.9105
R11405 VPWR.n136 VPWR.n135 7.9105
R11406 VPWR.n1727 VPWR.n1726 7.9105
R11407 VPWR.n1715 VPWR.n1714 7.9105
R11408 VPWR.n1701 VPWR.n1068 7.9105
R11409 VPWR.n1690 VPWR.n1689 7.9105
R11410 VPWR.n1688 VPWR.n1687 7.9105
R11411 VPWR.n1674 VPWR.n1079 7.9105
R11412 VPWR.n1663 VPWR.n1662 7.9105
R11413 VPWR.n1661 VPWR.n1660 7.9105
R11414 VPWR.n1647 VPWR.n1089 7.9105
R11415 VPWR.n1636 VPWR.n1635 7.9105
R11416 VPWR.n1634 VPWR.n1633 7.9105
R11417 VPWR.n1620 VPWR.n1099 7.9105
R11418 VPWR.n1609 VPWR.n1608 7.9105
R11419 VPWR.n1607 VPWR.n1606 7.9105
R11420 VPWR.n26 VPWR.n24 7.8627
R11421 VPWR.n7 VPWR.n6 7.56315
R11422 VPWR.n1242 VPWR.n1241 7.56315
R11423 VPWR.n1265 VPWR.n1264 7.56315
R11424 VPWR.n1289 VPWR.n1288 7.56315
R11425 VPWR.n2805 VPWR.n2803 6.4511
R11426 VPWR.n2788 VPWR.n2785 6.4511
R11427 VPWR.n2768 VPWR.n2765 6.4511
R11428 VPWR.n2749 VPWR.n2746 6.4511
R11429 VPWR.n1362 VPWR.n1339 6.4005
R11430 VPWR.n1401 VPWR.n1378 6.4005
R11431 VPWR.n1438 VPWR.n1415 6.4005
R11432 VPWR.n2723 VPWR.n2722 6.4005
R11433 VPWR.n2693 VPWR.n2692 6.4005
R11434 VPWR.n2656 VPWR.n2655 6.4005
R11435 VPWR.n2622 VPWR.n2599 6.4005
R11436 VPWR.n1595 VPWR.n1122 6.04494
R11437 VPWR.n2505 VPWR.n99 6.04494
R11438 VPWR.n1467 VPWR.n1231 6.04494
R11439 VPWR.n351 VPWR.n290 6.04494
R11440 VPWR.n2568 VPWR.n68 6.04494
R11441 VPWR.n1534 VPWR.n1153 6.04494
R11442 VPWR.n348 VPWR.n346 6.04494
R11443 VPWR.n2508 VPWR.n98 6.04494
R11444 VPWR.n965 VPWR.n963 6.04494
R11445 VPWR.n2478 VPWR.n356 6.04494
R11446 VPWR.n2475 VPWR.n357 6.04494
R11447 VPWR.n320 VPWR.n318 6.04494
R11448 VPWR.n2553 VPWR.n75 6.04494
R11449 VPWR.n973 VPWR.n971 6.04494
R11450 VPWR.n2445 VPWR.n369 6.04494
R11451 VPWR.n324 VPWR.n322 6.04494
R11452 VPWR.n2544 VPWR.n80 6.04494
R11453 VPWR.n1890 VPWR.n932 6.04494
R11454 VPWR.n1887 VPWR.n933 6.04494
R11455 VPWR.n1880 VPWR.n936 6.04494
R11456 VPWR.n389 VPWR.n387 6.04494
R11457 VPWR.n393 VPWR.n391 6.04494
R11458 VPWR.n397 VPWR.n395 6.04494
R11459 VPWR.n2455 VPWR.n365 6.04494
R11460 VPWR.n332 VPWR.n330 6.04494
R11461 VPWR.n2532 VPWR.n86 6.04494
R11462 VPWR.n1877 VPWR.n937 6.04494
R11463 VPWR.n405 VPWR.n403 6.04494
R11464 VPWR.n2458 VPWR.n364 6.04494
R11465 VPWR.n336 VPWR.n334 6.04494
R11466 VPWR.n2529 VPWR.n87 6.04494
R11467 VPWR.n2308 VPWR.n481 6.04494
R11468 VPWR.n2311 VPWR.n480 6.04494
R11469 VPWR.n2318 VPWR.n477 6.04494
R11470 VPWR.n2321 VPWR.n476 6.04494
R11471 VPWR.n2331 VPWR.n472 6.04494
R11472 VPWR.n2338 VPWR.n469 6.04494
R11473 VPWR.n2341 VPWR.n468 6.04494
R11474 VPWR.n2348 VPWR.n465 6.04494
R11475 VPWR.n2351 VPWR.n464 6.04494
R11476 VPWR.n2358 VPWR.n461 6.04494
R11477 VPWR.n2361 VPWR.n460 6.04494
R11478 VPWR.n2368 VPWR.n457 6.04494
R11479 VPWR.n2371 VPWR.n456 6.04494
R11480 VPWR.n2378 VPWR.n453 6.04494
R11481 VPWR.n2380 VPWR.n452 6.04494
R11482 VPWR.n2328 VPWR.n473 6.04494
R11483 VPWR.n543 VPWR.n482 6.04494
R11484 VPWR.n540 VPWR.n538 6.04494
R11485 VPWR.n536 VPWR.n534 6.04494
R11486 VPWR.n532 VPWR.n530 6.04494
R11487 VPWR.n524 VPWR.n522 6.04494
R11488 VPWR.n520 VPWR.n518 6.04494
R11489 VPWR.n516 VPWR.n514 6.04494
R11490 VPWR.n512 VPWR.n510 6.04494
R11491 VPWR.n508 VPWR.n506 6.04494
R11492 VPWR.n504 VPWR.n502 6.04494
R11493 VPWR.n500 VPWR.n498 6.04494
R11494 VPWR.n496 VPWR.n494 6.04494
R11495 VPWR.n492 VPWR.n490 6.04494
R11496 VPWR.n488 VPWR.n486 6.04494
R11497 VPWR.n485 VPWR.n483 6.04494
R11498 VPWR.n528 VPWR.n526 6.04494
R11499 VPWR.n2282 VPWR.n548 6.04494
R11500 VPWR.n2279 VPWR.n549 6.04494
R11501 VPWR.n2272 VPWR.n552 6.04494
R11502 VPWR.n2269 VPWR.n553 6.04494
R11503 VPWR.n2259 VPWR.n557 6.04494
R11504 VPWR.n2252 VPWR.n560 6.04494
R11505 VPWR.n2249 VPWR.n561 6.04494
R11506 VPWR.n2242 VPWR.n564 6.04494
R11507 VPWR.n2239 VPWR.n565 6.04494
R11508 VPWR.n2232 VPWR.n568 6.04494
R11509 VPWR.n2229 VPWR.n569 6.04494
R11510 VPWR.n2222 VPWR.n572 6.04494
R11511 VPWR.n2219 VPWR.n573 6.04494
R11512 VPWR.n2212 VPWR.n576 6.04494
R11513 VPWR.n2210 VPWR.n577 6.04494
R11514 VPWR.n2262 VPWR.n556 6.04494
R11515 VPWR.n581 VPWR.n579 6.04494
R11516 VPWR.n585 VPWR.n583 6.04494
R11517 VPWR.n589 VPWR.n587 6.04494
R11518 VPWR.n593 VPWR.n591 6.04494
R11519 VPWR.n601 VPWR.n599 6.04494
R11520 VPWR.n605 VPWR.n603 6.04494
R11521 VPWR.n609 VPWR.n607 6.04494
R11522 VPWR.n613 VPWR.n611 6.04494
R11523 VPWR.n617 VPWR.n615 6.04494
R11524 VPWR.n621 VPWR.n619 6.04494
R11525 VPWR.n625 VPWR.n623 6.04494
R11526 VPWR.n629 VPWR.n627 6.04494
R11527 VPWR.n633 VPWR.n631 6.04494
R11528 VPWR.n637 VPWR.n635 6.04494
R11529 VPWR.n639 VPWR.n578 6.04494
R11530 VPWR.n597 VPWR.n595 6.04494
R11531 VPWR.n2112 VPWR.n673 6.04494
R11532 VPWR.n2115 VPWR.n672 6.04494
R11533 VPWR.n2122 VPWR.n669 6.04494
R11534 VPWR.n2125 VPWR.n668 6.04494
R11535 VPWR.n2135 VPWR.n664 6.04494
R11536 VPWR.n2142 VPWR.n661 6.04494
R11537 VPWR.n2145 VPWR.n660 6.04494
R11538 VPWR.n2152 VPWR.n657 6.04494
R11539 VPWR.n2155 VPWR.n656 6.04494
R11540 VPWR.n2162 VPWR.n653 6.04494
R11541 VPWR.n2165 VPWR.n652 6.04494
R11542 VPWR.n2172 VPWR.n649 6.04494
R11543 VPWR.n2175 VPWR.n648 6.04494
R11544 VPWR.n2182 VPWR.n645 6.04494
R11545 VPWR.n2184 VPWR.n644 6.04494
R11546 VPWR.n2132 VPWR.n665 6.04494
R11547 VPWR.n735 VPWR.n674 6.04494
R11548 VPWR.n732 VPWR.n730 6.04494
R11549 VPWR.n728 VPWR.n726 6.04494
R11550 VPWR.n724 VPWR.n722 6.04494
R11551 VPWR.n716 VPWR.n714 6.04494
R11552 VPWR.n712 VPWR.n710 6.04494
R11553 VPWR.n708 VPWR.n706 6.04494
R11554 VPWR.n704 VPWR.n702 6.04494
R11555 VPWR.n700 VPWR.n698 6.04494
R11556 VPWR.n696 VPWR.n694 6.04494
R11557 VPWR.n692 VPWR.n690 6.04494
R11558 VPWR.n688 VPWR.n686 6.04494
R11559 VPWR.n684 VPWR.n682 6.04494
R11560 VPWR.n680 VPWR.n678 6.04494
R11561 VPWR.n677 VPWR.n675 6.04494
R11562 VPWR.n720 VPWR.n718 6.04494
R11563 VPWR.n2086 VPWR.n740 6.04494
R11564 VPWR.n2083 VPWR.n741 6.04494
R11565 VPWR.n2076 VPWR.n744 6.04494
R11566 VPWR.n2073 VPWR.n745 6.04494
R11567 VPWR.n2063 VPWR.n749 6.04494
R11568 VPWR.n2056 VPWR.n752 6.04494
R11569 VPWR.n2053 VPWR.n753 6.04494
R11570 VPWR.n2046 VPWR.n756 6.04494
R11571 VPWR.n2043 VPWR.n757 6.04494
R11572 VPWR.n2036 VPWR.n760 6.04494
R11573 VPWR.n2033 VPWR.n761 6.04494
R11574 VPWR.n2026 VPWR.n764 6.04494
R11575 VPWR.n2023 VPWR.n765 6.04494
R11576 VPWR.n2016 VPWR.n768 6.04494
R11577 VPWR.n2014 VPWR.n769 6.04494
R11578 VPWR.n2066 VPWR.n748 6.04494
R11579 VPWR.n773 VPWR.n771 6.04494
R11580 VPWR.n777 VPWR.n775 6.04494
R11581 VPWR.n781 VPWR.n779 6.04494
R11582 VPWR.n785 VPWR.n783 6.04494
R11583 VPWR.n793 VPWR.n791 6.04494
R11584 VPWR.n797 VPWR.n795 6.04494
R11585 VPWR.n801 VPWR.n799 6.04494
R11586 VPWR.n805 VPWR.n803 6.04494
R11587 VPWR.n809 VPWR.n807 6.04494
R11588 VPWR.n813 VPWR.n811 6.04494
R11589 VPWR.n817 VPWR.n815 6.04494
R11590 VPWR.n821 VPWR.n819 6.04494
R11591 VPWR.n825 VPWR.n823 6.04494
R11592 VPWR.n829 VPWR.n827 6.04494
R11593 VPWR.n831 VPWR.n770 6.04494
R11594 VPWR.n789 VPWR.n787 6.04494
R11595 VPWR.n1916 VPWR.n865 6.04494
R11596 VPWR.n1919 VPWR.n864 6.04494
R11597 VPWR.n1926 VPWR.n861 6.04494
R11598 VPWR.n1929 VPWR.n860 6.04494
R11599 VPWR.n1939 VPWR.n856 6.04494
R11600 VPWR.n1946 VPWR.n853 6.04494
R11601 VPWR.n1949 VPWR.n852 6.04494
R11602 VPWR.n1956 VPWR.n849 6.04494
R11603 VPWR.n1959 VPWR.n848 6.04494
R11604 VPWR.n1966 VPWR.n845 6.04494
R11605 VPWR.n1969 VPWR.n844 6.04494
R11606 VPWR.n1976 VPWR.n841 6.04494
R11607 VPWR.n1979 VPWR.n840 6.04494
R11608 VPWR.n1986 VPWR.n837 6.04494
R11609 VPWR.n1988 VPWR.n836 6.04494
R11610 VPWR.n1936 VPWR.n857 6.04494
R11611 VPWR.n927 VPWR.n866 6.04494
R11612 VPWR.n924 VPWR.n922 6.04494
R11613 VPWR.n920 VPWR.n918 6.04494
R11614 VPWR.n916 VPWR.n914 6.04494
R11615 VPWR.n908 VPWR.n906 6.04494
R11616 VPWR.n904 VPWR.n902 6.04494
R11617 VPWR.n900 VPWR.n898 6.04494
R11618 VPWR.n896 VPWR.n894 6.04494
R11619 VPWR.n892 VPWR.n890 6.04494
R11620 VPWR.n888 VPWR.n886 6.04494
R11621 VPWR.n884 VPWR.n882 6.04494
R11622 VPWR.n880 VPWR.n878 6.04494
R11623 VPWR.n876 VPWR.n874 6.04494
R11624 VPWR.n872 VPWR.n870 6.04494
R11625 VPWR.n869 VPWR.n867 6.04494
R11626 VPWR.n912 VPWR.n910 6.04494
R11627 VPWR.n1870 VPWR.n940 6.04494
R11628 VPWR.n981 VPWR.n979 6.04494
R11629 VPWR.n1494 VPWR.n1227 6.04494
R11630 VPWR.n1221 VPWR.n1179 6.04494
R11631 VPWR.n401 VPWR.n399 6.04494
R11632 VPWR.n2465 VPWR.n361 6.04494
R11633 VPWR.n340 VPWR.n338 6.04494
R11634 VPWR.n2520 VPWR.n92 6.04494
R11635 VPWR.n977 VPWR.n975 6.04494
R11636 VPWR.n1491 VPWR.n1485 6.04494
R11637 VPWR.n1184 VPWR.n1183 6.04494
R11638 VPWR.n1867 VPWR.n941 6.04494
R11639 VPWR.n985 VPWR.n983 6.04494
R11640 VPWR.n1505 VPWR.n1173 6.04494
R11641 VPWR.n1218 VPWR.n1217 6.04494
R11642 VPWR.n409 VPWR.n407 6.04494
R11643 VPWR.n417 VPWR.n415 6.04494
R11644 VPWR.n421 VPWR.n419 6.04494
R11645 VPWR.n425 VPWR.n423 6.04494
R11646 VPWR.n429 VPWR.n427 6.04494
R11647 VPWR.n433 VPWR.n431 6.04494
R11648 VPWR.n437 VPWR.n435 6.04494
R11649 VPWR.n441 VPWR.n439 6.04494
R11650 VPWR.n445 VPWR.n443 6.04494
R11651 VPWR.n447 VPWR.n386 6.04494
R11652 VPWR.n413 VPWR.n411 6.04494
R11653 VPWR.n2448 VPWR.n368 6.04494
R11654 VPWR.n328 VPWR.n326 6.04494
R11655 VPWR.n2541 VPWR.n81 6.04494
R11656 VPWR.n989 VPWR.n987 6.04494
R11657 VPWR.n1508 VPWR.n1169 6.04494
R11658 VPWR.n1215 VPWR.n1214 6.04494
R11659 VPWR.n1860 VPWR.n944 6.04494
R11660 VPWR.n1850 VPWR.n948 6.04494
R11661 VPWR.n1847 VPWR.n949 6.04494
R11662 VPWR.n1840 VPWR.n952 6.04494
R11663 VPWR.n1837 VPWR.n953 6.04494
R11664 VPWR.n1830 VPWR.n956 6.04494
R11665 VPWR.n1827 VPWR.n957 6.04494
R11666 VPWR.n1820 VPWR.n960 6.04494
R11667 VPWR.n1818 VPWR.n961 6.04494
R11668 VPWR.n1857 VPWR.n945 6.04494
R11669 VPWR.n993 VPWR.n991 6.04494
R11670 VPWR.n1519 VPWR.n1163 6.04494
R11671 VPWR.n1212 VPWR.n1206 6.04494
R11672 VPWR.n2468 VPWR.n360 6.04494
R11673 VPWR.n344 VPWR.n342 6.04494
R11674 VPWR.n2517 VPWR.n93 6.04494
R11675 VPWR.n1480 VPWR.n1479 6.04494
R11676 VPWR.n1181 VPWR.n1180 6.04494
R11677 VPWR.n997 VPWR.n995 6.04494
R11678 VPWR.n1522 VPWR.n1159 6.04494
R11679 VPWR.n1204 VPWR.n1203 6.04494
R11680 VPWR.n2438 VPWR.n372 6.04494
R11681 VPWR.n2428 VPWR.n376 6.04494
R11682 VPWR.n2425 VPWR.n377 6.04494
R11683 VPWR.n2418 VPWR.n380 6.04494
R11684 VPWR.n2415 VPWR.n381 6.04494
R11685 VPWR.n2408 VPWR.n384 6.04494
R11686 VPWR.n2406 VPWR.n385 6.04494
R11687 VPWR.n2435 VPWR.n373 6.04494
R11688 VPWR.n316 VPWR.n314 6.04494
R11689 VPWR.n2556 VPWR.n74 6.04494
R11690 VPWR.n1537 VPWR.n1149 6.04494
R11691 VPWR.n1201 VPWR.n1200 6.04494
R11692 VPWR.n1001 VPWR.n999 6.04494
R11693 VPWR.n1005 VPWR.n1003 6.04494
R11694 VPWR.n1009 VPWR.n1007 6.04494
R11695 VPWR.n1013 VPWR.n1011 6.04494
R11696 VPWR.n1017 VPWR.n1015 6.04494
R11697 VPWR.n1021 VPWR.n1019 6.04494
R11698 VPWR.n1023 VPWR.n962 6.04494
R11699 VPWR.n969 VPWR.n967 6.04494
R11700 VPWR.n1474 VPWR.n1472 6.04494
R11701 VPWR.n1592 VPWR.n1123 6.04494
R11702 VPWR.n312 VPWR.n310 6.04494
R11703 VPWR.n2565 VPWR.n69 6.04494
R11704 VPWR.n1198 VPWR.n1192 6.04494
R11705 VPWR.n1762 VPWR.n1049 6.04494
R11706 VPWR.n1190 VPWR.n1189 6.04494
R11707 VPWR.n308 VPWR.n306 6.04494
R11708 VPWR.n304 VPWR.n302 6.04494
R11709 VPWR.n296 VPWR.n294 6.04494
R11710 VPWR.n293 VPWR.n291 6.04494
R11711 VPWR.n300 VPWR.n298 6.04494
R11712 VPWR.n1741 VPWR.n1058 6.04494
R11713 VPWR.n1750 VPWR.n1748 6.04494
R11714 VPWR.n1790 VPWR.n1036 6.04494
R11715 VPWR.n1792 VPWR.n1032 6.04494
R11716 VPWR.n1759 VPWR.n1053 6.04494
R11717 VPWR.n1187 VPWR.n1186 6.04494
R11718 VPWR.n2577 VPWR.n63 6.04494
R11719 VPWR.n2580 VPWR.n62 6.04494
R11720 VPWR.n2589 VPWR.n57 6.04494
R11721 VPWR.n2591 VPWR.n56 6.04494
R11722 VPWR.n1738 VPWR.n1059 6.04494
R11723 VPWR.n1062 VPWR.n1061 6.04494
R11724 VPWR.n2785 VPWR.n2784 5.39628
R11725 VPWR.n2765 VPWR.n2764 5.39628
R11726 VPWR.n2746 VPWR.n2745 5.39628
R11727 VPWR.n54 VPWR 4.72593
R11728 VPWR.n52 VPWR 4.72593
R11729 VPWR.n50 VPWR 4.72593
R11730 VPWR.n48 VPWR 4.72593
R11731 VPWR.n46 VPWR 4.72593
R11732 VPWR.n44 VPWR 4.72593
R11733 VPWR.n42 VPWR 4.72593
R11734 VPWR.n40 VPWR 4.72593
R11735 VPWR.n38 VPWR 4.72593
R11736 VPWR.n36 VPWR 4.72593
R11737 VPWR.n34 VPWR 4.72593
R11738 VPWR.n32 VPWR 4.72593
R11739 VPWR.n30 VPWR 4.72593
R11740 VPWR.n28 VPWR 4.72593
R11741 VPWR.n26 VPWR 4.72593
R11742 VPWR.n1446 VPWR.n1445 4.55954
R11743 VPWR.n2571 VPWR.n2570 4.5005
R11744 VPWR.n2511 VPWR.n2510 4.5005
R11745 VPWR.n2551 VPWR.n2550 4.5005
R11746 VPWR.n319 VPWR.n77 4.5005
R11747 VPWR.n2547 VPWR.n2546 4.5005
R11748 VPWR.n323 VPWR.n78 4.5005
R11749 VPWR.n2535 VPWR.n2534 4.5005
R11750 VPWR.n331 VPWR.n84 4.5005
R11751 VPWR.n2454 VPWR.n2453 4.5005
R11752 VPWR.n2527 VPWR.n2526 4.5005
R11753 VPWR.n335 VPWR.n89 4.5005
R11754 VPWR.n2460 VPWR.n2459 4.5005
R11755 VPWR.n1498 VPWR.n1223 4.5005
R11756 VPWR.n1497 VPWR.n1495 4.5005
R11757 VPWR.n980 VPWR.n939 4.5005
R11758 VPWR.n1872 VPWR.n1871 4.5005
R11759 VPWR.n911 VPWR.n858 4.5005
R11760 VPWR.n1935 VPWR.n1934 4.5005
R11761 VPWR.n788 VPWR.n747 4.5005
R11762 VPWR.n2068 VPWR.n2067 4.5005
R11763 VPWR.n719 VPWR.n666 4.5005
R11764 VPWR.n2131 VPWR.n2130 4.5005
R11765 VPWR.n596 VPWR.n555 4.5005
R11766 VPWR.n2264 VPWR.n2263 4.5005
R11767 VPWR.n527 VPWR.n474 4.5005
R11768 VPWR.n2327 VPWR.n2326 4.5005
R11769 VPWR.n404 VPWR.n363 4.5005
R11770 VPWR.n2523 VPWR.n2522 4.5005
R11771 VPWR.n339 VPWR.n90 4.5005
R11772 VPWR.n2464 VPWR.n2463 4.5005
R11773 VPWR.n400 VPWR.n362 4.5005
R11774 VPWR.n2323 VPWR.n2322 4.5005
R11775 VPWR.n531 VPWR.n475 4.5005
R11776 VPWR.n2268 VPWR.n2267 4.5005
R11777 VPWR.n592 VPWR.n554 4.5005
R11778 VPWR.n2127 VPWR.n2126 4.5005
R11779 VPWR.n723 VPWR.n667 4.5005
R11780 VPWR.n2072 VPWR.n2071 4.5005
R11781 VPWR.n784 VPWR.n746 4.5005
R11782 VPWR.n1931 VPWR.n1930 4.5005
R11783 VPWR.n915 VPWR.n859 4.5005
R11784 VPWR.n1488 VPWR.n1486 4.5005
R11785 VPWR.n1490 VPWR.n1489 4.5005
R11786 VPWR.n976 VPWR.n938 4.5005
R11787 VPWR.n1876 VPWR.n1875 4.5005
R11788 VPWR.n1501 VPWR.n1174 4.5005
R11789 VPWR.n1504 VPWR.n1503 4.5005
R11790 VPWR.n984 VPWR.n942 4.5005
R11791 VPWR.n1866 VPWR.n1865 4.5005
R11792 VPWR.n907 VPWR.n855 4.5005
R11793 VPWR.n1941 VPWR.n1940 4.5005
R11794 VPWR.n792 VPWR.n750 4.5005
R11795 VPWR.n2062 VPWR.n2061 4.5005
R11796 VPWR.n715 VPWR.n663 4.5005
R11797 VPWR.n2137 VPWR.n2136 4.5005
R11798 VPWR.n600 VPWR.n558 4.5005
R11799 VPWR.n2258 VPWR.n2257 4.5005
R11800 VPWR.n523 VPWR.n471 4.5005
R11801 VPWR.n2333 VPWR.n2332 4.5005
R11802 VPWR.n408 VPWR.n366 4.5005
R11803 VPWR.n2539 VPWR.n2538 4.5005
R11804 VPWR.n327 VPWR.n83 4.5005
R11805 VPWR.n2450 VPWR.n2449 4.5005
R11806 VPWR.n412 VPWR.n367 4.5005
R11807 VPWR.n2337 VPWR.n2336 4.5005
R11808 VPWR.n519 VPWR.n470 4.5005
R11809 VPWR.n2254 VPWR.n2253 4.5005
R11810 VPWR.n604 VPWR.n559 4.5005
R11811 VPWR.n2141 VPWR.n2140 4.5005
R11812 VPWR.n711 VPWR.n662 4.5005
R11813 VPWR.n2058 VPWR.n2057 4.5005
R11814 VPWR.n796 VPWR.n751 4.5005
R11815 VPWR.n1945 VPWR.n1944 4.5005
R11816 VPWR.n903 VPWR.n854 4.5005
R11817 VPWR.n1512 VPWR.n1165 4.5005
R11818 VPWR.n1511 VPWR.n1509 4.5005
R11819 VPWR.n988 VPWR.n943 4.5005
R11820 VPWR.n1862 VPWR.n1861 4.5005
R11821 VPWR.n1515 VPWR.n1164 4.5005
R11822 VPWR.n1518 VPWR.n1517 4.5005
R11823 VPWR.n992 VPWR.n946 4.5005
R11824 VPWR.n1856 VPWR.n1855 4.5005
R11825 VPWR.n899 VPWR.n851 4.5005
R11826 VPWR.n1951 VPWR.n1950 4.5005
R11827 VPWR.n800 VPWR.n754 4.5005
R11828 VPWR.n2052 VPWR.n2051 4.5005
R11829 VPWR.n707 VPWR.n659 4.5005
R11830 VPWR.n2147 VPWR.n2146 4.5005
R11831 VPWR.n608 VPWR.n562 4.5005
R11832 VPWR.n2248 VPWR.n2247 4.5005
R11833 VPWR.n515 VPWR.n467 4.5005
R11834 VPWR.n2343 VPWR.n2342 4.5005
R11835 VPWR.n416 VPWR.n370 4.5005
R11836 VPWR.n2444 VPWR.n2443 4.5005
R11837 VPWR.n2515 VPWR.n2514 4.5005
R11838 VPWR.n343 VPWR.n95 4.5005
R11839 VPWR.n2470 VPWR.n2469 4.5005
R11840 VPWR.n396 VPWR.n359 4.5005
R11841 VPWR.n2317 VPWR.n2316 4.5005
R11842 VPWR.n535 VPWR.n478 4.5005
R11843 VPWR.n2274 VPWR.n2273 4.5005
R11844 VPWR.n588 VPWR.n551 4.5005
R11845 VPWR.n2121 VPWR.n2120 4.5005
R11846 VPWR.n727 VPWR.n670 4.5005
R11847 VPWR.n2078 VPWR.n2077 4.5005
R11848 VPWR.n780 VPWR.n743 4.5005
R11849 VPWR.n1925 VPWR.n1924 4.5005
R11850 VPWR.n919 VPWR.n862 4.5005
R11851 VPWR.n1882 VPWR.n1881 4.5005
R11852 VPWR.n1586 VPWR.n1129 4.5005
R11853 VPWR.n1585 VPWR.n1130 4.5005
R11854 VPWR.n972 VPWR.n935 4.5005
R11855 VPWR.n1526 VPWR.n1155 4.5005
R11856 VPWR.n1525 VPWR.n1523 4.5005
R11857 VPWR.n996 VPWR.n947 4.5005
R11858 VPWR.n1852 VPWR.n1851 4.5005
R11859 VPWR.n895 VPWR.n850 4.5005
R11860 VPWR.n1955 VPWR.n1954 4.5005
R11861 VPWR.n804 VPWR.n755 4.5005
R11862 VPWR.n2048 VPWR.n2047 4.5005
R11863 VPWR.n703 VPWR.n658 4.5005
R11864 VPWR.n2151 VPWR.n2150 4.5005
R11865 VPWR.n612 VPWR.n563 4.5005
R11866 VPWR.n2244 VPWR.n2243 4.5005
R11867 VPWR.n511 VPWR.n466 4.5005
R11868 VPWR.n2347 VPWR.n2346 4.5005
R11869 VPWR.n420 VPWR.n371 4.5005
R11870 VPWR.n2440 VPWR.n2439 4.5005
R11871 VPWR.n2559 VPWR.n2558 4.5005
R11872 VPWR.n315 VPWR.n72 4.5005
R11873 VPWR.n2434 VPWR.n2433 4.5005
R11874 VPWR.n424 VPWR.n374 4.5005
R11875 VPWR.n2353 VPWR.n2352 4.5005
R11876 VPWR.n507 VPWR.n463 4.5005
R11877 VPWR.n2238 VPWR.n2237 4.5005
R11878 VPWR.n616 VPWR.n566 4.5005
R11879 VPWR.n2157 VPWR.n2156 4.5005
R11880 VPWR.n699 VPWR.n655 4.5005
R11881 VPWR.n2042 VPWR.n2041 4.5005
R11882 VPWR.n808 VPWR.n758 4.5005
R11883 VPWR.n1961 VPWR.n1960 4.5005
R11884 VPWR.n891 VPWR.n847 4.5005
R11885 VPWR.n1846 VPWR.n1845 4.5005
R11886 VPWR.n1145 VPWR.n1144 4.5005
R11887 VPWR.n1539 VPWR.n1538 4.5005
R11888 VPWR.n1000 VPWR.n950 4.5005
R11889 VPWR.n1590 VPWR.n1589 4.5005
R11890 VPWR.n1473 VPWR.n1128 4.5005
R11891 VPWR.n968 VPWR.n934 4.5005
R11892 VPWR.n1886 VPWR.n1885 4.5005
R11893 VPWR.n923 VPWR.n863 4.5005
R11894 VPWR.n1921 VPWR.n1920 4.5005
R11895 VPWR.n776 VPWR.n742 4.5005
R11896 VPWR.n2082 VPWR.n2081 4.5005
R11897 VPWR.n731 VPWR.n671 4.5005
R11898 VPWR.n2117 VPWR.n2116 4.5005
R11899 VPWR.n584 VPWR.n550 4.5005
R11900 VPWR.n2278 VPWR.n2277 4.5005
R11901 VPWR.n539 VPWR.n479 4.5005
R11902 VPWR.n2313 VPWR.n2312 4.5005
R11903 VPWR.n392 VPWR.n358 4.5005
R11904 VPWR.n2474 VPWR.n2473 4.5005
R11905 VPWR.n347 VPWR.n96 4.5005
R11906 VPWR.n2563 VPWR.n2562 4.5005
R11907 VPWR.n311 VPWR.n71 4.5005
R11908 VPWR.n2430 VPWR.n2429 4.5005
R11909 VPWR.n428 VPWR.n375 4.5005
R11910 VPWR.n2357 VPWR.n2356 4.5005
R11911 VPWR.n503 VPWR.n462 4.5005
R11912 VPWR.n2234 VPWR.n2233 4.5005
R11913 VPWR.n620 VPWR.n567 4.5005
R11914 VPWR.n2161 VPWR.n2160 4.5005
R11915 VPWR.n695 VPWR.n654 4.5005
R11916 VPWR.n2038 VPWR.n2037 4.5005
R11917 VPWR.n812 VPWR.n759 4.5005
R11918 VPWR.n1965 VPWR.n1964 4.5005
R11919 VPWR.n887 VPWR.n846 4.5005
R11920 VPWR.n1842 VPWR.n1841 4.5005
R11921 VPWR.n1004 VPWR.n951 4.5005
R11922 VPWR.n1531 VPWR.n1154 4.5005
R11923 VPWR.n1533 VPWR.n1532 4.5005
R11924 VPWR.n1073 VPWR.n1045 4.5005
R11925 VPWR.n1764 VPWR.n1763 4.5005
R11926 VPWR.n1008 VPWR.n954 4.5005
R11927 VPWR.n1836 VPWR.n1835 4.5005
R11928 VPWR.n883 VPWR.n843 4.5005
R11929 VPWR.n1971 VPWR.n1970 4.5005
R11930 VPWR.n816 VPWR.n762 4.5005
R11931 VPWR.n2032 VPWR.n2031 4.5005
R11932 VPWR.n691 VPWR.n651 4.5005
R11933 VPWR.n2167 VPWR.n2166 4.5005
R11934 VPWR.n624 VPWR.n570 4.5005
R11935 VPWR.n2228 VPWR.n2227 4.5005
R11936 VPWR.n499 VPWR.n459 4.5005
R11937 VPWR.n2363 VPWR.n2362 4.5005
R11938 VPWR.n432 VPWR.n378 4.5005
R11939 VPWR.n2424 VPWR.n2423 4.5005
R11940 VPWR.n307 VPWR.n66 4.5005
R11941 VPWR.n299 VPWR.n60 4.5005
R11942 VPWR.n2414 VPWR.n2413 4.5005
R11943 VPWR.n440 VPWR.n382 4.5005
R11944 VPWR.n2373 VPWR.n2372 4.5005
R11945 VPWR.n491 VPWR.n455 4.5005
R11946 VPWR.n2218 VPWR.n2217 4.5005
R11947 VPWR.n632 VPWR.n574 4.5005
R11948 VPWR.n2177 VPWR.n2176 4.5005
R11949 VPWR.n683 VPWR.n647 4.5005
R11950 VPWR.n2022 VPWR.n2021 4.5005
R11951 VPWR.n824 VPWR.n766 4.5005
R11952 VPWR.n1981 VPWR.n1980 4.5005
R11953 VPWR.n875 VPWR.n839 4.5005
R11954 VPWR.n1826 VPWR.n1825 4.5005
R11955 VPWR.n1016 VPWR.n958 4.5005
R11956 VPWR.n1753 VPWR.n1743 4.5005
R11957 VPWR.n1752 VPWR.n1751 4.5005
R11958 VPWR.n1756 VPWR.n1054 4.5005
R11959 VPWR.n1758 VPWR.n1757 4.5005
R11960 VPWR.n1012 VPWR.n955 4.5005
R11961 VPWR.n1832 VPWR.n1831 4.5005
R11962 VPWR.n879 VPWR.n842 4.5005
R11963 VPWR.n1975 VPWR.n1974 4.5005
R11964 VPWR.n820 VPWR.n763 4.5005
R11965 VPWR.n2028 VPWR.n2027 4.5005
R11966 VPWR.n687 VPWR.n650 4.5005
R11967 VPWR.n2171 VPWR.n2170 4.5005
R11968 VPWR.n628 VPWR.n571 4.5005
R11969 VPWR.n2224 VPWR.n2223 4.5005
R11970 VPWR.n495 VPWR.n458 4.5005
R11971 VPWR.n2367 VPWR.n2366 4.5005
R11972 VPWR.n436 VPWR.n379 4.5005
R11973 VPWR.n2420 VPWR.n2419 4.5005
R11974 VPWR.n303 VPWR.n65 4.5005
R11975 VPWR.n2575 VPWR.n2574 4.5005
R11976 VPWR.n2583 VPWR.n2582 4.5005
R11977 VPWR.n2587 VPWR.n2586 4.5005
R11978 VPWR.n295 VPWR.n59 4.5005
R11979 VPWR.n2410 VPWR.n2409 4.5005
R11980 VPWR.n444 VPWR.n383 4.5005
R11981 VPWR.n2377 VPWR.n2376 4.5005
R11982 VPWR.n487 VPWR.n454 4.5005
R11983 VPWR.n2214 VPWR.n2213 4.5005
R11984 VPWR.n636 VPWR.n575 4.5005
R11985 VPWR.n2181 VPWR.n2180 4.5005
R11986 VPWR.n679 VPWR.n646 4.5005
R11987 VPWR.n2018 VPWR.n2017 4.5005
R11988 VPWR.n828 VPWR.n767 4.5005
R11989 VPWR.n1985 VPWR.n1984 4.5005
R11990 VPWR.n871 VPWR.n838 4.5005
R11991 VPWR.n1822 VPWR.n1821 4.5005
R11992 VPWR.n1020 VPWR.n959 4.5005
R11993 VPWR.n1789 VPWR.n1788 4.5005
R11994 VPWR.n1736 VPWR.n1037 4.5005
R11995 VPWR.n1232 VPWR.n1121 4.5005
R11996 VPWR.n1466 VPWR.n1465 4.5005
R11997 VPWR.n964 VPWR.n931 4.5005
R11998 VPWR.n1892 VPWR.n1891 4.5005
R11999 VPWR.n929 VPWR.n928 4.5005
R12000 VPWR.n1915 VPWR.n1914 4.5005
R12001 VPWR.n772 VPWR.n739 4.5005
R12002 VPWR.n2088 VPWR.n2087 4.5005
R12003 VPWR.n737 VPWR.n736 4.5005
R12004 VPWR.n2111 VPWR.n2110 4.5005
R12005 VPWR.n580 VPWR.n547 4.5005
R12006 VPWR.n2284 VPWR.n2283 4.5005
R12007 VPWR.n545 VPWR.n544 4.5005
R12008 VPWR.n2307 VPWR.n2306 4.5005
R12009 VPWR.n388 VPWR.n355 4.5005
R12010 VPWR.n2480 VPWR.n2479 4.5005
R12011 VPWR.n353 VPWR.n352 4.5005
R12012 VPWR.n2503 VPWR.n2502 4.5005
R12013 VPWR.n2594 VPWR.n2593 4.5005
R12014 VPWR.n292 VPWR.n22 4.5005
R12015 VPWR.n2405 VPWR.n2404 4.5005
R12016 VPWR.n449 VPWR.n448 4.5005
R12017 VPWR.n2382 VPWR.n2381 4.5005
R12018 VPWR.n484 VPWR.n451 4.5005
R12019 VPWR.n2209 VPWR.n2208 4.5005
R12020 VPWR.n641 VPWR.n640 4.5005
R12021 VPWR.n2186 VPWR.n2185 4.5005
R12022 VPWR.n676 VPWR.n643 4.5005
R12023 VPWR.n2013 VPWR.n2012 4.5005
R12024 VPWR.n833 VPWR.n832 4.5005
R12025 VPWR.n1990 VPWR.n1989 4.5005
R12026 VPWR.n868 VPWR.n835 4.5005
R12027 VPWR.n1817 VPWR.n1816 4.5005
R12028 VPWR.n1025 VPWR.n1024 4.5005
R12029 VPWR.n1794 VPWR.n1793 4.5005
R12030 VPWR.n1060 VPWR.n1028 4.5005
R12031 VPWR.n2628 VPWR 4.49965
R12032 VPWR.n19 VPWR.n18 4.20017
R12033 VPWR.n1255 VPWR.n1254 4.20017
R12034 VPWR.n1279 VPWR.n1278 4.20017
R12035 VPWR.n1302 VPWR.n1301 4.20017
R12036 VPWR.n1337 VPWR.n1336 4.20017
R12037 VPWR.n1376 VPWR.n1375 4.20017
R12038 VPWR.n1414 VPWR.n1413 4.20017
R12039 VPWR.n2813 VPWR 4.14027
R12040 VPWR.n2797 VPWR 4.14027
R12041 VPWR.n2778 VPWR 4.14027
R12042 VPWR.n2758 VPWR 4.14027
R12043 VPWR.n2739 VPWR 4.14027
R12044 VPWR.n2703 VPWR 4.14027
R12045 VPWR.n2665 VPWR 4.14027
R12046 VPWR.n55 VPWR.n54 4.0005
R12047 VPWR.n2716 VPWR.n2713 3.76521
R12048 VPWR.n2680 VPWR.n2676 3.76521
R12049 VPWR.n2643 VPWR.n2639 3.76521
R12050 VPWR.n2611 VPWR.n2610 3.76521
R12051 VPWR.n1906 VPWR.n858 3.4105
R12052 VPWR.n1934 VPWR.n1933 3.4105
R12053 VPWR.n1997 VPWR.n747 3.4105
R12054 VPWR.n2069 VPWR.n2068 3.4105
R12055 VPWR.n2102 VPWR.n666 3.4105
R12056 VPWR.n2130 VPWR.n2129 3.4105
R12057 VPWR.n2193 VPWR.n555 3.4105
R12058 VPWR.n2265 VPWR.n2264 3.4105
R12059 VPWR.n2298 VPWR.n474 3.4105
R12060 VPWR.n2326 VPWR.n2325 3.4105
R12061 VPWR.n2389 VPWR.n363 3.4105
R12062 VPWR.n2388 VPWR.n362 3.4105
R12063 VPWR.n2324 VPWR.n2323 3.4105
R12064 VPWR.n2299 VPWR.n475 3.4105
R12065 VPWR.n2267 VPWR.n2266 3.4105
R12066 VPWR.n2192 VPWR.n554 3.4105
R12067 VPWR.n2128 VPWR.n2127 3.4105
R12068 VPWR.n2103 VPWR.n667 3.4105
R12069 VPWR.n2071 VPWR.n2070 3.4105
R12070 VPWR.n1996 VPWR.n746 3.4105
R12071 VPWR.n1932 VPWR.n1931 3.4105
R12072 VPWR.n1907 VPWR.n859 3.4105
R12073 VPWR.n1875 VPWR.n1874 3.4105
R12074 VPWR.n1873 VPWR.n1872 3.4105
R12075 VPWR.n1865 VPWR.n1864 3.4105
R12076 VPWR.n1905 VPWR.n855 3.4105
R12077 VPWR.n1942 VPWR.n1941 3.4105
R12078 VPWR.n1998 VPWR.n750 3.4105
R12079 VPWR.n2061 VPWR.n2060 3.4105
R12080 VPWR.n2101 VPWR.n663 3.4105
R12081 VPWR.n2138 VPWR.n2137 3.4105
R12082 VPWR.n2194 VPWR.n558 3.4105
R12083 VPWR.n2257 VPWR.n2256 3.4105
R12084 VPWR.n2297 VPWR.n471 3.4105
R12085 VPWR.n2334 VPWR.n2333 3.4105
R12086 VPWR.n2390 VPWR.n366 3.4105
R12087 VPWR.n2391 VPWR.n367 3.4105
R12088 VPWR.n2336 VPWR.n2335 3.4105
R12089 VPWR.n2296 VPWR.n470 3.4105
R12090 VPWR.n2255 VPWR.n2254 3.4105
R12091 VPWR.n2195 VPWR.n559 3.4105
R12092 VPWR.n2140 VPWR.n2139 3.4105
R12093 VPWR.n2100 VPWR.n662 3.4105
R12094 VPWR.n2059 VPWR.n2058 3.4105
R12095 VPWR.n1999 VPWR.n751 3.4105
R12096 VPWR.n1944 VPWR.n1943 3.4105
R12097 VPWR.n1904 VPWR.n854 3.4105
R12098 VPWR.n1863 VPWR.n1862 3.4105
R12099 VPWR.n1855 VPWR.n1854 3.4105
R12100 VPWR.n1903 VPWR.n851 3.4105
R12101 VPWR.n1952 VPWR.n1951 3.4105
R12102 VPWR.n2000 VPWR.n754 3.4105
R12103 VPWR.n2051 VPWR.n2050 3.4105
R12104 VPWR.n2099 VPWR.n659 3.4105
R12105 VPWR.n2148 VPWR.n2147 3.4105
R12106 VPWR.n2196 VPWR.n562 3.4105
R12107 VPWR.n2247 VPWR.n2246 3.4105
R12108 VPWR.n2295 VPWR.n467 3.4105
R12109 VPWR.n2344 VPWR.n2343 3.4105
R12110 VPWR.n2392 VPWR.n370 3.4105
R12111 VPWR.n2443 VPWR.n2442 3.4105
R12112 VPWR.n2451 VPWR.n2450 3.4105
R12113 VPWR.n2453 VPWR.n2452 3.4105
R12114 VPWR.n2461 VPWR.n2460 3.4105
R12115 VPWR.n2463 VPWR.n2462 3.4105
R12116 VPWR.n2471 VPWR.n2470 3.4105
R12117 VPWR.n2387 VPWR.n359 3.4105
R12118 VPWR.n2316 VPWR.n2315 3.4105
R12119 VPWR.n2300 VPWR.n478 3.4105
R12120 VPWR.n2275 VPWR.n2274 3.4105
R12121 VPWR.n2191 VPWR.n551 3.4105
R12122 VPWR.n2120 VPWR.n2119 3.4105
R12123 VPWR.n2104 VPWR.n670 3.4105
R12124 VPWR.n2079 VPWR.n2078 3.4105
R12125 VPWR.n1995 VPWR.n743 3.4105
R12126 VPWR.n1924 VPWR.n1923 3.4105
R12127 VPWR.n1908 VPWR.n862 3.4105
R12128 VPWR.n1883 VPWR.n1882 3.4105
R12129 VPWR.n1799 VPWR.n935 3.4105
R12130 VPWR.n1800 VPWR.n938 3.4105
R12131 VPWR.n1801 VPWR.n939 3.4105
R12132 VPWR.n1802 VPWR.n942 3.4105
R12133 VPWR.n1803 VPWR.n943 3.4105
R12134 VPWR.n1804 VPWR.n946 3.4105
R12135 VPWR.n1805 VPWR.n947 3.4105
R12136 VPWR.n1853 VPWR.n1852 3.4105
R12137 VPWR.n1902 VPWR.n850 3.4105
R12138 VPWR.n1954 VPWR.n1953 3.4105
R12139 VPWR.n2001 VPWR.n755 3.4105
R12140 VPWR.n2049 VPWR.n2048 3.4105
R12141 VPWR.n2098 VPWR.n658 3.4105
R12142 VPWR.n2150 VPWR.n2149 3.4105
R12143 VPWR.n2197 VPWR.n563 3.4105
R12144 VPWR.n2245 VPWR.n2244 3.4105
R12145 VPWR.n2294 VPWR.n466 3.4105
R12146 VPWR.n2346 VPWR.n2345 3.4105
R12147 VPWR.n2393 VPWR.n371 3.4105
R12148 VPWR.n2441 VPWR.n2440 3.4105
R12149 VPWR.n2433 VPWR.n2432 3.4105
R12150 VPWR.n2394 VPWR.n374 3.4105
R12151 VPWR.n2354 VPWR.n2353 3.4105
R12152 VPWR.n2293 VPWR.n463 3.4105
R12153 VPWR.n2237 VPWR.n2236 3.4105
R12154 VPWR.n2198 VPWR.n566 3.4105
R12155 VPWR.n2158 VPWR.n2157 3.4105
R12156 VPWR.n2097 VPWR.n655 3.4105
R12157 VPWR.n2041 VPWR.n2040 3.4105
R12158 VPWR.n2002 VPWR.n758 3.4105
R12159 VPWR.n1962 VPWR.n1961 3.4105
R12160 VPWR.n1901 VPWR.n847 3.4105
R12161 VPWR.n1845 VPWR.n1844 3.4105
R12162 VPWR.n1806 VPWR.n950 3.4105
R12163 VPWR.n1798 VPWR.n934 3.4105
R12164 VPWR.n1885 VPWR.n1884 3.4105
R12165 VPWR.n1909 VPWR.n863 3.4105
R12166 VPWR.n1922 VPWR.n1921 3.4105
R12167 VPWR.n1994 VPWR.n742 3.4105
R12168 VPWR.n2081 VPWR.n2080 3.4105
R12169 VPWR.n2105 VPWR.n671 3.4105
R12170 VPWR.n2118 VPWR.n2117 3.4105
R12171 VPWR.n2190 VPWR.n550 3.4105
R12172 VPWR.n2277 VPWR.n2276 3.4105
R12173 VPWR.n2301 VPWR.n479 3.4105
R12174 VPWR.n2314 VPWR.n2313 3.4105
R12175 VPWR.n2386 VPWR.n358 3.4105
R12176 VPWR.n2473 VPWR.n2472 3.4105
R12177 VPWR.n2497 VPWR.n96 3.4105
R12178 VPWR.n2496 VPWR.n95 3.4105
R12179 VPWR.n2495 VPWR.n90 3.4105
R12180 VPWR.n2494 VPWR.n89 3.4105
R12181 VPWR.n2493 VPWR.n84 3.4105
R12182 VPWR.n2492 VPWR.n83 3.4105
R12183 VPWR.n2491 VPWR.n78 3.4105
R12184 VPWR.n2490 VPWR.n77 3.4105
R12185 VPWR.n2489 VPWR.n72 3.4105
R12186 VPWR.n2488 VPWR.n71 3.4105
R12187 VPWR.n2431 VPWR.n2430 3.4105
R12188 VPWR.n2395 VPWR.n375 3.4105
R12189 VPWR.n2356 VPWR.n2355 3.4105
R12190 VPWR.n2292 VPWR.n462 3.4105
R12191 VPWR.n2235 VPWR.n2234 3.4105
R12192 VPWR.n2199 VPWR.n567 3.4105
R12193 VPWR.n2160 VPWR.n2159 3.4105
R12194 VPWR.n2096 VPWR.n654 3.4105
R12195 VPWR.n2039 VPWR.n2038 3.4105
R12196 VPWR.n2003 VPWR.n759 3.4105
R12197 VPWR.n1964 VPWR.n1963 3.4105
R12198 VPWR.n1900 VPWR.n846 3.4105
R12199 VPWR.n1843 VPWR.n1842 3.4105
R12200 VPWR.n1807 VPWR.n951 3.4105
R12201 VPWR.n1532 VPWR.n1143 3.4105
R12202 VPWR.n1540 VPWR.n1539 3.4105
R12203 VPWR.n1525 VPWR.n1524 3.4105
R12204 VPWR.n1517 VPWR.n1516 3.4105
R12205 VPWR.n1511 VPWR.n1510 3.4105
R12206 VPWR.n1503 VPWR.n1502 3.4105
R12207 VPWR.n1497 VPWR.n1496 3.4105
R12208 VPWR.n1489 VPWR.n1132 3.4105
R12209 VPWR.n1585 VPWR.n1584 3.4105
R12210 VPWR.n1452 VPWR.n1128 3.4105
R12211 VPWR.n1765 VPWR.n1764 3.4105
R12212 VPWR.n1808 VPWR.n954 3.4105
R12213 VPWR.n1835 VPWR.n1834 3.4105
R12214 VPWR.n1899 VPWR.n843 3.4105
R12215 VPWR.n1972 VPWR.n1971 3.4105
R12216 VPWR.n2004 VPWR.n762 3.4105
R12217 VPWR.n2031 VPWR.n2030 3.4105
R12218 VPWR.n2095 VPWR.n651 3.4105
R12219 VPWR.n2168 VPWR.n2167 3.4105
R12220 VPWR.n2200 VPWR.n570 3.4105
R12221 VPWR.n2227 VPWR.n2226 3.4105
R12222 VPWR.n2291 VPWR.n459 3.4105
R12223 VPWR.n2364 VPWR.n2363 3.4105
R12224 VPWR.n2396 VPWR.n378 3.4105
R12225 VPWR.n2423 VPWR.n2422 3.4105
R12226 VPWR.n2487 VPWR.n66 3.4105
R12227 VPWR.n2485 VPWR.n60 3.4105
R12228 VPWR.n2413 VPWR.n2412 3.4105
R12229 VPWR.n2398 VPWR.n382 3.4105
R12230 VPWR.n2374 VPWR.n2373 3.4105
R12231 VPWR.n2289 VPWR.n455 3.4105
R12232 VPWR.n2217 VPWR.n2216 3.4105
R12233 VPWR.n2202 VPWR.n574 3.4105
R12234 VPWR.n2178 VPWR.n2177 3.4105
R12235 VPWR.n2093 VPWR.n647 3.4105
R12236 VPWR.n2021 VPWR.n2020 3.4105
R12237 VPWR.n2006 VPWR.n766 3.4105
R12238 VPWR.n1982 VPWR.n1981 3.4105
R12239 VPWR.n1897 VPWR.n839 3.4105
R12240 VPWR.n1825 VPWR.n1824 3.4105
R12241 VPWR.n1810 VPWR.n958 3.4105
R12242 VPWR.n1752 VPWR.n1744 3.4105
R12243 VPWR.n1757 VPWR.n1043 3.4105
R12244 VPWR.n1809 VPWR.n955 3.4105
R12245 VPWR.n1833 VPWR.n1832 3.4105
R12246 VPWR.n1898 VPWR.n842 3.4105
R12247 VPWR.n1974 VPWR.n1973 3.4105
R12248 VPWR.n2005 VPWR.n763 3.4105
R12249 VPWR.n2029 VPWR.n2028 3.4105
R12250 VPWR.n2094 VPWR.n650 3.4105
R12251 VPWR.n2170 VPWR.n2169 3.4105
R12252 VPWR.n2201 VPWR.n571 3.4105
R12253 VPWR.n2225 VPWR.n2224 3.4105
R12254 VPWR.n2290 VPWR.n458 3.4105
R12255 VPWR.n2366 VPWR.n2365 3.4105
R12256 VPWR.n2397 VPWR.n379 3.4105
R12257 VPWR.n2421 VPWR.n2420 3.4105
R12258 VPWR.n2486 VPWR.n65 3.4105
R12259 VPWR.n2484 VPWR.n59 3.4105
R12260 VPWR.n2411 VPWR.n2410 3.4105
R12261 VPWR.n2399 VPWR.n383 3.4105
R12262 VPWR.n2376 VPWR.n2375 3.4105
R12263 VPWR.n2288 VPWR.n454 3.4105
R12264 VPWR.n2215 VPWR.n2214 3.4105
R12265 VPWR.n2203 VPWR.n575 3.4105
R12266 VPWR.n2180 VPWR.n2179 3.4105
R12267 VPWR.n2092 VPWR.n646 3.4105
R12268 VPWR.n2019 VPWR.n2018 3.4105
R12269 VPWR.n2007 VPWR.n767 3.4105
R12270 VPWR.n1984 VPWR.n1983 3.4105
R12271 VPWR.n1896 VPWR.n838 3.4105
R12272 VPWR.n1823 VPWR.n1822 3.4105
R12273 VPWR.n1811 VPWR.n959 3.4105
R12274 VPWR.n1788 VPWR.n1787 3.4105
R12275 VPWR.n1465 VPWR.n1464 3.4105
R12276 VPWR.n1797 VPWR.n931 3.4105
R12277 VPWR.n1893 VPWR.n1892 3.4105
R12278 VPWR.n1910 VPWR.n929 3.4105
R12279 VPWR.n1914 VPWR.n1913 3.4105
R12280 VPWR.n1993 VPWR.n739 3.4105
R12281 VPWR.n2089 VPWR.n2088 3.4105
R12282 VPWR.n2106 VPWR.n737 3.4105
R12283 VPWR.n2110 VPWR.n2109 3.4105
R12284 VPWR.n2189 VPWR.n547 3.4105
R12285 VPWR.n2285 VPWR.n2284 3.4105
R12286 VPWR.n2302 VPWR.n545 3.4105
R12287 VPWR.n2306 VPWR.n2305 3.4105
R12288 VPWR.n2385 VPWR.n355 3.4105
R12289 VPWR.n2481 VPWR.n2480 3.4105
R12290 VPWR.n2498 VPWR.n353 3.4105
R12291 VPWR.n2502 VPWR.n2501 3.4105
R12292 VPWR.n2512 VPWR.n2511 3.4105
R12293 VPWR.n2514 VPWR.n2513 3.4105
R12294 VPWR.n2524 VPWR.n2523 3.4105
R12295 VPWR.n2526 VPWR.n2525 3.4105
R12296 VPWR.n2536 VPWR.n2535 3.4105
R12297 VPWR.n2538 VPWR.n2537 3.4105
R12298 VPWR.n2548 VPWR.n2547 3.4105
R12299 VPWR.n2550 VPWR.n2549 3.4105
R12300 VPWR.n2560 VPWR.n2559 3.4105
R12301 VPWR.n2562 VPWR.n2561 3.4105
R12302 VPWR.n2572 VPWR.n2571 3.4105
R12303 VPWR.n2574 VPWR.n2573 3.4105
R12304 VPWR.n2584 VPWR.n2583 3.4105
R12305 VPWR.n2586 VPWR.n2585 3.4105
R12306 VPWR.n2595 VPWR.n2594 3.4105
R12307 VPWR.n2483 VPWR.n22 3.4105
R12308 VPWR.n2404 VPWR.n2403 3.4105
R12309 VPWR.n2400 VPWR.n449 3.4105
R12310 VPWR.n2383 VPWR.n2382 3.4105
R12311 VPWR.n2287 VPWR.n451 3.4105
R12312 VPWR.n2208 VPWR.n2207 3.4105
R12313 VPWR.n2204 VPWR.n641 3.4105
R12314 VPWR.n2187 VPWR.n2186 3.4105
R12315 VPWR.n2091 VPWR.n643 3.4105
R12316 VPWR.n2012 VPWR.n2011 3.4105
R12317 VPWR.n2008 VPWR.n833 3.4105
R12318 VPWR.n1991 VPWR.n1990 3.4105
R12319 VPWR.n1895 VPWR.n835 3.4105
R12320 VPWR.n1816 VPWR.n1815 3.4105
R12321 VPWR.n1812 VPWR.n1025 3.4105
R12322 VPWR.n1795 VPWR.n1794 3.4105
R12323 VPWR.n1055 VPWR.n1028 3.4105
R12324 VPWR.n1056 VPWR.n1037 3.4105
R12325 VPWR.n1754 VPWR.n1753 3.4105
R12326 VPWR.n1756 VPWR.n1755 3.4105
R12327 VPWR.n1529 VPWR.n1045 3.4105
R12328 VPWR.n1531 VPWR.n1530 3.4105
R12329 VPWR.n1528 VPWR.n1145 3.4105
R12330 VPWR.n1527 VPWR.n1526 3.4105
R12331 VPWR.n1515 VPWR.n1514 3.4105
R12332 VPWR.n1513 VPWR.n1512 3.4105
R12333 VPWR.n1501 VPWR.n1500 3.4105
R12334 VPWR.n1499 VPWR.n1498 3.4105
R12335 VPWR.n1488 VPWR.n1487 3.4105
R12336 VPWR.n1587 VPWR.n1586 3.4105
R12337 VPWR.n1589 VPWR.n1588 3.4105
R12338 VPWR.n1448 VPWR.n1232 3.4105
R12339 VPWR.n1345 VPWR.n1341 3.38874
R12340 VPWR.n1384 VPWR.n1380 3.38874
R12341 VPWR.n1421 VPWR.n1417 3.38874
R12342 VPWR.n28 VPWR.n26 3.36211
R12343 VPWR.n30 VPWR.n28 3.36211
R12344 VPWR.n32 VPWR.n30 3.36211
R12345 VPWR.n34 VPWR.n32 3.36211
R12346 VPWR.n36 VPWR.n34 3.36211
R12347 VPWR.n38 VPWR.n36 3.36211
R12348 VPWR.n40 VPWR.n38 3.36211
R12349 VPWR.n42 VPWR.n40 3.36211
R12350 VPWR.n44 VPWR.n42 3.36211
R12351 VPWR.n46 VPWR.n44 3.36211
R12352 VPWR.n48 VPWR.n46 3.36211
R12353 VPWR.n50 VPWR.n48 3.36211
R12354 VPWR.n52 VPWR.n50 3.36211
R12355 VPWR.n54 VPWR.n52 3.36211
R12356 VPWR.t1198 VPWR.t1232 3.35739
R12357 VPWR.t189 VPWR.t1235 3.35739
R12358 VPWR.n2571 VPWR.n66 3.28012
R12359 VPWR.n2511 VPWR.n96 3.28012
R12360 VPWR.n2550 VPWR.n77 3.28012
R12361 VPWR.n2440 VPWR.n77 3.28012
R12362 VPWR.n2547 VPWR.n78 3.28012
R12363 VPWR.n2443 VPWR.n78 3.28012
R12364 VPWR.n2535 VPWR.n84 3.28012
R12365 VPWR.n2453 VPWR.n84 3.28012
R12366 VPWR.n2453 VPWR.n366 3.28012
R12367 VPWR.n2526 VPWR.n89 3.28012
R12368 VPWR.n2460 VPWR.n89 3.28012
R12369 VPWR.n2460 VPWR.n363 3.28012
R12370 VPWR.n1498 VPWR.n1497 3.28012
R12371 VPWR.n1497 VPWR.n939 3.28012
R12372 VPWR.n1872 VPWR.n939 3.28012
R12373 VPWR.n1872 VPWR.n858 3.28012
R12374 VPWR.n1934 VPWR.n858 3.28012
R12375 VPWR.n1934 VPWR.n747 3.28012
R12376 VPWR.n2068 VPWR.n747 3.28012
R12377 VPWR.n2068 VPWR.n666 3.28012
R12378 VPWR.n2130 VPWR.n666 3.28012
R12379 VPWR.n2130 VPWR.n555 3.28012
R12380 VPWR.n2264 VPWR.n555 3.28012
R12381 VPWR.n2264 VPWR.n474 3.28012
R12382 VPWR.n2326 VPWR.n474 3.28012
R12383 VPWR.n2326 VPWR.n363 3.28012
R12384 VPWR.n2523 VPWR.n90 3.28012
R12385 VPWR.n2463 VPWR.n90 3.28012
R12386 VPWR.n2463 VPWR.n362 3.28012
R12387 VPWR.n2323 VPWR.n362 3.28012
R12388 VPWR.n2323 VPWR.n475 3.28012
R12389 VPWR.n2267 VPWR.n475 3.28012
R12390 VPWR.n2267 VPWR.n554 3.28012
R12391 VPWR.n2127 VPWR.n554 3.28012
R12392 VPWR.n2127 VPWR.n667 3.28012
R12393 VPWR.n2071 VPWR.n667 3.28012
R12394 VPWR.n2071 VPWR.n746 3.28012
R12395 VPWR.n1931 VPWR.n746 3.28012
R12396 VPWR.n1931 VPWR.n859 3.28012
R12397 VPWR.n1875 VPWR.n859 3.28012
R12398 VPWR.n1489 VPWR.n1488 3.28012
R12399 VPWR.n1489 VPWR.n938 3.28012
R12400 VPWR.n1875 VPWR.n938 3.28012
R12401 VPWR.n1503 VPWR.n1501 3.28012
R12402 VPWR.n1503 VPWR.n942 3.28012
R12403 VPWR.n1865 VPWR.n942 3.28012
R12404 VPWR.n1865 VPWR.n855 3.28012
R12405 VPWR.n1941 VPWR.n855 3.28012
R12406 VPWR.n1941 VPWR.n750 3.28012
R12407 VPWR.n2061 VPWR.n750 3.28012
R12408 VPWR.n2061 VPWR.n663 3.28012
R12409 VPWR.n2137 VPWR.n663 3.28012
R12410 VPWR.n2137 VPWR.n558 3.28012
R12411 VPWR.n2257 VPWR.n558 3.28012
R12412 VPWR.n2257 VPWR.n471 3.28012
R12413 VPWR.n2333 VPWR.n471 3.28012
R12414 VPWR.n2333 VPWR.n366 3.28012
R12415 VPWR.n2538 VPWR.n83 3.28012
R12416 VPWR.n2450 VPWR.n83 3.28012
R12417 VPWR.n2450 VPWR.n367 3.28012
R12418 VPWR.n2336 VPWR.n367 3.28012
R12419 VPWR.n2336 VPWR.n470 3.28012
R12420 VPWR.n2254 VPWR.n470 3.28012
R12421 VPWR.n2254 VPWR.n559 3.28012
R12422 VPWR.n2140 VPWR.n559 3.28012
R12423 VPWR.n2140 VPWR.n662 3.28012
R12424 VPWR.n2058 VPWR.n662 3.28012
R12425 VPWR.n2058 VPWR.n751 3.28012
R12426 VPWR.n1944 VPWR.n751 3.28012
R12427 VPWR.n1944 VPWR.n854 3.28012
R12428 VPWR.n1862 VPWR.n854 3.28012
R12429 VPWR.n1512 VPWR.n1511 3.28012
R12430 VPWR.n1511 VPWR.n943 3.28012
R12431 VPWR.n1862 VPWR.n943 3.28012
R12432 VPWR.n1517 VPWR.n1515 3.28012
R12433 VPWR.n1517 VPWR.n946 3.28012
R12434 VPWR.n1855 VPWR.n946 3.28012
R12435 VPWR.n1855 VPWR.n851 3.28012
R12436 VPWR.n1951 VPWR.n851 3.28012
R12437 VPWR.n1951 VPWR.n754 3.28012
R12438 VPWR.n2051 VPWR.n754 3.28012
R12439 VPWR.n2051 VPWR.n659 3.28012
R12440 VPWR.n2147 VPWR.n659 3.28012
R12441 VPWR.n2147 VPWR.n562 3.28012
R12442 VPWR.n2247 VPWR.n562 3.28012
R12443 VPWR.n2247 VPWR.n467 3.28012
R12444 VPWR.n2343 VPWR.n467 3.28012
R12445 VPWR.n2343 VPWR.n370 3.28012
R12446 VPWR.n2443 VPWR.n370 3.28012
R12447 VPWR.n2514 VPWR.n95 3.28012
R12448 VPWR.n2470 VPWR.n95 3.28012
R12449 VPWR.n2470 VPWR.n359 3.28012
R12450 VPWR.n2316 VPWR.n359 3.28012
R12451 VPWR.n2316 VPWR.n478 3.28012
R12452 VPWR.n2274 VPWR.n478 3.28012
R12453 VPWR.n2274 VPWR.n551 3.28012
R12454 VPWR.n2120 VPWR.n551 3.28012
R12455 VPWR.n2120 VPWR.n670 3.28012
R12456 VPWR.n2078 VPWR.n670 3.28012
R12457 VPWR.n2078 VPWR.n743 3.28012
R12458 VPWR.n1924 VPWR.n743 3.28012
R12459 VPWR.n1924 VPWR.n862 3.28012
R12460 VPWR.n1882 VPWR.n862 3.28012
R12461 VPWR.n1882 VPWR.n935 3.28012
R12462 VPWR.n1586 VPWR.n1585 3.28012
R12463 VPWR.n1585 VPWR.n935 3.28012
R12464 VPWR.n1526 VPWR.n1525 3.28012
R12465 VPWR.n1525 VPWR.n947 3.28012
R12466 VPWR.n1852 VPWR.n947 3.28012
R12467 VPWR.n1852 VPWR.n850 3.28012
R12468 VPWR.n1954 VPWR.n850 3.28012
R12469 VPWR.n1954 VPWR.n755 3.28012
R12470 VPWR.n2048 VPWR.n755 3.28012
R12471 VPWR.n2048 VPWR.n658 3.28012
R12472 VPWR.n2150 VPWR.n658 3.28012
R12473 VPWR.n2150 VPWR.n563 3.28012
R12474 VPWR.n2244 VPWR.n563 3.28012
R12475 VPWR.n2244 VPWR.n466 3.28012
R12476 VPWR.n2346 VPWR.n466 3.28012
R12477 VPWR.n2346 VPWR.n371 3.28012
R12478 VPWR.n2440 VPWR.n371 3.28012
R12479 VPWR.n2559 VPWR.n72 3.28012
R12480 VPWR.n2433 VPWR.n72 3.28012
R12481 VPWR.n2433 VPWR.n374 3.28012
R12482 VPWR.n2353 VPWR.n374 3.28012
R12483 VPWR.n2353 VPWR.n463 3.28012
R12484 VPWR.n2237 VPWR.n463 3.28012
R12485 VPWR.n2237 VPWR.n566 3.28012
R12486 VPWR.n2157 VPWR.n566 3.28012
R12487 VPWR.n2157 VPWR.n655 3.28012
R12488 VPWR.n2041 VPWR.n655 3.28012
R12489 VPWR.n2041 VPWR.n758 3.28012
R12490 VPWR.n1961 VPWR.n758 3.28012
R12491 VPWR.n1961 VPWR.n847 3.28012
R12492 VPWR.n1845 VPWR.n847 3.28012
R12493 VPWR.n1845 VPWR.n950 3.28012
R12494 VPWR.n1539 VPWR.n1145 3.28012
R12495 VPWR.n1539 VPWR.n950 3.28012
R12496 VPWR.n1589 VPWR.n1128 3.28012
R12497 VPWR.n1128 VPWR.n934 3.28012
R12498 VPWR.n1885 VPWR.n934 3.28012
R12499 VPWR.n1885 VPWR.n863 3.28012
R12500 VPWR.n1921 VPWR.n863 3.28012
R12501 VPWR.n1921 VPWR.n742 3.28012
R12502 VPWR.n2081 VPWR.n742 3.28012
R12503 VPWR.n2081 VPWR.n671 3.28012
R12504 VPWR.n2117 VPWR.n671 3.28012
R12505 VPWR.n2117 VPWR.n550 3.28012
R12506 VPWR.n2277 VPWR.n550 3.28012
R12507 VPWR.n2277 VPWR.n479 3.28012
R12508 VPWR.n2313 VPWR.n479 3.28012
R12509 VPWR.n2313 VPWR.n358 3.28012
R12510 VPWR.n2473 VPWR.n358 3.28012
R12511 VPWR.n2473 VPWR.n96 3.28012
R12512 VPWR.n2562 VPWR.n71 3.28012
R12513 VPWR.n2430 VPWR.n71 3.28012
R12514 VPWR.n2430 VPWR.n375 3.28012
R12515 VPWR.n2356 VPWR.n375 3.28012
R12516 VPWR.n2356 VPWR.n462 3.28012
R12517 VPWR.n2234 VPWR.n462 3.28012
R12518 VPWR.n2234 VPWR.n567 3.28012
R12519 VPWR.n2160 VPWR.n567 3.28012
R12520 VPWR.n2160 VPWR.n654 3.28012
R12521 VPWR.n2038 VPWR.n654 3.28012
R12522 VPWR.n2038 VPWR.n759 3.28012
R12523 VPWR.n1964 VPWR.n759 3.28012
R12524 VPWR.n1964 VPWR.n846 3.28012
R12525 VPWR.n1842 VPWR.n846 3.28012
R12526 VPWR.n1842 VPWR.n951 3.28012
R12527 VPWR.n1532 VPWR.n951 3.28012
R12528 VPWR.n1532 VPWR.n1531 3.28012
R12529 VPWR.n1764 VPWR.n1045 3.28012
R12530 VPWR.n1764 VPWR.n954 3.28012
R12531 VPWR.n1835 VPWR.n954 3.28012
R12532 VPWR.n1835 VPWR.n843 3.28012
R12533 VPWR.n1971 VPWR.n843 3.28012
R12534 VPWR.n1971 VPWR.n762 3.28012
R12535 VPWR.n2031 VPWR.n762 3.28012
R12536 VPWR.n2031 VPWR.n651 3.28012
R12537 VPWR.n2167 VPWR.n651 3.28012
R12538 VPWR.n2167 VPWR.n570 3.28012
R12539 VPWR.n2227 VPWR.n570 3.28012
R12540 VPWR.n2227 VPWR.n459 3.28012
R12541 VPWR.n2363 VPWR.n459 3.28012
R12542 VPWR.n2363 VPWR.n378 3.28012
R12543 VPWR.n2423 VPWR.n378 3.28012
R12544 VPWR.n2423 VPWR.n66 3.28012
R12545 VPWR.n2583 VPWR.n60 3.28012
R12546 VPWR.n2413 VPWR.n60 3.28012
R12547 VPWR.n2413 VPWR.n382 3.28012
R12548 VPWR.n2373 VPWR.n382 3.28012
R12549 VPWR.n2373 VPWR.n455 3.28012
R12550 VPWR.n2217 VPWR.n455 3.28012
R12551 VPWR.n2217 VPWR.n574 3.28012
R12552 VPWR.n2177 VPWR.n574 3.28012
R12553 VPWR.n2177 VPWR.n647 3.28012
R12554 VPWR.n2021 VPWR.n647 3.28012
R12555 VPWR.n2021 VPWR.n766 3.28012
R12556 VPWR.n1981 VPWR.n766 3.28012
R12557 VPWR.n1981 VPWR.n839 3.28012
R12558 VPWR.n1825 VPWR.n839 3.28012
R12559 VPWR.n1825 VPWR.n958 3.28012
R12560 VPWR.n1752 VPWR.n958 3.28012
R12561 VPWR.n1753 VPWR.n1752 3.28012
R12562 VPWR.n1757 VPWR.n1756 3.28012
R12563 VPWR.n1757 VPWR.n955 3.28012
R12564 VPWR.n1832 VPWR.n955 3.28012
R12565 VPWR.n1832 VPWR.n842 3.28012
R12566 VPWR.n1974 VPWR.n842 3.28012
R12567 VPWR.n1974 VPWR.n763 3.28012
R12568 VPWR.n2028 VPWR.n763 3.28012
R12569 VPWR.n2028 VPWR.n650 3.28012
R12570 VPWR.n2170 VPWR.n650 3.28012
R12571 VPWR.n2170 VPWR.n571 3.28012
R12572 VPWR.n2224 VPWR.n571 3.28012
R12573 VPWR.n2224 VPWR.n458 3.28012
R12574 VPWR.n2366 VPWR.n458 3.28012
R12575 VPWR.n2366 VPWR.n379 3.28012
R12576 VPWR.n2420 VPWR.n379 3.28012
R12577 VPWR.n2420 VPWR.n65 3.28012
R12578 VPWR.n2574 VPWR.n65 3.28012
R12579 VPWR.n2586 VPWR.n59 3.28012
R12580 VPWR.n2410 VPWR.n59 3.28012
R12581 VPWR.n2410 VPWR.n383 3.28012
R12582 VPWR.n2376 VPWR.n383 3.28012
R12583 VPWR.n2376 VPWR.n454 3.28012
R12584 VPWR.n2214 VPWR.n454 3.28012
R12585 VPWR.n2214 VPWR.n575 3.28012
R12586 VPWR.n2180 VPWR.n575 3.28012
R12587 VPWR.n2180 VPWR.n646 3.28012
R12588 VPWR.n2018 VPWR.n646 3.28012
R12589 VPWR.n2018 VPWR.n767 3.28012
R12590 VPWR.n1984 VPWR.n767 3.28012
R12591 VPWR.n1984 VPWR.n838 3.28012
R12592 VPWR.n1822 VPWR.n838 3.28012
R12593 VPWR.n1822 VPWR.n959 3.28012
R12594 VPWR.n1788 VPWR.n959 3.28012
R12595 VPWR.n1788 VPWR.n1037 3.28012
R12596 VPWR.n1465 VPWR.n1232 3.28012
R12597 VPWR.n1465 VPWR.n931 3.28012
R12598 VPWR.n1892 VPWR.n931 3.28012
R12599 VPWR.n1892 VPWR.n929 3.28012
R12600 VPWR.n1914 VPWR.n929 3.28012
R12601 VPWR.n1914 VPWR.n739 3.28012
R12602 VPWR.n2088 VPWR.n739 3.28012
R12603 VPWR.n2088 VPWR.n737 3.28012
R12604 VPWR.n2110 VPWR.n737 3.28012
R12605 VPWR.n2110 VPWR.n547 3.28012
R12606 VPWR.n2284 VPWR.n547 3.28012
R12607 VPWR.n2284 VPWR.n545 3.28012
R12608 VPWR.n2306 VPWR.n545 3.28012
R12609 VPWR.n2306 VPWR.n355 3.28012
R12610 VPWR.n2480 VPWR.n355 3.28012
R12611 VPWR.n2480 VPWR.n353 3.28012
R12612 VPWR.n2502 VPWR.n353 3.28012
R12613 VPWR.n2404 VPWR.n22 3.28012
R12614 VPWR.n2404 VPWR.n449 3.28012
R12615 VPWR.n2382 VPWR.n449 3.28012
R12616 VPWR.n2382 VPWR.n451 3.28012
R12617 VPWR.n2208 VPWR.n451 3.28012
R12618 VPWR.n2208 VPWR.n641 3.28012
R12619 VPWR.n2186 VPWR.n641 3.28012
R12620 VPWR.n2186 VPWR.n643 3.28012
R12621 VPWR.n2012 VPWR.n643 3.28012
R12622 VPWR.n2012 VPWR.n833 3.28012
R12623 VPWR.n1990 VPWR.n833 3.28012
R12624 VPWR.n1990 VPWR.n835 3.28012
R12625 VPWR.n1816 VPWR.n835 3.28012
R12626 VPWR.n1816 VPWR.n1025 3.28012
R12627 VPWR.n1794 VPWR.n1025 3.28012
R12628 VPWR.n1794 VPWR.n1028 3.28012
R12629 VPWR.n2594 VPWR.n22 3.26393
R12630 VPWR.n2863 VPWR 3.18182
R12631 VPWR.n2832 VPWR.n2831 3.1005
R12632 VPWR.n2826 VPWR.n2825 3.1005
R12633 VPWR.n2846 VPWR.n2815 3.1005
R12634 VPWR.n1324 VPWR.n1322 3.01226
R12635 VPWR.n1328 VPWR.n1304 2.63579
R12636 VPWR.n2731 VPWR.n2730 2.25932
R12637 VPWR.n1447 VPWR.n1446 2.06026
R12638 VPWR.n1447 VPWR.n1026 1.78803
R12639 VPWR.n2384 VPWR.n2383 1.32852
R12640 VPWR.n2287 VPWR.n450 1.32852
R12641 VPWR.n2207 VPWR.n2206 1.32852
R12642 VPWR.n2205 VPWR.n2204 1.32852
R12643 VPWR.n2188 VPWR.n2187 1.32852
R12644 VPWR.n2091 VPWR.n642 1.32852
R12645 VPWR.n2011 VPWR.n2010 1.32852
R12646 VPWR.n2009 VPWR.n2008 1.32852
R12647 VPWR.n1992 VPWR.n1991 1.32852
R12648 VPWR.n1895 VPWR.n834 1.32852
R12649 VPWR.n2401 VPWR.n2400 1.32852
R12650 VPWR.n1815 VPWR.n1814 1.32852
R12651 VPWR.n2403 VPWR.n2402 1.32852
R12652 VPWR.n1813 VPWR.n1812 1.32852
R12653 VPWR.n2483 VPWR.n21 1.32852
R12654 VPWR.n1796 VPWR.n1795 1.32852
R12655 VPWR.n2596 VPWR.n2595 1.32852
R12656 VPWR.n1055 VPWR.n1026 1.32852
R12657 VPWR.n2482 VPWR 1.25994
R12658 VPWR VPWR.n354 1.25994
R12659 VPWR VPWR.n2304 1.25994
R12660 VPWR.n2303 VPWR 1.25994
R12661 VPWR.n2286 VPWR 1.25994
R12662 VPWR VPWR.n546 1.25994
R12663 VPWR VPWR.n2108 1.25994
R12664 VPWR.n2107 VPWR 1.25994
R12665 VPWR.n2090 VPWR 1.25994
R12666 VPWR VPWR.n738 1.25994
R12667 VPWR VPWR.n1912 1.25994
R12668 VPWR.n1911 VPWR 1.25994
R12669 VPWR.n1894 VPWR 1.25994
R12670 VPWR VPWR.n930 1.25994
R12671 VPWR.n2499 VPWR 1.25994
R12672 VPWR VPWR.n1450 1.25994
R12673 VPWR VPWR.n2500 1.25994
R12674 VPWR.n1449 VPWR 1.25994
R12675 VPWR.n2597 VPWR.n2596 1.144
R12676 VPWR.n2861 VPWR.n2860 0.936724
R12677 VPWR.n2592 VPWR 0.925943
R12678 VPWR VPWR.n1063 0.925943
R12679 VPWR.n2860 VPWR.n2816 0.925245
R12680 VPWR.n2569 VPWR.n67 0.904391
R12681 VPWR.n2509 VPWR.n97 0.904391
R12682 VPWR.n2552 VPWR.n76 0.904391
R12683 VPWR.n2545 VPWR.n79 0.904391
R12684 VPWR.n2533 VPWR.n85 0.904391
R12685 VPWR.n2528 VPWR.n88 0.904391
R12686 VPWR.n1222 VPWR.n1178 0.904391
R12687 VPWR.n2521 VPWR.n91 0.904391
R12688 VPWR.n1624 VPWR.n1102 0.904391
R12689 VPWR.n1640 VPWR.n1094 0.904391
R12690 VPWR.n2540 VPWR.n82 0.904391
R12691 VPWR.n1651 VPWR.n1092 0.904391
R12692 VPWR.n1211 VPWR.n1210 0.904391
R12693 VPWR.n2516 VPWR.n94 0.904391
R12694 VPWR.n1613 VPWR.n1104 0.904391
R12695 VPWR.n1667 VPWR.n1084 0.904391
R12696 VPWR.n2557 VPWR.n73 0.904391
R12697 VPWR.n1678 VPWR.n1082 0.904391
R12698 VPWR.n1591 VPWR.n1127 0.904391
R12699 VPWR.n2564 VPWR.n70 0.904391
R12700 VPWR.n1197 VPWR.n1196 0.904391
R12701 VPWR.n1694 VPWR.n1074 0.904391
R12702 VPWR.n1742 VPWR.n1057 0.904391
R12703 VPWR.n1705 VPWR.n1071 0.904391
R12704 VPWR.n2581 VPWR.n61 0.904391
R12705 VPWR.n2588 VPWR.n58 0.904391
R12706 VPWR.n1737 VPWR.n1735 0.904391
R12707 VPWR.n1597 VPWR.n1596 0.904391
R12708 VPWR.n2504 VPWR.n289 0.904391
R12709 VPWR.n2576 VPWR.n64 0.904391
R12710 VPWR VPWR.n2863 0.812229
R12711 VPWR.n140 VPWR.n64 0.675548
R12712 VPWR.n152 VPWR.n67 0.675548
R12713 VPWR.n164 VPWR.n70 0.675548
R12714 VPWR.n176 VPWR.n73 0.675548
R12715 VPWR.n188 VPWR.n76 0.675548
R12716 VPWR.n200 VPWR.n79 0.675548
R12717 VPWR.n212 VPWR.n82 0.675548
R12718 VPWR.n224 VPWR.n85 0.675548
R12719 VPWR.n236 VPWR.n88 0.675548
R12720 VPWR.n248 VPWR.n91 0.675548
R12721 VPWR.n260 VPWR.n94 0.675548
R12722 VPWR.n272 VPWR.n97 0.675548
R12723 VPWR.n289 VPWR.n288 0.675548
R12724 VPWR.n128 VPWR.n61 0.675548
R12725 VPWR.n117 VPWR.n58 0.675548
R12726 VPWR.n1735 VPWR.n1734 0.675548
R12727 VPWR.n1719 VPWR.n1057 0.675548
R12728 VPWR.n1707 VPWR.n1705 0.675548
R12729 VPWR.n1696 VPWR.n1694 0.675548
R12730 VPWR.n1196 VPWR.n1195 0.675548
R12731 VPWR.n1680 VPWR.n1678 0.675548
R12732 VPWR.n1669 VPWR.n1667 0.675548
R12733 VPWR.n1210 VPWR.n1209 0.675548
R12734 VPWR.n1653 VPWR.n1651 0.675548
R12735 VPWR.n1642 VPWR.n1640 0.675548
R12736 VPWR.n1178 VPWR.n1177 0.675548
R12737 VPWR.n1626 VPWR.n1624 0.675548
R12738 VPWR.n1615 VPWR.n1613 0.675548
R12739 VPWR.n1127 VPWR.n1126 0.675548
R12740 VPWR.n1599 VPWR.n1597 0.675548
R12741 VPWR.n2806 VPWR.n2805 0.672385
R12742 VPWR.n2790 VPWR.n2785 0.672385
R12743 VPWR.n2770 VPWR.n2765 0.672385
R12744 VPWR.n2751 VPWR.n2746 0.672385
R12745 VPWR.n7 VPWR 0.63497
R12746 VPWR.n1242 VPWR 0.63497
R12747 VPWR.n1265 VPWR 0.63497
R12748 VPWR.n1289 VPWR 0.63497
R12749 VPWR.n24 VPWR 0.499542
R12750 VPWR.n2814 VPWR.n2813 0.442692
R12751 VPWR.n1120 VPWR.n1118 0.404056
R12752 VPWR.n144 VPWR.n138 0.404056
R12753 VPWR.n156 VPWR.n150 0.404056
R12754 VPWR.n168 VPWR.n162 0.404056
R12755 VPWR.n180 VPWR.n174 0.404056
R12756 VPWR.n192 VPWR.n186 0.404056
R12757 VPWR.n204 VPWR.n198 0.404056
R12758 VPWR.n216 VPWR.n210 0.404056
R12759 VPWR.n228 VPWR.n222 0.404056
R12760 VPWR.n240 VPWR.n234 0.404056
R12761 VPWR.n252 VPWR.n246 0.404056
R12762 VPWR.n264 VPWR.n258 0.404056
R12763 VPWR.n276 VPWR.n270 0.404056
R12764 VPWR.n283 VPWR.n101 0.404056
R12765 VPWR.n110 VPWR.n105 0.404056
R12766 VPWR.n132 VPWR.n126 0.404056
R12767 VPWR.n121 VPWR.n115 0.404056
R12768 VPWR.n1729 VPWR.n1065 0.404056
R12769 VPWR.n1723 VPWR.n1717 0.404056
R12770 VPWR.n1711 VPWR.n1070 0.404056
R12771 VPWR.n1704 VPWR.n1702 0.404056
R12772 VPWR.n1693 VPWR.n1691 0.404056
R12773 VPWR.n1684 VPWR.n1081 0.404056
R12774 VPWR.n1677 VPWR.n1675 0.404056
R12775 VPWR.n1666 VPWR.n1664 0.404056
R12776 VPWR.n1657 VPWR.n1091 0.404056
R12777 VPWR.n1650 VPWR.n1648 0.404056
R12778 VPWR.n1639 VPWR.n1637 0.404056
R12779 VPWR.n1630 VPWR.n1101 0.404056
R12780 VPWR.n1623 VPWR.n1621 0.404056
R12781 VPWR.n1612 VPWR.n1610 0.404056
R12782 VPWR.n1603 VPWR.n1111 0.404056
R12783 VPWR.n2860 VPWR.n2859 0.388
R12784 VPWR.n1608 VPWR.n1607 0.349144
R12785 VPWR.n1608 VPWR.n1099 0.349144
R12786 VPWR.n1634 VPWR.n1099 0.349144
R12787 VPWR.n1635 VPWR.n1634 0.349144
R12788 VPWR.n1635 VPWR.n1089 0.349144
R12789 VPWR.n1661 VPWR.n1089 0.349144
R12790 VPWR.n1662 VPWR.n1661 0.349144
R12791 VPWR.n1662 VPWR.n1079 0.349144
R12792 VPWR.n1688 VPWR.n1079 0.349144
R12793 VPWR.n1689 VPWR.n1688 0.349144
R12794 VPWR.n1689 VPWR.n1068 0.349144
R12795 VPWR.n1715 VPWR.n1068 0.349144
R12796 VPWR.n1727 VPWR.n1715 0.349144
R12797 VPWR.n281 VPWR.n280 0.349144
R12798 VPWR.n280 VPWR.n268 0.349144
R12799 VPWR.n268 VPWR.n256 0.349144
R12800 VPWR.n256 VPWR.n244 0.349144
R12801 VPWR.n244 VPWR.n232 0.349144
R12802 VPWR.n232 VPWR.n220 0.349144
R12803 VPWR.n220 VPWR.n208 0.349144
R12804 VPWR.n208 VPWR.n196 0.349144
R12805 VPWR.n196 VPWR.n184 0.349144
R12806 VPWR.n184 VPWR.n172 0.349144
R12807 VPWR.n172 VPWR.n160 0.349144
R12808 VPWR.n160 VPWR.n148 0.349144
R12809 VPWR.n148 VPWR.n136 0.349144
R12810 VPWR.n1462 VPWR.n1456 0.346131
R12811 VPWR.n1461 VPWR.n1457 0.346131
R12812 VPWR.n1582 VPWR.n1136 0.346131
R12813 VPWR.n1581 VPWR.n1577 0.346131
R12814 VPWR.n1576 VPWR.n1572 0.346131
R12815 VPWR.n1571 VPWR.n1567 0.346131
R12816 VPWR.n1566 VPWR.n1562 0.346131
R12817 VPWR.n1561 VPWR.n1557 0.346131
R12818 VPWR.n1556 VPWR.n1552 0.346131
R12819 VPWR.n1551 VPWR.n1547 0.346131
R12820 VPWR.n1546 VPWR.n1542 0.346131
R12821 VPWR.n1767 VPWR.n1042 0.346131
R12822 VPWR.n1784 VPWR.n1780 0.346131
R12823 VPWR.n1785 VPWR.n1776 0.346131
R12824 VPWR.n1772 VPWR.n1771 0.346131
R12825 VPWR.n2862 VPWR.n2861 0.304571
R12826 VPWR.n2594 VPWR.n55 0.300179
R12827 VPWR.n1118 VPWR.n1113 0.286958
R12828 VPWR.n145 VPWR.n144 0.286958
R12829 VPWR.n157 VPWR.n156 0.286958
R12830 VPWR.n169 VPWR.n168 0.286958
R12831 VPWR.n181 VPWR.n180 0.286958
R12832 VPWR.n193 VPWR.n192 0.286958
R12833 VPWR.n205 VPWR.n204 0.286958
R12834 VPWR.n217 VPWR.n216 0.286958
R12835 VPWR.n229 VPWR.n228 0.286958
R12836 VPWR.n241 VPWR.n240 0.286958
R12837 VPWR.n253 VPWR.n252 0.286958
R12838 VPWR.n265 VPWR.n264 0.286958
R12839 VPWR.n277 VPWR.n276 0.286958
R12840 VPWR.n283 VPWR.n102 0.286958
R12841 VPWR.n111 VPWR.n110 0.286958
R12842 VPWR.n133 VPWR.n132 0.286958
R12843 VPWR.n122 VPWR.n121 0.286958
R12844 VPWR.n1729 VPWR.n1066 0.286958
R12845 VPWR.n1724 VPWR.n1723 0.286958
R12846 VPWR.n1712 VPWR.n1711 0.286958
R12847 VPWR.n1702 VPWR.n1072 0.286958
R12848 VPWR.n1691 VPWR.n1075 0.286958
R12849 VPWR.n1685 VPWR.n1684 0.286958
R12850 VPWR.n1675 VPWR.n1083 0.286958
R12851 VPWR.n1664 VPWR.n1085 0.286958
R12852 VPWR.n1658 VPWR.n1657 0.286958
R12853 VPWR.n1648 VPWR.n1093 0.286958
R12854 VPWR.n1637 VPWR.n1095 0.286958
R12855 VPWR.n1631 VPWR.n1630 0.286958
R12856 VPWR.n1621 VPWR.n1103 0.286958
R12857 VPWR.n1610 VPWR.n1105 0.286958
R12858 VPWR.n1604 VPWR.n1603 0.286958
R12859 VPWR.n55 VPWR 0.2505
R12860 VPWR VPWR.n2481 0.249238
R12861 VPWR.n2472 VPWR 0.249238
R12862 VPWR VPWR.n2471 0.249238
R12863 VPWR.n2385 VPWR 0.249238
R12864 VPWR.n2386 VPWR 0.249238
R12865 VPWR.n2387 VPWR 0.249238
R12866 VPWR.n2388 VPWR 0.249238
R12867 VPWR.n2305 VPWR 0.249238
R12868 VPWR.n2314 VPWR 0.249238
R12869 VPWR.n2315 VPWR 0.249238
R12870 VPWR.n2324 VPWR 0.249238
R12871 VPWR.n2325 VPWR 0.249238
R12872 VPWR.n2383 VPWR 0.249238
R12873 VPWR.n2375 VPWR 0.249238
R12874 VPWR.n2374 VPWR 0.249238
R12875 VPWR.n2365 VPWR 0.249238
R12876 VPWR.n2364 VPWR 0.249238
R12877 VPWR.n2355 VPWR 0.249238
R12878 VPWR.n2354 VPWR 0.249238
R12879 VPWR.n2345 VPWR 0.249238
R12880 VPWR.n2344 VPWR 0.249238
R12881 VPWR.n2335 VPWR 0.249238
R12882 VPWR.n2334 VPWR 0.249238
R12883 VPWR VPWR.n2302 0.249238
R12884 VPWR VPWR.n2301 0.249238
R12885 VPWR VPWR.n2300 0.249238
R12886 VPWR VPWR.n2299 0.249238
R12887 VPWR VPWR.n2298 0.249238
R12888 VPWR VPWR.n2287 0.249238
R12889 VPWR VPWR.n2288 0.249238
R12890 VPWR VPWR.n2289 0.249238
R12891 VPWR VPWR.n2290 0.249238
R12892 VPWR VPWR.n2291 0.249238
R12893 VPWR VPWR.n2292 0.249238
R12894 VPWR VPWR.n2293 0.249238
R12895 VPWR VPWR.n2294 0.249238
R12896 VPWR VPWR.n2295 0.249238
R12897 VPWR VPWR.n2296 0.249238
R12898 VPWR VPWR.n2297 0.249238
R12899 VPWR VPWR.n2285 0.249238
R12900 VPWR.n2276 VPWR 0.249238
R12901 VPWR VPWR.n2275 0.249238
R12902 VPWR.n2266 VPWR 0.249238
R12903 VPWR VPWR.n2265 0.249238
R12904 VPWR.n2207 VPWR 0.249238
R12905 VPWR VPWR.n2215 0.249238
R12906 VPWR.n2216 VPWR 0.249238
R12907 VPWR VPWR.n2225 0.249238
R12908 VPWR.n2226 VPWR 0.249238
R12909 VPWR VPWR.n2235 0.249238
R12910 VPWR.n2236 VPWR 0.249238
R12911 VPWR VPWR.n2245 0.249238
R12912 VPWR.n2246 VPWR 0.249238
R12913 VPWR VPWR.n2255 0.249238
R12914 VPWR.n2256 VPWR 0.249238
R12915 VPWR.n2189 VPWR 0.249238
R12916 VPWR.n2190 VPWR 0.249238
R12917 VPWR.n2191 VPWR 0.249238
R12918 VPWR.n2192 VPWR 0.249238
R12919 VPWR.n2193 VPWR 0.249238
R12920 VPWR.n2204 VPWR 0.249238
R12921 VPWR.n2203 VPWR 0.249238
R12922 VPWR.n2202 VPWR 0.249238
R12923 VPWR.n2201 VPWR 0.249238
R12924 VPWR.n2200 VPWR 0.249238
R12925 VPWR.n2199 VPWR 0.249238
R12926 VPWR.n2198 VPWR 0.249238
R12927 VPWR.n2197 VPWR 0.249238
R12928 VPWR.n2196 VPWR 0.249238
R12929 VPWR.n2195 VPWR 0.249238
R12930 VPWR.n2194 VPWR 0.249238
R12931 VPWR.n2109 VPWR 0.249238
R12932 VPWR.n2118 VPWR 0.249238
R12933 VPWR.n2119 VPWR 0.249238
R12934 VPWR.n2128 VPWR 0.249238
R12935 VPWR.n2129 VPWR 0.249238
R12936 VPWR.n2187 VPWR 0.249238
R12937 VPWR.n2179 VPWR 0.249238
R12938 VPWR.n2178 VPWR 0.249238
R12939 VPWR.n2169 VPWR 0.249238
R12940 VPWR.n2168 VPWR 0.249238
R12941 VPWR.n2159 VPWR 0.249238
R12942 VPWR.n2158 VPWR 0.249238
R12943 VPWR.n2149 VPWR 0.249238
R12944 VPWR.n2148 VPWR 0.249238
R12945 VPWR.n2139 VPWR 0.249238
R12946 VPWR.n2138 VPWR 0.249238
R12947 VPWR VPWR.n2106 0.249238
R12948 VPWR VPWR.n2105 0.249238
R12949 VPWR VPWR.n2104 0.249238
R12950 VPWR VPWR.n2103 0.249238
R12951 VPWR VPWR.n2102 0.249238
R12952 VPWR VPWR.n2091 0.249238
R12953 VPWR VPWR.n2092 0.249238
R12954 VPWR VPWR.n2093 0.249238
R12955 VPWR VPWR.n2094 0.249238
R12956 VPWR VPWR.n2095 0.249238
R12957 VPWR VPWR.n2096 0.249238
R12958 VPWR VPWR.n2097 0.249238
R12959 VPWR VPWR.n2098 0.249238
R12960 VPWR VPWR.n2099 0.249238
R12961 VPWR VPWR.n2100 0.249238
R12962 VPWR VPWR.n2101 0.249238
R12963 VPWR VPWR.n2089 0.249238
R12964 VPWR.n2080 VPWR 0.249238
R12965 VPWR VPWR.n2079 0.249238
R12966 VPWR.n2070 VPWR 0.249238
R12967 VPWR VPWR.n2069 0.249238
R12968 VPWR.n2011 VPWR 0.249238
R12969 VPWR VPWR.n2019 0.249238
R12970 VPWR.n2020 VPWR 0.249238
R12971 VPWR VPWR.n2029 0.249238
R12972 VPWR.n2030 VPWR 0.249238
R12973 VPWR VPWR.n2039 0.249238
R12974 VPWR.n2040 VPWR 0.249238
R12975 VPWR VPWR.n2049 0.249238
R12976 VPWR.n2050 VPWR 0.249238
R12977 VPWR VPWR.n2059 0.249238
R12978 VPWR.n2060 VPWR 0.249238
R12979 VPWR.n1993 VPWR 0.249238
R12980 VPWR.n1994 VPWR 0.249238
R12981 VPWR.n1995 VPWR 0.249238
R12982 VPWR.n1996 VPWR 0.249238
R12983 VPWR.n1997 VPWR 0.249238
R12984 VPWR.n2008 VPWR 0.249238
R12985 VPWR.n2007 VPWR 0.249238
R12986 VPWR.n2006 VPWR 0.249238
R12987 VPWR.n2005 VPWR 0.249238
R12988 VPWR.n2004 VPWR 0.249238
R12989 VPWR.n2003 VPWR 0.249238
R12990 VPWR.n2002 VPWR 0.249238
R12991 VPWR.n2001 VPWR 0.249238
R12992 VPWR.n2000 VPWR 0.249238
R12993 VPWR.n1999 VPWR 0.249238
R12994 VPWR.n1998 VPWR 0.249238
R12995 VPWR.n1913 VPWR 0.249238
R12996 VPWR.n1922 VPWR 0.249238
R12997 VPWR.n1923 VPWR 0.249238
R12998 VPWR.n1932 VPWR 0.249238
R12999 VPWR.n1933 VPWR 0.249238
R13000 VPWR.n1991 VPWR 0.249238
R13001 VPWR.n1983 VPWR 0.249238
R13002 VPWR.n1982 VPWR 0.249238
R13003 VPWR.n1973 VPWR 0.249238
R13004 VPWR.n1972 VPWR 0.249238
R13005 VPWR.n1963 VPWR 0.249238
R13006 VPWR.n1962 VPWR 0.249238
R13007 VPWR.n1953 VPWR 0.249238
R13008 VPWR.n1952 VPWR 0.249238
R13009 VPWR.n1943 VPWR 0.249238
R13010 VPWR.n1942 VPWR 0.249238
R13011 VPWR VPWR.n1910 0.249238
R13012 VPWR VPWR.n1909 0.249238
R13013 VPWR VPWR.n1908 0.249238
R13014 VPWR VPWR.n1907 0.249238
R13015 VPWR VPWR.n1906 0.249238
R13016 VPWR VPWR.n1895 0.249238
R13017 VPWR VPWR.n1896 0.249238
R13018 VPWR VPWR.n1897 0.249238
R13019 VPWR VPWR.n1898 0.249238
R13020 VPWR VPWR.n1899 0.249238
R13021 VPWR VPWR.n1900 0.249238
R13022 VPWR VPWR.n1901 0.249238
R13023 VPWR VPWR.n1902 0.249238
R13024 VPWR VPWR.n1903 0.249238
R13025 VPWR VPWR.n1904 0.249238
R13026 VPWR VPWR.n1905 0.249238
R13027 VPWR.n2400 VPWR 0.249238
R13028 VPWR.n2399 VPWR 0.249238
R13029 VPWR.n2398 VPWR 0.249238
R13030 VPWR.n2397 VPWR 0.249238
R13031 VPWR.n2396 VPWR 0.249238
R13032 VPWR.n2395 VPWR 0.249238
R13033 VPWR.n2394 VPWR 0.249238
R13034 VPWR.n2393 VPWR 0.249238
R13035 VPWR.n2392 VPWR 0.249238
R13036 VPWR.n2391 VPWR 0.249238
R13037 VPWR.n2390 VPWR 0.249238
R13038 VPWR.n2389 VPWR 0.249238
R13039 VPWR VPWR.n1893 0.249238
R13040 VPWR.n1884 VPWR 0.249238
R13041 VPWR VPWR.n1883 0.249238
R13042 VPWR.n1874 VPWR 0.249238
R13043 VPWR VPWR.n1873 0.249238
R13044 VPWR.n1864 VPWR 0.249238
R13045 VPWR.n1815 VPWR 0.249238
R13046 VPWR VPWR.n1823 0.249238
R13047 VPWR.n1824 VPWR 0.249238
R13048 VPWR VPWR.n1833 0.249238
R13049 VPWR.n1834 VPWR 0.249238
R13050 VPWR VPWR.n1843 0.249238
R13051 VPWR.n1844 VPWR 0.249238
R13052 VPWR VPWR.n1853 0.249238
R13053 VPWR.n1854 VPWR 0.249238
R13054 VPWR VPWR.n1863 0.249238
R13055 VPWR.n2403 VPWR 0.249238
R13056 VPWR VPWR.n2411 0.249238
R13057 VPWR.n2412 VPWR 0.249238
R13058 VPWR VPWR.n2421 0.249238
R13059 VPWR.n2422 VPWR 0.249238
R13060 VPWR VPWR.n2431 0.249238
R13061 VPWR.n2432 VPWR 0.249238
R13062 VPWR VPWR.n2441 0.249238
R13063 VPWR.n2442 VPWR 0.249238
R13064 VPWR VPWR.n2451 0.249238
R13065 VPWR.n2452 VPWR 0.249238
R13066 VPWR VPWR.n2461 0.249238
R13067 VPWR.n2462 VPWR 0.249238
R13068 VPWR.n1797 VPWR 0.249238
R13069 VPWR.n1798 VPWR 0.249238
R13070 VPWR.n1799 VPWR 0.249238
R13071 VPWR.n1800 VPWR 0.249238
R13072 VPWR.n1801 VPWR 0.249238
R13073 VPWR.n1802 VPWR 0.249238
R13074 VPWR.n1803 VPWR 0.249238
R13075 VPWR.n1804 VPWR 0.249238
R13076 VPWR.n1805 VPWR 0.249238
R13077 VPWR.n1812 VPWR 0.249238
R13078 VPWR.n1811 VPWR 0.249238
R13079 VPWR.n1810 VPWR 0.249238
R13080 VPWR.n1809 VPWR 0.249238
R13081 VPWR.n1808 VPWR 0.249238
R13082 VPWR.n1807 VPWR 0.249238
R13083 VPWR.n1806 VPWR 0.249238
R13084 VPWR VPWR.n2498 0.249238
R13085 VPWR VPWR.n2497 0.249238
R13086 VPWR VPWR.n2496 0.249238
R13087 VPWR VPWR.n2495 0.249238
R13088 VPWR VPWR.n2494 0.249238
R13089 VPWR VPWR.n2493 0.249238
R13090 VPWR VPWR.n2492 0.249238
R13091 VPWR VPWR.n2491 0.249238
R13092 VPWR VPWR.n2490 0.249238
R13093 VPWR VPWR.n2489 0.249238
R13094 VPWR VPWR.n2488 0.249238
R13095 VPWR VPWR.n2483 0.249238
R13096 VPWR VPWR.n2484 0.249238
R13097 VPWR VPWR.n2485 0.249238
R13098 VPWR VPWR.n2486 0.249238
R13099 VPWR VPWR.n2487 0.249238
R13100 VPWR.n2501 VPWR 0.249238
R13101 VPWR.n2512 VPWR 0.249238
R13102 VPWR.n2513 VPWR 0.249238
R13103 VPWR.n2524 VPWR 0.249238
R13104 VPWR.n2525 VPWR 0.249238
R13105 VPWR.n2536 VPWR 0.249238
R13106 VPWR.n2537 VPWR 0.249238
R13107 VPWR.n2548 VPWR 0.249238
R13108 VPWR.n2549 VPWR 0.249238
R13109 VPWR.n2560 VPWR 0.249238
R13110 VPWR.n2561 VPWR 0.249238
R13111 VPWR.n2572 VPWR 0.249238
R13112 VPWR.n2573 VPWR 0.249238
R13113 VPWR.n2584 VPWR 0.249238
R13114 VPWR.n2585 VPWR 0.249238
R13115 VPWR.n2595 VPWR 0.249238
R13116 VPWR VPWR.n1055 0.249238
R13117 VPWR VPWR.n1056 0.249238
R13118 VPWR VPWR.n1754 0.249238
R13119 VPWR.n1755 VPWR 0.249238
R13120 VPWR VPWR.n1529 0.249238
R13121 VPWR.n1530 VPWR 0.249238
R13122 VPWR.n1528 VPWR 0.249238
R13123 VPWR.n1527 VPWR 0.249238
R13124 VPWR.n1514 VPWR 0.249238
R13125 VPWR.n1513 VPWR 0.249238
R13126 VPWR.n1500 VPWR 0.249238
R13127 VPWR.n1499 VPWR 0.249238
R13128 VPWR.n1487 VPWR 0.249238
R13129 VPWR VPWR.n1587 0.249238
R13130 VPWR.n1588 VPWR 0.249238
R13131 VPWR VPWR.n1448 0.249238
R13132 VPWR.n2861 VPWR.n2815 0.245065
R13133 VPWR.n2813 VPWR.n2797 0.213567
R13134 VPWR.n2797 VPWR.n2778 0.213567
R13135 VPWR.n2778 VPWR.n2758 0.213567
R13136 VPWR.n2758 VPWR.n2739 0.213567
R13137 VPWR.n2739 VPWR.n2703 0.213567
R13138 VPWR.n2703 VPWR.n2665 0.213567
R13139 VPWR.n2665 VPWR.n2628 0.213567
R13140 VPWR.n1446 VPWR.n1414 0.213567
R13141 VPWR.n1414 VPWR.n1376 0.213567
R13142 VPWR.n1376 VPWR.n1337 0.213567
R13143 VPWR.n1337 VPWR.n1302 0.213567
R13144 VPWR.n1302 VPWR.n1279 0.213567
R13145 VPWR.n1279 VPWR.n1255 0.213567
R13146 VPWR.n1255 VPWR.n19 0.213567
R13147 VPWR VPWR.n2862 0.204304
R13148 VPWR.n1449 VPWR.n1447 0.179202
R13149 VPWR.n1450 VPWR.n1449 0.154425
R13150 VPWR.n1450 VPWR.n930 0.154425
R13151 VPWR.n1894 VPWR.n930 0.154425
R13152 VPWR.n1911 VPWR.n1894 0.154425
R13153 VPWR.n1912 VPWR.n1911 0.154425
R13154 VPWR.n1912 VPWR.n738 0.154425
R13155 VPWR.n2090 VPWR.n738 0.154425
R13156 VPWR.n2107 VPWR.n2090 0.154425
R13157 VPWR.n2108 VPWR.n2107 0.154425
R13158 VPWR.n2108 VPWR.n546 0.154425
R13159 VPWR.n2286 VPWR.n546 0.154425
R13160 VPWR.n2303 VPWR.n2286 0.154425
R13161 VPWR.n2304 VPWR.n2303 0.154425
R13162 VPWR.n2304 VPWR.n354 0.154425
R13163 VPWR.n2482 VPWR.n354 0.154425
R13164 VPWR.n2499 VPWR.n2482 0.154425
R13165 VPWR.n2500 VPWR.n2499 0.154425
R13166 VPWR.n1796 VPWR.n1026 0.154425
R13167 VPWR.n1813 VPWR.n1796 0.154425
R13168 VPWR.n1814 VPWR.n1813 0.154425
R13169 VPWR.n1814 VPWR.n834 0.154425
R13170 VPWR.n1992 VPWR.n834 0.154425
R13171 VPWR.n2009 VPWR.n1992 0.154425
R13172 VPWR.n2010 VPWR.n2009 0.154425
R13173 VPWR.n2010 VPWR.n642 0.154425
R13174 VPWR.n2188 VPWR.n642 0.154425
R13175 VPWR.n2205 VPWR.n2188 0.154425
R13176 VPWR.n2206 VPWR.n2205 0.154425
R13177 VPWR.n2206 VPWR.n450 0.154425
R13178 VPWR.n2384 VPWR.n450 0.154425
R13179 VPWR.n2401 VPWR.n2384 0.154425
R13180 VPWR.n2402 VPWR.n2401 0.154425
R13181 VPWR.n2402 VPWR.n21 0.154425
R13182 VPWR.n2596 VPWR.n21 0.154425
R13183 VPWR.n8 VPWR.n7 0.147771
R13184 VPWR.n1243 VPWR.n1242 0.147771
R13185 VPWR.n1266 VPWR.n1265 0.147771
R13186 VPWR.n1290 VPWR.n1289 0.147771
R13187 VPWR.n1113 VPWR 0.135917
R13188 VPWR.n145 VPWR 0.135917
R13189 VPWR.n157 VPWR 0.135917
R13190 VPWR.n169 VPWR 0.135917
R13191 VPWR.n181 VPWR 0.135917
R13192 VPWR.n193 VPWR 0.135917
R13193 VPWR.n205 VPWR 0.135917
R13194 VPWR.n217 VPWR 0.135917
R13195 VPWR.n229 VPWR 0.135917
R13196 VPWR.n241 VPWR 0.135917
R13197 VPWR.n253 VPWR 0.135917
R13198 VPWR.n265 VPWR 0.135917
R13199 VPWR.n277 VPWR 0.135917
R13200 VPWR.n102 VPWR 0.135917
R13201 VPWR.n111 VPWR 0.135917
R13202 VPWR.n133 VPWR 0.135917
R13203 VPWR.n122 VPWR 0.135917
R13204 VPWR.n1066 VPWR 0.135917
R13205 VPWR.n1724 VPWR 0.135917
R13206 VPWR.n1712 VPWR 0.135917
R13207 VPWR.n1072 VPWR 0.135917
R13208 VPWR.n1075 VPWR 0.135917
R13209 VPWR.n1685 VPWR 0.135917
R13210 VPWR.n1083 VPWR 0.135917
R13211 VPWR.n1085 VPWR 0.135917
R13212 VPWR.n1658 VPWR 0.135917
R13213 VPWR.n1093 VPWR 0.135917
R13214 VPWR.n1095 VPWR 0.135917
R13215 VPWR.n1631 VPWR 0.135917
R13216 VPWR.n1103 VPWR 0.135917
R13217 VPWR.n1105 VPWR 0.135917
R13218 VPWR.n1604 VPWR 0.135917
R13219 VPWR.n2863 VPWR.n2814 0.127988
R13220 VPWR.n2825 VPWR.n2816 0.1255
R13221 VPWR.n2831 VPWR.n2816 0.1255
R13222 VPWR.n18 VPWR.n0 0.120292
R13223 VPWR.n14 VPWR.n0 0.120292
R13224 VPWR.n9 VPWR.n8 0.120292
R13225 VPWR.n1254 VPWR.n1233 0.120292
R13226 VPWR.n1250 VPWR.n1233 0.120292
R13227 VPWR.n1244 VPWR.n1243 0.120292
R13228 VPWR.n1278 VPWR.n1256 0.120292
R13229 VPWR.n1273 VPWR.n1256 0.120292
R13230 VPWR.n1267 VPWR.n1266 0.120292
R13231 VPWR.n1301 VPWR.n1280 0.120292
R13232 VPWR.n1297 VPWR.n1280 0.120292
R13233 VPWR.n1291 VPWR.n1290 0.120292
R13234 VPWR.n1333 VPWR.n1332 0.120292
R13235 VPWR.n1326 VPWR.n1305 0.120292
R13236 VPWR.n1319 VPWR.n1305 0.120292
R13237 VPWR.n1319 VPWR.n1318 0.120292
R13238 VPWR.n1317 VPWR.n1309 0.120292
R13239 VPWR.n1312 VPWR.n1309 0.120292
R13240 VPWR.n1312 VPWR.n1311 0.120292
R13241 VPWR.n1371 VPWR.n1370 0.120292
R13242 VPWR.n1364 VPWR.n1363 0.120292
R13243 VPWR.n1363 VPWR.n1340 0.120292
R13244 VPWR.n1356 VPWR.n1340 0.120292
R13245 VPWR.n1356 VPWR.n1355 0.120292
R13246 VPWR.n1355 VPWR.n1354 0.120292
R13247 VPWR.n1354 VPWR.n1342 0.120292
R13248 VPWR.n1348 VPWR.n1342 0.120292
R13249 VPWR.n1348 VPWR.n1347 0.120292
R13250 VPWR.n1410 VPWR.n1409 0.120292
R13251 VPWR.n1403 VPWR.n1402 0.120292
R13252 VPWR.n1402 VPWR.n1379 0.120292
R13253 VPWR.n1395 VPWR.n1379 0.120292
R13254 VPWR.n1395 VPWR.n1394 0.120292
R13255 VPWR.n1394 VPWR.n1393 0.120292
R13256 VPWR.n1393 VPWR.n1381 0.120292
R13257 VPWR.n1387 VPWR.n1381 0.120292
R13258 VPWR.n1387 VPWR.n1386 0.120292
R13259 VPWR.n1440 VPWR.n1439 0.120292
R13260 VPWR.n1439 VPWR.n1416 0.120292
R13261 VPWR.n1432 VPWR.n1416 0.120292
R13262 VPWR.n1432 VPWR.n1431 0.120292
R13263 VPWR.n1431 VPWR.n1430 0.120292
R13264 VPWR.n1430 VPWR.n1418 0.120292
R13265 VPWR.n1424 VPWR.n1418 0.120292
R13266 VPWR.n1424 VPWR.n1423 0.120292
R13267 VPWR.n2812 VPWR.n2798 0.120292
R13268 VPWR.n2796 VPWR.n2779 0.120292
R13269 VPWR.n2777 VPWR.n2759 0.120292
R13270 VPWR.n2757 VPWR.n2740 0.120292
R13271 VPWR.n2719 VPWR.n2718 0.120292
R13272 VPWR.n2720 VPWR.n2719 0.120292
R13273 VPWR.n2720 VPWR.n2711 0.120292
R13274 VPWR.n2725 VPWR.n2711 0.120292
R13275 VPWR.n2726 VPWR.n2725 0.120292
R13276 VPWR.n2726 VPWR.n2707 0.120292
R13277 VPWR.n2732 VPWR.n2707 0.120292
R13278 VPWR.n2734 VPWR.n2704 0.120292
R13279 VPWR.n2738 VPWR.n2704 0.120292
R13280 VPWR.n2683 VPWR.n2682 0.120292
R13281 VPWR.n2684 VPWR.n2683 0.120292
R13282 VPWR.n2684 VPWR.n2673 0.120292
R13283 VPWR.n2689 VPWR.n2673 0.120292
R13284 VPWR.n2690 VPWR.n2689 0.120292
R13285 VPWR.n2690 VPWR.n2669 0.120292
R13286 VPWR.n2695 VPWR.n2669 0.120292
R13287 VPWR.n2697 VPWR.n2666 0.120292
R13288 VPWR.n2702 VPWR.n2666 0.120292
R13289 VPWR.n2646 VPWR.n2645 0.120292
R13290 VPWR.n2647 VPWR.n2646 0.120292
R13291 VPWR.n2647 VPWR.n2636 0.120292
R13292 VPWR.n2652 VPWR.n2636 0.120292
R13293 VPWR.n2653 VPWR.n2652 0.120292
R13294 VPWR.n2653 VPWR.n2632 0.120292
R13295 VPWR.n2658 VPWR.n2632 0.120292
R13296 VPWR.n2660 VPWR.n2629 0.120292
R13297 VPWR.n2664 VPWR.n2629 0.120292
R13298 VPWR.n2608 VPWR.n2604 0.120292
R13299 VPWR.n2616 VPWR.n2604 0.120292
R13300 VPWR.n2617 VPWR.n2616 0.120292
R13301 VPWR.n2618 VPWR.n2617 0.120292
R13302 VPWR.n2618 VPWR.n2600 0.120292
R13303 VPWR.n2623 VPWR.n2600 0.120292
R13304 VPWR.n2624 VPWR.n2623 0.120292
R13305 VPWR.n1605 VPWR 0.118556
R13306 VPWR.n1108 VPWR 0.118556
R13307 VPWR.n1619 VPWR 0.118556
R13308 VPWR.n1632 VPWR 0.118556
R13309 VPWR.n1098 VPWR 0.118556
R13310 VPWR.n1646 VPWR 0.118556
R13311 VPWR.n1659 VPWR 0.118556
R13312 VPWR.n1088 VPWR 0.118556
R13313 VPWR.n1673 VPWR 0.118556
R13314 VPWR.n1686 VPWR 0.118556
R13315 VPWR.n1078 VPWR 0.118556
R13316 VPWR.n1700 VPWR 0.118556
R13317 VPWR.n1713 VPWR 0.118556
R13318 VPWR.n1725 VPWR 0.118556
R13319 VPWR VPWR.n1112 0.118556
R13320 VPWR.n1067 VPWR 0.118556
R13321 VPWR.n123 VPWR 0.118556
R13322 VPWR.n112 VPWR 0.118556
R13323 VPWR.n103 VPWR 0.118556
R13324 VPWR.n278 VPWR 0.118556
R13325 VPWR.n266 VPWR 0.118556
R13326 VPWR.n254 VPWR 0.118556
R13327 VPWR.n242 VPWR 0.118556
R13328 VPWR.n230 VPWR 0.118556
R13329 VPWR.n218 VPWR 0.118556
R13330 VPWR.n206 VPWR 0.118556
R13331 VPWR.n194 VPWR 0.118556
R13332 VPWR.n182 VPWR 0.118556
R13333 VPWR.n170 VPWR 0.118556
R13334 VPWR.n158 VPWR 0.118556
R13335 VPWR.n146 VPWR 0.118556
R13336 VPWR.n134 VPWR 0.118556
R13337 VPWR.n1765 VPWR.n1044 0.108238
R13338 VPWR.n1541 VPWR.n1143 0.108238
R13339 VPWR.n1540 VPWR.n1142 0.108238
R13340 VPWR.n1524 VPWR.n1141 0.108238
R13341 VPWR.n1516 VPWR.n1140 0.108238
R13342 VPWR.n1510 VPWR.n1139 0.108238
R13343 VPWR.n1502 VPWR.n1138 0.108238
R13344 VPWR.n1496 VPWR.n1137 0.108238
R13345 VPWR.n1583 VPWR.n1132 0.108238
R13346 VPWR.n1584 VPWR.n1131 0.108238
R13347 VPWR.n1463 VPWR.n1452 0.108238
R13348 VPWR.n1464 VPWR.n1451 0.108238
R13349 VPWR.n1795 VPWR.n1027 0.108238
R13350 VPWR.n1766 VPWR.n1043 0.108238
R13351 VPWR.n1744 VPWR.n1038 0.108238
R13352 VPWR.n1787 VPWR.n1786 0.108238
R13353 VPWR.n2481 VPWR 0.100405
R13354 VPWR.n2472 VPWR 0.100405
R13355 VPWR VPWR.n2385 0.100405
R13356 VPWR VPWR.n2386 0.100405
R13357 VPWR VPWR.n2387 0.100405
R13358 VPWR.n2305 VPWR 0.100405
R13359 VPWR VPWR.n2314 0.100405
R13360 VPWR.n2315 VPWR 0.100405
R13361 VPWR VPWR.n2324 0.100405
R13362 VPWR.n2375 VPWR 0.100405
R13363 VPWR VPWR.n2374 0.100405
R13364 VPWR.n2365 VPWR 0.100405
R13365 VPWR VPWR.n2364 0.100405
R13366 VPWR.n2355 VPWR 0.100405
R13367 VPWR VPWR.n2354 0.100405
R13368 VPWR.n2345 VPWR 0.100405
R13369 VPWR VPWR.n2344 0.100405
R13370 VPWR.n2335 VPWR 0.100405
R13371 VPWR VPWR.n2334 0.100405
R13372 VPWR.n2325 VPWR 0.100405
R13373 VPWR.n2302 VPWR 0.100405
R13374 VPWR.n2301 VPWR 0.100405
R13375 VPWR.n2300 VPWR 0.100405
R13376 VPWR.n2299 VPWR 0.100405
R13377 VPWR.n2288 VPWR 0.100405
R13378 VPWR.n2289 VPWR 0.100405
R13379 VPWR.n2290 VPWR 0.100405
R13380 VPWR.n2291 VPWR 0.100405
R13381 VPWR.n2292 VPWR 0.100405
R13382 VPWR.n2293 VPWR 0.100405
R13383 VPWR.n2294 VPWR 0.100405
R13384 VPWR.n2295 VPWR 0.100405
R13385 VPWR.n2296 VPWR 0.100405
R13386 VPWR.n2297 VPWR 0.100405
R13387 VPWR.n2298 VPWR 0.100405
R13388 VPWR.n2285 VPWR 0.100405
R13389 VPWR.n2276 VPWR 0.100405
R13390 VPWR.n2275 VPWR 0.100405
R13391 VPWR.n2266 VPWR 0.100405
R13392 VPWR.n2215 VPWR 0.100405
R13393 VPWR.n2216 VPWR 0.100405
R13394 VPWR.n2225 VPWR 0.100405
R13395 VPWR.n2226 VPWR 0.100405
R13396 VPWR.n2235 VPWR 0.100405
R13397 VPWR.n2236 VPWR 0.100405
R13398 VPWR.n2245 VPWR 0.100405
R13399 VPWR.n2246 VPWR 0.100405
R13400 VPWR.n2255 VPWR 0.100405
R13401 VPWR.n2256 VPWR 0.100405
R13402 VPWR.n2265 VPWR 0.100405
R13403 VPWR VPWR.n2189 0.100405
R13404 VPWR VPWR.n2190 0.100405
R13405 VPWR VPWR.n2191 0.100405
R13406 VPWR VPWR.n2192 0.100405
R13407 VPWR VPWR.n2203 0.100405
R13408 VPWR VPWR.n2202 0.100405
R13409 VPWR VPWR.n2201 0.100405
R13410 VPWR VPWR.n2200 0.100405
R13411 VPWR VPWR.n2199 0.100405
R13412 VPWR VPWR.n2198 0.100405
R13413 VPWR VPWR.n2197 0.100405
R13414 VPWR VPWR.n2196 0.100405
R13415 VPWR VPWR.n2195 0.100405
R13416 VPWR VPWR.n2194 0.100405
R13417 VPWR VPWR.n2193 0.100405
R13418 VPWR.n2109 VPWR 0.100405
R13419 VPWR VPWR.n2118 0.100405
R13420 VPWR.n2119 VPWR 0.100405
R13421 VPWR VPWR.n2128 0.100405
R13422 VPWR.n2179 VPWR 0.100405
R13423 VPWR VPWR.n2178 0.100405
R13424 VPWR.n2169 VPWR 0.100405
R13425 VPWR VPWR.n2168 0.100405
R13426 VPWR.n2159 VPWR 0.100405
R13427 VPWR VPWR.n2158 0.100405
R13428 VPWR.n2149 VPWR 0.100405
R13429 VPWR VPWR.n2148 0.100405
R13430 VPWR.n2139 VPWR 0.100405
R13431 VPWR VPWR.n2138 0.100405
R13432 VPWR.n2129 VPWR 0.100405
R13433 VPWR.n2106 VPWR 0.100405
R13434 VPWR.n2105 VPWR 0.100405
R13435 VPWR.n2104 VPWR 0.100405
R13436 VPWR.n2103 VPWR 0.100405
R13437 VPWR.n2092 VPWR 0.100405
R13438 VPWR.n2093 VPWR 0.100405
R13439 VPWR.n2094 VPWR 0.100405
R13440 VPWR.n2095 VPWR 0.100405
R13441 VPWR.n2096 VPWR 0.100405
R13442 VPWR.n2097 VPWR 0.100405
R13443 VPWR.n2098 VPWR 0.100405
R13444 VPWR.n2099 VPWR 0.100405
R13445 VPWR.n2100 VPWR 0.100405
R13446 VPWR.n2101 VPWR 0.100405
R13447 VPWR.n2102 VPWR 0.100405
R13448 VPWR.n2089 VPWR 0.100405
R13449 VPWR.n2080 VPWR 0.100405
R13450 VPWR.n2079 VPWR 0.100405
R13451 VPWR.n2070 VPWR 0.100405
R13452 VPWR.n2019 VPWR 0.100405
R13453 VPWR.n2020 VPWR 0.100405
R13454 VPWR.n2029 VPWR 0.100405
R13455 VPWR.n2030 VPWR 0.100405
R13456 VPWR.n2039 VPWR 0.100405
R13457 VPWR.n2040 VPWR 0.100405
R13458 VPWR.n2049 VPWR 0.100405
R13459 VPWR.n2050 VPWR 0.100405
R13460 VPWR.n2059 VPWR 0.100405
R13461 VPWR.n2060 VPWR 0.100405
R13462 VPWR.n2069 VPWR 0.100405
R13463 VPWR VPWR.n1993 0.100405
R13464 VPWR VPWR.n1994 0.100405
R13465 VPWR VPWR.n1995 0.100405
R13466 VPWR VPWR.n1996 0.100405
R13467 VPWR VPWR.n2007 0.100405
R13468 VPWR VPWR.n2006 0.100405
R13469 VPWR VPWR.n2005 0.100405
R13470 VPWR VPWR.n2004 0.100405
R13471 VPWR VPWR.n2003 0.100405
R13472 VPWR VPWR.n2002 0.100405
R13473 VPWR VPWR.n2001 0.100405
R13474 VPWR VPWR.n2000 0.100405
R13475 VPWR VPWR.n1999 0.100405
R13476 VPWR VPWR.n1998 0.100405
R13477 VPWR VPWR.n1997 0.100405
R13478 VPWR.n1913 VPWR 0.100405
R13479 VPWR VPWR.n1922 0.100405
R13480 VPWR.n1923 VPWR 0.100405
R13481 VPWR VPWR.n1932 0.100405
R13482 VPWR.n1983 VPWR 0.100405
R13483 VPWR VPWR.n1982 0.100405
R13484 VPWR.n1973 VPWR 0.100405
R13485 VPWR VPWR.n1972 0.100405
R13486 VPWR.n1963 VPWR 0.100405
R13487 VPWR VPWR.n1962 0.100405
R13488 VPWR.n1953 VPWR 0.100405
R13489 VPWR VPWR.n1952 0.100405
R13490 VPWR.n1943 VPWR 0.100405
R13491 VPWR VPWR.n1942 0.100405
R13492 VPWR.n1933 VPWR 0.100405
R13493 VPWR.n1910 VPWR 0.100405
R13494 VPWR.n1909 VPWR 0.100405
R13495 VPWR.n1908 VPWR 0.100405
R13496 VPWR.n1907 VPWR 0.100405
R13497 VPWR.n1896 VPWR 0.100405
R13498 VPWR.n1897 VPWR 0.100405
R13499 VPWR.n1898 VPWR 0.100405
R13500 VPWR.n1899 VPWR 0.100405
R13501 VPWR.n1900 VPWR 0.100405
R13502 VPWR.n1901 VPWR 0.100405
R13503 VPWR.n1902 VPWR 0.100405
R13504 VPWR.n1903 VPWR 0.100405
R13505 VPWR.n1904 VPWR 0.100405
R13506 VPWR.n1905 VPWR 0.100405
R13507 VPWR.n1906 VPWR 0.100405
R13508 VPWR VPWR.n2399 0.100405
R13509 VPWR VPWR.n2398 0.100405
R13510 VPWR VPWR.n2397 0.100405
R13511 VPWR VPWR.n2396 0.100405
R13512 VPWR VPWR.n2395 0.100405
R13513 VPWR VPWR.n2394 0.100405
R13514 VPWR VPWR.n2393 0.100405
R13515 VPWR VPWR.n2392 0.100405
R13516 VPWR VPWR.n2391 0.100405
R13517 VPWR VPWR.n2390 0.100405
R13518 VPWR VPWR.n2389 0.100405
R13519 VPWR VPWR.n2388 0.100405
R13520 VPWR.n1893 VPWR 0.100405
R13521 VPWR.n1884 VPWR 0.100405
R13522 VPWR.n1883 VPWR 0.100405
R13523 VPWR.n1874 VPWR 0.100405
R13524 VPWR.n1873 VPWR 0.100405
R13525 VPWR.n1823 VPWR 0.100405
R13526 VPWR.n1824 VPWR 0.100405
R13527 VPWR.n1833 VPWR 0.100405
R13528 VPWR.n1834 VPWR 0.100405
R13529 VPWR.n1843 VPWR 0.100405
R13530 VPWR.n1844 VPWR 0.100405
R13531 VPWR.n1853 VPWR 0.100405
R13532 VPWR.n1854 VPWR 0.100405
R13533 VPWR.n1863 VPWR 0.100405
R13534 VPWR.n1864 VPWR 0.100405
R13535 VPWR.n2411 VPWR 0.100405
R13536 VPWR.n2412 VPWR 0.100405
R13537 VPWR.n2421 VPWR 0.100405
R13538 VPWR.n2422 VPWR 0.100405
R13539 VPWR.n2431 VPWR 0.100405
R13540 VPWR.n2432 VPWR 0.100405
R13541 VPWR.n2441 VPWR 0.100405
R13542 VPWR.n2442 VPWR 0.100405
R13543 VPWR.n2451 VPWR 0.100405
R13544 VPWR.n2452 VPWR 0.100405
R13545 VPWR.n2461 VPWR 0.100405
R13546 VPWR.n2462 VPWR 0.100405
R13547 VPWR.n2471 VPWR 0.100405
R13548 VPWR VPWR.n1797 0.100405
R13549 VPWR VPWR.n1798 0.100405
R13550 VPWR VPWR.n1799 0.100405
R13551 VPWR VPWR.n1800 0.100405
R13552 VPWR VPWR.n1801 0.100405
R13553 VPWR VPWR.n1802 0.100405
R13554 VPWR VPWR.n1803 0.100405
R13555 VPWR VPWR.n1804 0.100405
R13556 VPWR VPWR.n1811 0.100405
R13557 VPWR VPWR.n1810 0.100405
R13558 VPWR VPWR.n1809 0.100405
R13559 VPWR VPWR.n1808 0.100405
R13560 VPWR VPWR.n1807 0.100405
R13561 VPWR VPWR.n1806 0.100405
R13562 VPWR VPWR.n1805 0.100405
R13563 VPWR.n2498 VPWR 0.100405
R13564 VPWR.n2497 VPWR 0.100405
R13565 VPWR.n2496 VPWR 0.100405
R13566 VPWR.n2495 VPWR 0.100405
R13567 VPWR.n2494 VPWR 0.100405
R13568 VPWR.n2493 VPWR 0.100405
R13569 VPWR.n2492 VPWR 0.100405
R13570 VPWR.n2491 VPWR 0.100405
R13571 VPWR.n2490 VPWR 0.100405
R13572 VPWR.n2489 VPWR 0.100405
R13573 VPWR.n2484 VPWR 0.100405
R13574 VPWR.n2485 VPWR 0.100405
R13575 VPWR.n2486 VPWR 0.100405
R13576 VPWR.n2487 VPWR 0.100405
R13577 VPWR.n2488 VPWR 0.100405
R13578 VPWR.n1143 VPWR 0.100405
R13579 VPWR VPWR.n1540 0.100405
R13580 VPWR.n1524 VPWR 0.100405
R13581 VPWR.n1516 VPWR 0.100405
R13582 VPWR.n1510 VPWR 0.100405
R13583 VPWR.n1502 VPWR 0.100405
R13584 VPWR.n1496 VPWR 0.100405
R13585 VPWR VPWR.n1132 0.100405
R13586 VPWR.n1584 VPWR 0.100405
R13587 VPWR.n1452 VPWR 0.100405
R13588 VPWR.n1464 VPWR 0.100405
R13589 VPWR.n1043 VPWR 0.100405
R13590 VPWR.n1744 VPWR 0.100405
R13591 VPWR.n1787 VPWR 0.100405
R13592 VPWR VPWR.n1765 0.100405
R13593 VPWR.n2501 VPWR 0.100405
R13594 VPWR VPWR.n2512 0.100405
R13595 VPWR.n2513 VPWR 0.100405
R13596 VPWR VPWR.n2524 0.100405
R13597 VPWR.n2525 VPWR 0.100405
R13598 VPWR VPWR.n2536 0.100405
R13599 VPWR.n2537 VPWR 0.100405
R13600 VPWR VPWR.n2548 0.100405
R13601 VPWR.n2549 VPWR 0.100405
R13602 VPWR VPWR.n2560 0.100405
R13603 VPWR.n2561 VPWR 0.100405
R13604 VPWR VPWR.n2572 0.100405
R13605 VPWR.n2573 VPWR 0.100405
R13606 VPWR VPWR.n2584 0.100405
R13607 VPWR.n2585 VPWR 0.100405
R13608 VPWR.n1056 VPWR 0.100405
R13609 VPWR.n1754 VPWR 0.100405
R13610 VPWR.n1755 VPWR 0.100405
R13611 VPWR.n1529 VPWR 0.100405
R13612 VPWR.n1530 VPWR 0.100405
R13613 VPWR VPWR.n1528 0.100405
R13614 VPWR VPWR.n1527 0.100405
R13615 VPWR.n1514 VPWR 0.100405
R13616 VPWR VPWR.n1513 0.100405
R13617 VPWR.n1500 VPWR 0.100405
R13618 VPWR VPWR.n1499 0.100405
R13619 VPWR.n1487 VPWR 0.100405
R13620 VPWR.n1587 VPWR 0.100405
R13621 VPWR.n1588 VPWR 0.100405
R13622 VPWR.n1448 VPWR 0.100405
R13623 VPWR VPWR.n2798 0.0994583
R13624 VPWR VPWR.n2779 0.0994583
R13625 VPWR VPWR.n1326 0.0981562
R13626 VPWR.n1371 VPWR 0.0981562
R13627 VPWR.n1410 VPWR 0.0981562
R13628 VPWR.n9 VPWR 0.0968542
R13629 VPWR.n1244 VPWR 0.0968542
R13630 VPWR.n1267 VPWR 0.0968542
R13631 VPWR.n1291 VPWR 0.0968542
R13632 VPWR.n1333 VPWR 0.0968542
R13633 VPWR VPWR.n2759 0.0968542
R13634 VPWR VPWR.n2740 0.0968542
R13635 VPWR.n2718 VPWR 0.0968542
R13636 VPWR.n2682 VPWR 0.0968542
R13637 VPWR.n2645 VPWR 0.0968542
R13638 VPWR.n2608 VPWR 0.0968542
R13639 VPWR VPWR.n1044 0.0945
R13640 VPWR.n1541 VPWR 0.0945
R13641 VPWR VPWR.n1142 0.0945
R13642 VPWR VPWR.n1141 0.0945
R13643 VPWR VPWR.n1140 0.0945
R13644 VPWR VPWR.n1139 0.0945
R13645 VPWR VPWR.n1138 0.0945
R13646 VPWR.n1137 VPWR 0.0945
R13647 VPWR VPWR.n1583 0.0945
R13648 VPWR VPWR.n1131 0.0945
R13649 VPWR VPWR.n1463 0.0945
R13650 VPWR.n1451 VPWR 0.0945
R13651 VPWR VPWR.n1038 0.0945
R13652 VPWR.n1786 VPWR 0.0945
R13653 VPWR VPWR.n1027 0.0945
R13654 VPWR.n1766 VPWR 0.0945
R13655 VPWR.n1117 VPWR 0.093504
R13656 VPWR.n109 VPWR 0.093504
R13657 VPWR.n143 VPWR 0.093504
R13658 VPWR.n155 VPWR 0.093504
R13659 VPWR.n167 VPWR 0.093504
R13660 VPWR.n179 VPWR 0.093504
R13661 VPWR.n191 VPWR 0.093504
R13662 VPWR.n203 VPWR 0.093504
R13663 VPWR.n215 VPWR 0.093504
R13664 VPWR.n227 VPWR 0.093504
R13665 VPWR.n239 VPWR 0.093504
R13666 VPWR.n251 VPWR 0.093504
R13667 VPWR.n263 VPWR 0.093504
R13668 VPWR.n275 VPWR 0.093504
R13669 VPWR VPWR.n285 0.093504
R13670 VPWR.n131 VPWR 0.093504
R13671 VPWR.n120 VPWR 0.093504
R13672 VPWR VPWR.n1731 0.093504
R13673 VPWR.n1722 VPWR 0.093504
R13674 VPWR.n1710 VPWR 0.093504
R13675 VPWR.n1699 VPWR 0.093504
R13676 VPWR VPWR.n1077 0.093504
R13677 VPWR.n1683 VPWR 0.093504
R13678 VPWR.n1672 VPWR 0.093504
R13679 VPWR VPWR.n1087 0.093504
R13680 VPWR.n1656 VPWR 0.093504
R13681 VPWR.n1645 VPWR 0.093504
R13682 VPWR VPWR.n1097 0.093504
R13683 VPWR.n1629 VPWR 0.093504
R13684 VPWR.n1618 VPWR 0.093504
R13685 VPWR VPWR.n1107 0.093504
R13686 VPWR.n1602 VPWR 0.093504
R13687 VPWR.n2598 VPWR 0.0849042
R13688 VPWR.n1112 VPWR.n1109 0.0845517
R13689 VPWR.n147 VPWR.n146 0.0845517
R13690 VPWR.n159 VPWR.n158 0.0845517
R13691 VPWR.n171 VPWR.n170 0.0845517
R13692 VPWR.n183 VPWR.n182 0.0845517
R13693 VPWR.n195 VPWR.n194 0.0845517
R13694 VPWR.n207 VPWR.n206 0.0845517
R13695 VPWR.n219 VPWR.n218 0.0845517
R13696 VPWR.n231 VPWR.n230 0.0845517
R13697 VPWR.n243 VPWR.n242 0.0845517
R13698 VPWR.n255 VPWR.n254 0.0845517
R13699 VPWR.n267 VPWR.n266 0.0845517
R13700 VPWR.n279 VPWR.n278 0.0845517
R13701 VPWR.n282 VPWR.n103 0.0845517
R13702 VPWR.n113 VPWR.n112 0.0845517
R13703 VPWR.n135 VPWR.n134 0.0845517
R13704 VPWR.n124 VPWR.n123 0.0845517
R13705 VPWR.n1728 VPWR.n1067 0.0845517
R13706 VPWR.n1726 VPWR.n1725 0.0845517
R13707 VPWR.n1714 VPWR.n1713 0.0845517
R13708 VPWR.n1701 VPWR.n1700 0.0845517
R13709 VPWR.n1690 VPWR.n1078 0.0845517
R13710 VPWR.n1687 VPWR.n1686 0.0845517
R13711 VPWR.n1674 VPWR.n1673 0.0845517
R13712 VPWR.n1663 VPWR.n1088 0.0845517
R13713 VPWR.n1660 VPWR.n1659 0.0845517
R13714 VPWR.n1647 VPWR.n1646 0.0845517
R13715 VPWR.n1636 VPWR.n1098 0.0845517
R13716 VPWR.n1633 VPWR.n1632 0.0845517
R13717 VPWR.n1620 VPWR.n1619 0.0845517
R13718 VPWR.n1609 VPWR.n1108 0.0845517
R13719 VPWR.n1606 VPWR.n1605 0.0845517
R13720 VPWR.n1456 VPWR.n1451 0.0740128
R13721 VPWR.n1542 VPWR.n1044 0.071
R13722 VPWR.n1547 VPWR.n1541 0.071
R13723 VPWR.n1552 VPWR.n1142 0.071
R13724 VPWR.n1557 VPWR.n1141 0.071
R13725 VPWR.n1562 VPWR.n1140 0.071
R13726 VPWR.n1567 VPWR.n1139 0.071
R13727 VPWR.n1572 VPWR.n1138 0.071
R13728 VPWR.n1577 VPWR.n1137 0.071
R13729 VPWR.n1583 VPWR.n1582 0.071
R13730 VPWR.n1457 VPWR.n1131 0.071
R13731 VPWR.n1463 VPWR.n1462 0.071
R13732 VPWR.n1772 VPWR.n1038 0.071
R13733 VPWR.n1786 VPWR.n1785 0.071
R13734 VPWR.n1780 VPWR.n1027 0.071
R13735 VPWR.n1767 VPWR.n1766 0.071
R13736 VPWR VPWR.n1115 0.0678077
R13737 VPWR VPWR.n107 0.0678077
R13738 VPWR VPWR.n141 0.0678077
R13739 VPWR VPWR.n153 0.0678077
R13740 VPWR VPWR.n165 0.0678077
R13741 VPWR VPWR.n177 0.0678077
R13742 VPWR VPWR.n189 0.0678077
R13743 VPWR VPWR.n201 0.0678077
R13744 VPWR VPWR.n213 0.0678077
R13745 VPWR VPWR.n225 0.0678077
R13746 VPWR VPWR.n237 0.0678077
R13747 VPWR VPWR.n249 0.0678077
R13748 VPWR VPWR.n261 0.0678077
R13749 VPWR VPWR.n273 0.0678077
R13750 VPWR.n286 VPWR 0.0678077
R13751 VPWR VPWR.n129 0.0678077
R13752 VPWR VPWR.n118 0.0678077
R13753 VPWR.n1732 VPWR 0.0678077
R13754 VPWR VPWR.n1720 0.0678077
R13755 VPWR VPWR.n1708 0.0678077
R13756 VPWR VPWR.n1697 0.0678077
R13757 VPWR.n1193 VPWR 0.0678077
R13758 VPWR VPWR.n1681 0.0678077
R13759 VPWR VPWR.n1670 0.0678077
R13760 VPWR.n1207 VPWR 0.0678077
R13761 VPWR VPWR.n1654 0.0678077
R13762 VPWR VPWR.n1643 0.0678077
R13763 VPWR.n1175 VPWR 0.0678077
R13764 VPWR VPWR.n1627 0.0678077
R13765 VPWR VPWR.n1616 0.0678077
R13766 VPWR.n1124 VPWR 0.0678077
R13767 VPWR VPWR.n1600 0.0678077
R13768 VPWR.n150 VPWR 0.063
R13769 VPWR.n162 VPWR 0.063
R13770 VPWR.n174 VPWR 0.063
R13771 VPWR.n186 VPWR 0.063
R13772 VPWR.n198 VPWR 0.063
R13773 VPWR.n210 VPWR 0.063
R13774 VPWR.n222 VPWR 0.063
R13775 VPWR.n234 VPWR 0.063
R13776 VPWR.n246 VPWR 0.063
R13777 VPWR.n258 VPWR 0.063
R13778 VPWR.n270 VPWR 0.063
R13779 VPWR.n101 VPWR 0.063
R13780 VPWR.n105 VPWR 0.063
R13781 VPWR.n138 VPWR 0.063
R13782 VPWR.n115 VPWR 0.063
R13783 VPWR.n126 VPWR 0.063
R13784 VPWR.n1065 VPWR 0.063
R13785 VPWR.n1717 VPWR 0.063
R13786 VPWR.n1070 VPWR 0.063
R13787 VPWR VPWR.n1704 0.063
R13788 VPWR VPWR.n1693 0.063
R13789 VPWR VPWR.n1081 0.063
R13790 VPWR VPWR.n1677 0.063
R13791 VPWR VPWR.n1666 0.063
R13792 VPWR VPWR.n1091 0.063
R13793 VPWR VPWR.n1650 0.063
R13794 VPWR VPWR.n1639 0.063
R13795 VPWR VPWR.n1101 0.063
R13796 VPWR VPWR.n1623 0.063
R13797 VPWR VPWR.n1612 0.063
R13798 VPWR VPWR.n1111 0.063
R13799 VPWR VPWR.n1120 0.063
R13800 VPWR.n1115 VPWR 0.0608448
R13801 VPWR.n107 VPWR 0.0608448
R13802 VPWR.n141 VPWR 0.0608448
R13803 VPWR.n153 VPWR 0.0608448
R13804 VPWR.n165 VPWR 0.0608448
R13805 VPWR.n177 VPWR 0.0608448
R13806 VPWR.n189 VPWR 0.0608448
R13807 VPWR.n201 VPWR 0.0608448
R13808 VPWR.n213 VPWR 0.0608448
R13809 VPWR.n225 VPWR 0.0608448
R13810 VPWR.n237 VPWR 0.0608448
R13811 VPWR.n249 VPWR 0.0608448
R13812 VPWR.n261 VPWR 0.0608448
R13813 VPWR.n273 VPWR 0.0608448
R13814 VPWR.n286 VPWR 0.0608448
R13815 VPWR.n129 VPWR 0.0608448
R13816 VPWR.n118 VPWR 0.0608448
R13817 VPWR.n1732 VPWR 0.0608448
R13818 VPWR.n1720 VPWR 0.0608448
R13819 VPWR.n1708 VPWR 0.0608448
R13820 VPWR.n1697 VPWR 0.0608448
R13821 VPWR.n1193 VPWR 0.0608448
R13822 VPWR.n1681 VPWR 0.0608448
R13823 VPWR.n1670 VPWR 0.0608448
R13824 VPWR.n1207 VPWR 0.0608448
R13825 VPWR.n1654 VPWR 0.0608448
R13826 VPWR.n1643 VPWR 0.0608448
R13827 VPWR.n1175 VPWR 0.0608448
R13828 VPWR.n1627 VPWR 0.0608448
R13829 VPWR.n1616 VPWR 0.0608448
R13830 VPWR.n1124 VPWR 0.0608448
R13831 VPWR.n1600 VPWR 0.0608448
R13832 VPWR VPWR.n13 0.0603958
R13833 VPWR VPWR.n12 0.0603958
R13834 VPWR VPWR.n1249 0.0603958
R13835 VPWR VPWR.n1248 0.0603958
R13836 VPWR VPWR.n1272 0.0603958
R13837 VPWR VPWR.n1271 0.0603958
R13838 VPWR VPWR.n1296 0.0603958
R13839 VPWR VPWR.n1295 0.0603958
R13840 VPWR.n1332 VPWR 0.0603958
R13841 VPWR VPWR.n1331 0.0603958
R13842 VPWR.n1327 VPWR 0.0603958
R13843 VPWR.n1318 VPWR 0.0603958
R13844 VPWR VPWR.n1317 0.0603958
R13845 VPWR.n1370 VPWR 0.0603958
R13846 VPWR VPWR.n1369 0.0603958
R13847 VPWR.n1364 VPWR 0.0603958
R13848 VPWR.n1409 VPWR 0.0603958
R13849 VPWR VPWR.n1408 0.0603958
R13850 VPWR.n1403 VPWR 0.0603958
R13851 VPWR.n1440 VPWR 0.0603958
R13852 VPWR VPWR.n2800 0.0603958
R13853 VPWR VPWR.n2799 0.0603958
R13854 VPWR VPWR.n2812 0.0603958
R13855 VPWR.n2791 VPWR 0.0603958
R13856 VPWR.n2792 VPWR 0.0603958
R13857 VPWR VPWR.n2796 0.0603958
R13858 VPWR.n2771 VPWR 0.0603958
R13859 VPWR.n2772 VPWR 0.0603958
R13860 VPWR VPWR.n2777 0.0603958
R13861 VPWR.n2752 VPWR 0.0603958
R13862 VPWR.n2753 VPWR 0.0603958
R13863 VPWR VPWR.n2757 0.0603958
R13864 VPWR.n2733 VPWR 0.0603958
R13865 VPWR.n2734 VPWR 0.0603958
R13866 VPWR VPWR.n2695 0.0603958
R13867 VPWR.n2696 VPWR 0.0603958
R13868 VPWR.n2697 VPWR 0.0603958
R13869 VPWR VPWR.n2658 0.0603958
R13870 VPWR.n2659 VPWR 0.0603958
R13871 VPWR.n2660 VPWR 0.0603958
R13872 VPWR.n2624 VPWR 0.0603958
R13873 VPWR.n2627 VPWR 0.0603958
R13874 VPWR.n1770 VPWR.n1769 0.0599512
R13875 VPWR.n1041 VPWR.n1040 0.0599512
R13876 VPWR.n1545 VPWR.n1544 0.0599512
R13877 VPWR.n1550 VPWR.n1549 0.0599512
R13878 VPWR.n1555 VPWR.n1554 0.0599512
R13879 VPWR.n1560 VPWR.n1559 0.0599512
R13880 VPWR.n1565 VPWR.n1564 0.0599512
R13881 VPWR.n1570 VPWR.n1569 0.0599512
R13882 VPWR.n1575 VPWR.n1574 0.0599512
R13883 VPWR.n1580 VPWR.n1579 0.0599512
R13884 VPWR.n1135 VPWR.n1134 0.0599512
R13885 VPWR.n1460 VPWR.n1459 0.0599512
R13886 VPWR.n1455 VPWR.n1454 0.0599512
R13887 VPWR.n1775 VPWR.n1774 0.0599512
R13888 VPWR.n1783 VPWR.n1782 0.0599512
R13889 VPWR.n1779 VPWR.n1778 0.0599512
R13890 VPWR.n1118 VPWR.n1117 0.0565345
R13891 VPWR.n1112 VPWR 0.0565345
R13892 VPWR.n144 VPWR.n143 0.0565345
R13893 VPWR.n146 VPWR 0.0565345
R13894 VPWR.n156 VPWR.n155 0.0565345
R13895 VPWR.n158 VPWR 0.0565345
R13896 VPWR.n168 VPWR.n167 0.0565345
R13897 VPWR.n170 VPWR 0.0565345
R13898 VPWR.n180 VPWR.n179 0.0565345
R13899 VPWR.n182 VPWR 0.0565345
R13900 VPWR.n192 VPWR.n191 0.0565345
R13901 VPWR.n194 VPWR 0.0565345
R13902 VPWR.n204 VPWR.n203 0.0565345
R13903 VPWR.n206 VPWR 0.0565345
R13904 VPWR.n216 VPWR.n215 0.0565345
R13905 VPWR.n218 VPWR 0.0565345
R13906 VPWR.n228 VPWR.n227 0.0565345
R13907 VPWR.n230 VPWR 0.0565345
R13908 VPWR.n240 VPWR.n239 0.0565345
R13909 VPWR.n242 VPWR 0.0565345
R13910 VPWR.n252 VPWR.n251 0.0565345
R13911 VPWR.n254 VPWR 0.0565345
R13912 VPWR.n264 VPWR.n263 0.0565345
R13913 VPWR.n266 VPWR 0.0565345
R13914 VPWR.n276 VPWR.n275 0.0565345
R13915 VPWR.n278 VPWR 0.0565345
R13916 VPWR.n285 VPWR.n283 0.0565345
R13917 VPWR.n103 VPWR 0.0565345
R13918 VPWR.n110 VPWR.n109 0.0565345
R13919 VPWR.n112 VPWR 0.0565345
R13920 VPWR.n132 VPWR.n131 0.0565345
R13921 VPWR.n134 VPWR 0.0565345
R13922 VPWR.n121 VPWR.n120 0.0565345
R13923 VPWR.n123 VPWR 0.0565345
R13924 VPWR.n1731 VPWR.n1729 0.0565345
R13925 VPWR.n1067 VPWR 0.0565345
R13926 VPWR.n1723 VPWR.n1722 0.0565345
R13927 VPWR.n1725 VPWR 0.0565345
R13928 VPWR.n1711 VPWR.n1710 0.0565345
R13929 VPWR.n1713 VPWR 0.0565345
R13930 VPWR.n1702 VPWR.n1699 0.0565345
R13931 VPWR.n1700 VPWR 0.0565345
R13932 VPWR.n1691 VPWR.n1077 0.0565345
R13933 VPWR.n1078 VPWR 0.0565345
R13934 VPWR.n1684 VPWR.n1683 0.0565345
R13935 VPWR.n1686 VPWR 0.0565345
R13936 VPWR.n1675 VPWR.n1672 0.0565345
R13937 VPWR.n1673 VPWR 0.0565345
R13938 VPWR.n1664 VPWR.n1087 0.0565345
R13939 VPWR.n1088 VPWR 0.0565345
R13940 VPWR.n1657 VPWR.n1656 0.0565345
R13941 VPWR.n1659 VPWR 0.0565345
R13942 VPWR.n1648 VPWR.n1645 0.0565345
R13943 VPWR.n1646 VPWR 0.0565345
R13944 VPWR.n1637 VPWR.n1097 0.0565345
R13945 VPWR.n1098 VPWR 0.0565345
R13946 VPWR.n1630 VPWR.n1629 0.0565345
R13947 VPWR.n1632 VPWR 0.0565345
R13948 VPWR.n1621 VPWR.n1618 0.0565345
R13949 VPWR.n1619 VPWR 0.0565345
R13950 VPWR.n1610 VPWR.n1107 0.0565345
R13951 VPWR.n1108 VPWR 0.0565345
R13952 VPWR.n1603 VPWR.n1602 0.0565345
R13953 VPWR.n1605 VPWR 0.0565345
R13954 VPWR.n1769 VPWR 0.0469286
R13955 VPWR.n1040 VPWR 0.0469286
R13956 VPWR.n1544 VPWR 0.0469286
R13957 VPWR.n1549 VPWR 0.0469286
R13958 VPWR.n1554 VPWR 0.0469286
R13959 VPWR.n1559 VPWR 0.0469286
R13960 VPWR.n1564 VPWR 0.0469286
R13961 VPWR.n1569 VPWR 0.0469286
R13962 VPWR.n1574 VPWR 0.0469286
R13963 VPWR.n1579 VPWR 0.0469286
R13964 VPWR.n1134 VPWR 0.0469286
R13965 VPWR.n1459 VPWR 0.0469286
R13966 VPWR.n1454 VPWR 0.0469286
R13967 VPWR.n1774 VPWR 0.0469286
R13968 VPWR.n1782 VPWR 0.0469286
R13969 VPWR.n1778 VPWR 0.0469286
R13970 VPWR.n1769 VPWR 0.0401341
R13971 VPWR.n1040 VPWR 0.0401341
R13972 VPWR.n1544 VPWR 0.0401341
R13973 VPWR.n1549 VPWR 0.0401341
R13974 VPWR.n1554 VPWR 0.0401341
R13975 VPWR.n1559 VPWR 0.0401341
R13976 VPWR.n1564 VPWR 0.0401341
R13977 VPWR.n1569 VPWR 0.0401341
R13978 VPWR.n1574 VPWR 0.0401341
R13979 VPWR.n1579 VPWR 0.0401341
R13980 VPWR.n1134 VPWR 0.0401341
R13981 VPWR.n1459 VPWR 0.0401341
R13982 VPWR.n1454 VPWR 0.0401341
R13983 VPWR.n1774 VPWR 0.0401341
R13984 VPWR.n1782 VPWR 0.0401341
R13985 VPWR.n1778 VPWR 0.0401341
R13986 VPWR.n13 VPWR 0.0382604
R13987 VPWR.n1249 VPWR 0.0382604
R13988 VPWR.n1272 VPWR 0.0382604
R13989 VPWR.n1296 VPWR 0.0382604
R13990 VPWR.n1331 VPWR 0.0382604
R13991 VPWR.n1369 VPWR 0.0382604
R13992 VPWR.n1408 VPWR 0.0382604
R13993 VPWR.n1445 VPWR 0.0382604
R13994 VPWR.n20 VPWR 0.0375125
R13995 VPWR.n20 VPWR 0.0373589
R13996 VPWR.n1118 VPWR.n1109 0.0349828
R13997 VPWR.n147 VPWR.n144 0.0349828
R13998 VPWR.n159 VPWR.n156 0.0349828
R13999 VPWR.n171 VPWR.n168 0.0349828
R14000 VPWR.n183 VPWR.n180 0.0349828
R14001 VPWR.n195 VPWR.n192 0.0349828
R14002 VPWR.n207 VPWR.n204 0.0349828
R14003 VPWR.n219 VPWR.n216 0.0349828
R14004 VPWR.n231 VPWR.n228 0.0349828
R14005 VPWR.n243 VPWR.n240 0.0349828
R14006 VPWR.n255 VPWR.n252 0.0349828
R14007 VPWR.n267 VPWR.n264 0.0349828
R14008 VPWR.n279 VPWR.n276 0.0349828
R14009 VPWR.n283 VPWR.n282 0.0349828
R14010 VPWR.n113 VPWR.n110 0.0349828
R14011 VPWR.n135 VPWR.n132 0.0349828
R14012 VPWR.n124 VPWR.n121 0.0349828
R14013 VPWR.n1729 VPWR.n1728 0.0349828
R14014 VPWR.n1726 VPWR.n1723 0.0349828
R14015 VPWR.n1714 VPWR.n1711 0.0349828
R14016 VPWR.n1702 VPWR.n1701 0.0349828
R14017 VPWR.n1691 VPWR.n1690 0.0349828
R14018 VPWR.n1687 VPWR.n1684 0.0349828
R14019 VPWR.n1675 VPWR.n1674 0.0349828
R14020 VPWR.n1664 VPWR.n1663 0.0349828
R14021 VPWR.n1660 VPWR.n1657 0.0349828
R14022 VPWR.n1648 VPWR.n1647 0.0349828
R14023 VPWR.n1637 VPWR.n1636 0.0349828
R14024 VPWR.n1633 VPWR.n1630 0.0349828
R14025 VPWR.n1621 VPWR.n1620 0.0349828
R14026 VPWR.n1610 VPWR.n1609 0.0349828
R14027 VPWR.n1606 VPWR.n1603 0.0349828
R14028 VPWR.n2504 VPWR.n2503 0.0340366
R14029 VPWR.n2570 VPWR.n2569 0.0340366
R14030 VPWR.n2510 VPWR.n2509 0.0340366
R14031 VPWR.n2552 VPWR.n2551 0.0340366
R14032 VPWR.n2546 VPWR.n2545 0.0340366
R14033 VPWR.n2534 VPWR.n2533 0.0340366
R14034 VPWR.n2528 VPWR.n2527 0.0340366
R14035 VPWR.n1223 VPWR.n1222 0.0340366
R14036 VPWR.n2522 VPWR.n2521 0.0340366
R14037 VPWR.n1486 VPWR.n1102 0.0340366
R14038 VPWR.n1174 VPWR.n1094 0.0340366
R14039 VPWR.n2540 VPWR.n2539 0.0340366
R14040 VPWR.n1165 VPWR.n1092 0.0340366
R14041 VPWR.n1211 VPWR.n1164 0.0340366
R14042 VPWR.n2516 VPWR.n2515 0.0340366
R14043 VPWR.n1129 VPWR.n1104 0.0340366
R14044 VPWR.n1155 VPWR.n1084 0.0340366
R14045 VPWR.n2558 VPWR.n2557 0.0340366
R14046 VPWR.n1144 VPWR.n1082 0.0340366
R14047 VPWR.n1591 VPWR.n1590 0.0340366
R14048 VPWR.n2564 VPWR.n2563 0.0340366
R14049 VPWR.n1197 VPWR.n1154 0.0340366
R14050 VPWR.n1074 VPWR.n1073 0.0340366
R14051 VPWR.n1743 VPWR.n1742 0.0340366
R14052 VPWR.n1071 VPWR.n1054 0.0340366
R14053 VPWR.n2576 VPWR.n2575 0.0340366
R14054 VPWR.n2582 VPWR.n2581 0.0340366
R14055 VPWR.n2593 VPWR.n2592 0.0340366
R14056 VPWR.n2588 VPWR.n2587 0.0340366
R14057 VPWR.n1737 VPWR.n1736 0.0340366
R14058 VPWR.n1063 VPWR.n1060 0.0340366
R14059 VPWR.n1596 VPWR.n1121 0.0340366
R14060 VPWR.n2628 VPWR.n2598 0.0320292
R14061 VPWR.n2800 VPWR 0.03175
R14062 VPWR VPWR.n2791 0.03175
R14063 VPWR VPWR.n2771 0.03175
R14064 VPWR VPWR.n2752 0.03175
R14065 VPWR VPWR.n2733 0.03175
R14066 VPWR VPWR.n2696 0.03175
R14067 VPWR VPWR.n2659 0.03175
R14068 VPWR VPWR.n2627 0.03175
R14069 VPWR.n2598 VPWR.n2597 0.0240975
R14070 VPWR.n2597 VPWR.n20 0.0240975
R14071 VPWR.n2814 VPWR 0.024
R14072 VPWR.n14 VPWR 0.0239375
R14073 VPWR.n12 VPWR 0.0239375
R14074 VPWR.n1250 VPWR 0.0239375
R14075 VPWR.n1248 VPWR 0.0239375
R14076 VPWR.n1271 VPWR 0.0239375
R14077 VPWR.n1295 VPWR 0.0239375
R14078 VPWR.n2753 VPWR 0.0239375
R14079 VPWR.n2503 VPWR 0.0233659
R14080 VPWR.n1466 VPWR 0.0233659
R14081 VPWR.n352 VPWR 0.0233659
R14082 VPWR.n2570 VPWR 0.0233659
R14083 VPWR.n1533 VPWR 0.0233659
R14084 VPWR.n347 VPWR 0.0233659
R14085 VPWR.n2510 VPWR 0.0233659
R14086 VPWR.n964 VPWR 0.0233659
R14087 VPWR.n2479 VPWR 0.0233659
R14088 VPWR.n2474 VPWR 0.0233659
R14089 VPWR.n319 VPWR 0.0233659
R14090 VPWR.n2551 VPWR 0.0233659
R14091 VPWR.n972 VPWR 0.0233659
R14092 VPWR.n2444 VPWR 0.0233659
R14093 VPWR.n323 VPWR 0.0233659
R14094 VPWR.n2546 VPWR 0.0233659
R14095 VPWR.n1891 VPWR 0.0233659
R14096 VPWR.n1886 VPWR 0.0233659
R14097 VPWR.n1881 VPWR 0.0233659
R14098 VPWR.n388 VPWR 0.0233659
R14099 VPWR.n392 VPWR 0.0233659
R14100 VPWR.n396 VPWR 0.0233659
R14101 VPWR.n2454 VPWR 0.0233659
R14102 VPWR.n331 VPWR 0.0233659
R14103 VPWR.n2534 VPWR 0.0233659
R14104 VPWR.n1876 VPWR 0.0233659
R14105 VPWR.n404 VPWR 0.0233659
R14106 VPWR.n2459 VPWR 0.0233659
R14107 VPWR.n335 VPWR 0.0233659
R14108 VPWR.n2527 VPWR 0.0233659
R14109 VPWR.n2307 VPWR 0.0233659
R14110 VPWR.n2312 VPWR 0.0233659
R14111 VPWR.n2317 VPWR 0.0233659
R14112 VPWR.n2322 VPWR 0.0233659
R14113 VPWR.n2332 VPWR 0.0233659
R14114 VPWR.n2337 VPWR 0.0233659
R14115 VPWR.n2342 VPWR 0.0233659
R14116 VPWR.n2347 VPWR 0.0233659
R14117 VPWR.n2352 VPWR 0.0233659
R14118 VPWR.n2357 VPWR 0.0233659
R14119 VPWR.n2362 VPWR 0.0233659
R14120 VPWR.n2367 VPWR 0.0233659
R14121 VPWR.n2372 VPWR 0.0233659
R14122 VPWR.n2377 VPWR 0.0233659
R14123 VPWR.n2381 VPWR 0.0233659
R14124 VPWR.n2327 VPWR 0.0233659
R14125 VPWR.n544 VPWR 0.0233659
R14126 VPWR.n539 VPWR 0.0233659
R14127 VPWR.n535 VPWR 0.0233659
R14128 VPWR.n531 VPWR 0.0233659
R14129 VPWR.n523 VPWR 0.0233659
R14130 VPWR.n519 VPWR 0.0233659
R14131 VPWR.n515 VPWR 0.0233659
R14132 VPWR.n511 VPWR 0.0233659
R14133 VPWR.n507 VPWR 0.0233659
R14134 VPWR.n503 VPWR 0.0233659
R14135 VPWR.n499 VPWR 0.0233659
R14136 VPWR.n495 VPWR 0.0233659
R14137 VPWR.n491 VPWR 0.0233659
R14138 VPWR.n487 VPWR 0.0233659
R14139 VPWR.n484 VPWR 0.0233659
R14140 VPWR.n527 VPWR 0.0233659
R14141 VPWR.n2283 VPWR 0.0233659
R14142 VPWR.n2278 VPWR 0.0233659
R14143 VPWR.n2273 VPWR 0.0233659
R14144 VPWR.n2268 VPWR 0.0233659
R14145 VPWR.n2258 VPWR 0.0233659
R14146 VPWR.n2253 VPWR 0.0233659
R14147 VPWR.n2248 VPWR 0.0233659
R14148 VPWR.n2243 VPWR 0.0233659
R14149 VPWR.n2238 VPWR 0.0233659
R14150 VPWR.n2233 VPWR 0.0233659
R14151 VPWR.n2228 VPWR 0.0233659
R14152 VPWR.n2223 VPWR 0.0233659
R14153 VPWR.n2218 VPWR 0.0233659
R14154 VPWR.n2213 VPWR 0.0233659
R14155 VPWR.n2209 VPWR 0.0233659
R14156 VPWR.n2263 VPWR 0.0233659
R14157 VPWR.n580 VPWR 0.0233659
R14158 VPWR.n584 VPWR 0.0233659
R14159 VPWR.n588 VPWR 0.0233659
R14160 VPWR.n592 VPWR 0.0233659
R14161 VPWR.n600 VPWR 0.0233659
R14162 VPWR.n604 VPWR 0.0233659
R14163 VPWR.n608 VPWR 0.0233659
R14164 VPWR.n612 VPWR 0.0233659
R14165 VPWR.n616 VPWR 0.0233659
R14166 VPWR.n620 VPWR 0.0233659
R14167 VPWR.n624 VPWR 0.0233659
R14168 VPWR.n628 VPWR 0.0233659
R14169 VPWR.n632 VPWR 0.0233659
R14170 VPWR.n636 VPWR 0.0233659
R14171 VPWR.n640 VPWR 0.0233659
R14172 VPWR.n596 VPWR 0.0233659
R14173 VPWR.n2111 VPWR 0.0233659
R14174 VPWR.n2116 VPWR 0.0233659
R14175 VPWR.n2121 VPWR 0.0233659
R14176 VPWR.n2126 VPWR 0.0233659
R14177 VPWR.n2136 VPWR 0.0233659
R14178 VPWR.n2141 VPWR 0.0233659
R14179 VPWR.n2146 VPWR 0.0233659
R14180 VPWR.n2151 VPWR 0.0233659
R14181 VPWR.n2156 VPWR 0.0233659
R14182 VPWR.n2161 VPWR 0.0233659
R14183 VPWR.n2166 VPWR 0.0233659
R14184 VPWR.n2171 VPWR 0.0233659
R14185 VPWR.n2176 VPWR 0.0233659
R14186 VPWR.n2181 VPWR 0.0233659
R14187 VPWR.n2185 VPWR 0.0233659
R14188 VPWR.n2131 VPWR 0.0233659
R14189 VPWR.n736 VPWR 0.0233659
R14190 VPWR.n731 VPWR 0.0233659
R14191 VPWR.n727 VPWR 0.0233659
R14192 VPWR.n723 VPWR 0.0233659
R14193 VPWR.n715 VPWR 0.0233659
R14194 VPWR.n711 VPWR 0.0233659
R14195 VPWR.n707 VPWR 0.0233659
R14196 VPWR.n703 VPWR 0.0233659
R14197 VPWR.n699 VPWR 0.0233659
R14198 VPWR.n695 VPWR 0.0233659
R14199 VPWR.n691 VPWR 0.0233659
R14200 VPWR.n687 VPWR 0.0233659
R14201 VPWR.n683 VPWR 0.0233659
R14202 VPWR.n679 VPWR 0.0233659
R14203 VPWR.n676 VPWR 0.0233659
R14204 VPWR.n719 VPWR 0.0233659
R14205 VPWR.n2087 VPWR 0.0233659
R14206 VPWR.n2082 VPWR 0.0233659
R14207 VPWR.n2077 VPWR 0.0233659
R14208 VPWR.n2072 VPWR 0.0233659
R14209 VPWR.n2062 VPWR 0.0233659
R14210 VPWR.n2057 VPWR 0.0233659
R14211 VPWR.n2052 VPWR 0.0233659
R14212 VPWR.n2047 VPWR 0.0233659
R14213 VPWR.n2042 VPWR 0.0233659
R14214 VPWR.n2037 VPWR 0.0233659
R14215 VPWR.n2032 VPWR 0.0233659
R14216 VPWR.n2027 VPWR 0.0233659
R14217 VPWR.n2022 VPWR 0.0233659
R14218 VPWR.n2017 VPWR 0.0233659
R14219 VPWR.n2013 VPWR 0.0233659
R14220 VPWR.n2067 VPWR 0.0233659
R14221 VPWR.n772 VPWR 0.0233659
R14222 VPWR.n776 VPWR 0.0233659
R14223 VPWR.n780 VPWR 0.0233659
R14224 VPWR.n784 VPWR 0.0233659
R14225 VPWR.n792 VPWR 0.0233659
R14226 VPWR.n796 VPWR 0.0233659
R14227 VPWR.n800 VPWR 0.0233659
R14228 VPWR.n804 VPWR 0.0233659
R14229 VPWR.n808 VPWR 0.0233659
R14230 VPWR.n812 VPWR 0.0233659
R14231 VPWR.n816 VPWR 0.0233659
R14232 VPWR.n820 VPWR 0.0233659
R14233 VPWR.n824 VPWR 0.0233659
R14234 VPWR.n828 VPWR 0.0233659
R14235 VPWR.n832 VPWR 0.0233659
R14236 VPWR.n788 VPWR 0.0233659
R14237 VPWR.n1915 VPWR 0.0233659
R14238 VPWR.n1920 VPWR 0.0233659
R14239 VPWR.n1925 VPWR 0.0233659
R14240 VPWR.n1930 VPWR 0.0233659
R14241 VPWR.n1940 VPWR 0.0233659
R14242 VPWR.n1945 VPWR 0.0233659
R14243 VPWR.n1950 VPWR 0.0233659
R14244 VPWR.n1955 VPWR 0.0233659
R14245 VPWR.n1960 VPWR 0.0233659
R14246 VPWR.n1965 VPWR 0.0233659
R14247 VPWR.n1970 VPWR 0.0233659
R14248 VPWR.n1975 VPWR 0.0233659
R14249 VPWR.n1980 VPWR 0.0233659
R14250 VPWR.n1985 VPWR 0.0233659
R14251 VPWR.n1989 VPWR 0.0233659
R14252 VPWR.n1935 VPWR 0.0233659
R14253 VPWR.n928 VPWR 0.0233659
R14254 VPWR.n923 VPWR 0.0233659
R14255 VPWR.n919 VPWR 0.0233659
R14256 VPWR.n915 VPWR 0.0233659
R14257 VPWR.n907 VPWR 0.0233659
R14258 VPWR.n903 VPWR 0.0233659
R14259 VPWR.n899 VPWR 0.0233659
R14260 VPWR.n895 VPWR 0.0233659
R14261 VPWR.n891 VPWR 0.0233659
R14262 VPWR.n887 VPWR 0.0233659
R14263 VPWR.n883 VPWR 0.0233659
R14264 VPWR.n879 VPWR 0.0233659
R14265 VPWR.n875 VPWR 0.0233659
R14266 VPWR.n871 VPWR 0.0233659
R14267 VPWR.n868 VPWR 0.0233659
R14268 VPWR.n911 VPWR 0.0233659
R14269 VPWR.n1871 VPWR 0.0233659
R14270 VPWR.n980 VPWR 0.0233659
R14271 VPWR.n1495 VPWR 0.0233659
R14272 VPWR.n1223 VPWR 0.0233659
R14273 VPWR.n400 VPWR 0.0233659
R14274 VPWR.n2464 VPWR 0.0233659
R14275 VPWR.n339 VPWR 0.0233659
R14276 VPWR.n2522 VPWR 0.0233659
R14277 VPWR.n976 VPWR 0.0233659
R14278 VPWR.n1490 VPWR 0.0233659
R14279 VPWR.n1486 VPWR 0.0233659
R14280 VPWR.n1866 VPWR 0.0233659
R14281 VPWR.n984 VPWR 0.0233659
R14282 VPWR.n1504 VPWR 0.0233659
R14283 VPWR.n1174 VPWR 0.0233659
R14284 VPWR.n408 VPWR 0.0233659
R14285 VPWR.n416 VPWR 0.0233659
R14286 VPWR.n420 VPWR 0.0233659
R14287 VPWR.n424 VPWR 0.0233659
R14288 VPWR.n428 VPWR 0.0233659
R14289 VPWR.n432 VPWR 0.0233659
R14290 VPWR.n436 VPWR 0.0233659
R14291 VPWR.n440 VPWR 0.0233659
R14292 VPWR.n444 VPWR 0.0233659
R14293 VPWR.n448 VPWR 0.0233659
R14294 VPWR.n412 VPWR 0.0233659
R14295 VPWR.n2449 VPWR 0.0233659
R14296 VPWR.n327 VPWR 0.0233659
R14297 VPWR.n2539 VPWR 0.0233659
R14298 VPWR.n988 VPWR 0.0233659
R14299 VPWR.n1509 VPWR 0.0233659
R14300 VPWR.n1165 VPWR 0.0233659
R14301 VPWR.n1861 VPWR 0.0233659
R14302 VPWR.n1851 VPWR 0.0233659
R14303 VPWR.n1846 VPWR 0.0233659
R14304 VPWR.n1841 VPWR 0.0233659
R14305 VPWR.n1836 VPWR 0.0233659
R14306 VPWR.n1831 VPWR 0.0233659
R14307 VPWR.n1826 VPWR 0.0233659
R14308 VPWR.n1821 VPWR 0.0233659
R14309 VPWR.n1817 VPWR 0.0233659
R14310 VPWR.n1856 VPWR 0.0233659
R14311 VPWR.n992 VPWR 0.0233659
R14312 VPWR.n1518 VPWR 0.0233659
R14313 VPWR.n1164 VPWR 0.0233659
R14314 VPWR.n2469 VPWR 0.0233659
R14315 VPWR.n343 VPWR 0.0233659
R14316 VPWR.n2515 VPWR 0.0233659
R14317 VPWR.n1130 VPWR 0.0233659
R14318 VPWR.n1129 VPWR 0.0233659
R14319 VPWR.n996 VPWR 0.0233659
R14320 VPWR.n1523 VPWR 0.0233659
R14321 VPWR.n1155 VPWR 0.0233659
R14322 VPWR.n2439 VPWR 0.0233659
R14323 VPWR.n2429 VPWR 0.0233659
R14324 VPWR.n2424 VPWR 0.0233659
R14325 VPWR.n2419 VPWR 0.0233659
R14326 VPWR.n2414 VPWR 0.0233659
R14327 VPWR.n2409 VPWR 0.0233659
R14328 VPWR.n2405 VPWR 0.0233659
R14329 VPWR.n2434 VPWR 0.0233659
R14330 VPWR.n315 VPWR 0.0233659
R14331 VPWR.n2558 VPWR 0.0233659
R14332 VPWR.n1538 VPWR 0.0233659
R14333 VPWR.n1144 VPWR 0.0233659
R14334 VPWR.n1000 VPWR 0.0233659
R14335 VPWR.n1004 VPWR 0.0233659
R14336 VPWR.n1008 VPWR 0.0233659
R14337 VPWR.n1012 VPWR 0.0233659
R14338 VPWR.n1016 VPWR 0.0233659
R14339 VPWR.n1020 VPWR 0.0233659
R14340 VPWR.n1024 VPWR 0.0233659
R14341 VPWR.n968 VPWR 0.0233659
R14342 VPWR.n1473 VPWR 0.0233659
R14343 VPWR.n1590 VPWR 0.0233659
R14344 VPWR.n311 VPWR 0.0233659
R14345 VPWR.n2563 VPWR 0.0233659
R14346 VPWR.n1154 VPWR 0.0233659
R14347 VPWR.n1763 VPWR 0.0233659
R14348 VPWR.n1073 VPWR 0.0233659
R14349 VPWR.n307 VPWR 0.0233659
R14350 VPWR.n303 VPWR 0.0233659
R14351 VPWR.n295 VPWR 0.0233659
R14352 VPWR.n292 VPWR 0.0233659
R14353 VPWR.n299 VPWR 0.0233659
R14354 VPWR.n1743 VPWR 0.0233659
R14355 VPWR.n1751 VPWR 0.0233659
R14356 VPWR.n1789 VPWR 0.0233659
R14357 VPWR.n1793 VPWR 0.0233659
R14358 VPWR.n1758 VPWR 0.0233659
R14359 VPWR.n1054 VPWR 0.0233659
R14360 VPWR.n2575 VPWR 0.0233659
R14361 VPWR.n2582 VPWR 0.0233659
R14362 VPWR.n2593 VPWR 0.0233659
R14363 VPWR.n2587 VPWR 0.0233659
R14364 VPWR.n1736 VPWR 0.0233659
R14365 VPWR.n1060 VPWR 0.0233659
R14366 VPWR.n1121 VPWR 0.0233659
R14367 VPWR.n1336 VPWR 0.0226354
R14368 VPWR.n1327 VPWR 0.0226354
R14369 VPWR.n1413 VPWR 0.0226354
R14370 VPWR.n2772 VPWR 0.0226354
R14371 VPWR VPWR.n2732 0.0226354
R14372 VPWR VPWR.n2702 0.0226354
R14373 VPWR VPWR.n2664 0.0226354
R14374 VPWR VPWR.n64 0.0220517
R14375 VPWR VPWR.n67 0.0220517
R14376 VPWR VPWR.n70 0.0220517
R14377 VPWR VPWR.n73 0.0220517
R14378 VPWR VPWR.n76 0.0220517
R14379 VPWR VPWR.n79 0.0220517
R14380 VPWR VPWR.n82 0.0220517
R14381 VPWR VPWR.n85 0.0220517
R14382 VPWR VPWR.n88 0.0220517
R14383 VPWR VPWR.n91 0.0220517
R14384 VPWR VPWR.n94 0.0220517
R14385 VPWR VPWR.n97 0.0220517
R14386 VPWR.n289 VPWR 0.0220517
R14387 VPWR VPWR.n61 0.0220517
R14388 VPWR VPWR.n58 0.0220517
R14389 VPWR.n1735 VPWR 0.0220517
R14390 VPWR VPWR.n1057 0.0220517
R14391 VPWR.n1705 VPWR 0.0220517
R14392 VPWR.n1694 VPWR 0.0220517
R14393 VPWR.n1196 VPWR 0.0220517
R14394 VPWR.n1678 VPWR 0.0220517
R14395 VPWR.n1667 VPWR 0.0220517
R14396 VPWR.n1210 VPWR 0.0220517
R14397 VPWR.n1651 VPWR 0.0220517
R14398 VPWR.n1640 VPWR 0.0220517
R14399 VPWR.n1178 VPWR 0.0220517
R14400 VPWR.n1624 VPWR 0.0220517
R14401 VPWR.n1613 VPWR 0.0220517
R14402 VPWR.n1127 VPWR 0.0220517
R14403 VPWR.n1597 VPWR 0.0220517
R14404 VPWR.n1273 VPWR 0.0213333
R14405 VPWR.n1297 VPWR 0.0213333
R14406 VPWR.n1311 VPWR 0.0213333
R14407 VPWR.n1375 VPWR 0.0213333
R14408 VPWR.n1347 VPWR 0.0213333
R14409 VPWR.n1386 VPWR 0.0213333
R14410 VPWR.n1423 VPWR 0.0213333
R14411 VPWR.n2806 VPWR 0.0213333
R14412 VPWR.n2799 VPWR 0.0213333
R14413 VPWR VPWR.n2790 0.0213333
R14414 VPWR.n2792 VPWR 0.0213333
R14415 VPWR VPWR.n2770 0.0213333
R14416 VPWR VPWR.n2751 0.0213333
R14417 VPWR VPWR.n2738 0.0213333
R14418 VPWR.n2500 VPWR 0.0196917
R14419 VPWR.n24 VPWR 0.0143889
R14420 VPWR VPWR.n19 0.0099
R14421 VPWR VPWR.n1604 0.00397222
R14422 VPWR VPWR.n1105 0.00397222
R14423 VPWR VPWR.n1103 0.00397222
R14424 VPWR VPWR.n1631 0.00397222
R14425 VPWR VPWR.n1095 0.00397222
R14426 VPWR VPWR.n1093 0.00397222
R14427 VPWR VPWR.n1658 0.00397222
R14428 VPWR VPWR.n1085 0.00397222
R14429 VPWR VPWR.n1083 0.00397222
R14430 VPWR VPWR.n1685 0.00397222
R14431 VPWR VPWR.n1075 0.00397222
R14432 VPWR VPWR.n1072 0.00397222
R14433 VPWR VPWR.n1712 0.00397222
R14434 VPWR VPWR.n1724 0.00397222
R14435 VPWR.n1113 VPWR 0.00397222
R14436 VPWR VPWR.n1066 0.00397222
R14437 VPWR VPWR.n122 0.00397222
R14438 VPWR VPWR.n111 0.00397222
R14439 VPWR VPWR.n102 0.00397222
R14440 VPWR VPWR.n277 0.00397222
R14441 VPWR VPWR.n265 0.00397222
R14442 VPWR VPWR.n253 0.00397222
R14443 VPWR VPWR.n241 0.00397222
R14444 VPWR VPWR.n229 0.00397222
R14445 VPWR VPWR.n217 0.00397222
R14446 VPWR VPWR.n205 0.00397222
R14447 VPWR VPWR.n193 0.00397222
R14448 VPWR VPWR.n181 0.00397222
R14449 VPWR VPWR.n169 0.00397222
R14450 VPWR VPWR.n157 0.00397222
R14451 VPWR VPWR.n145 0.00397222
R14452 VPWR VPWR.n133 0.00397222
R14453 VPWR.n1462 VPWR.n1461 0.00351282
R14454 VPWR.n1457 VPWR.n1136 0.00351282
R14455 VPWR.n1582 VPWR.n1581 0.00351282
R14456 VPWR.n1577 VPWR.n1576 0.00351282
R14457 VPWR.n1572 VPWR.n1571 0.00351282
R14458 VPWR.n1567 VPWR.n1566 0.00351282
R14459 VPWR.n1562 VPWR.n1561 0.00351282
R14460 VPWR.n1557 VPWR.n1556 0.00351282
R14461 VPWR.n1552 VPWR.n1551 0.00351282
R14462 VPWR.n1547 VPWR.n1546 0.00351282
R14463 VPWR.n1542 VPWR.n1042 0.00351282
R14464 VPWR.n1785 VPWR.n1784 0.00351282
R14465 VPWR.n1776 VPWR.n1772 0.00351282
R14466 VPWR.n1771 VPWR.n1767 0.00351282
R14467 VPWR.n141 VPWR.n140 0.00265517
R14468 VPWR.n153 VPWR.n152 0.00265517
R14469 VPWR.n165 VPWR.n164 0.00265517
R14470 VPWR.n177 VPWR.n176 0.00265517
R14471 VPWR.n189 VPWR.n188 0.00265517
R14472 VPWR.n201 VPWR.n200 0.00265517
R14473 VPWR.n213 VPWR.n212 0.00265517
R14474 VPWR.n225 VPWR.n224 0.00265517
R14475 VPWR.n237 VPWR.n236 0.00265517
R14476 VPWR.n249 VPWR.n248 0.00265517
R14477 VPWR.n261 VPWR.n260 0.00265517
R14478 VPWR.n273 VPWR.n272 0.00265517
R14479 VPWR.n288 VPWR.n286 0.00265517
R14480 VPWR.n129 VPWR.n128 0.00265517
R14481 VPWR.n118 VPWR.n117 0.00265517
R14482 VPWR.n1734 VPWR.n1732 0.00265517
R14483 VPWR.n1720 VPWR.n1719 0.00265517
R14484 VPWR.n1708 VPWR.n1707 0.00265517
R14485 VPWR.n1697 VPWR.n1696 0.00265517
R14486 VPWR.n1195 VPWR.n1193 0.00265517
R14487 VPWR.n1681 VPWR.n1680 0.00265517
R14488 VPWR.n1670 VPWR.n1669 0.00265517
R14489 VPWR.n1209 VPWR.n1207 0.00265517
R14490 VPWR.n1654 VPWR.n1653 0.00265517
R14491 VPWR.n1643 VPWR.n1642 0.00265517
R14492 VPWR.n1177 VPWR.n1175 0.00265517
R14493 VPWR.n1627 VPWR.n1626 0.00265517
R14494 VPWR.n1616 VPWR.n1615 0.00265517
R14495 VPWR.n1126 VPWR.n1124 0.00265517
R14496 VPWR.n1600 VPWR.n1599 0.00265517
R14497 Iout.n1020 Iout.t174 239.927
R14498 Iout.n509 Iout.t142 239.927
R14499 Iout.n513 Iout.t23 239.927
R14500 Iout.n507 Iout.t159 239.927
R14501 Iout.n504 Iout.t127 239.927
R14502 Iout.n500 Iout.t148 239.927
R14503 Iout.n192 Iout.t167 239.927
R14504 Iout.n195 Iout.t197 239.927
R14505 Iout.n199 Iout.t233 239.927
R14506 Iout.n202 Iout.t18 239.927
R14507 Iout.n206 Iout.t193 239.927
R14508 Iout.n210 Iout.t89 239.927
R14509 Iout.n214 Iout.t78 239.927
R14510 Iout.n218 Iout.t161 239.927
R14511 Iout.n222 Iout.t181 239.927
R14512 Iout.n226 Iout.t48 239.927
R14513 Iout.n232 Iout.t133 239.927
R14514 Iout.n235 Iout.t126 239.927
R14515 Iout.n238 Iout.t3 239.927
R14516 Iout.n241 Iout.t2 239.927
R14517 Iout.n244 Iout.t255 239.927
R14518 Iout.n247 Iout.t8 239.927
R14519 Iout.n250 Iout.t245 239.927
R14520 Iout.n255 Iout.t21 239.927
R14521 Iout.n252 Iout.t212 239.927
R14522 Iout.n489 Iout.t170 239.927
R14523 Iout.n494 Iout.t188 239.927
R14524 Iout.n491 Iout.t135 239.927
R14525 Iout.n519 Iout.t139 239.927
R14526 Iout.n149 Iout.t7 239.927
R14527 Iout.n146 Iout.t125 239.927
R14528 Iout.n1010 Iout.t106 239.927
R14529 Iout.n1007 Iout.t16 239.927
R14530 Iout.n140 Iout.t185 239.927
R14531 Iout.n143 Iout.t0 239.927
R14532 Iout.n525 Iout.t246 239.927
R14533 Iout.n480 Iout.t171 239.927
R14534 Iout.n483 Iout.t195 239.927
R14535 Iout.n478 Iout.t17 239.927
R14536 Iout.n259 Iout.t227 239.927
R14537 Iout.n186 Iout.t29 239.927
R14538 Iout.n271 Iout.t81 239.927
R14539 Iout.n180 Iout.t13 239.927
R14540 Iout.n283 Iout.t198 239.927
R14541 Iout.n174 Iout.t248 239.927
R14542 Iout.n168 Iout.t189 239.927
R14543 Iout.n301 Iout.t67 239.927
R14544 Iout.n289 Iout.t149 239.927
R14545 Iout.n177 Iout.t12 239.927
R14546 Iout.n277 Iout.t247 239.927
R14547 Iout.n183 Iout.t230 239.927
R14548 Iout.n265 Iout.t229 239.927
R14549 Iout.n189 Iout.t118 239.927
R14550 Iout.n472 Iout.t43 239.927
R14551 Iout.n469 Iout.t178 239.927
R14552 Iout.n156 Iout.t40 239.927
R14553 Iout.n531 Iout.t22 239.927
R14554 Iout.n534 Iout.t163 239.927
R14555 Iout.n536 Iout.t80 239.927
R14556 Iout.n133 Iout.t84 239.927
R14557 Iout.n136 Iout.t214 239.927
R14558 Iout.n542 Iout.t28 239.927
R14559 Iout.n460 Iout.t108 239.927
R14560 Iout.n463 Iout.t216 239.927
R14561 Iout.n458 Iout.t191 239.927
R14562 Iout.n305 Iout.t208 239.927
R14563 Iout.n308 Iout.t218 239.927
R14564 Iout.n311 Iout.t244 239.927
R14565 Iout.n314 Iout.t199 239.927
R14566 Iout.n317 Iout.t145 239.927
R14567 Iout.n320 Iout.t113 239.927
R14568 Iout.n392 Iout.t226 239.927
R14569 Iout.n378 Iout.t54 239.927
R14570 Iout.n376 Iout.t157 239.927
R14571 Iout.n394 Iout.t46 239.927
R14572 Iout.n408 Iout.t228 239.927
R14573 Iout.n410 Iout.t169 239.927
R14574 Iout.n424 Iout.t88 239.927
R14575 Iout.n426 Iout.t162 239.927
R14576 Iout.n447 Iout.t249 239.927
R14577 Iout.n452 Iout.t37 239.927
R14578 Iout.n449 Iout.t158 239.927
R14579 Iout.n548 Iout.t72 239.927
R14580 Iout.n130 Iout.t225 239.927
R14581 Iout.n559 Iout.t196 239.927
R14582 Iout.n557 Iout.t116 239.927
R14583 Iout.n554 Iout.t51 239.927
R14584 Iout.n434 Iout.t232 239.927
R14585 Iout.n438 Iout.t156 239.927
R14586 Iout.n441 Iout.t42 239.927
R14587 Iout.n432 Iout.t134 239.927
R14588 Iout.n418 Iout.t128 239.927
R14589 Iout.n416 Iout.t90 239.927
R14590 Iout.n402 Iout.t190 239.927
R14591 Iout.n357 Iout.t138 239.927
R14592 Iout.n360 Iout.t210 239.927
R14593 Iout.n363 Iout.t147 239.927
R14594 Iout.n366 Iout.t25 239.927
R14595 Iout.n354 Iout.t102 239.927
R14596 Iout.n351 Iout.t194 239.927
R14597 Iout.n348 Iout.t172 239.927
R14598 Iout.n345 Iout.t207 239.927
R14599 Iout.n342 Iout.t155 239.927
R14600 Iout.n339 Iout.t59 239.927
R14601 Iout.n336 Iout.t223 239.927
R14602 Iout.n333 Iout.t74 239.927
R14603 Iout.n117 Iout.t34 239.927
R14604 Iout.n582 Iout.t123 239.927
R14605 Iout.n111 Iout.t250 239.927
R14606 Iout.n594 Iout.t117 239.927
R14607 Iout.n105 Iout.t203 239.927
R14608 Iout.n606 Iout.t205 239.927
R14609 Iout.n99 Iout.t132 239.927
R14610 Iout.n618 Iout.t64 239.927
R14611 Iout.n624 Iout.t152 239.927
R14612 Iout.n90 Iout.t20 239.927
R14613 Iout.n636 Iout.t140 239.927
R14614 Iout.n81 Iout.t131 239.927
R14615 Iout.n648 Iout.t220 239.927
R14616 Iout.n96 Iout.t253 239.927
R14617 Iout.n612 Iout.t57 239.927
R14618 Iout.n102 Iout.t93 239.927
R14619 Iout.n600 Iout.t70 239.927
R14620 Iout.n108 Iout.t211 239.927
R14621 Iout.n588 Iout.t231 239.927
R14622 Iout.n687 Iout.t105 239.927
R14623 Iout.n684 Iout.t31 239.927
R14624 Iout.n681 Iout.t39 239.927
R14625 Iout.n678 Iout.t143 239.927
R14626 Iout.n675 Iout.t47 239.927
R14627 Iout.n672 Iout.t186 239.927
R14628 Iout.n747 Iout.t236 239.927
R14629 Iout.n50 Iout.t200 239.927
R14630 Iout.n759 Iout.t137 239.927
R14631 Iout.n44 Iout.t201 239.927
R14632 Iout.n771 Iout.t35 239.927
R14633 Iout.n42 Iout.t184 239.927
R14634 Iout.n56 Iout.t69 239.927
R14635 Iout.n735 Iout.t97 239.927
R14636 Iout.n62 Iout.t92 239.927
R14637 Iout.n723 Iout.t100 239.927
R14638 Iout.n717 Iout.t146 239.927
R14639 Iout.n65 Iout.t61 239.927
R14640 Iout.n729 Iout.t217 239.927
R14641 Iout.n59 Iout.t24 239.927
R14642 Iout.n805 Iout.t160 239.927
R14643 Iout.n808 Iout.t239 239.927
R14644 Iout.n811 Iout.t202 239.927
R14645 Iout.n814 Iout.t119 239.927
R14646 Iout.n817 Iout.t19 239.927
R14647 Iout.n820 Iout.t63 239.927
R14648 Iout.n823 Iout.t166 239.927
R14649 Iout.n802 Iout.t243 239.927
R14650 Iout.n799 Iout.t192 239.927
R14651 Iout.n890 Iout.t165 239.927
R14652 Iout.n888 Iout.t71 239.927
R14653 Iout.n881 Iout.t56 239.927
R14654 Iout.n869 Iout.t176 239.927
R14655 Iout.n867 Iout.t219 239.927
R14656 Iout.n855 Iout.t130 239.927
R14657 Iout.n853 Iout.t66 239.927
R14658 Iout.n841 Iout.t129 239.927
R14659 Iout.n839 Iout.t11 239.927
R14660 Iout.n827 Iout.t141 239.927
R14661 Iout.n883 Iout.t150 239.927
R14662 Iout.n895 Iout.t76 239.927
R14663 Iout.n897 Iout.t14 239.927
R14664 Iout.n909 Iout.t254 239.927
R14665 Iout.n911 Iout.t62 239.927
R14666 Iout.n923 Iout.t33 239.927
R14667 Iout.n926 Iout.t115 239.927
R14668 Iout.n22 Iout.t79 239.927
R14669 Iout.n876 Iout.t204 239.927
R14670 Iout.n874 Iout.t55 239.927
R14671 Iout.n862 Iout.t251 239.927
R14672 Iout.n860 Iout.t153 239.927
R14673 Iout.n848 Iout.t215 239.927
R14674 Iout.n846 Iout.t144 239.927
R14675 Iout.n834 Iout.t30 239.927
R14676 Iout.n832 Iout.t241 239.927
R14677 Iout.n902 Iout.t65 239.927
R14678 Iout.n904 Iout.t206 239.927
R14679 Iout.n916 Iout.t213 239.927
R14680 Iout.n918 Iout.t99 239.927
R14681 Iout.n931 Iout.t179 239.927
R14682 Iout.n934 Iout.t224 239.927
R14683 Iout.n796 Iout.t187 239.927
R14684 Iout.n793 Iout.t77 239.927
R14685 Iout.n790 Iout.t83 239.927
R14686 Iout.n787 Iout.t4 239.927
R14687 Iout.n784 Iout.t26 239.927
R14688 Iout.n781 Iout.t87 239.927
R14689 Iout.n938 Iout.t235 239.927
R14690 Iout.n741 Iout.t103 239.927
R14691 Iout.n53 Iout.t120 239.927
R14692 Iout.n753 Iout.t151 239.927
R14693 Iout.n47 Iout.t94 239.927
R14694 Iout.n765 Iout.t252 239.927
R14695 Iout.n38 Iout.t44 239.927
R14696 Iout.n777 Iout.t60 239.927
R14697 Iout.n71 Iout.t112 239.927
R14698 Iout.n705 Iout.t154 239.927
R14699 Iout.n77 Iout.t110 239.927
R14700 Iout.n944 Iout.t5 239.927
R14701 Iout.n19 Iout.t10 239.927
R14702 Iout.n68 Iout.t85 239.927
R14703 Iout.n711 Iout.t109 239.927
R14704 Iout.n74 Iout.t136 239.927
R14705 Iout.n699 Iout.t222 239.927
R14706 Iout.n950 Iout.t238 239.927
R14707 Iout.n953 Iout.t15 239.927
R14708 Iout.n669 Iout.t164 239.927
R14709 Iout.n666 Iout.t86 239.927
R14710 Iout.n663 Iout.t58 239.927
R14711 Iout.n660 Iout.t41 239.927
R14712 Iout.n657 Iout.t96 239.927
R14713 Iout.n654 Iout.t221 239.927
R14714 Iout.n690 Iout.t242 239.927
R14715 Iout.n695 Iout.t82 239.927
R14716 Iout.n692 Iout.t183 239.927
R14717 Iout.n957 Iout.t95 239.927
R14718 Iout.n114 Iout.t175 239.927
R14719 Iout.n576 Iout.t45 239.927
R14720 Iout.n573 Iout.t68 239.927
R14721 Iout.n963 Iout.t36 239.927
R14722 Iout.n14 Iout.t32 239.927
R14723 Iout.n93 Iout.t173 239.927
R14724 Iout.n630 Iout.t9 239.927
R14725 Iout.n87 Iout.t52 239.927
R14726 Iout.n642 Iout.t180 239.927
R14727 Iout.n85 Iout.t50 239.927
R14728 Iout.n563 Iout.t114 239.927
R14729 Iout.n969 Iout.t122 239.927
R14730 Iout.n972 Iout.t1 239.927
R14731 Iout.n569 Iout.t237 239.927
R14732 Iout.n123 Iout.t168 239.927
R14733 Iout.n120 Iout.t6 239.927
R14734 Iout.n976 Iout.t107 239.927
R14735 Iout.n400 Iout.t182 239.927
R14736 Iout.n386 Iout.t27 239.927
R14737 Iout.n384 Iout.t104 239.927
R14738 Iout.n370 Iout.t209 239.927
R14739 Iout.n982 Iout.t240 239.927
R14740 Iout.n9 Iout.t75 239.927
R14741 Iout.n127 Iout.t101 239.927
R14742 Iout.n988 Iout.t111 239.927
R14743 Iout.n991 Iout.t38 239.927
R14744 Iout.n323 Iout.t121 239.927
R14745 Iout.n326 Iout.t73 239.927
R14746 Iout.n329 Iout.t49 239.927
R14747 Iout.n995 Iout.t53 239.927
R14748 Iout.n1001 Iout.t124 239.927
R14749 Iout.n4 Iout.t234 239.927
R14750 Iout.n295 Iout.t177 239.927
R14751 Iout.n172 Iout.t91 239.927
R14752 Iout.n1014 Iout.t98 239.927
R14753 Iout.n1021 Iout.n1020 7.9105
R14754 Iout.n510 Iout.n509 7.9105
R14755 Iout.n514 Iout.n513 7.9105
R14756 Iout.n508 Iout.n507 7.9105
R14757 Iout.n505 Iout.n504 7.9105
R14758 Iout.n501 Iout.n500 7.9105
R14759 Iout.n193 Iout.n192 7.9105
R14760 Iout.n196 Iout.n195 7.9105
R14761 Iout.n200 Iout.n199 7.9105
R14762 Iout.n203 Iout.n202 7.9105
R14763 Iout.n207 Iout.n206 7.9105
R14764 Iout.n211 Iout.n210 7.9105
R14765 Iout.n215 Iout.n214 7.9105
R14766 Iout.n219 Iout.n218 7.9105
R14767 Iout.n223 Iout.n222 7.9105
R14768 Iout.n227 Iout.n226 7.9105
R14769 Iout.n233 Iout.n232 7.9105
R14770 Iout.n236 Iout.n235 7.9105
R14771 Iout.n239 Iout.n238 7.9105
R14772 Iout.n242 Iout.n241 7.9105
R14773 Iout.n245 Iout.n244 7.9105
R14774 Iout.n248 Iout.n247 7.9105
R14775 Iout.n251 Iout.n250 7.9105
R14776 Iout.n256 Iout.n255 7.9105
R14777 Iout.n253 Iout.n252 7.9105
R14778 Iout.n490 Iout.n489 7.9105
R14779 Iout.n495 Iout.n494 7.9105
R14780 Iout.n492 Iout.n491 7.9105
R14781 Iout.n520 Iout.n519 7.9105
R14782 Iout.n150 Iout.n149 7.9105
R14783 Iout.n147 Iout.n146 7.9105
R14784 Iout.n1011 Iout.n1010 7.9105
R14785 Iout.n1008 Iout.n1007 7.9105
R14786 Iout.n141 Iout.n140 7.9105
R14787 Iout.n144 Iout.n143 7.9105
R14788 Iout.n526 Iout.n525 7.9105
R14789 Iout.n481 Iout.n480 7.9105
R14790 Iout.n484 Iout.n483 7.9105
R14791 Iout.n479 Iout.n478 7.9105
R14792 Iout.n260 Iout.n259 7.9105
R14793 Iout.n187 Iout.n186 7.9105
R14794 Iout.n272 Iout.n271 7.9105
R14795 Iout.n181 Iout.n180 7.9105
R14796 Iout.n284 Iout.n283 7.9105
R14797 Iout.n175 Iout.n174 7.9105
R14798 Iout.n169 Iout.n168 7.9105
R14799 Iout.n302 Iout.n301 7.9105
R14800 Iout.n290 Iout.n289 7.9105
R14801 Iout.n178 Iout.n177 7.9105
R14802 Iout.n278 Iout.n277 7.9105
R14803 Iout.n184 Iout.n183 7.9105
R14804 Iout.n266 Iout.n265 7.9105
R14805 Iout.n190 Iout.n189 7.9105
R14806 Iout.n473 Iout.n472 7.9105
R14807 Iout.n470 Iout.n469 7.9105
R14808 Iout.n157 Iout.n156 7.9105
R14809 Iout.n532 Iout.n531 7.9105
R14810 Iout.n535 Iout.n534 7.9105
R14811 Iout.n537 Iout.n536 7.9105
R14812 Iout.n134 Iout.n133 7.9105
R14813 Iout.n137 Iout.n136 7.9105
R14814 Iout.n543 Iout.n542 7.9105
R14815 Iout.n461 Iout.n460 7.9105
R14816 Iout.n464 Iout.n463 7.9105
R14817 Iout.n459 Iout.n458 7.9105
R14818 Iout.n306 Iout.n305 7.9105
R14819 Iout.n309 Iout.n308 7.9105
R14820 Iout.n312 Iout.n311 7.9105
R14821 Iout.n315 Iout.n314 7.9105
R14822 Iout.n318 Iout.n317 7.9105
R14823 Iout.n321 Iout.n320 7.9105
R14824 Iout.n393 Iout.n392 7.9105
R14825 Iout.n379 Iout.n378 7.9105
R14826 Iout.n377 Iout.n376 7.9105
R14827 Iout.n395 Iout.n394 7.9105
R14828 Iout.n409 Iout.n408 7.9105
R14829 Iout.n411 Iout.n410 7.9105
R14830 Iout.n425 Iout.n424 7.9105
R14831 Iout.n427 Iout.n426 7.9105
R14832 Iout.n448 Iout.n447 7.9105
R14833 Iout.n453 Iout.n452 7.9105
R14834 Iout.n450 Iout.n449 7.9105
R14835 Iout.n549 Iout.n548 7.9105
R14836 Iout.n131 Iout.n130 7.9105
R14837 Iout.n560 Iout.n559 7.9105
R14838 Iout.n558 Iout.n557 7.9105
R14839 Iout.n555 Iout.n554 7.9105
R14840 Iout.n435 Iout.n434 7.9105
R14841 Iout.n439 Iout.n438 7.9105
R14842 Iout.n442 Iout.n441 7.9105
R14843 Iout.n433 Iout.n432 7.9105
R14844 Iout.n419 Iout.n418 7.9105
R14845 Iout.n417 Iout.n416 7.9105
R14846 Iout.n403 Iout.n402 7.9105
R14847 Iout.n358 Iout.n357 7.9105
R14848 Iout.n361 Iout.n360 7.9105
R14849 Iout.n364 Iout.n363 7.9105
R14850 Iout.n367 Iout.n366 7.9105
R14851 Iout.n355 Iout.n354 7.9105
R14852 Iout.n352 Iout.n351 7.9105
R14853 Iout.n349 Iout.n348 7.9105
R14854 Iout.n346 Iout.n345 7.9105
R14855 Iout.n343 Iout.n342 7.9105
R14856 Iout.n340 Iout.n339 7.9105
R14857 Iout.n337 Iout.n336 7.9105
R14858 Iout.n334 Iout.n333 7.9105
R14859 Iout.n118 Iout.n117 7.9105
R14860 Iout.n583 Iout.n582 7.9105
R14861 Iout.n112 Iout.n111 7.9105
R14862 Iout.n595 Iout.n594 7.9105
R14863 Iout.n106 Iout.n105 7.9105
R14864 Iout.n607 Iout.n606 7.9105
R14865 Iout.n100 Iout.n99 7.9105
R14866 Iout.n619 Iout.n618 7.9105
R14867 Iout.n625 Iout.n624 7.9105
R14868 Iout.n91 Iout.n90 7.9105
R14869 Iout.n637 Iout.n636 7.9105
R14870 Iout.n82 Iout.n81 7.9105
R14871 Iout.n649 Iout.n648 7.9105
R14872 Iout.n97 Iout.n96 7.9105
R14873 Iout.n613 Iout.n612 7.9105
R14874 Iout.n103 Iout.n102 7.9105
R14875 Iout.n601 Iout.n600 7.9105
R14876 Iout.n109 Iout.n108 7.9105
R14877 Iout.n589 Iout.n588 7.9105
R14878 Iout.n688 Iout.n687 7.9105
R14879 Iout.n685 Iout.n684 7.9105
R14880 Iout.n682 Iout.n681 7.9105
R14881 Iout.n679 Iout.n678 7.9105
R14882 Iout.n676 Iout.n675 7.9105
R14883 Iout.n673 Iout.n672 7.9105
R14884 Iout.n748 Iout.n747 7.9105
R14885 Iout.n51 Iout.n50 7.9105
R14886 Iout.n760 Iout.n759 7.9105
R14887 Iout.n45 Iout.n44 7.9105
R14888 Iout.n772 Iout.n771 7.9105
R14889 Iout.n43 Iout.n42 7.9105
R14890 Iout.n57 Iout.n56 7.9105
R14891 Iout.n736 Iout.n735 7.9105
R14892 Iout.n63 Iout.n62 7.9105
R14893 Iout.n724 Iout.n723 7.9105
R14894 Iout.n718 Iout.n717 7.9105
R14895 Iout.n66 Iout.n65 7.9105
R14896 Iout.n730 Iout.n729 7.9105
R14897 Iout.n60 Iout.n59 7.9105
R14898 Iout.n806 Iout.n805 7.9105
R14899 Iout.n809 Iout.n808 7.9105
R14900 Iout.n812 Iout.n811 7.9105
R14901 Iout.n815 Iout.n814 7.9105
R14902 Iout.n818 Iout.n817 7.9105
R14903 Iout.n821 Iout.n820 7.9105
R14904 Iout.n824 Iout.n823 7.9105
R14905 Iout.n803 Iout.n802 7.9105
R14906 Iout.n800 Iout.n799 7.9105
R14907 Iout.n891 Iout.n890 7.9105
R14908 Iout.n889 Iout.n888 7.9105
R14909 Iout.n882 Iout.n881 7.9105
R14910 Iout.n870 Iout.n869 7.9105
R14911 Iout.n868 Iout.n867 7.9105
R14912 Iout.n856 Iout.n855 7.9105
R14913 Iout.n854 Iout.n853 7.9105
R14914 Iout.n842 Iout.n841 7.9105
R14915 Iout.n840 Iout.n839 7.9105
R14916 Iout.n828 Iout.n827 7.9105
R14917 Iout.n884 Iout.n883 7.9105
R14918 Iout.n896 Iout.n895 7.9105
R14919 Iout.n898 Iout.n897 7.9105
R14920 Iout.n910 Iout.n909 7.9105
R14921 Iout.n912 Iout.n911 7.9105
R14922 Iout.n924 Iout.n923 7.9105
R14923 Iout.n927 Iout.n926 7.9105
R14924 Iout.n23 Iout.n22 7.9105
R14925 Iout.n877 Iout.n876 7.9105
R14926 Iout.n875 Iout.n874 7.9105
R14927 Iout.n863 Iout.n862 7.9105
R14928 Iout.n861 Iout.n860 7.9105
R14929 Iout.n849 Iout.n848 7.9105
R14930 Iout.n847 Iout.n846 7.9105
R14931 Iout.n835 Iout.n834 7.9105
R14932 Iout.n833 Iout.n832 7.9105
R14933 Iout.n903 Iout.n902 7.9105
R14934 Iout.n905 Iout.n904 7.9105
R14935 Iout.n917 Iout.n916 7.9105
R14936 Iout.n919 Iout.n918 7.9105
R14937 Iout.n932 Iout.n931 7.9105
R14938 Iout.n935 Iout.n934 7.9105
R14939 Iout.n797 Iout.n796 7.9105
R14940 Iout.n794 Iout.n793 7.9105
R14941 Iout.n791 Iout.n790 7.9105
R14942 Iout.n788 Iout.n787 7.9105
R14943 Iout.n785 Iout.n784 7.9105
R14944 Iout.n782 Iout.n781 7.9105
R14945 Iout.n939 Iout.n938 7.9105
R14946 Iout.n742 Iout.n741 7.9105
R14947 Iout.n54 Iout.n53 7.9105
R14948 Iout.n754 Iout.n753 7.9105
R14949 Iout.n48 Iout.n47 7.9105
R14950 Iout.n766 Iout.n765 7.9105
R14951 Iout.n39 Iout.n38 7.9105
R14952 Iout.n778 Iout.n777 7.9105
R14953 Iout.n72 Iout.n71 7.9105
R14954 Iout.n706 Iout.n705 7.9105
R14955 Iout.n78 Iout.n77 7.9105
R14956 Iout.n945 Iout.n944 7.9105
R14957 Iout.n20 Iout.n19 7.9105
R14958 Iout.n69 Iout.n68 7.9105
R14959 Iout.n712 Iout.n711 7.9105
R14960 Iout.n75 Iout.n74 7.9105
R14961 Iout.n700 Iout.n699 7.9105
R14962 Iout.n951 Iout.n950 7.9105
R14963 Iout.n954 Iout.n953 7.9105
R14964 Iout.n670 Iout.n669 7.9105
R14965 Iout.n667 Iout.n666 7.9105
R14966 Iout.n664 Iout.n663 7.9105
R14967 Iout.n661 Iout.n660 7.9105
R14968 Iout.n658 Iout.n657 7.9105
R14969 Iout.n655 Iout.n654 7.9105
R14970 Iout.n691 Iout.n690 7.9105
R14971 Iout.n696 Iout.n695 7.9105
R14972 Iout.n693 Iout.n692 7.9105
R14973 Iout.n958 Iout.n957 7.9105
R14974 Iout.n115 Iout.n114 7.9105
R14975 Iout.n577 Iout.n576 7.9105
R14976 Iout.n574 Iout.n573 7.9105
R14977 Iout.n964 Iout.n963 7.9105
R14978 Iout.n15 Iout.n14 7.9105
R14979 Iout.n94 Iout.n93 7.9105
R14980 Iout.n631 Iout.n630 7.9105
R14981 Iout.n88 Iout.n87 7.9105
R14982 Iout.n643 Iout.n642 7.9105
R14983 Iout.n86 Iout.n85 7.9105
R14984 Iout.n564 Iout.n563 7.9105
R14985 Iout.n970 Iout.n969 7.9105
R14986 Iout.n973 Iout.n972 7.9105
R14987 Iout.n570 Iout.n569 7.9105
R14988 Iout.n124 Iout.n123 7.9105
R14989 Iout.n121 Iout.n120 7.9105
R14990 Iout.n977 Iout.n976 7.9105
R14991 Iout.n401 Iout.n400 7.9105
R14992 Iout.n387 Iout.n386 7.9105
R14993 Iout.n385 Iout.n384 7.9105
R14994 Iout.n371 Iout.n370 7.9105
R14995 Iout.n983 Iout.n982 7.9105
R14996 Iout.n10 Iout.n9 7.9105
R14997 Iout.n128 Iout.n127 7.9105
R14998 Iout.n989 Iout.n988 7.9105
R14999 Iout.n992 Iout.n991 7.9105
R15000 Iout.n324 Iout.n323 7.9105
R15001 Iout.n327 Iout.n326 7.9105
R15002 Iout.n330 Iout.n329 7.9105
R15003 Iout.n996 Iout.n995 7.9105
R15004 Iout.n1002 Iout.n1001 7.9105
R15005 Iout.n5 Iout.n4 7.9105
R15006 Iout.n296 Iout.n295 7.9105
R15007 Iout.n173 Iout.n172 7.9105
R15008 Iout.n1015 Iout.n1014 7.9105
R15009 Iout.n886 Iout.n885 3.86101
R15010 Iout.n880 Iout.n879 3.86101
R15011 Iout.n894 Iout.n893 3.86101
R15012 Iout.n872 Iout.n871 3.86101
R15013 Iout.n900 Iout.n899 3.86101
R15014 Iout.n866 Iout.n865 3.86101
R15015 Iout.n908 Iout.n907 3.86101
R15016 Iout.n858 Iout.n857 3.86101
R15017 Iout.n914 Iout.n913 3.86101
R15018 Iout.n852 Iout.n851 3.86101
R15019 Iout.n922 Iout.n921 3.86101
R15020 Iout.n844 Iout.n843 3.86101
R15021 Iout.n929 Iout.n928 3.86101
R15022 Iout.n838 Iout.n837 3.86101
R15023 Iout.n925 Iout.n21 3.86101
R15024 Iout.n830 Iout.n829 3.86101
R15025 Iout.n879 Iout.n878 3.4105
R15026 Iout.n887 Iout.n886 3.4105
R15027 Iout.n893 Iout.n892 3.4105
R15028 Iout.n798 Iout.n28 3.4105
R15029 Iout.n801 Iout.n29 3.4105
R15030 Iout.n804 Iout.n30 3.4105
R15031 Iout.n807 Iout.n31 3.4105
R15032 Iout.n873 Iout.n872 3.4105
R15033 Iout.n744 Iout.n743 3.4105
R15034 Iout.n740 Iout.n739 3.4105
R15035 Iout.n732 Iout.n731 3.4105
R15036 Iout.n728 Iout.n727 3.4105
R15037 Iout.n720 Iout.n719 3.4105
R15038 Iout.n795 Iout.n27 3.4105
R15039 Iout.n901 Iout.n900 3.4105
R15040 Iout.n722 Iout.n721 3.4105
R15041 Iout.n726 Iout.n725 3.4105
R15042 Iout.n734 Iout.n733 3.4105
R15043 Iout.n738 Iout.n737 3.4105
R15044 Iout.n746 Iout.n745 3.4105
R15045 Iout.n750 Iout.n749 3.4105
R15046 Iout.n752 Iout.n751 3.4105
R15047 Iout.n810 Iout.n32 3.4105
R15048 Iout.n865 Iout.n864 3.4105
R15049 Iout.n668 Iout.n55 3.4105
R15050 Iout.n671 Iout.n58 3.4105
R15051 Iout.n674 Iout.n61 3.4105
R15052 Iout.n677 Iout.n64 3.4105
R15053 Iout.n680 Iout.n67 3.4105
R15054 Iout.n683 Iout.n70 3.4105
R15055 Iout.n686 Iout.n73 3.4105
R15056 Iout.n714 Iout.n713 3.4105
R15057 Iout.n716 Iout.n715 3.4105
R15058 Iout.n792 Iout.n26 3.4105
R15059 Iout.n907 Iout.n906 3.4105
R15060 Iout.n587 Iout.n586 3.4105
R15061 Iout.n591 Iout.n590 3.4105
R15062 Iout.n599 Iout.n598 3.4105
R15063 Iout.n603 Iout.n602 3.4105
R15064 Iout.n611 Iout.n610 3.4105
R15065 Iout.n615 Iout.n614 3.4105
R15066 Iout.n623 Iout.n622 3.4105
R15067 Iout.n627 Iout.n626 3.4105
R15068 Iout.n665 Iout.n52 3.4105
R15069 Iout.n758 Iout.n757 3.4105
R15070 Iout.n756 Iout.n755 3.4105
R15071 Iout.n813 Iout.n33 3.4105
R15072 Iout.n859 Iout.n858 3.4105
R15073 Iout.n629 Iout.n628 3.4105
R15074 Iout.n621 Iout.n620 3.4105
R15075 Iout.n617 Iout.n616 3.4105
R15076 Iout.n609 Iout.n608 3.4105
R15077 Iout.n605 Iout.n604 3.4105
R15078 Iout.n597 Iout.n596 3.4105
R15079 Iout.n593 Iout.n592 3.4105
R15080 Iout.n585 Iout.n584 3.4105
R15081 Iout.n581 Iout.n580 3.4105
R15082 Iout.n579 Iout.n578 3.4105
R15083 Iout.n689 Iout.n76 3.4105
R15084 Iout.n710 Iout.n709 3.4105
R15085 Iout.n708 Iout.n707 3.4105
R15086 Iout.n789 Iout.n25 3.4105
R15087 Iout.n915 Iout.n914 3.4105
R15088 Iout.n572 Iout.n571 3.4105
R15089 Iout.n335 Iout.n116 3.4105
R15090 Iout.n338 Iout.n113 3.4105
R15091 Iout.n341 Iout.n110 3.4105
R15092 Iout.n344 Iout.n107 3.4105
R15093 Iout.n347 Iout.n104 3.4105
R15094 Iout.n350 Iout.n101 3.4105
R15095 Iout.n353 Iout.n98 3.4105
R15096 Iout.n356 Iout.n95 3.4105
R15097 Iout.n359 Iout.n92 3.4105
R15098 Iout.n633 Iout.n632 3.4105
R15099 Iout.n635 Iout.n634 3.4105
R15100 Iout.n662 Iout.n49 3.4105
R15101 Iout.n762 Iout.n761 3.4105
R15102 Iout.n764 Iout.n763 3.4105
R15103 Iout.n816 Iout.n34 3.4105
R15104 Iout.n851 Iout.n850 3.4105
R15105 Iout.n399 Iout.n398 3.4105
R15106 Iout.n405 Iout.n404 3.4105
R15107 Iout.n415 Iout.n414 3.4105
R15108 Iout.n421 Iout.n420 3.4105
R15109 Iout.n431 Iout.n430 3.4105
R15110 Iout.n444 Iout.n443 3.4105
R15111 Iout.n440 Iout.n159 3.4105
R15112 Iout.n437 Iout.n436 3.4105
R15113 Iout.n553 Iout.n552 3.4105
R15114 Iout.n556 Iout.n119 3.4105
R15115 Iout.n562 Iout.n561 3.4105
R15116 Iout.n568 Iout.n567 3.4105
R15117 Iout.n566 Iout.n565 3.4105
R15118 Iout.n575 Iout.n79 3.4105
R15119 Iout.n698 Iout.n697 3.4105
R15120 Iout.n702 Iout.n701 3.4105
R15121 Iout.n704 Iout.n703 3.4105
R15122 Iout.n786 Iout.n24 3.4105
R15123 Iout.n921 Iout.n920 3.4105
R15124 Iout.n129 Iout.n125 3.4105
R15125 Iout.n547 Iout.n546 3.4105
R15126 Iout.n551 Iout.n550 3.4105
R15127 Iout.n451 Iout.n158 3.4105
R15128 Iout.n455 Iout.n454 3.4105
R15129 Iout.n446 Iout.n445 3.4105
R15130 Iout.n429 Iout.n428 3.4105
R15131 Iout.n423 Iout.n422 3.4105
R15132 Iout.n413 Iout.n412 3.4105
R15133 Iout.n407 Iout.n406 3.4105
R15134 Iout.n397 Iout.n396 3.4105
R15135 Iout.n391 Iout.n390 3.4105
R15136 Iout.n389 Iout.n388 3.4105
R15137 Iout.n362 Iout.n89 3.4105
R15138 Iout.n641 Iout.n640 3.4105
R15139 Iout.n639 Iout.n638 3.4105
R15140 Iout.n659 Iout.n46 3.4105
R15141 Iout.n770 Iout.n769 3.4105
R15142 Iout.n768 Iout.n767 3.4105
R15143 Iout.n819 Iout.n35 3.4105
R15144 Iout.n845 Iout.n844 3.4105
R15145 Iout.n325 Iout.n165 3.4105
R15146 Iout.n322 Iout.n164 3.4105
R15147 Iout.n319 Iout.n163 3.4105
R15148 Iout.n316 Iout.n162 3.4105
R15149 Iout.n313 Iout.n161 3.4105
R15150 Iout.n310 Iout.n160 3.4105
R15151 Iout.n307 Iout.n155 3.4105
R15152 Iout.n457 Iout.n456 3.4105
R15153 Iout.n466 Iout.n465 3.4105
R15154 Iout.n462 Iout.n126 3.4105
R15155 Iout.n545 Iout.n544 3.4105
R15156 Iout.n541 Iout.n540 3.4105
R15157 Iout.n135 Iout.n3 3.4105
R15158 Iout.n987 Iout.n986 3.4105
R15159 Iout.n985 Iout.n984 3.4105
R15160 Iout.n122 Iout.n8 3.4105
R15161 Iout.n968 Iout.n967 3.4105
R15162 Iout.n966 Iout.n965 3.4105
R15163 Iout.n694 Iout.n13 3.4105
R15164 Iout.n949 Iout.n948 3.4105
R15165 Iout.n947 Iout.n946 3.4105
R15166 Iout.n783 Iout.n18 3.4105
R15167 Iout.n930 Iout.n929 3.4105
R15168 Iout.n1004 Iout.n1003 3.4105
R15169 Iout.n539 Iout.n538 3.4105
R15170 Iout.n533 Iout.n132 3.4105
R15171 Iout.n530 Iout.n529 3.4105
R15172 Iout.n468 Iout.n467 3.4105
R15173 Iout.n471 Iout.n153 3.4105
R15174 Iout.n475 Iout.n474 3.4105
R15175 Iout.n264 Iout.n263 3.4105
R15176 Iout.n268 Iout.n267 3.4105
R15177 Iout.n276 Iout.n275 3.4105
R15178 Iout.n280 Iout.n279 3.4105
R15179 Iout.n288 Iout.n287 3.4105
R15180 Iout.n292 Iout.n291 3.4105
R15181 Iout.n300 Iout.n299 3.4105
R15182 Iout.n328 Iout.n166 3.4105
R15183 Iout.n381 Iout.n380 3.4105
R15184 Iout.n383 Iout.n382 3.4105
R15185 Iout.n365 Iout.n83 3.4105
R15186 Iout.n645 Iout.n644 3.4105
R15187 Iout.n647 Iout.n646 3.4105
R15188 Iout.n656 Iout.n40 3.4105
R15189 Iout.n774 Iout.n773 3.4105
R15190 Iout.n776 Iout.n775 3.4105
R15191 Iout.n822 Iout.n36 3.4105
R15192 Iout.n837 Iout.n836 3.4105
R15193 Iout.n298 Iout.n297 3.4105
R15194 Iout.n294 Iout.n293 3.4105
R15195 Iout.n286 Iout.n285 3.4105
R15196 Iout.n282 Iout.n281 3.4105
R15197 Iout.n274 Iout.n273 3.4105
R15198 Iout.n270 Iout.n269 3.4105
R15199 Iout.n262 Iout.n261 3.4105
R15200 Iout.n477 Iout.n476 3.4105
R15201 Iout.n486 Iout.n485 3.4105
R15202 Iout.n482 Iout.n151 3.4105
R15203 Iout.n528 Iout.n527 3.4105
R15204 Iout.n524 Iout.n523 3.4105
R15205 Iout.n142 Iout.n138 3.4105
R15206 Iout.n1006 Iout.n1005 3.4105
R15207 Iout.n1009 Iout.n0 3.4105
R15208 Iout.n1000 Iout.n999 3.4105
R15209 Iout.n998 Iout.n997 3.4105
R15210 Iout.n990 Iout.n6 3.4105
R15211 Iout.n981 Iout.n980 3.4105
R15212 Iout.n979 Iout.n978 3.4105
R15213 Iout.n971 Iout.n11 3.4105
R15214 Iout.n962 Iout.n961 3.4105
R15215 Iout.n960 Iout.n959 3.4105
R15216 Iout.n952 Iout.n16 3.4105
R15217 Iout.n943 Iout.n942 3.4105
R15218 Iout.n941 Iout.n940 3.4105
R15219 Iout.n933 Iout.n21 3.4105
R15220 Iout.n1017 Iout.n1016 3.4105
R15221 Iout.n148 Iout.n2 3.4105
R15222 Iout.n518 Iout.n517 3.4105
R15223 Iout.n522 Iout.n521 3.4105
R15224 Iout.n493 Iout.n139 3.4105
R15225 Iout.n497 Iout.n496 3.4105
R15226 Iout.n488 Iout.n487 3.4105
R15227 Iout.n254 Iout.n154 3.4105
R15228 Iout.n258 Iout.n257 3.4105
R15229 Iout.n249 Iout.n188 3.4105
R15230 Iout.n246 Iout.n185 3.4105
R15231 Iout.n243 Iout.n182 3.4105
R15232 Iout.n240 Iout.n179 3.4105
R15233 Iout.n237 Iout.n176 3.4105
R15234 Iout.n234 Iout.n170 3.4105
R15235 Iout.n231 Iout.n230 3.4105
R15236 Iout.n171 Iout.n167 3.4105
R15237 Iout.n304 Iout.n303 3.4105
R15238 Iout.n332 Iout.n331 3.4105
R15239 Iout.n375 Iout.n374 3.4105
R15240 Iout.n373 Iout.n372 3.4105
R15241 Iout.n369 Iout.n368 3.4105
R15242 Iout.n84 Iout.n80 3.4105
R15243 Iout.n651 Iout.n650 3.4105
R15244 Iout.n653 Iout.n652 3.4105
R15245 Iout.n41 Iout.n37 3.4105
R15246 Iout.n780 Iout.n779 3.4105
R15247 Iout.n826 Iout.n825 3.4105
R15248 Iout.n831 Iout.n830 3.4105
R15249 Iout.n229 Iout.n228 3.4105
R15250 Iout.n225 Iout.n224 3.4105
R15251 Iout.n221 Iout.n220 3.4105
R15252 Iout.n217 Iout.n216 3.4105
R15253 Iout.n213 Iout.n212 3.4105
R15254 Iout.n209 Iout.n208 3.4105
R15255 Iout.n205 Iout.n204 3.4105
R15256 Iout.n201 Iout.n191 3.4105
R15257 Iout.n198 Iout.n197 3.4105
R15258 Iout.n194 Iout.n152 3.4105
R15259 Iout.n499 Iout.n498 3.4105
R15260 Iout.n503 Iout.n502 3.4105
R15261 Iout.n506 Iout.n145 3.4105
R15262 Iout.n516 Iout.n515 3.4105
R15263 Iout.n512 Iout.n511 3.4105
R15264 Iout.n1019 Iout.n1018 3.4105
R15265 Iout.n936 Iout.n23 1.43848
R15266 Iout.n936 Iout.n935 1.34612
R15267 Iout.n939 Iout.n937 1.34612
R15268 Iout.n20 Iout.n17 1.34612
R15269 Iout.n955 Iout.n954 1.34612
R15270 Iout.n958 Iout.n956 1.34612
R15271 Iout.n15 Iout.n12 1.34612
R15272 Iout.n974 Iout.n973 1.34612
R15273 Iout.n977 Iout.n975 1.34612
R15274 Iout.n10 Iout.n7 1.34612
R15275 Iout.n993 Iout.n992 1.34612
R15276 Iout.n996 Iout.n994 1.34612
R15277 Iout.n5 Iout.n1 1.34612
R15278 Iout.n1012 Iout.n1011 1.34612
R15279 Iout.n1015 Iout.n1013 1.34612
R15280 Iout.n1022 Iout.n1021 1.34612
R15281 Iout.n197 Iout.n154 0.451012
R15282 Iout.n476 Iout.n154 0.451012
R15283 Iout.n476 Iout.n475 0.451012
R15284 Iout.n475 Iout.n155 0.451012
R15285 Iout.n445 Iout.n155 0.451012
R15286 Iout.n445 Iout.n444 0.451012
R15287 Iout.n444 Iout.n107 0.451012
R15288 Iout.n604 Iout.n107 0.451012
R15289 Iout.n604 Iout.n603 0.451012
R15290 Iout.n603 Iout.n64 0.451012
R15291 Iout.n733 Iout.n64 0.451012
R15292 Iout.n733 Iout.n732 0.451012
R15293 Iout.n732 Iout.n29 0.451012
R15294 Iout.n886 Iout.n29 0.451012
R15295 Iout.n258 Iout.n191 0.451012
R15296 Iout.n262 Iout.n258 0.451012
R15297 Iout.n263 Iout.n262 0.451012
R15298 Iout.n263 Iout.n160 0.451012
R15299 Iout.n429 Iout.n160 0.451012
R15300 Iout.n430 Iout.n429 0.451012
R15301 Iout.n430 Iout.n104 0.451012
R15302 Iout.n609 Iout.n104 0.451012
R15303 Iout.n610 Iout.n609 0.451012
R15304 Iout.n610 Iout.n61 0.451012
R15305 Iout.n738 Iout.n61 0.451012
R15306 Iout.n739 Iout.n738 0.451012
R15307 Iout.n739 Iout.n30 0.451012
R15308 Iout.n879 Iout.n30 0.451012
R15309 Iout.n487 Iout.n152 0.451012
R15310 Iout.n487 Iout.n486 0.451012
R15311 Iout.n486 Iout.n153 0.451012
R15312 Iout.n456 Iout.n153 0.451012
R15313 Iout.n456 Iout.n455 0.451012
R15314 Iout.n455 Iout.n159 0.451012
R15315 Iout.n159 Iout.n110 0.451012
R15316 Iout.n597 Iout.n110 0.451012
R15317 Iout.n598 Iout.n597 0.451012
R15318 Iout.n598 Iout.n67 0.451012
R15319 Iout.n726 Iout.n67 0.451012
R15320 Iout.n727 Iout.n726 0.451012
R15321 Iout.n727 Iout.n28 0.451012
R15322 Iout.n893 Iout.n28 0.451012
R15323 Iout.n204 Iout.n188 0.451012
R15324 Iout.n269 Iout.n188 0.451012
R15325 Iout.n269 Iout.n268 0.451012
R15326 Iout.n268 Iout.n161 0.451012
R15327 Iout.n422 Iout.n161 0.451012
R15328 Iout.n422 Iout.n421 0.451012
R15329 Iout.n421 Iout.n101 0.451012
R15330 Iout.n616 Iout.n101 0.451012
R15331 Iout.n616 Iout.n615 0.451012
R15332 Iout.n615 Iout.n58 0.451012
R15333 Iout.n745 Iout.n58 0.451012
R15334 Iout.n745 Iout.n744 0.451012
R15335 Iout.n744 Iout.n31 0.451012
R15336 Iout.n872 Iout.n31 0.451012
R15337 Iout.n498 Iout.n497 0.451012
R15338 Iout.n497 Iout.n151 0.451012
R15339 Iout.n467 Iout.n151 0.451012
R15340 Iout.n467 Iout.n466 0.451012
R15341 Iout.n466 Iout.n158 0.451012
R15342 Iout.n436 Iout.n158 0.451012
R15343 Iout.n436 Iout.n113 0.451012
R15344 Iout.n592 Iout.n113 0.451012
R15345 Iout.n592 Iout.n591 0.451012
R15346 Iout.n591 Iout.n70 0.451012
R15347 Iout.n721 Iout.n70 0.451012
R15348 Iout.n721 Iout.n720 0.451012
R15349 Iout.n720 Iout.n27 0.451012
R15350 Iout.n900 Iout.n27 0.451012
R15351 Iout.n208 Iout.n185 0.451012
R15352 Iout.n274 Iout.n185 0.451012
R15353 Iout.n275 Iout.n274 0.451012
R15354 Iout.n275 Iout.n162 0.451012
R15355 Iout.n413 Iout.n162 0.451012
R15356 Iout.n414 Iout.n413 0.451012
R15357 Iout.n414 Iout.n98 0.451012
R15358 Iout.n621 Iout.n98 0.451012
R15359 Iout.n622 Iout.n621 0.451012
R15360 Iout.n622 Iout.n55 0.451012
R15361 Iout.n750 Iout.n55 0.451012
R15362 Iout.n751 Iout.n750 0.451012
R15363 Iout.n751 Iout.n32 0.451012
R15364 Iout.n865 Iout.n32 0.451012
R15365 Iout.n502 Iout.n139 0.451012
R15366 Iout.n528 Iout.n139 0.451012
R15367 Iout.n529 Iout.n528 0.451012
R15368 Iout.n529 Iout.n126 0.451012
R15369 Iout.n551 Iout.n126 0.451012
R15370 Iout.n552 Iout.n551 0.451012
R15371 Iout.n552 Iout.n116 0.451012
R15372 Iout.n585 Iout.n116 0.451012
R15373 Iout.n586 Iout.n585 0.451012
R15374 Iout.n586 Iout.n73 0.451012
R15375 Iout.n714 Iout.n73 0.451012
R15376 Iout.n715 Iout.n714 0.451012
R15377 Iout.n715 Iout.n26 0.451012
R15378 Iout.n907 Iout.n26 0.451012
R15379 Iout.n212 Iout.n182 0.451012
R15380 Iout.n281 Iout.n182 0.451012
R15381 Iout.n281 Iout.n280 0.451012
R15382 Iout.n280 Iout.n163 0.451012
R15383 Iout.n406 Iout.n163 0.451012
R15384 Iout.n406 Iout.n405 0.451012
R15385 Iout.n405 Iout.n95 0.451012
R15386 Iout.n628 Iout.n95 0.451012
R15387 Iout.n628 Iout.n627 0.451012
R15388 Iout.n627 Iout.n52 0.451012
R15389 Iout.n757 Iout.n52 0.451012
R15390 Iout.n757 Iout.n756 0.451012
R15391 Iout.n756 Iout.n33 0.451012
R15392 Iout.n858 Iout.n33 0.451012
R15393 Iout.n522 Iout.n145 0.451012
R15394 Iout.n523 Iout.n522 0.451012
R15395 Iout.n523 Iout.n132 0.451012
R15396 Iout.n545 Iout.n132 0.451012
R15397 Iout.n546 Iout.n545 0.451012
R15398 Iout.n546 Iout.n119 0.451012
R15399 Iout.n572 Iout.n119 0.451012
R15400 Iout.n580 Iout.n572 0.451012
R15401 Iout.n580 Iout.n579 0.451012
R15402 Iout.n579 Iout.n76 0.451012
R15403 Iout.n709 Iout.n76 0.451012
R15404 Iout.n709 Iout.n708 0.451012
R15405 Iout.n708 Iout.n25 0.451012
R15406 Iout.n914 Iout.n25 0.451012
R15407 Iout.n216 Iout.n179 0.451012
R15408 Iout.n286 Iout.n179 0.451012
R15409 Iout.n287 Iout.n286 0.451012
R15410 Iout.n287 Iout.n164 0.451012
R15411 Iout.n397 Iout.n164 0.451012
R15412 Iout.n398 Iout.n397 0.451012
R15413 Iout.n398 Iout.n92 0.451012
R15414 Iout.n633 Iout.n92 0.451012
R15415 Iout.n634 Iout.n633 0.451012
R15416 Iout.n634 Iout.n49 0.451012
R15417 Iout.n762 Iout.n49 0.451012
R15418 Iout.n763 Iout.n762 0.451012
R15419 Iout.n763 Iout.n34 0.451012
R15420 Iout.n851 Iout.n34 0.451012
R15421 Iout.n517 Iout.n516 0.451012
R15422 Iout.n517 Iout.n138 0.451012
R15423 Iout.n539 Iout.n138 0.451012
R15424 Iout.n540 Iout.n539 0.451012
R15425 Iout.n540 Iout.n125 0.451012
R15426 Iout.n562 Iout.n125 0.451012
R15427 Iout.n567 Iout.n562 0.451012
R15428 Iout.n567 Iout.n566 0.451012
R15429 Iout.n566 Iout.n79 0.451012
R15430 Iout.n698 Iout.n79 0.451012
R15431 Iout.n702 Iout.n698 0.451012
R15432 Iout.n703 Iout.n702 0.451012
R15433 Iout.n703 Iout.n24 0.451012
R15434 Iout.n921 Iout.n24 0.451012
R15435 Iout.n220 Iout.n176 0.451012
R15436 Iout.n293 Iout.n176 0.451012
R15437 Iout.n293 Iout.n292 0.451012
R15438 Iout.n292 Iout.n165 0.451012
R15439 Iout.n390 Iout.n165 0.451012
R15440 Iout.n390 Iout.n389 0.451012
R15441 Iout.n389 Iout.n89 0.451012
R15442 Iout.n640 Iout.n89 0.451012
R15443 Iout.n640 Iout.n639 0.451012
R15444 Iout.n639 Iout.n46 0.451012
R15445 Iout.n769 Iout.n46 0.451012
R15446 Iout.n769 Iout.n768 0.451012
R15447 Iout.n768 Iout.n35 0.451012
R15448 Iout.n844 Iout.n35 0.451012
R15449 Iout.n511 Iout.n2 0.451012
R15450 Iout.n1005 Iout.n2 0.451012
R15451 Iout.n1005 Iout.n1004 0.451012
R15452 Iout.n1004 Iout.n3 0.451012
R15453 Iout.n986 Iout.n3 0.451012
R15454 Iout.n986 Iout.n985 0.451012
R15455 Iout.n985 Iout.n8 0.451012
R15456 Iout.n967 Iout.n8 0.451012
R15457 Iout.n967 Iout.n966 0.451012
R15458 Iout.n966 Iout.n13 0.451012
R15459 Iout.n948 Iout.n13 0.451012
R15460 Iout.n948 Iout.n947 0.451012
R15461 Iout.n947 Iout.n18 0.451012
R15462 Iout.n929 Iout.n18 0.451012
R15463 Iout.n224 Iout.n170 0.451012
R15464 Iout.n298 Iout.n170 0.451012
R15465 Iout.n299 Iout.n298 0.451012
R15466 Iout.n299 Iout.n166 0.451012
R15467 Iout.n381 Iout.n166 0.451012
R15468 Iout.n382 Iout.n381 0.451012
R15469 Iout.n382 Iout.n83 0.451012
R15470 Iout.n645 Iout.n83 0.451012
R15471 Iout.n646 Iout.n645 0.451012
R15472 Iout.n646 Iout.n40 0.451012
R15473 Iout.n774 Iout.n40 0.451012
R15474 Iout.n775 Iout.n774 0.451012
R15475 Iout.n775 Iout.n36 0.451012
R15476 Iout.n837 Iout.n36 0.451012
R15477 Iout.n1018 Iout.n1017 0.451012
R15478 Iout.n1017 Iout.n0 0.451012
R15479 Iout.n999 Iout.n0 0.451012
R15480 Iout.n999 Iout.n998 0.451012
R15481 Iout.n998 Iout.n6 0.451012
R15482 Iout.n980 Iout.n6 0.451012
R15483 Iout.n980 Iout.n979 0.451012
R15484 Iout.n979 Iout.n11 0.451012
R15485 Iout.n961 Iout.n11 0.451012
R15486 Iout.n961 Iout.n960 0.451012
R15487 Iout.n960 Iout.n16 0.451012
R15488 Iout.n942 Iout.n16 0.451012
R15489 Iout.n942 Iout.n941 0.451012
R15490 Iout.n941 Iout.n21 0.451012
R15491 Iout.n230 Iout.n229 0.451012
R15492 Iout.n230 Iout.n167 0.451012
R15493 Iout.n304 Iout.n167 0.451012
R15494 Iout.n332 Iout.n304 0.451012
R15495 Iout.n374 Iout.n332 0.451012
R15496 Iout.n374 Iout.n373 0.451012
R15497 Iout.n373 Iout.n369 0.451012
R15498 Iout.n369 Iout.n80 0.451012
R15499 Iout.n651 Iout.n80 0.451012
R15500 Iout.n652 Iout.n651 0.451012
R15501 Iout.n652 Iout.n37 0.451012
R15502 Iout.n780 Iout.n37 0.451012
R15503 Iout.n826 Iout.n780 0.451012
R15504 Iout.n830 Iout.n826 0.451012
R15505 Iout.n231 Iout 0.2919
R15506 Iout.n303 Iout 0.2919
R15507 Iout Iout.n300 0.2919
R15508 Iout.n375 Iout 0.2919
R15509 Iout.n380 Iout 0.2919
R15510 Iout.n391 Iout 0.2919
R15511 Iout.n368 Iout 0.2919
R15512 Iout Iout.n365 0.2919
R15513 Iout Iout.n362 0.2919
R15514 Iout Iout.n359 0.2919
R15515 Iout.n650 Iout 0.2919
R15516 Iout Iout.n647 0.2919
R15517 Iout.n638 Iout 0.2919
R15518 Iout Iout.n635 0.2919
R15519 Iout.n626 Iout 0.2919
R15520 Iout.n41 Iout 0.2919
R15521 Iout.n773 Iout 0.2919
R15522 Iout Iout.n770 0.2919
R15523 Iout.n761 Iout 0.2919
R15524 Iout Iout.n758 0.2919
R15525 Iout.n749 Iout 0.2919
R15526 Iout.n825 Iout 0.2919
R15527 Iout Iout.n822 0.2919
R15528 Iout Iout.n819 0.2919
R15529 Iout Iout.n816 0.2919
R15530 Iout Iout.n813 0.2919
R15531 Iout Iout.n810 0.2919
R15532 Iout Iout.n807 0.2919
R15533 Iout.n829 Iout 0.2919
R15534 Iout.n838 Iout 0.2919
R15535 Iout.n843 Iout 0.2919
R15536 Iout.n852 Iout 0.2919
R15537 Iout.n857 Iout 0.2919
R15538 Iout.n866 Iout 0.2919
R15539 Iout.n871 Iout 0.2919
R15540 Iout.n880 Iout 0.2919
R15541 Iout Iout.n925 0.2919
R15542 Iout.n928 Iout 0.2919
R15543 Iout.n922 Iout 0.2919
R15544 Iout.n913 Iout 0.2919
R15545 Iout.n908 Iout 0.2919
R15546 Iout.n899 Iout 0.2919
R15547 Iout.n894 Iout 0.2919
R15548 Iout.n885 Iout 0.2919
R15549 Iout.n831 Iout 0.2919
R15550 Iout.n836 Iout 0.2919
R15551 Iout.n845 Iout 0.2919
R15552 Iout.n850 Iout 0.2919
R15553 Iout.n859 Iout 0.2919
R15554 Iout.n864 Iout 0.2919
R15555 Iout.n873 Iout 0.2919
R15556 Iout.n878 Iout 0.2919
R15557 Iout.n887 Iout 0.2919
R15558 Iout.n892 Iout 0.2919
R15559 Iout.n933 Iout 0.2919
R15560 Iout.n930 Iout 0.2919
R15561 Iout.n920 Iout 0.2919
R15562 Iout.n915 Iout 0.2919
R15563 Iout.n906 Iout 0.2919
R15564 Iout.n901 Iout 0.2919
R15565 Iout.n940 Iout 0.2919
R15566 Iout Iout.n783 0.2919
R15567 Iout Iout.n786 0.2919
R15568 Iout Iout.n789 0.2919
R15569 Iout Iout.n792 0.2919
R15570 Iout Iout.n795 0.2919
R15571 Iout Iout.n798 0.2919
R15572 Iout Iout.n801 0.2919
R15573 Iout Iout.n804 0.2919
R15574 Iout.n779 Iout 0.2919
R15575 Iout Iout.n776 0.2919
R15576 Iout.n767 Iout 0.2919
R15577 Iout Iout.n764 0.2919
R15578 Iout.n755 Iout 0.2919
R15579 Iout Iout.n752 0.2919
R15580 Iout.n743 Iout 0.2919
R15581 Iout Iout.n740 0.2919
R15582 Iout.n731 Iout 0.2919
R15583 Iout Iout.n728 0.2919
R15584 Iout.n719 Iout 0.2919
R15585 Iout Iout.n943 0.2919
R15586 Iout.n946 Iout 0.2919
R15587 Iout Iout.n704 0.2919
R15588 Iout.n707 Iout 0.2919
R15589 Iout Iout.n716 0.2919
R15590 Iout.n952 Iout 0.2919
R15591 Iout.n949 Iout 0.2919
R15592 Iout.n701 Iout 0.2919
R15593 Iout Iout.n710 0.2919
R15594 Iout.n713 Iout 0.2919
R15595 Iout Iout.n722 0.2919
R15596 Iout.n725 Iout 0.2919
R15597 Iout Iout.n734 0.2919
R15598 Iout.n737 Iout 0.2919
R15599 Iout Iout.n746 0.2919
R15600 Iout.n653 Iout 0.2919
R15601 Iout.n656 Iout 0.2919
R15602 Iout.n659 Iout 0.2919
R15603 Iout.n662 Iout 0.2919
R15604 Iout.n665 Iout 0.2919
R15605 Iout.n668 Iout 0.2919
R15606 Iout.n671 Iout 0.2919
R15607 Iout.n674 Iout 0.2919
R15608 Iout.n677 Iout 0.2919
R15609 Iout.n680 Iout 0.2919
R15610 Iout.n683 Iout 0.2919
R15611 Iout.n686 Iout 0.2919
R15612 Iout.n959 Iout 0.2919
R15613 Iout Iout.n694 0.2919
R15614 Iout.n697 Iout 0.2919
R15615 Iout.n689 Iout 0.2919
R15616 Iout Iout.n962 0.2919
R15617 Iout.n965 Iout 0.2919
R15618 Iout Iout.n575 0.2919
R15619 Iout.n578 Iout 0.2919
R15620 Iout Iout.n587 0.2919
R15621 Iout.n590 Iout 0.2919
R15622 Iout Iout.n599 0.2919
R15623 Iout.n602 Iout 0.2919
R15624 Iout Iout.n611 0.2919
R15625 Iout.n614 Iout 0.2919
R15626 Iout Iout.n623 0.2919
R15627 Iout.n84 Iout 0.2919
R15628 Iout.n644 Iout 0.2919
R15629 Iout Iout.n641 0.2919
R15630 Iout.n632 Iout 0.2919
R15631 Iout Iout.n629 0.2919
R15632 Iout.n620 Iout 0.2919
R15633 Iout Iout.n617 0.2919
R15634 Iout.n608 Iout 0.2919
R15635 Iout Iout.n605 0.2919
R15636 Iout.n596 Iout 0.2919
R15637 Iout Iout.n593 0.2919
R15638 Iout.n584 Iout 0.2919
R15639 Iout Iout.n581 0.2919
R15640 Iout.n971 Iout 0.2919
R15641 Iout.n968 Iout 0.2919
R15642 Iout.n565 Iout 0.2919
R15643 Iout.n978 Iout 0.2919
R15644 Iout Iout.n122 0.2919
R15645 Iout Iout.n568 0.2919
R15646 Iout.n571 Iout 0.2919
R15647 Iout Iout.n335 0.2919
R15648 Iout Iout.n338 0.2919
R15649 Iout Iout.n341 0.2919
R15650 Iout Iout.n344 0.2919
R15651 Iout Iout.n347 0.2919
R15652 Iout Iout.n350 0.2919
R15653 Iout Iout.n353 0.2919
R15654 Iout Iout.n356 0.2919
R15655 Iout.n372 Iout 0.2919
R15656 Iout.n383 Iout 0.2919
R15657 Iout.n388 Iout 0.2919
R15658 Iout.n399 Iout 0.2919
R15659 Iout.n404 Iout 0.2919
R15660 Iout.n415 Iout 0.2919
R15661 Iout.n420 Iout 0.2919
R15662 Iout.n431 Iout 0.2919
R15663 Iout.n443 Iout 0.2919
R15664 Iout Iout.n440 0.2919
R15665 Iout Iout.n437 0.2919
R15666 Iout.n553 Iout 0.2919
R15667 Iout.n556 Iout 0.2919
R15668 Iout.n561 Iout 0.2919
R15669 Iout Iout.n981 0.2919
R15670 Iout.n984 Iout 0.2919
R15671 Iout.n990 Iout 0.2919
R15672 Iout.n987 Iout 0.2919
R15673 Iout Iout.n129 0.2919
R15674 Iout Iout.n547 0.2919
R15675 Iout.n550 Iout 0.2919
R15676 Iout Iout.n451 0.2919
R15677 Iout.n454 Iout 0.2919
R15678 Iout.n446 Iout 0.2919
R15679 Iout.n428 Iout 0.2919
R15680 Iout.n423 Iout 0.2919
R15681 Iout.n412 Iout 0.2919
R15682 Iout.n407 Iout 0.2919
R15683 Iout.n396 Iout 0.2919
R15684 Iout.n331 Iout 0.2919
R15685 Iout Iout.n328 0.2919
R15686 Iout Iout.n325 0.2919
R15687 Iout Iout.n322 0.2919
R15688 Iout Iout.n319 0.2919
R15689 Iout Iout.n316 0.2919
R15690 Iout Iout.n313 0.2919
R15691 Iout Iout.n310 0.2919
R15692 Iout Iout.n307 0.2919
R15693 Iout.n457 Iout 0.2919
R15694 Iout.n465 Iout 0.2919
R15695 Iout Iout.n462 0.2919
R15696 Iout.n544 Iout 0.2919
R15697 Iout Iout.n541 0.2919
R15698 Iout Iout.n135 0.2919
R15699 Iout.n997 Iout 0.2919
R15700 Iout Iout.n1000 0.2919
R15701 Iout.n1003 Iout 0.2919
R15702 Iout.n538 Iout 0.2919
R15703 Iout.n533 Iout 0.2919
R15704 Iout.n530 Iout 0.2919
R15705 Iout Iout.n468 0.2919
R15706 Iout Iout.n471 0.2919
R15707 Iout.n474 Iout 0.2919
R15708 Iout Iout.n264 0.2919
R15709 Iout.n267 Iout 0.2919
R15710 Iout Iout.n276 0.2919
R15711 Iout.n279 Iout 0.2919
R15712 Iout Iout.n288 0.2919
R15713 Iout.n291 Iout 0.2919
R15714 Iout.n171 Iout 0.2919
R15715 Iout.n297 Iout 0.2919
R15716 Iout Iout.n294 0.2919
R15717 Iout.n285 Iout 0.2919
R15718 Iout Iout.n282 0.2919
R15719 Iout.n273 Iout 0.2919
R15720 Iout Iout.n270 0.2919
R15721 Iout.n261 Iout 0.2919
R15722 Iout.n477 Iout 0.2919
R15723 Iout.n485 Iout 0.2919
R15724 Iout Iout.n482 0.2919
R15725 Iout.n527 Iout 0.2919
R15726 Iout Iout.n524 0.2919
R15727 Iout Iout.n142 0.2919
R15728 Iout.n1006 Iout 0.2919
R15729 Iout.n1009 Iout 0.2919
R15730 Iout.n1016 Iout 0.2919
R15731 Iout Iout.n148 0.2919
R15732 Iout Iout.n518 0.2919
R15733 Iout.n521 Iout 0.2919
R15734 Iout Iout.n493 0.2919
R15735 Iout.n496 Iout 0.2919
R15736 Iout.n488 Iout 0.2919
R15737 Iout Iout.n254 0.2919
R15738 Iout.n257 Iout 0.2919
R15739 Iout.n249 Iout 0.2919
R15740 Iout.n246 Iout 0.2919
R15741 Iout.n243 Iout 0.2919
R15742 Iout.n240 Iout 0.2919
R15743 Iout.n237 Iout 0.2919
R15744 Iout.n234 Iout 0.2919
R15745 Iout.n228 Iout 0.2919
R15746 Iout Iout.n225 0.2919
R15747 Iout Iout.n221 0.2919
R15748 Iout Iout.n217 0.2919
R15749 Iout Iout.n213 0.2919
R15750 Iout Iout.n209 0.2919
R15751 Iout Iout.n205 0.2919
R15752 Iout Iout.n201 0.2919
R15753 Iout Iout.n198 0.2919
R15754 Iout Iout.n194 0.2919
R15755 Iout.n499 Iout 0.2919
R15756 Iout.n503 Iout 0.2919
R15757 Iout.n506 Iout 0.2919
R15758 Iout.n515 Iout 0.2919
R15759 Iout Iout.n512 0.2919
R15760 Iout.n1019 Iout 0.2919
R15761 Iout.n1013 Iout.n1012 0.092855
R15762 Iout.n1012 Iout.n1 0.092855
R15763 Iout.n994 Iout.n1 0.092855
R15764 Iout.n994 Iout.n993 0.092855
R15765 Iout.n993 Iout.n7 0.092855
R15766 Iout.n975 Iout.n7 0.092855
R15767 Iout.n975 Iout.n974 0.092855
R15768 Iout.n974 Iout.n12 0.092855
R15769 Iout.n956 Iout.n12 0.092855
R15770 Iout.n956 Iout.n955 0.092855
R15771 Iout.n955 Iout.n17 0.092855
R15772 Iout.n937 Iout.n17 0.092855
R15773 Iout.n937 Iout.n936 0.092855
R15774 Iout.n197 Iout 0.0818902
R15775 Iout.n191 Iout 0.0818902
R15776 Iout.n152 Iout 0.0818902
R15777 Iout.n204 Iout 0.0818902
R15778 Iout.n498 Iout 0.0818902
R15779 Iout.n208 Iout 0.0818902
R15780 Iout.n502 Iout 0.0818902
R15781 Iout.n212 Iout 0.0818902
R15782 Iout.n145 Iout 0.0818902
R15783 Iout.n216 Iout 0.0818902
R15784 Iout.n516 Iout 0.0818902
R15785 Iout.n220 Iout 0.0818902
R15786 Iout.n511 Iout 0.0818902
R15787 Iout.n224 Iout 0.0818902
R15788 Iout.n1018 Iout 0.0818902
R15789 Iout.n229 Iout 0.0818902
R15790 Iout.n1013 Iout 0.072645
R15791 Iout.n302 Iout 0.0532071
R15792 Iout Iout.n377 0.0532071
R15793 Iout.n379 Iout 0.0532071
R15794 Iout.n367 Iout 0.0532071
R15795 Iout.n364 Iout 0.0532071
R15796 Iout.n361 Iout 0.0532071
R15797 Iout.n649 Iout 0.0532071
R15798 Iout Iout.n82 0.0532071
R15799 Iout.n637 Iout 0.0532071
R15800 Iout Iout.n91 0.0532071
R15801 Iout Iout.n43 0.0532071
R15802 Iout.n772 Iout 0.0532071
R15803 Iout Iout.n45 0.0532071
R15804 Iout.n760 Iout 0.0532071
R15805 Iout Iout.n51 0.0532071
R15806 Iout.n824 Iout 0.0532071
R15807 Iout.n821 Iout 0.0532071
R15808 Iout.n818 Iout 0.0532071
R15809 Iout.n815 Iout 0.0532071
R15810 Iout.n812 Iout 0.0532071
R15811 Iout.n809 Iout 0.0532071
R15812 Iout.n828 Iout 0.0532071
R15813 Iout Iout.n840 0.0532071
R15814 Iout.n842 Iout 0.0532071
R15815 Iout Iout.n854 0.0532071
R15816 Iout.n856 Iout 0.0532071
R15817 Iout Iout.n868 0.0532071
R15818 Iout.n870 Iout 0.0532071
R15819 Iout.n927 Iout 0.0532071
R15820 Iout Iout.n924 0.0532071
R15821 Iout.n912 Iout 0.0532071
R15822 Iout Iout.n910 0.0532071
R15823 Iout.n898 Iout 0.0532071
R15824 Iout Iout.n896 0.0532071
R15825 Iout.n884 Iout 0.0532071
R15826 Iout Iout.n882 0.0532071
R15827 Iout Iout.n833 0.0532071
R15828 Iout.n835 Iout 0.0532071
R15829 Iout Iout.n847 0.0532071
R15830 Iout.n849 Iout 0.0532071
R15831 Iout Iout.n861 0.0532071
R15832 Iout.n863 Iout 0.0532071
R15833 Iout Iout.n875 0.0532071
R15834 Iout.n877 Iout 0.0532071
R15835 Iout Iout.n889 0.0532071
R15836 Iout Iout.n932 0.0532071
R15837 Iout.n919 Iout 0.0532071
R15838 Iout Iout.n917 0.0532071
R15839 Iout.n905 Iout 0.0532071
R15840 Iout Iout.n903 0.0532071
R15841 Iout.n891 Iout 0.0532071
R15842 Iout.n782 Iout 0.0532071
R15843 Iout.n785 Iout 0.0532071
R15844 Iout.n788 Iout 0.0532071
R15845 Iout.n791 Iout 0.0532071
R15846 Iout.n794 Iout 0.0532071
R15847 Iout.n797 Iout 0.0532071
R15848 Iout.n800 Iout 0.0532071
R15849 Iout.n803 Iout 0.0532071
R15850 Iout.n806 Iout 0.0532071
R15851 Iout.n778 Iout 0.0532071
R15852 Iout Iout.n39 0.0532071
R15853 Iout.n766 Iout 0.0532071
R15854 Iout Iout.n48 0.0532071
R15855 Iout.n754 Iout 0.0532071
R15856 Iout Iout.n54 0.0532071
R15857 Iout.n742 Iout 0.0532071
R15858 Iout Iout.n60 0.0532071
R15859 Iout.n730 Iout 0.0532071
R15860 Iout Iout.n66 0.0532071
R15861 Iout.n945 Iout 0.0532071
R15862 Iout.n78 Iout 0.0532071
R15863 Iout.n706 Iout 0.0532071
R15864 Iout Iout.n72 0.0532071
R15865 Iout.n718 Iout 0.0532071
R15866 Iout Iout.n951 0.0532071
R15867 Iout.n700 Iout 0.0532071
R15868 Iout Iout.n75 0.0532071
R15869 Iout.n712 Iout 0.0532071
R15870 Iout Iout.n69 0.0532071
R15871 Iout.n724 Iout 0.0532071
R15872 Iout Iout.n63 0.0532071
R15873 Iout.n736 Iout 0.0532071
R15874 Iout Iout.n57 0.0532071
R15875 Iout.n748 Iout 0.0532071
R15876 Iout Iout.n655 0.0532071
R15877 Iout Iout.n658 0.0532071
R15878 Iout Iout.n661 0.0532071
R15879 Iout Iout.n664 0.0532071
R15880 Iout Iout.n667 0.0532071
R15881 Iout Iout.n670 0.0532071
R15882 Iout Iout.n673 0.0532071
R15883 Iout Iout.n676 0.0532071
R15884 Iout Iout.n679 0.0532071
R15885 Iout Iout.n682 0.0532071
R15886 Iout Iout.n685 0.0532071
R15887 Iout.n693 Iout 0.0532071
R15888 Iout.n696 Iout 0.0532071
R15889 Iout Iout.n691 0.0532071
R15890 Iout Iout.n688 0.0532071
R15891 Iout.n964 Iout 0.0532071
R15892 Iout.n574 Iout 0.0532071
R15893 Iout.n577 Iout 0.0532071
R15894 Iout Iout.n115 0.0532071
R15895 Iout.n589 Iout 0.0532071
R15896 Iout Iout.n109 0.0532071
R15897 Iout.n601 Iout 0.0532071
R15898 Iout Iout.n103 0.0532071
R15899 Iout.n613 Iout 0.0532071
R15900 Iout Iout.n97 0.0532071
R15901 Iout.n625 Iout 0.0532071
R15902 Iout Iout.n86 0.0532071
R15903 Iout.n643 Iout 0.0532071
R15904 Iout Iout.n88 0.0532071
R15905 Iout.n631 Iout 0.0532071
R15906 Iout Iout.n94 0.0532071
R15907 Iout.n619 Iout 0.0532071
R15908 Iout Iout.n100 0.0532071
R15909 Iout.n607 Iout 0.0532071
R15910 Iout Iout.n106 0.0532071
R15911 Iout.n595 Iout 0.0532071
R15912 Iout Iout.n112 0.0532071
R15913 Iout.n583 Iout 0.0532071
R15914 Iout Iout.n970 0.0532071
R15915 Iout.n564 Iout 0.0532071
R15916 Iout Iout.n118 0.0532071
R15917 Iout.n121 Iout 0.0532071
R15918 Iout.n124 Iout 0.0532071
R15919 Iout.n570 Iout 0.0532071
R15920 Iout.n334 Iout 0.0532071
R15921 Iout.n337 Iout 0.0532071
R15922 Iout.n340 Iout 0.0532071
R15923 Iout.n343 Iout 0.0532071
R15924 Iout.n346 Iout 0.0532071
R15925 Iout.n349 Iout 0.0532071
R15926 Iout.n352 Iout 0.0532071
R15927 Iout.n355 Iout 0.0532071
R15928 Iout.n358 Iout 0.0532071
R15929 Iout.n371 Iout 0.0532071
R15930 Iout Iout.n385 0.0532071
R15931 Iout.n387 Iout 0.0532071
R15932 Iout Iout.n401 0.0532071
R15933 Iout.n403 Iout 0.0532071
R15934 Iout Iout.n417 0.0532071
R15935 Iout.n419 Iout 0.0532071
R15936 Iout Iout.n433 0.0532071
R15937 Iout.n442 Iout 0.0532071
R15938 Iout.n439 Iout 0.0532071
R15939 Iout.n435 Iout 0.0532071
R15940 Iout Iout.n555 0.0532071
R15941 Iout Iout.n558 0.0532071
R15942 Iout.n983 Iout 0.0532071
R15943 Iout.n560 Iout 0.0532071
R15944 Iout Iout.n989 0.0532071
R15945 Iout.n128 Iout 0.0532071
R15946 Iout.n131 Iout 0.0532071
R15947 Iout.n549 Iout 0.0532071
R15948 Iout.n450 Iout 0.0532071
R15949 Iout.n453 Iout 0.0532071
R15950 Iout Iout.n448 0.0532071
R15951 Iout.n427 Iout 0.0532071
R15952 Iout Iout.n425 0.0532071
R15953 Iout.n411 Iout 0.0532071
R15954 Iout Iout.n409 0.0532071
R15955 Iout.n395 Iout 0.0532071
R15956 Iout Iout.n393 0.0532071
R15957 Iout.n330 Iout 0.0532071
R15958 Iout.n327 Iout 0.0532071
R15959 Iout.n324 Iout 0.0532071
R15960 Iout.n321 Iout 0.0532071
R15961 Iout.n318 Iout 0.0532071
R15962 Iout.n315 Iout 0.0532071
R15963 Iout.n312 Iout 0.0532071
R15964 Iout.n309 Iout 0.0532071
R15965 Iout.n306 Iout 0.0532071
R15966 Iout Iout.n459 0.0532071
R15967 Iout.n464 Iout 0.0532071
R15968 Iout.n461 Iout 0.0532071
R15969 Iout.n543 Iout 0.0532071
R15970 Iout.n137 Iout 0.0532071
R15971 Iout.n134 Iout 0.0532071
R15972 Iout.n1002 Iout 0.0532071
R15973 Iout.n537 Iout 0.0532071
R15974 Iout Iout.n535 0.0532071
R15975 Iout Iout.n532 0.0532071
R15976 Iout.n157 Iout 0.0532071
R15977 Iout.n470 Iout 0.0532071
R15978 Iout.n473 Iout 0.0532071
R15979 Iout.n190 Iout 0.0532071
R15980 Iout.n266 Iout 0.0532071
R15981 Iout Iout.n184 0.0532071
R15982 Iout.n278 Iout 0.0532071
R15983 Iout Iout.n178 0.0532071
R15984 Iout.n290 Iout 0.0532071
R15985 Iout Iout.n169 0.0532071
R15986 Iout Iout.n173 0.0532071
R15987 Iout.n296 Iout 0.0532071
R15988 Iout Iout.n175 0.0532071
R15989 Iout.n284 Iout 0.0532071
R15990 Iout Iout.n181 0.0532071
R15991 Iout.n272 Iout 0.0532071
R15992 Iout Iout.n187 0.0532071
R15993 Iout.n260 Iout 0.0532071
R15994 Iout Iout.n479 0.0532071
R15995 Iout.n484 Iout 0.0532071
R15996 Iout.n481 Iout 0.0532071
R15997 Iout.n526 Iout 0.0532071
R15998 Iout.n144 Iout 0.0532071
R15999 Iout.n141 Iout 0.0532071
R16000 Iout Iout.n1008 0.0532071
R16001 Iout.n147 Iout 0.0532071
R16002 Iout.n150 Iout 0.0532071
R16003 Iout.n520 Iout 0.0532071
R16004 Iout.n492 Iout 0.0532071
R16005 Iout.n495 Iout 0.0532071
R16006 Iout Iout.n490 0.0532071
R16007 Iout.n253 Iout 0.0532071
R16008 Iout.n256 Iout 0.0532071
R16009 Iout Iout.n251 0.0532071
R16010 Iout Iout.n248 0.0532071
R16011 Iout Iout.n245 0.0532071
R16012 Iout Iout.n242 0.0532071
R16013 Iout Iout.n239 0.0532071
R16014 Iout Iout.n236 0.0532071
R16015 Iout Iout.n233 0.0532071
R16016 Iout.n227 Iout 0.0532071
R16017 Iout.n223 Iout 0.0532071
R16018 Iout.n219 Iout 0.0532071
R16019 Iout.n215 Iout 0.0532071
R16020 Iout.n211 Iout 0.0532071
R16021 Iout.n207 Iout 0.0532071
R16022 Iout.n203 Iout 0.0532071
R16023 Iout.n200 Iout 0.0532071
R16024 Iout.n196 Iout 0.0532071
R16025 Iout.n193 Iout 0.0532071
R16026 Iout Iout.n501 0.0532071
R16027 Iout Iout.n505 0.0532071
R16028 Iout Iout.n508 0.0532071
R16029 Iout.n514 Iout 0.0532071
R16030 Iout.n510 Iout 0.0532071
R16031 Iout.n1020 Iout 0.03925
R16032 Iout.n509 Iout 0.03925
R16033 Iout.n513 Iout 0.03925
R16034 Iout.n507 Iout 0.03925
R16035 Iout.n504 Iout 0.03925
R16036 Iout.n500 Iout 0.03925
R16037 Iout.n192 Iout 0.03925
R16038 Iout.n195 Iout 0.03925
R16039 Iout.n199 Iout 0.03925
R16040 Iout.n202 Iout 0.03925
R16041 Iout.n206 Iout 0.03925
R16042 Iout.n210 Iout 0.03925
R16043 Iout.n214 Iout 0.03925
R16044 Iout.n218 Iout 0.03925
R16045 Iout.n222 Iout 0.03925
R16046 Iout.n226 Iout 0.03925
R16047 Iout.n232 Iout 0.03925
R16048 Iout.n235 Iout 0.03925
R16049 Iout.n238 Iout 0.03925
R16050 Iout.n241 Iout 0.03925
R16051 Iout.n244 Iout 0.03925
R16052 Iout.n247 Iout 0.03925
R16053 Iout.n250 Iout 0.03925
R16054 Iout.n255 Iout 0.03925
R16055 Iout.n252 Iout 0.03925
R16056 Iout.n489 Iout 0.03925
R16057 Iout.n494 Iout 0.03925
R16058 Iout.n491 Iout 0.03925
R16059 Iout.n519 Iout 0.03925
R16060 Iout.n149 Iout 0.03925
R16061 Iout.n146 Iout 0.03925
R16062 Iout.n1010 Iout 0.03925
R16063 Iout.n1007 Iout 0.03925
R16064 Iout.n140 Iout 0.03925
R16065 Iout.n143 Iout 0.03925
R16066 Iout.n525 Iout 0.03925
R16067 Iout.n480 Iout 0.03925
R16068 Iout.n483 Iout 0.03925
R16069 Iout.n478 Iout 0.03925
R16070 Iout.n259 Iout 0.03925
R16071 Iout.n186 Iout 0.03925
R16072 Iout.n271 Iout 0.03925
R16073 Iout.n180 Iout 0.03925
R16074 Iout.n283 Iout 0.03925
R16075 Iout.n174 Iout 0.03925
R16076 Iout.n168 Iout 0.03925
R16077 Iout.n301 Iout 0.03925
R16078 Iout.n289 Iout 0.03925
R16079 Iout.n177 Iout 0.03925
R16080 Iout.n277 Iout 0.03925
R16081 Iout.n183 Iout 0.03925
R16082 Iout.n265 Iout 0.03925
R16083 Iout.n189 Iout 0.03925
R16084 Iout.n472 Iout 0.03925
R16085 Iout.n469 Iout 0.03925
R16086 Iout.n156 Iout 0.03925
R16087 Iout.n531 Iout 0.03925
R16088 Iout.n534 Iout 0.03925
R16089 Iout.n536 Iout 0.03925
R16090 Iout.n133 Iout 0.03925
R16091 Iout.n136 Iout 0.03925
R16092 Iout.n542 Iout 0.03925
R16093 Iout.n460 Iout 0.03925
R16094 Iout.n463 Iout 0.03925
R16095 Iout.n458 Iout 0.03925
R16096 Iout.n305 Iout 0.03925
R16097 Iout.n308 Iout 0.03925
R16098 Iout.n311 Iout 0.03925
R16099 Iout.n314 Iout 0.03925
R16100 Iout.n317 Iout 0.03925
R16101 Iout.n320 Iout 0.03925
R16102 Iout.n392 Iout 0.03925
R16103 Iout.n378 Iout 0.03925
R16104 Iout.n376 Iout 0.03925
R16105 Iout.n394 Iout 0.03925
R16106 Iout.n408 Iout 0.03925
R16107 Iout.n410 Iout 0.03925
R16108 Iout.n424 Iout 0.03925
R16109 Iout.n426 Iout 0.03925
R16110 Iout.n447 Iout 0.03925
R16111 Iout.n452 Iout 0.03925
R16112 Iout.n449 Iout 0.03925
R16113 Iout.n548 Iout 0.03925
R16114 Iout.n130 Iout 0.03925
R16115 Iout.n559 Iout 0.03925
R16116 Iout.n557 Iout 0.03925
R16117 Iout.n554 Iout 0.03925
R16118 Iout.n434 Iout 0.03925
R16119 Iout.n438 Iout 0.03925
R16120 Iout.n441 Iout 0.03925
R16121 Iout.n432 Iout 0.03925
R16122 Iout.n418 Iout 0.03925
R16123 Iout.n416 Iout 0.03925
R16124 Iout.n402 Iout 0.03925
R16125 Iout.n357 Iout 0.03925
R16126 Iout.n360 Iout 0.03925
R16127 Iout.n363 Iout 0.03925
R16128 Iout.n366 Iout 0.03925
R16129 Iout.n354 Iout 0.03925
R16130 Iout.n351 Iout 0.03925
R16131 Iout.n348 Iout 0.03925
R16132 Iout.n345 Iout 0.03925
R16133 Iout.n342 Iout 0.03925
R16134 Iout.n339 Iout 0.03925
R16135 Iout.n336 Iout 0.03925
R16136 Iout.n333 Iout 0.03925
R16137 Iout.n117 Iout 0.03925
R16138 Iout.n582 Iout 0.03925
R16139 Iout.n111 Iout 0.03925
R16140 Iout.n594 Iout 0.03925
R16141 Iout.n105 Iout 0.03925
R16142 Iout.n606 Iout 0.03925
R16143 Iout.n99 Iout 0.03925
R16144 Iout.n618 Iout 0.03925
R16145 Iout.n624 Iout 0.03925
R16146 Iout.n90 Iout 0.03925
R16147 Iout.n636 Iout 0.03925
R16148 Iout.n81 Iout 0.03925
R16149 Iout.n648 Iout 0.03925
R16150 Iout.n96 Iout 0.03925
R16151 Iout.n612 Iout 0.03925
R16152 Iout.n102 Iout 0.03925
R16153 Iout.n600 Iout 0.03925
R16154 Iout.n108 Iout 0.03925
R16155 Iout.n588 Iout 0.03925
R16156 Iout.n687 Iout 0.03925
R16157 Iout.n684 Iout 0.03925
R16158 Iout.n681 Iout 0.03925
R16159 Iout.n678 Iout 0.03925
R16160 Iout.n675 Iout 0.03925
R16161 Iout.n672 Iout 0.03925
R16162 Iout.n747 Iout 0.03925
R16163 Iout.n50 Iout 0.03925
R16164 Iout.n759 Iout 0.03925
R16165 Iout.n44 Iout 0.03925
R16166 Iout.n771 Iout 0.03925
R16167 Iout.n42 Iout 0.03925
R16168 Iout.n56 Iout 0.03925
R16169 Iout.n735 Iout 0.03925
R16170 Iout.n62 Iout 0.03925
R16171 Iout.n723 Iout 0.03925
R16172 Iout.n717 Iout 0.03925
R16173 Iout.n65 Iout 0.03925
R16174 Iout.n729 Iout 0.03925
R16175 Iout.n59 Iout 0.03925
R16176 Iout.n805 Iout 0.03925
R16177 Iout.n808 Iout 0.03925
R16178 Iout.n811 Iout 0.03925
R16179 Iout.n814 Iout 0.03925
R16180 Iout.n817 Iout 0.03925
R16181 Iout.n820 Iout 0.03925
R16182 Iout.n823 Iout 0.03925
R16183 Iout.n802 Iout 0.03925
R16184 Iout.n799 Iout 0.03925
R16185 Iout.n890 Iout 0.03925
R16186 Iout.n888 Iout 0.03925
R16187 Iout.n881 Iout 0.03925
R16188 Iout.n869 Iout 0.03925
R16189 Iout.n867 Iout 0.03925
R16190 Iout.n855 Iout 0.03925
R16191 Iout.n853 Iout 0.03925
R16192 Iout.n841 Iout 0.03925
R16193 Iout.n839 Iout 0.03925
R16194 Iout.n827 Iout 0.03925
R16195 Iout.n883 Iout 0.03925
R16196 Iout.n895 Iout 0.03925
R16197 Iout.n897 Iout 0.03925
R16198 Iout.n909 Iout 0.03925
R16199 Iout.n911 Iout 0.03925
R16200 Iout.n923 Iout 0.03925
R16201 Iout.n926 Iout 0.03925
R16202 Iout.n22 Iout 0.03925
R16203 Iout.n876 Iout 0.03925
R16204 Iout.n874 Iout 0.03925
R16205 Iout.n862 Iout 0.03925
R16206 Iout.n860 Iout 0.03925
R16207 Iout.n848 Iout 0.03925
R16208 Iout.n846 Iout 0.03925
R16209 Iout.n834 Iout 0.03925
R16210 Iout.n832 Iout 0.03925
R16211 Iout.n902 Iout 0.03925
R16212 Iout.n904 Iout 0.03925
R16213 Iout.n916 Iout 0.03925
R16214 Iout.n918 Iout 0.03925
R16215 Iout.n931 Iout 0.03925
R16216 Iout.n934 Iout 0.03925
R16217 Iout.n796 Iout 0.03925
R16218 Iout.n793 Iout 0.03925
R16219 Iout.n790 Iout 0.03925
R16220 Iout.n787 Iout 0.03925
R16221 Iout.n784 Iout 0.03925
R16222 Iout.n781 Iout 0.03925
R16223 Iout.n938 Iout 0.03925
R16224 Iout.n741 Iout 0.03925
R16225 Iout.n53 Iout 0.03925
R16226 Iout.n753 Iout 0.03925
R16227 Iout.n47 Iout 0.03925
R16228 Iout.n765 Iout 0.03925
R16229 Iout.n38 Iout 0.03925
R16230 Iout.n777 Iout 0.03925
R16231 Iout.n71 Iout 0.03925
R16232 Iout.n705 Iout 0.03925
R16233 Iout.n77 Iout 0.03925
R16234 Iout.n944 Iout 0.03925
R16235 Iout.n19 Iout 0.03925
R16236 Iout.n68 Iout 0.03925
R16237 Iout.n711 Iout 0.03925
R16238 Iout.n74 Iout 0.03925
R16239 Iout.n699 Iout 0.03925
R16240 Iout.n950 Iout 0.03925
R16241 Iout.n953 Iout 0.03925
R16242 Iout.n669 Iout 0.03925
R16243 Iout.n666 Iout 0.03925
R16244 Iout.n663 Iout 0.03925
R16245 Iout.n660 Iout 0.03925
R16246 Iout.n657 Iout 0.03925
R16247 Iout.n654 Iout 0.03925
R16248 Iout.n690 Iout 0.03925
R16249 Iout.n695 Iout 0.03925
R16250 Iout.n692 Iout 0.03925
R16251 Iout.n957 Iout 0.03925
R16252 Iout.n114 Iout 0.03925
R16253 Iout.n576 Iout 0.03925
R16254 Iout.n573 Iout 0.03925
R16255 Iout.n963 Iout 0.03925
R16256 Iout.n14 Iout 0.03925
R16257 Iout.n93 Iout 0.03925
R16258 Iout.n630 Iout 0.03925
R16259 Iout.n87 Iout 0.03925
R16260 Iout.n642 Iout 0.03925
R16261 Iout.n85 Iout 0.03925
R16262 Iout.n563 Iout 0.03925
R16263 Iout.n969 Iout 0.03925
R16264 Iout.n972 Iout 0.03925
R16265 Iout.n569 Iout 0.03925
R16266 Iout.n123 Iout 0.03925
R16267 Iout.n120 Iout 0.03925
R16268 Iout.n976 Iout 0.03925
R16269 Iout.n400 Iout 0.03925
R16270 Iout.n386 Iout 0.03925
R16271 Iout.n384 Iout 0.03925
R16272 Iout.n370 Iout 0.03925
R16273 Iout.n982 Iout 0.03925
R16274 Iout.n9 Iout 0.03925
R16275 Iout.n127 Iout 0.03925
R16276 Iout.n988 Iout 0.03925
R16277 Iout.n991 Iout 0.03925
R16278 Iout.n323 Iout 0.03925
R16279 Iout.n326 Iout 0.03925
R16280 Iout.n329 Iout 0.03925
R16281 Iout.n995 Iout 0.03925
R16282 Iout.n1001 Iout 0.03925
R16283 Iout.n4 Iout 0.03925
R16284 Iout.n295 Iout 0.03925
R16285 Iout.n172 Iout 0.03925
R16286 Iout.n1014 Iout 0.03925
R16287 Iout.n1022 Iout 0.02071
R16288 Iout Iout.n1022 0.00379
R16289 Iout.n303 Iout.n302 0.00105952
R16290 Iout.n377 Iout.n375 0.00105952
R16291 Iout.n380 Iout.n379 0.00105952
R16292 Iout.n368 Iout.n367 0.00105952
R16293 Iout.n365 Iout.n364 0.00105952
R16294 Iout.n362 Iout.n361 0.00105952
R16295 Iout.n650 Iout.n649 0.00105952
R16296 Iout.n647 Iout.n82 0.00105952
R16297 Iout.n638 Iout.n637 0.00105952
R16298 Iout.n635 Iout.n91 0.00105952
R16299 Iout.n43 Iout.n41 0.00105952
R16300 Iout.n773 Iout.n772 0.00105952
R16301 Iout.n770 Iout.n45 0.00105952
R16302 Iout.n761 Iout.n760 0.00105952
R16303 Iout.n758 Iout.n51 0.00105952
R16304 Iout.n825 Iout.n824 0.00105952
R16305 Iout.n822 Iout.n821 0.00105952
R16306 Iout.n819 Iout.n818 0.00105952
R16307 Iout.n816 Iout.n815 0.00105952
R16308 Iout.n813 Iout.n812 0.00105952
R16309 Iout.n810 Iout.n809 0.00105952
R16310 Iout.n829 Iout.n828 0.00105952
R16311 Iout.n840 Iout.n838 0.00105952
R16312 Iout.n843 Iout.n842 0.00105952
R16313 Iout.n854 Iout.n852 0.00105952
R16314 Iout.n857 Iout.n856 0.00105952
R16315 Iout.n868 Iout.n866 0.00105952
R16316 Iout.n871 Iout.n870 0.00105952
R16317 Iout.n925 Iout.n23 0.00105952
R16318 Iout.n928 Iout.n927 0.00105952
R16319 Iout.n924 Iout.n922 0.00105952
R16320 Iout.n913 Iout.n912 0.00105952
R16321 Iout.n910 Iout.n908 0.00105952
R16322 Iout.n899 Iout.n898 0.00105952
R16323 Iout.n896 Iout.n894 0.00105952
R16324 Iout.n885 Iout.n884 0.00105952
R16325 Iout.n882 Iout.n880 0.00105952
R16326 Iout.n833 Iout.n831 0.00105952
R16327 Iout.n836 Iout.n835 0.00105952
R16328 Iout.n847 Iout.n845 0.00105952
R16329 Iout.n850 Iout.n849 0.00105952
R16330 Iout.n861 Iout.n859 0.00105952
R16331 Iout.n864 Iout.n863 0.00105952
R16332 Iout.n875 Iout.n873 0.00105952
R16333 Iout.n878 Iout.n877 0.00105952
R16334 Iout.n889 Iout.n887 0.00105952
R16335 Iout.n935 Iout.n933 0.00105952
R16336 Iout.n932 Iout.n930 0.00105952
R16337 Iout.n920 Iout.n919 0.00105952
R16338 Iout.n917 Iout.n915 0.00105952
R16339 Iout.n906 Iout.n905 0.00105952
R16340 Iout.n903 Iout.n901 0.00105952
R16341 Iout.n892 Iout.n891 0.00105952
R16342 Iout.n940 Iout.n939 0.00105952
R16343 Iout.n783 Iout.n782 0.00105952
R16344 Iout.n786 Iout.n785 0.00105952
R16345 Iout.n789 Iout.n788 0.00105952
R16346 Iout.n792 Iout.n791 0.00105952
R16347 Iout.n795 Iout.n794 0.00105952
R16348 Iout.n798 Iout.n797 0.00105952
R16349 Iout.n801 Iout.n800 0.00105952
R16350 Iout.n804 Iout.n803 0.00105952
R16351 Iout.n807 Iout.n806 0.00105952
R16352 Iout.n779 Iout.n778 0.00105952
R16353 Iout.n776 Iout.n39 0.00105952
R16354 Iout.n767 Iout.n766 0.00105952
R16355 Iout.n764 Iout.n48 0.00105952
R16356 Iout.n755 Iout.n754 0.00105952
R16357 Iout.n752 Iout.n54 0.00105952
R16358 Iout.n743 Iout.n742 0.00105952
R16359 Iout.n740 Iout.n60 0.00105952
R16360 Iout.n731 Iout.n730 0.00105952
R16361 Iout.n728 Iout.n66 0.00105952
R16362 Iout.n943 Iout.n20 0.00105952
R16363 Iout.n946 Iout.n945 0.00105952
R16364 Iout.n704 Iout.n78 0.00105952
R16365 Iout.n707 Iout.n706 0.00105952
R16366 Iout.n716 Iout.n72 0.00105952
R16367 Iout.n719 Iout.n718 0.00105952
R16368 Iout.n954 Iout.n952 0.00105952
R16369 Iout.n951 Iout.n949 0.00105952
R16370 Iout.n701 Iout.n700 0.00105952
R16371 Iout.n710 Iout.n75 0.00105952
R16372 Iout.n713 Iout.n712 0.00105952
R16373 Iout.n722 Iout.n69 0.00105952
R16374 Iout.n725 Iout.n724 0.00105952
R16375 Iout.n734 Iout.n63 0.00105952
R16376 Iout.n737 Iout.n736 0.00105952
R16377 Iout.n746 Iout.n57 0.00105952
R16378 Iout.n749 Iout.n748 0.00105952
R16379 Iout.n655 Iout.n653 0.00105952
R16380 Iout.n658 Iout.n656 0.00105952
R16381 Iout.n661 Iout.n659 0.00105952
R16382 Iout.n664 Iout.n662 0.00105952
R16383 Iout.n667 Iout.n665 0.00105952
R16384 Iout.n670 Iout.n668 0.00105952
R16385 Iout.n673 Iout.n671 0.00105952
R16386 Iout.n676 Iout.n674 0.00105952
R16387 Iout.n679 Iout.n677 0.00105952
R16388 Iout.n682 Iout.n680 0.00105952
R16389 Iout.n685 Iout.n683 0.00105952
R16390 Iout.n959 Iout.n958 0.00105952
R16391 Iout.n694 Iout.n693 0.00105952
R16392 Iout.n697 Iout.n696 0.00105952
R16393 Iout.n691 Iout.n689 0.00105952
R16394 Iout.n688 Iout.n686 0.00105952
R16395 Iout.n962 Iout.n15 0.00105952
R16396 Iout.n965 Iout.n964 0.00105952
R16397 Iout.n575 Iout.n574 0.00105952
R16398 Iout.n578 Iout.n577 0.00105952
R16399 Iout.n587 Iout.n115 0.00105952
R16400 Iout.n590 Iout.n589 0.00105952
R16401 Iout.n599 Iout.n109 0.00105952
R16402 Iout.n602 Iout.n601 0.00105952
R16403 Iout.n611 Iout.n103 0.00105952
R16404 Iout.n614 Iout.n613 0.00105952
R16405 Iout.n623 Iout.n97 0.00105952
R16406 Iout.n626 Iout.n625 0.00105952
R16407 Iout.n86 Iout.n84 0.00105952
R16408 Iout.n644 Iout.n643 0.00105952
R16409 Iout.n641 Iout.n88 0.00105952
R16410 Iout.n632 Iout.n631 0.00105952
R16411 Iout.n629 Iout.n94 0.00105952
R16412 Iout.n620 Iout.n619 0.00105952
R16413 Iout.n617 Iout.n100 0.00105952
R16414 Iout.n608 Iout.n607 0.00105952
R16415 Iout.n605 Iout.n106 0.00105952
R16416 Iout.n596 Iout.n595 0.00105952
R16417 Iout.n593 Iout.n112 0.00105952
R16418 Iout.n584 Iout.n583 0.00105952
R16419 Iout.n973 Iout.n971 0.00105952
R16420 Iout.n970 Iout.n968 0.00105952
R16421 Iout.n565 Iout.n564 0.00105952
R16422 Iout.n581 Iout.n118 0.00105952
R16423 Iout.n978 Iout.n977 0.00105952
R16424 Iout.n122 Iout.n121 0.00105952
R16425 Iout.n568 Iout.n124 0.00105952
R16426 Iout.n571 Iout.n570 0.00105952
R16427 Iout.n335 Iout.n334 0.00105952
R16428 Iout.n338 Iout.n337 0.00105952
R16429 Iout.n341 Iout.n340 0.00105952
R16430 Iout.n344 Iout.n343 0.00105952
R16431 Iout.n347 Iout.n346 0.00105952
R16432 Iout.n350 Iout.n349 0.00105952
R16433 Iout.n353 Iout.n352 0.00105952
R16434 Iout.n356 Iout.n355 0.00105952
R16435 Iout.n359 Iout.n358 0.00105952
R16436 Iout.n372 Iout.n371 0.00105952
R16437 Iout.n385 Iout.n383 0.00105952
R16438 Iout.n388 Iout.n387 0.00105952
R16439 Iout.n401 Iout.n399 0.00105952
R16440 Iout.n404 Iout.n403 0.00105952
R16441 Iout.n417 Iout.n415 0.00105952
R16442 Iout.n420 Iout.n419 0.00105952
R16443 Iout.n433 Iout.n431 0.00105952
R16444 Iout.n443 Iout.n442 0.00105952
R16445 Iout.n440 Iout.n439 0.00105952
R16446 Iout.n437 Iout.n435 0.00105952
R16447 Iout.n555 Iout.n553 0.00105952
R16448 Iout.n558 Iout.n556 0.00105952
R16449 Iout.n981 Iout.n10 0.00105952
R16450 Iout.n984 Iout.n983 0.00105952
R16451 Iout.n561 Iout.n560 0.00105952
R16452 Iout.n992 Iout.n990 0.00105952
R16453 Iout.n989 Iout.n987 0.00105952
R16454 Iout.n129 Iout.n128 0.00105952
R16455 Iout.n547 Iout.n131 0.00105952
R16456 Iout.n550 Iout.n549 0.00105952
R16457 Iout.n451 Iout.n450 0.00105952
R16458 Iout.n454 Iout.n453 0.00105952
R16459 Iout.n448 Iout.n446 0.00105952
R16460 Iout.n428 Iout.n427 0.00105952
R16461 Iout.n425 Iout.n423 0.00105952
R16462 Iout.n412 Iout.n411 0.00105952
R16463 Iout.n409 Iout.n407 0.00105952
R16464 Iout.n396 Iout.n395 0.00105952
R16465 Iout.n393 Iout.n391 0.00105952
R16466 Iout.n331 Iout.n330 0.00105952
R16467 Iout.n328 Iout.n327 0.00105952
R16468 Iout.n325 Iout.n324 0.00105952
R16469 Iout.n322 Iout.n321 0.00105952
R16470 Iout.n319 Iout.n318 0.00105952
R16471 Iout.n316 Iout.n315 0.00105952
R16472 Iout.n313 Iout.n312 0.00105952
R16473 Iout.n310 Iout.n309 0.00105952
R16474 Iout.n307 Iout.n306 0.00105952
R16475 Iout.n459 Iout.n457 0.00105952
R16476 Iout.n465 Iout.n464 0.00105952
R16477 Iout.n462 Iout.n461 0.00105952
R16478 Iout.n544 Iout.n543 0.00105952
R16479 Iout.n541 Iout.n137 0.00105952
R16480 Iout.n997 Iout.n996 0.00105952
R16481 Iout.n135 Iout.n134 0.00105952
R16482 Iout.n1000 Iout.n5 0.00105952
R16483 Iout.n1003 Iout.n1002 0.00105952
R16484 Iout.n538 Iout.n537 0.00105952
R16485 Iout.n535 Iout.n533 0.00105952
R16486 Iout.n532 Iout.n530 0.00105952
R16487 Iout.n468 Iout.n157 0.00105952
R16488 Iout.n471 Iout.n470 0.00105952
R16489 Iout.n474 Iout.n473 0.00105952
R16490 Iout.n264 Iout.n190 0.00105952
R16491 Iout.n267 Iout.n266 0.00105952
R16492 Iout.n276 Iout.n184 0.00105952
R16493 Iout.n279 Iout.n278 0.00105952
R16494 Iout.n288 Iout.n178 0.00105952
R16495 Iout.n291 Iout.n290 0.00105952
R16496 Iout.n300 Iout.n169 0.00105952
R16497 Iout.n173 Iout.n171 0.00105952
R16498 Iout.n297 Iout.n296 0.00105952
R16499 Iout.n294 Iout.n175 0.00105952
R16500 Iout.n285 Iout.n284 0.00105952
R16501 Iout.n282 Iout.n181 0.00105952
R16502 Iout.n273 Iout.n272 0.00105952
R16503 Iout.n270 Iout.n187 0.00105952
R16504 Iout.n261 Iout.n260 0.00105952
R16505 Iout.n479 Iout.n477 0.00105952
R16506 Iout.n485 Iout.n484 0.00105952
R16507 Iout.n482 Iout.n481 0.00105952
R16508 Iout.n527 Iout.n526 0.00105952
R16509 Iout.n524 Iout.n144 0.00105952
R16510 Iout.n142 Iout.n141 0.00105952
R16511 Iout.n1008 Iout.n1006 0.00105952
R16512 Iout.n1011 Iout.n1009 0.00105952
R16513 Iout.n1016 Iout.n1015 0.00105952
R16514 Iout.n148 Iout.n147 0.00105952
R16515 Iout.n518 Iout.n150 0.00105952
R16516 Iout.n521 Iout.n520 0.00105952
R16517 Iout.n493 Iout.n492 0.00105952
R16518 Iout.n496 Iout.n495 0.00105952
R16519 Iout.n490 Iout.n488 0.00105952
R16520 Iout.n254 Iout.n253 0.00105952
R16521 Iout.n257 Iout.n256 0.00105952
R16522 Iout.n251 Iout.n249 0.00105952
R16523 Iout.n248 Iout.n246 0.00105952
R16524 Iout.n245 Iout.n243 0.00105952
R16525 Iout.n242 Iout.n240 0.00105952
R16526 Iout.n239 Iout.n237 0.00105952
R16527 Iout.n236 Iout.n234 0.00105952
R16528 Iout.n233 Iout.n231 0.00105952
R16529 Iout.n228 Iout.n227 0.00105952
R16530 Iout.n225 Iout.n223 0.00105952
R16531 Iout.n221 Iout.n219 0.00105952
R16532 Iout.n217 Iout.n215 0.00105952
R16533 Iout.n213 Iout.n211 0.00105952
R16534 Iout.n209 Iout.n207 0.00105952
R16535 Iout.n205 Iout.n203 0.00105952
R16536 Iout.n201 Iout.n200 0.00105952
R16537 Iout.n198 Iout.n196 0.00105952
R16538 Iout.n194 Iout.n193 0.00105952
R16539 Iout.n501 Iout.n499 0.00105952
R16540 Iout.n505 Iout.n503 0.00105952
R16541 Iout.n508 Iout.n506 0.00105952
R16542 Iout.n515 Iout.n514 0.00105952
R16543 Iout.n512 Iout.n510 0.00105952
R16544 Iout.n1021 Iout.n1019 0.00105952
R16545 XThC.Tn[10].n55 XThC.Tn[10].n54 256.104
R16546 XThC.Tn[10].n59 XThC.Tn[10].n58 243.679
R16547 XThC.Tn[10].n2 XThC.Tn[10].n0 241.847
R16548 XThC.Tn[10].n59 XThC.Tn[10].n57 205.28
R16549 XThC.Tn[10].n55 XThC.Tn[10].n53 202.095
R16550 XThC.Tn[10].n2 XThC.Tn[10].n1 185
R16551 XThC.Tn[10].n5 XThC.Tn[10].n3 161.406
R16552 XThC.Tn[10].n8 XThC.Tn[10].n6 161.406
R16553 XThC.Tn[10].n11 XThC.Tn[10].n9 161.406
R16554 XThC.Tn[10].n14 XThC.Tn[10].n12 161.406
R16555 XThC.Tn[10].n17 XThC.Tn[10].n15 161.406
R16556 XThC.Tn[10].n20 XThC.Tn[10].n18 161.406
R16557 XThC.Tn[10].n23 XThC.Tn[10].n21 161.406
R16558 XThC.Tn[10].n26 XThC.Tn[10].n24 161.406
R16559 XThC.Tn[10].n29 XThC.Tn[10].n27 161.406
R16560 XThC.Tn[10].n32 XThC.Tn[10].n30 161.406
R16561 XThC.Tn[10].n35 XThC.Tn[10].n33 161.406
R16562 XThC.Tn[10].n38 XThC.Tn[10].n36 161.406
R16563 XThC.Tn[10].n41 XThC.Tn[10].n39 161.406
R16564 XThC.Tn[10].n44 XThC.Tn[10].n42 161.406
R16565 XThC.Tn[10].n47 XThC.Tn[10].n45 161.406
R16566 XThC.Tn[10].n50 XThC.Tn[10].n48 161.406
R16567 XThC.Tn[10].n3 XThC.Tn[10].t36 161.202
R16568 XThC.Tn[10].n6 XThC.Tn[10].t21 161.202
R16569 XThC.Tn[10].n9 XThC.Tn[10].t23 161.202
R16570 XThC.Tn[10].n12 XThC.Tn[10].t25 161.202
R16571 XThC.Tn[10].n15 XThC.Tn[10].t14 161.202
R16572 XThC.Tn[10].n18 XThC.Tn[10].t15 161.202
R16573 XThC.Tn[10].n21 XThC.Tn[10].t28 161.202
R16574 XThC.Tn[10].n24 XThC.Tn[10].t37 161.202
R16575 XThC.Tn[10].n27 XThC.Tn[10].t39 161.202
R16576 XThC.Tn[10].n30 XThC.Tn[10].t26 161.202
R16577 XThC.Tn[10].n33 XThC.Tn[10].t27 161.202
R16578 XThC.Tn[10].n36 XThC.Tn[10].t40 161.202
R16579 XThC.Tn[10].n39 XThC.Tn[10].t16 161.202
R16580 XThC.Tn[10].n42 XThC.Tn[10].t19 161.202
R16581 XThC.Tn[10].n45 XThC.Tn[10].t32 161.202
R16582 XThC.Tn[10].n48 XThC.Tn[10].t42 161.202
R16583 XThC.Tn[10].n3 XThC.Tn[10].t38 145.137
R16584 XThC.Tn[10].n6 XThC.Tn[10].t24 145.137
R16585 XThC.Tn[10].n9 XThC.Tn[10].t29 145.137
R16586 XThC.Tn[10].n12 XThC.Tn[10].t30 145.137
R16587 XThC.Tn[10].n15 XThC.Tn[10].t17 145.137
R16588 XThC.Tn[10].n18 XThC.Tn[10].t18 145.137
R16589 XThC.Tn[10].n21 XThC.Tn[10].t34 145.137
R16590 XThC.Tn[10].n24 XThC.Tn[10].t41 145.137
R16591 XThC.Tn[10].n27 XThC.Tn[10].t43 145.137
R16592 XThC.Tn[10].n30 XThC.Tn[10].t31 145.137
R16593 XThC.Tn[10].n33 XThC.Tn[10].t33 145.137
R16594 XThC.Tn[10].n36 XThC.Tn[10].t12 145.137
R16595 XThC.Tn[10].n39 XThC.Tn[10].t20 145.137
R16596 XThC.Tn[10].n42 XThC.Tn[10].t22 145.137
R16597 XThC.Tn[10].n45 XThC.Tn[10].t35 145.137
R16598 XThC.Tn[10].n48 XThC.Tn[10].t13 145.137
R16599 XThC.Tn[10].n53 XThC.Tn[10].t2 26.5955
R16600 XThC.Tn[10].n53 XThC.Tn[10].t1 26.5955
R16601 XThC.Tn[10].n54 XThC.Tn[10].t5 26.5955
R16602 XThC.Tn[10].n54 XThC.Tn[10].t9 26.5955
R16603 XThC.Tn[10].n57 XThC.Tn[10].t7 26.5955
R16604 XThC.Tn[10].n57 XThC.Tn[10].t8 26.5955
R16605 XThC.Tn[10].n58 XThC.Tn[10].t0 26.5955
R16606 XThC.Tn[10].n58 XThC.Tn[10].t4 26.5955
R16607 XThC.Tn[10].n1 XThC.Tn[10].t6 24.9236
R16608 XThC.Tn[10].n1 XThC.Tn[10].t11 24.9236
R16609 XThC.Tn[10].n0 XThC.Tn[10].t10 24.9236
R16610 XThC.Tn[10].n0 XThC.Tn[10].t3 24.9236
R16611 XThC.Tn[10] XThC.Tn[10].n59 22.9652
R16612 XThC.Tn[10] XThC.Tn[10].n2 22.9615
R16613 XThC.Tn[10].n56 XThC.Tn[10].n55 13.9299
R16614 XThC.Tn[10] XThC.Tn[10].n56 13.9299
R16615 XThC.Tn[10].n52 XThC.Tn[10].n51 5.13256
R16616 XThC.Tn[10].n56 XThC.Tn[10].n52 2.99115
R16617 XThC.Tn[10].n56 XThC.Tn[10] 2.87153
R16618 XThC.Tn[10].n52 XThC.Tn[10] 2.2734
R16619 XThC.Tn[10].n51 XThC.Tn[10] 2.26343
R16620 XThC.Tn[10].n8 XThC.Tn[10] 0.931056
R16621 XThC.Tn[10].n11 XThC.Tn[10] 0.931056
R16622 XThC.Tn[10].n14 XThC.Tn[10] 0.931056
R16623 XThC.Tn[10].n17 XThC.Tn[10] 0.931056
R16624 XThC.Tn[10].n20 XThC.Tn[10] 0.931056
R16625 XThC.Tn[10].n23 XThC.Tn[10] 0.931056
R16626 XThC.Tn[10].n26 XThC.Tn[10] 0.931056
R16627 XThC.Tn[10].n29 XThC.Tn[10] 0.931056
R16628 XThC.Tn[10].n32 XThC.Tn[10] 0.931056
R16629 XThC.Tn[10].n35 XThC.Tn[10] 0.931056
R16630 XThC.Tn[10].n38 XThC.Tn[10] 0.931056
R16631 XThC.Tn[10].n41 XThC.Tn[10] 0.931056
R16632 XThC.Tn[10].n44 XThC.Tn[10] 0.931056
R16633 XThC.Tn[10].n47 XThC.Tn[10] 0.931056
R16634 XThC.Tn[10].n50 XThC.Tn[10] 0.931056
R16635 XThC.Tn[10] XThC.Tn[10].n5 0.396333
R16636 XThC.Tn[10] XThC.Tn[10].n8 0.396333
R16637 XThC.Tn[10] XThC.Tn[10].n11 0.396333
R16638 XThC.Tn[10] XThC.Tn[10].n14 0.396333
R16639 XThC.Tn[10] XThC.Tn[10].n17 0.396333
R16640 XThC.Tn[10] XThC.Tn[10].n20 0.396333
R16641 XThC.Tn[10] XThC.Tn[10].n23 0.396333
R16642 XThC.Tn[10] XThC.Tn[10].n26 0.396333
R16643 XThC.Tn[10] XThC.Tn[10].n29 0.396333
R16644 XThC.Tn[10] XThC.Tn[10].n32 0.396333
R16645 XThC.Tn[10] XThC.Tn[10].n35 0.396333
R16646 XThC.Tn[10] XThC.Tn[10].n38 0.396333
R16647 XThC.Tn[10] XThC.Tn[10].n41 0.396333
R16648 XThC.Tn[10] XThC.Tn[10].n44 0.396333
R16649 XThC.Tn[10] XThC.Tn[10].n47 0.396333
R16650 XThC.Tn[10] XThC.Tn[10].n50 0.396333
R16651 XThC.Tn[10].n4 XThC.Tn[10] 0.104667
R16652 XThC.Tn[10].n7 XThC.Tn[10] 0.104667
R16653 XThC.Tn[10].n10 XThC.Tn[10] 0.104667
R16654 XThC.Tn[10].n13 XThC.Tn[10] 0.104667
R16655 XThC.Tn[10].n16 XThC.Tn[10] 0.104667
R16656 XThC.Tn[10].n19 XThC.Tn[10] 0.104667
R16657 XThC.Tn[10].n22 XThC.Tn[10] 0.104667
R16658 XThC.Tn[10].n25 XThC.Tn[10] 0.104667
R16659 XThC.Tn[10].n28 XThC.Tn[10] 0.104667
R16660 XThC.Tn[10].n31 XThC.Tn[10] 0.104667
R16661 XThC.Tn[10].n34 XThC.Tn[10] 0.104667
R16662 XThC.Tn[10].n37 XThC.Tn[10] 0.104667
R16663 XThC.Tn[10].n40 XThC.Tn[10] 0.104667
R16664 XThC.Tn[10].n43 XThC.Tn[10] 0.104667
R16665 XThC.Tn[10].n46 XThC.Tn[10] 0.104667
R16666 XThC.Tn[10].n49 XThC.Tn[10] 0.104667
R16667 XThC.Tn[10].n4 XThC.Tn[10] 0.0309878
R16668 XThC.Tn[10].n7 XThC.Tn[10] 0.0309878
R16669 XThC.Tn[10].n10 XThC.Tn[10] 0.0309878
R16670 XThC.Tn[10].n13 XThC.Tn[10] 0.0309878
R16671 XThC.Tn[10].n16 XThC.Tn[10] 0.0309878
R16672 XThC.Tn[10].n19 XThC.Tn[10] 0.0309878
R16673 XThC.Tn[10].n22 XThC.Tn[10] 0.0309878
R16674 XThC.Tn[10].n25 XThC.Tn[10] 0.0309878
R16675 XThC.Tn[10].n28 XThC.Tn[10] 0.0309878
R16676 XThC.Tn[10].n31 XThC.Tn[10] 0.0309878
R16677 XThC.Tn[10].n34 XThC.Tn[10] 0.0309878
R16678 XThC.Tn[10].n37 XThC.Tn[10] 0.0309878
R16679 XThC.Tn[10].n40 XThC.Tn[10] 0.0309878
R16680 XThC.Tn[10].n43 XThC.Tn[10] 0.0309878
R16681 XThC.Tn[10].n46 XThC.Tn[10] 0.0309878
R16682 XThC.Tn[10].n49 XThC.Tn[10] 0.0309878
R16683 XThC.Tn[10].n5 XThC.Tn[10].n4 0.027939
R16684 XThC.Tn[10].n8 XThC.Tn[10].n7 0.027939
R16685 XThC.Tn[10].n11 XThC.Tn[10].n10 0.027939
R16686 XThC.Tn[10].n14 XThC.Tn[10].n13 0.027939
R16687 XThC.Tn[10].n17 XThC.Tn[10].n16 0.027939
R16688 XThC.Tn[10].n20 XThC.Tn[10].n19 0.027939
R16689 XThC.Tn[10].n23 XThC.Tn[10].n22 0.027939
R16690 XThC.Tn[10].n26 XThC.Tn[10].n25 0.027939
R16691 XThC.Tn[10].n29 XThC.Tn[10].n28 0.027939
R16692 XThC.Tn[10].n32 XThC.Tn[10].n31 0.027939
R16693 XThC.Tn[10].n35 XThC.Tn[10].n34 0.027939
R16694 XThC.Tn[10].n38 XThC.Tn[10].n37 0.027939
R16695 XThC.Tn[10].n41 XThC.Tn[10].n40 0.027939
R16696 XThC.Tn[10].n44 XThC.Tn[10].n43 0.027939
R16697 XThC.Tn[10].n47 XThC.Tn[10].n46 0.027939
R16698 XThC.Tn[10].n50 XThC.Tn[10].n49 0.027939
R16699 XThC.Tn[10].n51 XThC.Tn[10] 0.00285068
R16700 XThR.XTBN.Y.n1 XThR.XTBN.Y.t60 212.081
R16701 XThR.XTBN.Y.n8 XThR.XTBN.Y.t12 212.081
R16702 XThR.XTBN.Y.n2 XThR.XTBN.Y.t81 212.081
R16703 XThR.XTBN.Y.n3 XThR.XTBN.Y.t121 212.081
R16704 XThR.XTBN.Y.n12 XThR.XTBN.Y.t115 212.081
R16705 XThR.XTBN.Y.n19 XThR.XTBN.Y.t65 212.081
R16706 XThR.XTBN.Y.n13 XThR.XTBN.Y.t21 212.081
R16707 XThR.XTBN.Y.n14 XThR.XTBN.Y.t57 212.081
R16708 XThR.XTBN.Y.n24 XThR.XTBN.Y.t27 212.081
R16709 XThR.XTBN.Y.n31 XThR.XTBN.Y.t96 212.081
R16710 XThR.XTBN.Y.n25 XThR.XTBN.Y.t46 212.081
R16711 XThR.XTBN.Y.n26 XThR.XTBN.Y.t89 212.081
R16712 XThR.XTBN.Y.n36 XThR.XTBN.Y.t80 212.081
R16713 XThR.XTBN.Y.n43 XThR.XTBN.Y.t31 212.081
R16714 XThR.XTBN.Y.n37 XThR.XTBN.Y.t102 212.081
R16715 XThR.XTBN.Y.n38 XThR.XTBN.Y.t25 212.081
R16716 XThR.XTBN.Y.n48 XThR.XTBN.Y.t85 212.081
R16717 XThR.XTBN.Y.n55 XThR.XTBN.Y.t33 212.081
R16718 XThR.XTBN.Y.n49 XThR.XTBN.Y.t105 212.081
R16719 XThR.XTBN.Y.n50 XThR.XTBN.Y.t26 212.081
R16720 XThR.XTBN.Y.n60 XThR.XTBN.Y.t54 212.081
R16721 XThR.XTBN.Y.n67 XThR.XTBN.Y.t5 212.081
R16722 XThR.XTBN.Y.n61 XThR.XTBN.Y.t73 212.081
R16723 XThR.XTBN.Y.n62 XThR.XTBN.Y.t114 212.081
R16724 XThR.XTBN.Y.n72 XThR.XTBN.Y.t49 212.081
R16725 XThR.XTBN.Y.n79 XThR.XTBN.Y.t119 212.081
R16726 XThR.XTBN.Y.n73 XThR.XTBN.Y.t69 212.081
R16727 XThR.XTBN.Y.n74 XThR.XTBN.Y.t108 212.081
R16728 XThR.XTBN.Y.n163 XThR.XTBN.Y.t41 212.081
R16729 XThR.XTBN.Y.n154 XThR.XTBN.Y.t113 212.081
R16730 XThR.XTBN.Y.n158 XThR.XTBN.Y.t34 212.081
R16731 XThR.XTBN.Y.n155 XThR.XTBN.Y.t72 212.081
R16732 XThR.XTBN.Y.n151 XThR.XTBN.Y.t19 212.081
R16733 XThR.XTBN.Y.n142 XThR.XTBN.Y.t86 212.081
R16734 XThR.XTBN.Y.n146 XThR.XTBN.Y.t6 212.081
R16735 XThR.XTBN.Y.n143 XThR.XTBN.Y.t43 212.081
R16736 XThR.XTBN.Y.n139 XThR.XTBN.Y.t45 212.081
R16737 XThR.XTBN.Y.n130 XThR.XTBN.Y.t117 212.081
R16738 XThR.XTBN.Y.n134 XThR.XTBN.Y.t36 212.081
R16739 XThR.XTBN.Y.n131 XThR.XTBN.Y.t75 212.081
R16740 XThR.XTBN.Y.n127 XThR.XTBN.Y.t100 212.081
R16741 XThR.XTBN.Y.n118 XThR.XTBN.Y.t50 212.081
R16742 XThR.XTBN.Y.n122 XThR.XTBN.Y.t92 212.081
R16743 XThR.XTBN.Y.n119 XThR.XTBN.Y.t13 212.081
R16744 XThR.XTBN.Y.n115 XThR.XTBN.Y.t15 212.081
R16745 XThR.XTBN.Y.n106 XThR.XTBN.Y.t83 212.081
R16746 XThR.XTBN.Y.n110 XThR.XTBN.Y.t123 212.081
R16747 XThR.XTBN.Y.n107 XThR.XTBN.Y.t39 212.081
R16748 XThR.XTBN.Y.n103 XThR.XTBN.Y.t66 212.081
R16749 XThR.XTBN.Y.n94 XThR.XTBN.Y.t23 212.081
R16750 XThR.XTBN.Y.n98 XThR.XTBN.Y.t59 212.081
R16751 XThR.XTBN.Y.n95 XThR.XTBN.Y.t97 212.081
R16752 XThR.XTBN.Y.n92 XThR.XTBN.Y.t99 212.081
R16753 XThR.XTBN.Y.n83 XThR.XTBN.Y.t87 212.081
R16754 XThR.XTBN.Y.n87 XThR.XTBN.Y.t77 212.081
R16755 XThR.XTBN.Y.n84 XThR.XTBN.Y.t68 212.081
R16756 XThR.XTBN.Y.n167 XThR.XTBN.Y.t63 212.081
R16757 XThR.XTBN.Y.n169 XThR.XTBN.Y.t106 212.081
R16758 XThR.XTBN.Y.n174 XThR.XTBN.Y.t56 212.081
R16759 XThR.XTBN.Y.n170 XThR.XTBN.Y.t7 212.081
R16760 XThR.XTBN.Y XThR.XTBN.Y.n180 203.923
R16761 XThR.XTBN.Y.n171 XThR.XTBN.Y.n170 188.516
R16762 XThR.XTBN.Y.n164 XThR.XTBN.Y.n163 180.482
R16763 XThR.XTBN.Y.n152 XThR.XTBN.Y.n151 180.482
R16764 XThR.XTBN.Y.n140 XThR.XTBN.Y.n139 180.482
R16765 XThR.XTBN.Y.n128 XThR.XTBN.Y.n127 180.482
R16766 XThR.XTBN.Y.n116 XThR.XTBN.Y.n115 180.482
R16767 XThR.XTBN.Y.n104 XThR.XTBN.Y.n103 180.482
R16768 XThR.XTBN.Y.n93 XThR.XTBN.Y.n92 180.482
R16769 XThR.XTBN.Y.n5 XThR.XTBN.Y.n4 173.761
R16770 XThR.XTBN.Y.n16 XThR.XTBN.Y.n15 173.761
R16771 XThR.XTBN.Y.n28 XThR.XTBN.Y.n27 173.761
R16772 XThR.XTBN.Y.n40 XThR.XTBN.Y.n39 173.761
R16773 XThR.XTBN.Y.n52 XThR.XTBN.Y.n51 173.761
R16774 XThR.XTBN.Y.n64 XThR.XTBN.Y.n63 173.761
R16775 XThR.XTBN.Y.n76 XThR.XTBN.Y.n75 173.761
R16776 XThR.XTBN.Y.n168 XThR.XTBN.Y 154.304
R16777 XThR.XTBN.Y.n10 XThR.XTBN.Y.n9 152
R16778 XThR.XTBN.Y.n7 XThR.XTBN.Y.n0 152
R16779 XThR.XTBN.Y.n6 XThR.XTBN.Y.n5 152
R16780 XThR.XTBN.Y.n17 XThR.XTBN.Y.n16 152
R16781 XThR.XTBN.Y.n18 XThR.XTBN.Y.n11 152
R16782 XThR.XTBN.Y.n21 XThR.XTBN.Y.n20 152
R16783 XThR.XTBN.Y.n29 XThR.XTBN.Y.n28 152
R16784 XThR.XTBN.Y.n30 XThR.XTBN.Y.n23 152
R16785 XThR.XTBN.Y.n33 XThR.XTBN.Y.n32 152
R16786 XThR.XTBN.Y.n41 XThR.XTBN.Y.n40 152
R16787 XThR.XTBN.Y.n42 XThR.XTBN.Y.n35 152
R16788 XThR.XTBN.Y.n45 XThR.XTBN.Y.n44 152
R16789 XThR.XTBN.Y.n53 XThR.XTBN.Y.n52 152
R16790 XThR.XTBN.Y.n54 XThR.XTBN.Y.n47 152
R16791 XThR.XTBN.Y.n57 XThR.XTBN.Y.n56 152
R16792 XThR.XTBN.Y.n65 XThR.XTBN.Y.n64 152
R16793 XThR.XTBN.Y.n66 XThR.XTBN.Y.n59 152
R16794 XThR.XTBN.Y.n69 XThR.XTBN.Y.n68 152
R16795 XThR.XTBN.Y.n77 XThR.XTBN.Y.n76 152
R16796 XThR.XTBN.Y.n78 XThR.XTBN.Y.n71 152
R16797 XThR.XTBN.Y.n81 XThR.XTBN.Y.n80 152
R16798 XThR.XTBN.Y.n157 XThR.XTBN.Y.n156 152
R16799 XThR.XTBN.Y.n160 XThR.XTBN.Y.n159 152
R16800 XThR.XTBN.Y.n162 XThR.XTBN.Y.n161 152
R16801 XThR.XTBN.Y.n145 XThR.XTBN.Y.n144 152
R16802 XThR.XTBN.Y.n148 XThR.XTBN.Y.n147 152
R16803 XThR.XTBN.Y.n150 XThR.XTBN.Y.n149 152
R16804 XThR.XTBN.Y.n133 XThR.XTBN.Y.n132 152
R16805 XThR.XTBN.Y.n136 XThR.XTBN.Y.n135 152
R16806 XThR.XTBN.Y.n138 XThR.XTBN.Y.n137 152
R16807 XThR.XTBN.Y.n121 XThR.XTBN.Y.n120 152
R16808 XThR.XTBN.Y.n124 XThR.XTBN.Y.n123 152
R16809 XThR.XTBN.Y.n126 XThR.XTBN.Y.n125 152
R16810 XThR.XTBN.Y.n109 XThR.XTBN.Y.n108 152
R16811 XThR.XTBN.Y.n112 XThR.XTBN.Y.n111 152
R16812 XThR.XTBN.Y.n114 XThR.XTBN.Y.n113 152
R16813 XThR.XTBN.Y.n97 XThR.XTBN.Y.n96 152
R16814 XThR.XTBN.Y.n100 XThR.XTBN.Y.n99 152
R16815 XThR.XTBN.Y.n102 XThR.XTBN.Y.n101 152
R16816 XThR.XTBN.Y.n86 XThR.XTBN.Y.n85 152
R16817 XThR.XTBN.Y.n89 XThR.XTBN.Y.n88 152
R16818 XThR.XTBN.Y.n91 XThR.XTBN.Y.n90 152
R16819 XThR.XTBN.Y.n173 XThR.XTBN.Y.n172 152
R16820 XThR.XTBN.Y.n176 XThR.XTBN.Y.n175 152
R16821 XThR.XTBN.Y.n1 XThR.XTBN.Y.t95 139.78
R16822 XThR.XTBN.Y.n8 XThR.XTBN.Y.t44 139.78
R16823 XThR.XTBN.Y.n2 XThR.XTBN.Y.t116 139.78
R16824 XThR.XTBN.Y.n3 XThR.XTBN.Y.t35 139.78
R16825 XThR.XTBN.Y.n12 XThR.XTBN.Y.t42 139.78
R16826 XThR.XTBN.Y.n19 XThR.XTBN.Y.t112 139.78
R16827 XThR.XTBN.Y.n13 XThR.XTBN.Y.t64 139.78
R16828 XThR.XTBN.Y.n14 XThR.XTBN.Y.t107 139.78
R16829 XThR.XTBN.Y.n24 XThR.XTBN.Y.t61 139.78
R16830 XThR.XTBN.Y.n31 XThR.XTBN.Y.t14 139.78
R16831 XThR.XTBN.Y.n25 XThR.XTBN.Y.t82 139.78
R16832 XThR.XTBN.Y.n26 XThR.XTBN.Y.t122 139.78
R16833 XThR.XTBN.Y.n36 XThR.XTBN.Y.t11 139.78
R16834 XThR.XTBN.Y.n43 XThR.XTBN.Y.t79 139.78
R16835 XThR.XTBN.Y.n37 XThR.XTBN.Y.t32 139.78
R16836 XThR.XTBN.Y.n38 XThR.XTBN.Y.t71 139.78
R16837 XThR.XTBN.Y.n48 XThR.XTBN.Y.t29 139.78
R16838 XThR.XTBN.Y.n55 XThR.XTBN.Y.t98 139.78
R16839 XThR.XTBN.Y.n49 XThR.XTBN.Y.t47 139.78
R16840 XThR.XTBN.Y.n50 XThR.XTBN.Y.t90 139.78
R16841 XThR.XTBN.Y.n60 XThR.XTBN.Y.t8 139.78
R16842 XThR.XTBN.Y.n67 XThR.XTBN.Y.t74 139.78
R16843 XThR.XTBN.Y.n61 XThR.XTBN.Y.t28 139.78
R16844 XThR.XTBN.Y.n62 XThR.XTBN.Y.t67 139.78
R16845 XThR.XTBN.Y.n72 XThR.XTBN.Y.t111 139.78
R16846 XThR.XTBN.Y.n79 XThR.XTBN.Y.t62 139.78
R16847 XThR.XTBN.Y.n73 XThR.XTBN.Y.t18 139.78
R16848 XThR.XTBN.Y.n74 XThR.XTBN.Y.t53 139.78
R16849 XThR.XTBN.Y.n163 XThR.XTBN.Y.t101 139.78
R16850 XThR.XTBN.Y.n154 XThR.XTBN.Y.t52 139.78
R16851 XThR.XTBN.Y.n158 XThR.XTBN.Y.t93 139.78
R16852 XThR.XTBN.Y.n155 XThR.XTBN.Y.t16 139.78
R16853 XThR.XTBN.Y.n151 XThR.XTBN.Y.t88 139.78
R16854 XThR.XTBN.Y.n142 XThR.XTBN.Y.t37 139.78
R16855 XThR.XTBN.Y.n146 XThR.XTBN.Y.t76 139.78
R16856 XThR.XTBN.Y.n143 XThR.XTBN.Y.t118 139.78
R16857 XThR.XTBN.Y.n139 XThR.XTBN.Y.t104 139.78
R16858 XThR.XTBN.Y.n130 XThR.XTBN.Y.t55 139.78
R16859 XThR.XTBN.Y.n134 XThR.XTBN.Y.t94 139.78
R16860 XThR.XTBN.Y.n131 XThR.XTBN.Y.t17 139.78
R16861 XThR.XTBN.Y.n127 XThR.XTBN.Y.t51 139.78
R16862 XThR.XTBN.Y.n118 XThR.XTBN.Y.t4 139.78
R16863 XThR.XTBN.Y.n122 XThR.XTBN.Y.t40 139.78
R16864 XThR.XTBN.Y.n119 XThR.XTBN.Y.t84 139.78
R16865 XThR.XTBN.Y.n115 XThR.XTBN.Y.t38 139.78
R16866 XThR.XTBN.Y.n106 XThR.XTBN.Y.t109 139.78
R16867 XThR.XTBN.Y.n110 XThR.XTBN.Y.t30 139.78
R16868 XThR.XTBN.Y.n107 XThR.XTBN.Y.t70 139.78
R16869 XThR.XTBN.Y.n103 XThR.XTBN.Y.t24 139.78
R16870 XThR.XTBN.Y.n94 XThR.XTBN.Y.t91 139.78
R16871 XThR.XTBN.Y.n98 XThR.XTBN.Y.t10 139.78
R16872 XThR.XTBN.Y.n95 XThR.XTBN.Y.t48 139.78
R16873 XThR.XTBN.Y.n92 XThR.XTBN.Y.t20 139.78
R16874 XThR.XTBN.Y.n83 XThR.XTBN.Y.t120 139.78
R16875 XThR.XTBN.Y.n87 XThR.XTBN.Y.t110 139.78
R16876 XThR.XTBN.Y.n84 XThR.XTBN.Y.t103 139.78
R16877 XThR.XTBN.Y.n167 XThR.XTBN.Y.t22 139.78
R16878 XThR.XTBN.Y.n169 XThR.XTBN.Y.t58 139.78
R16879 XThR.XTBN.Y.n174 XThR.XTBN.Y.t9 139.78
R16880 XThR.XTBN.Y.n170 XThR.XTBN.Y.t78 139.78
R16881 XThR.XTBN.Y.n184 XThR.XTBN.Y.n183 101.489
R16882 XThR.XTBN.Y.n179 XThR.XTBN.Y 58.2909
R16883 XThR.XTBN.Y.n7 XThR.XTBN.Y.n6 49.6611
R16884 XThR.XTBN.Y.n18 XThR.XTBN.Y.n17 49.6611
R16885 XThR.XTBN.Y.n30 XThR.XTBN.Y.n29 49.6611
R16886 XThR.XTBN.Y.n42 XThR.XTBN.Y.n41 49.6611
R16887 XThR.XTBN.Y.n54 XThR.XTBN.Y.n53 49.6611
R16888 XThR.XTBN.Y.n66 XThR.XTBN.Y.n65 49.6611
R16889 XThR.XTBN.Y.n78 XThR.XTBN.Y.n77 49.6611
R16890 XThR.XTBN.Y.n9 XThR.XTBN.Y.n8 44.549
R16891 XThR.XTBN.Y.n20 XThR.XTBN.Y.n19 44.549
R16892 XThR.XTBN.Y.n32 XThR.XTBN.Y.n31 44.549
R16893 XThR.XTBN.Y.n44 XThR.XTBN.Y.n43 44.549
R16894 XThR.XTBN.Y.n56 XThR.XTBN.Y.n55 44.549
R16895 XThR.XTBN.Y.n68 XThR.XTBN.Y.n67 44.549
R16896 XThR.XTBN.Y.n80 XThR.XTBN.Y.n79 44.549
R16897 XThR.XTBN.Y.n4 XThR.XTBN.Y.n2 43.0884
R16898 XThR.XTBN.Y.n15 XThR.XTBN.Y.n13 43.0884
R16899 XThR.XTBN.Y.n27 XThR.XTBN.Y.n25 43.0884
R16900 XThR.XTBN.Y.n39 XThR.XTBN.Y.n37 43.0884
R16901 XThR.XTBN.Y.n51 XThR.XTBN.Y.n49 43.0884
R16902 XThR.XTBN.Y.n63 XThR.XTBN.Y.n61 43.0884
R16903 XThR.XTBN.Y.n75 XThR.XTBN.Y.n73 43.0884
R16904 XThR.XTBN.Y.n163 XThR.XTBN.Y.n162 30.6732
R16905 XThR.XTBN.Y.n162 XThR.XTBN.Y.n154 30.6732
R16906 XThR.XTBN.Y.n159 XThR.XTBN.Y.n154 30.6732
R16907 XThR.XTBN.Y.n159 XThR.XTBN.Y.n158 30.6732
R16908 XThR.XTBN.Y.n158 XThR.XTBN.Y.n157 30.6732
R16909 XThR.XTBN.Y.n157 XThR.XTBN.Y.n155 30.6732
R16910 XThR.XTBN.Y.n151 XThR.XTBN.Y.n150 30.6732
R16911 XThR.XTBN.Y.n150 XThR.XTBN.Y.n142 30.6732
R16912 XThR.XTBN.Y.n147 XThR.XTBN.Y.n142 30.6732
R16913 XThR.XTBN.Y.n147 XThR.XTBN.Y.n146 30.6732
R16914 XThR.XTBN.Y.n146 XThR.XTBN.Y.n145 30.6732
R16915 XThR.XTBN.Y.n145 XThR.XTBN.Y.n143 30.6732
R16916 XThR.XTBN.Y.n139 XThR.XTBN.Y.n138 30.6732
R16917 XThR.XTBN.Y.n138 XThR.XTBN.Y.n130 30.6732
R16918 XThR.XTBN.Y.n135 XThR.XTBN.Y.n130 30.6732
R16919 XThR.XTBN.Y.n135 XThR.XTBN.Y.n134 30.6732
R16920 XThR.XTBN.Y.n134 XThR.XTBN.Y.n133 30.6732
R16921 XThR.XTBN.Y.n133 XThR.XTBN.Y.n131 30.6732
R16922 XThR.XTBN.Y.n127 XThR.XTBN.Y.n126 30.6732
R16923 XThR.XTBN.Y.n126 XThR.XTBN.Y.n118 30.6732
R16924 XThR.XTBN.Y.n123 XThR.XTBN.Y.n118 30.6732
R16925 XThR.XTBN.Y.n123 XThR.XTBN.Y.n122 30.6732
R16926 XThR.XTBN.Y.n122 XThR.XTBN.Y.n121 30.6732
R16927 XThR.XTBN.Y.n121 XThR.XTBN.Y.n119 30.6732
R16928 XThR.XTBN.Y.n115 XThR.XTBN.Y.n114 30.6732
R16929 XThR.XTBN.Y.n114 XThR.XTBN.Y.n106 30.6732
R16930 XThR.XTBN.Y.n111 XThR.XTBN.Y.n106 30.6732
R16931 XThR.XTBN.Y.n111 XThR.XTBN.Y.n110 30.6732
R16932 XThR.XTBN.Y.n110 XThR.XTBN.Y.n109 30.6732
R16933 XThR.XTBN.Y.n109 XThR.XTBN.Y.n107 30.6732
R16934 XThR.XTBN.Y.n103 XThR.XTBN.Y.n102 30.6732
R16935 XThR.XTBN.Y.n102 XThR.XTBN.Y.n94 30.6732
R16936 XThR.XTBN.Y.n99 XThR.XTBN.Y.n94 30.6732
R16937 XThR.XTBN.Y.n99 XThR.XTBN.Y.n98 30.6732
R16938 XThR.XTBN.Y.n98 XThR.XTBN.Y.n97 30.6732
R16939 XThR.XTBN.Y.n97 XThR.XTBN.Y.n95 30.6732
R16940 XThR.XTBN.Y.n92 XThR.XTBN.Y.n91 30.6732
R16941 XThR.XTBN.Y.n91 XThR.XTBN.Y.n83 30.6732
R16942 XThR.XTBN.Y.n88 XThR.XTBN.Y.n83 30.6732
R16943 XThR.XTBN.Y.n88 XThR.XTBN.Y.n87 30.6732
R16944 XThR.XTBN.Y.n87 XThR.XTBN.Y.n86 30.6732
R16945 XThR.XTBN.Y.n86 XThR.XTBN.Y.n84 30.6732
R16946 XThR.XTBN.Y.n168 XThR.XTBN.Y.n167 30.6732
R16947 XThR.XTBN.Y.n169 XThR.XTBN.Y.n168 30.6732
R16948 XThR.XTBN.Y.n175 XThR.XTBN.Y.n169 30.6732
R16949 XThR.XTBN.Y.n175 XThR.XTBN.Y.n174 30.6732
R16950 XThR.XTBN.Y.n174 XThR.XTBN.Y.n173 30.6732
R16951 XThR.XTBN.Y.n173 XThR.XTBN.Y.n170 30.6732
R16952 XThR.XTBN.Y.n180 XThR.XTBN.Y.t3 26.5955
R16953 XThR.XTBN.Y.n180 XThR.XTBN.Y.t2 26.5955
R16954 XThR.XTBN.Y.n183 XThR.XTBN.Y.t0 24.9236
R16955 XThR.XTBN.Y.n183 XThR.XTBN.Y.t1 24.9236
R16956 XThR.XTBN.Y.n10 XThR.XTBN.Y.n0 21.7605
R16957 XThR.XTBN.Y.n21 XThR.XTBN.Y.n11 21.7605
R16958 XThR.XTBN.Y.n33 XThR.XTBN.Y.n23 21.7605
R16959 XThR.XTBN.Y.n45 XThR.XTBN.Y.n35 21.7605
R16960 XThR.XTBN.Y.n57 XThR.XTBN.Y.n47 21.7605
R16961 XThR.XTBN.Y.n69 XThR.XTBN.Y.n59 21.7605
R16962 XThR.XTBN.Y.n81 XThR.XTBN.Y.n71 21.7605
R16963 XThR.XTBN.Y.n161 XThR.XTBN.Y 18.4325
R16964 XThR.XTBN.Y.n149 XThR.XTBN.Y 18.4325
R16965 XThR.XTBN.Y.n137 XThR.XTBN.Y 18.4325
R16966 XThR.XTBN.Y.n125 XThR.XTBN.Y 18.4325
R16967 XThR.XTBN.Y.n113 XThR.XTBN.Y 18.4325
R16968 XThR.XTBN.Y.n101 XThR.XTBN.Y 18.4325
R16969 XThR.XTBN.Y.n90 XThR.XTBN.Y 18.4325
R16970 XThR.XTBN.Y.n4 XThR.XTBN.Y.n3 18.2581
R16971 XThR.XTBN.Y.n15 XThR.XTBN.Y.n14 18.2581
R16972 XThR.XTBN.Y.n27 XThR.XTBN.Y.n26 18.2581
R16973 XThR.XTBN.Y.n39 XThR.XTBN.Y.n38 18.2581
R16974 XThR.XTBN.Y.n51 XThR.XTBN.Y.n50 18.2581
R16975 XThR.XTBN.Y.n63 XThR.XTBN.Y.n62 18.2581
R16976 XThR.XTBN.Y.n75 XThR.XTBN.Y.n74 18.2581
R16977 XThR.XTBN.Y.n5 XThR.XTBN.Y 17.6005
R16978 XThR.XTBN.Y.n16 XThR.XTBN.Y 17.6005
R16979 XThR.XTBN.Y.n28 XThR.XTBN.Y 17.6005
R16980 XThR.XTBN.Y.n40 XThR.XTBN.Y 17.6005
R16981 XThR.XTBN.Y.n52 XThR.XTBN.Y 17.6005
R16982 XThR.XTBN.Y.n64 XThR.XTBN.Y 17.6005
R16983 XThR.XTBN.Y.n76 XThR.XTBN.Y 17.6005
R16984 XThR.XTBN.Y.n22 XThR.XTBN.Y.n10 17.1655
R16985 XThR.XTBN.Y.n172 XThR.XTBN.Y 17.1525
R16986 XThR.XTBN.Y XThR.XTBN.Y.n171 17.1525
R16987 XThR.XTBN.Y.n105 XThR.XTBN.Y.n93 17.054
R16988 XThR.XTBN.Y.n9 XThR.XTBN.Y.n1 16.7975
R16989 XThR.XTBN.Y.n20 XThR.XTBN.Y.n12 16.7975
R16990 XThR.XTBN.Y.n32 XThR.XTBN.Y.n24 16.7975
R16991 XThR.XTBN.Y.n44 XThR.XTBN.Y.n36 16.7975
R16992 XThR.XTBN.Y.n56 XThR.XTBN.Y.n48 16.7975
R16993 XThR.XTBN.Y.n68 XThR.XTBN.Y.n60 16.7975
R16994 XThR.XTBN.Y.n80 XThR.XTBN.Y.n72 16.7975
R16995 XThR.XTBN.Y XThR.XTBN.Y.n160 16.3845
R16996 XThR.XTBN.Y XThR.XTBN.Y.n148 16.3845
R16997 XThR.XTBN.Y XThR.XTBN.Y.n136 16.3845
R16998 XThR.XTBN.Y XThR.XTBN.Y.n124 16.3845
R16999 XThR.XTBN.Y XThR.XTBN.Y.n112 16.3845
R17000 XThR.XTBN.Y XThR.XTBN.Y.n100 16.3845
R17001 XThR.XTBN.Y XThR.XTBN.Y.n89 16.3845
R17002 XThR.XTBN.Y.n22 XThR.XTBN.Y.n21 16.0405
R17003 XThR.XTBN.Y.n34 XThR.XTBN.Y.n33 16.0405
R17004 XThR.XTBN.Y.n46 XThR.XTBN.Y.n45 16.0405
R17005 XThR.XTBN.Y.n58 XThR.XTBN.Y.n57 16.0405
R17006 XThR.XTBN.Y.n70 XThR.XTBN.Y.n69 16.0405
R17007 XThR.XTBN.Y.n82 XThR.XTBN.Y.n81 16.0405
R17008 XThR.XTBN.Y.n165 XThR.XTBN.Y.n164 15.5925
R17009 XThR.XTBN.Y.n153 XThR.XTBN.Y.n152 15.5925
R17010 XThR.XTBN.Y.n141 XThR.XTBN.Y.n140 15.5925
R17011 XThR.XTBN.Y.n129 XThR.XTBN.Y.n128 15.5925
R17012 XThR.XTBN.Y.n117 XThR.XTBN.Y.n116 15.5925
R17013 XThR.XTBN.Y.n105 XThR.XTBN.Y.n104 15.5925
R17014 XThR.XTBN.Y.n156 XThR.XTBN.Y 14.3365
R17015 XThR.XTBN.Y.n144 XThR.XTBN.Y 14.3365
R17016 XThR.XTBN.Y.n132 XThR.XTBN.Y 14.3365
R17017 XThR.XTBN.Y.n120 XThR.XTBN.Y 14.3365
R17018 XThR.XTBN.Y.n108 XThR.XTBN.Y 14.3365
R17019 XThR.XTBN.Y.n96 XThR.XTBN.Y 14.3365
R17020 XThR.XTBN.Y.n85 XThR.XTBN.Y 14.3365
R17021 XThR.XTBN.Y XThR.XTBN.Y.n182 13.5685
R17022 XThR.XTBN.Y.n177 XThR.XTBN.Y.n176 12.2885
R17023 XThR.XTBN.Y XThR.XTBN.Y.n181 10.7525
R17024 XThR.XTBN.Y.n156 XThR.XTBN.Y 9.2165
R17025 XThR.XTBN.Y.n144 XThR.XTBN.Y 9.2165
R17026 XThR.XTBN.Y.n132 XThR.XTBN.Y 9.2165
R17027 XThR.XTBN.Y.n120 XThR.XTBN.Y 9.2165
R17028 XThR.XTBN.Y.n108 XThR.XTBN.Y 9.2165
R17029 XThR.XTBN.Y.n96 XThR.XTBN.Y 9.2165
R17030 XThR.XTBN.Y.n85 XThR.XTBN.Y 9.2165
R17031 XThR.XTBN.Y.n160 XThR.XTBN.Y 7.1685
R17032 XThR.XTBN.Y.n148 XThR.XTBN.Y 7.1685
R17033 XThR.XTBN.Y.n136 XThR.XTBN.Y 7.1685
R17034 XThR.XTBN.Y.n124 XThR.XTBN.Y 7.1685
R17035 XThR.XTBN.Y.n112 XThR.XTBN.Y 7.1685
R17036 XThR.XTBN.Y.n100 XThR.XTBN.Y 7.1685
R17037 XThR.XTBN.Y.n89 XThR.XTBN.Y 7.1685
R17038 XThR.XTBN.Y.n177 XThR.XTBN.Y 6.9125
R17039 XThR.XTBN.Y.n181 XThR.XTBN.Y 6.6565
R17040 XThR.XTBN.Y.n6 XThR.XTBN.Y.n2 6.57323
R17041 XThR.XTBN.Y.n17 XThR.XTBN.Y.n13 6.57323
R17042 XThR.XTBN.Y.n29 XThR.XTBN.Y.n25 6.57323
R17043 XThR.XTBN.Y.n41 XThR.XTBN.Y.n37 6.57323
R17044 XThR.XTBN.Y.n53 XThR.XTBN.Y.n49 6.57323
R17045 XThR.XTBN.Y.n65 XThR.XTBN.Y.n61 6.57323
R17046 XThR.XTBN.Y.n77 XThR.XTBN.Y.n73 6.57323
R17047 XThR.XTBN.Y.n172 XThR.XTBN.Y 6.4005
R17048 XThR.XTBN.Y.n171 XThR.XTBN.Y 6.4005
R17049 XThR.XTBN.Y.n179 XThR.XTBN.Y.n178 5.74665
R17050 XThR.XTBN.Y.n178 XThR.XTBN.Y.n166 5.74569
R17051 XThR.XTBN.Y.n161 XThR.XTBN.Y 5.1205
R17052 XThR.XTBN.Y.n149 XThR.XTBN.Y 5.1205
R17053 XThR.XTBN.Y.n137 XThR.XTBN.Y 5.1205
R17054 XThR.XTBN.Y.n125 XThR.XTBN.Y 5.1205
R17055 XThR.XTBN.Y.n113 XThR.XTBN.Y 5.1205
R17056 XThR.XTBN.Y.n101 XThR.XTBN.Y 5.1205
R17057 XThR.XTBN.Y.n90 XThR.XTBN.Y 5.1205
R17058 XThR.XTBN.Y.n8 XThR.XTBN.Y.n7 5.11262
R17059 XThR.XTBN.Y.n19 XThR.XTBN.Y.n18 5.11262
R17060 XThR.XTBN.Y.n31 XThR.XTBN.Y.n30 5.11262
R17061 XThR.XTBN.Y.n43 XThR.XTBN.Y.n42 5.11262
R17062 XThR.XTBN.Y.n55 XThR.XTBN.Y.n54 5.11262
R17063 XThR.XTBN.Y.n67 XThR.XTBN.Y.n66 5.11262
R17064 XThR.XTBN.Y.n79 XThR.XTBN.Y.n78 5.11262
R17065 XThR.XTBN.Y.n182 XThR.XTBN.Y.n179 5.06717
R17066 XThR.XTBN.Y.n181 XThR.XTBN.Y 5.04292
R17067 XThR.XTBN.Y.n178 XThR.XTBN.Y.n177 4.6505
R17068 XThR.XTBN.Y.n176 XThR.XTBN.Y 4.3525
R17069 XThR.XTBN.Y XThR.XTBN.Y.n0 4.1605
R17070 XThR.XTBN.Y XThR.XTBN.Y.n11 4.1605
R17071 XThR.XTBN.Y XThR.XTBN.Y.n23 4.1605
R17072 XThR.XTBN.Y XThR.XTBN.Y.n35 4.1605
R17073 XThR.XTBN.Y XThR.XTBN.Y.n47 4.1605
R17074 XThR.XTBN.Y XThR.XTBN.Y.n59 4.1605
R17075 XThR.XTBN.Y XThR.XTBN.Y.n71 4.1605
R17076 XThR.XTBN.Y.n182 XThR.XTBN.Y 3.8405
R17077 XThR.XTBN.Y.n184 XThR.XTBN.Y 2.5605
R17078 XThR.XTBN.Y.n164 XThR.XTBN.Y 2.3045
R17079 XThR.XTBN.Y.n152 XThR.XTBN.Y 2.3045
R17080 XThR.XTBN.Y.n140 XThR.XTBN.Y 2.3045
R17081 XThR.XTBN.Y.n128 XThR.XTBN.Y 2.3045
R17082 XThR.XTBN.Y.n116 XThR.XTBN.Y 2.3045
R17083 XThR.XTBN.Y.n104 XThR.XTBN.Y 2.3045
R17084 XThR.XTBN.Y.n93 XThR.XTBN.Y 2.3045
R17085 XThR.XTBN.Y XThR.XTBN.Y.n184 1.93989
R17086 XThR.XTBN.Y.n166 XThR.XTBN.Y.n82 1.53415
R17087 XThR.XTBN.Y.n34 XThR.XTBN.Y.n22 1.49088
R17088 XThR.XTBN.Y.n58 XThR.XTBN.Y.n46 1.49088
R17089 XThR.XTBN.Y.n82 XThR.XTBN.Y.n70 1.48608
R17090 XThR.XTBN.Y.n153 XThR.XTBN.Y.n141 1.46204
R17091 XThR.XTBN.Y.n129 XThR.XTBN.Y.n117 1.46204
R17092 XThR.XTBN.Y.n166 XThR.XTBN.Y.n165 1.20723
R17093 XThR.XTBN.Y.n165 XThR.XTBN.Y.n153 1.15435
R17094 XThR.XTBN.Y.n141 XThR.XTBN.Y.n129 1.15435
R17095 XThR.XTBN.Y.n117 XThR.XTBN.Y.n105 1.15435
R17096 XThR.XTBN.Y.n70 XThR.XTBN.Y.n58 1.13031
R17097 XThR.XTBN.Y.n46 XThR.XTBN.Y.n34 1.1255
R17098 XThR.Tn[6].n2 XThR.Tn[6].n1 332.332
R17099 XThR.Tn[6].n2 XThR.Tn[6].n0 296.493
R17100 XThR.Tn[6] XThR.Tn[6].n82 161.363
R17101 XThR.Tn[6] XThR.Tn[6].n77 161.363
R17102 XThR.Tn[6] XThR.Tn[6].n72 161.363
R17103 XThR.Tn[6] XThR.Tn[6].n67 161.363
R17104 XThR.Tn[6] XThR.Tn[6].n62 161.363
R17105 XThR.Tn[6] XThR.Tn[6].n57 161.363
R17106 XThR.Tn[6] XThR.Tn[6].n52 161.363
R17107 XThR.Tn[6] XThR.Tn[6].n47 161.363
R17108 XThR.Tn[6] XThR.Tn[6].n42 161.363
R17109 XThR.Tn[6] XThR.Tn[6].n37 161.363
R17110 XThR.Tn[6] XThR.Tn[6].n32 161.363
R17111 XThR.Tn[6] XThR.Tn[6].n27 161.363
R17112 XThR.Tn[6] XThR.Tn[6].n22 161.363
R17113 XThR.Tn[6] XThR.Tn[6].n17 161.363
R17114 XThR.Tn[6] XThR.Tn[6].n12 161.363
R17115 XThR.Tn[6] XThR.Tn[6].n10 161.363
R17116 XThR.Tn[6].n84 XThR.Tn[6].n83 161.3
R17117 XThR.Tn[6].n79 XThR.Tn[6].n78 161.3
R17118 XThR.Tn[6].n74 XThR.Tn[6].n73 161.3
R17119 XThR.Tn[6].n69 XThR.Tn[6].n68 161.3
R17120 XThR.Tn[6].n64 XThR.Tn[6].n63 161.3
R17121 XThR.Tn[6].n59 XThR.Tn[6].n58 161.3
R17122 XThR.Tn[6].n54 XThR.Tn[6].n53 161.3
R17123 XThR.Tn[6].n49 XThR.Tn[6].n48 161.3
R17124 XThR.Tn[6].n44 XThR.Tn[6].n43 161.3
R17125 XThR.Tn[6].n39 XThR.Tn[6].n38 161.3
R17126 XThR.Tn[6].n34 XThR.Tn[6].n33 161.3
R17127 XThR.Tn[6].n29 XThR.Tn[6].n28 161.3
R17128 XThR.Tn[6].n24 XThR.Tn[6].n23 161.3
R17129 XThR.Tn[6].n19 XThR.Tn[6].n18 161.3
R17130 XThR.Tn[6].n14 XThR.Tn[6].n13 161.3
R17131 XThR.Tn[6].n82 XThR.Tn[6].t46 161.106
R17132 XThR.Tn[6].n77 XThR.Tn[6].t52 161.106
R17133 XThR.Tn[6].n72 XThR.Tn[6].t32 161.106
R17134 XThR.Tn[6].n67 XThR.Tn[6].t18 161.106
R17135 XThR.Tn[6].n62 XThR.Tn[6].t44 161.106
R17136 XThR.Tn[6].n57 XThR.Tn[6].t69 161.106
R17137 XThR.Tn[6].n52 XThR.Tn[6].t50 161.106
R17138 XThR.Tn[6].n47 XThR.Tn[6].t30 161.106
R17139 XThR.Tn[6].n42 XThR.Tn[6].t17 161.106
R17140 XThR.Tn[6].n37 XThR.Tn[6].t22 161.106
R17141 XThR.Tn[6].n32 XThR.Tn[6].t67 161.106
R17142 XThR.Tn[6].n27 XThR.Tn[6].t31 161.106
R17143 XThR.Tn[6].n22 XThR.Tn[6].t66 161.106
R17144 XThR.Tn[6].n17 XThR.Tn[6].t49 161.106
R17145 XThR.Tn[6].n12 XThR.Tn[6].t72 161.106
R17146 XThR.Tn[6].n10 XThR.Tn[6].t56 161.106
R17147 XThR.Tn[6].n83 XThR.Tn[6].t42 159.978
R17148 XThR.Tn[6].n78 XThR.Tn[6].t48 159.978
R17149 XThR.Tn[6].n73 XThR.Tn[6].t28 159.978
R17150 XThR.Tn[6].n68 XThR.Tn[6].t15 159.978
R17151 XThR.Tn[6].n63 XThR.Tn[6].t39 159.978
R17152 XThR.Tn[6].n58 XThR.Tn[6].t65 159.978
R17153 XThR.Tn[6].n53 XThR.Tn[6].t47 159.978
R17154 XThR.Tn[6].n48 XThR.Tn[6].t25 159.978
R17155 XThR.Tn[6].n43 XThR.Tn[6].t12 159.978
R17156 XThR.Tn[6].n38 XThR.Tn[6].t19 159.978
R17157 XThR.Tn[6].n33 XThR.Tn[6].t64 159.978
R17158 XThR.Tn[6].n28 XThR.Tn[6].t27 159.978
R17159 XThR.Tn[6].n23 XThR.Tn[6].t63 159.978
R17160 XThR.Tn[6].n18 XThR.Tn[6].t45 159.978
R17161 XThR.Tn[6].n13 XThR.Tn[6].t68 159.978
R17162 XThR.Tn[6].n82 XThR.Tn[6].t34 145.038
R17163 XThR.Tn[6].n77 XThR.Tn[6].t58 145.038
R17164 XThR.Tn[6].n72 XThR.Tn[6].t38 145.038
R17165 XThR.Tn[6].n67 XThR.Tn[6].t23 145.038
R17166 XThR.Tn[6].n62 XThR.Tn[6].t53 145.038
R17167 XThR.Tn[6].n57 XThR.Tn[6].t33 145.038
R17168 XThR.Tn[6].n52 XThR.Tn[6].t40 145.038
R17169 XThR.Tn[6].n47 XThR.Tn[6].t24 145.038
R17170 XThR.Tn[6].n42 XThR.Tn[6].t21 145.038
R17171 XThR.Tn[6].n37 XThR.Tn[6].t51 145.038
R17172 XThR.Tn[6].n32 XThR.Tn[6].t13 145.038
R17173 XThR.Tn[6].n27 XThR.Tn[6].t35 145.038
R17174 XThR.Tn[6].n22 XThR.Tn[6].t73 145.038
R17175 XThR.Tn[6].n17 XThR.Tn[6].t57 145.038
R17176 XThR.Tn[6].n12 XThR.Tn[6].t20 145.038
R17177 XThR.Tn[6].n10 XThR.Tn[6].t62 145.038
R17178 XThR.Tn[6].n83 XThR.Tn[6].t55 143.911
R17179 XThR.Tn[6].n78 XThR.Tn[6].t16 143.911
R17180 XThR.Tn[6].n73 XThR.Tn[6].t60 143.911
R17181 XThR.Tn[6].n68 XThR.Tn[6].t41 143.911
R17182 XThR.Tn[6].n63 XThR.Tn[6].t71 143.911
R17183 XThR.Tn[6].n58 XThR.Tn[6].t54 143.911
R17184 XThR.Tn[6].n53 XThR.Tn[6].t61 143.911
R17185 XThR.Tn[6].n48 XThR.Tn[6].t43 143.911
R17186 XThR.Tn[6].n43 XThR.Tn[6].t37 143.911
R17187 XThR.Tn[6].n38 XThR.Tn[6].t70 143.911
R17188 XThR.Tn[6].n33 XThR.Tn[6].t29 143.911
R17189 XThR.Tn[6].n28 XThR.Tn[6].t59 143.911
R17190 XThR.Tn[6].n23 XThR.Tn[6].t26 143.911
R17191 XThR.Tn[6].n18 XThR.Tn[6].t14 143.911
R17192 XThR.Tn[6].n13 XThR.Tn[6].t36 143.911
R17193 XThR.Tn[6].n7 XThR.Tn[6].n5 135.249
R17194 XThR.Tn[6].n9 XThR.Tn[6].n3 98.982
R17195 XThR.Tn[6].n8 XThR.Tn[6].n4 98.982
R17196 XThR.Tn[6].n7 XThR.Tn[6].n6 98.982
R17197 XThR.Tn[6].n9 XThR.Tn[6].n8 36.2672
R17198 XThR.Tn[6].n8 XThR.Tn[6].n7 36.2672
R17199 XThR.Tn[6].n88 XThR.Tn[6].n9 32.6405
R17200 XThR.Tn[6].n1 XThR.Tn[6].t6 26.5955
R17201 XThR.Tn[6].n1 XThR.Tn[6].t5 26.5955
R17202 XThR.Tn[6].n0 XThR.Tn[6].t7 26.5955
R17203 XThR.Tn[6].n0 XThR.Tn[6].t4 26.5955
R17204 XThR.Tn[6].n3 XThR.Tn[6].t8 24.9236
R17205 XThR.Tn[6].n3 XThR.Tn[6].t9 24.9236
R17206 XThR.Tn[6].n4 XThR.Tn[6].t11 24.9236
R17207 XThR.Tn[6].n4 XThR.Tn[6].t10 24.9236
R17208 XThR.Tn[6].n5 XThR.Tn[6].t0 24.9236
R17209 XThR.Tn[6].n5 XThR.Tn[6].t1 24.9236
R17210 XThR.Tn[6].n6 XThR.Tn[6].t3 24.9236
R17211 XThR.Tn[6].n6 XThR.Tn[6].t2 24.9236
R17212 XThR.Tn[6] XThR.Tn[6].n2 23.3605
R17213 XThR.Tn[6] XThR.Tn[6].n88 6.7205
R17214 XThR.Tn[6].n88 XThR.Tn[6] 5.37828
R17215 XThR.Tn[6] XThR.Tn[6].n11 5.34038
R17216 XThR.Tn[6].n16 XThR.Tn[6].n15 4.5005
R17217 XThR.Tn[6].n21 XThR.Tn[6].n20 4.5005
R17218 XThR.Tn[6].n26 XThR.Tn[6].n25 4.5005
R17219 XThR.Tn[6].n31 XThR.Tn[6].n30 4.5005
R17220 XThR.Tn[6].n36 XThR.Tn[6].n35 4.5005
R17221 XThR.Tn[6].n41 XThR.Tn[6].n40 4.5005
R17222 XThR.Tn[6].n46 XThR.Tn[6].n45 4.5005
R17223 XThR.Tn[6].n51 XThR.Tn[6].n50 4.5005
R17224 XThR.Tn[6].n56 XThR.Tn[6].n55 4.5005
R17225 XThR.Tn[6].n61 XThR.Tn[6].n60 4.5005
R17226 XThR.Tn[6].n66 XThR.Tn[6].n65 4.5005
R17227 XThR.Tn[6].n71 XThR.Tn[6].n70 4.5005
R17228 XThR.Tn[6].n76 XThR.Tn[6].n75 4.5005
R17229 XThR.Tn[6].n81 XThR.Tn[6].n80 4.5005
R17230 XThR.Tn[6].n86 XThR.Tn[6].n85 4.5005
R17231 XThR.Tn[6].n87 XThR.Tn[6] 3.70586
R17232 XThR.Tn[6].n16 XThR.Tn[6] 2.52282
R17233 XThR.Tn[6].n21 XThR.Tn[6] 2.52282
R17234 XThR.Tn[6].n26 XThR.Tn[6] 2.52282
R17235 XThR.Tn[6].n31 XThR.Tn[6] 2.52282
R17236 XThR.Tn[6].n36 XThR.Tn[6] 2.52282
R17237 XThR.Tn[6].n41 XThR.Tn[6] 2.52282
R17238 XThR.Tn[6].n46 XThR.Tn[6] 2.52282
R17239 XThR.Tn[6].n51 XThR.Tn[6] 2.52282
R17240 XThR.Tn[6].n56 XThR.Tn[6] 2.52282
R17241 XThR.Tn[6].n61 XThR.Tn[6] 2.52282
R17242 XThR.Tn[6].n66 XThR.Tn[6] 2.52282
R17243 XThR.Tn[6].n71 XThR.Tn[6] 2.52282
R17244 XThR.Tn[6].n76 XThR.Tn[6] 2.52282
R17245 XThR.Tn[6].n81 XThR.Tn[6] 2.52282
R17246 XThR.Tn[6].n86 XThR.Tn[6] 2.52282
R17247 XThR.Tn[6].n84 XThR.Tn[6] 1.08677
R17248 XThR.Tn[6].n79 XThR.Tn[6] 1.08677
R17249 XThR.Tn[6].n74 XThR.Tn[6] 1.08677
R17250 XThR.Tn[6].n69 XThR.Tn[6] 1.08677
R17251 XThR.Tn[6].n64 XThR.Tn[6] 1.08677
R17252 XThR.Tn[6].n59 XThR.Tn[6] 1.08677
R17253 XThR.Tn[6].n54 XThR.Tn[6] 1.08677
R17254 XThR.Tn[6].n49 XThR.Tn[6] 1.08677
R17255 XThR.Tn[6].n44 XThR.Tn[6] 1.08677
R17256 XThR.Tn[6].n39 XThR.Tn[6] 1.08677
R17257 XThR.Tn[6].n34 XThR.Tn[6] 1.08677
R17258 XThR.Tn[6].n29 XThR.Tn[6] 1.08677
R17259 XThR.Tn[6].n24 XThR.Tn[6] 1.08677
R17260 XThR.Tn[6].n19 XThR.Tn[6] 1.08677
R17261 XThR.Tn[6].n14 XThR.Tn[6] 1.08677
R17262 XThR.Tn[6] XThR.Tn[6].n16 0.839786
R17263 XThR.Tn[6] XThR.Tn[6].n21 0.839786
R17264 XThR.Tn[6] XThR.Tn[6].n26 0.839786
R17265 XThR.Tn[6] XThR.Tn[6].n31 0.839786
R17266 XThR.Tn[6] XThR.Tn[6].n36 0.839786
R17267 XThR.Tn[6] XThR.Tn[6].n41 0.839786
R17268 XThR.Tn[6] XThR.Tn[6].n46 0.839786
R17269 XThR.Tn[6] XThR.Tn[6].n51 0.839786
R17270 XThR.Tn[6] XThR.Tn[6].n56 0.839786
R17271 XThR.Tn[6] XThR.Tn[6].n61 0.839786
R17272 XThR.Tn[6] XThR.Tn[6].n66 0.839786
R17273 XThR.Tn[6] XThR.Tn[6].n71 0.839786
R17274 XThR.Tn[6] XThR.Tn[6].n76 0.839786
R17275 XThR.Tn[6] XThR.Tn[6].n81 0.839786
R17276 XThR.Tn[6] XThR.Tn[6].n86 0.839786
R17277 XThR.Tn[6].n11 XThR.Tn[6] 0.499542
R17278 XThR.Tn[6].n85 XThR.Tn[6] 0.063
R17279 XThR.Tn[6].n80 XThR.Tn[6] 0.063
R17280 XThR.Tn[6].n75 XThR.Tn[6] 0.063
R17281 XThR.Tn[6].n70 XThR.Tn[6] 0.063
R17282 XThR.Tn[6].n65 XThR.Tn[6] 0.063
R17283 XThR.Tn[6].n60 XThR.Tn[6] 0.063
R17284 XThR.Tn[6].n55 XThR.Tn[6] 0.063
R17285 XThR.Tn[6].n50 XThR.Tn[6] 0.063
R17286 XThR.Tn[6].n45 XThR.Tn[6] 0.063
R17287 XThR.Tn[6].n40 XThR.Tn[6] 0.063
R17288 XThR.Tn[6].n35 XThR.Tn[6] 0.063
R17289 XThR.Tn[6].n30 XThR.Tn[6] 0.063
R17290 XThR.Tn[6].n25 XThR.Tn[6] 0.063
R17291 XThR.Tn[6].n20 XThR.Tn[6] 0.063
R17292 XThR.Tn[6].n15 XThR.Tn[6] 0.063
R17293 XThR.Tn[6].n87 XThR.Tn[6] 0.0540714
R17294 XThR.Tn[6] XThR.Tn[6].n87 0.038
R17295 XThR.Tn[6].n11 XThR.Tn[6] 0.0143889
R17296 XThR.Tn[6].n85 XThR.Tn[6].n84 0.00771154
R17297 XThR.Tn[6].n80 XThR.Tn[6].n79 0.00771154
R17298 XThR.Tn[6].n75 XThR.Tn[6].n74 0.00771154
R17299 XThR.Tn[6].n70 XThR.Tn[6].n69 0.00771154
R17300 XThR.Tn[6].n65 XThR.Tn[6].n64 0.00771154
R17301 XThR.Tn[6].n60 XThR.Tn[6].n59 0.00771154
R17302 XThR.Tn[6].n55 XThR.Tn[6].n54 0.00771154
R17303 XThR.Tn[6].n50 XThR.Tn[6].n49 0.00771154
R17304 XThR.Tn[6].n45 XThR.Tn[6].n44 0.00771154
R17305 XThR.Tn[6].n40 XThR.Tn[6].n39 0.00771154
R17306 XThR.Tn[6].n35 XThR.Tn[6].n34 0.00771154
R17307 XThR.Tn[6].n30 XThR.Tn[6].n29 0.00771154
R17308 XThR.Tn[6].n25 XThR.Tn[6].n24 0.00771154
R17309 XThR.Tn[6].n20 XThR.Tn[6].n19 0.00771154
R17310 XThR.Tn[6].n15 XThR.Tn[6].n14 0.00771154
R17311 XThR.Tn[14].n5 XThR.Tn[14].n4 256.103
R17312 XThR.Tn[14].n2 XThR.Tn[14].n0 243.68
R17313 XThR.Tn[14].n88 XThR.Tn[14].n87 241.847
R17314 XThR.Tn[14].n2 XThR.Tn[14].n1 205.28
R17315 XThR.Tn[14].n5 XThR.Tn[14].n3 202.095
R17316 XThR.Tn[14].n88 XThR.Tn[14].n86 185
R17317 XThR.Tn[14] XThR.Tn[14].n79 161.363
R17318 XThR.Tn[14] XThR.Tn[14].n74 161.363
R17319 XThR.Tn[14] XThR.Tn[14].n69 161.363
R17320 XThR.Tn[14] XThR.Tn[14].n64 161.363
R17321 XThR.Tn[14] XThR.Tn[14].n59 161.363
R17322 XThR.Tn[14] XThR.Tn[14].n54 161.363
R17323 XThR.Tn[14] XThR.Tn[14].n49 161.363
R17324 XThR.Tn[14] XThR.Tn[14].n44 161.363
R17325 XThR.Tn[14] XThR.Tn[14].n39 161.363
R17326 XThR.Tn[14] XThR.Tn[14].n34 161.363
R17327 XThR.Tn[14] XThR.Tn[14].n29 161.363
R17328 XThR.Tn[14] XThR.Tn[14].n24 161.363
R17329 XThR.Tn[14] XThR.Tn[14].n19 161.363
R17330 XThR.Tn[14] XThR.Tn[14].n14 161.363
R17331 XThR.Tn[14] XThR.Tn[14].n9 161.363
R17332 XThR.Tn[14] XThR.Tn[14].n7 161.363
R17333 XThR.Tn[14].n81 XThR.Tn[14].n80 161.3
R17334 XThR.Tn[14].n76 XThR.Tn[14].n75 161.3
R17335 XThR.Tn[14].n71 XThR.Tn[14].n70 161.3
R17336 XThR.Tn[14].n66 XThR.Tn[14].n65 161.3
R17337 XThR.Tn[14].n61 XThR.Tn[14].n60 161.3
R17338 XThR.Tn[14].n56 XThR.Tn[14].n55 161.3
R17339 XThR.Tn[14].n51 XThR.Tn[14].n50 161.3
R17340 XThR.Tn[14].n46 XThR.Tn[14].n45 161.3
R17341 XThR.Tn[14].n41 XThR.Tn[14].n40 161.3
R17342 XThR.Tn[14].n36 XThR.Tn[14].n35 161.3
R17343 XThR.Tn[14].n31 XThR.Tn[14].n30 161.3
R17344 XThR.Tn[14].n26 XThR.Tn[14].n25 161.3
R17345 XThR.Tn[14].n21 XThR.Tn[14].n20 161.3
R17346 XThR.Tn[14].n16 XThR.Tn[14].n15 161.3
R17347 XThR.Tn[14].n11 XThR.Tn[14].n10 161.3
R17348 XThR.Tn[14].n79 XThR.Tn[14].t51 161.106
R17349 XThR.Tn[14].n74 XThR.Tn[14].t58 161.106
R17350 XThR.Tn[14].n69 XThR.Tn[14].t39 161.106
R17351 XThR.Tn[14].n64 XThR.Tn[14].t22 161.106
R17352 XThR.Tn[14].n59 XThR.Tn[14].t49 161.106
R17353 XThR.Tn[14].n54 XThR.Tn[14].t12 161.106
R17354 XThR.Tn[14].n49 XThR.Tn[14].t56 161.106
R17355 XThR.Tn[14].n44 XThR.Tn[14].t36 161.106
R17356 XThR.Tn[14].n39 XThR.Tn[14].t19 161.106
R17357 XThR.Tn[14].n34 XThR.Tn[14].t25 161.106
R17358 XThR.Tn[14].n29 XThR.Tn[14].t73 161.106
R17359 XThR.Tn[14].n24 XThR.Tn[14].t38 161.106
R17360 XThR.Tn[14].n19 XThR.Tn[14].t72 161.106
R17361 XThR.Tn[14].n14 XThR.Tn[14].t54 161.106
R17362 XThR.Tn[14].n9 XThR.Tn[14].t13 161.106
R17363 XThR.Tn[14].n7 XThR.Tn[14].t62 161.106
R17364 XThR.Tn[14].n80 XThR.Tn[14].t32 159.978
R17365 XThR.Tn[14].n75 XThR.Tn[14].t37 159.978
R17366 XThR.Tn[14].n70 XThR.Tn[14].t20 159.978
R17367 XThR.Tn[14].n65 XThR.Tn[14].t68 159.978
R17368 XThR.Tn[14].n60 XThR.Tn[14].t30 159.978
R17369 XThR.Tn[14].n55 XThR.Tn[14].t55 159.978
R17370 XThR.Tn[14].n50 XThR.Tn[14].t35 159.978
R17371 XThR.Tn[14].n45 XThR.Tn[14].t16 159.978
R17372 XThR.Tn[14].n40 XThR.Tn[14].t66 159.978
R17373 XThR.Tn[14].n35 XThR.Tn[14].t71 159.978
R17374 XThR.Tn[14].n30 XThR.Tn[14].t53 159.978
R17375 XThR.Tn[14].n25 XThR.Tn[14].t18 159.978
R17376 XThR.Tn[14].n20 XThR.Tn[14].t52 159.978
R17377 XThR.Tn[14].n15 XThR.Tn[14].t34 159.978
R17378 XThR.Tn[14].n10 XThR.Tn[14].t60 159.978
R17379 XThR.Tn[14].n79 XThR.Tn[14].t41 145.038
R17380 XThR.Tn[14].n74 XThR.Tn[14].t65 145.038
R17381 XThR.Tn[14].n69 XThR.Tn[14].t45 145.038
R17382 XThR.Tn[14].n64 XThR.Tn[14].t26 145.038
R17383 XThR.Tn[14].n59 XThR.Tn[14].t59 145.038
R17384 XThR.Tn[14].n54 XThR.Tn[14].t40 145.038
R17385 XThR.Tn[14].n49 XThR.Tn[14].t46 145.038
R17386 XThR.Tn[14].n44 XThR.Tn[14].t27 145.038
R17387 XThR.Tn[14].n39 XThR.Tn[14].t23 145.038
R17388 XThR.Tn[14].n34 XThR.Tn[14].t57 145.038
R17389 XThR.Tn[14].n29 XThR.Tn[14].t15 145.038
R17390 XThR.Tn[14].n24 XThR.Tn[14].t44 145.038
R17391 XThR.Tn[14].n19 XThR.Tn[14].t14 145.038
R17392 XThR.Tn[14].n14 XThR.Tn[14].t64 145.038
R17393 XThR.Tn[14].n9 XThR.Tn[14].t24 145.038
R17394 XThR.Tn[14].n7 XThR.Tn[14].t69 145.038
R17395 XThR.Tn[14].n80 XThR.Tn[14].t43 143.911
R17396 XThR.Tn[14].n75 XThR.Tn[14].t70 143.911
R17397 XThR.Tn[14].n70 XThR.Tn[14].t48 143.911
R17398 XThR.Tn[14].n65 XThR.Tn[14].t31 143.911
R17399 XThR.Tn[14].n60 XThR.Tn[14].t63 143.911
R17400 XThR.Tn[14].n55 XThR.Tn[14].t42 143.911
R17401 XThR.Tn[14].n50 XThR.Tn[14].t50 143.911
R17402 XThR.Tn[14].n45 XThR.Tn[14].t33 143.911
R17403 XThR.Tn[14].n40 XThR.Tn[14].t29 143.911
R17404 XThR.Tn[14].n35 XThR.Tn[14].t61 143.911
R17405 XThR.Tn[14].n30 XThR.Tn[14].t21 143.911
R17406 XThR.Tn[14].n25 XThR.Tn[14].t47 143.911
R17407 XThR.Tn[14].n20 XThR.Tn[14].t17 143.911
R17408 XThR.Tn[14].n15 XThR.Tn[14].t67 143.911
R17409 XThR.Tn[14].n10 XThR.Tn[14].t28 143.911
R17410 XThR.Tn[14] XThR.Tn[14].n2 35.7652
R17411 XThR.Tn[14].n3 XThR.Tn[14].t6 26.5955
R17412 XThR.Tn[14].n3 XThR.Tn[14].t7 26.5955
R17413 XThR.Tn[14].n4 XThR.Tn[14].t4 26.5955
R17414 XThR.Tn[14].n4 XThR.Tn[14].t5 26.5955
R17415 XThR.Tn[14].n0 XThR.Tn[14].t8 26.5955
R17416 XThR.Tn[14].n0 XThR.Tn[14].t9 26.5955
R17417 XThR.Tn[14].n1 XThR.Tn[14].t10 26.5955
R17418 XThR.Tn[14].n1 XThR.Tn[14].t11 26.5955
R17419 XThR.Tn[14].n86 XThR.Tn[14].t0 24.9236
R17420 XThR.Tn[14].n86 XThR.Tn[14].t1 24.9236
R17421 XThR.Tn[14].n87 XThR.Tn[14].t2 24.9236
R17422 XThR.Tn[14].n87 XThR.Tn[14].t3 24.9236
R17423 XThR.Tn[14] XThR.Tn[14].n88 18.8943
R17424 XThR.Tn[14].n6 XThR.Tn[14].n5 13.5534
R17425 XThR.Tn[14].n85 XThR.Tn[14] 8.47191
R17426 XThR.Tn[14] XThR.Tn[14].n85 6.34069
R17427 XThR.Tn[14] XThR.Tn[14].n8 5.34038
R17428 XThR.Tn[14].n13 XThR.Tn[14].n12 4.5005
R17429 XThR.Tn[14].n18 XThR.Tn[14].n17 4.5005
R17430 XThR.Tn[14].n23 XThR.Tn[14].n22 4.5005
R17431 XThR.Tn[14].n28 XThR.Tn[14].n27 4.5005
R17432 XThR.Tn[14].n33 XThR.Tn[14].n32 4.5005
R17433 XThR.Tn[14].n38 XThR.Tn[14].n37 4.5005
R17434 XThR.Tn[14].n43 XThR.Tn[14].n42 4.5005
R17435 XThR.Tn[14].n48 XThR.Tn[14].n47 4.5005
R17436 XThR.Tn[14].n53 XThR.Tn[14].n52 4.5005
R17437 XThR.Tn[14].n58 XThR.Tn[14].n57 4.5005
R17438 XThR.Tn[14].n63 XThR.Tn[14].n62 4.5005
R17439 XThR.Tn[14].n68 XThR.Tn[14].n67 4.5005
R17440 XThR.Tn[14].n73 XThR.Tn[14].n72 4.5005
R17441 XThR.Tn[14].n78 XThR.Tn[14].n77 4.5005
R17442 XThR.Tn[14].n83 XThR.Tn[14].n82 4.5005
R17443 XThR.Tn[14].n84 XThR.Tn[14] 3.70586
R17444 XThR.Tn[14].n13 XThR.Tn[14] 2.52282
R17445 XThR.Tn[14].n18 XThR.Tn[14] 2.52282
R17446 XThR.Tn[14].n23 XThR.Tn[14] 2.52282
R17447 XThR.Tn[14].n28 XThR.Tn[14] 2.52282
R17448 XThR.Tn[14].n33 XThR.Tn[14] 2.52282
R17449 XThR.Tn[14].n38 XThR.Tn[14] 2.52282
R17450 XThR.Tn[14].n43 XThR.Tn[14] 2.52282
R17451 XThR.Tn[14].n48 XThR.Tn[14] 2.52282
R17452 XThR.Tn[14].n53 XThR.Tn[14] 2.52282
R17453 XThR.Tn[14].n58 XThR.Tn[14] 2.52282
R17454 XThR.Tn[14].n63 XThR.Tn[14] 2.52282
R17455 XThR.Tn[14].n68 XThR.Tn[14] 2.52282
R17456 XThR.Tn[14].n73 XThR.Tn[14] 2.52282
R17457 XThR.Tn[14].n78 XThR.Tn[14] 2.52282
R17458 XThR.Tn[14].n83 XThR.Tn[14] 2.52282
R17459 XThR.Tn[14].n85 XThR.Tn[14] 1.79489
R17460 XThR.Tn[14].n6 XThR.Tn[14] 1.50638
R17461 XThR.Tn[14] XThR.Tn[14].n6 1.19676
R17462 XThR.Tn[14].n81 XThR.Tn[14] 1.08677
R17463 XThR.Tn[14].n76 XThR.Tn[14] 1.08677
R17464 XThR.Tn[14].n71 XThR.Tn[14] 1.08677
R17465 XThR.Tn[14].n66 XThR.Tn[14] 1.08677
R17466 XThR.Tn[14].n61 XThR.Tn[14] 1.08677
R17467 XThR.Tn[14].n56 XThR.Tn[14] 1.08677
R17468 XThR.Tn[14].n51 XThR.Tn[14] 1.08677
R17469 XThR.Tn[14].n46 XThR.Tn[14] 1.08677
R17470 XThR.Tn[14].n41 XThR.Tn[14] 1.08677
R17471 XThR.Tn[14].n36 XThR.Tn[14] 1.08677
R17472 XThR.Tn[14].n31 XThR.Tn[14] 1.08677
R17473 XThR.Tn[14].n26 XThR.Tn[14] 1.08677
R17474 XThR.Tn[14].n21 XThR.Tn[14] 1.08677
R17475 XThR.Tn[14].n16 XThR.Tn[14] 1.08677
R17476 XThR.Tn[14].n11 XThR.Tn[14] 1.08677
R17477 XThR.Tn[14] XThR.Tn[14].n13 0.839786
R17478 XThR.Tn[14] XThR.Tn[14].n18 0.839786
R17479 XThR.Tn[14] XThR.Tn[14].n23 0.839786
R17480 XThR.Tn[14] XThR.Tn[14].n28 0.839786
R17481 XThR.Tn[14] XThR.Tn[14].n33 0.839786
R17482 XThR.Tn[14] XThR.Tn[14].n38 0.839786
R17483 XThR.Tn[14] XThR.Tn[14].n43 0.839786
R17484 XThR.Tn[14] XThR.Tn[14].n48 0.839786
R17485 XThR.Tn[14] XThR.Tn[14].n53 0.839786
R17486 XThR.Tn[14] XThR.Tn[14].n58 0.839786
R17487 XThR.Tn[14] XThR.Tn[14].n63 0.839786
R17488 XThR.Tn[14] XThR.Tn[14].n68 0.839786
R17489 XThR.Tn[14] XThR.Tn[14].n73 0.839786
R17490 XThR.Tn[14] XThR.Tn[14].n78 0.839786
R17491 XThR.Tn[14] XThR.Tn[14].n83 0.839786
R17492 XThR.Tn[14].n8 XThR.Tn[14] 0.499542
R17493 XThR.Tn[14].n82 XThR.Tn[14] 0.063
R17494 XThR.Tn[14].n77 XThR.Tn[14] 0.063
R17495 XThR.Tn[14].n72 XThR.Tn[14] 0.063
R17496 XThR.Tn[14].n67 XThR.Tn[14] 0.063
R17497 XThR.Tn[14].n62 XThR.Tn[14] 0.063
R17498 XThR.Tn[14].n57 XThR.Tn[14] 0.063
R17499 XThR.Tn[14].n52 XThR.Tn[14] 0.063
R17500 XThR.Tn[14].n47 XThR.Tn[14] 0.063
R17501 XThR.Tn[14].n42 XThR.Tn[14] 0.063
R17502 XThR.Tn[14].n37 XThR.Tn[14] 0.063
R17503 XThR.Tn[14].n32 XThR.Tn[14] 0.063
R17504 XThR.Tn[14].n27 XThR.Tn[14] 0.063
R17505 XThR.Tn[14].n22 XThR.Tn[14] 0.063
R17506 XThR.Tn[14].n17 XThR.Tn[14] 0.063
R17507 XThR.Tn[14].n12 XThR.Tn[14] 0.063
R17508 XThR.Tn[14].n84 XThR.Tn[14] 0.0540714
R17509 XThR.Tn[14] XThR.Tn[14].n84 0.038
R17510 XThR.Tn[14].n8 XThR.Tn[14] 0.0143889
R17511 XThR.Tn[14].n82 XThR.Tn[14].n81 0.00771154
R17512 XThR.Tn[14].n77 XThR.Tn[14].n76 0.00771154
R17513 XThR.Tn[14].n72 XThR.Tn[14].n71 0.00771154
R17514 XThR.Tn[14].n67 XThR.Tn[14].n66 0.00771154
R17515 XThR.Tn[14].n62 XThR.Tn[14].n61 0.00771154
R17516 XThR.Tn[14].n57 XThR.Tn[14].n56 0.00771154
R17517 XThR.Tn[14].n52 XThR.Tn[14].n51 0.00771154
R17518 XThR.Tn[14].n47 XThR.Tn[14].n46 0.00771154
R17519 XThR.Tn[14].n42 XThR.Tn[14].n41 0.00771154
R17520 XThR.Tn[14].n37 XThR.Tn[14].n36 0.00771154
R17521 XThR.Tn[14].n32 XThR.Tn[14].n31 0.00771154
R17522 XThR.Tn[14].n27 XThR.Tn[14].n26 0.00771154
R17523 XThR.Tn[14].n22 XThR.Tn[14].n21 0.00771154
R17524 XThR.Tn[14].n17 XThR.Tn[14].n16 0.00771154
R17525 XThR.Tn[14].n12 XThR.Tn[14].n11 0.00771154
R17526 XThR.Tn[12].n5 XThR.Tn[12].n4 256.103
R17527 XThR.Tn[12].n2 XThR.Tn[12].n0 243.68
R17528 XThR.Tn[12].n88 XThR.Tn[12].n87 241.847
R17529 XThR.Tn[12].n2 XThR.Tn[12].n1 205.28
R17530 XThR.Tn[12].n5 XThR.Tn[12].n3 202.095
R17531 XThR.Tn[12].n88 XThR.Tn[12].n86 185
R17532 XThR.Tn[12] XThR.Tn[12].n79 161.363
R17533 XThR.Tn[12] XThR.Tn[12].n74 161.363
R17534 XThR.Tn[12] XThR.Tn[12].n69 161.363
R17535 XThR.Tn[12] XThR.Tn[12].n64 161.363
R17536 XThR.Tn[12] XThR.Tn[12].n59 161.363
R17537 XThR.Tn[12] XThR.Tn[12].n54 161.363
R17538 XThR.Tn[12] XThR.Tn[12].n49 161.363
R17539 XThR.Tn[12] XThR.Tn[12].n44 161.363
R17540 XThR.Tn[12] XThR.Tn[12].n39 161.363
R17541 XThR.Tn[12] XThR.Tn[12].n34 161.363
R17542 XThR.Tn[12] XThR.Tn[12].n29 161.363
R17543 XThR.Tn[12] XThR.Tn[12].n24 161.363
R17544 XThR.Tn[12] XThR.Tn[12].n19 161.363
R17545 XThR.Tn[12] XThR.Tn[12].n14 161.363
R17546 XThR.Tn[12] XThR.Tn[12].n9 161.363
R17547 XThR.Tn[12] XThR.Tn[12].n7 161.363
R17548 XThR.Tn[12].n81 XThR.Tn[12].n80 161.3
R17549 XThR.Tn[12].n76 XThR.Tn[12].n75 161.3
R17550 XThR.Tn[12].n71 XThR.Tn[12].n70 161.3
R17551 XThR.Tn[12].n66 XThR.Tn[12].n65 161.3
R17552 XThR.Tn[12].n61 XThR.Tn[12].n60 161.3
R17553 XThR.Tn[12].n56 XThR.Tn[12].n55 161.3
R17554 XThR.Tn[12].n51 XThR.Tn[12].n50 161.3
R17555 XThR.Tn[12].n46 XThR.Tn[12].n45 161.3
R17556 XThR.Tn[12].n41 XThR.Tn[12].n40 161.3
R17557 XThR.Tn[12].n36 XThR.Tn[12].n35 161.3
R17558 XThR.Tn[12].n31 XThR.Tn[12].n30 161.3
R17559 XThR.Tn[12].n26 XThR.Tn[12].n25 161.3
R17560 XThR.Tn[12].n21 XThR.Tn[12].n20 161.3
R17561 XThR.Tn[12].n16 XThR.Tn[12].n15 161.3
R17562 XThR.Tn[12].n11 XThR.Tn[12].n10 161.3
R17563 XThR.Tn[12].n79 XThR.Tn[12].t18 161.106
R17564 XThR.Tn[12].n74 XThR.Tn[12].t24 161.106
R17565 XThR.Tn[12].n69 XThR.Tn[12].t67 161.106
R17566 XThR.Tn[12].n64 XThR.Tn[12].t52 161.106
R17567 XThR.Tn[12].n59 XThR.Tn[12].t16 161.106
R17568 XThR.Tn[12].n54 XThR.Tn[12].t40 161.106
R17569 XThR.Tn[12].n49 XThR.Tn[12].t22 161.106
R17570 XThR.Tn[12].n44 XThR.Tn[12].t65 161.106
R17571 XThR.Tn[12].n39 XThR.Tn[12].t51 161.106
R17572 XThR.Tn[12].n34 XThR.Tn[12].t56 161.106
R17573 XThR.Tn[12].n29 XThR.Tn[12].t39 161.106
R17574 XThR.Tn[12].n24 XThR.Tn[12].t66 161.106
R17575 XThR.Tn[12].n19 XThR.Tn[12].t38 161.106
R17576 XThR.Tn[12].n14 XThR.Tn[12].t20 161.106
R17577 XThR.Tn[12].n9 XThR.Tn[12].t43 161.106
R17578 XThR.Tn[12].n7 XThR.Tn[12].t28 161.106
R17579 XThR.Tn[12].n80 XThR.Tn[12].t58 159.978
R17580 XThR.Tn[12].n75 XThR.Tn[12].t62 159.978
R17581 XThR.Tn[12].n70 XThR.Tn[12].t47 159.978
R17582 XThR.Tn[12].n65 XThR.Tn[12].t31 159.978
R17583 XThR.Tn[12].n60 XThR.Tn[12].t55 159.978
R17584 XThR.Tn[12].n55 XThR.Tn[12].t19 159.978
R17585 XThR.Tn[12].n50 XThR.Tn[12].t61 159.978
R17586 XThR.Tn[12].n45 XThR.Tn[12].t44 159.978
R17587 XThR.Tn[12].n40 XThR.Tn[12].t29 159.978
R17588 XThR.Tn[12].n35 XThR.Tn[12].t37 159.978
R17589 XThR.Tn[12].n30 XThR.Tn[12].t17 159.978
R17590 XThR.Tn[12].n25 XThR.Tn[12].t46 159.978
R17591 XThR.Tn[12].n20 XThR.Tn[12].t15 159.978
R17592 XThR.Tn[12].n15 XThR.Tn[12].t60 159.978
R17593 XThR.Tn[12].n10 XThR.Tn[12].t21 159.978
R17594 XThR.Tn[12].n79 XThR.Tn[12].t69 145.038
R17595 XThR.Tn[12].n74 XThR.Tn[12].t32 145.038
R17596 XThR.Tn[12].n69 XThR.Tn[12].t73 145.038
R17597 XThR.Tn[12].n64 XThR.Tn[12].t57 145.038
R17598 XThR.Tn[12].n59 XThR.Tn[12].t25 145.038
R17599 XThR.Tn[12].n54 XThR.Tn[12].t68 145.038
R17600 XThR.Tn[12].n49 XThR.Tn[12].t12 145.038
R17601 XThR.Tn[12].n44 XThR.Tn[12].t59 145.038
R17602 XThR.Tn[12].n39 XThR.Tn[12].t54 145.038
R17603 XThR.Tn[12].n34 XThR.Tn[12].t23 145.038
R17604 XThR.Tn[12].n29 XThR.Tn[12].t48 145.038
R17605 XThR.Tn[12].n24 XThR.Tn[12].t70 145.038
R17606 XThR.Tn[12].n19 XThR.Tn[12].t45 145.038
R17607 XThR.Tn[12].n14 XThR.Tn[12].t30 145.038
R17608 XThR.Tn[12].n9 XThR.Tn[12].t53 145.038
R17609 XThR.Tn[12].n7 XThR.Tn[12].t36 145.038
R17610 XThR.Tn[12].n80 XThR.Tn[12].t27 143.911
R17611 XThR.Tn[12].n75 XThR.Tn[12].t50 143.911
R17612 XThR.Tn[12].n70 XThR.Tn[12].t34 143.911
R17613 XThR.Tn[12].n65 XThR.Tn[12].t13 143.911
R17614 XThR.Tn[12].n60 XThR.Tn[12].t42 143.911
R17615 XThR.Tn[12].n55 XThR.Tn[12].t26 143.911
R17616 XThR.Tn[12].n50 XThR.Tn[12].t35 143.911
R17617 XThR.Tn[12].n45 XThR.Tn[12].t14 143.911
R17618 XThR.Tn[12].n40 XThR.Tn[12].t72 143.911
R17619 XThR.Tn[12].n35 XThR.Tn[12].t41 143.911
R17620 XThR.Tn[12].n30 XThR.Tn[12].t64 143.911
R17621 XThR.Tn[12].n25 XThR.Tn[12].t33 143.911
R17622 XThR.Tn[12].n20 XThR.Tn[12].t63 143.911
R17623 XThR.Tn[12].n15 XThR.Tn[12].t49 143.911
R17624 XThR.Tn[12].n10 XThR.Tn[12].t71 143.911
R17625 XThR.Tn[12] XThR.Tn[12].n2 35.7652
R17626 XThR.Tn[12].n3 XThR.Tn[12].t6 26.5955
R17627 XThR.Tn[12].n3 XThR.Tn[12].t4 26.5955
R17628 XThR.Tn[12].n4 XThR.Tn[12].t7 26.5955
R17629 XThR.Tn[12].n4 XThR.Tn[12].t5 26.5955
R17630 XThR.Tn[12].n0 XThR.Tn[12].t11 26.5955
R17631 XThR.Tn[12].n0 XThR.Tn[12].t9 26.5955
R17632 XThR.Tn[12].n1 XThR.Tn[12].t8 26.5955
R17633 XThR.Tn[12].n1 XThR.Tn[12].t10 26.5955
R17634 XThR.Tn[12].n86 XThR.Tn[12].t2 24.9236
R17635 XThR.Tn[12].n86 XThR.Tn[12].t0 24.9236
R17636 XThR.Tn[12].n87 XThR.Tn[12].t3 24.9236
R17637 XThR.Tn[12].n87 XThR.Tn[12].t1 24.9236
R17638 XThR.Tn[12] XThR.Tn[12].n88 18.8943
R17639 XThR.Tn[12].n6 XThR.Tn[12].n5 13.5534
R17640 XThR.Tn[12].n85 XThR.Tn[12] 8.18715
R17641 XThR.Tn[12] XThR.Tn[12].n85 6.34069
R17642 XThR.Tn[12] XThR.Tn[12].n8 5.34038
R17643 XThR.Tn[12].n13 XThR.Tn[12].n12 4.5005
R17644 XThR.Tn[12].n18 XThR.Tn[12].n17 4.5005
R17645 XThR.Tn[12].n23 XThR.Tn[12].n22 4.5005
R17646 XThR.Tn[12].n28 XThR.Tn[12].n27 4.5005
R17647 XThR.Tn[12].n33 XThR.Tn[12].n32 4.5005
R17648 XThR.Tn[12].n38 XThR.Tn[12].n37 4.5005
R17649 XThR.Tn[12].n43 XThR.Tn[12].n42 4.5005
R17650 XThR.Tn[12].n48 XThR.Tn[12].n47 4.5005
R17651 XThR.Tn[12].n53 XThR.Tn[12].n52 4.5005
R17652 XThR.Tn[12].n58 XThR.Tn[12].n57 4.5005
R17653 XThR.Tn[12].n63 XThR.Tn[12].n62 4.5005
R17654 XThR.Tn[12].n68 XThR.Tn[12].n67 4.5005
R17655 XThR.Tn[12].n73 XThR.Tn[12].n72 4.5005
R17656 XThR.Tn[12].n78 XThR.Tn[12].n77 4.5005
R17657 XThR.Tn[12].n83 XThR.Tn[12].n82 4.5005
R17658 XThR.Tn[12].n84 XThR.Tn[12] 3.70586
R17659 XThR.Tn[12].n13 XThR.Tn[12] 2.52282
R17660 XThR.Tn[12].n18 XThR.Tn[12] 2.52282
R17661 XThR.Tn[12].n23 XThR.Tn[12] 2.52282
R17662 XThR.Tn[12].n28 XThR.Tn[12] 2.52282
R17663 XThR.Tn[12].n33 XThR.Tn[12] 2.52282
R17664 XThR.Tn[12].n38 XThR.Tn[12] 2.52282
R17665 XThR.Tn[12].n43 XThR.Tn[12] 2.52282
R17666 XThR.Tn[12].n48 XThR.Tn[12] 2.52282
R17667 XThR.Tn[12].n53 XThR.Tn[12] 2.52282
R17668 XThR.Tn[12].n58 XThR.Tn[12] 2.52282
R17669 XThR.Tn[12].n63 XThR.Tn[12] 2.52282
R17670 XThR.Tn[12].n68 XThR.Tn[12] 2.52282
R17671 XThR.Tn[12].n73 XThR.Tn[12] 2.52282
R17672 XThR.Tn[12].n78 XThR.Tn[12] 2.52282
R17673 XThR.Tn[12].n83 XThR.Tn[12] 2.52282
R17674 XThR.Tn[12].n85 XThR.Tn[12] 1.79489
R17675 XThR.Tn[12].n6 XThR.Tn[12] 1.50638
R17676 XThR.Tn[12] XThR.Tn[12].n6 1.19676
R17677 XThR.Tn[12].n81 XThR.Tn[12] 1.08677
R17678 XThR.Tn[12].n76 XThR.Tn[12] 1.08677
R17679 XThR.Tn[12].n71 XThR.Tn[12] 1.08677
R17680 XThR.Tn[12].n66 XThR.Tn[12] 1.08677
R17681 XThR.Tn[12].n61 XThR.Tn[12] 1.08677
R17682 XThR.Tn[12].n56 XThR.Tn[12] 1.08677
R17683 XThR.Tn[12].n51 XThR.Tn[12] 1.08677
R17684 XThR.Tn[12].n46 XThR.Tn[12] 1.08677
R17685 XThR.Tn[12].n41 XThR.Tn[12] 1.08677
R17686 XThR.Tn[12].n36 XThR.Tn[12] 1.08677
R17687 XThR.Tn[12].n31 XThR.Tn[12] 1.08677
R17688 XThR.Tn[12].n26 XThR.Tn[12] 1.08677
R17689 XThR.Tn[12].n21 XThR.Tn[12] 1.08677
R17690 XThR.Tn[12].n16 XThR.Tn[12] 1.08677
R17691 XThR.Tn[12].n11 XThR.Tn[12] 1.08677
R17692 XThR.Tn[12] XThR.Tn[12].n13 0.839786
R17693 XThR.Tn[12] XThR.Tn[12].n18 0.839786
R17694 XThR.Tn[12] XThR.Tn[12].n23 0.839786
R17695 XThR.Tn[12] XThR.Tn[12].n28 0.839786
R17696 XThR.Tn[12] XThR.Tn[12].n33 0.839786
R17697 XThR.Tn[12] XThR.Tn[12].n38 0.839786
R17698 XThR.Tn[12] XThR.Tn[12].n43 0.839786
R17699 XThR.Tn[12] XThR.Tn[12].n48 0.839786
R17700 XThR.Tn[12] XThR.Tn[12].n53 0.839786
R17701 XThR.Tn[12] XThR.Tn[12].n58 0.839786
R17702 XThR.Tn[12] XThR.Tn[12].n63 0.839786
R17703 XThR.Tn[12] XThR.Tn[12].n68 0.839786
R17704 XThR.Tn[12] XThR.Tn[12].n73 0.839786
R17705 XThR.Tn[12] XThR.Tn[12].n78 0.839786
R17706 XThR.Tn[12] XThR.Tn[12].n83 0.839786
R17707 XThR.Tn[12].n8 XThR.Tn[12] 0.499542
R17708 XThR.Tn[12].n82 XThR.Tn[12] 0.063
R17709 XThR.Tn[12].n77 XThR.Tn[12] 0.063
R17710 XThR.Tn[12].n72 XThR.Tn[12] 0.063
R17711 XThR.Tn[12].n67 XThR.Tn[12] 0.063
R17712 XThR.Tn[12].n62 XThR.Tn[12] 0.063
R17713 XThR.Tn[12].n57 XThR.Tn[12] 0.063
R17714 XThR.Tn[12].n52 XThR.Tn[12] 0.063
R17715 XThR.Tn[12].n47 XThR.Tn[12] 0.063
R17716 XThR.Tn[12].n42 XThR.Tn[12] 0.063
R17717 XThR.Tn[12].n37 XThR.Tn[12] 0.063
R17718 XThR.Tn[12].n32 XThR.Tn[12] 0.063
R17719 XThR.Tn[12].n27 XThR.Tn[12] 0.063
R17720 XThR.Tn[12].n22 XThR.Tn[12] 0.063
R17721 XThR.Tn[12].n17 XThR.Tn[12] 0.063
R17722 XThR.Tn[12].n12 XThR.Tn[12] 0.063
R17723 XThR.Tn[12].n84 XThR.Tn[12] 0.0540714
R17724 XThR.Tn[12] XThR.Tn[12].n84 0.038
R17725 XThR.Tn[12].n8 XThR.Tn[12] 0.0143889
R17726 XThR.Tn[12].n82 XThR.Tn[12].n81 0.00771154
R17727 XThR.Tn[12].n77 XThR.Tn[12].n76 0.00771154
R17728 XThR.Tn[12].n72 XThR.Tn[12].n71 0.00771154
R17729 XThR.Tn[12].n67 XThR.Tn[12].n66 0.00771154
R17730 XThR.Tn[12].n62 XThR.Tn[12].n61 0.00771154
R17731 XThR.Tn[12].n57 XThR.Tn[12].n56 0.00771154
R17732 XThR.Tn[12].n52 XThR.Tn[12].n51 0.00771154
R17733 XThR.Tn[12].n47 XThR.Tn[12].n46 0.00771154
R17734 XThR.Tn[12].n42 XThR.Tn[12].n41 0.00771154
R17735 XThR.Tn[12].n37 XThR.Tn[12].n36 0.00771154
R17736 XThR.Tn[12].n32 XThR.Tn[12].n31 0.00771154
R17737 XThR.Tn[12].n27 XThR.Tn[12].n26 0.00771154
R17738 XThR.Tn[12].n22 XThR.Tn[12].n21 0.00771154
R17739 XThR.Tn[12].n17 XThR.Tn[12].n16 0.00771154
R17740 XThR.Tn[12].n12 XThR.Tn[12].n11 0.00771154
R17741 XThC.XTBN.Y.n182 XThC.XTBN.Y.t9 212.081
R17742 XThC.XTBN.Y.n181 XThC.XTBN.Y.t75 212.081
R17743 XThC.XTBN.Y.n175 XThC.XTBN.Y.t33 212.081
R17744 XThC.XTBN.Y.n176 XThC.XTBN.Y.t27 212.081
R17745 XThC.XTBN.Y.n87 XThC.XTBN.Y.t25 212.081
R17746 XThC.XTBN.Y.n78 XThC.XTBN.Y.t100 212.081
R17747 XThC.XTBN.Y.n82 XThC.XTBN.Y.t93 212.081
R17748 XThC.XTBN.Y.n80 XThC.XTBN.Y.t90 212.081
R17749 XThC.XTBN.Y.n61 XThC.XTBN.Y.t47 212.081
R17750 XThC.XTBN.Y.n52 XThC.XTBN.Y.t17 212.081
R17751 XThC.XTBN.Y.n56 XThC.XTBN.Y.t116 212.081
R17752 XThC.XTBN.Y.n54 XThC.XTBN.Y.t111 212.081
R17753 XThC.XTBN.Y.n35 XThC.XTBN.Y.t106 212.081
R17754 XThC.XTBN.Y.n26 XThC.XTBN.Y.t70 212.081
R17755 XThC.XTBN.Y.n30 XThC.XTBN.Y.t56 212.081
R17756 XThC.XTBN.Y.n28 XThC.XTBN.Y.t48 212.081
R17757 XThC.XTBN.Y.n10 XThC.XTBN.Y.t50 212.081
R17758 XThC.XTBN.Y.n1 XThC.XTBN.Y.t18 212.081
R17759 XThC.XTBN.Y.n5 XThC.XTBN.Y.t120 212.081
R17760 XThC.XTBN.Y.n3 XThC.XTBN.Y.t114 212.081
R17761 XThC.XTBN.Y.n74 XThC.XTBN.Y.t101 212.081
R17762 XThC.XTBN.Y.n65 XThC.XTBN.Y.t63 212.081
R17763 XThC.XTBN.Y.n69 XThC.XTBN.Y.t52 212.081
R17764 XThC.XTBN.Y.n67 XThC.XTBN.Y.t44 212.081
R17765 XThC.XTBN.Y.n48 XThC.XTBN.Y.t39 212.081
R17766 XThC.XTBN.Y.n39 XThC.XTBN.Y.t122 212.081
R17767 XThC.XTBN.Y.n43 XThC.XTBN.Y.t109 212.081
R17768 XThC.XTBN.Y.n41 XThC.XTBN.Y.t102 212.081
R17769 XThC.XTBN.Y.n22 XThC.XTBN.Y.t79 212.081
R17770 XThC.XTBN.Y.n13 XThC.XTBN.Y.t36 212.081
R17771 XThC.XTBN.Y.n17 XThC.XTBN.Y.t26 212.081
R17772 XThC.XTBN.Y.n15 XThC.XTBN.Y.t21 212.081
R17773 XThC.XTBN.Y.n99 XThC.XTBN.Y.t54 212.081
R17774 XThC.XTBN.Y.n98 XThC.XTBN.Y.t46 212.081
R17775 XThC.XTBN.Y.n93 XThC.XTBN.Y.t12 212.081
R17776 XThC.XTBN.Y.n92 XThC.XTBN.Y.t6 212.081
R17777 XThC.XTBN.Y.n122 XThC.XTBN.Y.t34 212.081
R17778 XThC.XTBN.Y.n121 XThC.XTBN.Y.t30 212.081
R17779 XThC.XTBN.Y.n116 XThC.XTBN.Y.t103 212.081
R17780 XThC.XTBN.Y.n115 XThC.XTBN.Y.t98 212.081
R17781 XThC.XTBN.Y.n146 XThC.XTBN.Y.t91 212.081
R17782 XThC.XTBN.Y.n145 XThC.XTBN.Y.t88 212.081
R17783 XThC.XTBN.Y.n140 XThC.XTBN.Y.t40 212.081
R17784 XThC.XTBN.Y.n139 XThC.XTBN.Y.t37 212.081
R17785 XThC.XTBN.Y.n170 XThC.XTBN.Y.t28 212.081
R17786 XThC.XTBN.Y.n169 XThC.XTBN.Y.t23 212.081
R17787 XThC.XTBN.Y.n164 XThC.XTBN.Y.t97 212.081
R17788 XThC.XTBN.Y.n163 XThC.XTBN.Y.t95 212.081
R17789 XThC.XTBN.Y.n110 XThC.XTBN.Y.t42 212.081
R17790 XThC.XTBN.Y.n109 XThC.XTBN.Y.t38 212.081
R17791 XThC.XTBN.Y.n104 XThC.XTBN.Y.t119 212.081
R17792 XThC.XTBN.Y.n103 XThC.XTBN.Y.t113 212.081
R17793 XThC.XTBN.Y.n134 XThC.XTBN.Y.t99 212.081
R17794 XThC.XTBN.Y.n133 XThC.XTBN.Y.t96 212.081
R17795 XThC.XTBN.Y.n128 XThC.XTBN.Y.t58 212.081
R17796 XThC.XTBN.Y.n127 XThC.XTBN.Y.t51 212.081
R17797 XThC.XTBN.Y.n158 XThC.XTBN.Y.t13 212.081
R17798 XThC.XTBN.Y.n157 XThC.XTBN.Y.t7 212.081
R17799 XThC.XTBN.Y.n152 XThC.XTBN.Y.t86 212.081
R17800 XThC.XTBN.Y.n151 XThC.XTBN.Y.t81 212.081
R17801 XThC.XTBN.Y.n189 XThC.XTBN.Y.n188 208.965
R17802 XThC.XTBN.Y.n176 XThC.XTBN.Y.n0 188.516
R17803 XThC.XTBN.Y.n88 XThC.XTBN.Y.n87 180.482
R17804 XThC.XTBN.Y.n62 XThC.XTBN.Y.n61 180.482
R17805 XThC.XTBN.Y.n36 XThC.XTBN.Y.n35 180.482
R17806 XThC.XTBN.Y.n11 XThC.XTBN.Y.n10 180.482
R17807 XThC.XTBN.Y.n75 XThC.XTBN.Y.n74 180.482
R17808 XThC.XTBN.Y.n49 XThC.XTBN.Y.n48 180.482
R17809 XThC.XTBN.Y.n23 XThC.XTBN.Y.n22 180.482
R17810 XThC.XTBN.Y.n95 XThC.XTBN.Y.n94 173.761
R17811 XThC.XTBN.Y.n118 XThC.XTBN.Y.n117 173.761
R17812 XThC.XTBN.Y.n142 XThC.XTBN.Y.n141 173.761
R17813 XThC.XTBN.Y.n166 XThC.XTBN.Y.n165 173.761
R17814 XThC.XTBN.Y.n106 XThC.XTBN.Y.n105 173.761
R17815 XThC.XTBN.Y.n130 XThC.XTBN.Y.n129 173.761
R17816 XThC.XTBN.Y.n154 XThC.XTBN.Y.n153 173.761
R17817 XThC.XTBN.Y.n81 XThC.XTBN.Y.n79 152
R17818 XThC.XTBN.Y.n84 XThC.XTBN.Y.n83 152
R17819 XThC.XTBN.Y.n86 XThC.XTBN.Y.n85 152
R17820 XThC.XTBN.Y.n55 XThC.XTBN.Y.n53 152
R17821 XThC.XTBN.Y.n58 XThC.XTBN.Y.n57 152
R17822 XThC.XTBN.Y.n60 XThC.XTBN.Y.n59 152
R17823 XThC.XTBN.Y.n29 XThC.XTBN.Y.n27 152
R17824 XThC.XTBN.Y.n32 XThC.XTBN.Y.n31 152
R17825 XThC.XTBN.Y.n34 XThC.XTBN.Y.n33 152
R17826 XThC.XTBN.Y.n4 XThC.XTBN.Y.n2 152
R17827 XThC.XTBN.Y.n7 XThC.XTBN.Y.n6 152
R17828 XThC.XTBN.Y.n9 XThC.XTBN.Y.n8 152
R17829 XThC.XTBN.Y.n68 XThC.XTBN.Y.n66 152
R17830 XThC.XTBN.Y.n71 XThC.XTBN.Y.n70 152
R17831 XThC.XTBN.Y.n73 XThC.XTBN.Y.n72 152
R17832 XThC.XTBN.Y.n42 XThC.XTBN.Y.n40 152
R17833 XThC.XTBN.Y.n45 XThC.XTBN.Y.n44 152
R17834 XThC.XTBN.Y.n47 XThC.XTBN.Y.n46 152
R17835 XThC.XTBN.Y.n16 XThC.XTBN.Y.n14 152
R17836 XThC.XTBN.Y.n19 XThC.XTBN.Y.n18 152
R17837 XThC.XTBN.Y.n21 XThC.XTBN.Y.n20 152
R17838 XThC.XTBN.Y.n95 XThC.XTBN.Y.n91 152
R17839 XThC.XTBN.Y.n97 XThC.XTBN.Y.n96 152
R17840 XThC.XTBN.Y.n101 XThC.XTBN.Y.n100 152
R17841 XThC.XTBN.Y.n118 XThC.XTBN.Y.n114 152
R17842 XThC.XTBN.Y.n120 XThC.XTBN.Y.n119 152
R17843 XThC.XTBN.Y.n124 XThC.XTBN.Y.n123 152
R17844 XThC.XTBN.Y.n142 XThC.XTBN.Y.n138 152
R17845 XThC.XTBN.Y.n144 XThC.XTBN.Y.n143 152
R17846 XThC.XTBN.Y.n148 XThC.XTBN.Y.n147 152
R17847 XThC.XTBN.Y.n166 XThC.XTBN.Y.n162 152
R17848 XThC.XTBN.Y.n168 XThC.XTBN.Y.n167 152
R17849 XThC.XTBN.Y.n172 XThC.XTBN.Y.n171 152
R17850 XThC.XTBN.Y.n106 XThC.XTBN.Y.n102 152
R17851 XThC.XTBN.Y.n108 XThC.XTBN.Y.n107 152
R17852 XThC.XTBN.Y.n112 XThC.XTBN.Y.n111 152
R17853 XThC.XTBN.Y.n130 XThC.XTBN.Y.n126 152
R17854 XThC.XTBN.Y.n132 XThC.XTBN.Y.n131 152
R17855 XThC.XTBN.Y.n136 XThC.XTBN.Y.n135 152
R17856 XThC.XTBN.Y.n154 XThC.XTBN.Y.n150 152
R17857 XThC.XTBN.Y.n156 XThC.XTBN.Y.n155 152
R17858 XThC.XTBN.Y.n160 XThC.XTBN.Y.n159 152
R17859 XThC.XTBN.Y.n178 XThC.XTBN.Y.n177 152
R17860 XThC.XTBN.Y.n180 XThC.XTBN.Y.n179 152
R17861 XThC.XTBN.Y.n184 XThC.XTBN.Y.n183 152
R17862 XThC.XTBN.Y.n182 XThC.XTBN.Y.t14 139.78
R17863 XThC.XTBN.Y.n181 XThC.XTBN.Y.t105 139.78
R17864 XThC.XTBN.Y.n175 XThC.XTBN.Y.t69 139.78
R17865 XThC.XTBN.Y.n176 XThC.XTBN.Y.t61 139.78
R17866 XThC.XTBN.Y.n87 XThC.XTBN.Y.t123 139.78
R17867 XThC.XTBN.Y.n78 XThC.XTBN.Y.t85 139.78
R17868 XThC.XTBN.Y.n82 XThC.XTBN.Y.t74 139.78
R17869 XThC.XTBN.Y.n80 XThC.XTBN.Y.t65 139.78
R17870 XThC.XTBN.Y.n61 XThC.XTBN.Y.t31 139.78
R17871 XThC.XTBN.Y.n52 XThC.XTBN.Y.t104 139.78
R17872 XThC.XTBN.Y.n56 XThC.XTBN.Y.t94 139.78
R17873 XThC.XTBN.Y.n54 XThC.XTBN.Y.t92 139.78
R17874 XThC.XTBN.Y.n35 XThC.XTBN.Y.t89 139.78
R17875 XThC.XTBN.Y.n26 XThC.XTBN.Y.t41 139.78
R17876 XThC.XTBN.Y.n30 XThC.XTBN.Y.t35 139.78
R17877 XThC.XTBN.Y.n28 XThC.XTBN.Y.t32 139.78
R17878 XThC.XTBN.Y.n10 XThC.XTBN.Y.t118 139.78
R17879 XThC.XTBN.Y.n1 XThC.XTBN.Y.t83 139.78
R17880 XThC.XTBN.Y.n5 XThC.XTBN.Y.t71 139.78
R17881 XThC.XTBN.Y.n3 XThC.XTBN.Y.t62 139.78
R17882 XThC.XTBN.Y.n74 XThC.XTBN.Y.t107 139.78
R17883 XThC.XTBN.Y.n65 XThC.XTBN.Y.t72 139.78
R17884 XThC.XTBN.Y.n69 XThC.XTBN.Y.t57 139.78
R17885 XThC.XTBN.Y.n67 XThC.XTBN.Y.t49 139.78
R17886 XThC.XTBN.Y.n48 XThC.XTBN.Y.t43 139.78
R17887 XThC.XTBN.Y.n39 XThC.XTBN.Y.t10 139.78
R17888 XThC.XTBN.Y.n43 XThC.XTBN.Y.t112 139.78
R17889 XThC.XTBN.Y.n41 XThC.XTBN.Y.t108 139.78
R17890 XThC.XTBN.Y.n22 XThC.XTBN.Y.t121 139.78
R17891 XThC.XTBN.Y.n13 XThC.XTBN.Y.t84 139.78
R17892 XThC.XTBN.Y.n17 XThC.XTBN.Y.t73 139.78
R17893 XThC.XTBN.Y.n15 XThC.XTBN.Y.t64 139.78
R17894 XThC.XTBN.Y.n99 XThC.XTBN.Y.t76 139.78
R17895 XThC.XTBN.Y.n98 XThC.XTBN.Y.t67 139.78
R17896 XThC.XTBN.Y.n93 XThC.XTBN.Y.t29 139.78
R17897 XThC.XTBN.Y.n92 XThC.XTBN.Y.t24 139.78
R17898 XThC.XTBN.Y.n122 XThC.XTBN.Y.t15 139.78
R17899 XThC.XTBN.Y.n121 XThC.XTBN.Y.t8 139.78
R17900 XThC.XTBN.Y.n116 XThC.XTBN.Y.t87 139.78
R17901 XThC.XTBN.Y.n115 XThC.XTBN.Y.t82 139.78
R17902 XThC.XTBN.Y.n146 XThC.XTBN.Y.t66 139.78
R17903 XThC.XTBN.Y.n145 XThC.XTBN.Y.t60 139.78
R17904 XThC.XTBN.Y.n140 XThC.XTBN.Y.t22 139.78
R17905 XThC.XTBN.Y.n139 XThC.XTBN.Y.t20 139.78
R17906 XThC.XTBN.Y.n170 XThC.XTBN.Y.t4 139.78
R17907 XThC.XTBN.Y.n169 XThC.XTBN.Y.t117 139.78
R17908 XThC.XTBN.Y.n164 XThC.XTBN.Y.t80 139.78
R17909 XThC.XTBN.Y.n163 XThC.XTBN.Y.t78 139.78
R17910 XThC.XTBN.Y.n110 XThC.XTBN.Y.t59 139.78
R17911 XThC.XTBN.Y.n109 XThC.XTBN.Y.t55 139.78
R17912 XThC.XTBN.Y.n104 XThC.XTBN.Y.t19 139.78
R17913 XThC.XTBN.Y.n103 XThC.XTBN.Y.t16 139.78
R17914 XThC.XTBN.Y.n134 XThC.XTBN.Y.t115 139.78
R17915 XThC.XTBN.Y.n133 XThC.XTBN.Y.t110 139.78
R17916 XThC.XTBN.Y.n128 XThC.XTBN.Y.t77 139.78
R17917 XThC.XTBN.Y.n127 XThC.XTBN.Y.t68 139.78
R17918 XThC.XTBN.Y.n158 XThC.XTBN.Y.t53 139.78
R17919 XThC.XTBN.Y.n157 XThC.XTBN.Y.t45 139.78
R17920 XThC.XTBN.Y.n152 XThC.XTBN.Y.t11 139.78
R17921 XThC.XTBN.Y.n151 XThC.XTBN.Y.t5 139.78
R17922 XThC.XTBN.Y XThC.XTBN.Y.n192 96.8352
R17923 XThC.XTBN.Y.n187 XThC.XTBN.Y.n0 64.6909
R17924 XThC.XTBN.Y.n97 XThC.XTBN.Y.n91 49.6611
R17925 XThC.XTBN.Y.n120 XThC.XTBN.Y.n114 49.6611
R17926 XThC.XTBN.Y.n144 XThC.XTBN.Y.n138 49.6611
R17927 XThC.XTBN.Y.n168 XThC.XTBN.Y.n162 49.6611
R17928 XThC.XTBN.Y.n108 XThC.XTBN.Y.n102 49.6611
R17929 XThC.XTBN.Y.n132 XThC.XTBN.Y.n126 49.6611
R17930 XThC.XTBN.Y.n156 XThC.XTBN.Y.n150 49.6611
R17931 XThC.XTBN.Y.n100 XThC.XTBN.Y.n98 44.549
R17932 XThC.XTBN.Y.n123 XThC.XTBN.Y.n121 44.549
R17933 XThC.XTBN.Y.n147 XThC.XTBN.Y.n145 44.549
R17934 XThC.XTBN.Y.n171 XThC.XTBN.Y.n169 44.549
R17935 XThC.XTBN.Y.n111 XThC.XTBN.Y.n109 44.549
R17936 XThC.XTBN.Y.n135 XThC.XTBN.Y.n133 44.549
R17937 XThC.XTBN.Y.n159 XThC.XTBN.Y.n157 44.549
R17938 XThC.XTBN.Y.n94 XThC.XTBN.Y.n93 43.0884
R17939 XThC.XTBN.Y.n117 XThC.XTBN.Y.n116 43.0884
R17940 XThC.XTBN.Y.n141 XThC.XTBN.Y.n140 43.0884
R17941 XThC.XTBN.Y.n165 XThC.XTBN.Y.n164 43.0884
R17942 XThC.XTBN.Y.n105 XThC.XTBN.Y.n104 43.0884
R17943 XThC.XTBN.Y.n129 XThC.XTBN.Y.n128 43.0884
R17944 XThC.XTBN.Y.n153 XThC.XTBN.Y.n152 43.0884
R17945 XThC.XTBN.Y.n177 XThC.XTBN.Y.n176 30.6732
R17946 XThC.XTBN.Y.n177 XThC.XTBN.Y.n175 30.6732
R17947 XThC.XTBN.Y.n180 XThC.XTBN.Y.n175 30.6732
R17948 XThC.XTBN.Y.n181 XThC.XTBN.Y.n180 30.6732
R17949 XThC.XTBN.Y.n183 XThC.XTBN.Y.n181 30.6732
R17950 XThC.XTBN.Y.n183 XThC.XTBN.Y.n182 30.6732
R17951 XThC.XTBN.Y.n81 XThC.XTBN.Y.n80 30.6732
R17952 XThC.XTBN.Y.n82 XThC.XTBN.Y.n81 30.6732
R17953 XThC.XTBN.Y.n83 XThC.XTBN.Y.n82 30.6732
R17954 XThC.XTBN.Y.n83 XThC.XTBN.Y.n78 30.6732
R17955 XThC.XTBN.Y.n86 XThC.XTBN.Y.n78 30.6732
R17956 XThC.XTBN.Y.n87 XThC.XTBN.Y.n86 30.6732
R17957 XThC.XTBN.Y.n55 XThC.XTBN.Y.n54 30.6732
R17958 XThC.XTBN.Y.n56 XThC.XTBN.Y.n55 30.6732
R17959 XThC.XTBN.Y.n57 XThC.XTBN.Y.n56 30.6732
R17960 XThC.XTBN.Y.n57 XThC.XTBN.Y.n52 30.6732
R17961 XThC.XTBN.Y.n60 XThC.XTBN.Y.n52 30.6732
R17962 XThC.XTBN.Y.n61 XThC.XTBN.Y.n60 30.6732
R17963 XThC.XTBN.Y.n29 XThC.XTBN.Y.n28 30.6732
R17964 XThC.XTBN.Y.n30 XThC.XTBN.Y.n29 30.6732
R17965 XThC.XTBN.Y.n31 XThC.XTBN.Y.n30 30.6732
R17966 XThC.XTBN.Y.n31 XThC.XTBN.Y.n26 30.6732
R17967 XThC.XTBN.Y.n34 XThC.XTBN.Y.n26 30.6732
R17968 XThC.XTBN.Y.n35 XThC.XTBN.Y.n34 30.6732
R17969 XThC.XTBN.Y.n4 XThC.XTBN.Y.n3 30.6732
R17970 XThC.XTBN.Y.n5 XThC.XTBN.Y.n4 30.6732
R17971 XThC.XTBN.Y.n6 XThC.XTBN.Y.n5 30.6732
R17972 XThC.XTBN.Y.n6 XThC.XTBN.Y.n1 30.6732
R17973 XThC.XTBN.Y.n9 XThC.XTBN.Y.n1 30.6732
R17974 XThC.XTBN.Y.n10 XThC.XTBN.Y.n9 30.6732
R17975 XThC.XTBN.Y.n68 XThC.XTBN.Y.n67 30.6732
R17976 XThC.XTBN.Y.n69 XThC.XTBN.Y.n68 30.6732
R17977 XThC.XTBN.Y.n70 XThC.XTBN.Y.n69 30.6732
R17978 XThC.XTBN.Y.n70 XThC.XTBN.Y.n65 30.6732
R17979 XThC.XTBN.Y.n73 XThC.XTBN.Y.n65 30.6732
R17980 XThC.XTBN.Y.n74 XThC.XTBN.Y.n73 30.6732
R17981 XThC.XTBN.Y.n42 XThC.XTBN.Y.n41 30.6732
R17982 XThC.XTBN.Y.n43 XThC.XTBN.Y.n42 30.6732
R17983 XThC.XTBN.Y.n44 XThC.XTBN.Y.n43 30.6732
R17984 XThC.XTBN.Y.n44 XThC.XTBN.Y.n39 30.6732
R17985 XThC.XTBN.Y.n47 XThC.XTBN.Y.n39 30.6732
R17986 XThC.XTBN.Y.n48 XThC.XTBN.Y.n47 30.6732
R17987 XThC.XTBN.Y.n16 XThC.XTBN.Y.n15 30.6732
R17988 XThC.XTBN.Y.n17 XThC.XTBN.Y.n16 30.6732
R17989 XThC.XTBN.Y.n18 XThC.XTBN.Y.n17 30.6732
R17990 XThC.XTBN.Y.n18 XThC.XTBN.Y.n13 30.6732
R17991 XThC.XTBN.Y.n21 XThC.XTBN.Y.n13 30.6732
R17992 XThC.XTBN.Y.n22 XThC.XTBN.Y.n21 30.6732
R17993 XThC.XTBN.Y.n188 XThC.XTBN.Y.t2 26.5955
R17994 XThC.XTBN.Y.n188 XThC.XTBN.Y.t3 26.5955
R17995 XThC.XTBN.Y.n192 XThC.XTBN.Y.t1 24.9236
R17996 XThC.XTBN.Y.n192 XThC.XTBN.Y.t0 24.9236
R17997 XThC.XTBN.Y.n96 XThC.XTBN.Y.n95 21.7605
R17998 XThC.XTBN.Y.n119 XThC.XTBN.Y.n118 21.7605
R17999 XThC.XTBN.Y.n143 XThC.XTBN.Y.n142 21.7605
R18000 XThC.XTBN.Y.n167 XThC.XTBN.Y.n166 21.7605
R18001 XThC.XTBN.Y.n107 XThC.XTBN.Y.n106 21.7605
R18002 XThC.XTBN.Y.n131 XThC.XTBN.Y.n130 21.7605
R18003 XThC.XTBN.Y.n155 XThC.XTBN.Y.n154 21.7605
R18004 XThC.XTBN.Y.n84 XThC.XTBN.Y.n79 21.5045
R18005 XThC.XTBN.Y.n58 XThC.XTBN.Y.n53 21.5045
R18006 XThC.XTBN.Y.n32 XThC.XTBN.Y.n27 21.5045
R18007 XThC.XTBN.Y.n7 XThC.XTBN.Y.n2 21.5045
R18008 XThC.XTBN.Y.n71 XThC.XTBN.Y.n66 21.5045
R18009 XThC.XTBN.Y.n45 XThC.XTBN.Y.n40 21.5045
R18010 XThC.XTBN.Y.n19 XThC.XTBN.Y.n14 21.5045
R18011 XThC.XTBN.Y.n178 XThC.XTBN.Y 21.2485
R18012 XThC.XTBN.Y.n85 XThC.XTBN.Y 19.9685
R18013 XThC.XTBN.Y.n59 XThC.XTBN.Y 19.9685
R18014 XThC.XTBN.Y.n33 XThC.XTBN.Y 19.9685
R18015 XThC.XTBN.Y.n8 XThC.XTBN.Y 19.9685
R18016 XThC.XTBN.Y.n72 XThC.XTBN.Y 19.9685
R18017 XThC.XTBN.Y.n46 XThC.XTBN.Y 19.9685
R18018 XThC.XTBN.Y.n20 XThC.XTBN.Y 19.9685
R18019 XThC.XTBN.Y.n179 XThC.XTBN.Y 19.2005
R18020 XThC.XTBN.Y.n94 XThC.XTBN.Y.n92 18.2581
R18021 XThC.XTBN.Y.n117 XThC.XTBN.Y.n115 18.2581
R18022 XThC.XTBN.Y.n141 XThC.XTBN.Y.n139 18.2581
R18023 XThC.XTBN.Y.n165 XThC.XTBN.Y.n163 18.2581
R18024 XThC.XTBN.Y.n105 XThC.XTBN.Y.n103 18.2581
R18025 XThC.XTBN.Y.n129 XThC.XTBN.Y.n127 18.2581
R18026 XThC.XTBN.Y.n153 XThC.XTBN.Y.n151 18.2581
R18027 XThC.XTBN.Y.n113 XThC.XTBN.Y.n101 17.1655
R18028 XThC.XTBN.Y.n88 XThC.XTBN.Y 17.1525
R18029 XThC.XTBN.Y.n62 XThC.XTBN.Y 17.1525
R18030 XThC.XTBN.Y.n36 XThC.XTBN.Y 17.1525
R18031 XThC.XTBN.Y.n11 XThC.XTBN.Y 17.1525
R18032 XThC.XTBN.Y.n75 XThC.XTBN.Y 17.1525
R18033 XThC.XTBN.Y.n49 XThC.XTBN.Y 17.1525
R18034 XThC.XTBN.Y.n23 XThC.XTBN.Y 17.1525
R18035 XThC.XTBN.Y.n100 XThC.XTBN.Y.n99 16.7975
R18036 XThC.XTBN.Y.n123 XThC.XTBN.Y.n122 16.7975
R18037 XThC.XTBN.Y.n147 XThC.XTBN.Y.n146 16.7975
R18038 XThC.XTBN.Y.n171 XThC.XTBN.Y.n170 16.7975
R18039 XThC.XTBN.Y.n111 XThC.XTBN.Y.n110 16.7975
R18040 XThC.XTBN.Y.n135 XThC.XTBN.Y.n134 16.7975
R18041 XThC.XTBN.Y.n159 XThC.XTBN.Y.n158 16.7975
R18042 XThC.XTBN.Y.n125 XThC.XTBN.Y.n124 16.0405
R18043 XThC.XTBN.Y.n149 XThC.XTBN.Y.n148 16.0405
R18044 XThC.XTBN.Y.n173 XThC.XTBN.Y.n172 16.0405
R18045 XThC.XTBN.Y.n113 XThC.XTBN.Y.n112 16.0405
R18046 XThC.XTBN.Y.n137 XThC.XTBN.Y.n136 16.0405
R18047 XThC.XTBN.Y.n161 XThC.XTBN.Y.n160 16.0405
R18048 XThC.XTBN.Y.n25 XThC.XTBN.Y.n12 15.262
R18049 XThC.XTBN.Y.n101 XThC.XTBN.Y 15.0405
R18050 XThC.XTBN.Y.n124 XThC.XTBN.Y 15.0405
R18051 XThC.XTBN.Y.n148 XThC.XTBN.Y 15.0405
R18052 XThC.XTBN.Y.n172 XThC.XTBN.Y 15.0405
R18053 XThC.XTBN.Y.n112 XThC.XTBN.Y 15.0405
R18054 XThC.XTBN.Y.n136 XThC.XTBN.Y 15.0405
R18055 XThC.XTBN.Y.n160 XThC.XTBN.Y 15.0405
R18056 XThC.XTBN.Y.n90 XThC.XTBN.Y.n89 13.8005
R18057 XThC.XTBN.Y.n64 XThC.XTBN.Y.n63 13.8005
R18058 XThC.XTBN.Y.n38 XThC.XTBN.Y.n37 13.8005
R18059 XThC.XTBN.Y.n77 XThC.XTBN.Y.n76 13.8005
R18060 XThC.XTBN.Y.n51 XThC.XTBN.Y.n50 13.8005
R18061 XThC.XTBN.Y.n25 XThC.XTBN.Y.n24 13.8005
R18062 XThC.XTBN.Y.n190 XThC.XTBN.Y 12.5445
R18063 XThC.XTBN.Y.n191 XThC.XTBN.Y 11.2645
R18064 XThC.XTBN.Y.n185 XThC.XTBN.Y.n184 9.2165
R18065 XThC.XTBN.Y.n185 XThC.XTBN.Y 7.9365
R18066 XThC.XTBN.Y.n96 XThC.XTBN.Y 6.7205
R18067 XThC.XTBN.Y.n119 XThC.XTBN.Y 6.7205
R18068 XThC.XTBN.Y.n143 XThC.XTBN.Y 6.7205
R18069 XThC.XTBN.Y.n167 XThC.XTBN.Y 6.7205
R18070 XThC.XTBN.Y.n107 XThC.XTBN.Y 6.7205
R18071 XThC.XTBN.Y.n131 XThC.XTBN.Y 6.7205
R18072 XThC.XTBN.Y.n155 XThC.XTBN.Y 6.7205
R18073 XThC.XTBN.Y.n93 XThC.XTBN.Y.n91 6.57323
R18074 XThC.XTBN.Y.n116 XThC.XTBN.Y.n114 6.57323
R18075 XThC.XTBN.Y.n140 XThC.XTBN.Y.n138 6.57323
R18076 XThC.XTBN.Y.n164 XThC.XTBN.Y.n162 6.57323
R18077 XThC.XTBN.Y.n104 XThC.XTBN.Y.n102 6.57323
R18078 XThC.XTBN.Y.n128 XThC.XTBN.Y.n126 6.57323
R18079 XThC.XTBN.Y.n152 XThC.XTBN.Y.n150 6.57323
R18080 XThC.XTBN.Y.n184 XThC.XTBN.Y 6.4005
R18081 XThC.XTBN.Y.n191 XThC.XTBN.Y 6.1445
R18082 XThC.XTBN.Y.n187 XThC.XTBN.Y.n186 5.74665
R18083 XThC.XTBN.Y.n186 XThC.XTBN.Y.n174 5.68319
R18084 XThC.XTBN.Y.n98 XThC.XTBN.Y.n97 5.11262
R18085 XThC.XTBN.Y.n121 XThC.XTBN.Y.n120 5.11262
R18086 XThC.XTBN.Y.n145 XThC.XTBN.Y.n144 5.11262
R18087 XThC.XTBN.Y.n169 XThC.XTBN.Y.n168 5.11262
R18088 XThC.XTBN.Y.n109 XThC.XTBN.Y.n108 5.11262
R18089 XThC.XTBN.Y.n133 XThC.XTBN.Y.n132 5.11262
R18090 XThC.XTBN.Y.n157 XThC.XTBN.Y.n156 5.11262
R18091 XThC.XTBN.Y.n190 XThC.XTBN.Y.n187 5.06717
R18092 XThC.XTBN.Y XThC.XTBN.Y.n190 4.8645
R18093 XThC.XTBN.Y XThC.XTBN.Y.n191 4.65505
R18094 XThC.XTBN.Y.n186 XThC.XTBN.Y.n185 4.6505
R18095 XThC.XTBN.Y.n89 XThC.XTBN.Y 4.6085
R18096 XThC.XTBN.Y.n63 XThC.XTBN.Y 4.6085
R18097 XThC.XTBN.Y.n37 XThC.XTBN.Y 4.6085
R18098 XThC.XTBN.Y.n12 XThC.XTBN.Y 4.6085
R18099 XThC.XTBN.Y.n76 XThC.XTBN.Y 4.6085
R18100 XThC.XTBN.Y.n50 XThC.XTBN.Y 4.6085
R18101 XThC.XTBN.Y.n24 XThC.XTBN.Y 4.6085
R18102 XThC.XTBN.Y.n179 XThC.XTBN.Y 4.3525
R18103 XThC.XTBN.Y.n85 XThC.XTBN.Y 3.5845
R18104 XThC.XTBN.Y.n59 XThC.XTBN.Y 3.5845
R18105 XThC.XTBN.Y.n33 XThC.XTBN.Y 3.5845
R18106 XThC.XTBN.Y.n8 XThC.XTBN.Y 3.5845
R18107 XThC.XTBN.Y.n72 XThC.XTBN.Y 3.5845
R18108 XThC.XTBN.Y.n46 XThC.XTBN.Y 3.5845
R18109 XThC.XTBN.Y.n20 XThC.XTBN.Y 3.5845
R18110 XThC.XTBN.Y XThC.XTBN.Y.n0 2.3045
R18111 XThC.XTBN.Y XThC.XTBN.Y.n178 2.3045
R18112 XThC.XTBN.Y XThC.XTBN.Y.n189 2.0485
R18113 XThC.XTBN.Y.n89 XThC.XTBN.Y.n88 1.7925
R18114 XThC.XTBN.Y.n63 XThC.XTBN.Y.n62 1.7925
R18115 XThC.XTBN.Y.n37 XThC.XTBN.Y.n36 1.7925
R18116 XThC.XTBN.Y.n12 XThC.XTBN.Y.n11 1.7925
R18117 XThC.XTBN.Y.n76 XThC.XTBN.Y.n75 1.7925
R18118 XThC.XTBN.Y.n50 XThC.XTBN.Y.n49 1.7925
R18119 XThC.XTBN.Y.n24 XThC.XTBN.Y.n23 1.7925
R18120 XThC.XTBN.Y.n174 XThC.XTBN.Y.n173 1.59665
R18121 XThC.XTBN.Y.n189 XThC.XTBN.Y 1.55202
R18122 XThC.XTBN.Y XThC.XTBN.Y.n84 1.5365
R18123 XThC.XTBN.Y XThC.XTBN.Y.n58 1.5365
R18124 XThC.XTBN.Y XThC.XTBN.Y.n32 1.5365
R18125 XThC.XTBN.Y XThC.XTBN.Y.n7 1.5365
R18126 XThC.XTBN.Y XThC.XTBN.Y.n71 1.5365
R18127 XThC.XTBN.Y XThC.XTBN.Y.n45 1.5365
R18128 XThC.XTBN.Y XThC.XTBN.Y.n19 1.5365
R18129 XThC.XTBN.Y.n149 XThC.XTBN.Y.n137 1.49088
R18130 XThC.XTBN.Y.n125 XThC.XTBN.Y.n113 1.49088
R18131 XThC.XTBN.Y.n173 XThC.XTBN.Y.n161 1.48608
R18132 XThC.XTBN.Y.n51 XThC.XTBN.Y.n38 1.46204
R18133 XThC.XTBN.Y.n77 XThC.XTBN.Y.n64 1.46204
R18134 XThC.XTBN.Y.n38 XThC.XTBN.Y.n25 1.15435
R18135 XThC.XTBN.Y.n64 XThC.XTBN.Y.n51 1.15435
R18136 XThC.XTBN.Y.n90 XThC.XTBN.Y.n77 1.15435
R18137 XThC.XTBN.Y.n174 XThC.XTBN.Y.n90 1.14473
R18138 XThC.XTBN.Y.n161 XThC.XTBN.Y.n149 1.13031
R18139 XThC.XTBN.Y.n137 XThC.XTBN.Y.n125 1.1255
R18140 XThC.XTBN.Y.n79 XThC.XTBN.Y 0.5125
R18141 XThC.XTBN.Y.n53 XThC.XTBN.Y 0.5125
R18142 XThC.XTBN.Y.n27 XThC.XTBN.Y 0.5125
R18143 XThC.XTBN.Y.n2 XThC.XTBN.Y 0.5125
R18144 XThC.XTBN.Y.n66 XThC.XTBN.Y 0.5125
R18145 XThC.XTBN.Y.n40 XThC.XTBN.Y 0.5125
R18146 XThC.XTBN.Y.n14 XThC.XTBN.Y 0.5125
R18147 XThC.Tn[6].n2 XThC.Tn[6].n1 332.332
R18148 XThC.Tn[6].n2 XThC.Tn[6].n0 296.493
R18149 XThC.Tn[6].n12 XThC.Tn[6].n10 161.406
R18150 XThC.Tn[6].n15 XThC.Tn[6].n13 161.406
R18151 XThC.Tn[6].n18 XThC.Tn[6].n16 161.406
R18152 XThC.Tn[6].n21 XThC.Tn[6].n19 161.406
R18153 XThC.Tn[6].n24 XThC.Tn[6].n22 161.406
R18154 XThC.Tn[6].n27 XThC.Tn[6].n25 161.406
R18155 XThC.Tn[6].n30 XThC.Tn[6].n28 161.406
R18156 XThC.Tn[6].n33 XThC.Tn[6].n31 161.406
R18157 XThC.Tn[6].n36 XThC.Tn[6].n34 161.406
R18158 XThC.Tn[6].n39 XThC.Tn[6].n37 161.406
R18159 XThC.Tn[6].n42 XThC.Tn[6].n40 161.406
R18160 XThC.Tn[6].n45 XThC.Tn[6].n43 161.406
R18161 XThC.Tn[6].n48 XThC.Tn[6].n46 161.406
R18162 XThC.Tn[6].n51 XThC.Tn[6].n49 161.406
R18163 XThC.Tn[6].n54 XThC.Tn[6].n52 161.406
R18164 XThC.Tn[6].n57 XThC.Tn[6].n55 161.406
R18165 XThC.Tn[6].n10 XThC.Tn[6].t26 161.202
R18166 XThC.Tn[6].n13 XThC.Tn[6].t13 161.202
R18167 XThC.Tn[6].n16 XThC.Tn[6].t17 161.202
R18168 XThC.Tn[6].n19 XThC.Tn[6].t18 161.202
R18169 XThC.Tn[6].n22 XThC.Tn[6].t37 161.202
R18170 XThC.Tn[6].n25 XThC.Tn[6].t38 161.202
R18171 XThC.Tn[6].n28 XThC.Tn[6].t22 161.202
R18172 XThC.Tn[6].n31 XThC.Tn[6].t29 161.202
R18173 XThC.Tn[6].n34 XThC.Tn[6].t31 161.202
R18174 XThC.Tn[6].n37 XThC.Tn[6].t19 161.202
R18175 XThC.Tn[6].n40 XThC.Tn[6].t21 161.202
R18176 XThC.Tn[6].n43 XThC.Tn[6].t32 161.202
R18177 XThC.Tn[6].n46 XThC.Tn[6].t41 161.202
R18178 XThC.Tn[6].n49 XThC.Tn[6].t43 161.202
R18179 XThC.Tn[6].n52 XThC.Tn[6].t24 161.202
R18180 XThC.Tn[6].n55 XThC.Tn[6].t34 161.202
R18181 XThC.Tn[6].n10 XThC.Tn[6].t23 145.137
R18182 XThC.Tn[6].n13 XThC.Tn[6].t40 145.137
R18183 XThC.Tn[6].n16 XThC.Tn[6].t42 145.137
R18184 XThC.Tn[6].n19 XThC.Tn[6].t12 145.137
R18185 XThC.Tn[6].n22 XThC.Tn[6].t33 145.137
R18186 XThC.Tn[6].n25 XThC.Tn[6].t35 145.137
R18187 XThC.Tn[6].n28 XThC.Tn[6].t16 145.137
R18188 XThC.Tn[6].n31 XThC.Tn[6].t25 145.137
R18189 XThC.Tn[6].n34 XThC.Tn[6].t27 145.137
R18190 XThC.Tn[6].n37 XThC.Tn[6].t14 145.137
R18191 XThC.Tn[6].n40 XThC.Tn[6].t15 145.137
R18192 XThC.Tn[6].n43 XThC.Tn[6].t28 145.137
R18193 XThC.Tn[6].n46 XThC.Tn[6].t36 145.137
R18194 XThC.Tn[6].n49 XThC.Tn[6].t39 145.137
R18195 XThC.Tn[6].n52 XThC.Tn[6].t20 145.137
R18196 XThC.Tn[6].n55 XThC.Tn[6].t30 145.137
R18197 XThC.Tn[6].n7 XThC.Tn[6].n6 135.248
R18198 XThC.Tn[6].n9 XThC.Tn[6].n3 98.982
R18199 XThC.Tn[6].n8 XThC.Tn[6].n4 98.982
R18200 XThC.Tn[6].n7 XThC.Tn[6].n5 98.982
R18201 XThC.Tn[6].n9 XThC.Tn[6].n8 36.2672
R18202 XThC.Tn[6].n8 XThC.Tn[6].n7 36.2672
R18203 XThC.Tn[6].n59 XThC.Tn[6].n9 32.6405
R18204 XThC.Tn[6].n1 XThC.Tn[6].t5 26.5955
R18205 XThC.Tn[6].n1 XThC.Tn[6].t4 26.5955
R18206 XThC.Tn[6].n0 XThC.Tn[6].t7 26.5955
R18207 XThC.Tn[6].n0 XThC.Tn[6].t6 26.5955
R18208 XThC.Tn[6].n3 XThC.Tn[6].t8 24.9236
R18209 XThC.Tn[6].n3 XThC.Tn[6].t11 24.9236
R18210 XThC.Tn[6].n4 XThC.Tn[6].t10 24.9236
R18211 XThC.Tn[6].n4 XThC.Tn[6].t9 24.9236
R18212 XThC.Tn[6].n5 XThC.Tn[6].t1 24.9236
R18213 XThC.Tn[6].n5 XThC.Tn[6].t0 24.9236
R18214 XThC.Tn[6].n6 XThC.Tn[6].t3 24.9236
R18215 XThC.Tn[6].n6 XThC.Tn[6].t2 24.9236
R18216 XThC.Tn[6].n60 XThC.Tn[6].n2 18.5605
R18217 XThC.Tn[6].n60 XThC.Tn[6].n59 11.5205
R18218 XThC.Tn[6].n59 XThC.Tn[6].n58 3.18344
R18219 XThC.Tn[6].n58 XThC.Tn[6] 3.09179
R18220 XThC.Tn[6].n15 XThC.Tn[6] 0.931056
R18221 XThC.Tn[6].n18 XThC.Tn[6] 0.931056
R18222 XThC.Tn[6].n21 XThC.Tn[6] 0.931056
R18223 XThC.Tn[6].n24 XThC.Tn[6] 0.931056
R18224 XThC.Tn[6].n27 XThC.Tn[6] 0.931056
R18225 XThC.Tn[6].n30 XThC.Tn[6] 0.931056
R18226 XThC.Tn[6].n33 XThC.Tn[6] 0.931056
R18227 XThC.Tn[6].n36 XThC.Tn[6] 0.931056
R18228 XThC.Tn[6].n39 XThC.Tn[6] 0.931056
R18229 XThC.Tn[6].n42 XThC.Tn[6] 0.931056
R18230 XThC.Tn[6].n45 XThC.Tn[6] 0.931056
R18231 XThC.Tn[6].n48 XThC.Tn[6] 0.931056
R18232 XThC.Tn[6].n51 XThC.Tn[6] 0.931056
R18233 XThC.Tn[6].n54 XThC.Tn[6] 0.931056
R18234 XThC.Tn[6].n57 XThC.Tn[6] 0.931056
R18235 XThC.Tn[6] XThC.Tn[6].n60 0.6405
R18236 XThC.Tn[6] XThC.Tn[6].n12 0.396333
R18237 XThC.Tn[6] XThC.Tn[6].n15 0.396333
R18238 XThC.Tn[6] XThC.Tn[6].n18 0.396333
R18239 XThC.Tn[6] XThC.Tn[6].n21 0.396333
R18240 XThC.Tn[6] XThC.Tn[6].n24 0.396333
R18241 XThC.Tn[6] XThC.Tn[6].n27 0.396333
R18242 XThC.Tn[6] XThC.Tn[6].n30 0.396333
R18243 XThC.Tn[6] XThC.Tn[6].n33 0.396333
R18244 XThC.Tn[6] XThC.Tn[6].n36 0.396333
R18245 XThC.Tn[6] XThC.Tn[6].n39 0.396333
R18246 XThC.Tn[6] XThC.Tn[6].n42 0.396333
R18247 XThC.Tn[6] XThC.Tn[6].n45 0.396333
R18248 XThC.Tn[6] XThC.Tn[6].n48 0.396333
R18249 XThC.Tn[6] XThC.Tn[6].n51 0.396333
R18250 XThC.Tn[6] XThC.Tn[6].n54 0.396333
R18251 XThC.Tn[6] XThC.Tn[6].n57 0.396333
R18252 XThC.Tn[6].n11 XThC.Tn[6] 0.104667
R18253 XThC.Tn[6].n14 XThC.Tn[6] 0.104667
R18254 XThC.Tn[6].n17 XThC.Tn[6] 0.104667
R18255 XThC.Tn[6].n20 XThC.Tn[6] 0.104667
R18256 XThC.Tn[6].n23 XThC.Tn[6] 0.104667
R18257 XThC.Tn[6].n26 XThC.Tn[6] 0.104667
R18258 XThC.Tn[6].n29 XThC.Tn[6] 0.104667
R18259 XThC.Tn[6].n32 XThC.Tn[6] 0.104667
R18260 XThC.Tn[6].n35 XThC.Tn[6] 0.104667
R18261 XThC.Tn[6].n38 XThC.Tn[6] 0.104667
R18262 XThC.Tn[6].n41 XThC.Tn[6] 0.104667
R18263 XThC.Tn[6].n44 XThC.Tn[6] 0.104667
R18264 XThC.Tn[6].n47 XThC.Tn[6] 0.104667
R18265 XThC.Tn[6].n50 XThC.Tn[6] 0.104667
R18266 XThC.Tn[6].n53 XThC.Tn[6] 0.104667
R18267 XThC.Tn[6].n56 XThC.Tn[6] 0.104667
R18268 XThC.Tn[6].n11 XThC.Tn[6] 0.0309878
R18269 XThC.Tn[6].n14 XThC.Tn[6] 0.0309878
R18270 XThC.Tn[6].n17 XThC.Tn[6] 0.0309878
R18271 XThC.Tn[6].n20 XThC.Tn[6] 0.0309878
R18272 XThC.Tn[6].n23 XThC.Tn[6] 0.0309878
R18273 XThC.Tn[6].n26 XThC.Tn[6] 0.0309878
R18274 XThC.Tn[6].n29 XThC.Tn[6] 0.0309878
R18275 XThC.Tn[6].n32 XThC.Tn[6] 0.0309878
R18276 XThC.Tn[6].n35 XThC.Tn[6] 0.0309878
R18277 XThC.Tn[6].n38 XThC.Tn[6] 0.0309878
R18278 XThC.Tn[6].n41 XThC.Tn[6] 0.0309878
R18279 XThC.Tn[6].n44 XThC.Tn[6] 0.0309878
R18280 XThC.Tn[6].n47 XThC.Tn[6] 0.0309878
R18281 XThC.Tn[6].n50 XThC.Tn[6] 0.0309878
R18282 XThC.Tn[6].n53 XThC.Tn[6] 0.0309878
R18283 XThC.Tn[6].n56 XThC.Tn[6] 0.0309878
R18284 XThC.Tn[6].n12 XThC.Tn[6].n11 0.027939
R18285 XThC.Tn[6].n15 XThC.Tn[6].n14 0.027939
R18286 XThC.Tn[6].n18 XThC.Tn[6].n17 0.027939
R18287 XThC.Tn[6].n21 XThC.Tn[6].n20 0.027939
R18288 XThC.Tn[6].n24 XThC.Tn[6].n23 0.027939
R18289 XThC.Tn[6].n27 XThC.Tn[6].n26 0.027939
R18290 XThC.Tn[6].n30 XThC.Tn[6].n29 0.027939
R18291 XThC.Tn[6].n33 XThC.Tn[6].n32 0.027939
R18292 XThC.Tn[6].n36 XThC.Tn[6].n35 0.027939
R18293 XThC.Tn[6].n39 XThC.Tn[6].n38 0.027939
R18294 XThC.Tn[6].n42 XThC.Tn[6].n41 0.027939
R18295 XThC.Tn[6].n45 XThC.Tn[6].n44 0.027939
R18296 XThC.Tn[6].n48 XThC.Tn[6].n47 0.027939
R18297 XThC.Tn[6].n51 XThC.Tn[6].n50 0.027939
R18298 XThC.Tn[6].n54 XThC.Tn[6].n53 0.027939
R18299 XThC.Tn[6].n57 XThC.Tn[6].n56 0.027939
R18300 XThC.Tn[6].n58 XThC.Tn[6] 0.0140108
R18301 XThR.Tn[9].n8 XThR.Tn[9].n7 256.104
R18302 XThR.Tn[9].n5 XThR.Tn[9].n3 243.68
R18303 XThR.Tn[9].n2 XThR.Tn[9].n1 241.847
R18304 XThR.Tn[9].n5 XThR.Tn[9].n4 205.28
R18305 XThR.Tn[9].n8 XThR.Tn[9].n6 202.094
R18306 XThR.Tn[9].n2 XThR.Tn[9].n0 185
R18307 XThR.Tn[9] XThR.Tn[9].n82 161.363
R18308 XThR.Tn[9] XThR.Tn[9].n77 161.363
R18309 XThR.Tn[9] XThR.Tn[9].n72 161.363
R18310 XThR.Tn[9] XThR.Tn[9].n67 161.363
R18311 XThR.Tn[9] XThR.Tn[9].n62 161.363
R18312 XThR.Tn[9] XThR.Tn[9].n57 161.363
R18313 XThR.Tn[9] XThR.Tn[9].n52 161.363
R18314 XThR.Tn[9] XThR.Tn[9].n47 161.363
R18315 XThR.Tn[9] XThR.Tn[9].n42 161.363
R18316 XThR.Tn[9] XThR.Tn[9].n37 161.363
R18317 XThR.Tn[9] XThR.Tn[9].n32 161.363
R18318 XThR.Tn[9] XThR.Tn[9].n27 161.363
R18319 XThR.Tn[9] XThR.Tn[9].n22 161.363
R18320 XThR.Tn[9] XThR.Tn[9].n17 161.363
R18321 XThR.Tn[9] XThR.Tn[9].n12 161.363
R18322 XThR.Tn[9] XThR.Tn[9].n10 161.363
R18323 XThR.Tn[9].n84 XThR.Tn[9].n83 161.3
R18324 XThR.Tn[9].n79 XThR.Tn[9].n78 161.3
R18325 XThR.Tn[9].n74 XThR.Tn[9].n73 161.3
R18326 XThR.Tn[9].n69 XThR.Tn[9].n68 161.3
R18327 XThR.Tn[9].n64 XThR.Tn[9].n63 161.3
R18328 XThR.Tn[9].n59 XThR.Tn[9].n58 161.3
R18329 XThR.Tn[9].n54 XThR.Tn[9].n53 161.3
R18330 XThR.Tn[9].n49 XThR.Tn[9].n48 161.3
R18331 XThR.Tn[9].n44 XThR.Tn[9].n43 161.3
R18332 XThR.Tn[9].n39 XThR.Tn[9].n38 161.3
R18333 XThR.Tn[9].n34 XThR.Tn[9].n33 161.3
R18334 XThR.Tn[9].n29 XThR.Tn[9].n28 161.3
R18335 XThR.Tn[9].n24 XThR.Tn[9].n23 161.3
R18336 XThR.Tn[9].n19 XThR.Tn[9].n18 161.3
R18337 XThR.Tn[9].n14 XThR.Tn[9].n13 161.3
R18338 XThR.Tn[9].n82 XThR.Tn[9].t63 161.106
R18339 XThR.Tn[9].n77 XThR.Tn[9].t69 161.106
R18340 XThR.Tn[9].n72 XThR.Tn[9].t47 161.106
R18341 XThR.Tn[9].n67 XThR.Tn[9].t34 161.106
R18342 XThR.Tn[9].n62 XThR.Tn[9].t62 161.106
R18343 XThR.Tn[9].n57 XThR.Tn[9].t24 161.106
R18344 XThR.Tn[9].n52 XThR.Tn[9].t66 161.106
R18345 XThR.Tn[9].n47 XThR.Tn[9].t45 161.106
R18346 XThR.Tn[9].n42 XThR.Tn[9].t32 161.106
R18347 XThR.Tn[9].n37 XThR.Tn[9].t37 161.106
R18348 XThR.Tn[9].n32 XThR.Tn[9].t23 161.106
R18349 XThR.Tn[9].n27 XThR.Tn[9].t46 161.106
R18350 XThR.Tn[9].n22 XThR.Tn[9].t21 161.106
R18351 XThR.Tn[9].n17 XThR.Tn[9].t64 161.106
R18352 XThR.Tn[9].n12 XThR.Tn[9].t28 161.106
R18353 XThR.Tn[9].n10 XThR.Tn[9].t71 161.106
R18354 XThR.Tn[9].n83 XThR.Tn[9].t54 159.978
R18355 XThR.Tn[9].n78 XThR.Tn[9].t61 159.978
R18356 XThR.Tn[9].n73 XThR.Tn[9].t43 159.978
R18357 XThR.Tn[9].n68 XThR.Tn[9].t27 159.978
R18358 XThR.Tn[9].n63 XThR.Tn[9].t52 159.978
R18359 XThR.Tn[9].n58 XThR.Tn[9].t18 159.978
R18360 XThR.Tn[9].n53 XThR.Tn[9].t60 159.978
R18361 XThR.Tn[9].n48 XThR.Tn[9].t40 159.978
R18362 XThR.Tn[9].n43 XThR.Tn[9].t25 159.978
R18363 XThR.Tn[9].n38 XThR.Tn[9].t33 159.978
R18364 XThR.Tn[9].n33 XThR.Tn[9].t16 159.978
R18365 XThR.Tn[9].n28 XThR.Tn[9].t42 159.978
R18366 XThR.Tn[9].n23 XThR.Tn[9].t15 159.978
R18367 XThR.Tn[9].n18 XThR.Tn[9].t59 159.978
R18368 XThR.Tn[9].n13 XThR.Tn[9].t19 159.978
R18369 XThR.Tn[9].n82 XThR.Tn[9].t49 145.038
R18370 XThR.Tn[9].n77 XThR.Tn[9].t14 145.038
R18371 XThR.Tn[9].n72 XThR.Tn[9].t57 145.038
R18372 XThR.Tn[9].n67 XThR.Tn[9].t38 145.038
R18373 XThR.Tn[9].n62 XThR.Tn[9].t70 145.038
R18374 XThR.Tn[9].n57 XThR.Tn[9].t48 145.038
R18375 XThR.Tn[9].n52 XThR.Tn[9].t58 145.038
R18376 XThR.Tn[9].n47 XThR.Tn[9].t39 145.038
R18377 XThR.Tn[9].n42 XThR.Tn[9].t36 145.038
R18378 XThR.Tn[9].n37 XThR.Tn[9].t67 145.038
R18379 XThR.Tn[9].n32 XThR.Tn[9].t31 145.038
R18380 XThR.Tn[9].n27 XThR.Tn[9].t56 145.038
R18381 XThR.Tn[9].n22 XThR.Tn[9].t29 145.038
R18382 XThR.Tn[9].n17 XThR.Tn[9].t72 145.038
R18383 XThR.Tn[9].n12 XThR.Tn[9].t35 145.038
R18384 XThR.Tn[9].n10 XThR.Tn[9].t17 145.038
R18385 XThR.Tn[9].n83 XThR.Tn[9].t68 143.911
R18386 XThR.Tn[9].n78 XThR.Tn[9].t30 143.911
R18387 XThR.Tn[9].n73 XThR.Tn[9].t12 143.911
R18388 XThR.Tn[9].n68 XThR.Tn[9].t53 143.911
R18389 XThR.Tn[9].n63 XThR.Tn[9].t22 143.911
R18390 XThR.Tn[9].n58 XThR.Tn[9].t65 143.911
R18391 XThR.Tn[9].n53 XThR.Tn[9].t13 143.911
R18392 XThR.Tn[9].n48 XThR.Tn[9].t55 143.911
R18393 XThR.Tn[9].n43 XThR.Tn[9].t51 143.911
R18394 XThR.Tn[9].n38 XThR.Tn[9].t20 143.911
R18395 XThR.Tn[9].n33 XThR.Tn[9].t44 143.911
R18396 XThR.Tn[9].n28 XThR.Tn[9].t73 143.911
R18397 XThR.Tn[9].n23 XThR.Tn[9].t41 143.911
R18398 XThR.Tn[9].n18 XThR.Tn[9].t26 143.911
R18399 XThR.Tn[9].n13 XThR.Tn[9].t50 143.911
R18400 XThR.Tn[9] XThR.Tn[9].n5 35.7652
R18401 XThR.Tn[9].n6 XThR.Tn[9].t6 26.5955
R18402 XThR.Tn[9].n6 XThR.Tn[9].t4 26.5955
R18403 XThR.Tn[9].n7 XThR.Tn[9].t7 26.5955
R18404 XThR.Tn[9].n7 XThR.Tn[9].t5 26.5955
R18405 XThR.Tn[9].n3 XThR.Tn[9].t10 26.5955
R18406 XThR.Tn[9].n3 XThR.Tn[9].t8 26.5955
R18407 XThR.Tn[9].n4 XThR.Tn[9].t11 26.5955
R18408 XThR.Tn[9].n4 XThR.Tn[9].t9 26.5955
R18409 XThR.Tn[9].n0 XThR.Tn[9].t0 24.9236
R18410 XThR.Tn[9].n0 XThR.Tn[9].t2 24.9236
R18411 XThR.Tn[9].n1 XThR.Tn[9].t1 24.9236
R18412 XThR.Tn[9].n1 XThR.Tn[9].t3 24.9236
R18413 XThR.Tn[9] XThR.Tn[9].n2 22.9615
R18414 XThR.Tn[9].n9 XThR.Tn[9].n8 13.5534
R18415 XThR.Tn[9].n88 XThR.Tn[9] 7.97984
R18416 XThR.Tn[9] XThR.Tn[9].n11 5.34038
R18417 XThR.Tn[9].n16 XThR.Tn[9].n15 4.5005
R18418 XThR.Tn[9].n21 XThR.Tn[9].n20 4.5005
R18419 XThR.Tn[9].n26 XThR.Tn[9].n25 4.5005
R18420 XThR.Tn[9].n31 XThR.Tn[9].n30 4.5005
R18421 XThR.Tn[9].n36 XThR.Tn[9].n35 4.5005
R18422 XThR.Tn[9].n41 XThR.Tn[9].n40 4.5005
R18423 XThR.Tn[9].n46 XThR.Tn[9].n45 4.5005
R18424 XThR.Tn[9].n51 XThR.Tn[9].n50 4.5005
R18425 XThR.Tn[9].n56 XThR.Tn[9].n55 4.5005
R18426 XThR.Tn[9].n61 XThR.Tn[9].n60 4.5005
R18427 XThR.Tn[9].n66 XThR.Tn[9].n65 4.5005
R18428 XThR.Tn[9].n71 XThR.Tn[9].n70 4.5005
R18429 XThR.Tn[9].n76 XThR.Tn[9].n75 4.5005
R18430 XThR.Tn[9].n81 XThR.Tn[9].n80 4.5005
R18431 XThR.Tn[9].n86 XThR.Tn[9].n85 4.5005
R18432 XThR.Tn[9].n87 XThR.Tn[9] 3.70586
R18433 XThR.Tn[9].n88 XThR.Tn[9].n9 2.99115
R18434 XThR.Tn[9].n9 XThR.Tn[9] 2.87153
R18435 XThR.Tn[9].n16 XThR.Tn[9] 2.52282
R18436 XThR.Tn[9].n21 XThR.Tn[9] 2.52282
R18437 XThR.Tn[9].n26 XThR.Tn[9] 2.52282
R18438 XThR.Tn[9].n31 XThR.Tn[9] 2.52282
R18439 XThR.Tn[9].n36 XThR.Tn[9] 2.52282
R18440 XThR.Tn[9].n41 XThR.Tn[9] 2.52282
R18441 XThR.Tn[9].n46 XThR.Tn[9] 2.52282
R18442 XThR.Tn[9].n51 XThR.Tn[9] 2.52282
R18443 XThR.Tn[9].n56 XThR.Tn[9] 2.52282
R18444 XThR.Tn[9].n61 XThR.Tn[9] 2.52282
R18445 XThR.Tn[9].n66 XThR.Tn[9] 2.52282
R18446 XThR.Tn[9].n71 XThR.Tn[9] 2.52282
R18447 XThR.Tn[9].n76 XThR.Tn[9] 2.52282
R18448 XThR.Tn[9].n81 XThR.Tn[9] 2.52282
R18449 XThR.Tn[9].n86 XThR.Tn[9] 2.52282
R18450 XThR.Tn[9] XThR.Tn[9].n88 2.2734
R18451 XThR.Tn[9].n9 XThR.Tn[9] 1.50638
R18452 XThR.Tn[9].n84 XThR.Tn[9] 1.08677
R18453 XThR.Tn[9].n79 XThR.Tn[9] 1.08677
R18454 XThR.Tn[9].n74 XThR.Tn[9] 1.08677
R18455 XThR.Tn[9].n69 XThR.Tn[9] 1.08677
R18456 XThR.Tn[9].n64 XThR.Tn[9] 1.08677
R18457 XThR.Tn[9].n59 XThR.Tn[9] 1.08677
R18458 XThR.Tn[9].n54 XThR.Tn[9] 1.08677
R18459 XThR.Tn[9].n49 XThR.Tn[9] 1.08677
R18460 XThR.Tn[9].n44 XThR.Tn[9] 1.08677
R18461 XThR.Tn[9].n39 XThR.Tn[9] 1.08677
R18462 XThR.Tn[9].n34 XThR.Tn[9] 1.08677
R18463 XThR.Tn[9].n29 XThR.Tn[9] 1.08677
R18464 XThR.Tn[9].n24 XThR.Tn[9] 1.08677
R18465 XThR.Tn[9].n19 XThR.Tn[9] 1.08677
R18466 XThR.Tn[9].n14 XThR.Tn[9] 1.08677
R18467 XThR.Tn[9] XThR.Tn[9].n16 0.839786
R18468 XThR.Tn[9] XThR.Tn[9].n21 0.839786
R18469 XThR.Tn[9] XThR.Tn[9].n26 0.839786
R18470 XThR.Tn[9] XThR.Tn[9].n31 0.839786
R18471 XThR.Tn[9] XThR.Tn[9].n36 0.839786
R18472 XThR.Tn[9] XThR.Tn[9].n41 0.839786
R18473 XThR.Tn[9] XThR.Tn[9].n46 0.839786
R18474 XThR.Tn[9] XThR.Tn[9].n51 0.839786
R18475 XThR.Tn[9] XThR.Tn[9].n56 0.839786
R18476 XThR.Tn[9] XThR.Tn[9].n61 0.839786
R18477 XThR.Tn[9] XThR.Tn[9].n66 0.839786
R18478 XThR.Tn[9] XThR.Tn[9].n71 0.839786
R18479 XThR.Tn[9] XThR.Tn[9].n76 0.839786
R18480 XThR.Tn[9] XThR.Tn[9].n81 0.839786
R18481 XThR.Tn[9] XThR.Tn[9].n86 0.839786
R18482 XThR.Tn[9].n11 XThR.Tn[9] 0.499542
R18483 XThR.Tn[9].n85 XThR.Tn[9] 0.063
R18484 XThR.Tn[9].n80 XThR.Tn[9] 0.063
R18485 XThR.Tn[9].n75 XThR.Tn[9] 0.063
R18486 XThR.Tn[9].n70 XThR.Tn[9] 0.063
R18487 XThR.Tn[9].n65 XThR.Tn[9] 0.063
R18488 XThR.Tn[9].n60 XThR.Tn[9] 0.063
R18489 XThR.Tn[9].n55 XThR.Tn[9] 0.063
R18490 XThR.Tn[9].n50 XThR.Tn[9] 0.063
R18491 XThR.Tn[9].n45 XThR.Tn[9] 0.063
R18492 XThR.Tn[9].n40 XThR.Tn[9] 0.063
R18493 XThR.Tn[9].n35 XThR.Tn[9] 0.063
R18494 XThR.Tn[9].n30 XThR.Tn[9] 0.063
R18495 XThR.Tn[9].n25 XThR.Tn[9] 0.063
R18496 XThR.Tn[9].n20 XThR.Tn[9] 0.063
R18497 XThR.Tn[9].n15 XThR.Tn[9] 0.063
R18498 XThR.Tn[9].n87 XThR.Tn[9] 0.0540714
R18499 XThR.Tn[9] XThR.Tn[9].n87 0.038
R18500 XThR.Tn[9].n11 XThR.Tn[9] 0.0143889
R18501 XThR.Tn[9].n85 XThR.Tn[9].n84 0.00771154
R18502 XThR.Tn[9].n80 XThR.Tn[9].n79 0.00771154
R18503 XThR.Tn[9].n75 XThR.Tn[9].n74 0.00771154
R18504 XThR.Tn[9].n70 XThR.Tn[9].n69 0.00771154
R18505 XThR.Tn[9].n65 XThR.Tn[9].n64 0.00771154
R18506 XThR.Tn[9].n60 XThR.Tn[9].n59 0.00771154
R18507 XThR.Tn[9].n55 XThR.Tn[9].n54 0.00771154
R18508 XThR.Tn[9].n50 XThR.Tn[9].n49 0.00771154
R18509 XThR.Tn[9].n45 XThR.Tn[9].n44 0.00771154
R18510 XThR.Tn[9].n40 XThR.Tn[9].n39 0.00771154
R18511 XThR.Tn[9].n35 XThR.Tn[9].n34 0.00771154
R18512 XThR.Tn[9].n30 XThR.Tn[9].n29 0.00771154
R18513 XThR.Tn[9].n25 XThR.Tn[9].n24 0.00771154
R18514 XThR.Tn[9].n20 XThR.Tn[9].n19 0.00771154
R18515 XThR.Tn[9].n15 XThR.Tn[9].n14 0.00771154
R18516 XThC.Tn[5].n2 XThC.Tn[5].n1 332.332
R18517 XThC.Tn[5].n2 XThC.Tn[5].n0 296.493
R18518 XThC.Tn[5].n12 XThC.Tn[5].n10 161.406
R18519 XThC.Tn[5].n15 XThC.Tn[5].n13 161.406
R18520 XThC.Tn[5].n18 XThC.Tn[5].n16 161.406
R18521 XThC.Tn[5].n21 XThC.Tn[5].n19 161.406
R18522 XThC.Tn[5].n24 XThC.Tn[5].n22 161.406
R18523 XThC.Tn[5].n27 XThC.Tn[5].n25 161.406
R18524 XThC.Tn[5].n30 XThC.Tn[5].n28 161.406
R18525 XThC.Tn[5].n33 XThC.Tn[5].n31 161.406
R18526 XThC.Tn[5].n36 XThC.Tn[5].n34 161.406
R18527 XThC.Tn[5].n39 XThC.Tn[5].n37 161.406
R18528 XThC.Tn[5].n42 XThC.Tn[5].n40 161.406
R18529 XThC.Tn[5].n45 XThC.Tn[5].n43 161.406
R18530 XThC.Tn[5].n48 XThC.Tn[5].n46 161.406
R18531 XThC.Tn[5].n51 XThC.Tn[5].n49 161.406
R18532 XThC.Tn[5].n54 XThC.Tn[5].n52 161.406
R18533 XThC.Tn[5].n57 XThC.Tn[5].n55 161.406
R18534 XThC.Tn[5].n10 XThC.Tn[5].t33 161.202
R18535 XThC.Tn[5].n13 XThC.Tn[5].t19 161.202
R18536 XThC.Tn[5].n16 XThC.Tn[5].t23 161.202
R18537 XThC.Tn[5].n19 XThC.Tn[5].t24 161.202
R18538 XThC.Tn[5].n22 XThC.Tn[5].t13 161.202
R18539 XThC.Tn[5].n25 XThC.Tn[5].t14 161.202
R18540 XThC.Tn[5].n28 XThC.Tn[5].t27 161.202
R18541 XThC.Tn[5].n31 XThC.Tn[5].t35 161.202
R18542 XThC.Tn[5].n34 XThC.Tn[5].t37 161.202
R18543 XThC.Tn[5].n37 XThC.Tn[5].t25 161.202
R18544 XThC.Tn[5].n40 XThC.Tn[5].t26 161.202
R18545 XThC.Tn[5].n43 XThC.Tn[5].t39 161.202
R18546 XThC.Tn[5].n46 XThC.Tn[5].t16 161.202
R18547 XThC.Tn[5].n49 XThC.Tn[5].t18 161.202
R18548 XThC.Tn[5].n52 XThC.Tn[5].t30 161.202
R18549 XThC.Tn[5].n55 XThC.Tn[5].t41 161.202
R18550 XThC.Tn[5].n10 XThC.Tn[5].t15 145.137
R18551 XThC.Tn[5].n13 XThC.Tn[5].t34 145.137
R18552 XThC.Tn[5].n16 XThC.Tn[5].t36 145.137
R18553 XThC.Tn[5].n19 XThC.Tn[5].t38 145.137
R18554 XThC.Tn[5].n22 XThC.Tn[5].t28 145.137
R18555 XThC.Tn[5].n25 XThC.Tn[5].t29 145.137
R18556 XThC.Tn[5].n28 XThC.Tn[5].t43 145.137
R18557 XThC.Tn[5].n31 XThC.Tn[5].t17 145.137
R18558 XThC.Tn[5].n34 XThC.Tn[5].t20 145.137
R18559 XThC.Tn[5].n37 XThC.Tn[5].t40 145.137
R18560 XThC.Tn[5].n40 XThC.Tn[5].t42 145.137
R18561 XThC.Tn[5].n43 XThC.Tn[5].t21 145.137
R18562 XThC.Tn[5].n46 XThC.Tn[5].t31 145.137
R18563 XThC.Tn[5].n49 XThC.Tn[5].t32 145.137
R18564 XThC.Tn[5].n52 XThC.Tn[5].t12 145.137
R18565 XThC.Tn[5].n55 XThC.Tn[5].t22 145.137
R18566 XThC.Tn[5].n7 XThC.Tn[5].n6 135.249
R18567 XThC.Tn[5].n9 XThC.Tn[5].n3 98.981
R18568 XThC.Tn[5].n8 XThC.Tn[5].n4 98.981
R18569 XThC.Tn[5].n7 XThC.Tn[5].n5 98.981
R18570 XThC.Tn[5].n9 XThC.Tn[5].n8 36.2672
R18571 XThC.Tn[5].n8 XThC.Tn[5].n7 36.2672
R18572 XThC.Tn[5].n59 XThC.Tn[5].n9 32.6405
R18573 XThC.Tn[5].n1 XThC.Tn[5].t5 26.5955
R18574 XThC.Tn[5].n1 XThC.Tn[5].t4 26.5955
R18575 XThC.Tn[5].n0 XThC.Tn[5].t7 26.5955
R18576 XThC.Tn[5].n0 XThC.Tn[5].t6 26.5955
R18577 XThC.Tn[5].n3 XThC.Tn[5].t9 24.9236
R18578 XThC.Tn[5].n3 XThC.Tn[5].t8 24.9236
R18579 XThC.Tn[5].n4 XThC.Tn[5].t11 24.9236
R18580 XThC.Tn[5].n4 XThC.Tn[5].t10 24.9236
R18581 XThC.Tn[5].n5 XThC.Tn[5].t2 24.9236
R18582 XThC.Tn[5].n5 XThC.Tn[5].t1 24.9236
R18583 XThC.Tn[5].n6 XThC.Tn[5].t0 24.9236
R18584 XThC.Tn[5].n6 XThC.Tn[5].t3 24.9236
R18585 XThC.Tn[5] XThC.Tn[5].n2 23.3605
R18586 XThC.Tn[5] XThC.Tn[5].n59 6.7205
R18587 XThC.Tn[5].n58 XThC.Tn[5] 3.62266
R18588 XThC.Tn[5].n59 XThC.Tn[5].n58 3.18437
R18589 XThC.Tn[5].n15 XThC.Tn[5] 0.931056
R18590 XThC.Tn[5].n18 XThC.Tn[5] 0.931056
R18591 XThC.Tn[5].n21 XThC.Tn[5] 0.931056
R18592 XThC.Tn[5].n24 XThC.Tn[5] 0.931056
R18593 XThC.Tn[5].n27 XThC.Tn[5] 0.931056
R18594 XThC.Tn[5].n30 XThC.Tn[5] 0.931056
R18595 XThC.Tn[5].n33 XThC.Tn[5] 0.931056
R18596 XThC.Tn[5].n36 XThC.Tn[5] 0.931056
R18597 XThC.Tn[5].n39 XThC.Tn[5] 0.931056
R18598 XThC.Tn[5].n42 XThC.Tn[5] 0.931056
R18599 XThC.Tn[5].n45 XThC.Tn[5] 0.931056
R18600 XThC.Tn[5].n48 XThC.Tn[5] 0.931056
R18601 XThC.Tn[5].n51 XThC.Tn[5] 0.931056
R18602 XThC.Tn[5].n54 XThC.Tn[5] 0.931056
R18603 XThC.Tn[5].n57 XThC.Tn[5] 0.931056
R18604 XThC.Tn[5] XThC.Tn[5].n12 0.396333
R18605 XThC.Tn[5] XThC.Tn[5].n15 0.396333
R18606 XThC.Tn[5] XThC.Tn[5].n18 0.396333
R18607 XThC.Tn[5] XThC.Tn[5].n21 0.396333
R18608 XThC.Tn[5] XThC.Tn[5].n24 0.396333
R18609 XThC.Tn[5] XThC.Tn[5].n27 0.396333
R18610 XThC.Tn[5] XThC.Tn[5].n30 0.396333
R18611 XThC.Tn[5] XThC.Tn[5].n33 0.396333
R18612 XThC.Tn[5] XThC.Tn[5].n36 0.396333
R18613 XThC.Tn[5] XThC.Tn[5].n39 0.396333
R18614 XThC.Tn[5] XThC.Tn[5].n42 0.396333
R18615 XThC.Tn[5] XThC.Tn[5].n45 0.396333
R18616 XThC.Tn[5] XThC.Tn[5].n48 0.396333
R18617 XThC.Tn[5] XThC.Tn[5].n51 0.396333
R18618 XThC.Tn[5] XThC.Tn[5].n54 0.396333
R18619 XThC.Tn[5] XThC.Tn[5].n57 0.396333
R18620 XThC.Tn[5].n11 XThC.Tn[5] 0.104667
R18621 XThC.Tn[5].n14 XThC.Tn[5] 0.104667
R18622 XThC.Tn[5].n17 XThC.Tn[5] 0.104667
R18623 XThC.Tn[5].n20 XThC.Tn[5] 0.104667
R18624 XThC.Tn[5].n23 XThC.Tn[5] 0.104667
R18625 XThC.Tn[5].n26 XThC.Tn[5] 0.104667
R18626 XThC.Tn[5].n29 XThC.Tn[5] 0.104667
R18627 XThC.Tn[5].n32 XThC.Tn[5] 0.104667
R18628 XThC.Tn[5].n35 XThC.Tn[5] 0.104667
R18629 XThC.Tn[5].n38 XThC.Tn[5] 0.104667
R18630 XThC.Tn[5].n41 XThC.Tn[5] 0.104667
R18631 XThC.Tn[5].n44 XThC.Tn[5] 0.104667
R18632 XThC.Tn[5].n47 XThC.Tn[5] 0.104667
R18633 XThC.Tn[5].n50 XThC.Tn[5] 0.104667
R18634 XThC.Tn[5].n53 XThC.Tn[5] 0.104667
R18635 XThC.Tn[5].n56 XThC.Tn[5] 0.104667
R18636 XThC.Tn[5].n11 XThC.Tn[5] 0.0309878
R18637 XThC.Tn[5].n14 XThC.Tn[5] 0.0309878
R18638 XThC.Tn[5].n17 XThC.Tn[5] 0.0309878
R18639 XThC.Tn[5].n20 XThC.Tn[5] 0.0309878
R18640 XThC.Tn[5].n23 XThC.Tn[5] 0.0309878
R18641 XThC.Tn[5].n26 XThC.Tn[5] 0.0309878
R18642 XThC.Tn[5].n29 XThC.Tn[5] 0.0309878
R18643 XThC.Tn[5].n32 XThC.Tn[5] 0.0309878
R18644 XThC.Tn[5].n35 XThC.Tn[5] 0.0309878
R18645 XThC.Tn[5].n38 XThC.Tn[5] 0.0309878
R18646 XThC.Tn[5].n41 XThC.Tn[5] 0.0309878
R18647 XThC.Tn[5].n44 XThC.Tn[5] 0.0309878
R18648 XThC.Tn[5].n47 XThC.Tn[5] 0.0309878
R18649 XThC.Tn[5].n50 XThC.Tn[5] 0.0309878
R18650 XThC.Tn[5].n53 XThC.Tn[5] 0.0309878
R18651 XThC.Tn[5].n56 XThC.Tn[5] 0.0309878
R18652 XThC.Tn[5].n12 XThC.Tn[5].n11 0.027939
R18653 XThC.Tn[5].n15 XThC.Tn[5].n14 0.027939
R18654 XThC.Tn[5].n18 XThC.Tn[5].n17 0.027939
R18655 XThC.Tn[5].n21 XThC.Tn[5].n20 0.027939
R18656 XThC.Tn[5].n24 XThC.Tn[5].n23 0.027939
R18657 XThC.Tn[5].n27 XThC.Tn[5].n26 0.027939
R18658 XThC.Tn[5].n30 XThC.Tn[5].n29 0.027939
R18659 XThC.Tn[5].n33 XThC.Tn[5].n32 0.027939
R18660 XThC.Tn[5].n36 XThC.Tn[5].n35 0.027939
R18661 XThC.Tn[5].n39 XThC.Tn[5].n38 0.027939
R18662 XThC.Tn[5].n42 XThC.Tn[5].n41 0.027939
R18663 XThC.Tn[5].n45 XThC.Tn[5].n44 0.027939
R18664 XThC.Tn[5].n48 XThC.Tn[5].n47 0.027939
R18665 XThC.Tn[5].n51 XThC.Tn[5].n50 0.027939
R18666 XThC.Tn[5].n54 XThC.Tn[5].n53 0.027939
R18667 XThC.Tn[5].n57 XThC.Tn[5].n56 0.027939
R18668 XThC.Tn[5].n58 XThC.Tn[5] 0.0129681
R18669 XThC.Tn[9].n2 XThC.Tn[9].n1 265.341
R18670 XThC.Tn[9].n5 XThC.Tn[9].n3 243.68
R18671 XThC.Tn[9].n58 XThC.Tn[9].n56 241.847
R18672 XThC.Tn[9].n5 XThC.Tn[9].n4 205.28
R18673 XThC.Tn[9].n2 XThC.Tn[9].n0 202.094
R18674 XThC.Tn[9].n58 XThC.Tn[9].n57 185
R18675 XThC.Tn[9].n9 XThC.Tn[9].n7 161.406
R18676 XThC.Tn[9].n12 XThC.Tn[9].n10 161.406
R18677 XThC.Tn[9].n15 XThC.Tn[9].n13 161.406
R18678 XThC.Tn[9].n18 XThC.Tn[9].n16 161.406
R18679 XThC.Tn[9].n21 XThC.Tn[9].n19 161.406
R18680 XThC.Tn[9].n24 XThC.Tn[9].n22 161.406
R18681 XThC.Tn[9].n27 XThC.Tn[9].n25 161.406
R18682 XThC.Tn[9].n30 XThC.Tn[9].n28 161.406
R18683 XThC.Tn[9].n33 XThC.Tn[9].n31 161.406
R18684 XThC.Tn[9].n36 XThC.Tn[9].n34 161.406
R18685 XThC.Tn[9].n39 XThC.Tn[9].n37 161.406
R18686 XThC.Tn[9].n42 XThC.Tn[9].n40 161.406
R18687 XThC.Tn[9].n45 XThC.Tn[9].n43 161.406
R18688 XThC.Tn[9].n48 XThC.Tn[9].n46 161.406
R18689 XThC.Tn[9].n51 XThC.Tn[9].n49 161.406
R18690 XThC.Tn[9].n54 XThC.Tn[9].n52 161.406
R18691 XThC.Tn[9].n7 XThC.Tn[9].t12 161.202
R18692 XThC.Tn[9].n10 XThC.Tn[9].t30 161.202
R18693 XThC.Tn[9].n13 XThC.Tn[9].t34 161.202
R18694 XThC.Tn[9].n16 XThC.Tn[9].t35 161.202
R18695 XThC.Tn[9].n19 XThC.Tn[9].t24 161.202
R18696 XThC.Tn[9].n22 XThC.Tn[9].t25 161.202
R18697 XThC.Tn[9].n25 XThC.Tn[9].t38 161.202
R18698 XThC.Tn[9].n28 XThC.Tn[9].t14 161.202
R18699 XThC.Tn[9].n31 XThC.Tn[9].t16 161.202
R18700 XThC.Tn[9].n34 XThC.Tn[9].t36 161.202
R18701 XThC.Tn[9].n37 XThC.Tn[9].t37 161.202
R18702 XThC.Tn[9].n40 XThC.Tn[9].t18 161.202
R18703 XThC.Tn[9].n43 XThC.Tn[9].t27 161.202
R18704 XThC.Tn[9].n46 XThC.Tn[9].t29 161.202
R18705 XThC.Tn[9].n49 XThC.Tn[9].t41 161.202
R18706 XThC.Tn[9].n52 XThC.Tn[9].t20 161.202
R18707 XThC.Tn[9].n7 XThC.Tn[9].t26 145.137
R18708 XThC.Tn[9].n10 XThC.Tn[9].t13 145.137
R18709 XThC.Tn[9].n13 XThC.Tn[9].t15 145.137
R18710 XThC.Tn[9].n16 XThC.Tn[9].t17 145.137
R18711 XThC.Tn[9].n19 XThC.Tn[9].t39 145.137
R18712 XThC.Tn[9].n22 XThC.Tn[9].t40 145.137
R18713 XThC.Tn[9].n25 XThC.Tn[9].t22 145.137
R18714 XThC.Tn[9].n28 XThC.Tn[9].t28 145.137
R18715 XThC.Tn[9].n31 XThC.Tn[9].t31 145.137
R18716 XThC.Tn[9].n34 XThC.Tn[9].t19 145.137
R18717 XThC.Tn[9].n37 XThC.Tn[9].t21 145.137
R18718 XThC.Tn[9].n40 XThC.Tn[9].t32 145.137
R18719 XThC.Tn[9].n43 XThC.Tn[9].t42 145.137
R18720 XThC.Tn[9].n46 XThC.Tn[9].t43 145.137
R18721 XThC.Tn[9].n49 XThC.Tn[9].t23 145.137
R18722 XThC.Tn[9].n52 XThC.Tn[9].t33 145.137
R18723 XThC.Tn[9].n1 XThC.Tn[9].t6 26.5955
R18724 XThC.Tn[9].n1 XThC.Tn[9].t5 26.5955
R18725 XThC.Tn[9].n0 XThC.Tn[9].t4 26.5955
R18726 XThC.Tn[9].n0 XThC.Tn[9].t7 26.5955
R18727 XThC.Tn[9].n3 XThC.Tn[9].t9 26.5955
R18728 XThC.Tn[9].n3 XThC.Tn[9].t8 26.5955
R18729 XThC.Tn[9].n4 XThC.Tn[9].t11 26.5955
R18730 XThC.Tn[9].n4 XThC.Tn[9].t10 26.5955
R18731 XThC.Tn[9].n56 XThC.Tn[9].t1 24.9236
R18732 XThC.Tn[9].n56 XThC.Tn[9].t0 24.9236
R18733 XThC.Tn[9].n57 XThC.Tn[9].t2 24.9236
R18734 XThC.Tn[9].n57 XThC.Tn[9].t3 24.9236
R18735 XThC.Tn[9] XThC.Tn[9].n5 22.9652
R18736 XThC.Tn[9] XThC.Tn[9].n58 18.8943
R18737 XThC.Tn[9].n6 XThC.Tn[9].n2 13.9299
R18738 XThC.Tn[9].n6 XThC.Tn[9] 13.9299
R18739 XThC.Tn[9] XThC.Tn[9].n55 6.34069
R18740 XThC.Tn[9].n55 XThC.Tn[9] 5.13485
R18741 XThC.Tn[9].n55 XThC.Tn[9] 1.79489
R18742 XThC.Tn[9] XThC.Tn[9].n6 1.19676
R18743 XThC.Tn[9].n12 XThC.Tn[9] 0.931056
R18744 XThC.Tn[9].n15 XThC.Tn[9] 0.931056
R18745 XThC.Tn[9].n18 XThC.Tn[9] 0.931056
R18746 XThC.Tn[9].n21 XThC.Tn[9] 0.931056
R18747 XThC.Tn[9].n24 XThC.Tn[9] 0.931056
R18748 XThC.Tn[9].n27 XThC.Tn[9] 0.931056
R18749 XThC.Tn[9].n30 XThC.Tn[9] 0.931056
R18750 XThC.Tn[9].n33 XThC.Tn[9] 0.931056
R18751 XThC.Tn[9].n36 XThC.Tn[9] 0.931056
R18752 XThC.Tn[9].n39 XThC.Tn[9] 0.931056
R18753 XThC.Tn[9].n42 XThC.Tn[9] 0.931056
R18754 XThC.Tn[9].n45 XThC.Tn[9] 0.931056
R18755 XThC.Tn[9].n48 XThC.Tn[9] 0.931056
R18756 XThC.Tn[9].n51 XThC.Tn[9] 0.931056
R18757 XThC.Tn[9].n54 XThC.Tn[9] 0.931056
R18758 XThC.Tn[9] XThC.Tn[9].n9 0.396333
R18759 XThC.Tn[9] XThC.Tn[9].n12 0.396333
R18760 XThC.Tn[9] XThC.Tn[9].n15 0.396333
R18761 XThC.Tn[9] XThC.Tn[9].n18 0.396333
R18762 XThC.Tn[9] XThC.Tn[9].n21 0.396333
R18763 XThC.Tn[9] XThC.Tn[9].n24 0.396333
R18764 XThC.Tn[9] XThC.Tn[9].n27 0.396333
R18765 XThC.Tn[9] XThC.Tn[9].n30 0.396333
R18766 XThC.Tn[9] XThC.Tn[9].n33 0.396333
R18767 XThC.Tn[9] XThC.Tn[9].n36 0.396333
R18768 XThC.Tn[9] XThC.Tn[9].n39 0.396333
R18769 XThC.Tn[9] XThC.Tn[9].n42 0.396333
R18770 XThC.Tn[9] XThC.Tn[9].n45 0.396333
R18771 XThC.Tn[9] XThC.Tn[9].n48 0.396333
R18772 XThC.Tn[9] XThC.Tn[9].n51 0.396333
R18773 XThC.Tn[9] XThC.Tn[9].n54 0.396333
R18774 XThC.Tn[9].n8 XThC.Tn[9] 0.104667
R18775 XThC.Tn[9].n11 XThC.Tn[9] 0.104667
R18776 XThC.Tn[9].n14 XThC.Tn[9] 0.104667
R18777 XThC.Tn[9].n17 XThC.Tn[9] 0.104667
R18778 XThC.Tn[9].n20 XThC.Tn[9] 0.104667
R18779 XThC.Tn[9].n23 XThC.Tn[9] 0.104667
R18780 XThC.Tn[9].n26 XThC.Tn[9] 0.104667
R18781 XThC.Tn[9].n29 XThC.Tn[9] 0.104667
R18782 XThC.Tn[9].n32 XThC.Tn[9] 0.104667
R18783 XThC.Tn[9].n35 XThC.Tn[9] 0.104667
R18784 XThC.Tn[9].n38 XThC.Tn[9] 0.104667
R18785 XThC.Tn[9].n41 XThC.Tn[9] 0.104667
R18786 XThC.Tn[9].n44 XThC.Tn[9] 0.104667
R18787 XThC.Tn[9].n47 XThC.Tn[9] 0.104667
R18788 XThC.Tn[9].n50 XThC.Tn[9] 0.104667
R18789 XThC.Tn[9].n53 XThC.Tn[9] 0.104667
R18790 XThC.Tn[9].n8 XThC.Tn[9] 0.0309878
R18791 XThC.Tn[9].n11 XThC.Tn[9] 0.0309878
R18792 XThC.Tn[9].n14 XThC.Tn[9] 0.0309878
R18793 XThC.Tn[9].n17 XThC.Tn[9] 0.0309878
R18794 XThC.Tn[9].n20 XThC.Tn[9] 0.0309878
R18795 XThC.Tn[9].n23 XThC.Tn[9] 0.0309878
R18796 XThC.Tn[9].n26 XThC.Tn[9] 0.0309878
R18797 XThC.Tn[9].n29 XThC.Tn[9] 0.0309878
R18798 XThC.Tn[9].n32 XThC.Tn[9] 0.0309878
R18799 XThC.Tn[9].n35 XThC.Tn[9] 0.0309878
R18800 XThC.Tn[9].n38 XThC.Tn[9] 0.0309878
R18801 XThC.Tn[9].n41 XThC.Tn[9] 0.0309878
R18802 XThC.Tn[9].n44 XThC.Tn[9] 0.0309878
R18803 XThC.Tn[9].n47 XThC.Tn[9] 0.0309878
R18804 XThC.Tn[9].n50 XThC.Tn[9] 0.0309878
R18805 XThC.Tn[9].n53 XThC.Tn[9] 0.0309878
R18806 XThC.Tn[9].n9 XThC.Tn[9].n8 0.027939
R18807 XThC.Tn[9].n12 XThC.Tn[9].n11 0.027939
R18808 XThC.Tn[9].n15 XThC.Tn[9].n14 0.027939
R18809 XThC.Tn[9].n18 XThC.Tn[9].n17 0.027939
R18810 XThC.Tn[9].n21 XThC.Tn[9].n20 0.027939
R18811 XThC.Tn[9].n24 XThC.Tn[9].n23 0.027939
R18812 XThC.Tn[9].n27 XThC.Tn[9].n26 0.027939
R18813 XThC.Tn[9].n30 XThC.Tn[9].n29 0.027939
R18814 XThC.Tn[9].n33 XThC.Tn[9].n32 0.027939
R18815 XThC.Tn[9].n36 XThC.Tn[9].n35 0.027939
R18816 XThC.Tn[9].n39 XThC.Tn[9].n38 0.027939
R18817 XThC.Tn[9].n42 XThC.Tn[9].n41 0.027939
R18818 XThC.Tn[9].n45 XThC.Tn[9].n44 0.027939
R18819 XThC.Tn[9].n48 XThC.Tn[9].n47 0.027939
R18820 XThC.Tn[9].n51 XThC.Tn[9].n50 0.027939
R18821 XThC.Tn[9].n54 XThC.Tn[9].n53 0.027939
R18822 XThC.Tn[11].n54 XThC.Tn[11].n53 265.341
R18823 XThC.Tn[11].n58 XThC.Tn[11].n56 243.68
R18824 XThC.Tn[11].n2 XThC.Tn[11].n0 241.847
R18825 XThC.Tn[11].n58 XThC.Tn[11].n57 205.28
R18826 XThC.Tn[11].n54 XThC.Tn[11].n52 202.094
R18827 XThC.Tn[11].n2 XThC.Tn[11].n1 185
R18828 XThC.Tn[11].n5 XThC.Tn[11].n3 161.406
R18829 XThC.Tn[11].n8 XThC.Tn[11].n6 161.406
R18830 XThC.Tn[11].n11 XThC.Tn[11].n9 161.406
R18831 XThC.Tn[11].n14 XThC.Tn[11].n12 161.406
R18832 XThC.Tn[11].n17 XThC.Tn[11].n15 161.406
R18833 XThC.Tn[11].n20 XThC.Tn[11].n18 161.406
R18834 XThC.Tn[11].n23 XThC.Tn[11].n21 161.406
R18835 XThC.Tn[11].n26 XThC.Tn[11].n24 161.406
R18836 XThC.Tn[11].n29 XThC.Tn[11].n27 161.406
R18837 XThC.Tn[11].n32 XThC.Tn[11].n30 161.406
R18838 XThC.Tn[11].n35 XThC.Tn[11].n33 161.406
R18839 XThC.Tn[11].n38 XThC.Tn[11].n36 161.406
R18840 XThC.Tn[11].n41 XThC.Tn[11].n39 161.406
R18841 XThC.Tn[11].n44 XThC.Tn[11].n42 161.406
R18842 XThC.Tn[11].n47 XThC.Tn[11].n45 161.406
R18843 XThC.Tn[11].n50 XThC.Tn[11].n48 161.406
R18844 XThC.Tn[11].n3 XThC.Tn[11].t18 161.202
R18845 XThC.Tn[11].n6 XThC.Tn[11].t35 161.202
R18846 XThC.Tn[11].n9 XThC.Tn[11].t37 161.202
R18847 XThC.Tn[11].n12 XThC.Tn[11].t39 161.202
R18848 XThC.Tn[11].n15 XThC.Tn[11].t28 161.202
R18849 XThC.Tn[11].n18 XThC.Tn[11].t29 161.202
R18850 XThC.Tn[11].n21 XThC.Tn[11].t42 161.202
R18851 XThC.Tn[11].n24 XThC.Tn[11].t19 161.202
R18852 XThC.Tn[11].n27 XThC.Tn[11].t21 161.202
R18853 XThC.Tn[11].n30 XThC.Tn[11].t40 161.202
R18854 XThC.Tn[11].n33 XThC.Tn[11].t41 161.202
R18855 XThC.Tn[11].n36 XThC.Tn[11].t22 161.202
R18856 XThC.Tn[11].n39 XThC.Tn[11].t30 161.202
R18857 XThC.Tn[11].n42 XThC.Tn[11].t33 161.202
R18858 XThC.Tn[11].n45 XThC.Tn[11].t14 161.202
R18859 XThC.Tn[11].n48 XThC.Tn[11].t24 161.202
R18860 XThC.Tn[11].n3 XThC.Tn[11].t20 145.137
R18861 XThC.Tn[11].n6 XThC.Tn[11].t38 145.137
R18862 XThC.Tn[11].n9 XThC.Tn[11].t43 145.137
R18863 XThC.Tn[11].n12 XThC.Tn[11].t12 145.137
R18864 XThC.Tn[11].n15 XThC.Tn[11].t31 145.137
R18865 XThC.Tn[11].n18 XThC.Tn[11].t32 145.137
R18866 XThC.Tn[11].n21 XThC.Tn[11].t16 145.137
R18867 XThC.Tn[11].n24 XThC.Tn[11].t23 145.137
R18868 XThC.Tn[11].n27 XThC.Tn[11].t25 145.137
R18869 XThC.Tn[11].n30 XThC.Tn[11].t13 145.137
R18870 XThC.Tn[11].n33 XThC.Tn[11].t15 145.137
R18871 XThC.Tn[11].n36 XThC.Tn[11].t26 145.137
R18872 XThC.Tn[11].n39 XThC.Tn[11].t34 145.137
R18873 XThC.Tn[11].n42 XThC.Tn[11].t36 145.137
R18874 XThC.Tn[11].n45 XThC.Tn[11].t17 145.137
R18875 XThC.Tn[11].n48 XThC.Tn[11].t27 145.137
R18876 XThC.Tn[11].n52 XThC.Tn[11].t8 26.5955
R18877 XThC.Tn[11].n52 XThC.Tn[11].t5 26.5955
R18878 XThC.Tn[11].n56 XThC.Tn[11].t1 26.5955
R18879 XThC.Tn[11].n56 XThC.Tn[11].t4 26.5955
R18880 XThC.Tn[11].n57 XThC.Tn[11].t3 26.5955
R18881 XThC.Tn[11].n57 XThC.Tn[11].t2 26.5955
R18882 XThC.Tn[11].n53 XThC.Tn[11].t0 26.5955
R18883 XThC.Tn[11].n53 XThC.Tn[11].t11 26.5955
R18884 XThC.Tn[11].n1 XThC.Tn[11].t9 24.9236
R18885 XThC.Tn[11].n1 XThC.Tn[11].t7 24.9236
R18886 XThC.Tn[11].n0 XThC.Tn[11].t10 24.9236
R18887 XThC.Tn[11].n0 XThC.Tn[11].t6 24.9236
R18888 XThC.Tn[11] XThC.Tn[11].n58 22.9652
R18889 XThC.Tn[11] XThC.Tn[11].n2 18.8943
R18890 XThC.Tn[11].n55 XThC.Tn[11].n54 13.9299
R18891 XThC.Tn[11] XThC.Tn[11].n55 13.9299
R18892 XThC.Tn[11].n51 XThC.Tn[11] 6.34069
R18893 XThC.Tn[11].n51 XThC.Tn[11] 5.13485
R18894 XThC.Tn[11] XThC.Tn[11].n51 1.79489
R18895 XThC.Tn[11].n55 XThC.Tn[11] 1.19676
R18896 XThC.Tn[11].n8 XThC.Tn[11] 0.931056
R18897 XThC.Tn[11].n11 XThC.Tn[11] 0.931056
R18898 XThC.Tn[11].n14 XThC.Tn[11] 0.931056
R18899 XThC.Tn[11].n17 XThC.Tn[11] 0.931056
R18900 XThC.Tn[11].n20 XThC.Tn[11] 0.931056
R18901 XThC.Tn[11].n23 XThC.Tn[11] 0.931056
R18902 XThC.Tn[11].n26 XThC.Tn[11] 0.931056
R18903 XThC.Tn[11].n29 XThC.Tn[11] 0.931056
R18904 XThC.Tn[11].n32 XThC.Tn[11] 0.931056
R18905 XThC.Tn[11].n35 XThC.Tn[11] 0.931056
R18906 XThC.Tn[11].n38 XThC.Tn[11] 0.931056
R18907 XThC.Tn[11].n41 XThC.Tn[11] 0.931056
R18908 XThC.Tn[11].n44 XThC.Tn[11] 0.931056
R18909 XThC.Tn[11].n47 XThC.Tn[11] 0.931056
R18910 XThC.Tn[11].n50 XThC.Tn[11] 0.931056
R18911 XThC.Tn[11] XThC.Tn[11].n5 0.396333
R18912 XThC.Tn[11] XThC.Tn[11].n8 0.396333
R18913 XThC.Tn[11] XThC.Tn[11].n11 0.396333
R18914 XThC.Tn[11] XThC.Tn[11].n14 0.396333
R18915 XThC.Tn[11] XThC.Tn[11].n17 0.396333
R18916 XThC.Tn[11] XThC.Tn[11].n20 0.396333
R18917 XThC.Tn[11] XThC.Tn[11].n23 0.396333
R18918 XThC.Tn[11] XThC.Tn[11].n26 0.396333
R18919 XThC.Tn[11] XThC.Tn[11].n29 0.396333
R18920 XThC.Tn[11] XThC.Tn[11].n32 0.396333
R18921 XThC.Tn[11] XThC.Tn[11].n35 0.396333
R18922 XThC.Tn[11] XThC.Tn[11].n38 0.396333
R18923 XThC.Tn[11] XThC.Tn[11].n41 0.396333
R18924 XThC.Tn[11] XThC.Tn[11].n44 0.396333
R18925 XThC.Tn[11] XThC.Tn[11].n47 0.396333
R18926 XThC.Tn[11] XThC.Tn[11].n50 0.396333
R18927 XThC.Tn[11].n4 XThC.Tn[11] 0.104667
R18928 XThC.Tn[11].n7 XThC.Tn[11] 0.104667
R18929 XThC.Tn[11].n10 XThC.Tn[11] 0.104667
R18930 XThC.Tn[11].n13 XThC.Tn[11] 0.104667
R18931 XThC.Tn[11].n16 XThC.Tn[11] 0.104667
R18932 XThC.Tn[11].n19 XThC.Tn[11] 0.104667
R18933 XThC.Tn[11].n22 XThC.Tn[11] 0.104667
R18934 XThC.Tn[11].n25 XThC.Tn[11] 0.104667
R18935 XThC.Tn[11].n28 XThC.Tn[11] 0.104667
R18936 XThC.Tn[11].n31 XThC.Tn[11] 0.104667
R18937 XThC.Tn[11].n34 XThC.Tn[11] 0.104667
R18938 XThC.Tn[11].n37 XThC.Tn[11] 0.104667
R18939 XThC.Tn[11].n40 XThC.Tn[11] 0.104667
R18940 XThC.Tn[11].n43 XThC.Tn[11] 0.104667
R18941 XThC.Tn[11].n46 XThC.Tn[11] 0.104667
R18942 XThC.Tn[11].n49 XThC.Tn[11] 0.104667
R18943 XThC.Tn[11].n4 XThC.Tn[11] 0.0309878
R18944 XThC.Tn[11].n7 XThC.Tn[11] 0.0309878
R18945 XThC.Tn[11].n10 XThC.Tn[11] 0.0309878
R18946 XThC.Tn[11].n13 XThC.Tn[11] 0.0309878
R18947 XThC.Tn[11].n16 XThC.Tn[11] 0.0309878
R18948 XThC.Tn[11].n19 XThC.Tn[11] 0.0309878
R18949 XThC.Tn[11].n22 XThC.Tn[11] 0.0309878
R18950 XThC.Tn[11].n25 XThC.Tn[11] 0.0309878
R18951 XThC.Tn[11].n28 XThC.Tn[11] 0.0309878
R18952 XThC.Tn[11].n31 XThC.Tn[11] 0.0309878
R18953 XThC.Tn[11].n34 XThC.Tn[11] 0.0309878
R18954 XThC.Tn[11].n37 XThC.Tn[11] 0.0309878
R18955 XThC.Tn[11].n40 XThC.Tn[11] 0.0309878
R18956 XThC.Tn[11].n43 XThC.Tn[11] 0.0309878
R18957 XThC.Tn[11].n46 XThC.Tn[11] 0.0309878
R18958 XThC.Tn[11].n49 XThC.Tn[11] 0.0309878
R18959 XThC.Tn[11].n5 XThC.Tn[11].n4 0.027939
R18960 XThC.Tn[11].n8 XThC.Tn[11].n7 0.027939
R18961 XThC.Tn[11].n11 XThC.Tn[11].n10 0.027939
R18962 XThC.Tn[11].n14 XThC.Tn[11].n13 0.027939
R18963 XThC.Tn[11].n17 XThC.Tn[11].n16 0.027939
R18964 XThC.Tn[11].n20 XThC.Tn[11].n19 0.027939
R18965 XThC.Tn[11].n23 XThC.Tn[11].n22 0.027939
R18966 XThC.Tn[11].n26 XThC.Tn[11].n25 0.027939
R18967 XThC.Tn[11].n29 XThC.Tn[11].n28 0.027939
R18968 XThC.Tn[11].n32 XThC.Tn[11].n31 0.027939
R18969 XThC.Tn[11].n35 XThC.Tn[11].n34 0.027939
R18970 XThC.Tn[11].n38 XThC.Tn[11].n37 0.027939
R18971 XThC.Tn[11].n41 XThC.Tn[11].n40 0.027939
R18972 XThC.Tn[11].n44 XThC.Tn[11].n43 0.027939
R18973 XThC.Tn[11].n47 XThC.Tn[11].n46 0.027939
R18974 XThC.Tn[11].n50 XThC.Tn[11].n49 0.027939
R18975 XThC.Tn[12].n5 XThC.Tn[12].n4 256.104
R18976 XThC.Tn[12].n8 XThC.Tn[12].n6 243.68
R18977 XThC.Tn[12].n2 XThC.Tn[12].n1 241.847
R18978 XThC.Tn[12].n8 XThC.Tn[12].n7 205.28
R18979 XThC.Tn[12].n5 XThC.Tn[12].n3 202.095
R18980 XThC.Tn[12].n2 XThC.Tn[12].n0 185
R18981 XThC.Tn[12].n12 XThC.Tn[12].n10 161.406
R18982 XThC.Tn[12].n15 XThC.Tn[12].n13 161.406
R18983 XThC.Tn[12].n18 XThC.Tn[12].n16 161.406
R18984 XThC.Tn[12].n21 XThC.Tn[12].n19 161.406
R18985 XThC.Tn[12].n24 XThC.Tn[12].n22 161.406
R18986 XThC.Tn[12].n27 XThC.Tn[12].n25 161.406
R18987 XThC.Tn[12].n30 XThC.Tn[12].n28 161.406
R18988 XThC.Tn[12].n33 XThC.Tn[12].n31 161.406
R18989 XThC.Tn[12].n36 XThC.Tn[12].n34 161.406
R18990 XThC.Tn[12].n39 XThC.Tn[12].n37 161.406
R18991 XThC.Tn[12].n42 XThC.Tn[12].n40 161.406
R18992 XThC.Tn[12].n45 XThC.Tn[12].n43 161.406
R18993 XThC.Tn[12].n48 XThC.Tn[12].n46 161.406
R18994 XThC.Tn[12].n51 XThC.Tn[12].n49 161.406
R18995 XThC.Tn[12].n54 XThC.Tn[12].n52 161.406
R18996 XThC.Tn[12].n57 XThC.Tn[12].n55 161.406
R18997 XThC.Tn[12].n10 XThC.Tn[12].t35 161.202
R18998 XThC.Tn[12].n13 XThC.Tn[12].t20 161.202
R18999 XThC.Tn[12].n16 XThC.Tn[12].t22 161.202
R19000 XThC.Tn[12].n19 XThC.Tn[12].t24 161.202
R19001 XThC.Tn[12].n22 XThC.Tn[12].t13 161.202
R19002 XThC.Tn[12].n25 XThC.Tn[12].t14 161.202
R19003 XThC.Tn[12].n28 XThC.Tn[12].t27 161.202
R19004 XThC.Tn[12].n31 XThC.Tn[12].t36 161.202
R19005 XThC.Tn[12].n34 XThC.Tn[12].t38 161.202
R19006 XThC.Tn[12].n37 XThC.Tn[12].t25 161.202
R19007 XThC.Tn[12].n40 XThC.Tn[12].t26 161.202
R19008 XThC.Tn[12].n43 XThC.Tn[12].t39 161.202
R19009 XThC.Tn[12].n46 XThC.Tn[12].t15 161.202
R19010 XThC.Tn[12].n49 XThC.Tn[12].t18 161.202
R19011 XThC.Tn[12].n52 XThC.Tn[12].t31 161.202
R19012 XThC.Tn[12].n55 XThC.Tn[12].t41 161.202
R19013 XThC.Tn[12].n10 XThC.Tn[12].t37 145.137
R19014 XThC.Tn[12].n13 XThC.Tn[12].t23 145.137
R19015 XThC.Tn[12].n16 XThC.Tn[12].t28 145.137
R19016 XThC.Tn[12].n19 XThC.Tn[12].t29 145.137
R19017 XThC.Tn[12].n22 XThC.Tn[12].t16 145.137
R19018 XThC.Tn[12].n25 XThC.Tn[12].t17 145.137
R19019 XThC.Tn[12].n28 XThC.Tn[12].t33 145.137
R19020 XThC.Tn[12].n31 XThC.Tn[12].t40 145.137
R19021 XThC.Tn[12].n34 XThC.Tn[12].t42 145.137
R19022 XThC.Tn[12].n37 XThC.Tn[12].t30 145.137
R19023 XThC.Tn[12].n40 XThC.Tn[12].t32 145.137
R19024 XThC.Tn[12].n43 XThC.Tn[12].t43 145.137
R19025 XThC.Tn[12].n46 XThC.Tn[12].t19 145.137
R19026 XThC.Tn[12].n49 XThC.Tn[12].t21 145.137
R19027 XThC.Tn[12].n52 XThC.Tn[12].t34 145.137
R19028 XThC.Tn[12].n55 XThC.Tn[12].t12 145.137
R19029 XThC.Tn[12].n3 XThC.Tn[12].t5 26.5955
R19030 XThC.Tn[12].n3 XThC.Tn[12].t6 26.5955
R19031 XThC.Tn[12].n4 XThC.Tn[12].t4 26.5955
R19032 XThC.Tn[12].n4 XThC.Tn[12].t7 26.5955
R19033 XThC.Tn[12].n6 XThC.Tn[12].t9 26.5955
R19034 XThC.Tn[12].n6 XThC.Tn[12].t8 26.5955
R19035 XThC.Tn[12].n7 XThC.Tn[12].t11 26.5955
R19036 XThC.Tn[12].n7 XThC.Tn[12].t10 26.5955
R19037 XThC.Tn[12].n0 XThC.Tn[12].t1 24.9236
R19038 XThC.Tn[12].n0 XThC.Tn[12].t0 24.9236
R19039 XThC.Tn[12].n1 XThC.Tn[12].t3 24.9236
R19040 XThC.Tn[12].n1 XThC.Tn[12].t2 24.9236
R19041 XThC.Tn[12] XThC.Tn[12].n8 22.9652
R19042 XThC.Tn[12] XThC.Tn[12].n2 22.9615
R19043 XThC.Tn[12].n9 XThC.Tn[12].n5 13.9299
R19044 XThC.Tn[12].n9 XThC.Tn[12] 13.9299
R19045 XThC.Tn[12].n59 XThC.Tn[12].n58 5.13244
R19046 XThC.Tn[12].n58 XThC.Tn[12] 3.8444
R19047 XThC.Tn[12].n59 XThC.Tn[12].n9 2.99115
R19048 XThC.Tn[12].n9 XThC.Tn[12] 2.87153
R19049 XThC.Tn[12] XThC.Tn[12].n59 2.2734
R19050 XThC.Tn[12].n15 XThC.Tn[12] 0.931056
R19051 XThC.Tn[12].n18 XThC.Tn[12] 0.931056
R19052 XThC.Tn[12].n21 XThC.Tn[12] 0.931056
R19053 XThC.Tn[12].n24 XThC.Tn[12] 0.931056
R19054 XThC.Tn[12].n27 XThC.Tn[12] 0.931056
R19055 XThC.Tn[12].n30 XThC.Tn[12] 0.931056
R19056 XThC.Tn[12].n33 XThC.Tn[12] 0.931056
R19057 XThC.Tn[12].n36 XThC.Tn[12] 0.931056
R19058 XThC.Tn[12].n39 XThC.Tn[12] 0.931056
R19059 XThC.Tn[12].n42 XThC.Tn[12] 0.931056
R19060 XThC.Tn[12].n45 XThC.Tn[12] 0.931056
R19061 XThC.Tn[12].n48 XThC.Tn[12] 0.931056
R19062 XThC.Tn[12].n51 XThC.Tn[12] 0.931056
R19063 XThC.Tn[12].n54 XThC.Tn[12] 0.931056
R19064 XThC.Tn[12].n57 XThC.Tn[12] 0.931056
R19065 XThC.Tn[12] XThC.Tn[12].n12 0.396333
R19066 XThC.Tn[12] XThC.Tn[12].n15 0.396333
R19067 XThC.Tn[12] XThC.Tn[12].n18 0.396333
R19068 XThC.Tn[12] XThC.Tn[12].n21 0.396333
R19069 XThC.Tn[12] XThC.Tn[12].n24 0.396333
R19070 XThC.Tn[12] XThC.Tn[12].n27 0.396333
R19071 XThC.Tn[12] XThC.Tn[12].n30 0.396333
R19072 XThC.Tn[12] XThC.Tn[12].n33 0.396333
R19073 XThC.Tn[12] XThC.Tn[12].n36 0.396333
R19074 XThC.Tn[12] XThC.Tn[12].n39 0.396333
R19075 XThC.Tn[12] XThC.Tn[12].n42 0.396333
R19076 XThC.Tn[12] XThC.Tn[12].n45 0.396333
R19077 XThC.Tn[12] XThC.Tn[12].n48 0.396333
R19078 XThC.Tn[12] XThC.Tn[12].n51 0.396333
R19079 XThC.Tn[12] XThC.Tn[12].n54 0.396333
R19080 XThC.Tn[12] XThC.Tn[12].n57 0.396333
R19081 XThC.Tn[12].n11 XThC.Tn[12] 0.104667
R19082 XThC.Tn[12].n14 XThC.Tn[12] 0.104667
R19083 XThC.Tn[12].n17 XThC.Tn[12] 0.104667
R19084 XThC.Tn[12].n20 XThC.Tn[12] 0.104667
R19085 XThC.Tn[12].n23 XThC.Tn[12] 0.104667
R19086 XThC.Tn[12].n26 XThC.Tn[12] 0.104667
R19087 XThC.Tn[12].n29 XThC.Tn[12] 0.104667
R19088 XThC.Tn[12].n32 XThC.Tn[12] 0.104667
R19089 XThC.Tn[12].n35 XThC.Tn[12] 0.104667
R19090 XThC.Tn[12].n38 XThC.Tn[12] 0.104667
R19091 XThC.Tn[12].n41 XThC.Tn[12] 0.104667
R19092 XThC.Tn[12].n44 XThC.Tn[12] 0.104667
R19093 XThC.Tn[12].n47 XThC.Tn[12] 0.104667
R19094 XThC.Tn[12].n50 XThC.Tn[12] 0.104667
R19095 XThC.Tn[12].n53 XThC.Tn[12] 0.104667
R19096 XThC.Tn[12].n56 XThC.Tn[12] 0.104667
R19097 XThC.Tn[12].n11 XThC.Tn[12] 0.0309878
R19098 XThC.Tn[12].n14 XThC.Tn[12] 0.0309878
R19099 XThC.Tn[12].n17 XThC.Tn[12] 0.0309878
R19100 XThC.Tn[12].n20 XThC.Tn[12] 0.0309878
R19101 XThC.Tn[12].n23 XThC.Tn[12] 0.0309878
R19102 XThC.Tn[12].n26 XThC.Tn[12] 0.0309878
R19103 XThC.Tn[12].n29 XThC.Tn[12] 0.0309878
R19104 XThC.Tn[12].n32 XThC.Tn[12] 0.0309878
R19105 XThC.Tn[12].n35 XThC.Tn[12] 0.0309878
R19106 XThC.Tn[12].n38 XThC.Tn[12] 0.0309878
R19107 XThC.Tn[12].n41 XThC.Tn[12] 0.0309878
R19108 XThC.Tn[12].n44 XThC.Tn[12] 0.0309878
R19109 XThC.Tn[12].n47 XThC.Tn[12] 0.0309878
R19110 XThC.Tn[12].n50 XThC.Tn[12] 0.0309878
R19111 XThC.Tn[12].n53 XThC.Tn[12] 0.0309878
R19112 XThC.Tn[12].n56 XThC.Tn[12] 0.0309878
R19113 XThC.Tn[12].n12 XThC.Tn[12].n11 0.027939
R19114 XThC.Tn[12].n15 XThC.Tn[12].n14 0.027939
R19115 XThC.Tn[12].n18 XThC.Tn[12].n17 0.027939
R19116 XThC.Tn[12].n21 XThC.Tn[12].n20 0.027939
R19117 XThC.Tn[12].n24 XThC.Tn[12].n23 0.027939
R19118 XThC.Tn[12].n27 XThC.Tn[12].n26 0.027939
R19119 XThC.Tn[12].n30 XThC.Tn[12].n29 0.027939
R19120 XThC.Tn[12].n33 XThC.Tn[12].n32 0.027939
R19121 XThC.Tn[12].n36 XThC.Tn[12].n35 0.027939
R19122 XThC.Tn[12].n39 XThC.Tn[12].n38 0.027939
R19123 XThC.Tn[12].n42 XThC.Tn[12].n41 0.027939
R19124 XThC.Tn[12].n45 XThC.Tn[12].n44 0.027939
R19125 XThC.Tn[12].n48 XThC.Tn[12].n47 0.027939
R19126 XThC.Tn[12].n51 XThC.Tn[12].n50 0.027939
R19127 XThC.Tn[12].n54 XThC.Tn[12].n53 0.027939
R19128 XThC.Tn[12].n57 XThC.Tn[12].n56 0.027939
R19129 XThC.Tn[12].n58 XThC.Tn[12] 0.00316553
R19130 XThC.Tn[13].n2 XThC.Tn[13].n1 265.341
R19131 XThC.Tn[13].n5 XThC.Tn[13].n3 243.68
R19132 XThC.Tn[13].n59 XThC.Tn[13].n58 241.847
R19133 XThC.Tn[13].n5 XThC.Tn[13].n4 205.28
R19134 XThC.Tn[13].n2 XThC.Tn[13].n0 202.094
R19135 XThC.Tn[13].n59 XThC.Tn[13].n57 185
R19136 XThC.Tn[13].n9 XThC.Tn[13].n7 161.406
R19137 XThC.Tn[13].n12 XThC.Tn[13].n10 161.406
R19138 XThC.Tn[13].n15 XThC.Tn[13].n13 161.406
R19139 XThC.Tn[13].n18 XThC.Tn[13].n16 161.406
R19140 XThC.Tn[13].n21 XThC.Tn[13].n19 161.406
R19141 XThC.Tn[13].n24 XThC.Tn[13].n22 161.406
R19142 XThC.Tn[13].n27 XThC.Tn[13].n25 161.406
R19143 XThC.Tn[13].n30 XThC.Tn[13].n28 161.406
R19144 XThC.Tn[13].n33 XThC.Tn[13].n31 161.406
R19145 XThC.Tn[13].n36 XThC.Tn[13].n34 161.406
R19146 XThC.Tn[13].n39 XThC.Tn[13].n37 161.406
R19147 XThC.Tn[13].n42 XThC.Tn[13].n40 161.406
R19148 XThC.Tn[13].n45 XThC.Tn[13].n43 161.406
R19149 XThC.Tn[13].n48 XThC.Tn[13].n46 161.406
R19150 XThC.Tn[13].n51 XThC.Tn[13].n49 161.406
R19151 XThC.Tn[13].n54 XThC.Tn[13].n52 161.406
R19152 XThC.Tn[13].n7 XThC.Tn[13].t27 161.202
R19153 XThC.Tn[13].n10 XThC.Tn[13].t12 161.202
R19154 XThC.Tn[13].n13 XThC.Tn[13].t14 161.202
R19155 XThC.Tn[13].n16 XThC.Tn[13].t16 161.202
R19156 XThC.Tn[13].n19 XThC.Tn[13].t37 161.202
R19157 XThC.Tn[13].n22 XThC.Tn[13].t38 161.202
R19158 XThC.Tn[13].n25 XThC.Tn[13].t19 161.202
R19159 XThC.Tn[13].n28 XThC.Tn[13].t28 161.202
R19160 XThC.Tn[13].n31 XThC.Tn[13].t30 161.202
R19161 XThC.Tn[13].n34 XThC.Tn[13].t17 161.202
R19162 XThC.Tn[13].n37 XThC.Tn[13].t18 161.202
R19163 XThC.Tn[13].n40 XThC.Tn[13].t31 161.202
R19164 XThC.Tn[13].n43 XThC.Tn[13].t39 161.202
R19165 XThC.Tn[13].n46 XThC.Tn[13].t42 161.202
R19166 XThC.Tn[13].n49 XThC.Tn[13].t23 161.202
R19167 XThC.Tn[13].n52 XThC.Tn[13].t33 161.202
R19168 XThC.Tn[13].n7 XThC.Tn[13].t29 145.137
R19169 XThC.Tn[13].n10 XThC.Tn[13].t15 145.137
R19170 XThC.Tn[13].n13 XThC.Tn[13].t20 145.137
R19171 XThC.Tn[13].n16 XThC.Tn[13].t21 145.137
R19172 XThC.Tn[13].n19 XThC.Tn[13].t40 145.137
R19173 XThC.Tn[13].n22 XThC.Tn[13].t41 145.137
R19174 XThC.Tn[13].n25 XThC.Tn[13].t25 145.137
R19175 XThC.Tn[13].n28 XThC.Tn[13].t32 145.137
R19176 XThC.Tn[13].n31 XThC.Tn[13].t34 145.137
R19177 XThC.Tn[13].n34 XThC.Tn[13].t22 145.137
R19178 XThC.Tn[13].n37 XThC.Tn[13].t24 145.137
R19179 XThC.Tn[13].n40 XThC.Tn[13].t35 145.137
R19180 XThC.Tn[13].n43 XThC.Tn[13].t43 145.137
R19181 XThC.Tn[13].n46 XThC.Tn[13].t13 145.137
R19182 XThC.Tn[13].n49 XThC.Tn[13].t26 145.137
R19183 XThC.Tn[13].n52 XThC.Tn[13].t36 145.137
R19184 XThC.Tn[13].n1 XThC.Tn[13].t4 26.5955
R19185 XThC.Tn[13].n1 XThC.Tn[13].t7 26.5955
R19186 XThC.Tn[13].n0 XThC.Tn[13].t6 26.5955
R19187 XThC.Tn[13].n0 XThC.Tn[13].t5 26.5955
R19188 XThC.Tn[13].n3 XThC.Tn[13].t9 26.5955
R19189 XThC.Tn[13].n3 XThC.Tn[13].t8 26.5955
R19190 XThC.Tn[13].n4 XThC.Tn[13].t11 26.5955
R19191 XThC.Tn[13].n4 XThC.Tn[13].t10 26.5955
R19192 XThC.Tn[13].n57 XThC.Tn[13].t0 24.9236
R19193 XThC.Tn[13].n57 XThC.Tn[13].t2 24.9236
R19194 XThC.Tn[13].n58 XThC.Tn[13].t3 24.9236
R19195 XThC.Tn[13].n58 XThC.Tn[13].t1 24.9236
R19196 XThC.Tn[13] XThC.Tn[13].n5 22.9652
R19197 XThC.Tn[13] XThC.Tn[13].n59 18.8943
R19198 XThC.Tn[13].n6 XThC.Tn[13].n2 13.9299
R19199 XThC.Tn[13].n6 XThC.Tn[13] 13.9299
R19200 XThC.Tn[13] XThC.Tn[13].n56 6.34069
R19201 XThC.Tn[13].n56 XThC.Tn[13].n55 5.13021
R19202 XThC.Tn[13].n55 XThC.Tn[13] 4.03795
R19203 XThC.Tn[13].n56 XThC.Tn[13] 1.79489
R19204 XThC.Tn[13] XThC.Tn[13].n6 1.19676
R19205 XThC.Tn[13].n12 XThC.Tn[13] 0.931056
R19206 XThC.Tn[13].n15 XThC.Tn[13] 0.931056
R19207 XThC.Tn[13].n18 XThC.Tn[13] 0.931056
R19208 XThC.Tn[13].n21 XThC.Tn[13] 0.931056
R19209 XThC.Tn[13].n24 XThC.Tn[13] 0.931056
R19210 XThC.Tn[13].n27 XThC.Tn[13] 0.931056
R19211 XThC.Tn[13].n30 XThC.Tn[13] 0.931056
R19212 XThC.Tn[13].n33 XThC.Tn[13] 0.931056
R19213 XThC.Tn[13].n36 XThC.Tn[13] 0.931056
R19214 XThC.Tn[13].n39 XThC.Tn[13] 0.931056
R19215 XThC.Tn[13].n42 XThC.Tn[13] 0.931056
R19216 XThC.Tn[13].n45 XThC.Tn[13] 0.931056
R19217 XThC.Tn[13].n48 XThC.Tn[13] 0.931056
R19218 XThC.Tn[13].n51 XThC.Tn[13] 0.931056
R19219 XThC.Tn[13].n54 XThC.Tn[13] 0.931056
R19220 XThC.Tn[13] XThC.Tn[13].n9 0.396333
R19221 XThC.Tn[13] XThC.Tn[13].n12 0.396333
R19222 XThC.Tn[13] XThC.Tn[13].n15 0.396333
R19223 XThC.Tn[13] XThC.Tn[13].n18 0.396333
R19224 XThC.Tn[13] XThC.Tn[13].n21 0.396333
R19225 XThC.Tn[13] XThC.Tn[13].n24 0.396333
R19226 XThC.Tn[13] XThC.Tn[13].n27 0.396333
R19227 XThC.Tn[13] XThC.Tn[13].n30 0.396333
R19228 XThC.Tn[13] XThC.Tn[13].n33 0.396333
R19229 XThC.Tn[13] XThC.Tn[13].n36 0.396333
R19230 XThC.Tn[13] XThC.Tn[13].n39 0.396333
R19231 XThC.Tn[13] XThC.Tn[13].n42 0.396333
R19232 XThC.Tn[13] XThC.Tn[13].n45 0.396333
R19233 XThC.Tn[13] XThC.Tn[13].n48 0.396333
R19234 XThC.Tn[13] XThC.Tn[13].n51 0.396333
R19235 XThC.Tn[13] XThC.Tn[13].n54 0.396333
R19236 XThC.Tn[13].n8 XThC.Tn[13] 0.104667
R19237 XThC.Tn[13].n11 XThC.Tn[13] 0.104667
R19238 XThC.Tn[13].n14 XThC.Tn[13] 0.104667
R19239 XThC.Tn[13].n17 XThC.Tn[13] 0.104667
R19240 XThC.Tn[13].n20 XThC.Tn[13] 0.104667
R19241 XThC.Tn[13].n23 XThC.Tn[13] 0.104667
R19242 XThC.Tn[13].n26 XThC.Tn[13] 0.104667
R19243 XThC.Tn[13].n29 XThC.Tn[13] 0.104667
R19244 XThC.Tn[13].n32 XThC.Tn[13] 0.104667
R19245 XThC.Tn[13].n35 XThC.Tn[13] 0.104667
R19246 XThC.Tn[13].n38 XThC.Tn[13] 0.104667
R19247 XThC.Tn[13].n41 XThC.Tn[13] 0.104667
R19248 XThC.Tn[13].n44 XThC.Tn[13] 0.104667
R19249 XThC.Tn[13].n47 XThC.Tn[13] 0.104667
R19250 XThC.Tn[13].n50 XThC.Tn[13] 0.104667
R19251 XThC.Tn[13].n53 XThC.Tn[13] 0.104667
R19252 XThC.Tn[13].n8 XThC.Tn[13] 0.0309878
R19253 XThC.Tn[13].n11 XThC.Tn[13] 0.0309878
R19254 XThC.Tn[13].n14 XThC.Tn[13] 0.0309878
R19255 XThC.Tn[13].n17 XThC.Tn[13] 0.0309878
R19256 XThC.Tn[13].n20 XThC.Tn[13] 0.0309878
R19257 XThC.Tn[13].n23 XThC.Tn[13] 0.0309878
R19258 XThC.Tn[13].n26 XThC.Tn[13] 0.0309878
R19259 XThC.Tn[13].n29 XThC.Tn[13] 0.0309878
R19260 XThC.Tn[13].n32 XThC.Tn[13] 0.0309878
R19261 XThC.Tn[13].n35 XThC.Tn[13] 0.0309878
R19262 XThC.Tn[13].n38 XThC.Tn[13] 0.0309878
R19263 XThC.Tn[13].n41 XThC.Tn[13] 0.0309878
R19264 XThC.Tn[13].n44 XThC.Tn[13] 0.0309878
R19265 XThC.Tn[13].n47 XThC.Tn[13] 0.0309878
R19266 XThC.Tn[13].n50 XThC.Tn[13] 0.0309878
R19267 XThC.Tn[13].n53 XThC.Tn[13] 0.0309878
R19268 XThC.Tn[13].n9 XThC.Tn[13].n8 0.027939
R19269 XThC.Tn[13].n12 XThC.Tn[13].n11 0.027939
R19270 XThC.Tn[13].n15 XThC.Tn[13].n14 0.027939
R19271 XThC.Tn[13].n18 XThC.Tn[13].n17 0.027939
R19272 XThC.Tn[13].n21 XThC.Tn[13].n20 0.027939
R19273 XThC.Tn[13].n24 XThC.Tn[13].n23 0.027939
R19274 XThC.Tn[13].n27 XThC.Tn[13].n26 0.027939
R19275 XThC.Tn[13].n30 XThC.Tn[13].n29 0.027939
R19276 XThC.Tn[13].n33 XThC.Tn[13].n32 0.027939
R19277 XThC.Tn[13].n36 XThC.Tn[13].n35 0.027939
R19278 XThC.Tn[13].n39 XThC.Tn[13].n38 0.027939
R19279 XThC.Tn[13].n42 XThC.Tn[13].n41 0.027939
R19280 XThC.Tn[13].n45 XThC.Tn[13].n44 0.027939
R19281 XThC.Tn[13].n48 XThC.Tn[13].n47 0.027939
R19282 XThC.Tn[13].n51 XThC.Tn[13].n50 0.027939
R19283 XThC.Tn[13].n54 XThC.Tn[13].n53 0.027939
R19284 XThC.Tn[13].n55 XThC.Tn[13] 0.00548355
R19285 XThC.Tn[0].n59 XThC.Tn[0].n58 332.332
R19286 XThC.Tn[0].n59 XThC.Tn[0].n57 296.493
R19287 XThC.Tn[0].n9 XThC.Tn[0].n7 161.406
R19288 XThC.Tn[0].n12 XThC.Tn[0].n10 161.406
R19289 XThC.Tn[0].n15 XThC.Tn[0].n13 161.406
R19290 XThC.Tn[0].n18 XThC.Tn[0].n16 161.406
R19291 XThC.Tn[0].n21 XThC.Tn[0].n19 161.406
R19292 XThC.Tn[0].n24 XThC.Tn[0].n22 161.406
R19293 XThC.Tn[0].n27 XThC.Tn[0].n25 161.406
R19294 XThC.Tn[0].n30 XThC.Tn[0].n28 161.406
R19295 XThC.Tn[0].n33 XThC.Tn[0].n31 161.406
R19296 XThC.Tn[0].n36 XThC.Tn[0].n34 161.406
R19297 XThC.Tn[0].n39 XThC.Tn[0].n37 161.406
R19298 XThC.Tn[0].n42 XThC.Tn[0].n40 161.406
R19299 XThC.Tn[0].n45 XThC.Tn[0].n43 161.406
R19300 XThC.Tn[0].n48 XThC.Tn[0].n46 161.406
R19301 XThC.Tn[0].n51 XThC.Tn[0].n49 161.406
R19302 XThC.Tn[0].n54 XThC.Tn[0].n52 161.406
R19303 XThC.Tn[0].n7 XThC.Tn[0].t22 161.202
R19304 XThC.Tn[0].n10 XThC.Tn[0].t41 161.202
R19305 XThC.Tn[0].n13 XThC.Tn[0].t12 161.202
R19306 XThC.Tn[0].n16 XThC.Tn[0].t13 161.202
R19307 XThC.Tn[0].n19 XThC.Tn[0].t32 161.202
R19308 XThC.Tn[0].n22 XThC.Tn[0].t34 161.202
R19309 XThC.Tn[0].n25 XThC.Tn[0].t17 161.202
R19310 XThC.Tn[0].n28 XThC.Tn[0].t25 161.202
R19311 XThC.Tn[0].n31 XThC.Tn[0].t26 161.202
R19312 XThC.Tn[0].n34 XThC.Tn[0].t15 161.202
R19313 XThC.Tn[0].n37 XThC.Tn[0].t16 161.202
R19314 XThC.Tn[0].n40 XThC.Tn[0].t27 161.202
R19315 XThC.Tn[0].n43 XThC.Tn[0].t36 161.202
R19316 XThC.Tn[0].n46 XThC.Tn[0].t38 161.202
R19317 XThC.Tn[0].n49 XThC.Tn[0].t19 161.202
R19318 XThC.Tn[0].n52 XThC.Tn[0].t29 161.202
R19319 XThC.Tn[0].n7 XThC.Tn[0].t18 145.137
R19320 XThC.Tn[0].n10 XThC.Tn[0].t35 145.137
R19321 XThC.Tn[0].n13 XThC.Tn[0].t37 145.137
R19322 XThC.Tn[0].n16 XThC.Tn[0].t39 145.137
R19323 XThC.Tn[0].n19 XThC.Tn[0].t28 145.137
R19324 XThC.Tn[0].n22 XThC.Tn[0].t30 145.137
R19325 XThC.Tn[0].n25 XThC.Tn[0].t43 145.137
R19326 XThC.Tn[0].n28 XThC.Tn[0].t20 145.137
R19327 XThC.Tn[0].n31 XThC.Tn[0].t21 145.137
R19328 XThC.Tn[0].n34 XThC.Tn[0].t40 145.137
R19329 XThC.Tn[0].n37 XThC.Tn[0].t42 145.137
R19330 XThC.Tn[0].n40 XThC.Tn[0].t23 145.137
R19331 XThC.Tn[0].n43 XThC.Tn[0].t31 145.137
R19332 XThC.Tn[0].n46 XThC.Tn[0].t33 145.137
R19333 XThC.Tn[0].n49 XThC.Tn[0].t14 145.137
R19334 XThC.Tn[0].n52 XThC.Tn[0].t24 145.137
R19335 XThC.Tn[0].n2 XThC.Tn[0].n0 135.248
R19336 XThC.Tn[0].n2 XThC.Tn[0].n1 98.982
R19337 XThC.Tn[0].n4 XThC.Tn[0].n3 98.982
R19338 XThC.Tn[0].n6 XThC.Tn[0].n5 98.982
R19339 XThC.Tn[0].n4 XThC.Tn[0].n2 36.2672
R19340 XThC.Tn[0].n6 XThC.Tn[0].n4 36.2672
R19341 XThC.Tn[0].n56 XThC.Tn[0].n6 32.6405
R19342 XThC.Tn[0].n57 XThC.Tn[0].t1 26.5955
R19343 XThC.Tn[0].n57 XThC.Tn[0].t0 26.5955
R19344 XThC.Tn[0].n58 XThC.Tn[0].t3 26.5955
R19345 XThC.Tn[0].n58 XThC.Tn[0].t2 26.5955
R19346 XThC.Tn[0].n0 XThC.Tn[0].t8 24.9236
R19347 XThC.Tn[0].n0 XThC.Tn[0].t9 24.9236
R19348 XThC.Tn[0].n1 XThC.Tn[0].t10 24.9236
R19349 XThC.Tn[0].n1 XThC.Tn[0].t11 24.9236
R19350 XThC.Tn[0].n3 XThC.Tn[0].t7 24.9236
R19351 XThC.Tn[0].n3 XThC.Tn[0].t6 24.9236
R19352 XThC.Tn[0].n5 XThC.Tn[0].t5 24.9236
R19353 XThC.Tn[0].n5 XThC.Tn[0].t4 24.9236
R19354 XThC.Tn[0].n60 XThC.Tn[0].n59 18.5605
R19355 XThC.Tn[0].n60 XThC.Tn[0].n56 11.5205
R19356 XThC.Tn[0].n56 XThC.Tn[0].n55 3.16389
R19357 XThC.Tn[0].n12 XThC.Tn[0] 0.931056
R19358 XThC.Tn[0].n15 XThC.Tn[0] 0.931056
R19359 XThC.Tn[0].n18 XThC.Tn[0] 0.931056
R19360 XThC.Tn[0].n21 XThC.Tn[0] 0.931056
R19361 XThC.Tn[0].n24 XThC.Tn[0] 0.931056
R19362 XThC.Tn[0].n27 XThC.Tn[0] 0.931056
R19363 XThC.Tn[0].n30 XThC.Tn[0] 0.931056
R19364 XThC.Tn[0].n33 XThC.Tn[0] 0.931056
R19365 XThC.Tn[0].n36 XThC.Tn[0] 0.931056
R19366 XThC.Tn[0].n39 XThC.Tn[0] 0.931056
R19367 XThC.Tn[0].n42 XThC.Tn[0] 0.931056
R19368 XThC.Tn[0].n45 XThC.Tn[0] 0.931056
R19369 XThC.Tn[0].n48 XThC.Tn[0] 0.931056
R19370 XThC.Tn[0].n51 XThC.Tn[0] 0.931056
R19371 XThC.Tn[0].n54 XThC.Tn[0] 0.931056
R19372 XThC.Tn[0] XThC.Tn[0].n60 0.6405
R19373 XThC.Tn[0] XThC.Tn[0].n9 0.396333
R19374 XThC.Tn[0] XThC.Tn[0].n12 0.396333
R19375 XThC.Tn[0] XThC.Tn[0].n15 0.396333
R19376 XThC.Tn[0] XThC.Tn[0].n18 0.396333
R19377 XThC.Tn[0] XThC.Tn[0].n21 0.396333
R19378 XThC.Tn[0] XThC.Tn[0].n24 0.396333
R19379 XThC.Tn[0] XThC.Tn[0].n27 0.396333
R19380 XThC.Tn[0] XThC.Tn[0].n30 0.396333
R19381 XThC.Tn[0] XThC.Tn[0].n33 0.396333
R19382 XThC.Tn[0] XThC.Tn[0].n36 0.396333
R19383 XThC.Tn[0] XThC.Tn[0].n39 0.396333
R19384 XThC.Tn[0] XThC.Tn[0].n42 0.396333
R19385 XThC.Tn[0] XThC.Tn[0].n45 0.396333
R19386 XThC.Tn[0] XThC.Tn[0].n48 0.396333
R19387 XThC.Tn[0] XThC.Tn[0].n51 0.396333
R19388 XThC.Tn[0] XThC.Tn[0].n54 0.396333
R19389 XThC.Tn[0].n55 XThC.Tn[0] 0.243556
R19390 XThC.Tn[0].n8 XThC.Tn[0] 0.104667
R19391 XThC.Tn[0].n11 XThC.Tn[0] 0.104667
R19392 XThC.Tn[0].n14 XThC.Tn[0] 0.104667
R19393 XThC.Tn[0].n17 XThC.Tn[0] 0.104667
R19394 XThC.Tn[0].n20 XThC.Tn[0] 0.104667
R19395 XThC.Tn[0].n23 XThC.Tn[0] 0.104667
R19396 XThC.Tn[0].n26 XThC.Tn[0] 0.104667
R19397 XThC.Tn[0].n29 XThC.Tn[0] 0.104667
R19398 XThC.Tn[0].n32 XThC.Tn[0] 0.104667
R19399 XThC.Tn[0].n35 XThC.Tn[0] 0.104667
R19400 XThC.Tn[0].n38 XThC.Tn[0] 0.104667
R19401 XThC.Tn[0].n41 XThC.Tn[0] 0.104667
R19402 XThC.Tn[0].n44 XThC.Tn[0] 0.104667
R19403 XThC.Tn[0].n47 XThC.Tn[0] 0.104667
R19404 XThC.Tn[0].n50 XThC.Tn[0] 0.104667
R19405 XThC.Tn[0].n53 XThC.Tn[0] 0.104667
R19406 XThC.Tn[0].n55 XThC.Tn[0] 0.0326429
R19407 XThC.Tn[0].n8 XThC.Tn[0] 0.0309878
R19408 XThC.Tn[0].n11 XThC.Tn[0] 0.0309878
R19409 XThC.Tn[0].n14 XThC.Tn[0] 0.0309878
R19410 XThC.Tn[0].n17 XThC.Tn[0] 0.0309878
R19411 XThC.Tn[0].n20 XThC.Tn[0] 0.0309878
R19412 XThC.Tn[0].n23 XThC.Tn[0] 0.0309878
R19413 XThC.Tn[0].n26 XThC.Tn[0] 0.0309878
R19414 XThC.Tn[0].n29 XThC.Tn[0] 0.0309878
R19415 XThC.Tn[0].n32 XThC.Tn[0] 0.0309878
R19416 XThC.Tn[0].n35 XThC.Tn[0] 0.0309878
R19417 XThC.Tn[0].n38 XThC.Tn[0] 0.0309878
R19418 XThC.Tn[0].n41 XThC.Tn[0] 0.0309878
R19419 XThC.Tn[0].n44 XThC.Tn[0] 0.0309878
R19420 XThC.Tn[0].n47 XThC.Tn[0] 0.0309878
R19421 XThC.Tn[0].n50 XThC.Tn[0] 0.0309878
R19422 XThC.Tn[0].n53 XThC.Tn[0] 0.0309878
R19423 XThC.Tn[0].n9 XThC.Tn[0].n8 0.027939
R19424 XThC.Tn[0].n12 XThC.Tn[0].n11 0.027939
R19425 XThC.Tn[0].n15 XThC.Tn[0].n14 0.027939
R19426 XThC.Tn[0].n18 XThC.Tn[0].n17 0.027939
R19427 XThC.Tn[0].n21 XThC.Tn[0].n20 0.027939
R19428 XThC.Tn[0].n24 XThC.Tn[0].n23 0.027939
R19429 XThC.Tn[0].n27 XThC.Tn[0].n26 0.027939
R19430 XThC.Tn[0].n30 XThC.Tn[0].n29 0.027939
R19431 XThC.Tn[0].n33 XThC.Tn[0].n32 0.027939
R19432 XThC.Tn[0].n36 XThC.Tn[0].n35 0.027939
R19433 XThC.Tn[0].n39 XThC.Tn[0].n38 0.027939
R19434 XThC.Tn[0].n42 XThC.Tn[0].n41 0.027939
R19435 XThC.Tn[0].n45 XThC.Tn[0].n44 0.027939
R19436 XThC.Tn[0].n48 XThC.Tn[0].n47 0.027939
R19437 XThC.Tn[0].n51 XThC.Tn[0].n50 0.027939
R19438 XThC.Tn[0].n54 XThC.Tn[0].n53 0.027939
R19439 XThC.XTB4.Y.t0 XThC.XTB4.Y.n21 268.738
R19440 XThC.XTB4.Y.n22 XThC.XTB4.Y.t0 268.077
R19441 XThC.XTB4.Y.n0 XThC.XTB4.Y.t1 235.56
R19442 XThC.XTB4.Y.n4 XThC.XTB4.Y.t3 212.081
R19443 XThC.XTB4.Y.n3 XThC.XTB4.Y.t2 212.081
R19444 XThC.XTB4.Y.n9 XThC.XTB4.Y.t17 212.081
R19445 XThC.XTB4.Y.n1 XThC.XTB4.Y.t13 212.081
R19446 XThC.XTB4.Y.n13 XThC.XTB4.Y.t8 212.081
R19447 XThC.XTB4.Y.n14 XThC.XTB4.Y.t12 212.081
R19448 XThC.XTB4.Y.n16 XThC.XTB4.Y.t6 212.081
R19449 XThC.XTB4.Y.n12 XThC.XTB4.Y.t16 212.081
R19450 XThC.XTB4.Y.n6 XThC.XTB4.Y.n5 173.761
R19451 XThC.XTB4.Y.n15 XThC.XTB4.Y 158.656
R19452 XThC.XTB4.Y.n8 XThC.XTB4.Y.n7 152
R19453 XThC.XTB4.Y.n6 XThC.XTB4.Y.n2 152
R19454 XThC.XTB4.Y.n11 XThC.XTB4.Y.n10 152
R19455 XThC.XTB4.Y.n18 XThC.XTB4.Y.n17 152
R19456 XThC.XTB4.Y.n4 XThC.XTB4.Y.t14 139.78
R19457 XThC.XTB4.Y.n3 XThC.XTB4.Y.t10 139.78
R19458 XThC.XTB4.Y.n9 XThC.XTB4.Y.t7 139.78
R19459 XThC.XTB4.Y.n1 XThC.XTB4.Y.t4 139.78
R19460 XThC.XTB4.Y.n13 XThC.XTB4.Y.t11 139.78
R19461 XThC.XTB4.Y.n14 XThC.XTB4.Y.t15 139.78
R19462 XThC.XTB4.Y.n16 XThC.XTB4.Y.t9 139.78
R19463 XThC.XTB4.Y.n12 XThC.XTB4.Y.t5 139.78
R19464 XThC.XTB4.Y.n20 XThC.XTB4.Y.n11 72.9296
R19465 XThC.XTB4.Y.n14 XThC.XTB4.Y.n13 61.346
R19466 XThC.XTB4.Y.n8 XThC.XTB4.Y.n2 49.6611
R19467 XThC.XTB4.Y.n10 XThC.XTB4.Y.n9 45.2793
R19468 XThC.XTB4.Y.n5 XThC.XTB4.Y.n3 42.3581
R19469 XThC.XTB4.Y.n20 XThC.XTB4.Y.n19 38.1854
R19470 XThC.XTB4.Y.n17 XThC.XTB4.Y.n12 30.6732
R19471 XThC.XTB4.Y.n17 XThC.XTB4.Y.n16 30.6732
R19472 XThC.XTB4.Y.n16 XThC.XTB4.Y.n15 30.6732
R19473 XThC.XTB4.Y.n15 XThC.XTB4.Y.n14 30.6732
R19474 XThC.XTB4.Y.n7 XThC.XTB4.Y.n6 21.7605
R19475 XThC.XTB4.Y.n5 XThC.XTB4.Y.n4 18.9884
R19476 XThC.XTB4.Y XThC.XTB4.Y.n22 17.8682
R19477 XThC.XTB4.Y.n10 XThC.XTB4.Y.n1 16.0672
R19478 XThC.XTB4.Y.n18 XThC.XTB4.Y 14.7905
R19479 XThC.XTB4.Y.n11 XThC.XTB4.Y 11.5205
R19480 XThC.XTB4.Y.n21 XThC.XTB4.Y.n20 10.353
R19481 XThC.XTB4.Y.n7 XThC.XTB4.Y 10.2405
R19482 XThC.XTB4.Y.n3 XThC.XTB4.Y.n2 7.30353
R19483 XThC.XTB4.Y.n19 XThC.XTB4.Y.n18 7.24578
R19484 XThC.XTB4.Y.n9 XThC.XTB4.Y.n8 4.38232
R19485 XThC.XTB4.Y.n22 XThC.XTB4.Y.n21 3.29747
R19486 XThC.XTB4.Y XThC.XTB4.Y.n0 2.22659
R19487 XThC.XTB4.Y.n0 XThC.XTB4.Y 1.55202
R19488 XThC.XTB4.Y.n19 XThC.XTB4.Y 0.966538
R19489 XThR.Tn[3].n2 XThR.Tn[3].n1 332.332
R19490 XThR.Tn[3].n2 XThR.Tn[3].n0 296.493
R19491 XThR.Tn[3] XThR.Tn[3].n82 161.363
R19492 XThR.Tn[3] XThR.Tn[3].n77 161.363
R19493 XThR.Tn[3] XThR.Tn[3].n72 161.363
R19494 XThR.Tn[3] XThR.Tn[3].n67 161.363
R19495 XThR.Tn[3] XThR.Tn[3].n62 161.363
R19496 XThR.Tn[3] XThR.Tn[3].n57 161.363
R19497 XThR.Tn[3] XThR.Tn[3].n52 161.363
R19498 XThR.Tn[3] XThR.Tn[3].n47 161.363
R19499 XThR.Tn[3] XThR.Tn[3].n42 161.363
R19500 XThR.Tn[3] XThR.Tn[3].n37 161.363
R19501 XThR.Tn[3] XThR.Tn[3].n32 161.363
R19502 XThR.Tn[3] XThR.Tn[3].n27 161.363
R19503 XThR.Tn[3] XThR.Tn[3].n22 161.363
R19504 XThR.Tn[3] XThR.Tn[3].n17 161.363
R19505 XThR.Tn[3] XThR.Tn[3].n12 161.363
R19506 XThR.Tn[3] XThR.Tn[3].n10 161.363
R19507 XThR.Tn[3].n84 XThR.Tn[3].n83 161.3
R19508 XThR.Tn[3].n79 XThR.Tn[3].n78 161.3
R19509 XThR.Tn[3].n74 XThR.Tn[3].n73 161.3
R19510 XThR.Tn[3].n69 XThR.Tn[3].n68 161.3
R19511 XThR.Tn[3].n64 XThR.Tn[3].n63 161.3
R19512 XThR.Tn[3].n59 XThR.Tn[3].n58 161.3
R19513 XThR.Tn[3].n54 XThR.Tn[3].n53 161.3
R19514 XThR.Tn[3].n49 XThR.Tn[3].n48 161.3
R19515 XThR.Tn[3].n44 XThR.Tn[3].n43 161.3
R19516 XThR.Tn[3].n39 XThR.Tn[3].n38 161.3
R19517 XThR.Tn[3].n34 XThR.Tn[3].n33 161.3
R19518 XThR.Tn[3].n29 XThR.Tn[3].n28 161.3
R19519 XThR.Tn[3].n24 XThR.Tn[3].n23 161.3
R19520 XThR.Tn[3].n19 XThR.Tn[3].n18 161.3
R19521 XThR.Tn[3].n14 XThR.Tn[3].n13 161.3
R19522 XThR.Tn[3].n82 XThR.Tn[3].t46 161.106
R19523 XThR.Tn[3].n77 XThR.Tn[3].t53 161.106
R19524 XThR.Tn[3].n72 XThR.Tn[3].t34 161.106
R19525 XThR.Tn[3].n67 XThR.Tn[3].t17 161.106
R19526 XThR.Tn[3].n62 XThR.Tn[3].t44 161.106
R19527 XThR.Tn[3].n57 XThR.Tn[3].t69 161.106
R19528 XThR.Tn[3].n52 XThR.Tn[3].t51 161.106
R19529 XThR.Tn[3].n47 XThR.Tn[3].t31 161.106
R19530 XThR.Tn[3].n42 XThR.Tn[3].t14 161.106
R19531 XThR.Tn[3].n37 XThR.Tn[3].t20 161.106
R19532 XThR.Tn[3].n32 XThR.Tn[3].t68 161.106
R19533 XThR.Tn[3].n27 XThR.Tn[3].t33 161.106
R19534 XThR.Tn[3].n22 XThR.Tn[3].t67 161.106
R19535 XThR.Tn[3].n17 XThR.Tn[3].t49 161.106
R19536 XThR.Tn[3].n12 XThR.Tn[3].t70 161.106
R19537 XThR.Tn[3].n10 XThR.Tn[3].t57 161.106
R19538 XThR.Tn[3].n83 XThR.Tn[3].t27 159.978
R19539 XThR.Tn[3].n78 XThR.Tn[3].t32 159.978
R19540 XThR.Tn[3].n73 XThR.Tn[3].t15 159.978
R19541 XThR.Tn[3].n68 XThR.Tn[3].t63 159.978
R19542 XThR.Tn[3].n63 XThR.Tn[3].t25 159.978
R19543 XThR.Tn[3].n58 XThR.Tn[3].t50 159.978
R19544 XThR.Tn[3].n53 XThR.Tn[3].t30 159.978
R19545 XThR.Tn[3].n48 XThR.Tn[3].t73 159.978
R19546 XThR.Tn[3].n43 XThR.Tn[3].t61 159.978
R19547 XThR.Tn[3].n38 XThR.Tn[3].t66 159.978
R19548 XThR.Tn[3].n33 XThR.Tn[3].t48 159.978
R19549 XThR.Tn[3].n28 XThR.Tn[3].t13 159.978
R19550 XThR.Tn[3].n23 XThR.Tn[3].t47 159.978
R19551 XThR.Tn[3].n18 XThR.Tn[3].t29 159.978
R19552 XThR.Tn[3].n13 XThR.Tn[3].t55 159.978
R19553 XThR.Tn[3].n82 XThR.Tn[3].t36 145.038
R19554 XThR.Tn[3].n77 XThR.Tn[3].t60 145.038
R19555 XThR.Tn[3].n72 XThR.Tn[3].t40 145.038
R19556 XThR.Tn[3].n67 XThR.Tn[3].t21 145.038
R19557 XThR.Tn[3].n62 XThR.Tn[3].t54 145.038
R19558 XThR.Tn[3].n57 XThR.Tn[3].t35 145.038
R19559 XThR.Tn[3].n52 XThR.Tn[3].t41 145.038
R19560 XThR.Tn[3].n47 XThR.Tn[3].t22 145.038
R19561 XThR.Tn[3].n42 XThR.Tn[3].t19 145.038
R19562 XThR.Tn[3].n37 XThR.Tn[3].t52 145.038
R19563 XThR.Tn[3].n32 XThR.Tn[3].t72 145.038
R19564 XThR.Tn[3].n27 XThR.Tn[3].t39 145.038
R19565 XThR.Tn[3].n22 XThR.Tn[3].t71 145.038
R19566 XThR.Tn[3].n17 XThR.Tn[3].t59 145.038
R19567 XThR.Tn[3].n12 XThR.Tn[3].t18 145.038
R19568 XThR.Tn[3].n10 XThR.Tn[3].t64 145.038
R19569 XThR.Tn[3].n83 XThR.Tn[3].t38 143.911
R19570 XThR.Tn[3].n78 XThR.Tn[3].t65 143.911
R19571 XThR.Tn[3].n73 XThR.Tn[3].t43 143.911
R19572 XThR.Tn[3].n68 XThR.Tn[3].t26 143.911
R19573 XThR.Tn[3].n63 XThR.Tn[3].t58 143.911
R19574 XThR.Tn[3].n58 XThR.Tn[3].t37 143.911
R19575 XThR.Tn[3].n53 XThR.Tn[3].t45 143.911
R19576 XThR.Tn[3].n48 XThR.Tn[3].t28 143.911
R19577 XThR.Tn[3].n43 XThR.Tn[3].t23 143.911
R19578 XThR.Tn[3].n38 XThR.Tn[3].t56 143.911
R19579 XThR.Tn[3].n33 XThR.Tn[3].t16 143.911
R19580 XThR.Tn[3].n28 XThR.Tn[3].t42 143.911
R19581 XThR.Tn[3].n23 XThR.Tn[3].t12 143.911
R19582 XThR.Tn[3].n18 XThR.Tn[3].t62 143.911
R19583 XThR.Tn[3].n13 XThR.Tn[3].t24 143.911
R19584 XThR.Tn[3].n7 XThR.Tn[3].n5 135.249
R19585 XThR.Tn[3].n9 XThR.Tn[3].n3 98.981
R19586 XThR.Tn[3].n8 XThR.Tn[3].n4 98.981
R19587 XThR.Tn[3].n7 XThR.Tn[3].n6 98.981
R19588 XThR.Tn[3].n9 XThR.Tn[3].n8 36.2672
R19589 XThR.Tn[3].n8 XThR.Tn[3].n7 36.2672
R19590 XThR.Tn[3].n88 XThR.Tn[3].n9 32.6405
R19591 XThR.Tn[3].n1 XThR.Tn[3].t4 26.5955
R19592 XThR.Tn[3].n1 XThR.Tn[3].t7 26.5955
R19593 XThR.Tn[3].n0 XThR.Tn[3].t5 26.5955
R19594 XThR.Tn[3].n0 XThR.Tn[3].t6 26.5955
R19595 XThR.Tn[3].n3 XThR.Tn[3].t11 24.9236
R19596 XThR.Tn[3].n3 XThR.Tn[3].t8 24.9236
R19597 XThR.Tn[3].n4 XThR.Tn[3].t10 24.9236
R19598 XThR.Tn[3].n4 XThR.Tn[3].t9 24.9236
R19599 XThR.Tn[3].n5 XThR.Tn[3].t0 24.9236
R19600 XThR.Tn[3].n5 XThR.Tn[3].t1 24.9236
R19601 XThR.Tn[3].n6 XThR.Tn[3].t3 24.9236
R19602 XThR.Tn[3].n6 XThR.Tn[3].t2 24.9236
R19603 XThR.Tn[3].n89 XThR.Tn[3].n2 18.5605
R19604 XThR.Tn[3].n89 XThR.Tn[3].n88 11.5205
R19605 XThR.Tn[3].n88 XThR.Tn[3] 6.21508
R19606 XThR.Tn[3] XThR.Tn[3].n11 5.34038
R19607 XThR.Tn[3].n16 XThR.Tn[3].n15 4.5005
R19608 XThR.Tn[3].n21 XThR.Tn[3].n20 4.5005
R19609 XThR.Tn[3].n26 XThR.Tn[3].n25 4.5005
R19610 XThR.Tn[3].n31 XThR.Tn[3].n30 4.5005
R19611 XThR.Tn[3].n36 XThR.Tn[3].n35 4.5005
R19612 XThR.Tn[3].n41 XThR.Tn[3].n40 4.5005
R19613 XThR.Tn[3].n46 XThR.Tn[3].n45 4.5005
R19614 XThR.Tn[3].n51 XThR.Tn[3].n50 4.5005
R19615 XThR.Tn[3].n56 XThR.Tn[3].n55 4.5005
R19616 XThR.Tn[3].n61 XThR.Tn[3].n60 4.5005
R19617 XThR.Tn[3].n66 XThR.Tn[3].n65 4.5005
R19618 XThR.Tn[3].n71 XThR.Tn[3].n70 4.5005
R19619 XThR.Tn[3].n76 XThR.Tn[3].n75 4.5005
R19620 XThR.Tn[3].n81 XThR.Tn[3].n80 4.5005
R19621 XThR.Tn[3].n86 XThR.Tn[3].n85 4.5005
R19622 XThR.Tn[3].n87 XThR.Tn[3] 3.70586
R19623 XThR.Tn[3].n16 XThR.Tn[3] 2.52282
R19624 XThR.Tn[3].n21 XThR.Tn[3] 2.52282
R19625 XThR.Tn[3].n26 XThR.Tn[3] 2.52282
R19626 XThR.Tn[3].n31 XThR.Tn[3] 2.52282
R19627 XThR.Tn[3].n36 XThR.Tn[3] 2.52282
R19628 XThR.Tn[3].n41 XThR.Tn[3] 2.52282
R19629 XThR.Tn[3].n46 XThR.Tn[3] 2.52282
R19630 XThR.Tn[3].n51 XThR.Tn[3] 2.52282
R19631 XThR.Tn[3].n56 XThR.Tn[3] 2.52282
R19632 XThR.Tn[3].n61 XThR.Tn[3] 2.52282
R19633 XThR.Tn[3].n66 XThR.Tn[3] 2.52282
R19634 XThR.Tn[3].n71 XThR.Tn[3] 2.52282
R19635 XThR.Tn[3].n76 XThR.Tn[3] 2.52282
R19636 XThR.Tn[3].n81 XThR.Tn[3] 2.52282
R19637 XThR.Tn[3].n86 XThR.Tn[3] 2.52282
R19638 XThR.Tn[3].n84 XThR.Tn[3] 1.08677
R19639 XThR.Tn[3].n79 XThR.Tn[3] 1.08677
R19640 XThR.Tn[3].n74 XThR.Tn[3] 1.08677
R19641 XThR.Tn[3].n69 XThR.Tn[3] 1.08677
R19642 XThR.Tn[3].n64 XThR.Tn[3] 1.08677
R19643 XThR.Tn[3].n59 XThR.Tn[3] 1.08677
R19644 XThR.Tn[3].n54 XThR.Tn[3] 1.08677
R19645 XThR.Tn[3].n49 XThR.Tn[3] 1.08677
R19646 XThR.Tn[3].n44 XThR.Tn[3] 1.08677
R19647 XThR.Tn[3].n39 XThR.Tn[3] 1.08677
R19648 XThR.Tn[3].n34 XThR.Tn[3] 1.08677
R19649 XThR.Tn[3].n29 XThR.Tn[3] 1.08677
R19650 XThR.Tn[3].n24 XThR.Tn[3] 1.08677
R19651 XThR.Tn[3].n19 XThR.Tn[3] 1.08677
R19652 XThR.Tn[3].n14 XThR.Tn[3] 1.08677
R19653 XThR.Tn[3] XThR.Tn[3].n16 0.839786
R19654 XThR.Tn[3] XThR.Tn[3].n21 0.839786
R19655 XThR.Tn[3] XThR.Tn[3].n26 0.839786
R19656 XThR.Tn[3] XThR.Tn[3].n31 0.839786
R19657 XThR.Tn[3] XThR.Tn[3].n36 0.839786
R19658 XThR.Tn[3] XThR.Tn[3].n41 0.839786
R19659 XThR.Tn[3] XThR.Tn[3].n46 0.839786
R19660 XThR.Tn[3] XThR.Tn[3].n51 0.839786
R19661 XThR.Tn[3] XThR.Tn[3].n56 0.839786
R19662 XThR.Tn[3] XThR.Tn[3].n61 0.839786
R19663 XThR.Tn[3] XThR.Tn[3].n66 0.839786
R19664 XThR.Tn[3] XThR.Tn[3].n71 0.839786
R19665 XThR.Tn[3] XThR.Tn[3].n76 0.839786
R19666 XThR.Tn[3] XThR.Tn[3].n81 0.839786
R19667 XThR.Tn[3] XThR.Tn[3].n86 0.839786
R19668 XThR.Tn[3] XThR.Tn[3].n89 0.6405
R19669 XThR.Tn[3].n11 XThR.Tn[3] 0.499542
R19670 XThR.Tn[3].n85 XThR.Tn[3] 0.063
R19671 XThR.Tn[3].n80 XThR.Tn[3] 0.063
R19672 XThR.Tn[3].n75 XThR.Tn[3] 0.063
R19673 XThR.Tn[3].n70 XThR.Tn[3] 0.063
R19674 XThR.Tn[3].n65 XThR.Tn[3] 0.063
R19675 XThR.Tn[3].n60 XThR.Tn[3] 0.063
R19676 XThR.Tn[3].n55 XThR.Tn[3] 0.063
R19677 XThR.Tn[3].n50 XThR.Tn[3] 0.063
R19678 XThR.Tn[3].n45 XThR.Tn[3] 0.063
R19679 XThR.Tn[3].n40 XThR.Tn[3] 0.063
R19680 XThR.Tn[3].n35 XThR.Tn[3] 0.063
R19681 XThR.Tn[3].n30 XThR.Tn[3] 0.063
R19682 XThR.Tn[3].n25 XThR.Tn[3] 0.063
R19683 XThR.Tn[3].n20 XThR.Tn[3] 0.063
R19684 XThR.Tn[3].n15 XThR.Tn[3] 0.063
R19685 XThR.Tn[3].n87 XThR.Tn[3] 0.0540714
R19686 XThR.Tn[3] XThR.Tn[3].n87 0.038
R19687 XThR.Tn[3].n11 XThR.Tn[3] 0.0143889
R19688 XThR.Tn[3].n85 XThR.Tn[3].n84 0.00771154
R19689 XThR.Tn[3].n80 XThR.Tn[3].n79 0.00771154
R19690 XThR.Tn[3].n75 XThR.Tn[3].n74 0.00771154
R19691 XThR.Tn[3].n70 XThR.Tn[3].n69 0.00771154
R19692 XThR.Tn[3].n65 XThR.Tn[3].n64 0.00771154
R19693 XThR.Tn[3].n60 XThR.Tn[3].n59 0.00771154
R19694 XThR.Tn[3].n55 XThR.Tn[3].n54 0.00771154
R19695 XThR.Tn[3].n50 XThR.Tn[3].n49 0.00771154
R19696 XThR.Tn[3].n45 XThR.Tn[3].n44 0.00771154
R19697 XThR.Tn[3].n40 XThR.Tn[3].n39 0.00771154
R19698 XThR.Tn[3].n35 XThR.Tn[3].n34 0.00771154
R19699 XThR.Tn[3].n30 XThR.Tn[3].n29 0.00771154
R19700 XThR.Tn[3].n25 XThR.Tn[3].n24 0.00771154
R19701 XThR.Tn[3].n20 XThR.Tn[3].n19 0.00771154
R19702 XThR.Tn[3].n15 XThR.Tn[3].n14 0.00771154
R19703 XThR.Tn[5].n2 XThR.Tn[5].n1 332.332
R19704 XThR.Tn[5].n2 XThR.Tn[5].n0 296.493
R19705 XThR.Tn[5] XThR.Tn[5].n82 161.363
R19706 XThR.Tn[5] XThR.Tn[5].n77 161.363
R19707 XThR.Tn[5] XThR.Tn[5].n72 161.363
R19708 XThR.Tn[5] XThR.Tn[5].n67 161.363
R19709 XThR.Tn[5] XThR.Tn[5].n62 161.363
R19710 XThR.Tn[5] XThR.Tn[5].n57 161.363
R19711 XThR.Tn[5] XThR.Tn[5].n52 161.363
R19712 XThR.Tn[5] XThR.Tn[5].n47 161.363
R19713 XThR.Tn[5] XThR.Tn[5].n42 161.363
R19714 XThR.Tn[5] XThR.Tn[5].n37 161.363
R19715 XThR.Tn[5] XThR.Tn[5].n32 161.363
R19716 XThR.Tn[5] XThR.Tn[5].n27 161.363
R19717 XThR.Tn[5] XThR.Tn[5].n22 161.363
R19718 XThR.Tn[5] XThR.Tn[5].n17 161.363
R19719 XThR.Tn[5] XThR.Tn[5].n12 161.363
R19720 XThR.Tn[5] XThR.Tn[5].n10 161.363
R19721 XThR.Tn[5].n84 XThR.Tn[5].n83 161.3
R19722 XThR.Tn[5].n79 XThR.Tn[5].n78 161.3
R19723 XThR.Tn[5].n74 XThR.Tn[5].n73 161.3
R19724 XThR.Tn[5].n69 XThR.Tn[5].n68 161.3
R19725 XThR.Tn[5].n64 XThR.Tn[5].n63 161.3
R19726 XThR.Tn[5].n59 XThR.Tn[5].n58 161.3
R19727 XThR.Tn[5].n54 XThR.Tn[5].n53 161.3
R19728 XThR.Tn[5].n49 XThR.Tn[5].n48 161.3
R19729 XThR.Tn[5].n44 XThR.Tn[5].n43 161.3
R19730 XThR.Tn[5].n39 XThR.Tn[5].n38 161.3
R19731 XThR.Tn[5].n34 XThR.Tn[5].n33 161.3
R19732 XThR.Tn[5].n29 XThR.Tn[5].n28 161.3
R19733 XThR.Tn[5].n24 XThR.Tn[5].n23 161.3
R19734 XThR.Tn[5].n19 XThR.Tn[5].n18 161.3
R19735 XThR.Tn[5].n14 XThR.Tn[5].n13 161.3
R19736 XThR.Tn[5].n82 XThR.Tn[5].t62 161.106
R19737 XThR.Tn[5].n77 XThR.Tn[5].t70 161.106
R19738 XThR.Tn[5].n72 XThR.Tn[5].t52 161.106
R19739 XThR.Tn[5].n67 XThR.Tn[5].t35 161.106
R19740 XThR.Tn[5].n62 XThR.Tn[5].t60 161.106
R19741 XThR.Tn[5].n57 XThR.Tn[5].t24 161.106
R19742 XThR.Tn[5].n52 XThR.Tn[5].t68 161.106
R19743 XThR.Tn[5].n47 XThR.Tn[5].t49 161.106
R19744 XThR.Tn[5].n42 XThR.Tn[5].t32 161.106
R19745 XThR.Tn[5].n37 XThR.Tn[5].t40 161.106
R19746 XThR.Tn[5].n32 XThR.Tn[5].t22 161.106
R19747 XThR.Tn[5].n27 XThR.Tn[5].t51 161.106
R19748 XThR.Tn[5].n22 XThR.Tn[5].t21 161.106
R19749 XThR.Tn[5].n17 XThR.Tn[5].t66 161.106
R19750 XThR.Tn[5].n12 XThR.Tn[5].t26 161.106
R19751 XThR.Tn[5].n10 XThR.Tn[5].t72 161.106
R19752 XThR.Tn[5].n83 XThR.Tn[5].t59 159.978
R19753 XThR.Tn[5].n78 XThR.Tn[5].t64 159.978
R19754 XThR.Tn[5].n73 XThR.Tn[5].t47 159.978
R19755 XThR.Tn[5].n68 XThR.Tn[5].t31 159.978
R19756 XThR.Tn[5].n63 XThR.Tn[5].t57 159.978
R19757 XThR.Tn[5].n58 XThR.Tn[5].t20 159.978
R19758 XThR.Tn[5].n53 XThR.Tn[5].t63 159.978
R19759 XThR.Tn[5].n48 XThR.Tn[5].t45 159.978
R19760 XThR.Tn[5].n43 XThR.Tn[5].t29 159.978
R19761 XThR.Tn[5].n38 XThR.Tn[5].t37 159.978
R19762 XThR.Tn[5].n33 XThR.Tn[5].t19 159.978
R19763 XThR.Tn[5].n28 XThR.Tn[5].t46 159.978
R19764 XThR.Tn[5].n23 XThR.Tn[5].t18 159.978
R19765 XThR.Tn[5].n18 XThR.Tn[5].t61 159.978
R19766 XThR.Tn[5].n13 XThR.Tn[5].t23 159.978
R19767 XThR.Tn[5].n82 XThR.Tn[5].t54 145.038
R19768 XThR.Tn[5].n77 XThR.Tn[5].t12 145.038
R19769 XThR.Tn[5].n72 XThR.Tn[5].t56 145.038
R19770 XThR.Tn[5].n67 XThR.Tn[5].t41 145.038
R19771 XThR.Tn[5].n62 XThR.Tn[5].t71 145.038
R19772 XThR.Tn[5].n57 XThR.Tn[5].t53 145.038
R19773 XThR.Tn[5].n52 XThR.Tn[5].t58 145.038
R19774 XThR.Tn[5].n47 XThR.Tn[5].t42 145.038
R19775 XThR.Tn[5].n42 XThR.Tn[5].t38 145.038
R19776 XThR.Tn[5].n37 XThR.Tn[5].t69 145.038
R19777 XThR.Tn[5].n32 XThR.Tn[5].t30 145.038
R19778 XThR.Tn[5].n27 XThR.Tn[5].t55 145.038
R19779 XThR.Tn[5].n22 XThR.Tn[5].t28 145.038
R19780 XThR.Tn[5].n17 XThR.Tn[5].t73 145.038
R19781 XThR.Tn[5].n12 XThR.Tn[5].t39 145.038
R19782 XThR.Tn[5].n10 XThR.Tn[5].t17 145.038
R19783 XThR.Tn[5].n83 XThR.Tn[5].t27 143.911
R19784 XThR.Tn[5].n78 XThR.Tn[5].t50 143.911
R19785 XThR.Tn[5].n73 XThR.Tn[5].t34 143.911
R19786 XThR.Tn[5].n68 XThR.Tn[5].t15 143.911
R19787 XThR.Tn[5].n63 XThR.Tn[5].t44 143.911
R19788 XThR.Tn[5].n58 XThR.Tn[5].t25 143.911
R19789 XThR.Tn[5].n53 XThR.Tn[5].t36 143.911
R19790 XThR.Tn[5].n48 XThR.Tn[5].t16 143.911
R19791 XThR.Tn[5].n43 XThR.Tn[5].t14 143.911
R19792 XThR.Tn[5].n38 XThR.Tn[5].t43 143.911
R19793 XThR.Tn[5].n33 XThR.Tn[5].t67 143.911
R19794 XThR.Tn[5].n28 XThR.Tn[5].t33 143.911
R19795 XThR.Tn[5].n23 XThR.Tn[5].t65 143.911
R19796 XThR.Tn[5].n18 XThR.Tn[5].t48 143.911
R19797 XThR.Tn[5].n13 XThR.Tn[5].t13 143.911
R19798 XThR.Tn[5].n7 XThR.Tn[5].n5 135.249
R19799 XThR.Tn[5].n9 XThR.Tn[5].n3 98.981
R19800 XThR.Tn[5].n8 XThR.Tn[5].n4 98.981
R19801 XThR.Tn[5].n7 XThR.Tn[5].n6 98.981
R19802 XThR.Tn[5].n9 XThR.Tn[5].n8 36.2672
R19803 XThR.Tn[5].n8 XThR.Tn[5].n7 36.2672
R19804 XThR.Tn[5].n88 XThR.Tn[5].n9 32.6405
R19805 XThR.Tn[5].n1 XThR.Tn[5].t9 26.5955
R19806 XThR.Tn[5].n1 XThR.Tn[5].t8 26.5955
R19807 XThR.Tn[5].n0 XThR.Tn[5].t10 26.5955
R19808 XThR.Tn[5].n0 XThR.Tn[5].t11 26.5955
R19809 XThR.Tn[5].n3 XThR.Tn[5].t7 24.9236
R19810 XThR.Tn[5].n3 XThR.Tn[5].t4 24.9236
R19811 XThR.Tn[5].n4 XThR.Tn[5].t6 24.9236
R19812 XThR.Tn[5].n4 XThR.Tn[5].t5 24.9236
R19813 XThR.Tn[5].n5 XThR.Tn[5].t0 24.9236
R19814 XThR.Tn[5].n5 XThR.Tn[5].t1 24.9236
R19815 XThR.Tn[5].n6 XThR.Tn[5].t3 24.9236
R19816 XThR.Tn[5].n6 XThR.Tn[5].t2 24.9236
R19817 XThR.Tn[5].n89 XThR.Tn[5].n2 18.5605
R19818 XThR.Tn[5].n89 XThR.Tn[5].n88 11.5205
R19819 XThR.Tn[5].n88 XThR.Tn[5] 5.71508
R19820 XThR.Tn[5] XThR.Tn[5].n11 5.34038
R19821 XThR.Tn[5].n16 XThR.Tn[5].n15 4.5005
R19822 XThR.Tn[5].n21 XThR.Tn[5].n20 4.5005
R19823 XThR.Tn[5].n26 XThR.Tn[5].n25 4.5005
R19824 XThR.Tn[5].n31 XThR.Tn[5].n30 4.5005
R19825 XThR.Tn[5].n36 XThR.Tn[5].n35 4.5005
R19826 XThR.Tn[5].n41 XThR.Tn[5].n40 4.5005
R19827 XThR.Tn[5].n46 XThR.Tn[5].n45 4.5005
R19828 XThR.Tn[5].n51 XThR.Tn[5].n50 4.5005
R19829 XThR.Tn[5].n56 XThR.Tn[5].n55 4.5005
R19830 XThR.Tn[5].n61 XThR.Tn[5].n60 4.5005
R19831 XThR.Tn[5].n66 XThR.Tn[5].n65 4.5005
R19832 XThR.Tn[5].n71 XThR.Tn[5].n70 4.5005
R19833 XThR.Tn[5].n76 XThR.Tn[5].n75 4.5005
R19834 XThR.Tn[5].n81 XThR.Tn[5].n80 4.5005
R19835 XThR.Tn[5].n86 XThR.Tn[5].n85 4.5005
R19836 XThR.Tn[5].n87 XThR.Tn[5] 3.70586
R19837 XThR.Tn[5].n16 XThR.Tn[5] 2.52282
R19838 XThR.Tn[5].n21 XThR.Tn[5] 2.52282
R19839 XThR.Tn[5].n26 XThR.Tn[5] 2.52282
R19840 XThR.Tn[5].n31 XThR.Tn[5] 2.52282
R19841 XThR.Tn[5].n36 XThR.Tn[5] 2.52282
R19842 XThR.Tn[5].n41 XThR.Tn[5] 2.52282
R19843 XThR.Tn[5].n46 XThR.Tn[5] 2.52282
R19844 XThR.Tn[5].n51 XThR.Tn[5] 2.52282
R19845 XThR.Tn[5].n56 XThR.Tn[5] 2.52282
R19846 XThR.Tn[5].n61 XThR.Tn[5] 2.52282
R19847 XThR.Tn[5].n66 XThR.Tn[5] 2.52282
R19848 XThR.Tn[5].n71 XThR.Tn[5] 2.52282
R19849 XThR.Tn[5].n76 XThR.Tn[5] 2.52282
R19850 XThR.Tn[5].n81 XThR.Tn[5] 2.52282
R19851 XThR.Tn[5].n86 XThR.Tn[5] 2.52282
R19852 XThR.Tn[5].n84 XThR.Tn[5] 1.08677
R19853 XThR.Tn[5].n79 XThR.Tn[5] 1.08677
R19854 XThR.Tn[5].n74 XThR.Tn[5] 1.08677
R19855 XThR.Tn[5].n69 XThR.Tn[5] 1.08677
R19856 XThR.Tn[5].n64 XThR.Tn[5] 1.08677
R19857 XThR.Tn[5].n59 XThR.Tn[5] 1.08677
R19858 XThR.Tn[5].n54 XThR.Tn[5] 1.08677
R19859 XThR.Tn[5].n49 XThR.Tn[5] 1.08677
R19860 XThR.Tn[5].n44 XThR.Tn[5] 1.08677
R19861 XThR.Tn[5].n39 XThR.Tn[5] 1.08677
R19862 XThR.Tn[5].n34 XThR.Tn[5] 1.08677
R19863 XThR.Tn[5].n29 XThR.Tn[5] 1.08677
R19864 XThR.Tn[5].n24 XThR.Tn[5] 1.08677
R19865 XThR.Tn[5].n19 XThR.Tn[5] 1.08677
R19866 XThR.Tn[5].n14 XThR.Tn[5] 1.08677
R19867 XThR.Tn[5] XThR.Tn[5].n16 0.839786
R19868 XThR.Tn[5] XThR.Tn[5].n21 0.839786
R19869 XThR.Tn[5] XThR.Tn[5].n26 0.839786
R19870 XThR.Tn[5] XThR.Tn[5].n31 0.839786
R19871 XThR.Tn[5] XThR.Tn[5].n36 0.839786
R19872 XThR.Tn[5] XThR.Tn[5].n41 0.839786
R19873 XThR.Tn[5] XThR.Tn[5].n46 0.839786
R19874 XThR.Tn[5] XThR.Tn[5].n51 0.839786
R19875 XThR.Tn[5] XThR.Tn[5].n56 0.839786
R19876 XThR.Tn[5] XThR.Tn[5].n61 0.839786
R19877 XThR.Tn[5] XThR.Tn[5].n66 0.839786
R19878 XThR.Tn[5] XThR.Tn[5].n71 0.839786
R19879 XThR.Tn[5] XThR.Tn[5].n76 0.839786
R19880 XThR.Tn[5] XThR.Tn[5].n81 0.839786
R19881 XThR.Tn[5] XThR.Tn[5].n86 0.839786
R19882 XThR.Tn[5] XThR.Tn[5].n89 0.6405
R19883 XThR.Tn[5].n11 XThR.Tn[5] 0.499542
R19884 XThR.Tn[5].n85 XThR.Tn[5] 0.063
R19885 XThR.Tn[5].n80 XThR.Tn[5] 0.063
R19886 XThR.Tn[5].n75 XThR.Tn[5] 0.063
R19887 XThR.Tn[5].n70 XThR.Tn[5] 0.063
R19888 XThR.Tn[5].n65 XThR.Tn[5] 0.063
R19889 XThR.Tn[5].n60 XThR.Tn[5] 0.063
R19890 XThR.Tn[5].n55 XThR.Tn[5] 0.063
R19891 XThR.Tn[5].n50 XThR.Tn[5] 0.063
R19892 XThR.Tn[5].n45 XThR.Tn[5] 0.063
R19893 XThR.Tn[5].n40 XThR.Tn[5] 0.063
R19894 XThR.Tn[5].n35 XThR.Tn[5] 0.063
R19895 XThR.Tn[5].n30 XThR.Tn[5] 0.063
R19896 XThR.Tn[5].n25 XThR.Tn[5] 0.063
R19897 XThR.Tn[5].n20 XThR.Tn[5] 0.063
R19898 XThR.Tn[5].n15 XThR.Tn[5] 0.063
R19899 XThR.Tn[5].n87 XThR.Tn[5] 0.0540714
R19900 XThR.Tn[5] XThR.Tn[5].n87 0.038
R19901 XThR.Tn[5].n11 XThR.Tn[5] 0.0143889
R19902 XThR.Tn[5].n85 XThR.Tn[5].n84 0.00771154
R19903 XThR.Tn[5].n80 XThR.Tn[5].n79 0.00771154
R19904 XThR.Tn[5].n75 XThR.Tn[5].n74 0.00771154
R19905 XThR.Tn[5].n70 XThR.Tn[5].n69 0.00771154
R19906 XThR.Tn[5].n65 XThR.Tn[5].n64 0.00771154
R19907 XThR.Tn[5].n60 XThR.Tn[5].n59 0.00771154
R19908 XThR.Tn[5].n55 XThR.Tn[5].n54 0.00771154
R19909 XThR.Tn[5].n50 XThR.Tn[5].n49 0.00771154
R19910 XThR.Tn[5].n45 XThR.Tn[5].n44 0.00771154
R19911 XThR.Tn[5].n40 XThR.Tn[5].n39 0.00771154
R19912 XThR.Tn[5].n35 XThR.Tn[5].n34 0.00771154
R19913 XThR.Tn[5].n30 XThR.Tn[5].n29 0.00771154
R19914 XThR.Tn[5].n25 XThR.Tn[5].n24 0.00771154
R19915 XThR.Tn[5].n20 XThR.Tn[5].n19 0.00771154
R19916 XThR.Tn[5].n15 XThR.Tn[5].n14 0.00771154
R19917 XThC.Tn[4].n2 XThC.Tn[4].n1 332.332
R19918 XThC.Tn[4].n2 XThC.Tn[4].n0 296.493
R19919 XThC.Tn[4].n12 XThC.Tn[4].n10 161.406
R19920 XThC.Tn[4].n15 XThC.Tn[4].n13 161.406
R19921 XThC.Tn[4].n18 XThC.Tn[4].n16 161.406
R19922 XThC.Tn[4].n21 XThC.Tn[4].n19 161.406
R19923 XThC.Tn[4].n24 XThC.Tn[4].n22 161.406
R19924 XThC.Tn[4].n27 XThC.Tn[4].n25 161.406
R19925 XThC.Tn[4].n30 XThC.Tn[4].n28 161.406
R19926 XThC.Tn[4].n33 XThC.Tn[4].n31 161.406
R19927 XThC.Tn[4].n36 XThC.Tn[4].n34 161.406
R19928 XThC.Tn[4].n39 XThC.Tn[4].n37 161.406
R19929 XThC.Tn[4].n42 XThC.Tn[4].n40 161.406
R19930 XThC.Tn[4].n45 XThC.Tn[4].n43 161.406
R19931 XThC.Tn[4].n48 XThC.Tn[4].n46 161.406
R19932 XThC.Tn[4].n51 XThC.Tn[4].n49 161.406
R19933 XThC.Tn[4].n54 XThC.Tn[4].n52 161.406
R19934 XThC.Tn[4].n57 XThC.Tn[4].n55 161.406
R19935 XThC.Tn[4].n10 XThC.Tn[4].t26 161.202
R19936 XThC.Tn[4].n13 XThC.Tn[4].t43 161.202
R19937 XThC.Tn[4].n16 XThC.Tn[4].t13 161.202
R19938 XThC.Tn[4].n19 XThC.Tn[4].t15 161.202
R19939 XThC.Tn[4].n22 XThC.Tn[4].t36 161.202
R19940 XThC.Tn[4].n25 XThC.Tn[4].t37 161.202
R19941 XThC.Tn[4].n28 XThC.Tn[4].t18 161.202
R19942 XThC.Tn[4].n31 XThC.Tn[4].t27 161.202
R19943 XThC.Tn[4].n34 XThC.Tn[4].t29 161.202
R19944 XThC.Tn[4].n37 XThC.Tn[4].t16 161.202
R19945 XThC.Tn[4].n40 XThC.Tn[4].t17 161.202
R19946 XThC.Tn[4].n43 XThC.Tn[4].t30 161.202
R19947 XThC.Tn[4].n46 XThC.Tn[4].t38 161.202
R19948 XThC.Tn[4].n49 XThC.Tn[4].t41 161.202
R19949 XThC.Tn[4].n52 XThC.Tn[4].t22 161.202
R19950 XThC.Tn[4].n55 XThC.Tn[4].t32 161.202
R19951 XThC.Tn[4].n10 XThC.Tn[4].t28 145.137
R19952 XThC.Tn[4].n13 XThC.Tn[4].t14 145.137
R19953 XThC.Tn[4].n16 XThC.Tn[4].t19 145.137
R19954 XThC.Tn[4].n19 XThC.Tn[4].t20 145.137
R19955 XThC.Tn[4].n22 XThC.Tn[4].t39 145.137
R19956 XThC.Tn[4].n25 XThC.Tn[4].t40 145.137
R19957 XThC.Tn[4].n28 XThC.Tn[4].t24 145.137
R19958 XThC.Tn[4].n31 XThC.Tn[4].t31 145.137
R19959 XThC.Tn[4].n34 XThC.Tn[4].t33 145.137
R19960 XThC.Tn[4].n37 XThC.Tn[4].t21 145.137
R19961 XThC.Tn[4].n40 XThC.Tn[4].t23 145.137
R19962 XThC.Tn[4].n43 XThC.Tn[4].t34 145.137
R19963 XThC.Tn[4].n46 XThC.Tn[4].t42 145.137
R19964 XThC.Tn[4].n49 XThC.Tn[4].t12 145.137
R19965 XThC.Tn[4].n52 XThC.Tn[4].t25 145.137
R19966 XThC.Tn[4].n55 XThC.Tn[4].t35 145.137
R19967 XThC.Tn[4].n7 XThC.Tn[4].n6 135.248
R19968 XThC.Tn[4].n9 XThC.Tn[4].n3 98.982
R19969 XThC.Tn[4].n8 XThC.Tn[4].n4 98.982
R19970 XThC.Tn[4].n7 XThC.Tn[4].n5 98.982
R19971 XThC.Tn[4].n9 XThC.Tn[4].n8 36.2672
R19972 XThC.Tn[4].n8 XThC.Tn[4].n7 36.2672
R19973 XThC.Tn[4].n59 XThC.Tn[4].n9 32.6405
R19974 XThC.Tn[4].n1 XThC.Tn[4].t7 26.5955
R19975 XThC.Tn[4].n1 XThC.Tn[4].t6 26.5955
R19976 XThC.Tn[4].n0 XThC.Tn[4].t5 26.5955
R19977 XThC.Tn[4].n0 XThC.Tn[4].t4 26.5955
R19978 XThC.Tn[4].n3 XThC.Tn[4].t9 24.9236
R19979 XThC.Tn[4].n3 XThC.Tn[4].t8 24.9236
R19980 XThC.Tn[4].n4 XThC.Tn[4].t11 24.9236
R19981 XThC.Tn[4].n4 XThC.Tn[4].t10 24.9236
R19982 XThC.Tn[4].n5 XThC.Tn[4].t2 24.9236
R19983 XThC.Tn[4].n5 XThC.Tn[4].t1 24.9236
R19984 XThC.Tn[4].n6 XThC.Tn[4].t0 24.9236
R19985 XThC.Tn[4].n6 XThC.Tn[4].t3 24.9236
R19986 XThC.Tn[4].n60 XThC.Tn[4].n2 18.5605
R19987 XThC.Tn[4].n60 XThC.Tn[4].n59 11.5205
R19988 XThC.Tn[4].n58 XThC.Tn[4] 4.63701
R19989 XThC.Tn[4].n59 XThC.Tn[4].n58 3.1844
R19990 XThC.Tn[4].n15 XThC.Tn[4] 0.931056
R19991 XThC.Tn[4].n18 XThC.Tn[4] 0.931056
R19992 XThC.Tn[4].n21 XThC.Tn[4] 0.931056
R19993 XThC.Tn[4].n24 XThC.Tn[4] 0.931056
R19994 XThC.Tn[4].n27 XThC.Tn[4] 0.931056
R19995 XThC.Tn[4].n30 XThC.Tn[4] 0.931056
R19996 XThC.Tn[4].n33 XThC.Tn[4] 0.931056
R19997 XThC.Tn[4].n36 XThC.Tn[4] 0.931056
R19998 XThC.Tn[4].n39 XThC.Tn[4] 0.931056
R19999 XThC.Tn[4].n42 XThC.Tn[4] 0.931056
R20000 XThC.Tn[4].n45 XThC.Tn[4] 0.931056
R20001 XThC.Tn[4].n48 XThC.Tn[4] 0.931056
R20002 XThC.Tn[4].n51 XThC.Tn[4] 0.931056
R20003 XThC.Tn[4].n54 XThC.Tn[4] 0.931056
R20004 XThC.Tn[4].n57 XThC.Tn[4] 0.931056
R20005 XThC.Tn[4] XThC.Tn[4].n60 0.6405
R20006 XThC.Tn[4] XThC.Tn[4].n12 0.396333
R20007 XThC.Tn[4] XThC.Tn[4].n15 0.396333
R20008 XThC.Tn[4] XThC.Tn[4].n18 0.396333
R20009 XThC.Tn[4] XThC.Tn[4].n21 0.396333
R20010 XThC.Tn[4] XThC.Tn[4].n24 0.396333
R20011 XThC.Tn[4] XThC.Tn[4].n27 0.396333
R20012 XThC.Tn[4] XThC.Tn[4].n30 0.396333
R20013 XThC.Tn[4] XThC.Tn[4].n33 0.396333
R20014 XThC.Tn[4] XThC.Tn[4].n36 0.396333
R20015 XThC.Tn[4] XThC.Tn[4].n39 0.396333
R20016 XThC.Tn[4] XThC.Tn[4].n42 0.396333
R20017 XThC.Tn[4] XThC.Tn[4].n45 0.396333
R20018 XThC.Tn[4] XThC.Tn[4].n48 0.396333
R20019 XThC.Tn[4] XThC.Tn[4].n51 0.396333
R20020 XThC.Tn[4] XThC.Tn[4].n54 0.396333
R20021 XThC.Tn[4] XThC.Tn[4].n57 0.396333
R20022 XThC.Tn[4].n11 XThC.Tn[4] 0.104667
R20023 XThC.Tn[4].n14 XThC.Tn[4] 0.104667
R20024 XThC.Tn[4].n17 XThC.Tn[4] 0.104667
R20025 XThC.Tn[4].n20 XThC.Tn[4] 0.104667
R20026 XThC.Tn[4].n23 XThC.Tn[4] 0.104667
R20027 XThC.Tn[4].n26 XThC.Tn[4] 0.104667
R20028 XThC.Tn[4].n29 XThC.Tn[4] 0.104667
R20029 XThC.Tn[4].n32 XThC.Tn[4] 0.104667
R20030 XThC.Tn[4].n35 XThC.Tn[4] 0.104667
R20031 XThC.Tn[4].n38 XThC.Tn[4] 0.104667
R20032 XThC.Tn[4].n41 XThC.Tn[4] 0.104667
R20033 XThC.Tn[4].n44 XThC.Tn[4] 0.104667
R20034 XThC.Tn[4].n47 XThC.Tn[4] 0.104667
R20035 XThC.Tn[4].n50 XThC.Tn[4] 0.104667
R20036 XThC.Tn[4].n53 XThC.Tn[4] 0.104667
R20037 XThC.Tn[4].n56 XThC.Tn[4] 0.104667
R20038 XThC.Tn[4].n11 XThC.Tn[4] 0.0309878
R20039 XThC.Tn[4].n14 XThC.Tn[4] 0.0309878
R20040 XThC.Tn[4].n17 XThC.Tn[4] 0.0309878
R20041 XThC.Tn[4].n20 XThC.Tn[4] 0.0309878
R20042 XThC.Tn[4].n23 XThC.Tn[4] 0.0309878
R20043 XThC.Tn[4].n26 XThC.Tn[4] 0.0309878
R20044 XThC.Tn[4].n29 XThC.Tn[4] 0.0309878
R20045 XThC.Tn[4].n32 XThC.Tn[4] 0.0309878
R20046 XThC.Tn[4].n35 XThC.Tn[4] 0.0309878
R20047 XThC.Tn[4].n38 XThC.Tn[4] 0.0309878
R20048 XThC.Tn[4].n41 XThC.Tn[4] 0.0309878
R20049 XThC.Tn[4].n44 XThC.Tn[4] 0.0309878
R20050 XThC.Tn[4].n47 XThC.Tn[4] 0.0309878
R20051 XThC.Tn[4].n50 XThC.Tn[4] 0.0309878
R20052 XThC.Tn[4].n53 XThC.Tn[4] 0.0309878
R20053 XThC.Tn[4].n56 XThC.Tn[4] 0.0309878
R20054 XThC.Tn[4].n12 XThC.Tn[4].n11 0.027939
R20055 XThC.Tn[4].n15 XThC.Tn[4].n14 0.027939
R20056 XThC.Tn[4].n18 XThC.Tn[4].n17 0.027939
R20057 XThC.Tn[4].n21 XThC.Tn[4].n20 0.027939
R20058 XThC.Tn[4].n24 XThC.Tn[4].n23 0.027939
R20059 XThC.Tn[4].n27 XThC.Tn[4].n26 0.027939
R20060 XThC.Tn[4].n30 XThC.Tn[4].n29 0.027939
R20061 XThC.Tn[4].n33 XThC.Tn[4].n32 0.027939
R20062 XThC.Tn[4].n36 XThC.Tn[4].n35 0.027939
R20063 XThC.Tn[4].n39 XThC.Tn[4].n38 0.027939
R20064 XThC.Tn[4].n42 XThC.Tn[4].n41 0.027939
R20065 XThC.Tn[4].n45 XThC.Tn[4].n44 0.027939
R20066 XThC.Tn[4].n48 XThC.Tn[4].n47 0.027939
R20067 XThC.Tn[4].n51 XThC.Tn[4].n50 0.027939
R20068 XThC.Tn[4].n54 XThC.Tn[4].n53 0.027939
R20069 XThC.Tn[4].n57 XThC.Tn[4].n56 0.027939
R20070 XThC.Tn[4].n58 XThC.Tn[4] 0.0129465
R20071 XThC.Tn[2].n2 XThC.Tn[2].n1 332.332
R20072 XThC.Tn[2].n2 XThC.Tn[2].n0 296.493
R20073 XThC.Tn[2].n12 XThC.Tn[2].n10 161.406
R20074 XThC.Tn[2].n15 XThC.Tn[2].n13 161.406
R20075 XThC.Tn[2].n18 XThC.Tn[2].n16 161.406
R20076 XThC.Tn[2].n21 XThC.Tn[2].n19 161.406
R20077 XThC.Tn[2].n24 XThC.Tn[2].n22 161.406
R20078 XThC.Tn[2].n27 XThC.Tn[2].n25 161.406
R20079 XThC.Tn[2].n30 XThC.Tn[2].n28 161.406
R20080 XThC.Tn[2].n33 XThC.Tn[2].n31 161.406
R20081 XThC.Tn[2].n36 XThC.Tn[2].n34 161.406
R20082 XThC.Tn[2].n39 XThC.Tn[2].n37 161.406
R20083 XThC.Tn[2].n42 XThC.Tn[2].n40 161.406
R20084 XThC.Tn[2].n45 XThC.Tn[2].n43 161.406
R20085 XThC.Tn[2].n48 XThC.Tn[2].n46 161.406
R20086 XThC.Tn[2].n51 XThC.Tn[2].n49 161.406
R20087 XThC.Tn[2].n54 XThC.Tn[2].n52 161.406
R20088 XThC.Tn[2].n57 XThC.Tn[2].n55 161.406
R20089 XThC.Tn[2].n10 XThC.Tn[2].t18 161.202
R20090 XThC.Tn[2].n13 XThC.Tn[2].t35 161.202
R20091 XThC.Tn[2].n16 XThC.Tn[2].t37 161.202
R20092 XThC.Tn[2].n19 XThC.Tn[2].t39 161.202
R20093 XThC.Tn[2].n22 XThC.Tn[2].t28 161.202
R20094 XThC.Tn[2].n25 XThC.Tn[2].t29 161.202
R20095 XThC.Tn[2].n28 XThC.Tn[2].t42 161.202
R20096 XThC.Tn[2].n31 XThC.Tn[2].t19 161.202
R20097 XThC.Tn[2].n34 XThC.Tn[2].t21 161.202
R20098 XThC.Tn[2].n37 XThC.Tn[2].t40 161.202
R20099 XThC.Tn[2].n40 XThC.Tn[2].t41 161.202
R20100 XThC.Tn[2].n43 XThC.Tn[2].t22 161.202
R20101 XThC.Tn[2].n46 XThC.Tn[2].t30 161.202
R20102 XThC.Tn[2].n49 XThC.Tn[2].t33 161.202
R20103 XThC.Tn[2].n52 XThC.Tn[2].t14 161.202
R20104 XThC.Tn[2].n55 XThC.Tn[2].t24 161.202
R20105 XThC.Tn[2].n10 XThC.Tn[2].t20 145.137
R20106 XThC.Tn[2].n13 XThC.Tn[2].t38 145.137
R20107 XThC.Tn[2].n16 XThC.Tn[2].t43 145.137
R20108 XThC.Tn[2].n19 XThC.Tn[2].t12 145.137
R20109 XThC.Tn[2].n22 XThC.Tn[2].t31 145.137
R20110 XThC.Tn[2].n25 XThC.Tn[2].t32 145.137
R20111 XThC.Tn[2].n28 XThC.Tn[2].t16 145.137
R20112 XThC.Tn[2].n31 XThC.Tn[2].t23 145.137
R20113 XThC.Tn[2].n34 XThC.Tn[2].t25 145.137
R20114 XThC.Tn[2].n37 XThC.Tn[2].t13 145.137
R20115 XThC.Tn[2].n40 XThC.Tn[2].t15 145.137
R20116 XThC.Tn[2].n43 XThC.Tn[2].t26 145.137
R20117 XThC.Tn[2].n46 XThC.Tn[2].t34 145.137
R20118 XThC.Tn[2].n49 XThC.Tn[2].t36 145.137
R20119 XThC.Tn[2].n52 XThC.Tn[2].t17 145.137
R20120 XThC.Tn[2].n55 XThC.Tn[2].t27 145.137
R20121 XThC.Tn[2].n7 XThC.Tn[2].n5 135.248
R20122 XThC.Tn[2].n9 XThC.Tn[2].n3 98.982
R20123 XThC.Tn[2].n8 XThC.Tn[2].n4 98.982
R20124 XThC.Tn[2].n7 XThC.Tn[2].n6 98.982
R20125 XThC.Tn[2].n9 XThC.Tn[2].n8 36.2672
R20126 XThC.Tn[2].n8 XThC.Tn[2].n7 36.2672
R20127 XThC.Tn[2].n59 XThC.Tn[2].n9 32.6405
R20128 XThC.Tn[2].n1 XThC.Tn[2].t2 26.5955
R20129 XThC.Tn[2].n1 XThC.Tn[2].t1 26.5955
R20130 XThC.Tn[2].n0 XThC.Tn[2].t4 26.5955
R20131 XThC.Tn[2].n0 XThC.Tn[2].t3 26.5955
R20132 XThC.Tn[2].n3 XThC.Tn[2].t8 24.9236
R20133 XThC.Tn[2].n3 XThC.Tn[2].t7 24.9236
R20134 XThC.Tn[2].n4 XThC.Tn[2].t6 24.9236
R20135 XThC.Tn[2].n4 XThC.Tn[2].t5 24.9236
R20136 XThC.Tn[2].n5 XThC.Tn[2].t9 24.9236
R20137 XThC.Tn[2].n5 XThC.Tn[2].t10 24.9236
R20138 XThC.Tn[2].n6 XThC.Tn[2].t11 24.9236
R20139 XThC.Tn[2].n6 XThC.Tn[2].t0 24.9236
R20140 XThC.Tn[2].n60 XThC.Tn[2].n2 18.5605
R20141 XThC.Tn[2].n60 XThC.Tn[2].n59 11.5205
R20142 XThC.Tn[2].n58 XThC.Tn[2] 6.32799
R20143 XThC.Tn[2].n59 XThC.Tn[2].n58 3.18175
R20144 XThC.Tn[2].n15 XThC.Tn[2] 0.931056
R20145 XThC.Tn[2].n18 XThC.Tn[2] 0.931056
R20146 XThC.Tn[2].n21 XThC.Tn[2] 0.931056
R20147 XThC.Tn[2].n24 XThC.Tn[2] 0.931056
R20148 XThC.Tn[2].n27 XThC.Tn[2] 0.931056
R20149 XThC.Tn[2].n30 XThC.Tn[2] 0.931056
R20150 XThC.Tn[2].n33 XThC.Tn[2] 0.931056
R20151 XThC.Tn[2].n36 XThC.Tn[2] 0.931056
R20152 XThC.Tn[2].n39 XThC.Tn[2] 0.931056
R20153 XThC.Tn[2].n42 XThC.Tn[2] 0.931056
R20154 XThC.Tn[2].n45 XThC.Tn[2] 0.931056
R20155 XThC.Tn[2].n48 XThC.Tn[2] 0.931056
R20156 XThC.Tn[2].n51 XThC.Tn[2] 0.931056
R20157 XThC.Tn[2].n54 XThC.Tn[2] 0.931056
R20158 XThC.Tn[2].n57 XThC.Tn[2] 0.931056
R20159 XThC.Tn[2] XThC.Tn[2].n60 0.6405
R20160 XThC.Tn[2] XThC.Tn[2].n12 0.396333
R20161 XThC.Tn[2] XThC.Tn[2].n15 0.396333
R20162 XThC.Tn[2] XThC.Tn[2].n18 0.396333
R20163 XThC.Tn[2] XThC.Tn[2].n21 0.396333
R20164 XThC.Tn[2] XThC.Tn[2].n24 0.396333
R20165 XThC.Tn[2] XThC.Tn[2].n27 0.396333
R20166 XThC.Tn[2] XThC.Tn[2].n30 0.396333
R20167 XThC.Tn[2] XThC.Tn[2].n33 0.396333
R20168 XThC.Tn[2] XThC.Tn[2].n36 0.396333
R20169 XThC.Tn[2] XThC.Tn[2].n39 0.396333
R20170 XThC.Tn[2] XThC.Tn[2].n42 0.396333
R20171 XThC.Tn[2] XThC.Tn[2].n45 0.396333
R20172 XThC.Tn[2] XThC.Tn[2].n48 0.396333
R20173 XThC.Tn[2] XThC.Tn[2].n51 0.396333
R20174 XThC.Tn[2] XThC.Tn[2].n54 0.396333
R20175 XThC.Tn[2] XThC.Tn[2].n57 0.396333
R20176 XThC.Tn[2].n11 XThC.Tn[2] 0.104667
R20177 XThC.Tn[2].n14 XThC.Tn[2] 0.104667
R20178 XThC.Tn[2].n17 XThC.Tn[2] 0.104667
R20179 XThC.Tn[2].n20 XThC.Tn[2] 0.104667
R20180 XThC.Tn[2].n23 XThC.Tn[2] 0.104667
R20181 XThC.Tn[2].n26 XThC.Tn[2] 0.104667
R20182 XThC.Tn[2].n29 XThC.Tn[2] 0.104667
R20183 XThC.Tn[2].n32 XThC.Tn[2] 0.104667
R20184 XThC.Tn[2].n35 XThC.Tn[2] 0.104667
R20185 XThC.Tn[2].n38 XThC.Tn[2] 0.104667
R20186 XThC.Tn[2].n41 XThC.Tn[2] 0.104667
R20187 XThC.Tn[2].n44 XThC.Tn[2] 0.104667
R20188 XThC.Tn[2].n47 XThC.Tn[2] 0.104667
R20189 XThC.Tn[2].n50 XThC.Tn[2] 0.104667
R20190 XThC.Tn[2].n53 XThC.Tn[2] 0.104667
R20191 XThC.Tn[2].n56 XThC.Tn[2] 0.104667
R20192 XThC.Tn[2].n11 XThC.Tn[2] 0.0309878
R20193 XThC.Tn[2].n14 XThC.Tn[2] 0.0309878
R20194 XThC.Tn[2].n17 XThC.Tn[2] 0.0309878
R20195 XThC.Tn[2].n20 XThC.Tn[2] 0.0309878
R20196 XThC.Tn[2].n23 XThC.Tn[2] 0.0309878
R20197 XThC.Tn[2].n26 XThC.Tn[2] 0.0309878
R20198 XThC.Tn[2].n29 XThC.Tn[2] 0.0309878
R20199 XThC.Tn[2].n32 XThC.Tn[2] 0.0309878
R20200 XThC.Tn[2].n35 XThC.Tn[2] 0.0309878
R20201 XThC.Tn[2].n38 XThC.Tn[2] 0.0309878
R20202 XThC.Tn[2].n41 XThC.Tn[2] 0.0309878
R20203 XThC.Tn[2].n44 XThC.Tn[2] 0.0309878
R20204 XThC.Tn[2].n47 XThC.Tn[2] 0.0309878
R20205 XThC.Tn[2].n50 XThC.Tn[2] 0.0309878
R20206 XThC.Tn[2].n53 XThC.Tn[2] 0.0309878
R20207 XThC.Tn[2].n56 XThC.Tn[2] 0.0309878
R20208 XThC.Tn[2].n12 XThC.Tn[2].n11 0.027939
R20209 XThC.Tn[2].n15 XThC.Tn[2].n14 0.027939
R20210 XThC.Tn[2].n18 XThC.Tn[2].n17 0.027939
R20211 XThC.Tn[2].n21 XThC.Tn[2].n20 0.027939
R20212 XThC.Tn[2].n24 XThC.Tn[2].n23 0.027939
R20213 XThC.Tn[2].n27 XThC.Tn[2].n26 0.027939
R20214 XThC.Tn[2].n30 XThC.Tn[2].n29 0.027939
R20215 XThC.Tn[2].n33 XThC.Tn[2].n32 0.027939
R20216 XThC.Tn[2].n36 XThC.Tn[2].n35 0.027939
R20217 XThC.Tn[2].n39 XThC.Tn[2].n38 0.027939
R20218 XThC.Tn[2].n42 XThC.Tn[2].n41 0.027939
R20219 XThC.Tn[2].n45 XThC.Tn[2].n44 0.027939
R20220 XThC.Tn[2].n48 XThC.Tn[2].n47 0.027939
R20221 XThC.Tn[2].n51 XThC.Tn[2].n50 0.027939
R20222 XThC.Tn[2].n54 XThC.Tn[2].n53 0.027939
R20223 XThC.Tn[2].n57 XThC.Tn[2].n56 0.027939
R20224 XThC.Tn[2].n58 XThC.Tn[2] 0.0156819
R20225 Vbias.n512 Vbias.t4 651.571
R20226 Vbias.n512 Vbias.t3 651.571
R20227 Vbias.n513 Vbias.t0 651.571
R20228 Vbias.n513 Vbias.t5 651.571
R20229 Vbias.n509 Vbias.t181 119.309
R20230 Vbias.n507 Vbias.t24 119.309
R20231 Vbias.n505 Vbias.t12 119.309
R20232 Vbias.n503 Vbias.t248 119.309
R20233 Vbias.n501 Vbias.t95 119.309
R20234 Vbias.n499 Vbias.t75 119.309
R20235 Vbias.n497 Vbias.t246 119.309
R20236 Vbias.n495 Vbias.t169 119.309
R20237 Vbias.n493 Vbias.t147 119.309
R20238 Vbias.n491 Vbias.t60 119.309
R20239 Vbias.n489 Vbias.t227 119.309
R20240 Vbias.n487 Vbias.t141 119.309
R20241 Vbias.n485 Vbias.t56 119.309
R20242 Vbias.n483 Vbias.t41 119.309
R20243 Vbias.n481 Vbias.t201 119.309
R20244 Vbias.n480 Vbias.t129 119.309
R20245 Vbias.n477 Vbias.t110 119.309
R20246 Vbias.n475 Vbias.t210 119.309
R20247 Vbias.n473 Vbias.t193 119.309
R20248 Vbias.n471 Vbias.t173 119.309
R20249 Vbias.n469 Vbias.t25 119.309
R20250 Vbias.n467 Vbias.t258 119.309
R20251 Vbias.n465 Vbias.t171 119.309
R20252 Vbias.n463 Vbias.t96 119.309
R20253 Vbias.n461 Vbias.t76 119.309
R20254 Vbias.n459 Vbias.t247 119.309
R20255 Vbias.n457 Vbias.t156 119.309
R20256 Vbias.n455 Vbias.t69 119.309
R20257 Vbias.n453 Vbias.t242 119.309
R20258 Vbias.n451 Vbias.t229 119.309
R20259 Vbias.n449 Vbias.t130 119.309
R20260 Vbias.n448 Vbias.t57 119.309
R20261 Vbias.n445 Vbias.t146 119.309
R20262 Vbias.n443 Vbias.t238 119.309
R20263 Vbias.n441 Vbias.t225 119.309
R20264 Vbias.n439 Vbias.t205 119.309
R20265 Vbias.n437 Vbias.t52 119.309
R20266 Vbias.n435 Vbias.t32 119.309
R20267 Vbias.n433 Vbias.t199 119.309
R20268 Vbias.n431 Vbias.t125 119.309
R20269 Vbias.n429 Vbias.t102 119.309
R20270 Vbias.n427 Vbias.t18 119.309
R20271 Vbias.n425 Vbias.t183 119.309
R20272 Vbias.n423 Vbias.t99 119.309
R20273 Vbias.n421 Vbias.t14 119.309
R20274 Vbias.n419 Vbias.t261 119.309
R20275 Vbias.n417 Vbias.t160 119.309
R20276 Vbias.n416 Vbias.t87 119.309
R20277 Vbias.n413 Vbias.t73 119.309
R20278 Vbias.n411 Vbias.t165 119.309
R20279 Vbias.n409 Vbias.t153 119.309
R20280 Vbias.n407 Vbias.t133 119.309
R20281 Vbias.n405 Vbias.t239 119.309
R20282 Vbias.n403 Vbias.t217 119.309
R20283 Vbias.n401 Vbias.t126 119.309
R20284 Vbias.n399 Vbias.t53 119.309
R20285 Vbias.n397 Vbias.t33 119.309
R20286 Vbias.n395 Vbias.t200 119.309
R20287 Vbias.n393 Vbias.t112 119.309
R20288 Vbias.n391 Vbias.t29 119.309
R20289 Vbias.n389 Vbias.t196 119.309
R20290 Vbias.n387 Vbias.t185 119.309
R20291 Vbias.n385 Vbias.t88 119.309
R20292 Vbias.n384 Vbias.t16 119.309
R20293 Vbias.n381 Vbias.t255 119.309
R20294 Vbias.n379 Vbias.t92 119.309
R20295 Vbias.n377 Vbias.t81 119.309
R20296 Vbias.n375 Vbias.t62 119.309
R20297 Vbias.n373 Vbias.t166 119.309
R20298 Vbias.n371 Vbias.t144 119.309
R20299 Vbias.n369 Vbias.t54 119.309
R20300 Vbias.n367 Vbias.t240 119.309
R20301 Vbias.n365 Vbias.t219 119.309
R20302 Vbias.n363 Vbias.t127 119.309
R20303 Vbias.n361 Vbias.t40 119.309
R20304 Vbias.n359 Vbias.t213 119.309
R20305 Vbias.n357 Vbias.t124 119.309
R20306 Vbias.n355 Vbias.t113 119.309
R20307 Vbias.n353 Vbias.t17 119.309
R20308 Vbias.n352 Vbias.t198 119.309
R20309 Vbias.n349 Vbias.t176 119.309
R20310 Vbias.n347 Vbias.t20 119.309
R20311 Vbias.n345 Vbias.t7 119.309
R20312 Vbias.n343 Vbias.t243 119.309
R20313 Vbias.n341 Vbias.t90 119.309
R20314 Vbias.n339 Vbias.t65 119.309
R20315 Vbias.n337 Vbias.t236 119.309
R20316 Vbias.n335 Vbias.t163 119.309
R20317 Vbias.n333 Vbias.t138 119.309
R20318 Vbias.n331 Vbias.t50 119.309
R20319 Vbias.n329 Vbias.t221 119.309
R20320 Vbias.n327 Vbias.t135 119.309
R20321 Vbias.n325 Vbias.t48 119.309
R20322 Vbias.n323 Vbias.t37 119.309
R20323 Vbias.n321 Vbias.t195 119.309
R20324 Vbias.n320 Vbias.t121 119.309
R20325 Vbias.n317 Vbias.t105 119.309
R20326 Vbias.n315 Vbias.t204 119.309
R20327 Vbias.n313 Vbias.t187 119.309
R20328 Vbias.n311 Vbias.t168 119.309
R20329 Vbias.n309 Vbias.t21 119.309
R20330 Vbias.n307 Vbias.t251 119.309
R20331 Vbias.n305 Vbias.t164 119.309
R20332 Vbias.n303 Vbias.t91 119.309
R20333 Vbias.n301 Vbias.t68 119.309
R20334 Vbias.n299 Vbias.t237 119.309
R20335 Vbias.n297 Vbias.t150 119.309
R20336 Vbias.n295 Vbias.t63 119.309
R20337 Vbias.n293 Vbias.t235 119.309
R20338 Vbias.n291 Vbias.t222 119.309
R20339 Vbias.n289 Vbias.t122 119.309
R20340 Vbias.n288 Vbias.t49 119.309
R20341 Vbias.n285 Vbias.t137 119.309
R20342 Vbias.n283 Vbias.t232 119.309
R20343 Vbias.n281 Vbias.t220 119.309
R20344 Vbias.n279 Vbias.t197 119.309
R20345 Vbias.n277 Vbias.t44 119.309
R20346 Vbias.n275 Vbias.t27 119.309
R20347 Vbias.n273 Vbias.t190 119.309
R20348 Vbias.n271 Vbias.t118 119.309
R20349 Vbias.n269 Vbias.t98 119.309
R20350 Vbias.n267 Vbias.t11 119.309
R20351 Vbias.n265 Vbias.t179 119.309
R20352 Vbias.n263 Vbias.t93 119.309
R20353 Vbias.n261 Vbias.t8 119.309
R20354 Vbias.n259 Vbias.t257 119.309
R20355 Vbias.n257 Vbias.t154 119.309
R20356 Vbias.n256 Vbias.t82 119.309
R20357 Vbias.n253 Vbias.t64 119.309
R20358 Vbias.n251 Vbias.t161 119.309
R20359 Vbias.n249 Vbias.t149 119.309
R20360 Vbias.n247 Vbias.t123 119.309
R20361 Vbias.n245 Vbias.t233 119.309
R20362 Vbias.n243 Vbias.t211 119.309
R20363 Vbias.n241 Vbias.t119 119.309
R20364 Vbias.n239 Vbias.t45 119.309
R20365 Vbias.n237 Vbias.t28 119.309
R20366 Vbias.n235 Vbias.t192 119.309
R20367 Vbias.n233 Vbias.t107 119.309
R20368 Vbias.n231 Vbias.t23 119.309
R20369 Vbias.n229 Vbias.t188 119.309
R20370 Vbias.n227 Vbias.t180 119.309
R20371 Vbias.n225 Vbias.t83 119.309
R20372 Vbias.n224 Vbias.t9 119.309
R20373 Vbias.n221 Vbias.t250 119.309
R20374 Vbias.n219 Vbias.t89 119.309
R20375 Vbias.n217 Vbias.t80 119.309
R20376 Vbias.n215 Vbias.t51 119.309
R20377 Vbias.n213 Vbias.t162 119.309
R20378 Vbias.n211 Vbias.t136 119.309
R20379 Vbias.n209 Vbias.t46 119.309
R20380 Vbias.n207 Vbias.t234 119.309
R20381 Vbias.n205 Vbias.t212 119.309
R20382 Vbias.n203 Vbias.t120 119.309
R20383 Vbias.n201 Vbias.t36 119.309
R20384 Vbias.n199 Vbias.t208 119.309
R20385 Vbias.n197 Vbias.t117 119.309
R20386 Vbias.n195 Vbias.t108 119.309
R20387 Vbias.n193 Vbias.t10 119.309
R20388 Vbias.n192 Vbias.t189 119.309
R20389 Vbias.n189 Vbias.t109 119.309
R20390 Vbias.n187 Vbias.t207 119.309
R20391 Vbias.n185 Vbias.t191 119.309
R20392 Vbias.n183 Vbias.t172 119.309
R20393 Vbias.n181 Vbias.t22 119.309
R20394 Vbias.n179 Vbias.t256 119.309
R20395 Vbias.n177 Vbias.t167 119.309
R20396 Vbias.n175 Vbias.t94 119.309
R20397 Vbias.n173 Vbias.t74 119.309
R20398 Vbias.n171 Vbias.t244 119.309
R20399 Vbias.n169 Vbias.t155 119.309
R20400 Vbias.n167 Vbias.t66 119.309
R20401 Vbias.n165 Vbias.t241 119.309
R20402 Vbias.n163 Vbias.t226 119.309
R20403 Vbias.n161 Vbias.t128 119.309
R20404 Vbias.n160 Vbias.t55 119.309
R20405 Vbias.n157 Vbias.t249 119.309
R20406 Vbias.n155 Vbias.t85 119.309
R20407 Vbias.n153 Vbias.t78 119.309
R20408 Vbias.n151 Vbias.t47 119.309
R20409 Vbias.n149 Vbias.t159 119.309
R20410 Vbias.n147 Vbias.t134 119.309
R20411 Vbias.n145 Vbias.t43 119.309
R20412 Vbias.n143 Vbias.t231 119.309
R20413 Vbias.n141 Vbias.t209 119.309
R20414 Vbias.n139 Vbias.t116 119.309
R20415 Vbias.n137 Vbias.t34 119.309
R20416 Vbias.n135 Vbias.t206 119.309
R20417 Vbias.n133 Vbias.t115 119.309
R20418 Vbias.n131 Vbias.t103 119.309
R20419 Vbias.n129 Vbias.t6 119.309
R20420 Vbias.n128 Vbias.t186 119.309
R20421 Vbias.n125 Vbias.t86 119.309
R20422 Vbias.n123 Vbias.t175 119.309
R20423 Vbias.n121 Vbias.t170 119.309
R20424 Vbias.n119 Vbias.t148 119.309
R20425 Vbias.n117 Vbias.t252 119.309
R20426 Vbias.n115 Vbias.t228 119.309
R20427 Vbias.n113 Vbias.t143 119.309
R20428 Vbias.n111 Vbias.t70 119.309
R20429 Vbias.n109 Vbias.t42 119.309
R20430 Vbias.n107 Vbias.t218 119.309
R20431 Vbias.n105 Vbias.t131 119.309
R20432 Vbias.n103 Vbias.t38 119.309
R20433 Vbias.n101 Vbias.t214 119.309
R20434 Vbias.n99 Vbias.t203 119.309
R20435 Vbias.n97 Vbias.t100 119.309
R20436 Vbias.n96 Vbias.t30 119.309
R20437 Vbias.n93 Vbias.t13 119.309
R20438 Vbias.n91 Vbias.t104 119.309
R20439 Vbias.n89 Vbias.t97 119.309
R20440 Vbias.n87 Vbias.t77 119.309
R20441 Vbias.n85 Vbias.t177 119.309
R20442 Vbias.n83 Vbias.t157 119.309
R20443 Vbias.n81 Vbias.t71 119.309
R20444 Vbias.n79 Vbias.t253 119.309
R20445 Vbias.n77 Vbias.t230 119.309
R20446 Vbias.n75 Vbias.t145 119.309
R20447 Vbias.n73 Vbias.t58 119.309
R20448 Vbias.n71 Vbias.t224 119.309
R20449 Vbias.n69 Vbias.t139 119.309
R20450 Vbias.n67 Vbias.t132 119.309
R20451 Vbias.n65 Vbias.t31 119.309
R20452 Vbias.n64 Vbias.t215 119.309
R20453 Vbias.n61 Vbias.t194 119.309
R20454 Vbias.n59 Vbias.t35 119.309
R20455 Vbias.n57 Vbias.t26 119.309
R20456 Vbias.n55 Vbias.t259 119.309
R20457 Vbias.n53 Vbias.t106 119.309
R20458 Vbias.n51 Vbias.t84 119.309
R20459 Vbias.n49 Vbias.t254 119.309
R20460 Vbias.n47 Vbias.t178 119.309
R20461 Vbias.n45 Vbias.t158 119.309
R20462 Vbias.n43 Vbias.t72 119.309
R20463 Vbias.n41 Vbias.t245 119.309
R20464 Vbias.n39 Vbias.t152 119.309
R20465 Vbias.n37 Vbias.t67 119.309
R20466 Vbias.n35 Vbias.t59 119.309
R20467 Vbias.n33 Vbias.t216 119.309
R20468 Vbias.n32 Vbias.t140 119.309
R20469 Vbias.n29 Vbias.t61 119.309
R20470 Vbias.n27 Vbias.t151 119.309
R20471 Vbias.n25 Vbias.t142 119.309
R20472 Vbias.n23 Vbias.t114 119.309
R20473 Vbias.n21 Vbias.t223 119.309
R20474 Vbias.n19 Vbias.t202 119.309
R20475 Vbias.n17 Vbias.t111 119.309
R20476 Vbias.n15 Vbias.t39 119.309
R20477 Vbias.n13 Vbias.t19 119.309
R20478 Vbias.n11 Vbias.t184 119.309
R20479 Vbias.n9 Vbias.t101 119.309
R20480 Vbias.n7 Vbias.t15 119.309
R20481 Vbias.n5 Vbias.t182 119.309
R20482 Vbias.n3 Vbias.t174 119.309
R20483 Vbias.n1 Vbias.t79 119.309
R20484 Vbias.n0 Vbias.t260 119.309
R20485 Vbias.n515 Vbias.t1 77.1775
R20486 Vbias.n515 Vbias.t2 34.3847
R20487 Vbias Vbias.n480 8.00727
R20488 Vbias Vbias.n448 8.00727
R20489 Vbias Vbias.n416 8.00727
R20490 Vbias Vbias.n384 8.00727
R20491 Vbias Vbias.n352 8.00727
R20492 Vbias Vbias.n320 8.00727
R20493 Vbias Vbias.n288 8.00727
R20494 Vbias Vbias.n256 8.00727
R20495 Vbias Vbias.n224 8.00727
R20496 Vbias Vbias.n192 8.00727
R20497 Vbias Vbias.n160 8.00727
R20498 Vbias Vbias.n128 8.00727
R20499 Vbias Vbias.n96 8.00727
R20500 Vbias Vbias.n64 8.00727
R20501 Vbias Vbias.n32 8.00727
R20502 Vbias Vbias.n0 8.00727
R20503 Vbias.n510 Vbias.n509 7.9105
R20504 Vbias.n508 Vbias.n507 7.9105
R20505 Vbias.n506 Vbias.n505 7.9105
R20506 Vbias.n504 Vbias.n503 7.9105
R20507 Vbias.n502 Vbias.n501 7.9105
R20508 Vbias.n500 Vbias.n499 7.9105
R20509 Vbias.n498 Vbias.n497 7.9105
R20510 Vbias.n496 Vbias.n495 7.9105
R20511 Vbias.n494 Vbias.n493 7.9105
R20512 Vbias.n492 Vbias.n491 7.9105
R20513 Vbias.n490 Vbias.n489 7.9105
R20514 Vbias.n488 Vbias.n487 7.9105
R20515 Vbias.n486 Vbias.n485 7.9105
R20516 Vbias.n484 Vbias.n483 7.9105
R20517 Vbias.n482 Vbias.n481 7.9105
R20518 Vbias.n478 Vbias.n477 7.9105
R20519 Vbias.n476 Vbias.n475 7.9105
R20520 Vbias.n474 Vbias.n473 7.9105
R20521 Vbias.n472 Vbias.n471 7.9105
R20522 Vbias.n470 Vbias.n469 7.9105
R20523 Vbias.n468 Vbias.n467 7.9105
R20524 Vbias.n466 Vbias.n465 7.9105
R20525 Vbias.n464 Vbias.n463 7.9105
R20526 Vbias.n462 Vbias.n461 7.9105
R20527 Vbias.n460 Vbias.n459 7.9105
R20528 Vbias.n458 Vbias.n457 7.9105
R20529 Vbias.n456 Vbias.n455 7.9105
R20530 Vbias.n454 Vbias.n453 7.9105
R20531 Vbias.n452 Vbias.n451 7.9105
R20532 Vbias.n450 Vbias.n449 7.9105
R20533 Vbias.n446 Vbias.n445 7.9105
R20534 Vbias.n444 Vbias.n443 7.9105
R20535 Vbias.n442 Vbias.n441 7.9105
R20536 Vbias.n440 Vbias.n439 7.9105
R20537 Vbias.n438 Vbias.n437 7.9105
R20538 Vbias.n436 Vbias.n435 7.9105
R20539 Vbias.n434 Vbias.n433 7.9105
R20540 Vbias.n432 Vbias.n431 7.9105
R20541 Vbias.n430 Vbias.n429 7.9105
R20542 Vbias.n428 Vbias.n427 7.9105
R20543 Vbias.n426 Vbias.n425 7.9105
R20544 Vbias.n424 Vbias.n423 7.9105
R20545 Vbias.n422 Vbias.n421 7.9105
R20546 Vbias.n420 Vbias.n419 7.9105
R20547 Vbias.n418 Vbias.n417 7.9105
R20548 Vbias.n414 Vbias.n413 7.9105
R20549 Vbias.n412 Vbias.n411 7.9105
R20550 Vbias.n410 Vbias.n409 7.9105
R20551 Vbias.n408 Vbias.n407 7.9105
R20552 Vbias.n406 Vbias.n405 7.9105
R20553 Vbias.n404 Vbias.n403 7.9105
R20554 Vbias.n402 Vbias.n401 7.9105
R20555 Vbias.n400 Vbias.n399 7.9105
R20556 Vbias.n398 Vbias.n397 7.9105
R20557 Vbias.n396 Vbias.n395 7.9105
R20558 Vbias.n394 Vbias.n393 7.9105
R20559 Vbias.n392 Vbias.n391 7.9105
R20560 Vbias.n390 Vbias.n389 7.9105
R20561 Vbias.n388 Vbias.n387 7.9105
R20562 Vbias.n386 Vbias.n385 7.9105
R20563 Vbias.n382 Vbias.n381 7.9105
R20564 Vbias.n380 Vbias.n379 7.9105
R20565 Vbias.n378 Vbias.n377 7.9105
R20566 Vbias.n376 Vbias.n375 7.9105
R20567 Vbias.n374 Vbias.n373 7.9105
R20568 Vbias.n372 Vbias.n371 7.9105
R20569 Vbias.n370 Vbias.n369 7.9105
R20570 Vbias.n368 Vbias.n367 7.9105
R20571 Vbias.n366 Vbias.n365 7.9105
R20572 Vbias.n364 Vbias.n363 7.9105
R20573 Vbias.n362 Vbias.n361 7.9105
R20574 Vbias.n360 Vbias.n359 7.9105
R20575 Vbias.n358 Vbias.n357 7.9105
R20576 Vbias.n356 Vbias.n355 7.9105
R20577 Vbias.n354 Vbias.n353 7.9105
R20578 Vbias.n350 Vbias.n349 7.9105
R20579 Vbias.n348 Vbias.n347 7.9105
R20580 Vbias.n346 Vbias.n345 7.9105
R20581 Vbias.n344 Vbias.n343 7.9105
R20582 Vbias.n342 Vbias.n341 7.9105
R20583 Vbias.n340 Vbias.n339 7.9105
R20584 Vbias.n338 Vbias.n337 7.9105
R20585 Vbias.n336 Vbias.n335 7.9105
R20586 Vbias.n334 Vbias.n333 7.9105
R20587 Vbias.n332 Vbias.n331 7.9105
R20588 Vbias.n330 Vbias.n329 7.9105
R20589 Vbias.n328 Vbias.n327 7.9105
R20590 Vbias.n326 Vbias.n325 7.9105
R20591 Vbias.n324 Vbias.n323 7.9105
R20592 Vbias.n322 Vbias.n321 7.9105
R20593 Vbias.n318 Vbias.n317 7.9105
R20594 Vbias.n316 Vbias.n315 7.9105
R20595 Vbias.n314 Vbias.n313 7.9105
R20596 Vbias.n312 Vbias.n311 7.9105
R20597 Vbias.n310 Vbias.n309 7.9105
R20598 Vbias.n308 Vbias.n307 7.9105
R20599 Vbias.n306 Vbias.n305 7.9105
R20600 Vbias.n304 Vbias.n303 7.9105
R20601 Vbias.n302 Vbias.n301 7.9105
R20602 Vbias.n300 Vbias.n299 7.9105
R20603 Vbias.n298 Vbias.n297 7.9105
R20604 Vbias.n296 Vbias.n295 7.9105
R20605 Vbias.n294 Vbias.n293 7.9105
R20606 Vbias.n292 Vbias.n291 7.9105
R20607 Vbias.n290 Vbias.n289 7.9105
R20608 Vbias.n286 Vbias.n285 7.9105
R20609 Vbias.n284 Vbias.n283 7.9105
R20610 Vbias.n282 Vbias.n281 7.9105
R20611 Vbias.n280 Vbias.n279 7.9105
R20612 Vbias.n278 Vbias.n277 7.9105
R20613 Vbias.n276 Vbias.n275 7.9105
R20614 Vbias.n274 Vbias.n273 7.9105
R20615 Vbias.n272 Vbias.n271 7.9105
R20616 Vbias.n270 Vbias.n269 7.9105
R20617 Vbias.n268 Vbias.n267 7.9105
R20618 Vbias.n266 Vbias.n265 7.9105
R20619 Vbias.n264 Vbias.n263 7.9105
R20620 Vbias.n262 Vbias.n261 7.9105
R20621 Vbias.n260 Vbias.n259 7.9105
R20622 Vbias.n258 Vbias.n257 7.9105
R20623 Vbias.n254 Vbias.n253 7.9105
R20624 Vbias.n252 Vbias.n251 7.9105
R20625 Vbias.n250 Vbias.n249 7.9105
R20626 Vbias.n248 Vbias.n247 7.9105
R20627 Vbias.n246 Vbias.n245 7.9105
R20628 Vbias.n244 Vbias.n243 7.9105
R20629 Vbias.n242 Vbias.n241 7.9105
R20630 Vbias.n240 Vbias.n239 7.9105
R20631 Vbias.n238 Vbias.n237 7.9105
R20632 Vbias.n236 Vbias.n235 7.9105
R20633 Vbias.n234 Vbias.n233 7.9105
R20634 Vbias.n232 Vbias.n231 7.9105
R20635 Vbias.n230 Vbias.n229 7.9105
R20636 Vbias.n228 Vbias.n227 7.9105
R20637 Vbias.n226 Vbias.n225 7.9105
R20638 Vbias.n222 Vbias.n221 7.9105
R20639 Vbias.n220 Vbias.n219 7.9105
R20640 Vbias.n218 Vbias.n217 7.9105
R20641 Vbias.n216 Vbias.n215 7.9105
R20642 Vbias.n214 Vbias.n213 7.9105
R20643 Vbias.n212 Vbias.n211 7.9105
R20644 Vbias.n210 Vbias.n209 7.9105
R20645 Vbias.n208 Vbias.n207 7.9105
R20646 Vbias.n206 Vbias.n205 7.9105
R20647 Vbias.n204 Vbias.n203 7.9105
R20648 Vbias.n202 Vbias.n201 7.9105
R20649 Vbias.n200 Vbias.n199 7.9105
R20650 Vbias.n198 Vbias.n197 7.9105
R20651 Vbias.n196 Vbias.n195 7.9105
R20652 Vbias.n194 Vbias.n193 7.9105
R20653 Vbias.n190 Vbias.n189 7.9105
R20654 Vbias.n188 Vbias.n187 7.9105
R20655 Vbias.n186 Vbias.n185 7.9105
R20656 Vbias.n184 Vbias.n183 7.9105
R20657 Vbias.n182 Vbias.n181 7.9105
R20658 Vbias.n180 Vbias.n179 7.9105
R20659 Vbias.n178 Vbias.n177 7.9105
R20660 Vbias.n176 Vbias.n175 7.9105
R20661 Vbias.n174 Vbias.n173 7.9105
R20662 Vbias.n172 Vbias.n171 7.9105
R20663 Vbias.n170 Vbias.n169 7.9105
R20664 Vbias.n168 Vbias.n167 7.9105
R20665 Vbias.n166 Vbias.n165 7.9105
R20666 Vbias.n164 Vbias.n163 7.9105
R20667 Vbias.n162 Vbias.n161 7.9105
R20668 Vbias.n158 Vbias.n157 7.9105
R20669 Vbias.n156 Vbias.n155 7.9105
R20670 Vbias.n154 Vbias.n153 7.9105
R20671 Vbias.n152 Vbias.n151 7.9105
R20672 Vbias.n150 Vbias.n149 7.9105
R20673 Vbias.n148 Vbias.n147 7.9105
R20674 Vbias.n146 Vbias.n145 7.9105
R20675 Vbias.n144 Vbias.n143 7.9105
R20676 Vbias.n142 Vbias.n141 7.9105
R20677 Vbias.n140 Vbias.n139 7.9105
R20678 Vbias.n138 Vbias.n137 7.9105
R20679 Vbias.n136 Vbias.n135 7.9105
R20680 Vbias.n134 Vbias.n133 7.9105
R20681 Vbias.n132 Vbias.n131 7.9105
R20682 Vbias.n130 Vbias.n129 7.9105
R20683 Vbias.n126 Vbias.n125 7.9105
R20684 Vbias.n124 Vbias.n123 7.9105
R20685 Vbias.n122 Vbias.n121 7.9105
R20686 Vbias.n120 Vbias.n119 7.9105
R20687 Vbias.n118 Vbias.n117 7.9105
R20688 Vbias.n116 Vbias.n115 7.9105
R20689 Vbias.n114 Vbias.n113 7.9105
R20690 Vbias.n112 Vbias.n111 7.9105
R20691 Vbias.n110 Vbias.n109 7.9105
R20692 Vbias.n108 Vbias.n107 7.9105
R20693 Vbias.n106 Vbias.n105 7.9105
R20694 Vbias.n104 Vbias.n103 7.9105
R20695 Vbias.n102 Vbias.n101 7.9105
R20696 Vbias.n100 Vbias.n99 7.9105
R20697 Vbias.n98 Vbias.n97 7.9105
R20698 Vbias.n94 Vbias.n93 7.9105
R20699 Vbias.n92 Vbias.n91 7.9105
R20700 Vbias.n90 Vbias.n89 7.9105
R20701 Vbias.n88 Vbias.n87 7.9105
R20702 Vbias.n86 Vbias.n85 7.9105
R20703 Vbias.n84 Vbias.n83 7.9105
R20704 Vbias.n82 Vbias.n81 7.9105
R20705 Vbias.n80 Vbias.n79 7.9105
R20706 Vbias.n78 Vbias.n77 7.9105
R20707 Vbias.n76 Vbias.n75 7.9105
R20708 Vbias.n74 Vbias.n73 7.9105
R20709 Vbias.n72 Vbias.n71 7.9105
R20710 Vbias.n70 Vbias.n69 7.9105
R20711 Vbias.n68 Vbias.n67 7.9105
R20712 Vbias.n66 Vbias.n65 7.9105
R20713 Vbias.n62 Vbias.n61 7.9105
R20714 Vbias.n60 Vbias.n59 7.9105
R20715 Vbias.n58 Vbias.n57 7.9105
R20716 Vbias.n56 Vbias.n55 7.9105
R20717 Vbias.n54 Vbias.n53 7.9105
R20718 Vbias.n52 Vbias.n51 7.9105
R20719 Vbias.n50 Vbias.n49 7.9105
R20720 Vbias.n48 Vbias.n47 7.9105
R20721 Vbias.n46 Vbias.n45 7.9105
R20722 Vbias.n44 Vbias.n43 7.9105
R20723 Vbias.n42 Vbias.n41 7.9105
R20724 Vbias.n40 Vbias.n39 7.9105
R20725 Vbias.n38 Vbias.n37 7.9105
R20726 Vbias.n36 Vbias.n35 7.9105
R20727 Vbias.n34 Vbias.n33 7.9105
R20728 Vbias.n30 Vbias.n29 7.9105
R20729 Vbias.n28 Vbias.n27 7.9105
R20730 Vbias.n26 Vbias.n25 7.9105
R20731 Vbias.n24 Vbias.n23 7.9105
R20732 Vbias.n22 Vbias.n21 7.9105
R20733 Vbias.n20 Vbias.n19 7.9105
R20734 Vbias.n18 Vbias.n17 7.9105
R20735 Vbias.n16 Vbias.n15 7.9105
R20736 Vbias.n14 Vbias.n13 7.9105
R20737 Vbias.n12 Vbias.n11 7.9105
R20738 Vbias.n10 Vbias.n9 7.9105
R20739 Vbias.n8 Vbias.n7 7.9105
R20740 Vbias.n6 Vbias.n5 7.9105
R20741 Vbias.n4 Vbias.n3 7.9105
R20742 Vbias.n2 Vbias.n1 7.9105
R20743 Vbias.n514 Vbias.n512 4.78773
R20744 Vbias.n514 Vbias.n513 4.78773
R20745 Vbias.n516 Vbias.n514 2.09636
R20746 Vbias.n511 Vbias 1.6647
R20747 Vbias.n479 Vbias 1.6647
R20748 Vbias.n447 Vbias 1.6647
R20749 Vbias.n415 Vbias 1.6647
R20750 Vbias.n383 Vbias 1.6647
R20751 Vbias.n351 Vbias 1.6647
R20752 Vbias.n319 Vbias 1.6647
R20753 Vbias.n287 Vbias 1.6647
R20754 Vbias.n255 Vbias 1.6647
R20755 Vbias.n223 Vbias 1.6647
R20756 Vbias.n191 Vbias 1.6647
R20757 Vbias.n159 Vbias 1.6647
R20758 Vbias.n127 Vbias 1.6647
R20759 Vbias.n95 Vbias 1.6647
R20760 Vbias.n63 Vbias 1.6647
R20761 Vbias.n31 Vbias 1.6647
R20762 Vbias.n517 Vbias 1.34721
R20763 Vbias Vbias.n516 0.752103
R20764 Vbias.n517 Vbias.n511 0.5692
R20765 Vbias.n516 Vbias.n515 0.515506
R20766 Vbias.n63 Vbias.n31 0.410967
R20767 Vbias.n95 Vbias.n63 0.410967
R20768 Vbias.n127 Vbias.n95 0.410967
R20769 Vbias.n159 Vbias.n127 0.410967
R20770 Vbias.n191 Vbias.n159 0.410967
R20771 Vbias.n223 Vbias.n191 0.410967
R20772 Vbias.n255 Vbias.n223 0.410967
R20773 Vbias.n287 Vbias.n255 0.410967
R20774 Vbias.n319 Vbias.n287 0.410967
R20775 Vbias.n351 Vbias.n319 0.410967
R20776 Vbias.n383 Vbias.n351 0.410967
R20777 Vbias.n415 Vbias.n383 0.410967
R20778 Vbias.n447 Vbias.n415 0.410967
R20779 Vbias.n479 Vbias.n447 0.410967
R20780 Vbias.n511 Vbias.n479 0.410967
R20781 Vbias.n31 Vbias 0.383811
R20782 Vbias.n482 Vbias 0.252372
R20783 Vbias.n484 Vbias 0.252372
R20784 Vbias.n486 Vbias 0.252372
R20785 Vbias.n488 Vbias 0.252372
R20786 Vbias.n490 Vbias 0.252372
R20787 Vbias.n492 Vbias 0.252372
R20788 Vbias.n494 Vbias 0.252372
R20789 Vbias.n496 Vbias 0.252372
R20790 Vbias.n498 Vbias 0.252372
R20791 Vbias.n500 Vbias 0.252372
R20792 Vbias.n502 Vbias 0.252372
R20793 Vbias.n504 Vbias 0.252372
R20794 Vbias.n506 Vbias 0.252372
R20795 Vbias.n508 Vbias 0.252372
R20796 Vbias.n510 Vbias 0.252372
R20797 Vbias.n450 Vbias 0.252372
R20798 Vbias.n452 Vbias 0.252372
R20799 Vbias.n454 Vbias 0.252372
R20800 Vbias.n456 Vbias 0.252372
R20801 Vbias.n458 Vbias 0.252372
R20802 Vbias.n460 Vbias 0.252372
R20803 Vbias.n462 Vbias 0.252372
R20804 Vbias.n464 Vbias 0.252372
R20805 Vbias.n466 Vbias 0.252372
R20806 Vbias.n468 Vbias 0.252372
R20807 Vbias.n470 Vbias 0.252372
R20808 Vbias.n472 Vbias 0.252372
R20809 Vbias.n474 Vbias 0.252372
R20810 Vbias.n476 Vbias 0.252372
R20811 Vbias.n478 Vbias 0.252372
R20812 Vbias.n418 Vbias 0.252372
R20813 Vbias.n420 Vbias 0.252372
R20814 Vbias.n422 Vbias 0.252372
R20815 Vbias.n424 Vbias 0.252372
R20816 Vbias.n426 Vbias 0.252372
R20817 Vbias.n428 Vbias 0.252372
R20818 Vbias.n430 Vbias 0.252372
R20819 Vbias.n432 Vbias 0.252372
R20820 Vbias.n434 Vbias 0.252372
R20821 Vbias.n436 Vbias 0.252372
R20822 Vbias.n438 Vbias 0.252372
R20823 Vbias.n440 Vbias 0.252372
R20824 Vbias.n442 Vbias 0.252372
R20825 Vbias.n444 Vbias 0.252372
R20826 Vbias.n446 Vbias 0.252372
R20827 Vbias.n386 Vbias 0.252372
R20828 Vbias.n388 Vbias 0.252372
R20829 Vbias.n390 Vbias 0.252372
R20830 Vbias.n392 Vbias 0.252372
R20831 Vbias.n394 Vbias 0.252372
R20832 Vbias.n396 Vbias 0.252372
R20833 Vbias.n398 Vbias 0.252372
R20834 Vbias.n400 Vbias 0.252372
R20835 Vbias.n402 Vbias 0.252372
R20836 Vbias.n404 Vbias 0.252372
R20837 Vbias.n406 Vbias 0.252372
R20838 Vbias.n408 Vbias 0.252372
R20839 Vbias.n410 Vbias 0.252372
R20840 Vbias.n412 Vbias 0.252372
R20841 Vbias.n414 Vbias 0.252372
R20842 Vbias.n354 Vbias 0.252372
R20843 Vbias.n356 Vbias 0.252372
R20844 Vbias.n358 Vbias 0.252372
R20845 Vbias.n360 Vbias 0.252372
R20846 Vbias.n362 Vbias 0.252372
R20847 Vbias.n364 Vbias 0.252372
R20848 Vbias.n366 Vbias 0.252372
R20849 Vbias.n368 Vbias 0.252372
R20850 Vbias.n370 Vbias 0.252372
R20851 Vbias.n372 Vbias 0.252372
R20852 Vbias.n374 Vbias 0.252372
R20853 Vbias.n376 Vbias 0.252372
R20854 Vbias.n378 Vbias 0.252372
R20855 Vbias.n380 Vbias 0.252372
R20856 Vbias.n382 Vbias 0.252372
R20857 Vbias.n322 Vbias 0.252372
R20858 Vbias.n324 Vbias 0.252372
R20859 Vbias.n326 Vbias 0.252372
R20860 Vbias.n328 Vbias 0.252372
R20861 Vbias.n330 Vbias 0.252372
R20862 Vbias.n332 Vbias 0.252372
R20863 Vbias.n334 Vbias 0.252372
R20864 Vbias.n336 Vbias 0.252372
R20865 Vbias.n338 Vbias 0.252372
R20866 Vbias.n340 Vbias 0.252372
R20867 Vbias.n342 Vbias 0.252372
R20868 Vbias.n344 Vbias 0.252372
R20869 Vbias.n346 Vbias 0.252372
R20870 Vbias.n348 Vbias 0.252372
R20871 Vbias.n350 Vbias 0.252372
R20872 Vbias.n290 Vbias 0.252372
R20873 Vbias.n292 Vbias 0.252372
R20874 Vbias.n294 Vbias 0.252372
R20875 Vbias.n296 Vbias 0.252372
R20876 Vbias.n298 Vbias 0.252372
R20877 Vbias.n300 Vbias 0.252372
R20878 Vbias.n302 Vbias 0.252372
R20879 Vbias.n304 Vbias 0.252372
R20880 Vbias.n306 Vbias 0.252372
R20881 Vbias.n308 Vbias 0.252372
R20882 Vbias.n310 Vbias 0.252372
R20883 Vbias.n312 Vbias 0.252372
R20884 Vbias.n314 Vbias 0.252372
R20885 Vbias.n316 Vbias 0.252372
R20886 Vbias.n318 Vbias 0.252372
R20887 Vbias.n258 Vbias 0.252372
R20888 Vbias.n260 Vbias 0.252372
R20889 Vbias.n262 Vbias 0.252372
R20890 Vbias.n264 Vbias 0.252372
R20891 Vbias.n266 Vbias 0.252372
R20892 Vbias.n268 Vbias 0.252372
R20893 Vbias.n270 Vbias 0.252372
R20894 Vbias.n272 Vbias 0.252372
R20895 Vbias.n274 Vbias 0.252372
R20896 Vbias.n276 Vbias 0.252372
R20897 Vbias.n278 Vbias 0.252372
R20898 Vbias.n280 Vbias 0.252372
R20899 Vbias.n282 Vbias 0.252372
R20900 Vbias.n284 Vbias 0.252372
R20901 Vbias.n286 Vbias 0.252372
R20902 Vbias.n226 Vbias 0.252372
R20903 Vbias.n228 Vbias 0.252372
R20904 Vbias.n230 Vbias 0.252372
R20905 Vbias.n232 Vbias 0.252372
R20906 Vbias.n234 Vbias 0.252372
R20907 Vbias.n236 Vbias 0.252372
R20908 Vbias.n238 Vbias 0.252372
R20909 Vbias.n240 Vbias 0.252372
R20910 Vbias.n242 Vbias 0.252372
R20911 Vbias.n244 Vbias 0.252372
R20912 Vbias.n246 Vbias 0.252372
R20913 Vbias.n248 Vbias 0.252372
R20914 Vbias.n250 Vbias 0.252372
R20915 Vbias.n252 Vbias 0.252372
R20916 Vbias.n254 Vbias 0.252372
R20917 Vbias.n194 Vbias 0.252372
R20918 Vbias.n196 Vbias 0.252372
R20919 Vbias.n198 Vbias 0.252372
R20920 Vbias.n200 Vbias 0.252372
R20921 Vbias.n202 Vbias 0.252372
R20922 Vbias.n204 Vbias 0.252372
R20923 Vbias.n206 Vbias 0.252372
R20924 Vbias.n208 Vbias 0.252372
R20925 Vbias.n210 Vbias 0.252372
R20926 Vbias.n212 Vbias 0.252372
R20927 Vbias.n214 Vbias 0.252372
R20928 Vbias.n216 Vbias 0.252372
R20929 Vbias.n218 Vbias 0.252372
R20930 Vbias.n220 Vbias 0.252372
R20931 Vbias.n222 Vbias 0.252372
R20932 Vbias.n162 Vbias 0.252372
R20933 Vbias.n164 Vbias 0.252372
R20934 Vbias.n166 Vbias 0.252372
R20935 Vbias.n168 Vbias 0.252372
R20936 Vbias.n170 Vbias 0.252372
R20937 Vbias.n172 Vbias 0.252372
R20938 Vbias.n174 Vbias 0.252372
R20939 Vbias.n176 Vbias 0.252372
R20940 Vbias.n178 Vbias 0.252372
R20941 Vbias.n180 Vbias 0.252372
R20942 Vbias.n182 Vbias 0.252372
R20943 Vbias.n184 Vbias 0.252372
R20944 Vbias.n186 Vbias 0.252372
R20945 Vbias.n188 Vbias 0.252372
R20946 Vbias.n190 Vbias 0.252372
R20947 Vbias.n130 Vbias 0.252372
R20948 Vbias.n132 Vbias 0.252372
R20949 Vbias.n134 Vbias 0.252372
R20950 Vbias.n136 Vbias 0.252372
R20951 Vbias.n138 Vbias 0.252372
R20952 Vbias.n140 Vbias 0.252372
R20953 Vbias.n142 Vbias 0.252372
R20954 Vbias.n144 Vbias 0.252372
R20955 Vbias.n146 Vbias 0.252372
R20956 Vbias.n148 Vbias 0.252372
R20957 Vbias.n150 Vbias 0.252372
R20958 Vbias.n152 Vbias 0.252372
R20959 Vbias.n154 Vbias 0.252372
R20960 Vbias.n156 Vbias 0.252372
R20961 Vbias.n158 Vbias 0.252372
R20962 Vbias.n98 Vbias 0.252372
R20963 Vbias.n100 Vbias 0.252372
R20964 Vbias.n102 Vbias 0.252372
R20965 Vbias.n104 Vbias 0.252372
R20966 Vbias.n106 Vbias 0.252372
R20967 Vbias.n108 Vbias 0.252372
R20968 Vbias.n110 Vbias 0.252372
R20969 Vbias.n112 Vbias 0.252372
R20970 Vbias.n114 Vbias 0.252372
R20971 Vbias.n116 Vbias 0.252372
R20972 Vbias.n118 Vbias 0.252372
R20973 Vbias.n120 Vbias 0.252372
R20974 Vbias.n122 Vbias 0.252372
R20975 Vbias.n124 Vbias 0.252372
R20976 Vbias.n126 Vbias 0.252372
R20977 Vbias.n66 Vbias 0.252372
R20978 Vbias.n68 Vbias 0.252372
R20979 Vbias.n70 Vbias 0.252372
R20980 Vbias.n72 Vbias 0.252372
R20981 Vbias.n74 Vbias 0.252372
R20982 Vbias.n76 Vbias 0.252372
R20983 Vbias.n78 Vbias 0.252372
R20984 Vbias.n80 Vbias 0.252372
R20985 Vbias.n82 Vbias 0.252372
R20986 Vbias.n84 Vbias 0.252372
R20987 Vbias.n86 Vbias 0.252372
R20988 Vbias.n88 Vbias 0.252372
R20989 Vbias.n90 Vbias 0.252372
R20990 Vbias.n92 Vbias 0.252372
R20991 Vbias.n94 Vbias 0.252372
R20992 Vbias.n34 Vbias 0.252372
R20993 Vbias.n36 Vbias 0.252372
R20994 Vbias.n38 Vbias 0.252372
R20995 Vbias.n40 Vbias 0.252372
R20996 Vbias.n42 Vbias 0.252372
R20997 Vbias.n44 Vbias 0.252372
R20998 Vbias.n46 Vbias 0.252372
R20999 Vbias.n48 Vbias 0.252372
R21000 Vbias.n50 Vbias 0.252372
R21001 Vbias.n52 Vbias 0.252372
R21002 Vbias.n54 Vbias 0.252372
R21003 Vbias.n56 Vbias 0.252372
R21004 Vbias.n58 Vbias 0.252372
R21005 Vbias.n60 Vbias 0.252372
R21006 Vbias.n62 Vbias 0.252372
R21007 Vbias.n2 Vbias 0.252372
R21008 Vbias.n4 Vbias 0.252372
R21009 Vbias.n6 Vbias 0.252372
R21010 Vbias.n8 Vbias 0.252372
R21011 Vbias.n10 Vbias 0.252372
R21012 Vbias.n12 Vbias 0.252372
R21013 Vbias.n14 Vbias 0.252372
R21014 Vbias.n16 Vbias 0.252372
R21015 Vbias.n18 Vbias 0.252372
R21016 Vbias.n20 Vbias 0.252372
R21017 Vbias.n22 Vbias 0.252372
R21018 Vbias.n24 Vbias 0.252372
R21019 Vbias.n26 Vbias 0.252372
R21020 Vbias.n28 Vbias 0.252372
R21021 Vbias.n30 Vbias 0.252372
R21022 Vbias Vbias.n517 0.237067
R21023 Vbias Vbias.n482 0.0972718
R21024 Vbias Vbias.n484 0.0972718
R21025 Vbias Vbias.n486 0.0972718
R21026 Vbias Vbias.n488 0.0972718
R21027 Vbias Vbias.n490 0.0972718
R21028 Vbias Vbias.n492 0.0972718
R21029 Vbias Vbias.n494 0.0972718
R21030 Vbias Vbias.n496 0.0972718
R21031 Vbias Vbias.n498 0.0972718
R21032 Vbias Vbias.n500 0.0972718
R21033 Vbias Vbias.n502 0.0972718
R21034 Vbias Vbias.n504 0.0972718
R21035 Vbias Vbias.n506 0.0972718
R21036 Vbias Vbias.n508 0.0972718
R21037 Vbias Vbias.n510 0.0972718
R21038 Vbias Vbias.n450 0.0972718
R21039 Vbias Vbias.n452 0.0972718
R21040 Vbias Vbias.n454 0.0972718
R21041 Vbias Vbias.n456 0.0972718
R21042 Vbias Vbias.n458 0.0972718
R21043 Vbias Vbias.n460 0.0972718
R21044 Vbias Vbias.n462 0.0972718
R21045 Vbias Vbias.n464 0.0972718
R21046 Vbias Vbias.n466 0.0972718
R21047 Vbias Vbias.n468 0.0972718
R21048 Vbias Vbias.n470 0.0972718
R21049 Vbias Vbias.n472 0.0972718
R21050 Vbias Vbias.n474 0.0972718
R21051 Vbias Vbias.n476 0.0972718
R21052 Vbias Vbias.n478 0.0972718
R21053 Vbias Vbias.n418 0.0972718
R21054 Vbias Vbias.n420 0.0972718
R21055 Vbias Vbias.n422 0.0972718
R21056 Vbias Vbias.n424 0.0972718
R21057 Vbias Vbias.n426 0.0972718
R21058 Vbias Vbias.n428 0.0972718
R21059 Vbias Vbias.n430 0.0972718
R21060 Vbias Vbias.n432 0.0972718
R21061 Vbias Vbias.n434 0.0972718
R21062 Vbias Vbias.n436 0.0972718
R21063 Vbias Vbias.n438 0.0972718
R21064 Vbias Vbias.n440 0.0972718
R21065 Vbias Vbias.n442 0.0972718
R21066 Vbias Vbias.n444 0.0972718
R21067 Vbias Vbias.n446 0.0972718
R21068 Vbias Vbias.n386 0.0972718
R21069 Vbias Vbias.n388 0.0972718
R21070 Vbias Vbias.n390 0.0972718
R21071 Vbias Vbias.n392 0.0972718
R21072 Vbias Vbias.n394 0.0972718
R21073 Vbias Vbias.n396 0.0972718
R21074 Vbias Vbias.n398 0.0972718
R21075 Vbias Vbias.n400 0.0972718
R21076 Vbias Vbias.n402 0.0972718
R21077 Vbias Vbias.n404 0.0972718
R21078 Vbias Vbias.n406 0.0972718
R21079 Vbias Vbias.n408 0.0972718
R21080 Vbias Vbias.n410 0.0972718
R21081 Vbias Vbias.n412 0.0972718
R21082 Vbias Vbias.n414 0.0972718
R21083 Vbias Vbias.n354 0.0972718
R21084 Vbias Vbias.n356 0.0972718
R21085 Vbias Vbias.n358 0.0972718
R21086 Vbias Vbias.n360 0.0972718
R21087 Vbias Vbias.n362 0.0972718
R21088 Vbias Vbias.n364 0.0972718
R21089 Vbias Vbias.n366 0.0972718
R21090 Vbias Vbias.n368 0.0972718
R21091 Vbias Vbias.n370 0.0972718
R21092 Vbias Vbias.n372 0.0972718
R21093 Vbias Vbias.n374 0.0972718
R21094 Vbias Vbias.n376 0.0972718
R21095 Vbias Vbias.n378 0.0972718
R21096 Vbias Vbias.n380 0.0972718
R21097 Vbias Vbias.n382 0.0972718
R21098 Vbias Vbias.n322 0.0972718
R21099 Vbias Vbias.n324 0.0972718
R21100 Vbias Vbias.n326 0.0972718
R21101 Vbias Vbias.n328 0.0972718
R21102 Vbias Vbias.n330 0.0972718
R21103 Vbias Vbias.n332 0.0972718
R21104 Vbias Vbias.n334 0.0972718
R21105 Vbias Vbias.n336 0.0972718
R21106 Vbias Vbias.n338 0.0972718
R21107 Vbias Vbias.n340 0.0972718
R21108 Vbias Vbias.n342 0.0972718
R21109 Vbias Vbias.n344 0.0972718
R21110 Vbias Vbias.n346 0.0972718
R21111 Vbias Vbias.n348 0.0972718
R21112 Vbias Vbias.n350 0.0972718
R21113 Vbias Vbias.n290 0.0972718
R21114 Vbias Vbias.n292 0.0972718
R21115 Vbias Vbias.n294 0.0972718
R21116 Vbias Vbias.n296 0.0972718
R21117 Vbias Vbias.n298 0.0972718
R21118 Vbias Vbias.n300 0.0972718
R21119 Vbias Vbias.n302 0.0972718
R21120 Vbias Vbias.n304 0.0972718
R21121 Vbias Vbias.n306 0.0972718
R21122 Vbias Vbias.n308 0.0972718
R21123 Vbias Vbias.n310 0.0972718
R21124 Vbias Vbias.n312 0.0972718
R21125 Vbias Vbias.n314 0.0972718
R21126 Vbias Vbias.n316 0.0972718
R21127 Vbias Vbias.n318 0.0972718
R21128 Vbias Vbias.n258 0.0972718
R21129 Vbias Vbias.n260 0.0972718
R21130 Vbias Vbias.n262 0.0972718
R21131 Vbias Vbias.n264 0.0972718
R21132 Vbias Vbias.n266 0.0972718
R21133 Vbias Vbias.n268 0.0972718
R21134 Vbias Vbias.n270 0.0972718
R21135 Vbias Vbias.n272 0.0972718
R21136 Vbias Vbias.n274 0.0972718
R21137 Vbias Vbias.n276 0.0972718
R21138 Vbias Vbias.n278 0.0972718
R21139 Vbias Vbias.n280 0.0972718
R21140 Vbias Vbias.n282 0.0972718
R21141 Vbias Vbias.n284 0.0972718
R21142 Vbias Vbias.n286 0.0972718
R21143 Vbias Vbias.n226 0.0972718
R21144 Vbias Vbias.n228 0.0972718
R21145 Vbias Vbias.n230 0.0972718
R21146 Vbias Vbias.n232 0.0972718
R21147 Vbias Vbias.n234 0.0972718
R21148 Vbias Vbias.n236 0.0972718
R21149 Vbias Vbias.n238 0.0972718
R21150 Vbias Vbias.n240 0.0972718
R21151 Vbias Vbias.n242 0.0972718
R21152 Vbias Vbias.n244 0.0972718
R21153 Vbias Vbias.n246 0.0972718
R21154 Vbias Vbias.n248 0.0972718
R21155 Vbias Vbias.n250 0.0972718
R21156 Vbias Vbias.n252 0.0972718
R21157 Vbias Vbias.n254 0.0972718
R21158 Vbias Vbias.n194 0.0972718
R21159 Vbias Vbias.n196 0.0972718
R21160 Vbias Vbias.n198 0.0972718
R21161 Vbias Vbias.n200 0.0972718
R21162 Vbias Vbias.n202 0.0972718
R21163 Vbias Vbias.n204 0.0972718
R21164 Vbias Vbias.n206 0.0972718
R21165 Vbias Vbias.n208 0.0972718
R21166 Vbias Vbias.n210 0.0972718
R21167 Vbias Vbias.n212 0.0972718
R21168 Vbias Vbias.n214 0.0972718
R21169 Vbias Vbias.n216 0.0972718
R21170 Vbias Vbias.n218 0.0972718
R21171 Vbias Vbias.n220 0.0972718
R21172 Vbias Vbias.n222 0.0972718
R21173 Vbias Vbias.n162 0.0972718
R21174 Vbias Vbias.n164 0.0972718
R21175 Vbias Vbias.n166 0.0972718
R21176 Vbias Vbias.n168 0.0972718
R21177 Vbias Vbias.n170 0.0972718
R21178 Vbias Vbias.n172 0.0972718
R21179 Vbias Vbias.n174 0.0972718
R21180 Vbias Vbias.n176 0.0972718
R21181 Vbias Vbias.n178 0.0972718
R21182 Vbias Vbias.n180 0.0972718
R21183 Vbias Vbias.n182 0.0972718
R21184 Vbias Vbias.n184 0.0972718
R21185 Vbias Vbias.n186 0.0972718
R21186 Vbias Vbias.n188 0.0972718
R21187 Vbias Vbias.n190 0.0972718
R21188 Vbias Vbias.n130 0.0972718
R21189 Vbias Vbias.n132 0.0972718
R21190 Vbias Vbias.n134 0.0972718
R21191 Vbias Vbias.n136 0.0972718
R21192 Vbias Vbias.n138 0.0972718
R21193 Vbias Vbias.n140 0.0972718
R21194 Vbias Vbias.n142 0.0972718
R21195 Vbias Vbias.n144 0.0972718
R21196 Vbias Vbias.n146 0.0972718
R21197 Vbias Vbias.n148 0.0972718
R21198 Vbias Vbias.n150 0.0972718
R21199 Vbias Vbias.n152 0.0972718
R21200 Vbias Vbias.n154 0.0972718
R21201 Vbias Vbias.n156 0.0972718
R21202 Vbias Vbias.n158 0.0972718
R21203 Vbias Vbias.n98 0.0972718
R21204 Vbias Vbias.n100 0.0972718
R21205 Vbias Vbias.n102 0.0972718
R21206 Vbias Vbias.n104 0.0972718
R21207 Vbias Vbias.n106 0.0972718
R21208 Vbias Vbias.n108 0.0972718
R21209 Vbias Vbias.n110 0.0972718
R21210 Vbias Vbias.n112 0.0972718
R21211 Vbias Vbias.n114 0.0972718
R21212 Vbias Vbias.n116 0.0972718
R21213 Vbias Vbias.n118 0.0972718
R21214 Vbias Vbias.n120 0.0972718
R21215 Vbias Vbias.n122 0.0972718
R21216 Vbias Vbias.n124 0.0972718
R21217 Vbias Vbias.n126 0.0972718
R21218 Vbias Vbias.n66 0.0972718
R21219 Vbias Vbias.n68 0.0972718
R21220 Vbias Vbias.n70 0.0972718
R21221 Vbias Vbias.n72 0.0972718
R21222 Vbias Vbias.n74 0.0972718
R21223 Vbias Vbias.n76 0.0972718
R21224 Vbias Vbias.n78 0.0972718
R21225 Vbias Vbias.n80 0.0972718
R21226 Vbias Vbias.n82 0.0972718
R21227 Vbias Vbias.n84 0.0972718
R21228 Vbias Vbias.n86 0.0972718
R21229 Vbias Vbias.n88 0.0972718
R21230 Vbias Vbias.n90 0.0972718
R21231 Vbias Vbias.n92 0.0972718
R21232 Vbias Vbias.n94 0.0972718
R21233 Vbias Vbias.n34 0.0972718
R21234 Vbias Vbias.n36 0.0972718
R21235 Vbias Vbias.n38 0.0972718
R21236 Vbias Vbias.n40 0.0972718
R21237 Vbias Vbias.n42 0.0972718
R21238 Vbias Vbias.n44 0.0972718
R21239 Vbias Vbias.n46 0.0972718
R21240 Vbias Vbias.n48 0.0972718
R21241 Vbias Vbias.n50 0.0972718
R21242 Vbias Vbias.n52 0.0972718
R21243 Vbias Vbias.n54 0.0972718
R21244 Vbias Vbias.n56 0.0972718
R21245 Vbias Vbias.n58 0.0972718
R21246 Vbias Vbias.n60 0.0972718
R21247 Vbias Vbias.n62 0.0972718
R21248 Vbias Vbias.n2 0.0972718
R21249 Vbias Vbias.n4 0.0972718
R21250 Vbias Vbias.n6 0.0972718
R21251 Vbias Vbias.n8 0.0972718
R21252 Vbias Vbias.n10 0.0972718
R21253 Vbias Vbias.n12 0.0972718
R21254 Vbias Vbias.n14 0.0972718
R21255 Vbias Vbias.n16 0.0972718
R21256 Vbias Vbias.n18 0.0972718
R21257 Vbias Vbias.n20 0.0972718
R21258 Vbias Vbias.n22 0.0972718
R21259 Vbias Vbias.n24 0.0972718
R21260 Vbias Vbias.n26 0.0972718
R21261 Vbias Vbias.n28 0.0972718
R21262 Vbias Vbias.n30 0.0972718
R21263 Vbias.n509 Vbias 0.0489375
R21264 Vbias.n507 Vbias 0.0489375
R21265 Vbias.n505 Vbias 0.0489375
R21266 Vbias.n503 Vbias 0.0489375
R21267 Vbias.n501 Vbias 0.0489375
R21268 Vbias.n499 Vbias 0.0489375
R21269 Vbias.n497 Vbias 0.0489375
R21270 Vbias.n495 Vbias 0.0489375
R21271 Vbias.n493 Vbias 0.0489375
R21272 Vbias.n491 Vbias 0.0489375
R21273 Vbias.n489 Vbias 0.0489375
R21274 Vbias.n487 Vbias 0.0489375
R21275 Vbias.n485 Vbias 0.0489375
R21276 Vbias.n483 Vbias 0.0489375
R21277 Vbias.n481 Vbias 0.0489375
R21278 Vbias.n480 Vbias 0.0489375
R21279 Vbias.n477 Vbias 0.0489375
R21280 Vbias.n475 Vbias 0.0489375
R21281 Vbias.n473 Vbias 0.0489375
R21282 Vbias.n471 Vbias 0.0489375
R21283 Vbias.n469 Vbias 0.0489375
R21284 Vbias.n467 Vbias 0.0489375
R21285 Vbias.n465 Vbias 0.0489375
R21286 Vbias.n463 Vbias 0.0489375
R21287 Vbias.n461 Vbias 0.0489375
R21288 Vbias.n459 Vbias 0.0489375
R21289 Vbias.n457 Vbias 0.0489375
R21290 Vbias.n455 Vbias 0.0489375
R21291 Vbias.n453 Vbias 0.0489375
R21292 Vbias.n451 Vbias 0.0489375
R21293 Vbias.n449 Vbias 0.0489375
R21294 Vbias.n448 Vbias 0.0489375
R21295 Vbias.n445 Vbias 0.0489375
R21296 Vbias.n443 Vbias 0.0489375
R21297 Vbias.n441 Vbias 0.0489375
R21298 Vbias.n439 Vbias 0.0489375
R21299 Vbias.n437 Vbias 0.0489375
R21300 Vbias.n435 Vbias 0.0489375
R21301 Vbias.n433 Vbias 0.0489375
R21302 Vbias.n431 Vbias 0.0489375
R21303 Vbias.n429 Vbias 0.0489375
R21304 Vbias.n427 Vbias 0.0489375
R21305 Vbias.n425 Vbias 0.0489375
R21306 Vbias.n423 Vbias 0.0489375
R21307 Vbias.n421 Vbias 0.0489375
R21308 Vbias.n419 Vbias 0.0489375
R21309 Vbias.n417 Vbias 0.0489375
R21310 Vbias.n416 Vbias 0.0489375
R21311 Vbias.n413 Vbias 0.0489375
R21312 Vbias.n411 Vbias 0.0489375
R21313 Vbias.n409 Vbias 0.0489375
R21314 Vbias.n407 Vbias 0.0489375
R21315 Vbias.n405 Vbias 0.0489375
R21316 Vbias.n403 Vbias 0.0489375
R21317 Vbias.n401 Vbias 0.0489375
R21318 Vbias.n399 Vbias 0.0489375
R21319 Vbias.n397 Vbias 0.0489375
R21320 Vbias.n395 Vbias 0.0489375
R21321 Vbias.n393 Vbias 0.0489375
R21322 Vbias.n391 Vbias 0.0489375
R21323 Vbias.n389 Vbias 0.0489375
R21324 Vbias.n387 Vbias 0.0489375
R21325 Vbias.n385 Vbias 0.0489375
R21326 Vbias.n384 Vbias 0.0489375
R21327 Vbias.n381 Vbias 0.0489375
R21328 Vbias.n379 Vbias 0.0489375
R21329 Vbias.n377 Vbias 0.0489375
R21330 Vbias.n375 Vbias 0.0489375
R21331 Vbias.n373 Vbias 0.0489375
R21332 Vbias.n371 Vbias 0.0489375
R21333 Vbias.n369 Vbias 0.0489375
R21334 Vbias.n367 Vbias 0.0489375
R21335 Vbias.n365 Vbias 0.0489375
R21336 Vbias.n363 Vbias 0.0489375
R21337 Vbias.n361 Vbias 0.0489375
R21338 Vbias.n359 Vbias 0.0489375
R21339 Vbias.n357 Vbias 0.0489375
R21340 Vbias.n355 Vbias 0.0489375
R21341 Vbias.n353 Vbias 0.0489375
R21342 Vbias.n352 Vbias 0.0489375
R21343 Vbias.n349 Vbias 0.0489375
R21344 Vbias.n347 Vbias 0.0489375
R21345 Vbias.n345 Vbias 0.0489375
R21346 Vbias.n343 Vbias 0.0489375
R21347 Vbias.n341 Vbias 0.0489375
R21348 Vbias.n339 Vbias 0.0489375
R21349 Vbias.n337 Vbias 0.0489375
R21350 Vbias.n335 Vbias 0.0489375
R21351 Vbias.n333 Vbias 0.0489375
R21352 Vbias.n331 Vbias 0.0489375
R21353 Vbias.n329 Vbias 0.0489375
R21354 Vbias.n327 Vbias 0.0489375
R21355 Vbias.n325 Vbias 0.0489375
R21356 Vbias.n323 Vbias 0.0489375
R21357 Vbias.n321 Vbias 0.0489375
R21358 Vbias.n320 Vbias 0.0489375
R21359 Vbias.n317 Vbias 0.0489375
R21360 Vbias.n315 Vbias 0.0489375
R21361 Vbias.n313 Vbias 0.0489375
R21362 Vbias.n311 Vbias 0.0489375
R21363 Vbias.n309 Vbias 0.0489375
R21364 Vbias.n307 Vbias 0.0489375
R21365 Vbias.n305 Vbias 0.0489375
R21366 Vbias.n303 Vbias 0.0489375
R21367 Vbias.n301 Vbias 0.0489375
R21368 Vbias.n299 Vbias 0.0489375
R21369 Vbias.n297 Vbias 0.0489375
R21370 Vbias.n295 Vbias 0.0489375
R21371 Vbias.n293 Vbias 0.0489375
R21372 Vbias.n291 Vbias 0.0489375
R21373 Vbias.n289 Vbias 0.0489375
R21374 Vbias.n288 Vbias 0.0489375
R21375 Vbias.n285 Vbias 0.0489375
R21376 Vbias.n283 Vbias 0.0489375
R21377 Vbias.n281 Vbias 0.0489375
R21378 Vbias.n279 Vbias 0.0489375
R21379 Vbias.n277 Vbias 0.0489375
R21380 Vbias.n275 Vbias 0.0489375
R21381 Vbias.n273 Vbias 0.0489375
R21382 Vbias.n271 Vbias 0.0489375
R21383 Vbias.n269 Vbias 0.0489375
R21384 Vbias.n267 Vbias 0.0489375
R21385 Vbias.n265 Vbias 0.0489375
R21386 Vbias.n263 Vbias 0.0489375
R21387 Vbias.n261 Vbias 0.0489375
R21388 Vbias.n259 Vbias 0.0489375
R21389 Vbias.n257 Vbias 0.0489375
R21390 Vbias.n256 Vbias 0.0489375
R21391 Vbias.n253 Vbias 0.0489375
R21392 Vbias.n251 Vbias 0.0489375
R21393 Vbias.n249 Vbias 0.0489375
R21394 Vbias.n247 Vbias 0.0489375
R21395 Vbias.n245 Vbias 0.0489375
R21396 Vbias.n243 Vbias 0.0489375
R21397 Vbias.n241 Vbias 0.0489375
R21398 Vbias.n239 Vbias 0.0489375
R21399 Vbias.n237 Vbias 0.0489375
R21400 Vbias.n235 Vbias 0.0489375
R21401 Vbias.n233 Vbias 0.0489375
R21402 Vbias.n231 Vbias 0.0489375
R21403 Vbias.n229 Vbias 0.0489375
R21404 Vbias.n227 Vbias 0.0489375
R21405 Vbias.n225 Vbias 0.0489375
R21406 Vbias.n224 Vbias 0.0489375
R21407 Vbias.n221 Vbias 0.0489375
R21408 Vbias.n219 Vbias 0.0489375
R21409 Vbias.n217 Vbias 0.0489375
R21410 Vbias.n215 Vbias 0.0489375
R21411 Vbias.n213 Vbias 0.0489375
R21412 Vbias.n211 Vbias 0.0489375
R21413 Vbias.n209 Vbias 0.0489375
R21414 Vbias.n207 Vbias 0.0489375
R21415 Vbias.n205 Vbias 0.0489375
R21416 Vbias.n203 Vbias 0.0489375
R21417 Vbias.n201 Vbias 0.0489375
R21418 Vbias.n199 Vbias 0.0489375
R21419 Vbias.n197 Vbias 0.0489375
R21420 Vbias.n195 Vbias 0.0489375
R21421 Vbias.n193 Vbias 0.0489375
R21422 Vbias.n192 Vbias 0.0489375
R21423 Vbias.n189 Vbias 0.0489375
R21424 Vbias.n187 Vbias 0.0489375
R21425 Vbias.n185 Vbias 0.0489375
R21426 Vbias.n183 Vbias 0.0489375
R21427 Vbias.n181 Vbias 0.0489375
R21428 Vbias.n179 Vbias 0.0489375
R21429 Vbias.n177 Vbias 0.0489375
R21430 Vbias.n175 Vbias 0.0489375
R21431 Vbias.n173 Vbias 0.0489375
R21432 Vbias.n171 Vbias 0.0489375
R21433 Vbias.n169 Vbias 0.0489375
R21434 Vbias.n167 Vbias 0.0489375
R21435 Vbias.n165 Vbias 0.0489375
R21436 Vbias.n163 Vbias 0.0489375
R21437 Vbias.n161 Vbias 0.0489375
R21438 Vbias.n160 Vbias 0.0489375
R21439 Vbias.n157 Vbias 0.0489375
R21440 Vbias.n155 Vbias 0.0489375
R21441 Vbias.n153 Vbias 0.0489375
R21442 Vbias.n151 Vbias 0.0489375
R21443 Vbias.n149 Vbias 0.0489375
R21444 Vbias.n147 Vbias 0.0489375
R21445 Vbias.n145 Vbias 0.0489375
R21446 Vbias.n143 Vbias 0.0489375
R21447 Vbias.n141 Vbias 0.0489375
R21448 Vbias.n139 Vbias 0.0489375
R21449 Vbias.n137 Vbias 0.0489375
R21450 Vbias.n135 Vbias 0.0489375
R21451 Vbias.n133 Vbias 0.0489375
R21452 Vbias.n131 Vbias 0.0489375
R21453 Vbias.n129 Vbias 0.0489375
R21454 Vbias.n128 Vbias 0.0489375
R21455 Vbias.n125 Vbias 0.0489375
R21456 Vbias.n123 Vbias 0.0489375
R21457 Vbias.n121 Vbias 0.0489375
R21458 Vbias.n119 Vbias 0.0489375
R21459 Vbias.n117 Vbias 0.0489375
R21460 Vbias.n115 Vbias 0.0489375
R21461 Vbias.n113 Vbias 0.0489375
R21462 Vbias.n111 Vbias 0.0489375
R21463 Vbias.n109 Vbias 0.0489375
R21464 Vbias.n107 Vbias 0.0489375
R21465 Vbias.n105 Vbias 0.0489375
R21466 Vbias.n103 Vbias 0.0489375
R21467 Vbias.n101 Vbias 0.0489375
R21468 Vbias.n99 Vbias 0.0489375
R21469 Vbias.n97 Vbias 0.0489375
R21470 Vbias.n96 Vbias 0.0489375
R21471 Vbias.n93 Vbias 0.0489375
R21472 Vbias.n91 Vbias 0.0489375
R21473 Vbias.n89 Vbias 0.0489375
R21474 Vbias.n87 Vbias 0.0489375
R21475 Vbias.n85 Vbias 0.0489375
R21476 Vbias.n83 Vbias 0.0489375
R21477 Vbias.n81 Vbias 0.0489375
R21478 Vbias.n79 Vbias 0.0489375
R21479 Vbias.n77 Vbias 0.0489375
R21480 Vbias.n75 Vbias 0.0489375
R21481 Vbias.n73 Vbias 0.0489375
R21482 Vbias.n71 Vbias 0.0489375
R21483 Vbias.n69 Vbias 0.0489375
R21484 Vbias.n67 Vbias 0.0489375
R21485 Vbias.n65 Vbias 0.0489375
R21486 Vbias.n64 Vbias 0.0489375
R21487 Vbias.n61 Vbias 0.0489375
R21488 Vbias.n59 Vbias 0.0489375
R21489 Vbias.n57 Vbias 0.0489375
R21490 Vbias.n55 Vbias 0.0489375
R21491 Vbias.n53 Vbias 0.0489375
R21492 Vbias.n51 Vbias 0.0489375
R21493 Vbias.n49 Vbias 0.0489375
R21494 Vbias.n47 Vbias 0.0489375
R21495 Vbias.n45 Vbias 0.0489375
R21496 Vbias.n43 Vbias 0.0489375
R21497 Vbias.n41 Vbias 0.0489375
R21498 Vbias.n39 Vbias 0.0489375
R21499 Vbias.n37 Vbias 0.0489375
R21500 Vbias.n35 Vbias 0.0489375
R21501 Vbias.n33 Vbias 0.0489375
R21502 Vbias.n32 Vbias 0.0489375
R21503 Vbias.n29 Vbias 0.0489375
R21504 Vbias.n27 Vbias 0.0489375
R21505 Vbias.n25 Vbias 0.0489375
R21506 Vbias.n23 Vbias 0.0489375
R21507 Vbias.n21 Vbias 0.0489375
R21508 Vbias.n19 Vbias 0.0489375
R21509 Vbias.n17 Vbias 0.0489375
R21510 Vbias.n15 Vbias 0.0489375
R21511 Vbias.n13 Vbias 0.0489375
R21512 Vbias.n11 Vbias 0.0489375
R21513 Vbias.n9 Vbias 0.0489375
R21514 Vbias.n7 Vbias 0.0489375
R21515 Vbias.n5 Vbias 0.0489375
R21516 Vbias.n3 Vbias 0.0489375
R21517 Vbias.n1 Vbias 0.0489375
R21518 Vbias.n0 Vbias 0.0489375
R21519 XThC.Tn[1].n2 XThC.Tn[1].n1 332.332
R21520 XThC.Tn[1].n2 XThC.Tn[1].n0 296.493
R21521 XThC.Tn[1].n12 XThC.Tn[1].n10 161.406
R21522 XThC.Tn[1].n15 XThC.Tn[1].n13 161.406
R21523 XThC.Tn[1].n18 XThC.Tn[1].n16 161.406
R21524 XThC.Tn[1].n21 XThC.Tn[1].n19 161.406
R21525 XThC.Tn[1].n24 XThC.Tn[1].n22 161.406
R21526 XThC.Tn[1].n27 XThC.Tn[1].n25 161.406
R21527 XThC.Tn[1].n30 XThC.Tn[1].n28 161.406
R21528 XThC.Tn[1].n33 XThC.Tn[1].n31 161.406
R21529 XThC.Tn[1].n36 XThC.Tn[1].n34 161.406
R21530 XThC.Tn[1].n39 XThC.Tn[1].n37 161.406
R21531 XThC.Tn[1].n42 XThC.Tn[1].n40 161.406
R21532 XThC.Tn[1].n45 XThC.Tn[1].n43 161.406
R21533 XThC.Tn[1].n48 XThC.Tn[1].n46 161.406
R21534 XThC.Tn[1].n51 XThC.Tn[1].n49 161.406
R21535 XThC.Tn[1].n54 XThC.Tn[1].n52 161.406
R21536 XThC.Tn[1].n57 XThC.Tn[1].n55 161.406
R21537 XThC.Tn[1].n10 XThC.Tn[1].t29 161.202
R21538 XThC.Tn[1].n13 XThC.Tn[1].t14 161.202
R21539 XThC.Tn[1].n16 XThC.Tn[1].t16 161.202
R21540 XThC.Tn[1].n19 XThC.Tn[1].t18 161.202
R21541 XThC.Tn[1].n22 XThC.Tn[1].t39 161.202
R21542 XThC.Tn[1].n25 XThC.Tn[1].t40 161.202
R21543 XThC.Tn[1].n28 XThC.Tn[1].t21 161.202
R21544 XThC.Tn[1].n31 XThC.Tn[1].t30 161.202
R21545 XThC.Tn[1].n34 XThC.Tn[1].t32 161.202
R21546 XThC.Tn[1].n37 XThC.Tn[1].t19 161.202
R21547 XThC.Tn[1].n40 XThC.Tn[1].t20 161.202
R21548 XThC.Tn[1].n43 XThC.Tn[1].t33 161.202
R21549 XThC.Tn[1].n46 XThC.Tn[1].t41 161.202
R21550 XThC.Tn[1].n49 XThC.Tn[1].t12 161.202
R21551 XThC.Tn[1].n52 XThC.Tn[1].t25 161.202
R21552 XThC.Tn[1].n55 XThC.Tn[1].t35 161.202
R21553 XThC.Tn[1].n10 XThC.Tn[1].t31 145.137
R21554 XThC.Tn[1].n13 XThC.Tn[1].t17 145.137
R21555 XThC.Tn[1].n16 XThC.Tn[1].t22 145.137
R21556 XThC.Tn[1].n19 XThC.Tn[1].t23 145.137
R21557 XThC.Tn[1].n22 XThC.Tn[1].t42 145.137
R21558 XThC.Tn[1].n25 XThC.Tn[1].t43 145.137
R21559 XThC.Tn[1].n28 XThC.Tn[1].t27 145.137
R21560 XThC.Tn[1].n31 XThC.Tn[1].t34 145.137
R21561 XThC.Tn[1].n34 XThC.Tn[1].t36 145.137
R21562 XThC.Tn[1].n37 XThC.Tn[1].t24 145.137
R21563 XThC.Tn[1].n40 XThC.Tn[1].t26 145.137
R21564 XThC.Tn[1].n43 XThC.Tn[1].t37 145.137
R21565 XThC.Tn[1].n46 XThC.Tn[1].t13 145.137
R21566 XThC.Tn[1].n49 XThC.Tn[1].t15 145.137
R21567 XThC.Tn[1].n52 XThC.Tn[1].t28 145.137
R21568 XThC.Tn[1].n55 XThC.Tn[1].t38 145.137
R21569 XThC.Tn[1].n7 XThC.Tn[1].n6 135.249
R21570 XThC.Tn[1].n9 XThC.Tn[1].n3 98.981
R21571 XThC.Tn[1].n8 XThC.Tn[1].n4 98.981
R21572 XThC.Tn[1].n7 XThC.Tn[1].n5 98.981
R21573 XThC.Tn[1].n9 XThC.Tn[1].n8 36.2672
R21574 XThC.Tn[1].n8 XThC.Tn[1].n7 36.2672
R21575 XThC.Tn[1].n59 XThC.Tn[1].n9 32.6405
R21576 XThC.Tn[1].n1 XThC.Tn[1].t5 26.5955
R21577 XThC.Tn[1].n1 XThC.Tn[1].t4 26.5955
R21578 XThC.Tn[1].n0 XThC.Tn[1].t7 26.5955
R21579 XThC.Tn[1].n0 XThC.Tn[1].t6 26.5955
R21580 XThC.Tn[1].n3 XThC.Tn[1].t9 24.9236
R21581 XThC.Tn[1].n3 XThC.Tn[1].t8 24.9236
R21582 XThC.Tn[1].n4 XThC.Tn[1].t11 24.9236
R21583 XThC.Tn[1].n4 XThC.Tn[1].t10 24.9236
R21584 XThC.Tn[1].n5 XThC.Tn[1].t1 24.9236
R21585 XThC.Tn[1].n5 XThC.Tn[1].t0 24.9236
R21586 XThC.Tn[1].n6 XThC.Tn[1].t3 24.9236
R21587 XThC.Tn[1].n6 XThC.Tn[1].t2 24.9236
R21588 XThC.Tn[1] XThC.Tn[1].n2 23.3605
R21589 XThC.Tn[1].n58 XThC.Tn[1] 7.29217
R21590 XThC.Tn[1] XThC.Tn[1].n59 6.7205
R21591 XThC.Tn[1].n59 XThC.Tn[1].n58 3.13711
R21592 XThC.Tn[1].n15 XThC.Tn[1] 0.931056
R21593 XThC.Tn[1].n18 XThC.Tn[1] 0.931056
R21594 XThC.Tn[1].n21 XThC.Tn[1] 0.931056
R21595 XThC.Tn[1].n24 XThC.Tn[1] 0.931056
R21596 XThC.Tn[1].n27 XThC.Tn[1] 0.931056
R21597 XThC.Tn[1].n30 XThC.Tn[1] 0.931056
R21598 XThC.Tn[1].n33 XThC.Tn[1] 0.931056
R21599 XThC.Tn[1].n36 XThC.Tn[1] 0.931056
R21600 XThC.Tn[1].n39 XThC.Tn[1] 0.931056
R21601 XThC.Tn[1].n42 XThC.Tn[1] 0.931056
R21602 XThC.Tn[1].n45 XThC.Tn[1] 0.931056
R21603 XThC.Tn[1].n48 XThC.Tn[1] 0.931056
R21604 XThC.Tn[1].n51 XThC.Tn[1] 0.931056
R21605 XThC.Tn[1].n54 XThC.Tn[1] 0.931056
R21606 XThC.Tn[1].n57 XThC.Tn[1] 0.931056
R21607 XThC.Tn[1] XThC.Tn[1].n12 0.396333
R21608 XThC.Tn[1] XThC.Tn[1].n15 0.396333
R21609 XThC.Tn[1] XThC.Tn[1].n18 0.396333
R21610 XThC.Tn[1] XThC.Tn[1].n21 0.396333
R21611 XThC.Tn[1] XThC.Tn[1].n24 0.396333
R21612 XThC.Tn[1] XThC.Tn[1].n27 0.396333
R21613 XThC.Tn[1] XThC.Tn[1].n30 0.396333
R21614 XThC.Tn[1] XThC.Tn[1].n33 0.396333
R21615 XThC.Tn[1] XThC.Tn[1].n36 0.396333
R21616 XThC.Tn[1] XThC.Tn[1].n39 0.396333
R21617 XThC.Tn[1] XThC.Tn[1].n42 0.396333
R21618 XThC.Tn[1] XThC.Tn[1].n45 0.396333
R21619 XThC.Tn[1] XThC.Tn[1].n48 0.396333
R21620 XThC.Tn[1] XThC.Tn[1].n51 0.396333
R21621 XThC.Tn[1] XThC.Tn[1].n54 0.396333
R21622 XThC.Tn[1] XThC.Tn[1].n57 0.396333
R21623 XThC.Tn[1].n11 XThC.Tn[1] 0.104667
R21624 XThC.Tn[1].n14 XThC.Tn[1] 0.104667
R21625 XThC.Tn[1].n17 XThC.Tn[1] 0.104667
R21626 XThC.Tn[1].n20 XThC.Tn[1] 0.104667
R21627 XThC.Tn[1].n23 XThC.Tn[1] 0.104667
R21628 XThC.Tn[1].n26 XThC.Tn[1] 0.104667
R21629 XThC.Tn[1].n29 XThC.Tn[1] 0.104667
R21630 XThC.Tn[1].n32 XThC.Tn[1] 0.104667
R21631 XThC.Tn[1].n35 XThC.Tn[1] 0.104667
R21632 XThC.Tn[1].n38 XThC.Tn[1] 0.104667
R21633 XThC.Tn[1].n41 XThC.Tn[1] 0.104667
R21634 XThC.Tn[1].n44 XThC.Tn[1] 0.104667
R21635 XThC.Tn[1].n47 XThC.Tn[1] 0.104667
R21636 XThC.Tn[1].n50 XThC.Tn[1] 0.104667
R21637 XThC.Tn[1].n53 XThC.Tn[1] 0.104667
R21638 XThC.Tn[1].n56 XThC.Tn[1] 0.104667
R21639 XThC.Tn[1].n58 XThC.Tn[1] 0.0594286
R21640 XThC.Tn[1].n11 XThC.Tn[1] 0.0309878
R21641 XThC.Tn[1].n14 XThC.Tn[1] 0.0309878
R21642 XThC.Tn[1].n17 XThC.Tn[1] 0.0309878
R21643 XThC.Tn[1].n20 XThC.Tn[1] 0.0309878
R21644 XThC.Tn[1].n23 XThC.Tn[1] 0.0309878
R21645 XThC.Tn[1].n26 XThC.Tn[1] 0.0309878
R21646 XThC.Tn[1].n29 XThC.Tn[1] 0.0309878
R21647 XThC.Tn[1].n32 XThC.Tn[1] 0.0309878
R21648 XThC.Tn[1].n35 XThC.Tn[1] 0.0309878
R21649 XThC.Tn[1].n38 XThC.Tn[1] 0.0309878
R21650 XThC.Tn[1].n41 XThC.Tn[1] 0.0309878
R21651 XThC.Tn[1].n44 XThC.Tn[1] 0.0309878
R21652 XThC.Tn[1].n47 XThC.Tn[1] 0.0309878
R21653 XThC.Tn[1].n50 XThC.Tn[1] 0.0309878
R21654 XThC.Tn[1].n53 XThC.Tn[1] 0.0309878
R21655 XThC.Tn[1].n56 XThC.Tn[1] 0.0309878
R21656 XThC.Tn[1].n12 XThC.Tn[1].n11 0.027939
R21657 XThC.Tn[1].n15 XThC.Tn[1].n14 0.027939
R21658 XThC.Tn[1].n18 XThC.Tn[1].n17 0.027939
R21659 XThC.Tn[1].n21 XThC.Tn[1].n20 0.027939
R21660 XThC.Tn[1].n24 XThC.Tn[1].n23 0.027939
R21661 XThC.Tn[1].n27 XThC.Tn[1].n26 0.027939
R21662 XThC.Tn[1].n30 XThC.Tn[1].n29 0.027939
R21663 XThC.Tn[1].n33 XThC.Tn[1].n32 0.027939
R21664 XThC.Tn[1].n36 XThC.Tn[1].n35 0.027939
R21665 XThC.Tn[1].n39 XThC.Tn[1].n38 0.027939
R21666 XThC.Tn[1].n42 XThC.Tn[1].n41 0.027939
R21667 XThC.Tn[1].n45 XThC.Tn[1].n44 0.027939
R21668 XThC.Tn[1].n48 XThC.Tn[1].n47 0.027939
R21669 XThC.Tn[1].n51 XThC.Tn[1].n50 0.027939
R21670 XThC.Tn[1].n54 XThC.Tn[1].n53 0.027939
R21671 XThC.Tn[1].n57 XThC.Tn[1].n56 0.027939
R21672 XThC.Tn[3].n2 XThC.Tn[3].n1 332.334
R21673 XThC.Tn[3].n2 XThC.Tn[3].n0 296.493
R21674 XThC.Tn[3].n12 XThC.Tn[3].n10 161.406
R21675 XThC.Tn[3].n15 XThC.Tn[3].n13 161.406
R21676 XThC.Tn[3].n18 XThC.Tn[3].n16 161.406
R21677 XThC.Tn[3].n21 XThC.Tn[3].n19 161.406
R21678 XThC.Tn[3].n24 XThC.Tn[3].n22 161.406
R21679 XThC.Tn[3].n27 XThC.Tn[3].n25 161.406
R21680 XThC.Tn[3].n30 XThC.Tn[3].n28 161.406
R21681 XThC.Tn[3].n33 XThC.Tn[3].n31 161.406
R21682 XThC.Tn[3].n36 XThC.Tn[3].n34 161.406
R21683 XThC.Tn[3].n39 XThC.Tn[3].n37 161.406
R21684 XThC.Tn[3].n42 XThC.Tn[3].n40 161.406
R21685 XThC.Tn[3].n45 XThC.Tn[3].n43 161.406
R21686 XThC.Tn[3].n48 XThC.Tn[3].n46 161.406
R21687 XThC.Tn[3].n51 XThC.Tn[3].n49 161.406
R21688 XThC.Tn[3].n54 XThC.Tn[3].n52 161.406
R21689 XThC.Tn[3].n57 XThC.Tn[3].n55 161.406
R21690 XThC.Tn[3].n10 XThC.Tn[3].t42 161.202
R21691 XThC.Tn[3].n13 XThC.Tn[3].t27 161.202
R21692 XThC.Tn[3].n16 XThC.Tn[3].t29 161.202
R21693 XThC.Tn[3].n19 XThC.Tn[3].t31 161.202
R21694 XThC.Tn[3].n22 XThC.Tn[3].t20 161.202
R21695 XThC.Tn[3].n25 XThC.Tn[3].t21 161.202
R21696 XThC.Tn[3].n28 XThC.Tn[3].t34 161.202
R21697 XThC.Tn[3].n31 XThC.Tn[3].t43 161.202
R21698 XThC.Tn[3].n34 XThC.Tn[3].t13 161.202
R21699 XThC.Tn[3].n37 XThC.Tn[3].t32 161.202
R21700 XThC.Tn[3].n40 XThC.Tn[3].t33 161.202
R21701 XThC.Tn[3].n43 XThC.Tn[3].t14 161.202
R21702 XThC.Tn[3].n46 XThC.Tn[3].t22 161.202
R21703 XThC.Tn[3].n49 XThC.Tn[3].t25 161.202
R21704 XThC.Tn[3].n52 XThC.Tn[3].t38 161.202
R21705 XThC.Tn[3].n55 XThC.Tn[3].t16 161.202
R21706 XThC.Tn[3].n10 XThC.Tn[3].t12 145.137
R21707 XThC.Tn[3].n13 XThC.Tn[3].t30 145.137
R21708 XThC.Tn[3].n16 XThC.Tn[3].t35 145.137
R21709 XThC.Tn[3].n19 XThC.Tn[3].t36 145.137
R21710 XThC.Tn[3].n22 XThC.Tn[3].t23 145.137
R21711 XThC.Tn[3].n25 XThC.Tn[3].t24 145.137
R21712 XThC.Tn[3].n28 XThC.Tn[3].t40 145.137
R21713 XThC.Tn[3].n31 XThC.Tn[3].t15 145.137
R21714 XThC.Tn[3].n34 XThC.Tn[3].t17 145.137
R21715 XThC.Tn[3].n37 XThC.Tn[3].t37 145.137
R21716 XThC.Tn[3].n40 XThC.Tn[3].t39 145.137
R21717 XThC.Tn[3].n43 XThC.Tn[3].t18 145.137
R21718 XThC.Tn[3].n46 XThC.Tn[3].t26 145.137
R21719 XThC.Tn[3].n49 XThC.Tn[3].t28 145.137
R21720 XThC.Tn[3].n52 XThC.Tn[3].t41 145.137
R21721 XThC.Tn[3].n55 XThC.Tn[3].t19 145.137
R21722 XThC.Tn[3].n5 XThC.Tn[3].n3 135.249
R21723 XThC.Tn[3].n5 XThC.Tn[3].n4 98.981
R21724 XThC.Tn[3].n7 XThC.Tn[3].n6 98.981
R21725 XThC.Tn[3].n9 XThC.Tn[3].n8 98.981
R21726 XThC.Tn[3].n7 XThC.Tn[3].n5 36.2672
R21727 XThC.Tn[3].n9 XThC.Tn[3].n7 36.2672
R21728 XThC.Tn[3].n58 XThC.Tn[3].n9 32.6405
R21729 XThC.Tn[3].n0 XThC.Tn[3].t1 26.5955
R21730 XThC.Tn[3].n0 XThC.Tn[3].t0 26.5955
R21731 XThC.Tn[3].n1 XThC.Tn[3].t3 26.5955
R21732 XThC.Tn[3].n1 XThC.Tn[3].t2 26.5955
R21733 XThC.Tn[3].n3 XThC.Tn[3].t11 24.9236
R21734 XThC.Tn[3].n3 XThC.Tn[3].t10 24.9236
R21735 XThC.Tn[3].n4 XThC.Tn[3].t9 24.9236
R21736 XThC.Tn[3].n4 XThC.Tn[3].t8 24.9236
R21737 XThC.Tn[3].n6 XThC.Tn[3].t7 24.9236
R21738 XThC.Tn[3].n6 XThC.Tn[3].t6 24.9236
R21739 XThC.Tn[3].n8 XThC.Tn[3].t5 24.9236
R21740 XThC.Tn[3].n8 XThC.Tn[3].t4 24.9236
R21741 XThC.Tn[3] XThC.Tn[3].n2 23.3605
R21742 XThC.Tn[3] XThC.Tn[3].n58 6.7205
R21743 XThC.Tn[3].n58 XThC.Tn[3] 3.19574
R21744 XThC.Tn[3].n15 XThC.Tn[3] 0.931056
R21745 XThC.Tn[3].n18 XThC.Tn[3] 0.931056
R21746 XThC.Tn[3].n21 XThC.Tn[3] 0.931056
R21747 XThC.Tn[3].n24 XThC.Tn[3] 0.931056
R21748 XThC.Tn[3].n27 XThC.Tn[3] 0.931056
R21749 XThC.Tn[3].n30 XThC.Tn[3] 0.931056
R21750 XThC.Tn[3].n33 XThC.Tn[3] 0.931056
R21751 XThC.Tn[3].n36 XThC.Tn[3] 0.931056
R21752 XThC.Tn[3].n39 XThC.Tn[3] 0.931056
R21753 XThC.Tn[3].n42 XThC.Tn[3] 0.931056
R21754 XThC.Tn[3].n45 XThC.Tn[3] 0.931056
R21755 XThC.Tn[3].n48 XThC.Tn[3] 0.931056
R21756 XThC.Tn[3].n51 XThC.Tn[3] 0.931056
R21757 XThC.Tn[3].n54 XThC.Tn[3] 0.931056
R21758 XThC.Tn[3].n57 XThC.Tn[3] 0.931056
R21759 XThC.Tn[3] XThC.Tn[3].n12 0.396333
R21760 XThC.Tn[3] XThC.Tn[3].n15 0.396333
R21761 XThC.Tn[3] XThC.Tn[3].n18 0.396333
R21762 XThC.Tn[3] XThC.Tn[3].n21 0.396333
R21763 XThC.Tn[3] XThC.Tn[3].n24 0.396333
R21764 XThC.Tn[3] XThC.Tn[3].n27 0.396333
R21765 XThC.Tn[3] XThC.Tn[3].n30 0.396333
R21766 XThC.Tn[3] XThC.Tn[3].n33 0.396333
R21767 XThC.Tn[3] XThC.Tn[3].n36 0.396333
R21768 XThC.Tn[3] XThC.Tn[3].n39 0.396333
R21769 XThC.Tn[3] XThC.Tn[3].n42 0.396333
R21770 XThC.Tn[3] XThC.Tn[3].n45 0.396333
R21771 XThC.Tn[3] XThC.Tn[3].n48 0.396333
R21772 XThC.Tn[3] XThC.Tn[3].n51 0.396333
R21773 XThC.Tn[3] XThC.Tn[3].n54 0.396333
R21774 XThC.Tn[3] XThC.Tn[3].n57 0.396333
R21775 XThC.Tn[3].n11 XThC.Tn[3] 0.104667
R21776 XThC.Tn[3].n14 XThC.Tn[3] 0.104667
R21777 XThC.Tn[3].n17 XThC.Tn[3] 0.104667
R21778 XThC.Tn[3].n20 XThC.Tn[3] 0.104667
R21779 XThC.Tn[3].n23 XThC.Tn[3] 0.104667
R21780 XThC.Tn[3].n26 XThC.Tn[3] 0.104667
R21781 XThC.Tn[3].n29 XThC.Tn[3] 0.104667
R21782 XThC.Tn[3].n32 XThC.Tn[3] 0.104667
R21783 XThC.Tn[3].n35 XThC.Tn[3] 0.104667
R21784 XThC.Tn[3].n38 XThC.Tn[3] 0.104667
R21785 XThC.Tn[3].n41 XThC.Tn[3] 0.104667
R21786 XThC.Tn[3].n44 XThC.Tn[3] 0.104667
R21787 XThC.Tn[3].n47 XThC.Tn[3] 0.104667
R21788 XThC.Tn[3].n50 XThC.Tn[3] 0.104667
R21789 XThC.Tn[3].n53 XThC.Tn[3] 0.104667
R21790 XThC.Tn[3].n56 XThC.Tn[3] 0.104667
R21791 XThC.Tn[3].n11 XThC.Tn[3] 0.0309878
R21792 XThC.Tn[3].n14 XThC.Tn[3] 0.0309878
R21793 XThC.Tn[3].n17 XThC.Tn[3] 0.0309878
R21794 XThC.Tn[3].n20 XThC.Tn[3] 0.0309878
R21795 XThC.Tn[3].n23 XThC.Tn[3] 0.0309878
R21796 XThC.Tn[3].n26 XThC.Tn[3] 0.0309878
R21797 XThC.Tn[3].n29 XThC.Tn[3] 0.0309878
R21798 XThC.Tn[3].n32 XThC.Tn[3] 0.0309878
R21799 XThC.Tn[3].n35 XThC.Tn[3] 0.0309878
R21800 XThC.Tn[3].n38 XThC.Tn[3] 0.0309878
R21801 XThC.Tn[3].n41 XThC.Tn[3] 0.0309878
R21802 XThC.Tn[3].n44 XThC.Tn[3] 0.0309878
R21803 XThC.Tn[3].n47 XThC.Tn[3] 0.0309878
R21804 XThC.Tn[3].n50 XThC.Tn[3] 0.0309878
R21805 XThC.Tn[3].n53 XThC.Tn[3] 0.0309878
R21806 XThC.Tn[3].n56 XThC.Tn[3] 0.0309878
R21807 XThC.Tn[3].n12 XThC.Tn[3].n11 0.027939
R21808 XThC.Tn[3].n15 XThC.Tn[3].n14 0.027939
R21809 XThC.Tn[3].n18 XThC.Tn[3].n17 0.027939
R21810 XThC.Tn[3].n21 XThC.Tn[3].n20 0.027939
R21811 XThC.Tn[3].n24 XThC.Tn[3].n23 0.027939
R21812 XThC.Tn[3].n27 XThC.Tn[3].n26 0.027939
R21813 XThC.Tn[3].n30 XThC.Tn[3].n29 0.027939
R21814 XThC.Tn[3].n33 XThC.Tn[3].n32 0.027939
R21815 XThC.Tn[3].n36 XThC.Tn[3].n35 0.027939
R21816 XThC.Tn[3].n39 XThC.Tn[3].n38 0.027939
R21817 XThC.Tn[3].n42 XThC.Tn[3].n41 0.027939
R21818 XThC.Tn[3].n45 XThC.Tn[3].n44 0.027939
R21819 XThC.Tn[3].n48 XThC.Tn[3].n47 0.027939
R21820 XThC.Tn[3].n51 XThC.Tn[3].n50 0.027939
R21821 XThC.Tn[3].n54 XThC.Tn[3].n53 0.027939
R21822 XThC.Tn[3].n57 XThC.Tn[3].n56 0.027939
R21823 XThR.Tn[10].n5 XThR.Tn[10].n4 256.103
R21824 XThR.Tn[10].n2 XThR.Tn[10].n0 243.68
R21825 XThR.Tn[10].n88 XThR.Tn[10].n87 241.847
R21826 XThR.Tn[10].n2 XThR.Tn[10].n1 205.28
R21827 XThR.Tn[10].n5 XThR.Tn[10].n3 202.095
R21828 XThR.Tn[10].n88 XThR.Tn[10].n86 185
R21829 XThR.Tn[10] XThR.Tn[10].n79 161.363
R21830 XThR.Tn[10] XThR.Tn[10].n74 161.363
R21831 XThR.Tn[10] XThR.Tn[10].n69 161.363
R21832 XThR.Tn[10] XThR.Tn[10].n64 161.363
R21833 XThR.Tn[10] XThR.Tn[10].n59 161.363
R21834 XThR.Tn[10] XThR.Tn[10].n54 161.363
R21835 XThR.Tn[10] XThR.Tn[10].n49 161.363
R21836 XThR.Tn[10] XThR.Tn[10].n44 161.363
R21837 XThR.Tn[10] XThR.Tn[10].n39 161.363
R21838 XThR.Tn[10] XThR.Tn[10].n34 161.363
R21839 XThR.Tn[10] XThR.Tn[10].n29 161.363
R21840 XThR.Tn[10] XThR.Tn[10].n24 161.363
R21841 XThR.Tn[10] XThR.Tn[10].n19 161.363
R21842 XThR.Tn[10] XThR.Tn[10].n14 161.363
R21843 XThR.Tn[10] XThR.Tn[10].n9 161.363
R21844 XThR.Tn[10] XThR.Tn[10].n7 161.363
R21845 XThR.Tn[10].n81 XThR.Tn[10].n80 161.3
R21846 XThR.Tn[10].n76 XThR.Tn[10].n75 161.3
R21847 XThR.Tn[10].n71 XThR.Tn[10].n70 161.3
R21848 XThR.Tn[10].n66 XThR.Tn[10].n65 161.3
R21849 XThR.Tn[10].n61 XThR.Tn[10].n60 161.3
R21850 XThR.Tn[10].n56 XThR.Tn[10].n55 161.3
R21851 XThR.Tn[10].n51 XThR.Tn[10].n50 161.3
R21852 XThR.Tn[10].n46 XThR.Tn[10].n45 161.3
R21853 XThR.Tn[10].n41 XThR.Tn[10].n40 161.3
R21854 XThR.Tn[10].n36 XThR.Tn[10].n35 161.3
R21855 XThR.Tn[10].n31 XThR.Tn[10].n30 161.3
R21856 XThR.Tn[10].n26 XThR.Tn[10].n25 161.3
R21857 XThR.Tn[10].n21 XThR.Tn[10].n20 161.3
R21858 XThR.Tn[10].n16 XThR.Tn[10].n15 161.3
R21859 XThR.Tn[10].n11 XThR.Tn[10].n10 161.3
R21860 XThR.Tn[10].n79 XThR.Tn[10].t37 161.106
R21861 XThR.Tn[10].n74 XThR.Tn[10].t45 161.106
R21862 XThR.Tn[10].n69 XThR.Tn[10].t27 161.106
R21863 XThR.Tn[10].n64 XThR.Tn[10].t72 161.106
R21864 XThR.Tn[10].n59 XThR.Tn[10].t35 161.106
R21865 XThR.Tn[10].n54 XThR.Tn[10].t61 161.106
R21866 XThR.Tn[10].n49 XThR.Tn[10].t43 161.106
R21867 XThR.Tn[10].n44 XThR.Tn[10].t24 161.106
R21868 XThR.Tn[10].n39 XThR.Tn[10].t69 161.106
R21869 XThR.Tn[10].n34 XThR.Tn[10].t15 161.106
R21870 XThR.Tn[10].n29 XThR.Tn[10].t59 161.106
R21871 XThR.Tn[10].n24 XThR.Tn[10].t26 161.106
R21872 XThR.Tn[10].n19 XThR.Tn[10].t58 161.106
R21873 XThR.Tn[10].n14 XThR.Tn[10].t41 161.106
R21874 XThR.Tn[10].n9 XThR.Tn[10].t63 161.106
R21875 XThR.Tn[10].n7 XThR.Tn[10].t47 161.106
R21876 XThR.Tn[10].n80 XThR.Tn[10].t34 159.978
R21877 XThR.Tn[10].n75 XThR.Tn[10].t39 159.978
R21878 XThR.Tn[10].n70 XThR.Tn[10].t22 159.978
R21879 XThR.Tn[10].n65 XThR.Tn[10].t68 159.978
R21880 XThR.Tn[10].n60 XThR.Tn[10].t32 159.978
R21881 XThR.Tn[10].n55 XThR.Tn[10].t57 159.978
R21882 XThR.Tn[10].n50 XThR.Tn[10].t38 159.978
R21883 XThR.Tn[10].n45 XThR.Tn[10].t20 159.978
R21884 XThR.Tn[10].n40 XThR.Tn[10].t66 159.978
R21885 XThR.Tn[10].n35 XThR.Tn[10].t12 159.978
R21886 XThR.Tn[10].n30 XThR.Tn[10].t56 159.978
R21887 XThR.Tn[10].n25 XThR.Tn[10].t21 159.978
R21888 XThR.Tn[10].n20 XThR.Tn[10].t55 159.978
R21889 XThR.Tn[10].n15 XThR.Tn[10].t36 159.978
R21890 XThR.Tn[10].n10 XThR.Tn[10].t60 159.978
R21891 XThR.Tn[10].n79 XThR.Tn[10].t29 145.038
R21892 XThR.Tn[10].n74 XThR.Tn[10].t49 145.038
R21893 XThR.Tn[10].n69 XThR.Tn[10].t31 145.038
R21894 XThR.Tn[10].n64 XThR.Tn[10].t16 145.038
R21895 XThR.Tn[10].n59 XThR.Tn[10].t46 145.038
R21896 XThR.Tn[10].n54 XThR.Tn[10].t28 145.038
R21897 XThR.Tn[10].n49 XThR.Tn[10].t33 145.038
R21898 XThR.Tn[10].n44 XThR.Tn[10].t17 145.038
R21899 XThR.Tn[10].n39 XThR.Tn[10].t14 145.038
R21900 XThR.Tn[10].n34 XThR.Tn[10].t44 145.038
R21901 XThR.Tn[10].n29 XThR.Tn[10].t67 145.038
R21902 XThR.Tn[10].n24 XThR.Tn[10].t30 145.038
R21903 XThR.Tn[10].n19 XThR.Tn[10].t65 145.038
R21904 XThR.Tn[10].n14 XThR.Tn[10].t48 145.038
R21905 XThR.Tn[10].n9 XThR.Tn[10].t13 145.038
R21906 XThR.Tn[10].n7 XThR.Tn[10].t54 145.038
R21907 XThR.Tn[10].n80 XThR.Tn[10].t64 143.911
R21908 XThR.Tn[10].n75 XThR.Tn[10].t25 143.911
R21909 XThR.Tn[10].n70 XThR.Tn[10].t71 143.911
R21910 XThR.Tn[10].n65 XThR.Tn[10].t52 143.911
R21911 XThR.Tn[10].n60 XThR.Tn[10].t19 143.911
R21912 XThR.Tn[10].n55 XThR.Tn[10].t62 143.911
R21913 XThR.Tn[10].n50 XThR.Tn[10].t73 143.911
R21914 XThR.Tn[10].n45 XThR.Tn[10].t53 143.911
R21915 XThR.Tn[10].n40 XThR.Tn[10].t51 143.911
R21916 XThR.Tn[10].n35 XThR.Tn[10].t18 143.911
R21917 XThR.Tn[10].n30 XThR.Tn[10].t42 143.911
R21918 XThR.Tn[10].n25 XThR.Tn[10].t70 143.911
R21919 XThR.Tn[10].n20 XThR.Tn[10].t40 143.911
R21920 XThR.Tn[10].n15 XThR.Tn[10].t23 143.911
R21921 XThR.Tn[10].n10 XThR.Tn[10].t50 143.911
R21922 XThR.Tn[10] XThR.Tn[10].n2 35.7652
R21923 XThR.Tn[10].n3 XThR.Tn[10].t6 26.5955
R21924 XThR.Tn[10].n3 XThR.Tn[10].t4 26.5955
R21925 XThR.Tn[10].n4 XThR.Tn[10].t7 26.5955
R21926 XThR.Tn[10].n4 XThR.Tn[10].t5 26.5955
R21927 XThR.Tn[10].n0 XThR.Tn[10].t10 26.5955
R21928 XThR.Tn[10].n0 XThR.Tn[10].t8 26.5955
R21929 XThR.Tn[10].n1 XThR.Tn[10].t11 26.5955
R21930 XThR.Tn[10].n1 XThR.Tn[10].t9 26.5955
R21931 XThR.Tn[10].n86 XThR.Tn[10].t0 24.9236
R21932 XThR.Tn[10].n86 XThR.Tn[10].t2 24.9236
R21933 XThR.Tn[10].n87 XThR.Tn[10].t1 24.9236
R21934 XThR.Tn[10].n87 XThR.Tn[10].t3 24.9236
R21935 XThR.Tn[10] XThR.Tn[10].n88 18.8943
R21936 XThR.Tn[10].n6 XThR.Tn[10].n5 13.5534
R21937 XThR.Tn[10].n85 XThR.Tn[10] 7.84567
R21938 XThR.Tn[10] XThR.Tn[10].n85 6.34069
R21939 XThR.Tn[10] XThR.Tn[10].n8 5.34038
R21940 XThR.Tn[10].n13 XThR.Tn[10].n12 4.5005
R21941 XThR.Tn[10].n18 XThR.Tn[10].n17 4.5005
R21942 XThR.Tn[10].n23 XThR.Tn[10].n22 4.5005
R21943 XThR.Tn[10].n28 XThR.Tn[10].n27 4.5005
R21944 XThR.Tn[10].n33 XThR.Tn[10].n32 4.5005
R21945 XThR.Tn[10].n38 XThR.Tn[10].n37 4.5005
R21946 XThR.Tn[10].n43 XThR.Tn[10].n42 4.5005
R21947 XThR.Tn[10].n48 XThR.Tn[10].n47 4.5005
R21948 XThR.Tn[10].n53 XThR.Tn[10].n52 4.5005
R21949 XThR.Tn[10].n58 XThR.Tn[10].n57 4.5005
R21950 XThR.Tn[10].n63 XThR.Tn[10].n62 4.5005
R21951 XThR.Tn[10].n68 XThR.Tn[10].n67 4.5005
R21952 XThR.Tn[10].n73 XThR.Tn[10].n72 4.5005
R21953 XThR.Tn[10].n78 XThR.Tn[10].n77 4.5005
R21954 XThR.Tn[10].n83 XThR.Tn[10].n82 4.5005
R21955 XThR.Tn[10].n84 XThR.Tn[10] 3.70586
R21956 XThR.Tn[10].n13 XThR.Tn[10] 2.52282
R21957 XThR.Tn[10].n18 XThR.Tn[10] 2.52282
R21958 XThR.Tn[10].n23 XThR.Tn[10] 2.52282
R21959 XThR.Tn[10].n28 XThR.Tn[10] 2.52282
R21960 XThR.Tn[10].n33 XThR.Tn[10] 2.52282
R21961 XThR.Tn[10].n38 XThR.Tn[10] 2.52282
R21962 XThR.Tn[10].n43 XThR.Tn[10] 2.52282
R21963 XThR.Tn[10].n48 XThR.Tn[10] 2.52282
R21964 XThR.Tn[10].n53 XThR.Tn[10] 2.52282
R21965 XThR.Tn[10].n58 XThR.Tn[10] 2.52282
R21966 XThR.Tn[10].n63 XThR.Tn[10] 2.52282
R21967 XThR.Tn[10].n68 XThR.Tn[10] 2.52282
R21968 XThR.Tn[10].n73 XThR.Tn[10] 2.52282
R21969 XThR.Tn[10].n78 XThR.Tn[10] 2.52282
R21970 XThR.Tn[10].n83 XThR.Tn[10] 2.52282
R21971 XThR.Tn[10].n85 XThR.Tn[10] 1.79489
R21972 XThR.Tn[10].n6 XThR.Tn[10] 1.50638
R21973 XThR.Tn[10] XThR.Tn[10].n6 1.19676
R21974 XThR.Tn[10].n81 XThR.Tn[10] 1.08677
R21975 XThR.Tn[10].n76 XThR.Tn[10] 1.08677
R21976 XThR.Tn[10].n71 XThR.Tn[10] 1.08677
R21977 XThR.Tn[10].n66 XThR.Tn[10] 1.08677
R21978 XThR.Tn[10].n61 XThR.Tn[10] 1.08677
R21979 XThR.Tn[10].n56 XThR.Tn[10] 1.08677
R21980 XThR.Tn[10].n51 XThR.Tn[10] 1.08677
R21981 XThR.Tn[10].n46 XThR.Tn[10] 1.08677
R21982 XThR.Tn[10].n41 XThR.Tn[10] 1.08677
R21983 XThR.Tn[10].n36 XThR.Tn[10] 1.08677
R21984 XThR.Tn[10].n31 XThR.Tn[10] 1.08677
R21985 XThR.Tn[10].n26 XThR.Tn[10] 1.08677
R21986 XThR.Tn[10].n21 XThR.Tn[10] 1.08677
R21987 XThR.Tn[10].n16 XThR.Tn[10] 1.08677
R21988 XThR.Tn[10].n11 XThR.Tn[10] 1.08677
R21989 XThR.Tn[10] XThR.Tn[10].n13 0.839786
R21990 XThR.Tn[10] XThR.Tn[10].n18 0.839786
R21991 XThR.Tn[10] XThR.Tn[10].n23 0.839786
R21992 XThR.Tn[10] XThR.Tn[10].n28 0.839786
R21993 XThR.Tn[10] XThR.Tn[10].n33 0.839786
R21994 XThR.Tn[10] XThR.Tn[10].n38 0.839786
R21995 XThR.Tn[10] XThR.Tn[10].n43 0.839786
R21996 XThR.Tn[10] XThR.Tn[10].n48 0.839786
R21997 XThR.Tn[10] XThR.Tn[10].n53 0.839786
R21998 XThR.Tn[10] XThR.Tn[10].n58 0.839786
R21999 XThR.Tn[10] XThR.Tn[10].n63 0.839786
R22000 XThR.Tn[10] XThR.Tn[10].n68 0.839786
R22001 XThR.Tn[10] XThR.Tn[10].n73 0.839786
R22002 XThR.Tn[10] XThR.Tn[10].n78 0.839786
R22003 XThR.Tn[10] XThR.Tn[10].n83 0.839786
R22004 XThR.Tn[10].n8 XThR.Tn[10] 0.499542
R22005 XThR.Tn[10].n82 XThR.Tn[10] 0.063
R22006 XThR.Tn[10].n77 XThR.Tn[10] 0.063
R22007 XThR.Tn[10].n72 XThR.Tn[10] 0.063
R22008 XThR.Tn[10].n67 XThR.Tn[10] 0.063
R22009 XThR.Tn[10].n62 XThR.Tn[10] 0.063
R22010 XThR.Tn[10].n57 XThR.Tn[10] 0.063
R22011 XThR.Tn[10].n52 XThR.Tn[10] 0.063
R22012 XThR.Tn[10].n47 XThR.Tn[10] 0.063
R22013 XThR.Tn[10].n42 XThR.Tn[10] 0.063
R22014 XThR.Tn[10].n37 XThR.Tn[10] 0.063
R22015 XThR.Tn[10].n32 XThR.Tn[10] 0.063
R22016 XThR.Tn[10].n27 XThR.Tn[10] 0.063
R22017 XThR.Tn[10].n22 XThR.Tn[10] 0.063
R22018 XThR.Tn[10].n17 XThR.Tn[10] 0.063
R22019 XThR.Tn[10].n12 XThR.Tn[10] 0.063
R22020 XThR.Tn[10].n84 XThR.Tn[10] 0.0540714
R22021 XThR.Tn[10] XThR.Tn[10].n84 0.038
R22022 XThR.Tn[10].n8 XThR.Tn[10] 0.0143889
R22023 XThR.Tn[10].n82 XThR.Tn[10].n81 0.00771154
R22024 XThR.Tn[10].n77 XThR.Tn[10].n76 0.00771154
R22025 XThR.Tn[10].n72 XThR.Tn[10].n71 0.00771154
R22026 XThR.Tn[10].n67 XThR.Tn[10].n66 0.00771154
R22027 XThR.Tn[10].n62 XThR.Tn[10].n61 0.00771154
R22028 XThR.Tn[10].n57 XThR.Tn[10].n56 0.00771154
R22029 XThR.Tn[10].n52 XThR.Tn[10].n51 0.00771154
R22030 XThR.Tn[10].n47 XThR.Tn[10].n46 0.00771154
R22031 XThR.Tn[10].n42 XThR.Tn[10].n41 0.00771154
R22032 XThR.Tn[10].n37 XThR.Tn[10].n36 0.00771154
R22033 XThR.Tn[10].n32 XThR.Tn[10].n31 0.00771154
R22034 XThR.Tn[10].n27 XThR.Tn[10].n26 0.00771154
R22035 XThR.Tn[10].n22 XThR.Tn[10].n21 0.00771154
R22036 XThR.Tn[10].n17 XThR.Tn[10].n16 0.00771154
R22037 XThR.Tn[10].n12 XThR.Tn[10].n11 0.00771154
R22038 XThC.Tn[14].n5 XThC.Tn[14].n4 256.104
R22039 XThC.Tn[14].n8 XThC.Tn[14].n6 243.68
R22040 XThC.Tn[14].n2 XThC.Tn[14].n0 241.847
R22041 XThC.Tn[14].n8 XThC.Tn[14].n7 205.28
R22042 XThC.Tn[14].n5 XThC.Tn[14].n3 202.095
R22043 XThC.Tn[14].n2 XThC.Tn[14].n1 185
R22044 XThC.Tn[14].n12 XThC.Tn[14].n10 161.406
R22045 XThC.Tn[14].n15 XThC.Tn[14].n13 161.406
R22046 XThC.Tn[14].n18 XThC.Tn[14].n16 161.406
R22047 XThC.Tn[14].n21 XThC.Tn[14].n19 161.406
R22048 XThC.Tn[14].n24 XThC.Tn[14].n22 161.406
R22049 XThC.Tn[14].n27 XThC.Tn[14].n25 161.406
R22050 XThC.Tn[14].n30 XThC.Tn[14].n28 161.406
R22051 XThC.Tn[14].n33 XThC.Tn[14].n31 161.406
R22052 XThC.Tn[14].n36 XThC.Tn[14].n34 161.406
R22053 XThC.Tn[14].n39 XThC.Tn[14].n37 161.406
R22054 XThC.Tn[14].n42 XThC.Tn[14].n40 161.406
R22055 XThC.Tn[14].n45 XThC.Tn[14].n43 161.406
R22056 XThC.Tn[14].n48 XThC.Tn[14].n46 161.406
R22057 XThC.Tn[14].n51 XThC.Tn[14].n49 161.406
R22058 XThC.Tn[14].n54 XThC.Tn[14].n52 161.406
R22059 XThC.Tn[14].n57 XThC.Tn[14].n55 161.406
R22060 XThC.Tn[14].n10 XThC.Tn[14].t38 161.202
R22061 XThC.Tn[14].n13 XThC.Tn[14].t22 161.202
R22062 XThC.Tn[14].n16 XThC.Tn[14].t25 161.202
R22063 XThC.Tn[14].n19 XThC.Tn[14].t26 161.202
R22064 XThC.Tn[14].n22 XThC.Tn[14].t14 161.202
R22065 XThC.Tn[14].n25 XThC.Tn[14].t17 161.202
R22066 XThC.Tn[14].n28 XThC.Tn[14].t31 161.202
R22067 XThC.Tn[14].n31 XThC.Tn[14].t39 161.202
R22068 XThC.Tn[14].n34 XThC.Tn[14].t41 161.202
R22069 XThC.Tn[14].n37 XThC.Tn[14].t27 161.202
R22070 XThC.Tn[14].n40 XThC.Tn[14].t30 161.202
R22071 XThC.Tn[14].n43 XThC.Tn[14].t42 161.202
R22072 XThC.Tn[14].n46 XThC.Tn[14].t19 161.202
R22073 XThC.Tn[14].n49 XThC.Tn[14].t21 161.202
R22074 XThC.Tn[14].n52 XThC.Tn[14].t33 161.202
R22075 XThC.Tn[14].n55 XThC.Tn[14].t12 161.202
R22076 XThC.Tn[14].n10 XThC.Tn[14].t43 145.137
R22077 XThC.Tn[14].n13 XThC.Tn[14].t29 145.137
R22078 XThC.Tn[14].n16 XThC.Tn[14].t32 145.137
R22079 XThC.Tn[14].n19 XThC.Tn[14].t34 145.137
R22080 XThC.Tn[14].n22 XThC.Tn[14].t20 145.137
R22081 XThC.Tn[14].n25 XThC.Tn[14].t23 145.137
R22082 XThC.Tn[14].n28 XThC.Tn[14].t37 145.137
R22083 XThC.Tn[14].n31 XThC.Tn[14].t13 145.137
R22084 XThC.Tn[14].n34 XThC.Tn[14].t15 145.137
R22085 XThC.Tn[14].n37 XThC.Tn[14].t35 145.137
R22086 XThC.Tn[14].n40 XThC.Tn[14].t36 145.137
R22087 XThC.Tn[14].n43 XThC.Tn[14].t16 145.137
R22088 XThC.Tn[14].n46 XThC.Tn[14].t24 145.137
R22089 XThC.Tn[14].n49 XThC.Tn[14].t28 145.137
R22090 XThC.Tn[14].n52 XThC.Tn[14].t40 145.137
R22091 XThC.Tn[14].n55 XThC.Tn[14].t18 145.137
R22092 XThC.Tn[14].n3 XThC.Tn[14].t4 26.5955
R22093 XThC.Tn[14].n3 XThC.Tn[14].t5 26.5955
R22094 XThC.Tn[14].n4 XThC.Tn[14].t7 26.5955
R22095 XThC.Tn[14].n4 XThC.Tn[14].t6 26.5955
R22096 XThC.Tn[14].n6 XThC.Tn[14].t11 26.5955
R22097 XThC.Tn[14].n6 XThC.Tn[14].t10 26.5955
R22098 XThC.Tn[14].n7 XThC.Tn[14].t9 26.5955
R22099 XThC.Tn[14].n7 XThC.Tn[14].t8 26.5955
R22100 XThC.Tn[14].n0 XThC.Tn[14].t0 24.9236
R22101 XThC.Tn[14].n0 XThC.Tn[14].t2 24.9236
R22102 XThC.Tn[14].n1 XThC.Tn[14].t1 24.9236
R22103 XThC.Tn[14].n1 XThC.Tn[14].t3 24.9236
R22104 XThC.Tn[14] XThC.Tn[14].n8 22.9652
R22105 XThC.Tn[14] XThC.Tn[14].n2 22.9615
R22106 XThC.Tn[14].n9 XThC.Tn[14].n5 13.9299
R22107 XThC.Tn[14].n9 XThC.Tn[14] 13.9299
R22108 XThC.Tn[14].n58 XThC.Tn[14] 5.65386
R22109 XThC.Tn[14].n59 XThC.Tn[14].n58 5.13312
R22110 XThC.Tn[14].n59 XThC.Tn[14].n9 2.99115
R22111 XThC.Tn[14].n9 XThC.Tn[14] 2.87153
R22112 XThC.Tn[14] XThC.Tn[14].n59 2.2734
R22113 XThC.Tn[14].n15 XThC.Tn[14] 0.931056
R22114 XThC.Tn[14].n18 XThC.Tn[14] 0.931056
R22115 XThC.Tn[14].n21 XThC.Tn[14] 0.931056
R22116 XThC.Tn[14].n24 XThC.Tn[14] 0.931056
R22117 XThC.Tn[14].n27 XThC.Tn[14] 0.931056
R22118 XThC.Tn[14].n30 XThC.Tn[14] 0.931056
R22119 XThC.Tn[14].n33 XThC.Tn[14] 0.931056
R22120 XThC.Tn[14].n36 XThC.Tn[14] 0.931056
R22121 XThC.Tn[14].n39 XThC.Tn[14] 0.931056
R22122 XThC.Tn[14].n42 XThC.Tn[14] 0.931056
R22123 XThC.Tn[14].n45 XThC.Tn[14] 0.931056
R22124 XThC.Tn[14].n48 XThC.Tn[14] 0.931056
R22125 XThC.Tn[14].n51 XThC.Tn[14] 0.931056
R22126 XThC.Tn[14].n54 XThC.Tn[14] 0.931056
R22127 XThC.Tn[14].n57 XThC.Tn[14] 0.931056
R22128 XThC.Tn[14] XThC.Tn[14].n12 0.396333
R22129 XThC.Tn[14] XThC.Tn[14].n15 0.396333
R22130 XThC.Tn[14] XThC.Tn[14].n18 0.396333
R22131 XThC.Tn[14] XThC.Tn[14].n21 0.396333
R22132 XThC.Tn[14] XThC.Tn[14].n24 0.396333
R22133 XThC.Tn[14] XThC.Tn[14].n27 0.396333
R22134 XThC.Tn[14] XThC.Tn[14].n30 0.396333
R22135 XThC.Tn[14] XThC.Tn[14].n33 0.396333
R22136 XThC.Tn[14] XThC.Tn[14].n36 0.396333
R22137 XThC.Tn[14] XThC.Tn[14].n39 0.396333
R22138 XThC.Tn[14] XThC.Tn[14].n42 0.396333
R22139 XThC.Tn[14] XThC.Tn[14].n45 0.396333
R22140 XThC.Tn[14] XThC.Tn[14].n48 0.396333
R22141 XThC.Tn[14] XThC.Tn[14].n51 0.396333
R22142 XThC.Tn[14] XThC.Tn[14].n54 0.396333
R22143 XThC.Tn[14] XThC.Tn[14].n57 0.396333
R22144 XThC.Tn[14].n11 XThC.Tn[14] 0.104667
R22145 XThC.Tn[14].n14 XThC.Tn[14] 0.104667
R22146 XThC.Tn[14].n17 XThC.Tn[14] 0.104667
R22147 XThC.Tn[14].n20 XThC.Tn[14] 0.104667
R22148 XThC.Tn[14].n23 XThC.Tn[14] 0.104667
R22149 XThC.Tn[14].n26 XThC.Tn[14] 0.104667
R22150 XThC.Tn[14].n29 XThC.Tn[14] 0.104667
R22151 XThC.Tn[14].n32 XThC.Tn[14] 0.104667
R22152 XThC.Tn[14].n35 XThC.Tn[14] 0.104667
R22153 XThC.Tn[14].n38 XThC.Tn[14] 0.104667
R22154 XThC.Tn[14].n41 XThC.Tn[14] 0.104667
R22155 XThC.Tn[14].n44 XThC.Tn[14] 0.104667
R22156 XThC.Tn[14].n47 XThC.Tn[14] 0.104667
R22157 XThC.Tn[14].n50 XThC.Tn[14] 0.104667
R22158 XThC.Tn[14].n53 XThC.Tn[14] 0.104667
R22159 XThC.Tn[14].n56 XThC.Tn[14] 0.104667
R22160 XThC.Tn[14].n11 XThC.Tn[14] 0.0309878
R22161 XThC.Tn[14].n14 XThC.Tn[14] 0.0309878
R22162 XThC.Tn[14].n17 XThC.Tn[14] 0.0309878
R22163 XThC.Tn[14].n20 XThC.Tn[14] 0.0309878
R22164 XThC.Tn[14].n23 XThC.Tn[14] 0.0309878
R22165 XThC.Tn[14].n26 XThC.Tn[14] 0.0309878
R22166 XThC.Tn[14].n29 XThC.Tn[14] 0.0309878
R22167 XThC.Tn[14].n32 XThC.Tn[14] 0.0309878
R22168 XThC.Tn[14].n35 XThC.Tn[14] 0.0309878
R22169 XThC.Tn[14].n38 XThC.Tn[14] 0.0309878
R22170 XThC.Tn[14].n41 XThC.Tn[14] 0.0309878
R22171 XThC.Tn[14].n44 XThC.Tn[14] 0.0309878
R22172 XThC.Tn[14].n47 XThC.Tn[14] 0.0309878
R22173 XThC.Tn[14].n50 XThC.Tn[14] 0.0309878
R22174 XThC.Tn[14].n53 XThC.Tn[14] 0.0309878
R22175 XThC.Tn[14].n56 XThC.Tn[14] 0.0309878
R22176 XThC.Tn[14].n12 XThC.Tn[14].n11 0.027939
R22177 XThC.Tn[14].n15 XThC.Tn[14].n14 0.027939
R22178 XThC.Tn[14].n18 XThC.Tn[14].n17 0.027939
R22179 XThC.Tn[14].n21 XThC.Tn[14].n20 0.027939
R22180 XThC.Tn[14].n24 XThC.Tn[14].n23 0.027939
R22181 XThC.Tn[14].n27 XThC.Tn[14].n26 0.027939
R22182 XThC.Tn[14].n30 XThC.Tn[14].n29 0.027939
R22183 XThC.Tn[14].n33 XThC.Tn[14].n32 0.027939
R22184 XThC.Tn[14].n36 XThC.Tn[14].n35 0.027939
R22185 XThC.Tn[14].n39 XThC.Tn[14].n38 0.027939
R22186 XThC.Tn[14].n42 XThC.Tn[14].n41 0.027939
R22187 XThC.Tn[14].n45 XThC.Tn[14].n44 0.027939
R22188 XThC.Tn[14].n48 XThC.Tn[14].n47 0.027939
R22189 XThC.Tn[14].n51 XThC.Tn[14].n50 0.027939
R22190 XThC.Tn[14].n54 XThC.Tn[14].n53 0.027939
R22191 XThC.Tn[14].n57 XThC.Tn[14].n56 0.027939
R22192 XThC.Tn[14].n58 XThC.Tn[14] 0.00250754
R22193 XThC.XTB1.Y.n6 XThC.XTB1.Y.t11 212.081
R22194 XThC.XTB1.Y.n5 XThC.XTB1.Y.t8 212.081
R22195 XThC.XTB1.Y.n11 XThC.XTB1.Y.t6 212.081
R22196 XThC.XTB1.Y.n3 XThC.XTB1.Y.t17 212.081
R22197 XThC.XTB1.Y.n15 XThC.XTB1.Y.t10 212.081
R22198 XThC.XTB1.Y.n16 XThC.XTB1.Y.t14 212.081
R22199 XThC.XTB1.Y.n18 XThC.XTB1.Y.t7 212.081
R22200 XThC.XTB1.Y.n14 XThC.XTB1.Y.t18 212.081
R22201 XThC.XTB1.Y.n22 XThC.XTB1.Y.n2 201.288
R22202 XThC.XTB1.Y.n8 XThC.XTB1.Y.n7 173.761
R22203 XThC.XTB1.Y.n17 XThC.XTB1.Y 158.656
R22204 XThC.XTB1.Y.n10 XThC.XTB1.Y.n9 152
R22205 XThC.XTB1.Y.n8 XThC.XTB1.Y.n4 152
R22206 XThC.XTB1.Y.n13 XThC.XTB1.Y.n12 152
R22207 XThC.XTB1.Y.n20 XThC.XTB1.Y.n19 152
R22208 XThC.XTB1.Y.n6 XThC.XTB1.Y.t16 139.78
R22209 XThC.XTB1.Y.n5 XThC.XTB1.Y.t13 139.78
R22210 XThC.XTB1.Y.n11 XThC.XTB1.Y.t12 139.78
R22211 XThC.XTB1.Y.n3 XThC.XTB1.Y.t5 139.78
R22212 XThC.XTB1.Y.n15 XThC.XTB1.Y.t4 139.78
R22213 XThC.XTB1.Y.n16 XThC.XTB1.Y.t3 139.78
R22214 XThC.XTB1.Y.n18 XThC.XTB1.Y.t15 139.78
R22215 XThC.XTB1.Y.n14 XThC.XTB1.Y.t9 139.78
R22216 XThC.XTB1.Y.n0 XThC.XTB1.Y.t1 132.067
R22217 XThC.XTB1.Y.n21 XThC.XTB1.Y 83.4676
R22218 XThC.XTB1.Y.n21 XThC.XTB1.Y.n13 61.4091
R22219 XThC.XTB1.Y.n16 XThC.XTB1.Y.n15 61.346
R22220 XThC.XTB1.Y.n10 XThC.XTB1.Y.n4 49.6611
R22221 XThC.XTB1.Y.n12 XThC.XTB1.Y.n11 45.2793
R22222 XThC.XTB1.Y.n7 XThC.XTB1.Y.n5 42.3581
R22223 XThC.XTB1.Y.n19 XThC.XTB1.Y.n14 30.6732
R22224 XThC.XTB1.Y.n19 XThC.XTB1.Y.n18 30.6732
R22225 XThC.XTB1.Y.n18 XThC.XTB1.Y.n17 30.6732
R22226 XThC.XTB1.Y.n17 XThC.XTB1.Y.n16 30.6732
R22227 XThC.XTB1.Y.n2 XThC.XTB1.Y.t0 26.5955
R22228 XThC.XTB1.Y.n2 XThC.XTB1.Y.t2 26.5955
R22229 XThC.XTB1.Y XThC.XTB1.Y.n22 23.489
R22230 XThC.XTB1.Y.n9 XThC.XTB1.Y.n8 21.7605
R22231 XThC.XTB1.Y.n7 XThC.XTB1.Y.n6 18.9884
R22232 XThC.XTB1.Y.n12 XThC.XTB1.Y.n3 16.0672
R22233 XThC.XTB1.Y.n20 XThC.XTB1.Y 14.8485
R22234 XThC.XTB1.Y.n13 XThC.XTB1.Y 11.5205
R22235 XThC.XTB1.Y.n22 XThC.XTB1.Y.n21 10.7939
R22236 XThC.XTB1.Y.n9 XThC.XTB1.Y 10.2405
R22237 XThC.XTB1.Y XThC.XTB1.Y.n20 8.7045
R22238 XThC.XTB1.Y.n5 XThC.XTB1.Y.n4 7.30353
R22239 XThC.XTB1.Y.n11 XThC.XTB1.Y.n10 4.38232
R22240 XThC.XTB1.Y.n1 XThC.XTB1.Y.n0 4.15748
R22241 XThC.XTB1.Y XThC.XTB1.Y.n1 3.76521
R22242 XThC.XTB1.Y.n0 XThC.XTB1.Y 1.17559
R22243 XThC.XTB1.Y.n1 XThC.XTB1.Y 0.921363
R22244 XThC.Tn[8].n5 XThC.Tn[8].n4 256.104
R22245 XThC.Tn[8].n8 XThC.Tn[8].n6 243.68
R22246 XThC.Tn[8].n2 XThC.Tn[8].n0 241.847
R22247 XThC.Tn[8].n8 XThC.Tn[8].n7 205.28
R22248 XThC.Tn[8].n5 XThC.Tn[8].n3 202.095
R22249 XThC.Tn[8].n2 XThC.Tn[8].n1 185
R22250 XThC.Tn[8].n12 XThC.Tn[8].n10 161.406
R22251 XThC.Tn[8].n15 XThC.Tn[8].n13 161.406
R22252 XThC.Tn[8].n18 XThC.Tn[8].n16 161.406
R22253 XThC.Tn[8].n21 XThC.Tn[8].n19 161.406
R22254 XThC.Tn[8].n24 XThC.Tn[8].n22 161.406
R22255 XThC.Tn[8].n27 XThC.Tn[8].n25 161.406
R22256 XThC.Tn[8].n30 XThC.Tn[8].n28 161.406
R22257 XThC.Tn[8].n33 XThC.Tn[8].n31 161.406
R22258 XThC.Tn[8].n36 XThC.Tn[8].n34 161.406
R22259 XThC.Tn[8].n39 XThC.Tn[8].n37 161.406
R22260 XThC.Tn[8].n42 XThC.Tn[8].n40 161.406
R22261 XThC.Tn[8].n45 XThC.Tn[8].n43 161.406
R22262 XThC.Tn[8].n48 XThC.Tn[8].n46 161.406
R22263 XThC.Tn[8].n51 XThC.Tn[8].n49 161.406
R22264 XThC.Tn[8].n54 XThC.Tn[8].n52 161.406
R22265 XThC.Tn[8].n57 XThC.Tn[8].n55 161.406
R22266 XThC.Tn[8].n10 XThC.Tn[8].t41 161.202
R22267 XThC.Tn[8].n13 XThC.Tn[8].t26 161.202
R22268 XThC.Tn[8].n16 XThC.Tn[8].t28 161.202
R22269 XThC.Tn[8].n19 XThC.Tn[8].t30 161.202
R22270 XThC.Tn[8].n22 XThC.Tn[8].t19 161.202
R22271 XThC.Tn[8].n25 XThC.Tn[8].t20 161.202
R22272 XThC.Tn[8].n28 XThC.Tn[8].t33 161.202
R22273 XThC.Tn[8].n31 XThC.Tn[8].t42 161.202
R22274 XThC.Tn[8].n34 XThC.Tn[8].t12 161.202
R22275 XThC.Tn[8].n37 XThC.Tn[8].t31 161.202
R22276 XThC.Tn[8].n40 XThC.Tn[8].t32 161.202
R22277 XThC.Tn[8].n43 XThC.Tn[8].t13 161.202
R22278 XThC.Tn[8].n46 XThC.Tn[8].t21 161.202
R22279 XThC.Tn[8].n49 XThC.Tn[8].t24 161.202
R22280 XThC.Tn[8].n52 XThC.Tn[8].t37 161.202
R22281 XThC.Tn[8].n55 XThC.Tn[8].t15 161.202
R22282 XThC.Tn[8].n10 XThC.Tn[8].t43 145.137
R22283 XThC.Tn[8].n13 XThC.Tn[8].t29 145.137
R22284 XThC.Tn[8].n16 XThC.Tn[8].t34 145.137
R22285 XThC.Tn[8].n19 XThC.Tn[8].t35 145.137
R22286 XThC.Tn[8].n22 XThC.Tn[8].t22 145.137
R22287 XThC.Tn[8].n25 XThC.Tn[8].t23 145.137
R22288 XThC.Tn[8].n28 XThC.Tn[8].t39 145.137
R22289 XThC.Tn[8].n31 XThC.Tn[8].t14 145.137
R22290 XThC.Tn[8].n34 XThC.Tn[8].t16 145.137
R22291 XThC.Tn[8].n37 XThC.Tn[8].t36 145.137
R22292 XThC.Tn[8].n40 XThC.Tn[8].t38 145.137
R22293 XThC.Tn[8].n43 XThC.Tn[8].t17 145.137
R22294 XThC.Tn[8].n46 XThC.Tn[8].t25 145.137
R22295 XThC.Tn[8].n49 XThC.Tn[8].t27 145.137
R22296 XThC.Tn[8].n52 XThC.Tn[8].t40 145.137
R22297 XThC.Tn[8].n55 XThC.Tn[8].t18 145.137
R22298 XThC.Tn[8].n3 XThC.Tn[8].t5 26.5955
R22299 XThC.Tn[8].n3 XThC.Tn[8].t6 26.5955
R22300 XThC.Tn[8].n4 XThC.Tn[8].t4 26.5955
R22301 XThC.Tn[8].n4 XThC.Tn[8].t7 26.5955
R22302 XThC.Tn[8].n6 XThC.Tn[8].t8 26.5955
R22303 XThC.Tn[8].n6 XThC.Tn[8].t11 26.5955
R22304 XThC.Tn[8].n7 XThC.Tn[8].t10 26.5955
R22305 XThC.Tn[8].n7 XThC.Tn[8].t9 26.5955
R22306 XThC.Tn[8].n0 XThC.Tn[8].t1 24.9236
R22307 XThC.Tn[8].n0 XThC.Tn[8].t0 24.9236
R22308 XThC.Tn[8].n1 XThC.Tn[8].t3 24.9236
R22309 XThC.Tn[8].n1 XThC.Tn[8].t2 24.9236
R22310 XThC.Tn[8] XThC.Tn[8].n8 22.9652
R22311 XThC.Tn[8] XThC.Tn[8].n2 22.9615
R22312 XThC.Tn[8].n9 XThC.Tn[8].n5 13.9299
R22313 XThC.Tn[8].n9 XThC.Tn[8] 13.9299
R22314 XThC.Tn[8].n60 XThC.Tn[8].n59 5.09639
R22315 XThC.Tn[8].n60 XThC.Tn[8].n9 2.99115
R22316 XThC.Tn[8].n9 XThC.Tn[8] 2.87153
R22317 XThC.Tn[8] XThC.Tn[8].n60 2.2734
R22318 XThC.Tn[8].n58 XThC.Tn[8] 1.14336
R22319 XThC.Tn[8].n15 XThC.Tn[8] 0.931056
R22320 XThC.Tn[8].n18 XThC.Tn[8] 0.931056
R22321 XThC.Tn[8].n21 XThC.Tn[8] 0.931056
R22322 XThC.Tn[8].n24 XThC.Tn[8] 0.931056
R22323 XThC.Tn[8].n27 XThC.Tn[8] 0.931056
R22324 XThC.Tn[8].n30 XThC.Tn[8] 0.931056
R22325 XThC.Tn[8].n33 XThC.Tn[8] 0.931056
R22326 XThC.Tn[8].n36 XThC.Tn[8] 0.931056
R22327 XThC.Tn[8].n39 XThC.Tn[8] 0.931056
R22328 XThC.Tn[8].n42 XThC.Tn[8] 0.931056
R22329 XThC.Tn[8].n45 XThC.Tn[8] 0.931056
R22330 XThC.Tn[8].n48 XThC.Tn[8] 0.931056
R22331 XThC.Tn[8].n51 XThC.Tn[8] 0.931056
R22332 XThC.Tn[8].n54 XThC.Tn[8] 0.931056
R22333 XThC.Tn[8].n57 XThC.Tn[8] 0.931056
R22334 XThC.Tn[8] XThC.Tn[8].n12 0.396333
R22335 XThC.Tn[8] XThC.Tn[8].n15 0.396333
R22336 XThC.Tn[8] XThC.Tn[8].n18 0.396333
R22337 XThC.Tn[8] XThC.Tn[8].n21 0.396333
R22338 XThC.Tn[8] XThC.Tn[8].n24 0.396333
R22339 XThC.Tn[8] XThC.Tn[8].n27 0.396333
R22340 XThC.Tn[8] XThC.Tn[8].n30 0.396333
R22341 XThC.Tn[8] XThC.Tn[8].n33 0.396333
R22342 XThC.Tn[8] XThC.Tn[8].n36 0.396333
R22343 XThC.Tn[8] XThC.Tn[8].n39 0.396333
R22344 XThC.Tn[8] XThC.Tn[8].n42 0.396333
R22345 XThC.Tn[8] XThC.Tn[8].n45 0.396333
R22346 XThC.Tn[8] XThC.Tn[8].n48 0.396333
R22347 XThC.Tn[8] XThC.Tn[8].n51 0.396333
R22348 XThC.Tn[8] XThC.Tn[8].n54 0.396333
R22349 XThC.Tn[8] XThC.Tn[8].n57 0.396333
R22350 XThC.Tn[8].n59 XThC.Tn[8].n58 0.166125
R22351 XThC.Tn[8].n11 XThC.Tn[8] 0.104667
R22352 XThC.Tn[8].n14 XThC.Tn[8] 0.104667
R22353 XThC.Tn[8].n17 XThC.Tn[8] 0.104667
R22354 XThC.Tn[8].n20 XThC.Tn[8] 0.104667
R22355 XThC.Tn[8].n23 XThC.Tn[8] 0.104667
R22356 XThC.Tn[8].n26 XThC.Tn[8] 0.104667
R22357 XThC.Tn[8].n29 XThC.Tn[8] 0.104667
R22358 XThC.Tn[8].n32 XThC.Tn[8] 0.104667
R22359 XThC.Tn[8].n35 XThC.Tn[8] 0.104667
R22360 XThC.Tn[8].n38 XThC.Tn[8] 0.104667
R22361 XThC.Tn[8].n41 XThC.Tn[8] 0.104667
R22362 XThC.Tn[8].n44 XThC.Tn[8] 0.104667
R22363 XThC.Tn[8].n47 XThC.Tn[8] 0.104667
R22364 XThC.Tn[8].n50 XThC.Tn[8] 0.104667
R22365 XThC.Tn[8].n53 XThC.Tn[8] 0.104667
R22366 XThC.Tn[8].n56 XThC.Tn[8] 0.104667
R22367 XThC.Tn[8].n59 XThC.Tn[8] 0.0389615
R22368 XThC.Tn[8].n58 XThC.Tn[8] 0.038
R22369 XThC.Tn[8].n11 XThC.Tn[8] 0.0309878
R22370 XThC.Tn[8].n14 XThC.Tn[8] 0.0309878
R22371 XThC.Tn[8].n17 XThC.Tn[8] 0.0309878
R22372 XThC.Tn[8].n20 XThC.Tn[8] 0.0309878
R22373 XThC.Tn[8].n23 XThC.Tn[8] 0.0309878
R22374 XThC.Tn[8].n26 XThC.Tn[8] 0.0309878
R22375 XThC.Tn[8].n29 XThC.Tn[8] 0.0309878
R22376 XThC.Tn[8].n32 XThC.Tn[8] 0.0309878
R22377 XThC.Tn[8].n35 XThC.Tn[8] 0.0309878
R22378 XThC.Tn[8].n38 XThC.Tn[8] 0.0309878
R22379 XThC.Tn[8].n41 XThC.Tn[8] 0.0309878
R22380 XThC.Tn[8].n44 XThC.Tn[8] 0.0309878
R22381 XThC.Tn[8].n47 XThC.Tn[8] 0.0309878
R22382 XThC.Tn[8].n50 XThC.Tn[8] 0.0309878
R22383 XThC.Tn[8].n53 XThC.Tn[8] 0.0309878
R22384 XThC.Tn[8].n56 XThC.Tn[8] 0.0309878
R22385 XThC.Tn[8].n12 XThC.Tn[8].n11 0.027939
R22386 XThC.Tn[8].n15 XThC.Tn[8].n14 0.027939
R22387 XThC.Tn[8].n18 XThC.Tn[8].n17 0.027939
R22388 XThC.Tn[8].n21 XThC.Tn[8].n20 0.027939
R22389 XThC.Tn[8].n24 XThC.Tn[8].n23 0.027939
R22390 XThC.Tn[8].n27 XThC.Tn[8].n26 0.027939
R22391 XThC.Tn[8].n30 XThC.Tn[8].n29 0.027939
R22392 XThC.Tn[8].n33 XThC.Tn[8].n32 0.027939
R22393 XThC.Tn[8].n36 XThC.Tn[8].n35 0.027939
R22394 XThC.Tn[8].n39 XThC.Tn[8].n38 0.027939
R22395 XThC.Tn[8].n42 XThC.Tn[8].n41 0.027939
R22396 XThC.Tn[8].n45 XThC.Tn[8].n44 0.027939
R22397 XThC.Tn[8].n48 XThC.Tn[8].n47 0.027939
R22398 XThC.Tn[8].n51 XThC.Tn[8].n50 0.027939
R22399 XThC.Tn[8].n54 XThC.Tn[8].n53 0.027939
R22400 XThC.Tn[8].n57 XThC.Tn[8].n56 0.027939
R22401 XThR.Tn[1].n2 XThR.Tn[1].n1 332.332
R22402 XThR.Tn[1].n2 XThR.Tn[1].n0 296.493
R22403 XThR.Tn[1] XThR.Tn[1].n82 161.363
R22404 XThR.Tn[1] XThR.Tn[1].n77 161.363
R22405 XThR.Tn[1] XThR.Tn[1].n72 161.363
R22406 XThR.Tn[1] XThR.Tn[1].n67 161.363
R22407 XThR.Tn[1] XThR.Tn[1].n62 161.363
R22408 XThR.Tn[1] XThR.Tn[1].n57 161.363
R22409 XThR.Tn[1] XThR.Tn[1].n52 161.363
R22410 XThR.Tn[1] XThR.Tn[1].n47 161.363
R22411 XThR.Tn[1] XThR.Tn[1].n42 161.363
R22412 XThR.Tn[1] XThR.Tn[1].n37 161.363
R22413 XThR.Tn[1] XThR.Tn[1].n32 161.363
R22414 XThR.Tn[1] XThR.Tn[1].n27 161.363
R22415 XThR.Tn[1] XThR.Tn[1].n22 161.363
R22416 XThR.Tn[1] XThR.Tn[1].n17 161.363
R22417 XThR.Tn[1] XThR.Tn[1].n12 161.363
R22418 XThR.Tn[1] XThR.Tn[1].n10 161.363
R22419 XThR.Tn[1].n84 XThR.Tn[1].n83 161.3
R22420 XThR.Tn[1].n79 XThR.Tn[1].n78 161.3
R22421 XThR.Tn[1].n74 XThR.Tn[1].n73 161.3
R22422 XThR.Tn[1].n69 XThR.Tn[1].n68 161.3
R22423 XThR.Tn[1].n64 XThR.Tn[1].n63 161.3
R22424 XThR.Tn[1].n59 XThR.Tn[1].n58 161.3
R22425 XThR.Tn[1].n54 XThR.Tn[1].n53 161.3
R22426 XThR.Tn[1].n49 XThR.Tn[1].n48 161.3
R22427 XThR.Tn[1].n44 XThR.Tn[1].n43 161.3
R22428 XThR.Tn[1].n39 XThR.Tn[1].n38 161.3
R22429 XThR.Tn[1].n34 XThR.Tn[1].n33 161.3
R22430 XThR.Tn[1].n29 XThR.Tn[1].n28 161.3
R22431 XThR.Tn[1].n24 XThR.Tn[1].n23 161.3
R22432 XThR.Tn[1].n19 XThR.Tn[1].n18 161.3
R22433 XThR.Tn[1].n14 XThR.Tn[1].n13 161.3
R22434 XThR.Tn[1].n82 XThR.Tn[1].t70 161.106
R22435 XThR.Tn[1].n77 XThR.Tn[1].t14 161.106
R22436 XThR.Tn[1].n72 XThR.Tn[1].t56 161.106
R22437 XThR.Tn[1].n67 XThR.Tn[1].t42 161.106
R22438 XThR.Tn[1].n62 XThR.Tn[1].t68 161.106
R22439 XThR.Tn[1].n57 XThR.Tn[1].t31 161.106
R22440 XThR.Tn[1].n52 XThR.Tn[1].t12 161.106
R22441 XThR.Tn[1].n47 XThR.Tn[1].t54 161.106
R22442 XThR.Tn[1].n42 XThR.Tn[1].t41 161.106
R22443 XThR.Tn[1].n37 XThR.Tn[1].t46 161.106
R22444 XThR.Tn[1].n32 XThR.Tn[1].t29 161.106
R22445 XThR.Tn[1].n27 XThR.Tn[1].t55 161.106
R22446 XThR.Tn[1].n22 XThR.Tn[1].t28 161.106
R22447 XThR.Tn[1].n17 XThR.Tn[1].t73 161.106
R22448 XThR.Tn[1].n12 XThR.Tn[1].t34 161.106
R22449 XThR.Tn[1].n10 XThR.Tn[1].t18 161.106
R22450 XThR.Tn[1].n83 XThR.Tn[1].t66 159.978
R22451 XThR.Tn[1].n78 XThR.Tn[1].t72 159.978
R22452 XThR.Tn[1].n73 XThR.Tn[1].t52 159.978
R22453 XThR.Tn[1].n68 XThR.Tn[1].t39 159.978
R22454 XThR.Tn[1].n63 XThR.Tn[1].t63 159.978
R22455 XThR.Tn[1].n58 XThR.Tn[1].t27 159.978
R22456 XThR.Tn[1].n53 XThR.Tn[1].t71 159.978
R22457 XThR.Tn[1].n48 XThR.Tn[1].t49 159.978
R22458 XThR.Tn[1].n43 XThR.Tn[1].t36 159.978
R22459 XThR.Tn[1].n38 XThR.Tn[1].t43 159.978
R22460 XThR.Tn[1].n33 XThR.Tn[1].t26 159.978
R22461 XThR.Tn[1].n28 XThR.Tn[1].t51 159.978
R22462 XThR.Tn[1].n23 XThR.Tn[1].t25 159.978
R22463 XThR.Tn[1].n18 XThR.Tn[1].t69 159.978
R22464 XThR.Tn[1].n13 XThR.Tn[1].t30 159.978
R22465 XThR.Tn[1].n82 XThR.Tn[1].t58 145.038
R22466 XThR.Tn[1].n77 XThR.Tn[1].t20 145.038
R22467 XThR.Tn[1].n72 XThR.Tn[1].t62 145.038
R22468 XThR.Tn[1].n67 XThR.Tn[1].t47 145.038
R22469 XThR.Tn[1].n62 XThR.Tn[1].t15 145.038
R22470 XThR.Tn[1].n57 XThR.Tn[1].t57 145.038
R22471 XThR.Tn[1].n52 XThR.Tn[1].t64 145.038
R22472 XThR.Tn[1].n47 XThR.Tn[1].t48 145.038
R22473 XThR.Tn[1].n42 XThR.Tn[1].t45 145.038
R22474 XThR.Tn[1].n37 XThR.Tn[1].t13 145.038
R22475 XThR.Tn[1].n32 XThR.Tn[1].t37 145.038
R22476 XThR.Tn[1].n27 XThR.Tn[1].t59 145.038
R22477 XThR.Tn[1].n22 XThR.Tn[1].t35 145.038
R22478 XThR.Tn[1].n17 XThR.Tn[1].t19 145.038
R22479 XThR.Tn[1].n12 XThR.Tn[1].t44 145.038
R22480 XThR.Tn[1].n10 XThR.Tn[1].t24 145.038
R22481 XThR.Tn[1].n83 XThR.Tn[1].t17 143.911
R22482 XThR.Tn[1].n78 XThR.Tn[1].t40 143.911
R22483 XThR.Tn[1].n73 XThR.Tn[1].t22 143.911
R22484 XThR.Tn[1].n68 XThR.Tn[1].t65 143.911
R22485 XThR.Tn[1].n63 XThR.Tn[1].t33 143.911
R22486 XThR.Tn[1].n58 XThR.Tn[1].t16 143.911
R22487 XThR.Tn[1].n53 XThR.Tn[1].t23 143.911
R22488 XThR.Tn[1].n48 XThR.Tn[1].t67 143.911
R22489 XThR.Tn[1].n43 XThR.Tn[1].t60 143.911
R22490 XThR.Tn[1].n38 XThR.Tn[1].t32 143.911
R22491 XThR.Tn[1].n33 XThR.Tn[1].t53 143.911
R22492 XThR.Tn[1].n28 XThR.Tn[1].t21 143.911
R22493 XThR.Tn[1].n23 XThR.Tn[1].t50 143.911
R22494 XThR.Tn[1].n18 XThR.Tn[1].t38 143.911
R22495 XThR.Tn[1].n13 XThR.Tn[1].t61 143.911
R22496 XThR.Tn[1].n7 XThR.Tn[1].n6 135.249
R22497 XThR.Tn[1].n9 XThR.Tn[1].n3 98.981
R22498 XThR.Tn[1].n8 XThR.Tn[1].n4 98.981
R22499 XThR.Tn[1].n7 XThR.Tn[1].n5 98.981
R22500 XThR.Tn[1].n9 XThR.Tn[1].n8 36.2672
R22501 XThR.Tn[1].n8 XThR.Tn[1].n7 36.2672
R22502 XThR.Tn[1].n88 XThR.Tn[1].n9 32.6405
R22503 XThR.Tn[1].n1 XThR.Tn[1].t7 26.5955
R22504 XThR.Tn[1].n1 XThR.Tn[1].t6 26.5955
R22505 XThR.Tn[1].n0 XThR.Tn[1].t4 26.5955
R22506 XThR.Tn[1].n0 XThR.Tn[1].t5 26.5955
R22507 XThR.Tn[1].n3 XThR.Tn[1].t11 24.9236
R22508 XThR.Tn[1].n3 XThR.Tn[1].t8 24.9236
R22509 XThR.Tn[1].n4 XThR.Tn[1].t10 24.9236
R22510 XThR.Tn[1].n4 XThR.Tn[1].t9 24.9236
R22511 XThR.Tn[1].n5 XThR.Tn[1].t2 24.9236
R22512 XThR.Tn[1].n5 XThR.Tn[1].t1 24.9236
R22513 XThR.Tn[1].n6 XThR.Tn[1].t3 24.9236
R22514 XThR.Tn[1].n6 XThR.Tn[1].t0 24.9236
R22515 XThR.Tn[1].n89 XThR.Tn[1].n2 18.5605
R22516 XThR.Tn[1].n89 XThR.Tn[1].n88 11.5205
R22517 XThR.Tn[1].n88 XThR.Tn[1] 6.42118
R22518 XThR.Tn[1] XThR.Tn[1].n11 5.34038
R22519 XThR.Tn[1].n16 XThR.Tn[1].n15 4.5005
R22520 XThR.Tn[1].n21 XThR.Tn[1].n20 4.5005
R22521 XThR.Tn[1].n26 XThR.Tn[1].n25 4.5005
R22522 XThR.Tn[1].n31 XThR.Tn[1].n30 4.5005
R22523 XThR.Tn[1].n36 XThR.Tn[1].n35 4.5005
R22524 XThR.Tn[1].n41 XThR.Tn[1].n40 4.5005
R22525 XThR.Tn[1].n46 XThR.Tn[1].n45 4.5005
R22526 XThR.Tn[1].n51 XThR.Tn[1].n50 4.5005
R22527 XThR.Tn[1].n56 XThR.Tn[1].n55 4.5005
R22528 XThR.Tn[1].n61 XThR.Tn[1].n60 4.5005
R22529 XThR.Tn[1].n66 XThR.Tn[1].n65 4.5005
R22530 XThR.Tn[1].n71 XThR.Tn[1].n70 4.5005
R22531 XThR.Tn[1].n76 XThR.Tn[1].n75 4.5005
R22532 XThR.Tn[1].n81 XThR.Tn[1].n80 4.5005
R22533 XThR.Tn[1].n86 XThR.Tn[1].n85 4.5005
R22534 XThR.Tn[1].n87 XThR.Tn[1] 3.70586
R22535 XThR.Tn[1].n16 XThR.Tn[1] 2.52282
R22536 XThR.Tn[1].n21 XThR.Tn[1] 2.52282
R22537 XThR.Tn[1].n26 XThR.Tn[1] 2.52282
R22538 XThR.Tn[1].n31 XThR.Tn[1] 2.52282
R22539 XThR.Tn[1].n36 XThR.Tn[1] 2.52282
R22540 XThR.Tn[1].n41 XThR.Tn[1] 2.52282
R22541 XThR.Tn[1].n46 XThR.Tn[1] 2.52282
R22542 XThR.Tn[1].n51 XThR.Tn[1] 2.52282
R22543 XThR.Tn[1].n56 XThR.Tn[1] 2.52282
R22544 XThR.Tn[1].n61 XThR.Tn[1] 2.52282
R22545 XThR.Tn[1].n66 XThR.Tn[1] 2.52282
R22546 XThR.Tn[1].n71 XThR.Tn[1] 2.52282
R22547 XThR.Tn[1].n76 XThR.Tn[1] 2.52282
R22548 XThR.Tn[1].n81 XThR.Tn[1] 2.52282
R22549 XThR.Tn[1].n86 XThR.Tn[1] 2.52282
R22550 XThR.Tn[1].n84 XThR.Tn[1] 1.08677
R22551 XThR.Tn[1].n79 XThR.Tn[1] 1.08677
R22552 XThR.Tn[1].n74 XThR.Tn[1] 1.08677
R22553 XThR.Tn[1].n69 XThR.Tn[1] 1.08677
R22554 XThR.Tn[1].n64 XThR.Tn[1] 1.08677
R22555 XThR.Tn[1].n59 XThR.Tn[1] 1.08677
R22556 XThR.Tn[1].n54 XThR.Tn[1] 1.08677
R22557 XThR.Tn[1].n49 XThR.Tn[1] 1.08677
R22558 XThR.Tn[1].n44 XThR.Tn[1] 1.08677
R22559 XThR.Tn[1].n39 XThR.Tn[1] 1.08677
R22560 XThR.Tn[1].n34 XThR.Tn[1] 1.08677
R22561 XThR.Tn[1].n29 XThR.Tn[1] 1.08677
R22562 XThR.Tn[1].n24 XThR.Tn[1] 1.08677
R22563 XThR.Tn[1].n19 XThR.Tn[1] 1.08677
R22564 XThR.Tn[1].n14 XThR.Tn[1] 1.08677
R22565 XThR.Tn[1] XThR.Tn[1].n16 0.839786
R22566 XThR.Tn[1] XThR.Tn[1].n21 0.839786
R22567 XThR.Tn[1] XThR.Tn[1].n26 0.839786
R22568 XThR.Tn[1] XThR.Tn[1].n31 0.839786
R22569 XThR.Tn[1] XThR.Tn[1].n36 0.839786
R22570 XThR.Tn[1] XThR.Tn[1].n41 0.839786
R22571 XThR.Tn[1] XThR.Tn[1].n46 0.839786
R22572 XThR.Tn[1] XThR.Tn[1].n51 0.839786
R22573 XThR.Tn[1] XThR.Tn[1].n56 0.839786
R22574 XThR.Tn[1] XThR.Tn[1].n61 0.839786
R22575 XThR.Tn[1] XThR.Tn[1].n66 0.839786
R22576 XThR.Tn[1] XThR.Tn[1].n71 0.839786
R22577 XThR.Tn[1] XThR.Tn[1].n76 0.839786
R22578 XThR.Tn[1] XThR.Tn[1].n81 0.839786
R22579 XThR.Tn[1] XThR.Tn[1].n86 0.839786
R22580 XThR.Tn[1] XThR.Tn[1].n89 0.6405
R22581 XThR.Tn[1].n11 XThR.Tn[1] 0.499542
R22582 XThR.Tn[1].n85 XThR.Tn[1] 0.063
R22583 XThR.Tn[1].n80 XThR.Tn[1] 0.063
R22584 XThR.Tn[1].n75 XThR.Tn[1] 0.063
R22585 XThR.Tn[1].n70 XThR.Tn[1] 0.063
R22586 XThR.Tn[1].n65 XThR.Tn[1] 0.063
R22587 XThR.Tn[1].n60 XThR.Tn[1] 0.063
R22588 XThR.Tn[1].n55 XThR.Tn[1] 0.063
R22589 XThR.Tn[1].n50 XThR.Tn[1] 0.063
R22590 XThR.Tn[1].n45 XThR.Tn[1] 0.063
R22591 XThR.Tn[1].n40 XThR.Tn[1] 0.063
R22592 XThR.Tn[1].n35 XThR.Tn[1] 0.063
R22593 XThR.Tn[1].n30 XThR.Tn[1] 0.063
R22594 XThR.Tn[1].n25 XThR.Tn[1] 0.063
R22595 XThR.Tn[1].n20 XThR.Tn[1] 0.063
R22596 XThR.Tn[1].n15 XThR.Tn[1] 0.063
R22597 XThR.Tn[1].n87 XThR.Tn[1] 0.0540714
R22598 XThR.Tn[1] XThR.Tn[1].n87 0.038
R22599 XThR.Tn[1].n11 XThR.Tn[1] 0.0143889
R22600 XThR.Tn[1].n85 XThR.Tn[1].n84 0.00771154
R22601 XThR.Tn[1].n80 XThR.Tn[1].n79 0.00771154
R22602 XThR.Tn[1].n75 XThR.Tn[1].n74 0.00771154
R22603 XThR.Tn[1].n70 XThR.Tn[1].n69 0.00771154
R22604 XThR.Tn[1].n65 XThR.Tn[1].n64 0.00771154
R22605 XThR.Tn[1].n60 XThR.Tn[1].n59 0.00771154
R22606 XThR.Tn[1].n55 XThR.Tn[1].n54 0.00771154
R22607 XThR.Tn[1].n50 XThR.Tn[1].n49 0.00771154
R22608 XThR.Tn[1].n45 XThR.Tn[1].n44 0.00771154
R22609 XThR.Tn[1].n40 XThR.Tn[1].n39 0.00771154
R22610 XThR.Tn[1].n35 XThR.Tn[1].n34 0.00771154
R22611 XThR.Tn[1].n30 XThR.Tn[1].n29 0.00771154
R22612 XThR.Tn[1].n25 XThR.Tn[1].n24 0.00771154
R22613 XThR.Tn[1].n20 XThR.Tn[1].n19 0.00771154
R22614 XThR.Tn[1].n15 XThR.Tn[1].n14 0.00771154
R22615 XThC.Tn[7].n2 XThC.Tn[7].n1 255.096
R22616 XThC.Tn[7].n55 XThC.Tn[7].n53 236.589
R22617 XThC.Tn[7].n2 XThC.Tn[7].n0 201.845
R22618 XThC.Tn[7].n55 XThC.Tn[7].n54 200.321
R22619 XThC.Tn[7].n5 XThC.Tn[7].n3 161.406
R22620 XThC.Tn[7].n8 XThC.Tn[7].n6 161.406
R22621 XThC.Tn[7].n11 XThC.Tn[7].n9 161.406
R22622 XThC.Tn[7].n14 XThC.Tn[7].n12 161.406
R22623 XThC.Tn[7].n17 XThC.Tn[7].n15 161.406
R22624 XThC.Tn[7].n20 XThC.Tn[7].n18 161.406
R22625 XThC.Tn[7].n23 XThC.Tn[7].n21 161.406
R22626 XThC.Tn[7].n26 XThC.Tn[7].n24 161.406
R22627 XThC.Tn[7].n29 XThC.Tn[7].n27 161.406
R22628 XThC.Tn[7].n32 XThC.Tn[7].n30 161.406
R22629 XThC.Tn[7].n35 XThC.Tn[7].n33 161.406
R22630 XThC.Tn[7].n38 XThC.Tn[7].n36 161.406
R22631 XThC.Tn[7].n41 XThC.Tn[7].n39 161.406
R22632 XThC.Tn[7].n44 XThC.Tn[7].n42 161.406
R22633 XThC.Tn[7].n47 XThC.Tn[7].n45 161.406
R22634 XThC.Tn[7].n50 XThC.Tn[7].n48 161.406
R22635 XThC.Tn[7].n3 XThC.Tn[7].t11 161.202
R22636 XThC.Tn[7].n6 XThC.Tn[7].t30 161.202
R22637 XThC.Tn[7].n9 XThC.Tn[7].t34 161.202
R22638 XThC.Tn[7].n12 XThC.Tn[7].t35 161.202
R22639 XThC.Tn[7].n15 XThC.Tn[7].t22 161.202
R22640 XThC.Tn[7].n18 XThC.Tn[7].t23 161.202
R22641 XThC.Tn[7].n21 XThC.Tn[7].t39 161.202
R22642 XThC.Tn[7].n24 XThC.Tn[7].t14 161.202
R22643 XThC.Tn[7].n27 XThC.Tn[7].t16 161.202
R22644 XThC.Tn[7].n30 XThC.Tn[7].t36 161.202
R22645 XThC.Tn[7].n33 XThC.Tn[7].t38 161.202
R22646 XThC.Tn[7].n36 XThC.Tn[7].t17 161.202
R22647 XThC.Tn[7].n39 XThC.Tn[7].t26 161.202
R22648 XThC.Tn[7].n42 XThC.Tn[7].t28 161.202
R22649 XThC.Tn[7].n45 XThC.Tn[7].t9 161.202
R22650 XThC.Tn[7].n48 XThC.Tn[7].t19 161.202
R22651 XThC.Tn[7].n3 XThC.Tn[7].t8 145.137
R22652 XThC.Tn[7].n6 XThC.Tn[7].t25 145.137
R22653 XThC.Tn[7].n9 XThC.Tn[7].t27 145.137
R22654 XThC.Tn[7].n12 XThC.Tn[7].t29 145.137
R22655 XThC.Tn[7].n15 XThC.Tn[7].t18 145.137
R22656 XThC.Tn[7].n18 XThC.Tn[7].t20 145.137
R22657 XThC.Tn[7].n21 XThC.Tn[7].t33 145.137
R22658 XThC.Tn[7].n24 XThC.Tn[7].t10 145.137
R22659 XThC.Tn[7].n27 XThC.Tn[7].t12 145.137
R22660 XThC.Tn[7].n30 XThC.Tn[7].t31 145.137
R22661 XThC.Tn[7].n33 XThC.Tn[7].t32 145.137
R22662 XThC.Tn[7].n36 XThC.Tn[7].t13 145.137
R22663 XThC.Tn[7].n39 XThC.Tn[7].t21 145.137
R22664 XThC.Tn[7].n42 XThC.Tn[7].t24 145.137
R22665 XThC.Tn[7].n45 XThC.Tn[7].t37 145.137
R22666 XThC.Tn[7].n48 XThC.Tn[7].t15 145.137
R22667 XThC.Tn[7].n0 XThC.Tn[7].t4 26.5955
R22668 XThC.Tn[7].n0 XThC.Tn[7].t7 26.5955
R22669 XThC.Tn[7].n1 XThC.Tn[7].t6 26.5955
R22670 XThC.Tn[7].n1 XThC.Tn[7].t5 26.5955
R22671 XThC.Tn[7] XThC.Tn[7].n2 26.5002
R22672 XThC.Tn[7].n53 XThC.Tn[7].t2 24.9236
R22673 XThC.Tn[7].n53 XThC.Tn[7].t1 24.9236
R22674 XThC.Tn[7].n54 XThC.Tn[7].t0 24.9236
R22675 XThC.Tn[7].n54 XThC.Tn[7].t3 24.9236
R22676 XThC.Tn[7].n56 XThC.Tn[7].n55 12.0894
R22677 XThC.Tn[7].n56 XThC.Tn[7] 9.64206
R22678 XThC.Tn[7].n52 XThC.Tn[7] 8.14595
R22679 XThC.Tn[7].n52 XThC.Tn[7].n51 3.36239
R22680 XThC.Tn[7] XThC.Tn[7].n52 3.15894
R22681 XThC.Tn[7].n51 XThC.Tn[7] 2.07622
R22682 XThC.Tn[7] XThC.Tn[7].n56 1.66284
R22683 XThC.Tn[7].n8 XThC.Tn[7] 0.931056
R22684 XThC.Tn[7].n11 XThC.Tn[7] 0.931056
R22685 XThC.Tn[7].n14 XThC.Tn[7] 0.931056
R22686 XThC.Tn[7].n17 XThC.Tn[7] 0.931056
R22687 XThC.Tn[7].n20 XThC.Tn[7] 0.931056
R22688 XThC.Tn[7].n23 XThC.Tn[7] 0.931056
R22689 XThC.Tn[7].n26 XThC.Tn[7] 0.931056
R22690 XThC.Tn[7].n29 XThC.Tn[7] 0.931056
R22691 XThC.Tn[7].n32 XThC.Tn[7] 0.931056
R22692 XThC.Tn[7].n35 XThC.Tn[7] 0.931056
R22693 XThC.Tn[7].n38 XThC.Tn[7] 0.931056
R22694 XThC.Tn[7].n41 XThC.Tn[7] 0.931056
R22695 XThC.Tn[7].n44 XThC.Tn[7] 0.931056
R22696 XThC.Tn[7].n47 XThC.Tn[7] 0.931056
R22697 XThC.Tn[7].n50 XThC.Tn[7] 0.931056
R22698 XThC.Tn[7] XThC.Tn[7].n5 0.396333
R22699 XThC.Tn[7] XThC.Tn[7].n8 0.396333
R22700 XThC.Tn[7] XThC.Tn[7].n11 0.396333
R22701 XThC.Tn[7] XThC.Tn[7].n14 0.396333
R22702 XThC.Tn[7] XThC.Tn[7].n17 0.396333
R22703 XThC.Tn[7] XThC.Tn[7].n20 0.396333
R22704 XThC.Tn[7] XThC.Tn[7].n23 0.396333
R22705 XThC.Tn[7] XThC.Tn[7].n26 0.396333
R22706 XThC.Tn[7] XThC.Tn[7].n29 0.396333
R22707 XThC.Tn[7] XThC.Tn[7].n32 0.396333
R22708 XThC.Tn[7] XThC.Tn[7].n35 0.396333
R22709 XThC.Tn[7] XThC.Tn[7].n38 0.396333
R22710 XThC.Tn[7] XThC.Tn[7].n41 0.396333
R22711 XThC.Tn[7] XThC.Tn[7].n44 0.396333
R22712 XThC.Tn[7] XThC.Tn[7].n47 0.396333
R22713 XThC.Tn[7] XThC.Tn[7].n50 0.396333
R22714 XThC.Tn[7].n4 XThC.Tn[7] 0.104667
R22715 XThC.Tn[7].n7 XThC.Tn[7] 0.104667
R22716 XThC.Tn[7].n10 XThC.Tn[7] 0.104667
R22717 XThC.Tn[7].n13 XThC.Tn[7] 0.104667
R22718 XThC.Tn[7].n16 XThC.Tn[7] 0.104667
R22719 XThC.Tn[7].n19 XThC.Tn[7] 0.104667
R22720 XThC.Tn[7].n22 XThC.Tn[7] 0.104667
R22721 XThC.Tn[7].n25 XThC.Tn[7] 0.104667
R22722 XThC.Tn[7].n28 XThC.Tn[7] 0.104667
R22723 XThC.Tn[7].n31 XThC.Tn[7] 0.104667
R22724 XThC.Tn[7].n34 XThC.Tn[7] 0.104667
R22725 XThC.Tn[7].n37 XThC.Tn[7] 0.104667
R22726 XThC.Tn[7].n40 XThC.Tn[7] 0.104667
R22727 XThC.Tn[7].n43 XThC.Tn[7] 0.104667
R22728 XThC.Tn[7].n46 XThC.Tn[7] 0.104667
R22729 XThC.Tn[7].n49 XThC.Tn[7] 0.104667
R22730 XThC.Tn[7].n4 XThC.Tn[7] 0.0309878
R22731 XThC.Tn[7].n7 XThC.Tn[7] 0.0309878
R22732 XThC.Tn[7].n10 XThC.Tn[7] 0.0309878
R22733 XThC.Tn[7].n13 XThC.Tn[7] 0.0309878
R22734 XThC.Tn[7].n16 XThC.Tn[7] 0.0309878
R22735 XThC.Tn[7].n19 XThC.Tn[7] 0.0309878
R22736 XThC.Tn[7].n22 XThC.Tn[7] 0.0309878
R22737 XThC.Tn[7].n25 XThC.Tn[7] 0.0309878
R22738 XThC.Tn[7].n28 XThC.Tn[7] 0.0309878
R22739 XThC.Tn[7].n31 XThC.Tn[7] 0.0309878
R22740 XThC.Tn[7].n34 XThC.Tn[7] 0.0309878
R22741 XThC.Tn[7].n37 XThC.Tn[7] 0.0309878
R22742 XThC.Tn[7].n40 XThC.Tn[7] 0.0309878
R22743 XThC.Tn[7].n43 XThC.Tn[7] 0.0309878
R22744 XThC.Tn[7].n46 XThC.Tn[7] 0.0309878
R22745 XThC.Tn[7].n49 XThC.Tn[7] 0.0309878
R22746 XThC.Tn[7].n5 XThC.Tn[7].n4 0.027939
R22747 XThC.Tn[7].n8 XThC.Tn[7].n7 0.027939
R22748 XThC.Tn[7].n11 XThC.Tn[7].n10 0.027939
R22749 XThC.Tn[7].n14 XThC.Tn[7].n13 0.027939
R22750 XThC.Tn[7].n17 XThC.Tn[7].n16 0.027939
R22751 XThC.Tn[7].n20 XThC.Tn[7].n19 0.027939
R22752 XThC.Tn[7].n23 XThC.Tn[7].n22 0.027939
R22753 XThC.Tn[7].n26 XThC.Tn[7].n25 0.027939
R22754 XThC.Tn[7].n29 XThC.Tn[7].n28 0.027939
R22755 XThC.Tn[7].n32 XThC.Tn[7].n31 0.027939
R22756 XThC.Tn[7].n35 XThC.Tn[7].n34 0.027939
R22757 XThC.Tn[7].n38 XThC.Tn[7].n37 0.027939
R22758 XThC.Tn[7].n41 XThC.Tn[7].n40 0.027939
R22759 XThC.Tn[7].n44 XThC.Tn[7].n43 0.027939
R22760 XThC.Tn[7].n47 XThC.Tn[7].n46 0.027939
R22761 XThC.Tn[7].n50 XThC.Tn[7].n49 0.027939
R22762 XThC.Tn[7].n51 XThC.Tn[7] 0.00240908
R22763 XThR.Tn[4].n2 XThR.Tn[4].n1 332.332
R22764 XThR.Tn[4].n2 XThR.Tn[4].n0 296.493
R22765 XThR.Tn[4] XThR.Tn[4].n82 161.363
R22766 XThR.Tn[4] XThR.Tn[4].n77 161.363
R22767 XThR.Tn[4] XThR.Tn[4].n72 161.363
R22768 XThR.Tn[4] XThR.Tn[4].n67 161.363
R22769 XThR.Tn[4] XThR.Tn[4].n62 161.363
R22770 XThR.Tn[4] XThR.Tn[4].n57 161.363
R22771 XThR.Tn[4] XThR.Tn[4].n52 161.363
R22772 XThR.Tn[4] XThR.Tn[4].n47 161.363
R22773 XThR.Tn[4] XThR.Tn[4].n42 161.363
R22774 XThR.Tn[4] XThR.Tn[4].n37 161.363
R22775 XThR.Tn[4] XThR.Tn[4].n32 161.363
R22776 XThR.Tn[4] XThR.Tn[4].n27 161.363
R22777 XThR.Tn[4] XThR.Tn[4].n22 161.363
R22778 XThR.Tn[4] XThR.Tn[4].n17 161.363
R22779 XThR.Tn[4] XThR.Tn[4].n12 161.363
R22780 XThR.Tn[4] XThR.Tn[4].n10 161.363
R22781 XThR.Tn[4].n84 XThR.Tn[4].n83 161.3
R22782 XThR.Tn[4].n79 XThR.Tn[4].n78 161.3
R22783 XThR.Tn[4].n74 XThR.Tn[4].n73 161.3
R22784 XThR.Tn[4].n69 XThR.Tn[4].n68 161.3
R22785 XThR.Tn[4].n64 XThR.Tn[4].n63 161.3
R22786 XThR.Tn[4].n59 XThR.Tn[4].n58 161.3
R22787 XThR.Tn[4].n54 XThR.Tn[4].n53 161.3
R22788 XThR.Tn[4].n49 XThR.Tn[4].n48 161.3
R22789 XThR.Tn[4].n44 XThR.Tn[4].n43 161.3
R22790 XThR.Tn[4].n39 XThR.Tn[4].n38 161.3
R22791 XThR.Tn[4].n34 XThR.Tn[4].n33 161.3
R22792 XThR.Tn[4].n29 XThR.Tn[4].n28 161.3
R22793 XThR.Tn[4].n24 XThR.Tn[4].n23 161.3
R22794 XThR.Tn[4].n19 XThR.Tn[4].n18 161.3
R22795 XThR.Tn[4].n14 XThR.Tn[4].n13 161.3
R22796 XThR.Tn[4].n82 XThR.Tn[4].t28 161.106
R22797 XThR.Tn[4].n77 XThR.Tn[4].t34 161.106
R22798 XThR.Tn[4].n72 XThR.Tn[4].t14 161.106
R22799 XThR.Tn[4].n67 XThR.Tn[4].t62 161.106
R22800 XThR.Tn[4].n62 XThR.Tn[4].t26 161.106
R22801 XThR.Tn[4].n57 XThR.Tn[4].t51 161.106
R22802 XThR.Tn[4].n52 XThR.Tn[4].t32 161.106
R22803 XThR.Tn[4].n47 XThR.Tn[4].t12 161.106
R22804 XThR.Tn[4].n42 XThR.Tn[4].t61 161.106
R22805 XThR.Tn[4].n37 XThR.Tn[4].t66 161.106
R22806 XThR.Tn[4].n32 XThR.Tn[4].t49 161.106
R22807 XThR.Tn[4].n27 XThR.Tn[4].t13 161.106
R22808 XThR.Tn[4].n22 XThR.Tn[4].t48 161.106
R22809 XThR.Tn[4].n17 XThR.Tn[4].t31 161.106
R22810 XThR.Tn[4].n12 XThR.Tn[4].t54 161.106
R22811 XThR.Tn[4].n10 XThR.Tn[4].t38 161.106
R22812 XThR.Tn[4].n83 XThR.Tn[4].t24 159.978
R22813 XThR.Tn[4].n78 XThR.Tn[4].t30 159.978
R22814 XThR.Tn[4].n73 XThR.Tn[4].t72 159.978
R22815 XThR.Tn[4].n68 XThR.Tn[4].t59 159.978
R22816 XThR.Tn[4].n63 XThR.Tn[4].t21 159.978
R22817 XThR.Tn[4].n58 XThR.Tn[4].t47 159.978
R22818 XThR.Tn[4].n53 XThR.Tn[4].t29 159.978
R22819 XThR.Tn[4].n48 XThR.Tn[4].t69 159.978
R22820 XThR.Tn[4].n43 XThR.Tn[4].t56 159.978
R22821 XThR.Tn[4].n38 XThR.Tn[4].t63 159.978
R22822 XThR.Tn[4].n33 XThR.Tn[4].t46 159.978
R22823 XThR.Tn[4].n28 XThR.Tn[4].t71 159.978
R22824 XThR.Tn[4].n23 XThR.Tn[4].t45 159.978
R22825 XThR.Tn[4].n18 XThR.Tn[4].t27 159.978
R22826 XThR.Tn[4].n13 XThR.Tn[4].t50 159.978
R22827 XThR.Tn[4].n82 XThR.Tn[4].t16 145.038
R22828 XThR.Tn[4].n77 XThR.Tn[4].t40 145.038
R22829 XThR.Tn[4].n72 XThR.Tn[4].t20 145.038
R22830 XThR.Tn[4].n67 XThR.Tn[4].t67 145.038
R22831 XThR.Tn[4].n62 XThR.Tn[4].t35 145.038
R22832 XThR.Tn[4].n57 XThR.Tn[4].t15 145.038
R22833 XThR.Tn[4].n52 XThR.Tn[4].t22 145.038
R22834 XThR.Tn[4].n47 XThR.Tn[4].t68 145.038
R22835 XThR.Tn[4].n42 XThR.Tn[4].t64 145.038
R22836 XThR.Tn[4].n37 XThR.Tn[4].t33 145.038
R22837 XThR.Tn[4].n32 XThR.Tn[4].t57 145.038
R22838 XThR.Tn[4].n27 XThR.Tn[4].t17 145.038
R22839 XThR.Tn[4].n22 XThR.Tn[4].t55 145.038
R22840 XThR.Tn[4].n17 XThR.Tn[4].t39 145.038
R22841 XThR.Tn[4].n12 XThR.Tn[4].t65 145.038
R22842 XThR.Tn[4].n10 XThR.Tn[4].t44 145.038
R22843 XThR.Tn[4].n83 XThR.Tn[4].t37 143.911
R22844 XThR.Tn[4].n78 XThR.Tn[4].t60 143.911
R22845 XThR.Tn[4].n73 XThR.Tn[4].t42 143.911
R22846 XThR.Tn[4].n68 XThR.Tn[4].t23 143.911
R22847 XThR.Tn[4].n63 XThR.Tn[4].t53 143.911
R22848 XThR.Tn[4].n58 XThR.Tn[4].t36 143.911
R22849 XThR.Tn[4].n53 XThR.Tn[4].t43 143.911
R22850 XThR.Tn[4].n48 XThR.Tn[4].t25 143.911
R22851 XThR.Tn[4].n43 XThR.Tn[4].t18 143.911
R22852 XThR.Tn[4].n38 XThR.Tn[4].t52 143.911
R22853 XThR.Tn[4].n33 XThR.Tn[4].t73 143.911
R22854 XThR.Tn[4].n28 XThR.Tn[4].t41 143.911
R22855 XThR.Tn[4].n23 XThR.Tn[4].t70 143.911
R22856 XThR.Tn[4].n18 XThR.Tn[4].t58 143.911
R22857 XThR.Tn[4].n13 XThR.Tn[4].t19 143.911
R22858 XThR.Tn[4].n7 XThR.Tn[4].n5 135.249
R22859 XThR.Tn[4].n9 XThR.Tn[4].n3 98.982
R22860 XThR.Tn[4].n8 XThR.Tn[4].n4 98.982
R22861 XThR.Tn[4].n7 XThR.Tn[4].n6 98.982
R22862 XThR.Tn[4].n9 XThR.Tn[4].n8 36.2672
R22863 XThR.Tn[4].n8 XThR.Tn[4].n7 36.2672
R22864 XThR.Tn[4].n88 XThR.Tn[4].n9 32.6405
R22865 XThR.Tn[4].n1 XThR.Tn[4].t4 26.5955
R22866 XThR.Tn[4].n1 XThR.Tn[4].t7 26.5955
R22867 XThR.Tn[4].n0 XThR.Tn[4].t5 26.5955
R22868 XThR.Tn[4].n0 XThR.Tn[4].t6 26.5955
R22869 XThR.Tn[4].n3 XThR.Tn[4].t11 24.9236
R22870 XThR.Tn[4].n3 XThR.Tn[4].t8 24.9236
R22871 XThR.Tn[4].n4 XThR.Tn[4].t10 24.9236
R22872 XThR.Tn[4].n4 XThR.Tn[4].t9 24.9236
R22873 XThR.Tn[4].n5 XThR.Tn[4].t0 24.9236
R22874 XThR.Tn[4].n5 XThR.Tn[4].t1 24.9236
R22875 XThR.Tn[4].n6 XThR.Tn[4].t3 24.9236
R22876 XThR.Tn[4].n6 XThR.Tn[4].t2 24.9236
R22877 XThR.Tn[4] XThR.Tn[4].n2 23.3605
R22878 XThR.Tn[4] XThR.Tn[4].n88 6.7205
R22879 XThR.Tn[4].n88 XThR.Tn[4] 5.80883
R22880 XThR.Tn[4] XThR.Tn[4].n11 5.34038
R22881 XThR.Tn[4].n16 XThR.Tn[4].n15 4.5005
R22882 XThR.Tn[4].n21 XThR.Tn[4].n20 4.5005
R22883 XThR.Tn[4].n26 XThR.Tn[4].n25 4.5005
R22884 XThR.Tn[4].n31 XThR.Tn[4].n30 4.5005
R22885 XThR.Tn[4].n36 XThR.Tn[4].n35 4.5005
R22886 XThR.Tn[4].n41 XThR.Tn[4].n40 4.5005
R22887 XThR.Tn[4].n46 XThR.Tn[4].n45 4.5005
R22888 XThR.Tn[4].n51 XThR.Tn[4].n50 4.5005
R22889 XThR.Tn[4].n56 XThR.Tn[4].n55 4.5005
R22890 XThR.Tn[4].n61 XThR.Tn[4].n60 4.5005
R22891 XThR.Tn[4].n66 XThR.Tn[4].n65 4.5005
R22892 XThR.Tn[4].n71 XThR.Tn[4].n70 4.5005
R22893 XThR.Tn[4].n76 XThR.Tn[4].n75 4.5005
R22894 XThR.Tn[4].n81 XThR.Tn[4].n80 4.5005
R22895 XThR.Tn[4].n86 XThR.Tn[4].n85 4.5005
R22896 XThR.Tn[4].n87 XThR.Tn[4] 3.70586
R22897 XThR.Tn[4].n16 XThR.Tn[4] 2.52282
R22898 XThR.Tn[4].n21 XThR.Tn[4] 2.52282
R22899 XThR.Tn[4].n26 XThR.Tn[4] 2.52282
R22900 XThR.Tn[4].n31 XThR.Tn[4] 2.52282
R22901 XThR.Tn[4].n36 XThR.Tn[4] 2.52282
R22902 XThR.Tn[4].n41 XThR.Tn[4] 2.52282
R22903 XThR.Tn[4].n46 XThR.Tn[4] 2.52282
R22904 XThR.Tn[4].n51 XThR.Tn[4] 2.52282
R22905 XThR.Tn[4].n56 XThR.Tn[4] 2.52282
R22906 XThR.Tn[4].n61 XThR.Tn[4] 2.52282
R22907 XThR.Tn[4].n66 XThR.Tn[4] 2.52282
R22908 XThR.Tn[4].n71 XThR.Tn[4] 2.52282
R22909 XThR.Tn[4].n76 XThR.Tn[4] 2.52282
R22910 XThR.Tn[4].n81 XThR.Tn[4] 2.52282
R22911 XThR.Tn[4].n86 XThR.Tn[4] 2.52282
R22912 XThR.Tn[4].n84 XThR.Tn[4] 1.08677
R22913 XThR.Tn[4].n79 XThR.Tn[4] 1.08677
R22914 XThR.Tn[4].n74 XThR.Tn[4] 1.08677
R22915 XThR.Tn[4].n69 XThR.Tn[4] 1.08677
R22916 XThR.Tn[4].n64 XThR.Tn[4] 1.08677
R22917 XThR.Tn[4].n59 XThR.Tn[4] 1.08677
R22918 XThR.Tn[4].n54 XThR.Tn[4] 1.08677
R22919 XThR.Tn[4].n49 XThR.Tn[4] 1.08677
R22920 XThR.Tn[4].n44 XThR.Tn[4] 1.08677
R22921 XThR.Tn[4].n39 XThR.Tn[4] 1.08677
R22922 XThR.Tn[4].n34 XThR.Tn[4] 1.08677
R22923 XThR.Tn[4].n29 XThR.Tn[4] 1.08677
R22924 XThR.Tn[4].n24 XThR.Tn[4] 1.08677
R22925 XThR.Tn[4].n19 XThR.Tn[4] 1.08677
R22926 XThR.Tn[4].n14 XThR.Tn[4] 1.08677
R22927 XThR.Tn[4] XThR.Tn[4].n16 0.839786
R22928 XThR.Tn[4] XThR.Tn[4].n21 0.839786
R22929 XThR.Tn[4] XThR.Tn[4].n26 0.839786
R22930 XThR.Tn[4] XThR.Tn[4].n31 0.839786
R22931 XThR.Tn[4] XThR.Tn[4].n36 0.839786
R22932 XThR.Tn[4] XThR.Tn[4].n41 0.839786
R22933 XThR.Tn[4] XThR.Tn[4].n46 0.839786
R22934 XThR.Tn[4] XThR.Tn[4].n51 0.839786
R22935 XThR.Tn[4] XThR.Tn[4].n56 0.839786
R22936 XThR.Tn[4] XThR.Tn[4].n61 0.839786
R22937 XThR.Tn[4] XThR.Tn[4].n66 0.839786
R22938 XThR.Tn[4] XThR.Tn[4].n71 0.839786
R22939 XThR.Tn[4] XThR.Tn[4].n76 0.839786
R22940 XThR.Tn[4] XThR.Tn[4].n81 0.839786
R22941 XThR.Tn[4] XThR.Tn[4].n86 0.839786
R22942 XThR.Tn[4].n11 XThR.Tn[4] 0.499542
R22943 XThR.Tn[4].n85 XThR.Tn[4] 0.063
R22944 XThR.Tn[4].n80 XThR.Tn[4] 0.063
R22945 XThR.Tn[4].n75 XThR.Tn[4] 0.063
R22946 XThR.Tn[4].n70 XThR.Tn[4] 0.063
R22947 XThR.Tn[4].n65 XThR.Tn[4] 0.063
R22948 XThR.Tn[4].n60 XThR.Tn[4] 0.063
R22949 XThR.Tn[4].n55 XThR.Tn[4] 0.063
R22950 XThR.Tn[4].n50 XThR.Tn[4] 0.063
R22951 XThR.Tn[4].n45 XThR.Tn[4] 0.063
R22952 XThR.Tn[4].n40 XThR.Tn[4] 0.063
R22953 XThR.Tn[4].n35 XThR.Tn[4] 0.063
R22954 XThR.Tn[4].n30 XThR.Tn[4] 0.063
R22955 XThR.Tn[4].n25 XThR.Tn[4] 0.063
R22956 XThR.Tn[4].n20 XThR.Tn[4] 0.063
R22957 XThR.Tn[4].n15 XThR.Tn[4] 0.063
R22958 XThR.Tn[4].n87 XThR.Tn[4] 0.0540714
R22959 XThR.Tn[4] XThR.Tn[4].n87 0.038
R22960 XThR.Tn[4].n11 XThR.Tn[4] 0.0143889
R22961 XThR.Tn[4].n85 XThR.Tn[4].n84 0.00771154
R22962 XThR.Tn[4].n80 XThR.Tn[4].n79 0.00771154
R22963 XThR.Tn[4].n75 XThR.Tn[4].n74 0.00771154
R22964 XThR.Tn[4].n70 XThR.Tn[4].n69 0.00771154
R22965 XThR.Tn[4].n65 XThR.Tn[4].n64 0.00771154
R22966 XThR.Tn[4].n60 XThR.Tn[4].n59 0.00771154
R22967 XThR.Tn[4].n55 XThR.Tn[4].n54 0.00771154
R22968 XThR.Tn[4].n50 XThR.Tn[4].n49 0.00771154
R22969 XThR.Tn[4].n45 XThR.Tn[4].n44 0.00771154
R22970 XThR.Tn[4].n40 XThR.Tn[4].n39 0.00771154
R22971 XThR.Tn[4].n35 XThR.Tn[4].n34 0.00771154
R22972 XThR.Tn[4].n30 XThR.Tn[4].n29 0.00771154
R22973 XThR.Tn[4].n25 XThR.Tn[4].n24 0.00771154
R22974 XThR.Tn[4].n20 XThR.Tn[4].n19 0.00771154
R22975 XThR.Tn[4].n15 XThR.Tn[4].n14 0.00771154
R22976 XThR.Tn[11].n8 XThR.Tn[11].n7 256.104
R22977 XThR.Tn[11].n5 XThR.Tn[11].n3 243.68
R22978 XThR.Tn[11].n2 XThR.Tn[11].n1 241.847
R22979 XThR.Tn[11].n5 XThR.Tn[11].n4 205.28
R22980 XThR.Tn[11].n8 XThR.Tn[11].n6 202.094
R22981 XThR.Tn[11].n2 XThR.Tn[11].n0 185
R22982 XThR.Tn[11] XThR.Tn[11].n82 161.363
R22983 XThR.Tn[11] XThR.Tn[11].n77 161.363
R22984 XThR.Tn[11] XThR.Tn[11].n72 161.363
R22985 XThR.Tn[11] XThR.Tn[11].n67 161.363
R22986 XThR.Tn[11] XThR.Tn[11].n62 161.363
R22987 XThR.Tn[11] XThR.Tn[11].n57 161.363
R22988 XThR.Tn[11] XThR.Tn[11].n52 161.363
R22989 XThR.Tn[11] XThR.Tn[11].n47 161.363
R22990 XThR.Tn[11] XThR.Tn[11].n42 161.363
R22991 XThR.Tn[11] XThR.Tn[11].n37 161.363
R22992 XThR.Tn[11] XThR.Tn[11].n32 161.363
R22993 XThR.Tn[11] XThR.Tn[11].n27 161.363
R22994 XThR.Tn[11] XThR.Tn[11].n22 161.363
R22995 XThR.Tn[11] XThR.Tn[11].n17 161.363
R22996 XThR.Tn[11] XThR.Tn[11].n12 161.363
R22997 XThR.Tn[11] XThR.Tn[11].n10 161.363
R22998 XThR.Tn[11].n84 XThR.Tn[11].n83 161.3
R22999 XThR.Tn[11].n79 XThR.Tn[11].n78 161.3
R23000 XThR.Tn[11].n74 XThR.Tn[11].n73 161.3
R23001 XThR.Tn[11].n69 XThR.Tn[11].n68 161.3
R23002 XThR.Tn[11].n64 XThR.Tn[11].n63 161.3
R23003 XThR.Tn[11].n59 XThR.Tn[11].n58 161.3
R23004 XThR.Tn[11].n54 XThR.Tn[11].n53 161.3
R23005 XThR.Tn[11].n49 XThR.Tn[11].n48 161.3
R23006 XThR.Tn[11].n44 XThR.Tn[11].n43 161.3
R23007 XThR.Tn[11].n39 XThR.Tn[11].n38 161.3
R23008 XThR.Tn[11].n34 XThR.Tn[11].n33 161.3
R23009 XThR.Tn[11].n29 XThR.Tn[11].n28 161.3
R23010 XThR.Tn[11].n24 XThR.Tn[11].n23 161.3
R23011 XThR.Tn[11].n19 XThR.Tn[11].n18 161.3
R23012 XThR.Tn[11].n14 XThR.Tn[11].n13 161.3
R23013 XThR.Tn[11].n82 XThR.Tn[11].t40 161.106
R23014 XThR.Tn[11].n77 XThR.Tn[11].t46 161.106
R23015 XThR.Tn[11].n72 XThR.Tn[11].t24 161.106
R23016 XThR.Tn[11].n67 XThR.Tn[11].t73 161.106
R23017 XThR.Tn[11].n62 XThR.Tn[11].t39 161.106
R23018 XThR.Tn[11].n57 XThR.Tn[11].t63 161.106
R23019 XThR.Tn[11].n52 XThR.Tn[11].t43 161.106
R23020 XThR.Tn[11].n47 XThR.Tn[11].t22 161.106
R23021 XThR.Tn[11].n42 XThR.Tn[11].t71 161.106
R23022 XThR.Tn[11].n37 XThR.Tn[11].t14 161.106
R23023 XThR.Tn[11].n32 XThR.Tn[11].t62 161.106
R23024 XThR.Tn[11].n27 XThR.Tn[11].t23 161.106
R23025 XThR.Tn[11].n22 XThR.Tn[11].t60 161.106
R23026 XThR.Tn[11].n17 XThR.Tn[11].t41 161.106
R23027 XThR.Tn[11].n12 XThR.Tn[11].t67 161.106
R23028 XThR.Tn[11].n10 XThR.Tn[11].t48 161.106
R23029 XThR.Tn[11].n83 XThR.Tn[11].t31 159.978
R23030 XThR.Tn[11].n78 XThR.Tn[11].t38 159.978
R23031 XThR.Tn[11].n73 XThR.Tn[11].t20 159.978
R23032 XThR.Tn[11].n68 XThR.Tn[11].t66 159.978
R23033 XThR.Tn[11].n63 XThR.Tn[11].t29 159.978
R23034 XThR.Tn[11].n58 XThR.Tn[11].t57 159.978
R23035 XThR.Tn[11].n53 XThR.Tn[11].t37 159.978
R23036 XThR.Tn[11].n48 XThR.Tn[11].t17 159.978
R23037 XThR.Tn[11].n43 XThR.Tn[11].t64 159.978
R23038 XThR.Tn[11].n38 XThR.Tn[11].t72 159.978
R23039 XThR.Tn[11].n33 XThR.Tn[11].t55 159.978
R23040 XThR.Tn[11].n28 XThR.Tn[11].t19 159.978
R23041 XThR.Tn[11].n23 XThR.Tn[11].t54 159.978
R23042 XThR.Tn[11].n18 XThR.Tn[11].t36 159.978
R23043 XThR.Tn[11].n13 XThR.Tn[11].t58 159.978
R23044 XThR.Tn[11].n82 XThR.Tn[11].t26 145.038
R23045 XThR.Tn[11].n77 XThR.Tn[11].t53 145.038
R23046 XThR.Tn[11].n72 XThR.Tn[11].t34 145.038
R23047 XThR.Tn[11].n67 XThR.Tn[11].t15 145.038
R23048 XThR.Tn[11].n62 XThR.Tn[11].t47 145.038
R23049 XThR.Tn[11].n57 XThR.Tn[11].t25 145.038
R23050 XThR.Tn[11].n52 XThR.Tn[11].t35 145.038
R23051 XThR.Tn[11].n47 XThR.Tn[11].t16 145.038
R23052 XThR.Tn[11].n42 XThR.Tn[11].t13 145.038
R23053 XThR.Tn[11].n37 XThR.Tn[11].t44 145.038
R23054 XThR.Tn[11].n32 XThR.Tn[11].t70 145.038
R23055 XThR.Tn[11].n27 XThR.Tn[11].t33 145.038
R23056 XThR.Tn[11].n22 XThR.Tn[11].t68 145.038
R23057 XThR.Tn[11].n17 XThR.Tn[11].t49 145.038
R23058 XThR.Tn[11].n12 XThR.Tn[11].t12 145.038
R23059 XThR.Tn[11].n10 XThR.Tn[11].t56 145.038
R23060 XThR.Tn[11].n83 XThR.Tn[11].t45 143.911
R23061 XThR.Tn[11].n78 XThR.Tn[11].t69 143.911
R23062 XThR.Tn[11].n73 XThR.Tn[11].t51 143.911
R23063 XThR.Tn[11].n68 XThR.Tn[11].t30 143.911
R23064 XThR.Tn[11].n63 XThR.Tn[11].t61 143.911
R23065 XThR.Tn[11].n58 XThR.Tn[11].t42 143.911
R23066 XThR.Tn[11].n53 XThR.Tn[11].t52 143.911
R23067 XThR.Tn[11].n48 XThR.Tn[11].t32 143.911
R23068 XThR.Tn[11].n43 XThR.Tn[11].t28 143.911
R23069 XThR.Tn[11].n38 XThR.Tn[11].t59 143.911
R23070 XThR.Tn[11].n33 XThR.Tn[11].t21 143.911
R23071 XThR.Tn[11].n28 XThR.Tn[11].t50 143.911
R23072 XThR.Tn[11].n23 XThR.Tn[11].t18 143.911
R23073 XThR.Tn[11].n18 XThR.Tn[11].t65 143.911
R23074 XThR.Tn[11].n13 XThR.Tn[11].t27 143.911
R23075 XThR.Tn[11] XThR.Tn[11].n5 35.7652
R23076 XThR.Tn[11].n6 XThR.Tn[11].t4 26.5955
R23077 XThR.Tn[11].n6 XThR.Tn[11].t6 26.5955
R23078 XThR.Tn[11].n7 XThR.Tn[11].t5 26.5955
R23079 XThR.Tn[11].n7 XThR.Tn[11].t7 26.5955
R23080 XThR.Tn[11].n3 XThR.Tn[11].t8 26.5955
R23081 XThR.Tn[11].n3 XThR.Tn[11].t10 26.5955
R23082 XThR.Tn[11].n4 XThR.Tn[11].t9 26.5955
R23083 XThR.Tn[11].n4 XThR.Tn[11].t11 26.5955
R23084 XThR.Tn[11].n0 XThR.Tn[11].t2 24.9236
R23085 XThR.Tn[11].n0 XThR.Tn[11].t0 24.9236
R23086 XThR.Tn[11].n1 XThR.Tn[11].t3 24.9236
R23087 XThR.Tn[11].n1 XThR.Tn[11].t1 24.9236
R23088 XThR.Tn[11] XThR.Tn[11].n2 22.9615
R23089 XThR.Tn[11].n9 XThR.Tn[11].n8 13.5534
R23090 XThR.Tn[11].n88 XThR.Tn[11] 8.41462
R23091 XThR.Tn[11] XThR.Tn[11].n11 5.34038
R23092 XThR.Tn[11].n16 XThR.Tn[11].n15 4.5005
R23093 XThR.Tn[11].n21 XThR.Tn[11].n20 4.5005
R23094 XThR.Tn[11].n26 XThR.Tn[11].n25 4.5005
R23095 XThR.Tn[11].n31 XThR.Tn[11].n30 4.5005
R23096 XThR.Tn[11].n36 XThR.Tn[11].n35 4.5005
R23097 XThR.Tn[11].n41 XThR.Tn[11].n40 4.5005
R23098 XThR.Tn[11].n46 XThR.Tn[11].n45 4.5005
R23099 XThR.Tn[11].n51 XThR.Tn[11].n50 4.5005
R23100 XThR.Tn[11].n56 XThR.Tn[11].n55 4.5005
R23101 XThR.Tn[11].n61 XThR.Tn[11].n60 4.5005
R23102 XThR.Tn[11].n66 XThR.Tn[11].n65 4.5005
R23103 XThR.Tn[11].n71 XThR.Tn[11].n70 4.5005
R23104 XThR.Tn[11].n76 XThR.Tn[11].n75 4.5005
R23105 XThR.Tn[11].n81 XThR.Tn[11].n80 4.5005
R23106 XThR.Tn[11].n86 XThR.Tn[11].n85 4.5005
R23107 XThR.Tn[11].n87 XThR.Tn[11] 3.70586
R23108 XThR.Tn[11].n88 XThR.Tn[11].n9 2.99115
R23109 XThR.Tn[11].n9 XThR.Tn[11] 2.87153
R23110 XThR.Tn[11].n16 XThR.Tn[11] 2.52282
R23111 XThR.Tn[11].n21 XThR.Tn[11] 2.52282
R23112 XThR.Tn[11].n26 XThR.Tn[11] 2.52282
R23113 XThR.Tn[11].n31 XThR.Tn[11] 2.52282
R23114 XThR.Tn[11].n36 XThR.Tn[11] 2.52282
R23115 XThR.Tn[11].n41 XThR.Tn[11] 2.52282
R23116 XThR.Tn[11].n46 XThR.Tn[11] 2.52282
R23117 XThR.Tn[11].n51 XThR.Tn[11] 2.52282
R23118 XThR.Tn[11].n56 XThR.Tn[11] 2.52282
R23119 XThR.Tn[11].n61 XThR.Tn[11] 2.52282
R23120 XThR.Tn[11].n66 XThR.Tn[11] 2.52282
R23121 XThR.Tn[11].n71 XThR.Tn[11] 2.52282
R23122 XThR.Tn[11].n76 XThR.Tn[11] 2.52282
R23123 XThR.Tn[11].n81 XThR.Tn[11] 2.52282
R23124 XThR.Tn[11].n86 XThR.Tn[11] 2.52282
R23125 XThR.Tn[11] XThR.Tn[11].n88 2.2734
R23126 XThR.Tn[11].n9 XThR.Tn[11] 1.50638
R23127 XThR.Tn[11].n84 XThR.Tn[11] 1.08677
R23128 XThR.Tn[11].n79 XThR.Tn[11] 1.08677
R23129 XThR.Tn[11].n74 XThR.Tn[11] 1.08677
R23130 XThR.Tn[11].n69 XThR.Tn[11] 1.08677
R23131 XThR.Tn[11].n64 XThR.Tn[11] 1.08677
R23132 XThR.Tn[11].n59 XThR.Tn[11] 1.08677
R23133 XThR.Tn[11].n54 XThR.Tn[11] 1.08677
R23134 XThR.Tn[11].n49 XThR.Tn[11] 1.08677
R23135 XThR.Tn[11].n44 XThR.Tn[11] 1.08677
R23136 XThR.Tn[11].n39 XThR.Tn[11] 1.08677
R23137 XThR.Tn[11].n34 XThR.Tn[11] 1.08677
R23138 XThR.Tn[11].n29 XThR.Tn[11] 1.08677
R23139 XThR.Tn[11].n24 XThR.Tn[11] 1.08677
R23140 XThR.Tn[11].n19 XThR.Tn[11] 1.08677
R23141 XThR.Tn[11].n14 XThR.Tn[11] 1.08677
R23142 XThR.Tn[11] XThR.Tn[11].n16 0.839786
R23143 XThR.Tn[11] XThR.Tn[11].n21 0.839786
R23144 XThR.Tn[11] XThR.Tn[11].n26 0.839786
R23145 XThR.Tn[11] XThR.Tn[11].n31 0.839786
R23146 XThR.Tn[11] XThR.Tn[11].n36 0.839786
R23147 XThR.Tn[11] XThR.Tn[11].n41 0.839786
R23148 XThR.Tn[11] XThR.Tn[11].n46 0.839786
R23149 XThR.Tn[11] XThR.Tn[11].n51 0.839786
R23150 XThR.Tn[11] XThR.Tn[11].n56 0.839786
R23151 XThR.Tn[11] XThR.Tn[11].n61 0.839786
R23152 XThR.Tn[11] XThR.Tn[11].n66 0.839786
R23153 XThR.Tn[11] XThR.Tn[11].n71 0.839786
R23154 XThR.Tn[11] XThR.Tn[11].n76 0.839786
R23155 XThR.Tn[11] XThR.Tn[11].n81 0.839786
R23156 XThR.Tn[11] XThR.Tn[11].n86 0.839786
R23157 XThR.Tn[11].n11 XThR.Tn[11] 0.499542
R23158 XThR.Tn[11].n85 XThR.Tn[11] 0.063
R23159 XThR.Tn[11].n80 XThR.Tn[11] 0.063
R23160 XThR.Tn[11].n75 XThR.Tn[11] 0.063
R23161 XThR.Tn[11].n70 XThR.Tn[11] 0.063
R23162 XThR.Tn[11].n65 XThR.Tn[11] 0.063
R23163 XThR.Tn[11].n60 XThR.Tn[11] 0.063
R23164 XThR.Tn[11].n55 XThR.Tn[11] 0.063
R23165 XThR.Tn[11].n50 XThR.Tn[11] 0.063
R23166 XThR.Tn[11].n45 XThR.Tn[11] 0.063
R23167 XThR.Tn[11].n40 XThR.Tn[11] 0.063
R23168 XThR.Tn[11].n35 XThR.Tn[11] 0.063
R23169 XThR.Tn[11].n30 XThR.Tn[11] 0.063
R23170 XThR.Tn[11].n25 XThR.Tn[11] 0.063
R23171 XThR.Tn[11].n20 XThR.Tn[11] 0.063
R23172 XThR.Tn[11].n15 XThR.Tn[11] 0.063
R23173 XThR.Tn[11].n87 XThR.Tn[11] 0.0540714
R23174 XThR.Tn[11] XThR.Tn[11].n87 0.038
R23175 XThR.Tn[11].n11 XThR.Tn[11] 0.0143889
R23176 XThR.Tn[11].n85 XThR.Tn[11].n84 0.00771154
R23177 XThR.Tn[11].n80 XThR.Tn[11].n79 0.00771154
R23178 XThR.Tn[11].n75 XThR.Tn[11].n74 0.00771154
R23179 XThR.Tn[11].n70 XThR.Tn[11].n69 0.00771154
R23180 XThR.Tn[11].n65 XThR.Tn[11].n64 0.00771154
R23181 XThR.Tn[11].n60 XThR.Tn[11].n59 0.00771154
R23182 XThR.Tn[11].n55 XThR.Tn[11].n54 0.00771154
R23183 XThR.Tn[11].n50 XThR.Tn[11].n49 0.00771154
R23184 XThR.Tn[11].n45 XThR.Tn[11].n44 0.00771154
R23185 XThR.Tn[11].n40 XThR.Tn[11].n39 0.00771154
R23186 XThR.Tn[11].n35 XThR.Tn[11].n34 0.00771154
R23187 XThR.Tn[11].n30 XThR.Tn[11].n29 0.00771154
R23188 XThR.Tn[11].n25 XThR.Tn[11].n24 0.00771154
R23189 XThR.Tn[11].n20 XThR.Tn[11].n19 0.00771154
R23190 XThR.Tn[11].n15 XThR.Tn[11].n14 0.00771154
R23191 XThR.Tn[7].n5 XThR.Tn[7].n3 244.069
R23192 XThR.Tn[7].n2 XThR.Tn[7].n1 236.589
R23193 XThR.Tn[7].n5 XThR.Tn[7].n4 204.893
R23194 XThR.Tn[7].n2 XThR.Tn[7].n0 200.321
R23195 XThR.Tn[7] XThR.Tn[7].n79 161.363
R23196 XThR.Tn[7] XThR.Tn[7].n74 161.363
R23197 XThR.Tn[7] XThR.Tn[7].n69 161.363
R23198 XThR.Tn[7] XThR.Tn[7].n64 161.363
R23199 XThR.Tn[7] XThR.Tn[7].n59 161.363
R23200 XThR.Tn[7] XThR.Tn[7].n54 161.363
R23201 XThR.Tn[7] XThR.Tn[7].n49 161.363
R23202 XThR.Tn[7] XThR.Tn[7].n44 161.363
R23203 XThR.Tn[7] XThR.Tn[7].n39 161.363
R23204 XThR.Tn[7] XThR.Tn[7].n34 161.363
R23205 XThR.Tn[7] XThR.Tn[7].n29 161.363
R23206 XThR.Tn[7] XThR.Tn[7].n24 161.363
R23207 XThR.Tn[7] XThR.Tn[7].n19 161.363
R23208 XThR.Tn[7] XThR.Tn[7].n14 161.363
R23209 XThR.Tn[7] XThR.Tn[7].n9 161.363
R23210 XThR.Tn[7] XThR.Tn[7].n7 161.363
R23211 XThR.Tn[7].n81 XThR.Tn[7].n80 161.3
R23212 XThR.Tn[7].n76 XThR.Tn[7].n75 161.3
R23213 XThR.Tn[7].n71 XThR.Tn[7].n70 161.3
R23214 XThR.Tn[7].n66 XThR.Tn[7].n65 161.3
R23215 XThR.Tn[7].n61 XThR.Tn[7].n60 161.3
R23216 XThR.Tn[7].n56 XThR.Tn[7].n55 161.3
R23217 XThR.Tn[7].n51 XThR.Tn[7].n50 161.3
R23218 XThR.Tn[7].n46 XThR.Tn[7].n45 161.3
R23219 XThR.Tn[7].n41 XThR.Tn[7].n40 161.3
R23220 XThR.Tn[7].n36 XThR.Tn[7].n35 161.3
R23221 XThR.Tn[7].n31 XThR.Tn[7].n30 161.3
R23222 XThR.Tn[7].n26 XThR.Tn[7].n25 161.3
R23223 XThR.Tn[7].n21 XThR.Tn[7].n20 161.3
R23224 XThR.Tn[7].n16 XThR.Tn[7].n15 161.3
R23225 XThR.Tn[7].n11 XThR.Tn[7].n10 161.3
R23226 XThR.Tn[7].n79 XThR.Tn[7].t35 161.106
R23227 XThR.Tn[7].n74 XThR.Tn[7].t41 161.106
R23228 XThR.Tn[7].n69 XThR.Tn[7].t22 161.106
R23229 XThR.Tn[7].n64 XThR.Tn[7].t69 161.106
R23230 XThR.Tn[7].n59 XThR.Tn[7].t33 161.106
R23231 XThR.Tn[7].n54 XThR.Tn[7].t57 161.106
R23232 XThR.Tn[7].n49 XThR.Tn[7].t39 161.106
R23233 XThR.Tn[7].n44 XThR.Tn[7].t20 161.106
R23234 XThR.Tn[7].n39 XThR.Tn[7].t68 161.106
R23235 XThR.Tn[7].n34 XThR.Tn[7].t11 161.106
R23236 XThR.Tn[7].n29 XThR.Tn[7].t56 161.106
R23237 XThR.Tn[7].n24 XThR.Tn[7].t21 161.106
R23238 XThR.Tn[7].n19 XThR.Tn[7].t55 161.106
R23239 XThR.Tn[7].n14 XThR.Tn[7].t37 161.106
R23240 XThR.Tn[7].n9 XThR.Tn[7].t60 161.106
R23241 XThR.Tn[7].n7 XThR.Tn[7].t45 161.106
R23242 XThR.Tn[7].n80 XThR.Tn[7].t13 159.978
R23243 XThR.Tn[7].n75 XThR.Tn[7].t17 159.978
R23244 XThR.Tn[7].n70 XThR.Tn[7].t64 159.978
R23245 XThR.Tn[7].n65 XThR.Tn[7].t48 159.978
R23246 XThR.Tn[7].n60 XThR.Tn[7].t10 159.978
R23247 XThR.Tn[7].n55 XThR.Tn[7].t36 159.978
R23248 XThR.Tn[7].n50 XThR.Tn[7].t16 159.978
R23249 XThR.Tn[7].n45 XThR.Tn[7].t61 159.978
R23250 XThR.Tn[7].n40 XThR.Tn[7].t46 159.978
R23251 XThR.Tn[7].n35 XThR.Tn[7].t54 159.978
R23252 XThR.Tn[7].n30 XThR.Tn[7].t34 159.978
R23253 XThR.Tn[7].n25 XThR.Tn[7].t63 159.978
R23254 XThR.Tn[7].n20 XThR.Tn[7].t32 159.978
R23255 XThR.Tn[7].n15 XThR.Tn[7].t15 159.978
R23256 XThR.Tn[7].n10 XThR.Tn[7].t38 159.978
R23257 XThR.Tn[7].n79 XThR.Tn[7].t24 145.038
R23258 XThR.Tn[7].n74 XThR.Tn[7].t49 145.038
R23259 XThR.Tn[7].n69 XThR.Tn[7].t28 145.038
R23260 XThR.Tn[7].n64 XThR.Tn[7].t12 145.038
R23261 XThR.Tn[7].n59 XThR.Tn[7].t42 145.038
R23262 XThR.Tn[7].n54 XThR.Tn[7].t23 145.038
R23263 XThR.Tn[7].n49 XThR.Tn[7].t29 145.038
R23264 XThR.Tn[7].n44 XThR.Tn[7].t14 145.038
R23265 XThR.Tn[7].n39 XThR.Tn[7].t9 145.038
R23266 XThR.Tn[7].n34 XThR.Tn[7].t40 145.038
R23267 XThR.Tn[7].n29 XThR.Tn[7].t65 145.038
R23268 XThR.Tn[7].n24 XThR.Tn[7].t25 145.038
R23269 XThR.Tn[7].n19 XThR.Tn[7].t62 145.038
R23270 XThR.Tn[7].n14 XThR.Tn[7].t47 145.038
R23271 XThR.Tn[7].n9 XThR.Tn[7].t8 145.038
R23272 XThR.Tn[7].n7 XThR.Tn[7].t53 145.038
R23273 XThR.Tn[7].n80 XThR.Tn[7].t44 143.911
R23274 XThR.Tn[7].n75 XThR.Tn[7].t67 143.911
R23275 XThR.Tn[7].n70 XThR.Tn[7].t51 143.911
R23276 XThR.Tn[7].n65 XThR.Tn[7].t30 143.911
R23277 XThR.Tn[7].n60 XThR.Tn[7].t59 143.911
R23278 XThR.Tn[7].n55 XThR.Tn[7].t43 143.911
R23279 XThR.Tn[7].n50 XThR.Tn[7].t52 143.911
R23280 XThR.Tn[7].n45 XThR.Tn[7].t31 143.911
R23281 XThR.Tn[7].n40 XThR.Tn[7].t27 143.911
R23282 XThR.Tn[7].n35 XThR.Tn[7].t58 143.911
R23283 XThR.Tn[7].n30 XThR.Tn[7].t19 143.911
R23284 XThR.Tn[7].n25 XThR.Tn[7].t50 143.911
R23285 XThR.Tn[7].n20 XThR.Tn[7].t18 143.911
R23286 XThR.Tn[7].n15 XThR.Tn[7].t66 143.911
R23287 XThR.Tn[7].n10 XThR.Tn[7].t26 143.911
R23288 XThR.Tn[7].n4 XThR.Tn[7].t5 26.5955
R23289 XThR.Tn[7].n4 XThR.Tn[7].t4 26.5955
R23290 XThR.Tn[7].n3 XThR.Tn[7].t6 26.5955
R23291 XThR.Tn[7].n3 XThR.Tn[7].t7 26.5955
R23292 XThR.Tn[7].n0 XThR.Tn[7].t2 24.9236
R23293 XThR.Tn[7].n0 XThR.Tn[7].t1 24.9236
R23294 XThR.Tn[7].n1 XThR.Tn[7].t3 24.9236
R23295 XThR.Tn[7].n1 XThR.Tn[7].t0 24.9236
R23296 XThR.Tn[7] XThR.Tn[7].n2 16.079
R23297 XThR.Tn[7].n6 XThR.Tn[7].n5 11.4531
R23298 XThR.Tn[7] XThR.Tn[7].n6 10.4732
R23299 XThR.Tn[7] XThR.Tn[7].n85 8.81089
R23300 XThR.Tn[7] XThR.Tn[7].n8 5.34038
R23301 XThR.Tn[7].n85 XThR.Tn[7] 5.25732
R23302 XThR.Tn[7].n13 XThR.Tn[7].n12 4.5005
R23303 XThR.Tn[7].n18 XThR.Tn[7].n17 4.5005
R23304 XThR.Tn[7].n23 XThR.Tn[7].n22 4.5005
R23305 XThR.Tn[7].n28 XThR.Tn[7].n27 4.5005
R23306 XThR.Tn[7].n33 XThR.Tn[7].n32 4.5005
R23307 XThR.Tn[7].n38 XThR.Tn[7].n37 4.5005
R23308 XThR.Tn[7].n43 XThR.Tn[7].n42 4.5005
R23309 XThR.Tn[7].n48 XThR.Tn[7].n47 4.5005
R23310 XThR.Tn[7].n53 XThR.Tn[7].n52 4.5005
R23311 XThR.Tn[7].n58 XThR.Tn[7].n57 4.5005
R23312 XThR.Tn[7].n63 XThR.Tn[7].n62 4.5005
R23313 XThR.Tn[7].n68 XThR.Tn[7].n67 4.5005
R23314 XThR.Tn[7].n73 XThR.Tn[7].n72 4.5005
R23315 XThR.Tn[7].n78 XThR.Tn[7].n77 4.5005
R23316 XThR.Tn[7].n83 XThR.Tn[7].n82 4.5005
R23317 XThR.Tn[7].n84 XThR.Tn[7] 3.70586
R23318 XThR.Tn[7].n13 XThR.Tn[7] 2.52282
R23319 XThR.Tn[7].n18 XThR.Tn[7] 2.52282
R23320 XThR.Tn[7].n23 XThR.Tn[7] 2.52282
R23321 XThR.Tn[7].n28 XThR.Tn[7] 2.52282
R23322 XThR.Tn[7].n33 XThR.Tn[7] 2.52282
R23323 XThR.Tn[7].n38 XThR.Tn[7] 2.52282
R23324 XThR.Tn[7].n43 XThR.Tn[7] 2.52282
R23325 XThR.Tn[7].n48 XThR.Tn[7] 2.52282
R23326 XThR.Tn[7].n53 XThR.Tn[7] 2.52282
R23327 XThR.Tn[7].n58 XThR.Tn[7] 2.52282
R23328 XThR.Tn[7].n63 XThR.Tn[7] 2.52282
R23329 XThR.Tn[7].n68 XThR.Tn[7] 2.52282
R23330 XThR.Tn[7].n73 XThR.Tn[7] 2.52282
R23331 XThR.Tn[7].n78 XThR.Tn[7] 2.52282
R23332 XThR.Tn[7].n83 XThR.Tn[7] 2.52282
R23333 XThR.Tn[7].n85 XThR.Tn[7] 2.49401
R23334 XThR.Tn[7].n81 XThR.Tn[7] 1.08677
R23335 XThR.Tn[7].n76 XThR.Tn[7] 1.08677
R23336 XThR.Tn[7].n71 XThR.Tn[7] 1.08677
R23337 XThR.Tn[7].n66 XThR.Tn[7] 1.08677
R23338 XThR.Tn[7].n61 XThR.Tn[7] 1.08677
R23339 XThR.Tn[7].n56 XThR.Tn[7] 1.08677
R23340 XThR.Tn[7].n51 XThR.Tn[7] 1.08677
R23341 XThR.Tn[7].n46 XThR.Tn[7] 1.08677
R23342 XThR.Tn[7].n41 XThR.Tn[7] 1.08677
R23343 XThR.Tn[7].n36 XThR.Tn[7] 1.08677
R23344 XThR.Tn[7].n31 XThR.Tn[7] 1.08677
R23345 XThR.Tn[7].n26 XThR.Tn[7] 1.08677
R23346 XThR.Tn[7].n21 XThR.Tn[7] 1.08677
R23347 XThR.Tn[7].n16 XThR.Tn[7] 1.08677
R23348 XThR.Tn[7].n11 XThR.Tn[7] 1.08677
R23349 XThR.Tn[7] XThR.Tn[7].n13 0.839786
R23350 XThR.Tn[7] XThR.Tn[7].n18 0.839786
R23351 XThR.Tn[7] XThR.Tn[7].n23 0.839786
R23352 XThR.Tn[7] XThR.Tn[7].n28 0.839786
R23353 XThR.Tn[7] XThR.Tn[7].n33 0.839786
R23354 XThR.Tn[7] XThR.Tn[7].n38 0.839786
R23355 XThR.Tn[7] XThR.Tn[7].n43 0.839786
R23356 XThR.Tn[7] XThR.Tn[7].n48 0.839786
R23357 XThR.Tn[7] XThR.Tn[7].n53 0.839786
R23358 XThR.Tn[7] XThR.Tn[7].n58 0.839786
R23359 XThR.Tn[7] XThR.Tn[7].n63 0.839786
R23360 XThR.Tn[7] XThR.Tn[7].n68 0.839786
R23361 XThR.Tn[7] XThR.Tn[7].n73 0.839786
R23362 XThR.Tn[7] XThR.Tn[7].n78 0.839786
R23363 XThR.Tn[7] XThR.Tn[7].n83 0.839786
R23364 XThR.Tn[7].n6 XThR.Tn[7] 0.829611
R23365 XThR.Tn[7].n8 XThR.Tn[7] 0.499542
R23366 XThR.Tn[7].n82 XThR.Tn[7] 0.063
R23367 XThR.Tn[7].n77 XThR.Tn[7] 0.063
R23368 XThR.Tn[7].n72 XThR.Tn[7] 0.063
R23369 XThR.Tn[7].n67 XThR.Tn[7] 0.063
R23370 XThR.Tn[7].n62 XThR.Tn[7] 0.063
R23371 XThR.Tn[7].n57 XThR.Tn[7] 0.063
R23372 XThR.Tn[7].n52 XThR.Tn[7] 0.063
R23373 XThR.Tn[7].n47 XThR.Tn[7] 0.063
R23374 XThR.Tn[7].n42 XThR.Tn[7] 0.063
R23375 XThR.Tn[7].n37 XThR.Tn[7] 0.063
R23376 XThR.Tn[7].n32 XThR.Tn[7] 0.063
R23377 XThR.Tn[7].n27 XThR.Tn[7] 0.063
R23378 XThR.Tn[7].n22 XThR.Tn[7] 0.063
R23379 XThR.Tn[7].n17 XThR.Tn[7] 0.063
R23380 XThR.Tn[7].n12 XThR.Tn[7] 0.063
R23381 XThR.Tn[7].n84 XThR.Tn[7] 0.0540714
R23382 XThR.Tn[7] XThR.Tn[7].n84 0.038
R23383 XThR.Tn[7].n8 XThR.Tn[7] 0.0143889
R23384 XThR.Tn[7].n82 XThR.Tn[7].n81 0.00771154
R23385 XThR.Tn[7].n77 XThR.Tn[7].n76 0.00771154
R23386 XThR.Tn[7].n72 XThR.Tn[7].n71 0.00771154
R23387 XThR.Tn[7].n67 XThR.Tn[7].n66 0.00771154
R23388 XThR.Tn[7].n62 XThR.Tn[7].n61 0.00771154
R23389 XThR.Tn[7].n57 XThR.Tn[7].n56 0.00771154
R23390 XThR.Tn[7].n52 XThR.Tn[7].n51 0.00771154
R23391 XThR.Tn[7].n47 XThR.Tn[7].n46 0.00771154
R23392 XThR.Tn[7].n42 XThR.Tn[7].n41 0.00771154
R23393 XThR.Tn[7].n37 XThR.Tn[7].n36 0.00771154
R23394 XThR.Tn[7].n32 XThR.Tn[7].n31 0.00771154
R23395 XThR.Tn[7].n27 XThR.Tn[7].n26 0.00771154
R23396 XThR.Tn[7].n22 XThR.Tn[7].n21 0.00771154
R23397 XThR.Tn[7].n17 XThR.Tn[7].n16 0.00771154
R23398 XThR.Tn[7].n12 XThR.Tn[7].n11 0.00771154
R23399 XThR.Tn[0].n2 XThR.Tn[0].n1 332.332
R23400 XThR.Tn[0].n2 XThR.Tn[0].n0 296.493
R23401 XThR.Tn[0] XThR.Tn[0].n82 161.363
R23402 XThR.Tn[0] XThR.Tn[0].n77 161.363
R23403 XThR.Tn[0] XThR.Tn[0].n72 161.363
R23404 XThR.Tn[0] XThR.Tn[0].n67 161.363
R23405 XThR.Tn[0] XThR.Tn[0].n62 161.363
R23406 XThR.Tn[0] XThR.Tn[0].n57 161.363
R23407 XThR.Tn[0] XThR.Tn[0].n52 161.363
R23408 XThR.Tn[0] XThR.Tn[0].n47 161.363
R23409 XThR.Tn[0] XThR.Tn[0].n42 161.363
R23410 XThR.Tn[0] XThR.Tn[0].n37 161.363
R23411 XThR.Tn[0] XThR.Tn[0].n32 161.363
R23412 XThR.Tn[0] XThR.Tn[0].n27 161.363
R23413 XThR.Tn[0] XThR.Tn[0].n22 161.363
R23414 XThR.Tn[0] XThR.Tn[0].n17 161.363
R23415 XThR.Tn[0] XThR.Tn[0].n12 161.363
R23416 XThR.Tn[0] XThR.Tn[0].n10 161.363
R23417 XThR.Tn[0].n84 XThR.Tn[0].n83 161.3
R23418 XThR.Tn[0].n79 XThR.Tn[0].n78 161.3
R23419 XThR.Tn[0].n74 XThR.Tn[0].n73 161.3
R23420 XThR.Tn[0].n69 XThR.Tn[0].n68 161.3
R23421 XThR.Tn[0].n64 XThR.Tn[0].n63 161.3
R23422 XThR.Tn[0].n59 XThR.Tn[0].n58 161.3
R23423 XThR.Tn[0].n54 XThR.Tn[0].n53 161.3
R23424 XThR.Tn[0].n49 XThR.Tn[0].n48 161.3
R23425 XThR.Tn[0].n44 XThR.Tn[0].n43 161.3
R23426 XThR.Tn[0].n39 XThR.Tn[0].n38 161.3
R23427 XThR.Tn[0].n34 XThR.Tn[0].n33 161.3
R23428 XThR.Tn[0].n29 XThR.Tn[0].n28 161.3
R23429 XThR.Tn[0].n24 XThR.Tn[0].n23 161.3
R23430 XThR.Tn[0].n19 XThR.Tn[0].n18 161.3
R23431 XThR.Tn[0].n14 XThR.Tn[0].n13 161.3
R23432 XThR.Tn[0].n82 XThR.Tn[0].t32 161.106
R23433 XThR.Tn[0].n77 XThR.Tn[0].t36 161.106
R23434 XThR.Tn[0].n72 XThR.Tn[0].t16 161.106
R23435 XThR.Tn[0].n67 XThR.Tn[0].t65 161.106
R23436 XThR.Tn[0].n62 XThR.Tn[0].t31 161.106
R23437 XThR.Tn[0].n57 XThR.Tn[0].t53 161.106
R23438 XThR.Tn[0].n52 XThR.Tn[0].t34 161.106
R23439 XThR.Tn[0].n47 XThR.Tn[0].t14 161.106
R23440 XThR.Tn[0].n42 XThR.Tn[0].t63 161.106
R23441 XThR.Tn[0].n37 XThR.Tn[0].t68 161.106
R23442 XThR.Tn[0].n32 XThR.Tn[0].t52 161.106
R23443 XThR.Tn[0].n27 XThR.Tn[0].t15 161.106
R23444 XThR.Tn[0].n22 XThR.Tn[0].t51 161.106
R23445 XThR.Tn[0].n17 XThR.Tn[0].t33 161.106
R23446 XThR.Tn[0].n12 XThR.Tn[0].t58 161.106
R23447 XThR.Tn[0].n10 XThR.Tn[0].t40 161.106
R23448 XThR.Tn[0].n83 XThR.Tn[0].t20 159.978
R23449 XThR.Tn[0].n78 XThR.Tn[0].t30 159.978
R23450 XThR.Tn[0].n73 XThR.Tn[0].t73 159.978
R23451 XThR.Tn[0].n68 XThR.Tn[0].t57 159.978
R23452 XThR.Tn[0].n63 XThR.Tn[0].t19 159.978
R23453 XThR.Tn[0].n58 XThR.Tn[0].t49 159.978
R23454 XThR.Tn[0].n53 XThR.Tn[0].t29 159.978
R23455 XThR.Tn[0].n48 XThR.Tn[0].t71 159.978
R23456 XThR.Tn[0].n43 XThR.Tn[0].t55 159.978
R23457 XThR.Tn[0].n38 XThR.Tn[0].t64 159.978
R23458 XThR.Tn[0].n33 XThR.Tn[0].t46 159.978
R23459 XThR.Tn[0].n28 XThR.Tn[0].t72 159.978
R23460 XThR.Tn[0].n23 XThR.Tn[0].t44 159.978
R23461 XThR.Tn[0].n18 XThR.Tn[0].t26 159.978
R23462 XThR.Tn[0].n13 XThR.Tn[0].t50 159.978
R23463 XThR.Tn[0].n82 XThR.Tn[0].t18 145.038
R23464 XThR.Tn[0].n77 XThR.Tn[0].t42 145.038
R23465 XThR.Tn[0].n72 XThR.Tn[0].t22 145.038
R23466 XThR.Tn[0].n67 XThR.Tn[0].t69 145.038
R23467 XThR.Tn[0].n62 XThR.Tn[0].t37 145.038
R23468 XThR.Tn[0].n57 XThR.Tn[0].t17 145.038
R23469 XThR.Tn[0].n52 XThR.Tn[0].t25 145.038
R23470 XThR.Tn[0].n47 XThR.Tn[0].t70 145.038
R23471 XThR.Tn[0].n42 XThR.Tn[0].t66 145.038
R23472 XThR.Tn[0].n37 XThR.Tn[0].t35 145.038
R23473 XThR.Tn[0].n32 XThR.Tn[0].t60 145.038
R23474 XThR.Tn[0].n27 XThR.Tn[0].t21 145.038
R23475 XThR.Tn[0].n22 XThR.Tn[0].t59 145.038
R23476 XThR.Tn[0].n17 XThR.Tn[0].t41 145.038
R23477 XThR.Tn[0].n12 XThR.Tn[0].t67 145.038
R23478 XThR.Tn[0].n10 XThR.Tn[0].t48 145.038
R23479 XThR.Tn[0].n83 XThR.Tn[0].t39 143.911
R23480 XThR.Tn[0].n78 XThR.Tn[0].t62 143.911
R23481 XThR.Tn[0].n73 XThR.Tn[0].t45 143.911
R23482 XThR.Tn[0].n68 XThR.Tn[0].t27 143.911
R23483 XThR.Tn[0].n63 XThR.Tn[0].t56 143.911
R23484 XThR.Tn[0].n58 XThR.Tn[0].t38 143.911
R23485 XThR.Tn[0].n53 XThR.Tn[0].t47 143.911
R23486 XThR.Tn[0].n48 XThR.Tn[0].t28 143.911
R23487 XThR.Tn[0].n43 XThR.Tn[0].t23 143.911
R23488 XThR.Tn[0].n38 XThR.Tn[0].t54 143.911
R23489 XThR.Tn[0].n33 XThR.Tn[0].t13 143.911
R23490 XThR.Tn[0].n28 XThR.Tn[0].t43 143.911
R23491 XThR.Tn[0].n23 XThR.Tn[0].t12 143.911
R23492 XThR.Tn[0].n18 XThR.Tn[0].t61 143.911
R23493 XThR.Tn[0].n13 XThR.Tn[0].t24 143.911
R23494 XThR.Tn[0].n7 XThR.Tn[0].n5 135.249
R23495 XThR.Tn[0].n9 XThR.Tn[0].n3 98.982
R23496 XThR.Tn[0].n8 XThR.Tn[0].n4 98.982
R23497 XThR.Tn[0].n7 XThR.Tn[0].n6 98.982
R23498 XThR.Tn[0].n9 XThR.Tn[0].n8 36.2672
R23499 XThR.Tn[0].n8 XThR.Tn[0].n7 36.2672
R23500 XThR.Tn[0].n88 XThR.Tn[0].n9 32.6405
R23501 XThR.Tn[0].n1 XThR.Tn[0].t5 26.5955
R23502 XThR.Tn[0].n1 XThR.Tn[0].t4 26.5955
R23503 XThR.Tn[0].n0 XThR.Tn[0].t6 26.5955
R23504 XThR.Tn[0].n0 XThR.Tn[0].t7 26.5955
R23505 XThR.Tn[0].n3 XThR.Tn[0].t9 24.9236
R23506 XThR.Tn[0].n3 XThR.Tn[0].t10 24.9236
R23507 XThR.Tn[0].n4 XThR.Tn[0].t8 24.9236
R23508 XThR.Tn[0].n4 XThR.Tn[0].t11 24.9236
R23509 XThR.Tn[0].n5 XThR.Tn[0].t1 24.9236
R23510 XThR.Tn[0].n5 XThR.Tn[0].t2 24.9236
R23511 XThR.Tn[0].n6 XThR.Tn[0].t0 24.9236
R23512 XThR.Tn[0].n6 XThR.Tn[0].t3 24.9236
R23513 XThR.Tn[0] XThR.Tn[0].n2 23.3605
R23514 XThR.Tn[0] XThR.Tn[0].n88 6.7205
R23515 XThR.Tn[0].n88 XThR.Tn[0] 6.36522
R23516 XThR.Tn[0] XThR.Tn[0].n11 5.34038
R23517 XThR.Tn[0].n16 XThR.Tn[0].n15 4.5005
R23518 XThR.Tn[0].n21 XThR.Tn[0].n20 4.5005
R23519 XThR.Tn[0].n26 XThR.Tn[0].n25 4.5005
R23520 XThR.Tn[0].n31 XThR.Tn[0].n30 4.5005
R23521 XThR.Tn[0].n36 XThR.Tn[0].n35 4.5005
R23522 XThR.Tn[0].n41 XThR.Tn[0].n40 4.5005
R23523 XThR.Tn[0].n46 XThR.Tn[0].n45 4.5005
R23524 XThR.Tn[0].n51 XThR.Tn[0].n50 4.5005
R23525 XThR.Tn[0].n56 XThR.Tn[0].n55 4.5005
R23526 XThR.Tn[0].n61 XThR.Tn[0].n60 4.5005
R23527 XThR.Tn[0].n66 XThR.Tn[0].n65 4.5005
R23528 XThR.Tn[0].n71 XThR.Tn[0].n70 4.5005
R23529 XThR.Tn[0].n76 XThR.Tn[0].n75 4.5005
R23530 XThR.Tn[0].n81 XThR.Tn[0].n80 4.5005
R23531 XThR.Tn[0].n86 XThR.Tn[0].n85 4.5005
R23532 XThR.Tn[0].n87 XThR.Tn[0] 3.70586
R23533 XThR.Tn[0].n16 XThR.Tn[0] 2.52282
R23534 XThR.Tn[0].n21 XThR.Tn[0] 2.52282
R23535 XThR.Tn[0].n26 XThR.Tn[0] 2.52282
R23536 XThR.Tn[0].n31 XThR.Tn[0] 2.52282
R23537 XThR.Tn[0].n36 XThR.Tn[0] 2.52282
R23538 XThR.Tn[0].n41 XThR.Tn[0] 2.52282
R23539 XThR.Tn[0].n46 XThR.Tn[0] 2.52282
R23540 XThR.Tn[0].n51 XThR.Tn[0] 2.52282
R23541 XThR.Tn[0].n56 XThR.Tn[0] 2.52282
R23542 XThR.Tn[0].n61 XThR.Tn[0] 2.52282
R23543 XThR.Tn[0].n66 XThR.Tn[0] 2.52282
R23544 XThR.Tn[0].n71 XThR.Tn[0] 2.52282
R23545 XThR.Tn[0].n76 XThR.Tn[0] 2.52282
R23546 XThR.Tn[0].n81 XThR.Tn[0] 2.52282
R23547 XThR.Tn[0].n86 XThR.Tn[0] 2.52282
R23548 XThR.Tn[0].n84 XThR.Tn[0] 1.08677
R23549 XThR.Tn[0].n79 XThR.Tn[0] 1.08677
R23550 XThR.Tn[0].n74 XThR.Tn[0] 1.08677
R23551 XThR.Tn[0].n69 XThR.Tn[0] 1.08677
R23552 XThR.Tn[0].n64 XThR.Tn[0] 1.08677
R23553 XThR.Tn[0].n59 XThR.Tn[0] 1.08677
R23554 XThR.Tn[0].n54 XThR.Tn[0] 1.08677
R23555 XThR.Tn[0].n49 XThR.Tn[0] 1.08677
R23556 XThR.Tn[0].n44 XThR.Tn[0] 1.08677
R23557 XThR.Tn[0].n39 XThR.Tn[0] 1.08677
R23558 XThR.Tn[0].n34 XThR.Tn[0] 1.08677
R23559 XThR.Tn[0].n29 XThR.Tn[0] 1.08677
R23560 XThR.Tn[0].n24 XThR.Tn[0] 1.08677
R23561 XThR.Tn[0].n19 XThR.Tn[0] 1.08677
R23562 XThR.Tn[0].n14 XThR.Tn[0] 1.08677
R23563 XThR.Tn[0] XThR.Tn[0].n16 0.839786
R23564 XThR.Tn[0] XThR.Tn[0].n21 0.839786
R23565 XThR.Tn[0] XThR.Tn[0].n26 0.839786
R23566 XThR.Tn[0] XThR.Tn[0].n31 0.839786
R23567 XThR.Tn[0] XThR.Tn[0].n36 0.839786
R23568 XThR.Tn[0] XThR.Tn[0].n41 0.839786
R23569 XThR.Tn[0] XThR.Tn[0].n46 0.839786
R23570 XThR.Tn[0] XThR.Tn[0].n51 0.839786
R23571 XThR.Tn[0] XThR.Tn[0].n56 0.839786
R23572 XThR.Tn[0] XThR.Tn[0].n61 0.839786
R23573 XThR.Tn[0] XThR.Tn[0].n66 0.839786
R23574 XThR.Tn[0] XThR.Tn[0].n71 0.839786
R23575 XThR.Tn[0] XThR.Tn[0].n76 0.839786
R23576 XThR.Tn[0] XThR.Tn[0].n81 0.839786
R23577 XThR.Tn[0] XThR.Tn[0].n86 0.839786
R23578 XThR.Tn[0].n11 XThR.Tn[0] 0.499542
R23579 XThR.Tn[0].n85 XThR.Tn[0] 0.063
R23580 XThR.Tn[0].n80 XThR.Tn[0] 0.063
R23581 XThR.Tn[0].n75 XThR.Tn[0] 0.063
R23582 XThR.Tn[0].n70 XThR.Tn[0] 0.063
R23583 XThR.Tn[0].n65 XThR.Tn[0] 0.063
R23584 XThR.Tn[0].n60 XThR.Tn[0] 0.063
R23585 XThR.Tn[0].n55 XThR.Tn[0] 0.063
R23586 XThR.Tn[0].n50 XThR.Tn[0] 0.063
R23587 XThR.Tn[0].n45 XThR.Tn[0] 0.063
R23588 XThR.Tn[0].n40 XThR.Tn[0] 0.063
R23589 XThR.Tn[0].n35 XThR.Tn[0] 0.063
R23590 XThR.Tn[0].n30 XThR.Tn[0] 0.063
R23591 XThR.Tn[0].n25 XThR.Tn[0] 0.063
R23592 XThR.Tn[0].n20 XThR.Tn[0] 0.063
R23593 XThR.Tn[0].n15 XThR.Tn[0] 0.063
R23594 XThR.Tn[0].n87 XThR.Tn[0] 0.0540714
R23595 XThR.Tn[0] XThR.Tn[0].n87 0.038
R23596 XThR.Tn[0].n11 XThR.Tn[0] 0.0143889
R23597 XThR.Tn[0].n85 XThR.Tn[0].n84 0.00771154
R23598 XThR.Tn[0].n80 XThR.Tn[0].n79 0.00771154
R23599 XThR.Tn[0].n75 XThR.Tn[0].n74 0.00771154
R23600 XThR.Tn[0].n70 XThR.Tn[0].n69 0.00771154
R23601 XThR.Tn[0].n65 XThR.Tn[0].n64 0.00771154
R23602 XThR.Tn[0].n60 XThR.Tn[0].n59 0.00771154
R23603 XThR.Tn[0].n55 XThR.Tn[0].n54 0.00771154
R23604 XThR.Tn[0].n50 XThR.Tn[0].n49 0.00771154
R23605 XThR.Tn[0].n45 XThR.Tn[0].n44 0.00771154
R23606 XThR.Tn[0].n40 XThR.Tn[0].n39 0.00771154
R23607 XThR.Tn[0].n35 XThR.Tn[0].n34 0.00771154
R23608 XThR.Tn[0].n30 XThR.Tn[0].n29 0.00771154
R23609 XThR.Tn[0].n25 XThR.Tn[0].n24 0.00771154
R23610 XThR.Tn[0].n20 XThR.Tn[0].n19 0.00771154
R23611 XThR.Tn[0].n15 XThR.Tn[0].n14 0.00771154
R23612 XThR.Tn[8].n5 XThR.Tn[8].n4 256.103
R23613 XThR.Tn[8].n2 XThR.Tn[8].n0 243.68
R23614 XThR.Tn[8].n88 XThR.Tn[8].n87 241.847
R23615 XThR.Tn[8].n2 XThR.Tn[8].n1 205.28
R23616 XThR.Tn[8].n5 XThR.Tn[8].n3 202.095
R23617 XThR.Tn[8].n88 XThR.Tn[8].n86 185
R23618 XThR.Tn[8] XThR.Tn[8].n79 161.363
R23619 XThR.Tn[8] XThR.Tn[8].n74 161.363
R23620 XThR.Tn[8] XThR.Tn[8].n69 161.363
R23621 XThR.Tn[8] XThR.Tn[8].n64 161.363
R23622 XThR.Tn[8] XThR.Tn[8].n59 161.363
R23623 XThR.Tn[8] XThR.Tn[8].n54 161.363
R23624 XThR.Tn[8] XThR.Tn[8].n49 161.363
R23625 XThR.Tn[8] XThR.Tn[8].n44 161.363
R23626 XThR.Tn[8] XThR.Tn[8].n39 161.363
R23627 XThR.Tn[8] XThR.Tn[8].n34 161.363
R23628 XThR.Tn[8] XThR.Tn[8].n29 161.363
R23629 XThR.Tn[8] XThR.Tn[8].n24 161.363
R23630 XThR.Tn[8] XThR.Tn[8].n19 161.363
R23631 XThR.Tn[8] XThR.Tn[8].n14 161.363
R23632 XThR.Tn[8] XThR.Tn[8].n9 161.363
R23633 XThR.Tn[8] XThR.Tn[8].n7 161.363
R23634 XThR.Tn[8].n81 XThR.Tn[8].n80 161.3
R23635 XThR.Tn[8].n76 XThR.Tn[8].n75 161.3
R23636 XThR.Tn[8].n71 XThR.Tn[8].n70 161.3
R23637 XThR.Tn[8].n66 XThR.Tn[8].n65 161.3
R23638 XThR.Tn[8].n61 XThR.Tn[8].n60 161.3
R23639 XThR.Tn[8].n56 XThR.Tn[8].n55 161.3
R23640 XThR.Tn[8].n51 XThR.Tn[8].n50 161.3
R23641 XThR.Tn[8].n46 XThR.Tn[8].n45 161.3
R23642 XThR.Tn[8].n41 XThR.Tn[8].n40 161.3
R23643 XThR.Tn[8].n36 XThR.Tn[8].n35 161.3
R23644 XThR.Tn[8].n31 XThR.Tn[8].n30 161.3
R23645 XThR.Tn[8].n26 XThR.Tn[8].n25 161.3
R23646 XThR.Tn[8].n21 XThR.Tn[8].n20 161.3
R23647 XThR.Tn[8].n16 XThR.Tn[8].n15 161.3
R23648 XThR.Tn[8].n11 XThR.Tn[8].n10 161.3
R23649 XThR.Tn[8].n79 XThR.Tn[8].t23 161.106
R23650 XThR.Tn[8].n74 XThR.Tn[8].t29 161.106
R23651 XThR.Tn[8].n69 XThR.Tn[8].t71 161.106
R23652 XThR.Tn[8].n64 XThR.Tn[8].t57 161.106
R23653 XThR.Tn[8].n59 XThR.Tn[8].t21 161.106
R23654 XThR.Tn[8].n54 XThR.Tn[8].t46 161.106
R23655 XThR.Tn[8].n49 XThR.Tn[8].t27 161.106
R23656 XThR.Tn[8].n44 XThR.Tn[8].t69 161.106
R23657 XThR.Tn[8].n39 XThR.Tn[8].t56 161.106
R23658 XThR.Tn[8].n34 XThR.Tn[8].t61 161.106
R23659 XThR.Tn[8].n29 XThR.Tn[8].t44 161.106
R23660 XThR.Tn[8].n24 XThR.Tn[8].t70 161.106
R23661 XThR.Tn[8].n19 XThR.Tn[8].t43 161.106
R23662 XThR.Tn[8].n14 XThR.Tn[8].t26 161.106
R23663 XThR.Tn[8].n9 XThR.Tn[8].t49 161.106
R23664 XThR.Tn[8].n7 XThR.Tn[8].t33 161.106
R23665 XThR.Tn[8].n80 XThR.Tn[8].t19 159.978
R23666 XThR.Tn[8].n75 XThR.Tn[8].t25 159.978
R23667 XThR.Tn[8].n70 XThR.Tn[8].t67 159.978
R23668 XThR.Tn[8].n65 XThR.Tn[8].t54 159.978
R23669 XThR.Tn[8].n60 XThR.Tn[8].t16 159.978
R23670 XThR.Tn[8].n55 XThR.Tn[8].t42 159.978
R23671 XThR.Tn[8].n50 XThR.Tn[8].t24 159.978
R23672 XThR.Tn[8].n45 XThR.Tn[8].t64 159.978
R23673 XThR.Tn[8].n40 XThR.Tn[8].t51 159.978
R23674 XThR.Tn[8].n35 XThR.Tn[8].t58 159.978
R23675 XThR.Tn[8].n30 XThR.Tn[8].t41 159.978
R23676 XThR.Tn[8].n25 XThR.Tn[8].t66 159.978
R23677 XThR.Tn[8].n20 XThR.Tn[8].t40 159.978
R23678 XThR.Tn[8].n15 XThR.Tn[8].t22 159.978
R23679 XThR.Tn[8].n10 XThR.Tn[8].t45 159.978
R23680 XThR.Tn[8].n79 XThR.Tn[8].t73 145.038
R23681 XThR.Tn[8].n74 XThR.Tn[8].t35 145.038
R23682 XThR.Tn[8].n69 XThR.Tn[8].t15 145.038
R23683 XThR.Tn[8].n64 XThR.Tn[8].t62 145.038
R23684 XThR.Tn[8].n59 XThR.Tn[8].t30 145.038
R23685 XThR.Tn[8].n54 XThR.Tn[8].t72 145.038
R23686 XThR.Tn[8].n49 XThR.Tn[8].t17 145.038
R23687 XThR.Tn[8].n44 XThR.Tn[8].t63 145.038
R23688 XThR.Tn[8].n39 XThR.Tn[8].t60 145.038
R23689 XThR.Tn[8].n34 XThR.Tn[8].t28 145.038
R23690 XThR.Tn[8].n29 XThR.Tn[8].t52 145.038
R23691 XThR.Tn[8].n24 XThR.Tn[8].t12 145.038
R23692 XThR.Tn[8].n19 XThR.Tn[8].t50 145.038
R23693 XThR.Tn[8].n14 XThR.Tn[8].t34 145.038
R23694 XThR.Tn[8].n9 XThR.Tn[8].t59 145.038
R23695 XThR.Tn[8].n7 XThR.Tn[8].t39 145.038
R23696 XThR.Tn[8].n80 XThR.Tn[8].t32 143.911
R23697 XThR.Tn[8].n75 XThR.Tn[8].t55 143.911
R23698 XThR.Tn[8].n70 XThR.Tn[8].t37 143.911
R23699 XThR.Tn[8].n65 XThR.Tn[8].t18 143.911
R23700 XThR.Tn[8].n60 XThR.Tn[8].t48 143.911
R23701 XThR.Tn[8].n55 XThR.Tn[8].t31 143.911
R23702 XThR.Tn[8].n50 XThR.Tn[8].t38 143.911
R23703 XThR.Tn[8].n45 XThR.Tn[8].t20 143.911
R23704 XThR.Tn[8].n40 XThR.Tn[8].t14 143.911
R23705 XThR.Tn[8].n35 XThR.Tn[8].t47 143.911
R23706 XThR.Tn[8].n30 XThR.Tn[8].t68 143.911
R23707 XThR.Tn[8].n25 XThR.Tn[8].t36 143.911
R23708 XThR.Tn[8].n20 XThR.Tn[8].t65 143.911
R23709 XThR.Tn[8].n15 XThR.Tn[8].t53 143.911
R23710 XThR.Tn[8].n10 XThR.Tn[8].t13 143.911
R23711 XThR.Tn[8] XThR.Tn[8].n2 35.7652
R23712 XThR.Tn[8].n3 XThR.Tn[8].t6 26.5955
R23713 XThR.Tn[8].n3 XThR.Tn[8].t4 26.5955
R23714 XThR.Tn[8].n4 XThR.Tn[8].t7 26.5955
R23715 XThR.Tn[8].n4 XThR.Tn[8].t5 26.5955
R23716 XThR.Tn[8].n0 XThR.Tn[8].t10 26.5955
R23717 XThR.Tn[8].n0 XThR.Tn[8].t8 26.5955
R23718 XThR.Tn[8].n1 XThR.Tn[8].t11 26.5955
R23719 XThR.Tn[8].n1 XThR.Tn[8].t9 26.5955
R23720 XThR.Tn[8].n86 XThR.Tn[8].t0 24.9236
R23721 XThR.Tn[8].n86 XThR.Tn[8].t2 24.9236
R23722 XThR.Tn[8].n87 XThR.Tn[8].t1 24.9236
R23723 XThR.Tn[8].n87 XThR.Tn[8].t3 24.9236
R23724 XThR.Tn[8] XThR.Tn[8].n88 18.8943
R23725 XThR.Tn[8].n6 XThR.Tn[8].n5 13.5534
R23726 XThR.Tn[8].n85 XThR.Tn[8] 7.82692
R23727 XThR.Tn[8] XThR.Tn[8].n85 6.34069
R23728 XThR.Tn[8] XThR.Tn[8].n8 5.34038
R23729 XThR.Tn[8].n13 XThR.Tn[8].n12 4.5005
R23730 XThR.Tn[8].n18 XThR.Tn[8].n17 4.5005
R23731 XThR.Tn[8].n23 XThR.Tn[8].n22 4.5005
R23732 XThR.Tn[8].n28 XThR.Tn[8].n27 4.5005
R23733 XThR.Tn[8].n33 XThR.Tn[8].n32 4.5005
R23734 XThR.Tn[8].n38 XThR.Tn[8].n37 4.5005
R23735 XThR.Tn[8].n43 XThR.Tn[8].n42 4.5005
R23736 XThR.Tn[8].n48 XThR.Tn[8].n47 4.5005
R23737 XThR.Tn[8].n53 XThR.Tn[8].n52 4.5005
R23738 XThR.Tn[8].n58 XThR.Tn[8].n57 4.5005
R23739 XThR.Tn[8].n63 XThR.Tn[8].n62 4.5005
R23740 XThR.Tn[8].n68 XThR.Tn[8].n67 4.5005
R23741 XThR.Tn[8].n73 XThR.Tn[8].n72 4.5005
R23742 XThR.Tn[8].n78 XThR.Tn[8].n77 4.5005
R23743 XThR.Tn[8].n83 XThR.Tn[8].n82 4.5005
R23744 XThR.Tn[8].n84 XThR.Tn[8] 3.70586
R23745 XThR.Tn[8].n13 XThR.Tn[8] 2.52282
R23746 XThR.Tn[8].n18 XThR.Tn[8] 2.52282
R23747 XThR.Tn[8].n23 XThR.Tn[8] 2.52282
R23748 XThR.Tn[8].n28 XThR.Tn[8] 2.52282
R23749 XThR.Tn[8].n33 XThR.Tn[8] 2.52282
R23750 XThR.Tn[8].n38 XThR.Tn[8] 2.52282
R23751 XThR.Tn[8].n43 XThR.Tn[8] 2.52282
R23752 XThR.Tn[8].n48 XThR.Tn[8] 2.52282
R23753 XThR.Tn[8].n53 XThR.Tn[8] 2.52282
R23754 XThR.Tn[8].n58 XThR.Tn[8] 2.52282
R23755 XThR.Tn[8].n63 XThR.Tn[8] 2.52282
R23756 XThR.Tn[8].n68 XThR.Tn[8] 2.52282
R23757 XThR.Tn[8].n73 XThR.Tn[8] 2.52282
R23758 XThR.Tn[8].n78 XThR.Tn[8] 2.52282
R23759 XThR.Tn[8].n83 XThR.Tn[8] 2.52282
R23760 XThR.Tn[8].n85 XThR.Tn[8] 1.79489
R23761 XThR.Tn[8].n6 XThR.Tn[8] 1.50638
R23762 XThR.Tn[8] XThR.Tn[8].n6 1.19676
R23763 XThR.Tn[8].n81 XThR.Tn[8] 1.08677
R23764 XThR.Tn[8].n76 XThR.Tn[8] 1.08677
R23765 XThR.Tn[8].n71 XThR.Tn[8] 1.08677
R23766 XThR.Tn[8].n66 XThR.Tn[8] 1.08677
R23767 XThR.Tn[8].n61 XThR.Tn[8] 1.08677
R23768 XThR.Tn[8].n56 XThR.Tn[8] 1.08677
R23769 XThR.Tn[8].n51 XThR.Tn[8] 1.08677
R23770 XThR.Tn[8].n46 XThR.Tn[8] 1.08677
R23771 XThR.Tn[8].n41 XThR.Tn[8] 1.08677
R23772 XThR.Tn[8].n36 XThR.Tn[8] 1.08677
R23773 XThR.Tn[8].n31 XThR.Tn[8] 1.08677
R23774 XThR.Tn[8].n26 XThR.Tn[8] 1.08677
R23775 XThR.Tn[8].n21 XThR.Tn[8] 1.08677
R23776 XThR.Tn[8].n16 XThR.Tn[8] 1.08677
R23777 XThR.Tn[8].n11 XThR.Tn[8] 1.08677
R23778 XThR.Tn[8] XThR.Tn[8].n13 0.839786
R23779 XThR.Tn[8] XThR.Tn[8].n18 0.839786
R23780 XThR.Tn[8] XThR.Tn[8].n23 0.839786
R23781 XThR.Tn[8] XThR.Tn[8].n28 0.839786
R23782 XThR.Tn[8] XThR.Tn[8].n33 0.839786
R23783 XThR.Tn[8] XThR.Tn[8].n38 0.839786
R23784 XThR.Tn[8] XThR.Tn[8].n43 0.839786
R23785 XThR.Tn[8] XThR.Tn[8].n48 0.839786
R23786 XThR.Tn[8] XThR.Tn[8].n53 0.839786
R23787 XThR.Tn[8] XThR.Tn[8].n58 0.839786
R23788 XThR.Tn[8] XThR.Tn[8].n63 0.839786
R23789 XThR.Tn[8] XThR.Tn[8].n68 0.839786
R23790 XThR.Tn[8] XThR.Tn[8].n73 0.839786
R23791 XThR.Tn[8] XThR.Tn[8].n78 0.839786
R23792 XThR.Tn[8] XThR.Tn[8].n83 0.839786
R23793 XThR.Tn[8].n8 XThR.Tn[8] 0.499542
R23794 XThR.Tn[8].n82 XThR.Tn[8] 0.063
R23795 XThR.Tn[8].n77 XThR.Tn[8] 0.063
R23796 XThR.Tn[8].n72 XThR.Tn[8] 0.063
R23797 XThR.Tn[8].n67 XThR.Tn[8] 0.063
R23798 XThR.Tn[8].n62 XThR.Tn[8] 0.063
R23799 XThR.Tn[8].n57 XThR.Tn[8] 0.063
R23800 XThR.Tn[8].n52 XThR.Tn[8] 0.063
R23801 XThR.Tn[8].n47 XThR.Tn[8] 0.063
R23802 XThR.Tn[8].n42 XThR.Tn[8] 0.063
R23803 XThR.Tn[8].n37 XThR.Tn[8] 0.063
R23804 XThR.Tn[8].n32 XThR.Tn[8] 0.063
R23805 XThR.Tn[8].n27 XThR.Tn[8] 0.063
R23806 XThR.Tn[8].n22 XThR.Tn[8] 0.063
R23807 XThR.Tn[8].n17 XThR.Tn[8] 0.063
R23808 XThR.Tn[8].n12 XThR.Tn[8] 0.063
R23809 XThR.Tn[8].n84 XThR.Tn[8] 0.0540714
R23810 XThR.Tn[8] XThR.Tn[8].n84 0.038
R23811 XThR.Tn[8].n8 XThR.Tn[8] 0.0143889
R23812 XThR.Tn[8].n82 XThR.Tn[8].n81 0.00771154
R23813 XThR.Tn[8].n77 XThR.Tn[8].n76 0.00771154
R23814 XThR.Tn[8].n72 XThR.Tn[8].n71 0.00771154
R23815 XThR.Tn[8].n67 XThR.Tn[8].n66 0.00771154
R23816 XThR.Tn[8].n62 XThR.Tn[8].n61 0.00771154
R23817 XThR.Tn[8].n57 XThR.Tn[8].n56 0.00771154
R23818 XThR.Tn[8].n52 XThR.Tn[8].n51 0.00771154
R23819 XThR.Tn[8].n47 XThR.Tn[8].n46 0.00771154
R23820 XThR.Tn[8].n42 XThR.Tn[8].n41 0.00771154
R23821 XThR.Tn[8].n37 XThR.Tn[8].n36 0.00771154
R23822 XThR.Tn[8].n32 XThR.Tn[8].n31 0.00771154
R23823 XThR.Tn[8].n27 XThR.Tn[8].n26 0.00771154
R23824 XThR.Tn[8].n22 XThR.Tn[8].n21 0.00771154
R23825 XThR.Tn[8].n17 XThR.Tn[8].n16 0.00771154
R23826 XThR.Tn[8].n12 XThR.Tn[8].n11 0.00771154
R23827 XThC.XTB3.Y.n6 XThC.XTB3.Y.t3 212.081
R23828 XThC.XTB3.Y.n5 XThC.XTB3.Y.t15 212.081
R23829 XThC.XTB3.Y.n11 XThC.XTB3.Y.t14 212.081
R23830 XThC.XTB3.Y.n3 XThC.XTB3.Y.t10 212.081
R23831 XThC.XTB3.Y.n15 XThC.XTB3.Y.t11 212.081
R23832 XThC.XTB3.Y.n16 XThC.XTB3.Y.t12 212.081
R23833 XThC.XTB3.Y.n18 XThC.XTB3.Y.t4 212.081
R23834 XThC.XTB3.Y.n14 XThC.XTB3.Y.t16 212.081
R23835 XThC.XTB3.Y.n22 XThC.XTB3.Y.n2 201.288
R23836 XThC.XTB3.Y.n8 XThC.XTB3.Y.n7 173.761
R23837 XThC.XTB3.Y.n17 XThC.XTB3.Y 158.656
R23838 XThC.XTB3.Y.n10 XThC.XTB3.Y.n9 152
R23839 XThC.XTB3.Y.n8 XThC.XTB3.Y.n4 152
R23840 XThC.XTB3.Y.n13 XThC.XTB3.Y.n12 152
R23841 XThC.XTB3.Y.n20 XThC.XTB3.Y.n19 152
R23842 XThC.XTB3.Y.n6 XThC.XTB3.Y.t9 139.78
R23843 XThC.XTB3.Y.n5 XThC.XTB3.Y.t6 139.78
R23844 XThC.XTB3.Y.n11 XThC.XTB3.Y.t5 139.78
R23845 XThC.XTB3.Y.n3 XThC.XTB3.Y.t17 139.78
R23846 XThC.XTB3.Y.n15 XThC.XTB3.Y.t8 139.78
R23847 XThC.XTB3.Y.n16 XThC.XTB3.Y.t18 139.78
R23848 XThC.XTB3.Y.n18 XThC.XTB3.Y.t13 139.78
R23849 XThC.XTB3.Y.n14 XThC.XTB3.Y.t7 139.78
R23850 XThC.XTB3.Y.n0 XThC.XTB3.Y.t1 132.067
R23851 XThC.XTB3.Y.n21 XThC.XTB3.Y.n13 61.4096
R23852 XThC.XTB3.Y.n16 XThC.XTB3.Y.n15 61.346
R23853 XThC.XTB3.Y.n21 XThC.XTB3.Y 54.2785
R23854 XThC.XTB3.Y.n10 XThC.XTB3.Y.n4 49.6611
R23855 XThC.XTB3.Y.n12 XThC.XTB3.Y.n11 45.2793
R23856 XThC.XTB3.Y.n7 XThC.XTB3.Y.n5 42.3581
R23857 XThC.XTB3.Y.n19 XThC.XTB3.Y.n14 30.6732
R23858 XThC.XTB3.Y.n19 XThC.XTB3.Y.n18 30.6732
R23859 XThC.XTB3.Y.n18 XThC.XTB3.Y.n17 30.6732
R23860 XThC.XTB3.Y.n17 XThC.XTB3.Y.n16 30.6732
R23861 XThC.XTB3.Y.n2 XThC.XTB3.Y.t2 26.5955
R23862 XThC.XTB3.Y.n2 XThC.XTB3.Y.t0 26.5955
R23863 XThC.XTB3.Y XThC.XTB3.Y.n22 23.489
R23864 XThC.XTB3.Y.n9 XThC.XTB3.Y.n8 21.7605
R23865 XThC.XTB3.Y.n7 XThC.XTB3.Y.n6 18.9884
R23866 XThC.XTB3.Y.n12 XThC.XTB3.Y.n3 16.0672
R23867 XThC.XTB3.Y.n20 XThC.XTB3.Y 14.8485
R23868 XThC.XTB3.Y.n13 XThC.XTB3.Y 11.5205
R23869 XThC.XTB3.Y.n22 XThC.XTB3.Y.n21 10.8207
R23870 XThC.XTB3.Y.n9 XThC.XTB3.Y 10.2405
R23871 XThC.XTB3.Y XThC.XTB3.Y.n20 8.7045
R23872 XThC.XTB3.Y.n5 XThC.XTB3.Y.n4 7.30353
R23873 XThC.XTB3.Y.n11 XThC.XTB3.Y.n10 4.38232
R23874 XThC.XTB3.Y.n1 XThC.XTB3.Y.n0 4.15748
R23875 XThC.XTB3.Y XThC.XTB3.Y.n1 3.76521
R23876 XThC.XTB3.Y.n0 XThC.XTB3.Y 1.17559
R23877 XThC.XTB3.Y.n1 XThC.XTB3.Y 0.921363
R23878 data[4].n3 data[4].t0 231.835
R23879 data[4].n0 data[4].t3 230.155
R23880 data[4].n0 data[4].t1 157.856
R23881 data[4].n3 data[4].t2 157.07
R23882 data[4].n1 data[4].n0 152
R23883 data[4].n4 data[4].n3 152
R23884 data[4].n2 data[4].n1 25.6681
R23885 data[4].n4 data[4].n2 10.7642
R23886 data[4].n2 data[4] 2.763
R23887 data[4].n1 data[4] 2.10199
R23888 data[4] data[4].n4 2.01193
R23889 XThR.Tn[13].n8 XThR.Tn[13].n7 256.104
R23890 XThR.Tn[13].n5 XThR.Tn[13].n3 243.68
R23891 XThR.Tn[13].n2 XThR.Tn[13].n1 241.847
R23892 XThR.Tn[13].n5 XThR.Tn[13].n4 205.28
R23893 XThR.Tn[13].n8 XThR.Tn[13].n6 202.094
R23894 XThR.Tn[13].n2 XThR.Tn[13].n0 185
R23895 XThR.Tn[13] XThR.Tn[13].n82 161.363
R23896 XThR.Tn[13] XThR.Tn[13].n77 161.363
R23897 XThR.Tn[13] XThR.Tn[13].n72 161.363
R23898 XThR.Tn[13] XThR.Tn[13].n67 161.363
R23899 XThR.Tn[13] XThR.Tn[13].n62 161.363
R23900 XThR.Tn[13] XThR.Tn[13].n57 161.363
R23901 XThR.Tn[13] XThR.Tn[13].n52 161.363
R23902 XThR.Tn[13] XThR.Tn[13].n47 161.363
R23903 XThR.Tn[13] XThR.Tn[13].n42 161.363
R23904 XThR.Tn[13] XThR.Tn[13].n37 161.363
R23905 XThR.Tn[13] XThR.Tn[13].n32 161.363
R23906 XThR.Tn[13] XThR.Tn[13].n27 161.363
R23907 XThR.Tn[13] XThR.Tn[13].n22 161.363
R23908 XThR.Tn[13] XThR.Tn[13].n17 161.363
R23909 XThR.Tn[13] XThR.Tn[13].n12 161.363
R23910 XThR.Tn[13] XThR.Tn[13].n10 161.363
R23911 XThR.Tn[13].n84 XThR.Tn[13].n83 161.3
R23912 XThR.Tn[13].n79 XThR.Tn[13].n78 161.3
R23913 XThR.Tn[13].n74 XThR.Tn[13].n73 161.3
R23914 XThR.Tn[13].n69 XThR.Tn[13].n68 161.3
R23915 XThR.Tn[13].n64 XThR.Tn[13].n63 161.3
R23916 XThR.Tn[13].n59 XThR.Tn[13].n58 161.3
R23917 XThR.Tn[13].n54 XThR.Tn[13].n53 161.3
R23918 XThR.Tn[13].n49 XThR.Tn[13].n48 161.3
R23919 XThR.Tn[13].n44 XThR.Tn[13].n43 161.3
R23920 XThR.Tn[13].n39 XThR.Tn[13].n38 161.3
R23921 XThR.Tn[13].n34 XThR.Tn[13].n33 161.3
R23922 XThR.Tn[13].n29 XThR.Tn[13].n28 161.3
R23923 XThR.Tn[13].n24 XThR.Tn[13].n23 161.3
R23924 XThR.Tn[13].n19 XThR.Tn[13].n18 161.3
R23925 XThR.Tn[13].n14 XThR.Tn[13].n13 161.3
R23926 XThR.Tn[13].n82 XThR.Tn[13].t56 161.106
R23927 XThR.Tn[13].n77 XThR.Tn[13].t62 161.106
R23928 XThR.Tn[13].n72 XThR.Tn[13].t40 161.106
R23929 XThR.Tn[13].n67 XThR.Tn[13].t27 161.106
R23930 XThR.Tn[13].n62 XThR.Tn[13].t55 161.106
R23931 XThR.Tn[13].n57 XThR.Tn[13].t17 161.106
R23932 XThR.Tn[13].n52 XThR.Tn[13].t59 161.106
R23933 XThR.Tn[13].n47 XThR.Tn[13].t38 161.106
R23934 XThR.Tn[13].n42 XThR.Tn[13].t25 161.106
R23935 XThR.Tn[13].n37 XThR.Tn[13].t30 161.106
R23936 XThR.Tn[13].n32 XThR.Tn[13].t16 161.106
R23937 XThR.Tn[13].n27 XThR.Tn[13].t39 161.106
R23938 XThR.Tn[13].n22 XThR.Tn[13].t14 161.106
R23939 XThR.Tn[13].n17 XThR.Tn[13].t57 161.106
R23940 XThR.Tn[13].n12 XThR.Tn[13].t21 161.106
R23941 XThR.Tn[13].n10 XThR.Tn[13].t64 161.106
R23942 XThR.Tn[13].n83 XThR.Tn[13].t47 159.978
R23943 XThR.Tn[13].n78 XThR.Tn[13].t54 159.978
R23944 XThR.Tn[13].n73 XThR.Tn[13].t36 159.978
R23945 XThR.Tn[13].n68 XThR.Tn[13].t20 159.978
R23946 XThR.Tn[13].n63 XThR.Tn[13].t45 159.978
R23947 XThR.Tn[13].n58 XThR.Tn[13].t73 159.978
R23948 XThR.Tn[13].n53 XThR.Tn[13].t53 159.978
R23949 XThR.Tn[13].n48 XThR.Tn[13].t33 159.978
R23950 XThR.Tn[13].n43 XThR.Tn[13].t18 159.978
R23951 XThR.Tn[13].n38 XThR.Tn[13].t26 159.978
R23952 XThR.Tn[13].n33 XThR.Tn[13].t71 159.978
R23953 XThR.Tn[13].n28 XThR.Tn[13].t35 159.978
R23954 XThR.Tn[13].n23 XThR.Tn[13].t70 159.978
R23955 XThR.Tn[13].n18 XThR.Tn[13].t52 159.978
R23956 XThR.Tn[13].n13 XThR.Tn[13].t12 159.978
R23957 XThR.Tn[13].n82 XThR.Tn[13].t42 145.038
R23958 XThR.Tn[13].n77 XThR.Tn[13].t69 145.038
R23959 XThR.Tn[13].n72 XThR.Tn[13].t50 145.038
R23960 XThR.Tn[13].n67 XThR.Tn[13].t31 145.038
R23961 XThR.Tn[13].n62 XThR.Tn[13].t63 145.038
R23962 XThR.Tn[13].n57 XThR.Tn[13].t41 145.038
R23963 XThR.Tn[13].n52 XThR.Tn[13].t51 145.038
R23964 XThR.Tn[13].n47 XThR.Tn[13].t32 145.038
R23965 XThR.Tn[13].n42 XThR.Tn[13].t29 145.038
R23966 XThR.Tn[13].n37 XThR.Tn[13].t60 145.038
R23967 XThR.Tn[13].n32 XThR.Tn[13].t24 145.038
R23968 XThR.Tn[13].n27 XThR.Tn[13].t49 145.038
R23969 XThR.Tn[13].n22 XThR.Tn[13].t22 145.038
R23970 XThR.Tn[13].n17 XThR.Tn[13].t65 145.038
R23971 XThR.Tn[13].n12 XThR.Tn[13].t28 145.038
R23972 XThR.Tn[13].n10 XThR.Tn[13].t72 145.038
R23973 XThR.Tn[13].n83 XThR.Tn[13].t61 143.911
R23974 XThR.Tn[13].n78 XThR.Tn[13].t23 143.911
R23975 XThR.Tn[13].n73 XThR.Tn[13].t67 143.911
R23976 XThR.Tn[13].n68 XThR.Tn[13].t46 143.911
R23977 XThR.Tn[13].n63 XThR.Tn[13].t15 143.911
R23978 XThR.Tn[13].n58 XThR.Tn[13].t58 143.911
R23979 XThR.Tn[13].n53 XThR.Tn[13].t68 143.911
R23980 XThR.Tn[13].n48 XThR.Tn[13].t48 143.911
R23981 XThR.Tn[13].n43 XThR.Tn[13].t43 143.911
R23982 XThR.Tn[13].n38 XThR.Tn[13].t13 143.911
R23983 XThR.Tn[13].n33 XThR.Tn[13].t37 143.911
R23984 XThR.Tn[13].n28 XThR.Tn[13].t66 143.911
R23985 XThR.Tn[13].n23 XThR.Tn[13].t34 143.911
R23986 XThR.Tn[13].n18 XThR.Tn[13].t19 143.911
R23987 XThR.Tn[13].n13 XThR.Tn[13].t44 143.911
R23988 XThR.Tn[13] XThR.Tn[13].n5 35.7652
R23989 XThR.Tn[13].n6 XThR.Tn[13].t6 26.5955
R23990 XThR.Tn[13].n6 XThR.Tn[13].t4 26.5955
R23991 XThR.Tn[13].n7 XThR.Tn[13].t7 26.5955
R23992 XThR.Tn[13].n7 XThR.Tn[13].t5 26.5955
R23993 XThR.Tn[13].n3 XThR.Tn[13].t9 26.5955
R23994 XThR.Tn[13].n3 XThR.Tn[13].t11 26.5955
R23995 XThR.Tn[13].n4 XThR.Tn[13].t10 26.5955
R23996 XThR.Tn[13].n4 XThR.Tn[13].t8 26.5955
R23997 XThR.Tn[13].n0 XThR.Tn[13].t2 24.9236
R23998 XThR.Tn[13].n0 XThR.Tn[13].t0 24.9236
R23999 XThR.Tn[13].n1 XThR.Tn[13].t3 24.9236
R24000 XThR.Tn[13].n1 XThR.Tn[13].t1 24.9236
R24001 XThR.Tn[13] XThR.Tn[13].n2 22.9615
R24002 XThR.Tn[13].n9 XThR.Tn[13].n8 13.5534
R24003 XThR.Tn[13].n88 XThR.Tn[13] 8.8494
R24004 XThR.Tn[13] XThR.Tn[13].n11 5.34038
R24005 XThR.Tn[13].n16 XThR.Tn[13].n15 4.5005
R24006 XThR.Tn[13].n21 XThR.Tn[13].n20 4.5005
R24007 XThR.Tn[13].n26 XThR.Tn[13].n25 4.5005
R24008 XThR.Tn[13].n31 XThR.Tn[13].n30 4.5005
R24009 XThR.Tn[13].n36 XThR.Tn[13].n35 4.5005
R24010 XThR.Tn[13].n41 XThR.Tn[13].n40 4.5005
R24011 XThR.Tn[13].n46 XThR.Tn[13].n45 4.5005
R24012 XThR.Tn[13].n51 XThR.Tn[13].n50 4.5005
R24013 XThR.Tn[13].n56 XThR.Tn[13].n55 4.5005
R24014 XThR.Tn[13].n61 XThR.Tn[13].n60 4.5005
R24015 XThR.Tn[13].n66 XThR.Tn[13].n65 4.5005
R24016 XThR.Tn[13].n71 XThR.Tn[13].n70 4.5005
R24017 XThR.Tn[13].n76 XThR.Tn[13].n75 4.5005
R24018 XThR.Tn[13].n81 XThR.Tn[13].n80 4.5005
R24019 XThR.Tn[13].n86 XThR.Tn[13].n85 4.5005
R24020 XThR.Tn[13].n87 XThR.Tn[13] 3.70586
R24021 XThR.Tn[13].n88 XThR.Tn[13].n9 2.99115
R24022 XThR.Tn[13].n9 XThR.Tn[13] 2.87153
R24023 XThR.Tn[13].n16 XThR.Tn[13] 2.52282
R24024 XThR.Tn[13].n21 XThR.Tn[13] 2.52282
R24025 XThR.Tn[13].n26 XThR.Tn[13] 2.52282
R24026 XThR.Tn[13].n31 XThR.Tn[13] 2.52282
R24027 XThR.Tn[13].n36 XThR.Tn[13] 2.52282
R24028 XThR.Tn[13].n41 XThR.Tn[13] 2.52282
R24029 XThR.Tn[13].n46 XThR.Tn[13] 2.52282
R24030 XThR.Tn[13].n51 XThR.Tn[13] 2.52282
R24031 XThR.Tn[13].n56 XThR.Tn[13] 2.52282
R24032 XThR.Tn[13].n61 XThR.Tn[13] 2.52282
R24033 XThR.Tn[13].n66 XThR.Tn[13] 2.52282
R24034 XThR.Tn[13].n71 XThR.Tn[13] 2.52282
R24035 XThR.Tn[13].n76 XThR.Tn[13] 2.52282
R24036 XThR.Tn[13].n81 XThR.Tn[13] 2.52282
R24037 XThR.Tn[13].n86 XThR.Tn[13] 2.52282
R24038 XThR.Tn[13] XThR.Tn[13].n88 2.2734
R24039 XThR.Tn[13].n9 XThR.Tn[13] 1.50638
R24040 XThR.Tn[13].n84 XThR.Tn[13] 1.08677
R24041 XThR.Tn[13].n79 XThR.Tn[13] 1.08677
R24042 XThR.Tn[13].n74 XThR.Tn[13] 1.08677
R24043 XThR.Tn[13].n69 XThR.Tn[13] 1.08677
R24044 XThR.Tn[13].n64 XThR.Tn[13] 1.08677
R24045 XThR.Tn[13].n59 XThR.Tn[13] 1.08677
R24046 XThR.Tn[13].n54 XThR.Tn[13] 1.08677
R24047 XThR.Tn[13].n49 XThR.Tn[13] 1.08677
R24048 XThR.Tn[13].n44 XThR.Tn[13] 1.08677
R24049 XThR.Tn[13].n39 XThR.Tn[13] 1.08677
R24050 XThR.Tn[13].n34 XThR.Tn[13] 1.08677
R24051 XThR.Tn[13].n29 XThR.Tn[13] 1.08677
R24052 XThR.Tn[13].n24 XThR.Tn[13] 1.08677
R24053 XThR.Tn[13].n19 XThR.Tn[13] 1.08677
R24054 XThR.Tn[13].n14 XThR.Tn[13] 1.08677
R24055 XThR.Tn[13] XThR.Tn[13].n16 0.839786
R24056 XThR.Tn[13] XThR.Tn[13].n21 0.839786
R24057 XThR.Tn[13] XThR.Tn[13].n26 0.839786
R24058 XThR.Tn[13] XThR.Tn[13].n31 0.839786
R24059 XThR.Tn[13] XThR.Tn[13].n36 0.839786
R24060 XThR.Tn[13] XThR.Tn[13].n41 0.839786
R24061 XThR.Tn[13] XThR.Tn[13].n46 0.839786
R24062 XThR.Tn[13] XThR.Tn[13].n51 0.839786
R24063 XThR.Tn[13] XThR.Tn[13].n56 0.839786
R24064 XThR.Tn[13] XThR.Tn[13].n61 0.839786
R24065 XThR.Tn[13] XThR.Tn[13].n66 0.839786
R24066 XThR.Tn[13] XThR.Tn[13].n71 0.839786
R24067 XThR.Tn[13] XThR.Tn[13].n76 0.839786
R24068 XThR.Tn[13] XThR.Tn[13].n81 0.839786
R24069 XThR.Tn[13] XThR.Tn[13].n86 0.839786
R24070 XThR.Tn[13].n11 XThR.Tn[13] 0.499542
R24071 XThR.Tn[13].n85 XThR.Tn[13] 0.063
R24072 XThR.Tn[13].n80 XThR.Tn[13] 0.063
R24073 XThR.Tn[13].n75 XThR.Tn[13] 0.063
R24074 XThR.Tn[13].n70 XThR.Tn[13] 0.063
R24075 XThR.Tn[13].n65 XThR.Tn[13] 0.063
R24076 XThR.Tn[13].n60 XThR.Tn[13] 0.063
R24077 XThR.Tn[13].n55 XThR.Tn[13] 0.063
R24078 XThR.Tn[13].n50 XThR.Tn[13] 0.063
R24079 XThR.Tn[13].n45 XThR.Tn[13] 0.063
R24080 XThR.Tn[13].n40 XThR.Tn[13] 0.063
R24081 XThR.Tn[13].n35 XThR.Tn[13] 0.063
R24082 XThR.Tn[13].n30 XThR.Tn[13] 0.063
R24083 XThR.Tn[13].n25 XThR.Tn[13] 0.063
R24084 XThR.Tn[13].n20 XThR.Tn[13] 0.063
R24085 XThR.Tn[13].n15 XThR.Tn[13] 0.063
R24086 XThR.Tn[13].n87 XThR.Tn[13] 0.0540714
R24087 XThR.Tn[13] XThR.Tn[13].n87 0.038
R24088 XThR.Tn[13].n11 XThR.Tn[13] 0.0143889
R24089 XThR.Tn[13].n85 XThR.Tn[13].n84 0.00771154
R24090 XThR.Tn[13].n80 XThR.Tn[13].n79 0.00771154
R24091 XThR.Tn[13].n75 XThR.Tn[13].n74 0.00771154
R24092 XThR.Tn[13].n70 XThR.Tn[13].n69 0.00771154
R24093 XThR.Tn[13].n65 XThR.Tn[13].n64 0.00771154
R24094 XThR.Tn[13].n60 XThR.Tn[13].n59 0.00771154
R24095 XThR.Tn[13].n55 XThR.Tn[13].n54 0.00771154
R24096 XThR.Tn[13].n50 XThR.Tn[13].n49 0.00771154
R24097 XThR.Tn[13].n45 XThR.Tn[13].n44 0.00771154
R24098 XThR.Tn[13].n40 XThR.Tn[13].n39 0.00771154
R24099 XThR.Tn[13].n35 XThR.Tn[13].n34 0.00771154
R24100 XThR.Tn[13].n30 XThR.Tn[13].n29 0.00771154
R24101 XThR.Tn[13].n25 XThR.Tn[13].n24 0.00771154
R24102 XThR.Tn[13].n20 XThR.Tn[13].n19 0.00771154
R24103 XThR.Tn[13].n15 XThR.Tn[13].n14 0.00771154
R24104 data[0].n1 data[0].t0 230.155
R24105 data[0].n0 data[0].t2 228.463
R24106 data[0].n1 data[0].t1 157.856
R24107 data[0].n0 data[0].t3 157.07
R24108 data[0].n2 data[0].n1 152.768
R24109 data[0].n4 data[0].n0 152.256
R24110 data[0].n3 data[0].n2 24.1398
R24111 data[0].n4 data[0].n3 9.48418
R24112 data[0] data[0].n4 6.1445
R24113 data[0].n2 data[0] 5.6325
R24114 data[0].n3 data[0] 2.638
R24115 data[6].n0 data[6].t0 230.576
R24116 data[6].n0 data[6].t1 158.275
R24117 data[6].n1 data[6].n0 152
R24118 data[6].n1 data[6] 11.9995
R24119 data[6] data[6].n1 6.66717
R24120 data[1].n4 data[1].t2 230.576
R24121 data[1].n1 data[1].t0 230.363
R24122 data[1].n0 data[1].t4 229.369
R24123 data[1].n4 data[1].t5 158.275
R24124 data[1].n1 data[1].t3 158.064
R24125 data[1].n0 data[1].t1 157.07
R24126 data[1].n2 data[1].n1 153.28
R24127 data[1].n7 data[1].n0 153.147
R24128 data[1].n5 data[1].n4 152
R24129 data[1].n7 data[1].n6 16.3874
R24130 data[1].n6 data[1].n5 14.9641
R24131 data[1].n3 data[1].n2 9.3005
R24132 data[1].n6 data[1].n3 6.49639
R24133 data[1] data[1].n7 3.24826
R24134 data[1].n2 data[1] 2.92621
R24135 data[1].n3 data[1] 2.15819
R24136 data[1].n5 data[1] 2.13383
R24137 data[2].n0 data[2].t0 230.576
R24138 data[2].n0 data[2].t1 158.275
R24139 data[2].n1 data[2].n0 152
R24140 data[2].n1 data[2] 12.7714
R24141 data[2] data[2].n1 2.13383
R24142 data[5].n4 data[5].t2 230.576
R24143 data[5].n1 data[5].t0 230.363
R24144 data[5].n0 data[5].t1 229.369
R24145 data[5].n4 data[5].t5 158.275
R24146 data[5].n1 data[5].t3 158.064
R24147 data[5].n0 data[5].t4 157.07
R24148 data[5].n2 data[5].n1 152.256
R24149 data[5].n7 data[5].n0 152.238
R24150 data[5].n5 data[5].n4 152
R24151 data[5].n7 data[5].n6 16.3874
R24152 data[5].n6 data[5].n5 14.6005
R24153 data[5].n3 data[5].n2 9.3005
R24154 data[5].n5 data[5] 6.66717
R24155 data[5].n6 data[5].n3 6.49639
R24156 data[5].n2 data[5] 6.1445
R24157 data[5] data[5].n7 5.68939
R24158 data[5].n3 data[5] 2.28319
R24159 bias[0] bias[0].t0 12.1467
R24160 bias[2].n0 bias[2].t0 56.8043
R24161 bias[2].n0 bias[2] 6.35112
R24162 bias[2] bias[2].n0 0.828709
R24163 data[3].n0 data[3].t1 230.576
R24164 data[3].n0 data[3].t0 158.275
R24165 data[3].n1 data[3].n0 153.553
R24166 data[3].n1 data[3] 11.6078
R24167 data[3] data[3].n1 2.90959
R24168 data[7].n0 data[7].t0 230.576
R24169 data[7].n0 data[7].t1 158.275
R24170 data[7].n1 data[7].n0 152
R24171 data[7].n1 data[7] 11.9995
R24172 data[7] data[7].n1 6.66717
R24173 bias[1] bias[1].t0 23.8076
C0 XA.XIR[15].XIC[8].icell.Ien Vbias 0.15966f
C1 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PDM 0.02601f
C2 XThC.XTB7.A data[0] 0.86893f
C3 XA.XIR[5].XIC[1].icell.Ien Iout 0.06801f
C4 XThC.Tn[7] XThC.Tn[8] 0.06603f
C5 XA.XIR[8].XIC[0].icell.PDM Vbias 0.03915f
C6 XA.XIR[4].XIC[11].icell.Ien Vbias 0.19161f
C7 XThR.Tn[14] Iout 1.12763f
C8 XThC.Tn[9] XA.XIR[7].XIC[9].icell.Ien 0.04604f
C9 XA.XIR[11].XIC[13].icell.PDM Vbias 0.03928f
C10 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout 0.06446f
C11 XA.XIR[2].XIC[4].icell.PDM Vbias 0.03928f
C12 XA.XIR[8].XIC[5].icell.Ien Vbias 0.19161f
C13 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PDM 0.04035f
C14 XA.XIR[10].XIC[12].icell.Ien Iout 0.06801f
C15 XThC.XTB6.Y VPWR 1.03165f
C16 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.Ien 0.04854f
C17 XA.XIR[14].XIC[14].icell.PDM Vbias 0.03928f
C18 XA.XIR[11].XIC_dummy_left.icell.Iout VPWR 0.10954f
C19 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.PDM 0.02104f
C20 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.02602f
C21 XA.XIR[5].XIC[10].icell.Ien VPWR 0.18829f
C22 XThC.XTBN.Y a_10051_9569# 0.23006f
C23 XThR.XTB7.A XThR.Tn[2] 0.12549f
C24 XA.XIR[9].XIC[14].icell.Ien Vbias 0.19161f
C25 XThR.XTB5.Y XThR.Tn[8] 0.01728f
C26 XThR.Tn[4] XA.XIR[4].XIC[1].icell.Ien 0.14211f
C27 XA.XIR[3].XIC[2].icell.PDM VPWR 0.01171f
C28 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.Ien 0.04854f
C29 XA.XIR[5].XIC[6].icell.Ien Iout 0.06801f
C30 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PDM 0.02601f
C31 XA.XIR[8].XIC[4].icell.PDM VPWR 0.01171f
C32 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10] 0.14211f
C33 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PDM 0.02601f
C34 XThR.Tn[3] XA.XIR[3].XIC[1].icell.Ien 0.14211f
C35 XA.XIR[2].XIC[8].icell.PDM VPWR 0.01171f
C36 XA.XIR[0].XIC[7].icell.Ien Vbias 0.19213f
C37 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PDM 0.0279f
C38 XA.XIR[12].XIC[5].icell.Ien VPWR 0.18829f
C39 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.Ien 0.04854f
C40 XThC.Tn[11] XA.XIR[9].XIC[11].icell.Ien 0.04604f
C41 XThC.Tn[4] XThR.Tn[14] 0.40738f
C42 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.Ien 0.04854f
C43 XA.XIR[7].XIC[10].icell.Ien Vbias 0.19161f
C44 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PDM 0.04035f
C45 XA.XIR[2].XIC_dummy_left.icell.Iout Iout 0.03553f
C46 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PDM 0.02601f
C47 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR 0.01691f
C48 XA.XIR[15].XIC[11].icell.Ien VPWR 0.31713f
C49 XThR.Tn[4] XA.XIR[4].XIC[6].icell.Ien 0.14211f
C50 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PDM 0.02601f
C51 XA.XIR[13].XIC[14].icell.Ien Iout 0.06801f
C52 XThC.XTB4.Y VPWR 0.91479f
C53 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.Ien 0.04854f
C54 XThC.Tn[12] XA.XIR[1].XIC[12].icell.Ien 0.04606f
C55 XA.XIR[8].XIC[0].icell.Ien Vbias 0.19149f
C56 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PDM 0.04035f
C57 XA.XIR[8].XIC_dummy_left.icell.Iout XA.XIR[9].XIC_dummy_left.icell.Iout 0.03665f
C58 XThC.XTB3.Y XThC.XTBN.A 0.03907f
C59 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout 0.06446f
C60 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PDM 0.04035f
C61 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Iout 0.03935f
C62 XThR.XTB5.A VPWR 0.83125f
C63 XThC.XTB5.A data[0] 0.14415f
C64 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PDM 0.04035f
C65 XA.XIR[7].XIC[4].icell.PDM Vbias 0.03928f
C66 XThR.XTB1.Y XThR.Tn[8] 0.29191f
C67 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PDM 0.0404f
C68 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR 0.08221f
C69 XA.XIR[15].XIC[2].icell.PDM Vbias 0.03928f
C70 XA.XIR[6].XIC[11].icell.PDM Vbias 0.03928f
C71 XA.XIR[10].XIC[10].icell.Ien Iout 0.06801f
C72 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.PDM 0.02104f
C73 XThR.Tn[12] XA.XIR[12].XIC[4].icell.Ien 0.14211f
C74 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PDM 0.02601f
C75 XThR.Tn[3] XA.XIR[3].XIC[9].icell.Ien 0.14211f
C76 XA.XIR[14].XIC[8].icell.PDM Vbias 0.03928f
C77 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PDM 0.02601f
C78 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PDM 0.02601f
C79 XThR.XTBN.Y XThR.XTB7.A 0.59539f
C80 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.Ien 0.04854f
C81 XA.XIR[9].XIC[0].icell.PDM Vbias 0.03915f
C82 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR 0.35722f
C83 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PDM 0.04035f
C84 XThC.Tn[9] XA.XIR[8].XIC[9].icell.Ien 0.04604f
C85 XA.XIR[7].XIC[8].icell.PDM VPWR 0.01171f
C86 XA.XIR[9].XIC[1].icell.Ien VPWR 0.18829f
C87 XThR.Tn[2] XA.XIR[2].XIC[4].icell.Ien 0.14211f
C88 XThC.Tn[6] XThR.Tn[13] 0.40738f
C89 XA.XIR[15].XIC[6].icell.PDM VPWR 0.01512f
C90 XA.XIR[4].XIC[3].icell.Ien VPWR 0.18829f
C91 VPWR data[5] 0.4402f
C92 XA.XIR[6].XIC_15.icell.PDM VPWR 0.07527f
C93 XThC.Tn[7] XA.XIR[15].XIC[7].icell.Ien 0.04292f
C94 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout 0.06446f
C95 XThC.Tn[0] Iout 0.07042f
C96 XA.XIR[11].XIC[12].icell.PDM Vbias 0.03928f
C97 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.PDM 0.02104f
C98 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.Ien 0.04854f
C99 XThC.Tn[0] XThR.Tn[9] 0.40738f
C100 XA.XIR[1].XIC[5].icell.PDM Vbias 0.03928f
C101 XA.XIR[3].XIC[7].icell.Ien Vbias 0.19161f
C102 XThC.Tn[5] XThR.Tn[8] 0.40738f
C103 XThR.XTB7.A XThR.XTB4.Y 0.14536f
C104 XThR.XTB2.Y XThR.XTB5.Y 0.0451f
C105 XA.XIR[14].XIC[13].icell.PDM Vbias 0.03928f
C106 XA.XIR[9].XIC[4].icell.PDM VPWR 0.01171f
C107 XThC.Tn[12] XA.XIR[6].XIC[12].icell.Ien 0.04604f
C108 XA.XIR[13].XIC[12].icell.Ien Iout 0.06801f
C109 XThC.Tn[3] XA.XIR[2].XIC[3].icell.Ien 0.04605f
C110 XThC.XTB2.Y VPWR 0.97668f
C111 XA.XIR[4].XIC[5].icell.PDM Vbias 0.03928f
C112 XThC.XTB5.Y XThC.XTB7.Y 0.036f
C113 XThC.XTB7.B XThC.XTB6.Y 0.30244f
C114 XA.XIR[9].XIC[6].icell.Ien VPWR 0.18829f
C115 XA.XIR[14].XIC_dummy_left.icell.Iout VPWR 0.10954f
C116 XA.XIR[1].XIC[2].icell.Ien Vbias 0.19173f
C117 XA.XIR[3].XIC[13].icell.PDM Vbias 0.03928f
C118 XA.XIR[8].XIC_15.icell.PDM Vbias 0.03927f
C119 XThC.Tn[0] XA.XIR[15].XIC[0].icell.Ien 0.04292f
C120 XA.XIR[9].XIC[2].icell.Ien Iout 0.06801f
C121 XThR.Tn[9] XA.XIR[9].XIC[2].icell.Ien 0.14211f
C122 XThC.XTB1.Y XThC.XTBN.A 0.12307f
C123 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.Ien 0.04854f
C124 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PDM 0.02601f
C125 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PDM 0.04035f
C126 XA.XIR[8].XIC[10].icell.Ien Vbias 0.19161f
C127 XThC.XTB3.Y XThC.Tn[2] 0.18399f
C128 XA.XIR[1].XIC[9].icell.PDM VPWR 0.01171f
C129 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PDM 0.02803f
C130 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.Ien 0.04854f
C131 XA.XIR[4].XIC[9].icell.PDM VPWR 0.01171f
C132 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PDM 0.02601f
C133 XA.XIR[5].XIC_15.icell.Ien VPWR 0.26829f
C134 XA.XIR[7].XIC[2].icell.Ien VPWR 0.18829f
C135 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PDM 0.04035f
C136 XThC.Tn[6] XThC.Tn[7] 0.0974f
C137 XA.XIR[5].XIC[11].icell.Ien Iout 0.06801f
C138 XThC.XTB7.Y XThC.XTBN.Y 0.50018f
C139 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.Ien 0.04854f
C140 XA.XIR[12].XIC_15.icell.PDM VPWR 0.07527f
C141 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR 0.01691f
C142 XA.XIR[0].XIC[12].icell.Ien Vbias 0.19213f
C143 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PDM 0.02601f
C144 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.04035f
C145 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.PDM 0.02104f
C146 XThC.XTB4.Y XThC.XTB7.B 0.33064f
C147 XThC.Tn[8] XThR.Tn[7] 0.40738f
C148 XThR.XTB1.Y XThR.XTB2.Y 2.14864f
C149 XA.XIR[12].XIC[6].icell.Ien Iout 0.06801f
C150 XA.XIR[7].XIC_15.icell.Ien Vbias 0.19195f
C151 XA.XIR[10].XIC_15.icell.Ien Iout 0.0694f
C152 VPWR Iout 57.8523f
C153 XA.XIR[5].XIC[0].icell.Ien Vbias 0.19149f
C154 XThC.XTB7.Y XThC.Tn[10] 0.07427f
C155 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PDM 0.04035f
C156 XThR.Tn[9] VPWR 8.97014f
C157 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.PDM 0.02104f
C158 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.04035f
C159 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.PDM 0.02104f
C160 XThR.Tn[4] XA.XIR[4].XIC[11].icell.Ien 0.14211f
C161 XA.XIR[5].XIC_dummy_right.icell.Iout VPWR 0.11567f
C162 XThC.Tn[14] Vbias 0.8291f
C163 XThR.Tn[0] XA.XIR[0].XIC[3].icell.Ien 0.14211f
C164 XThR.Tn[10] XA.XIR[10].XIC[2].icell.Ien 0.14211f
C165 XThR.XTB7.B XThR.XTBN.Y 0.3875f
C166 XA.XIR[13].XIC[10].icell.Ien Iout 0.06801f
C167 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PDM 0.04035f
C168 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.04056f
C169 XThR.Tn[7] XA.XIR[7].XIC[4].icell.Ien 0.14211f
C170 XA.XIR[6].XIC[2].icell.Ien Vbias 0.19161f
C171 XA.XIR[15].XIC[0].icell.Ien VPWR 0.31713f
C172 XThC.Tn[11] XA.XIR[10].XIC[11].icell.Ien 0.04604f
C173 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.PDM 0.02104f
C174 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.Ien 0.04854f
C175 XThC.XTB1.Y XThC.XTB3.Y 0.04033f
C176 XA.XIR[10].XIC_dummy_right.icell.Iout Iout 0.01732f
C177 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PDM 0.02601f
C178 XA.XIR[11].XIC[11].icell.PDM Vbias 0.03928f
C179 XThR.Tn[12] XA.XIR[12].XIC[9].icell.Ien 0.14211f
C180 XA.XIR[10].XIC[3].icell.PDM VPWR 0.01171f
C181 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.PDM 0.02104f
C182 XThC.Tn[4] VPWR 3.6464f
C183 XThR.Tn[3] XA.XIR[3].XIC[14].icell.Ien 0.144f
C184 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.Ien 0.04854f
C185 XThR.XTB7.B XThR.XTB4.Y 0.33064f
C186 XA.XIR[14].XIC[12].icell.PDM Vbias 0.03928f
C187 XA.XIR[9].XIC_15.icell.PDM Vbias 0.03927f
C188 XThR.XTBN.Y XThR.Tn[2] 0.6189f
C189 XThC.Tn[10] XThR.Tn[0] 0.40762f
C190 XA.XIR[15].XIC[5].icell.Ien VPWR 0.31713f
C191 XA.XIR[0].XIC[7].icell.PDM Vbias 0.03945f
C192 XThC.Tn[12] XThR.Tn[5] 0.40738f
C193 XThR.XTB7.B XThR.Tn[10] 0.06102f
C194 XThC.XTB7.B a_7875_9569# 0.01174f
C195 XThR.Tn[2] XA.XIR[2].XIC[9].icell.Ien 0.14211f
C196 XA.XIR[4].XIC[8].icell.Ien VPWR 0.18829f
C197 XA.XIR[10].XIC[3].icell.Ien Vbias 0.19161f
C198 XThC.XTB6.A XThC.XTB5.Y 0.01866f
C199 XThC.XTB2.Y XThC.XTB7.B 0.22599f
C200 XA.XIR[4].XIC[4].icell.Ien Iout 0.06801f
C201 a_8963_9569# XThC.Tn[11] 0.1927f
C202 XA.XIR[8].XIC[2].icell.Ien VPWR 0.18829f
C203 XA.XIR[3].XIC[12].icell.Ien Vbias 0.19161f
C204 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.Ien 0.04854f
C205 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13] 0.14211f
C206 XA.XIR[0].XIC[11].icell.PDM VPWR 0.01132f
C207 XThC.Tn[2] XA.XIR[0].XIC[2].icell.Ien 0.04658f
C208 XA.XIR[2].XIC[5].icell.Ien Vbias 0.19161f
C209 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.Ien 0.04854f
C210 XA.XIR[9].XIC[11].icell.Ien VPWR 0.18829f
C211 XA.XIR[1].XIC[7].icell.Ien Vbias 0.19173f
C212 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.PDM 0.02104f
C213 XA.XIR[12].XIC[14].icell.PDM VPWR 0.0118f
C214 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.PDM 0.02104f
C215 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PDM 0.02602f
C216 XA.XIR[9].XIC[7].icell.Ien Iout 0.06801f
C217 XThR.Tn[9] XA.XIR[9].XIC[7].icell.Ien 0.14211f
C218 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PDM 0.04035f
C219 XThC.XTB6.A XThC.XTBN.Y 0.03867f
C220 XA.XIR[0].XIC[4].icell.Ien VPWR 0.18788f
C221 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PDM 0.04035f
C222 XA.XIR[8].XIC_15.icell.Ien Vbias 0.19195f
C223 XThC.Tn[9] XThR.Tn[2] 0.40741f
C224 XA.XIR[15].XIC_15.icell.PDM VPWR 0.07867f
C225 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PDM 0.02601f
C226 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.PDM 0.02104f
C227 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.Ien 0.04854f
C228 XThC.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.04604f
C229 XA.XIR[7].XIC[7].icell.Ien VPWR 0.18829f
C230 XThR.XTB5.Y XThR.XTB7.Y 0.036f
C231 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.04035f
C232 XA.XIR[7].XIC[3].icell.Ien Iout 0.06801f
C233 XA.XIR[7].XIC_dummy_left.icell.Ien XThR.Tn[7] 0.01256f
C234 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.PDM 0.02104f
C235 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.Ien 0.04854f
C236 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PDM 0.02601f
C237 XA.XIR[13].XIC_15.icell.Ien Iout 0.0694f
C238 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.Ien 0.04854f
C239 XThC.XTB7.A XThC.Tn[5] 0.02777f
C240 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR 0.38922f
C241 XA.XIR[5].XIC[5].icell.PDM Vbias 0.03928f
C242 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.PDM 0.02104f
C243 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PDM 0.0404f
C244 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.Ien 0.04854f
C245 data[1] data[0] 0.64735f
C246 XThC.Tn[14] XA.XIR[11].XIC[14].icell.Ien 0.04604f
C247 XThR.Tn[11] XA.XIR[11].XIC[3].icell.Ien 0.14211f
C248 XThC.Tn[14] XThR.Tn[6] 0.40742f
C249 XA.XIR[12].XIC[4].icell.PDM Vbias 0.03928f
C250 XThR.Tn[12] XA.XIR[12].XIC[14].icell.Ien 0.144f
C251 XA.XIR[11].XIC[10].icell.PDM Vbias 0.03928f
C252 a_6243_9615# VPWR 0.7055f
C253 XA.XIR[6].XIC[2].icell.PDM VPWR 0.01171f
C254 XThR.Tn[0] XA.XIR[0].XIC[8].icell.Ien 0.14211f
C255 XThC.Tn[11] XA.XIR[13].XIC[11].icell.Ien 0.04604f
C256 XThR.Tn[10] XA.XIR[10].XIC[7].icell.Ien 0.14211f
C257 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.Ien 0.04854f
C258 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PDM 0.04035f
C259 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.Ien 0.04854f
C260 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PDM 0.02601f
C261 XA.XIR[5].XIC[9].icell.PDM VPWR 0.01171f
C262 XThR.Tn[6] XA.XIR[6].XIC[2].icell.Ien 0.14211f
C263 XThR.XTBN.Y XThR.XTB4.Y 0.15627f
C264 XA.XIR[13].XIC_dummy_right.icell.Iout Iout 0.01732f
C265 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.02601f
C266 XA.XIR[14].XIC[11].icell.PDM Vbias 0.03928f
C267 XThC.Tn[6] XThR.Tn[7] 0.40738f
C268 XA.XIR[11].XIC_dummy_left.icell.Iout XA.XIR[12].XIC_dummy_left.icell.Iout 0.03665f
C269 XA.XIR[13].XIC[3].icell.PDM VPWR 0.01171f
C270 XA.XIR[6].XIC[7].icell.Ien Vbias 0.19161f
C271 XThR.Tn[7] XA.XIR[7].XIC[9].icell.Ien 0.14211f
C272 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PDM 0.02805f
C273 XThR.XTBN.Y XThR.Tn[10] 0.46535f
C274 XThC.XTB5.Y XThC.Tn[8] 0.0173f
C275 XThR.XTB1.Y data[4] 0.06453f
C276 XA.XIR[12].XIC[8].icell.PDM VPWR 0.01171f
C277 XThR.XTB1.Y XThR.XTB7.Y 0.05211f
C278 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PDM 0.02601f
C279 XThC.Tn[3] Vbias 0.84088f
C280 XThC.XTB6.Y XThC.Tn[12] 0.0253f
C281 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.Ien 0.04854f
C282 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.Ien 0.04854f
C283 XA.XIR[15].XIC[1].icell.Ien Iout 0.07192f
C284 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.Ien 0.04854f
C285 XThC.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.04604f
C286 XA.XIR[5].XIC_dummy_left.icell.Iout Iout 0.03553f
C287 XA.XIR[3].XIC[0].icell.PDM Vbias 0.03915f
C288 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.Ien 0.04854f
C289 XA.XIR[8].XIC[2].icell.PDM Vbias 0.03928f
C290 XThC.Tn[10] XThR.Tn[1] 0.40744f
C291 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PDM 0.02601f
C292 XThC.Tn[9] XA.XIR[2].XIC[9].icell.Ien 0.04605f
C293 a_5949_9615# XThC.Tn[5] 0.26251f
C294 XA.XIR[2].XIC[6].icell.PDM Vbias 0.03928f
C295 XA.XIR[13].XIC[3].icell.Ien Vbias 0.19161f
C296 XA.XIR[10].XIC[13].icell.Ien VPWR 0.18829f
C297 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PDM 0.04035f
C298 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR 0.01691f
C299 XA.XIR[3].XIC[4].icell.Ien VPWR 0.18829f
C300 XThC.Tn[10] XThR.Tn[12] 0.40738f
C301 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.02601f
C302 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.PDM 0.02104f
C303 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.Ien 0.04854f
C304 XThR.XTB4.Y XThR.Tn[10] 0.01391f
C305 XA.XIR[11].XIC[6].icell.Ien Vbias 0.19161f
C306 XThC.Tn[5] XThR.Tn[3] 0.40738f
C307 XThR.Tn[2] XA.XIR[2].XIC[14].icell.Ien 0.144f
C308 XThC.XTBN.Y XThC.Tn[8] 0.41222f
C309 XA.XIR[6].XIC_dummy_right.icell.Iout XA.XIR[7].XIC_dummy_right.icell.Iout 0.04047f
C310 XA.XIR[15].XIC[6].icell.Ien Iout 0.07192f
C311 XA.XIR[4].XIC[13].icell.Ien VPWR 0.18829f
C312 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Iout 0.03908f
C313 XA.XIR[10].XIC[8].icell.Ien Vbias 0.19161f
C314 XA.XIR[3].XIC[4].icell.PDM VPWR 0.01171f
C315 XA.XIR[12].XIC[13].icell.PDM VPWR 0.01171f
C316 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.PDM 0.02104f
C317 XThC.XTB1.Y a_2979_9615# 0.21263f
C318 XA.XIR[8].XIC[6].icell.PDM VPWR 0.01171f
C319 XThC.Tn[14] XThR.Tn[4] 0.40742f
C320 XA.XIR[2].XIC[10].icell.PDM VPWR 0.01171f
C321 XA.XIR[4].XIC[9].icell.Ien Iout 0.06801f
C322 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Iout 0.03843f
C323 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.PDM 0.02104f
C324 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PDM 0.02602f
C325 XA.XIR[0].XIC[0].icell.Ien Iout 0.06743f
C326 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PDM 0.04041f
C327 XThR.XTB5.Y XThR.Tn[11] 0.02067f
C328 XA.XIR[15].XIC[14].icell.PDM VPWR 0.01521f
C329 XA.XIR[8].XIC[7].icell.Ien VPWR 0.18829f
C330 XThC.Tn[9] XThR.Tn[10] 0.40738f
C331 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.PDM 0.02104f
C332 XThC.Tn[1] XThR.Tn[5] 0.40738f
C333 XA.XIR[8].XIC[3].icell.Ien Iout 0.06801f
C334 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PDM 0.02601f
C335 XThR.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.14211f
C336 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.Ien 0.04854f
C337 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.Ien 0.04854f
C338 XA.XIR[2].XIC[10].icell.Ien Vbias 0.19161f
C339 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PDM 0.02601f
C340 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PDM 0.04035f
C341 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR 0.35722f
C342 XThC.Tn[13] XThC.Tn[14] 0.3543f
C343 XA.XIR[1].XIC[12].icell.Ien Vbias 0.19173f
C344 XA.XIR[9].XIC[12].icell.Ien Iout 0.06801f
C345 XThR.Tn[9] XA.XIR[9].XIC[12].icell.Ien 0.14211f
C346 XA.XIR[0].XIC[9].icell.Ien VPWR 0.18925f
C347 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR 0.01604f
C348 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PDM 0.02601f
C349 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.PDM 0.02104f
C350 XA.XIR[0].XIC[5].icell.Ien Iout 0.0675f
C351 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PDM 0.04035f
C352 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PDM 0.04035f
C353 XThR.XTBN.Y a_n997_1803# 0.22873f
C354 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PDM 0.04035f
C355 XA.XIR[7].XIC[12].icell.Ien VPWR 0.18829f
C356 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.PDM 0.02104f
C357 XThR.Tn[13] XA.XIR[13].XIC[2].icell.Ien 0.14211f
C358 XA.XIR[7].XIC[8].icell.Ien Iout 0.06801f
C359 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PDM 0.04035f
C360 XA.XIR[7].XIC[6].icell.PDM Vbias 0.03928f
C361 XThC.Tn[3] XA.XIR[5].XIC[3].icell.Ien 0.04604f
C362 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.Ien 0.04854f
C363 XThC.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.04604f
C364 XA.XIR[15].XIC[4].icell.PDM Vbias 0.03928f
C365 XThR.XTB6.A XThR.XTB2.Y 0.18237f
C366 XA.XIR[6].XIC[13].icell.PDM Vbias 0.03928f
C367 XA.XIR[10].XIC[11].icell.Ien VPWR 0.18829f
C368 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.Ien 0.04854f
C369 XThC.Tn[7] XThR.Tn[2] 0.40741f
C370 XA.XIR[3].XIC[1].icell.Ien VPWR 0.18829f
C371 XThC.XTB7.B a_6243_9615# 0.01743f
C372 XA.XIR[14].XIC[10].icell.PDM Vbias 0.03928f
C373 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PDM 0.02601f
C374 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.PDM 0.02104f
C375 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout 0.06446f
C376 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PDM 0.02601f
C377 XThR.Tn[11] XA.XIR[11].XIC[8].icell.Ien 0.14211f
C378 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PDM 0.0404f
C379 XA.XIR[9].XIC[2].icell.PDM Vbias 0.03928f
C380 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PDM 0.02804f
C381 XA.XIR[7].XIC[10].icell.PDM VPWR 0.01171f
C382 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.PDM 0.02104f
C383 XA.XIR[9].XIC_dummy_left.icell.Iout VPWR 0.10954f
C384 XThR.XTBN.Y XThR.Tn[13] 0.56841f
C385 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PDM 0.02601f
C386 XA.XIR[12].XIC[13].icell.Ien Vbias 0.19161f
C387 XA.XIR[15].XIC[8].icell.PDM VPWR 0.01512f
C388 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.PDM 0.02104f
C389 XThR.Tn[0] XA.XIR[0].XIC[13].icell.Ien 0.14211f
C390 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.PDM 0.02104f
C391 XA.XIR[10].XIC[0].icell.Ien Iout 0.06795f
C392 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.Ien 0.04854f
C393 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.PDM 0.02104f
C394 XThR.Tn[6] XA.XIR[6].XIC[7].icell.Ien 0.14211f
C395 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.PDM 0.02104f
C396 XThR.Tn[12] XA.XIR[12].XIC[10].icell.Ien 0.14211f
C397 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.PDM 0.02104f
C398 XA.XIR[0].XIC_dummy_left.icell.Iout XA.XIR[1].XIC_dummy_left.icell.Iout 0.03665f
C399 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PDM 0.02601f
C400 XThC.Tn[3] XThR.Tn[6] 0.40738f
C401 XA.XIR[1].XIC[7].icell.PDM Vbias 0.03928f
C402 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.PDM 0.02104f
C403 XA.XIR[6].XIC[12].icell.Ien Vbias 0.19161f
C404 XThR.Tn[7] XA.XIR[7].XIC[14].icell.Ien 0.144f
C405 XA.XIR[9].XIC[6].icell.PDM VPWR 0.01171f
C406 VPWR data[0] 0.52929f
C407 XA.XIR[13].XIC[13].icell.Ien VPWR 0.18829f
C408 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.Ien 0.04854f
C409 XA.XIR[4].XIC[7].icell.PDM Vbias 0.03928f
C410 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PDM 0.02601f
C411 XThC.Tn[5] XThR.Tn[11] 0.40738f
C412 XA.XIR[12].XIC[12].icell.PDM VPWR 0.01171f
C413 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.Ien 0.04854f
C414 XA.XIR[3].XIC_15.icell.PDM Vbias 0.03927f
C415 XA.XIR[14].XIC[6].icell.Ien Vbias 0.19161f
C416 XThC.XTB7.A XThC.XTB7.Y 0.37429f
C417 XThC.Tn[8] XA.XIR[0].XIC[8].icell.Ien 0.04654f
C418 XA.XIR[13].XIC[8].icell.Ien Vbias 0.19161f
C419 XA.XIR[15].XIC[13].icell.PDM VPWR 0.01512f
C420 XThC.Tn[7] XA.XIR[10].XIC[7].icell.Ien 0.04604f
C421 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PDM 0.04035f
C422 XA.XIR[3].XIC[9].icell.Ien VPWR 0.18829f
C423 XA.XIR[1].XIC[11].icell.PDM VPWR 0.01171f
C424 XThC.Tn[2] XA.XIR[1].XIC[2].icell.Ien 0.04606f
C425 XA.XIR[12].XIC_dummy_left.icell.Iout Iout 0.03553f
C426 XA.XIR[3].XIC[5].icell.Ien Iout 0.06801f
C427 XThC.Tn[9] XThR.Tn[13] 0.40738f
C428 XA.XIR[4].XIC[11].icell.PDM VPWR 0.01171f
C429 XA.XIR[2].XIC[2].icell.Ien VPWR 0.18829f
C430 XA.XIR[2].XIC_dummy_right.icell.Iout XA.XIR[3].XIC_dummy_right.icell.Iout 0.04047f
C431 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.PDM 0.02104f
C432 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PDM 0.04035f
C433 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PDM 0.02601f
C434 XA.XIR[1].XIC[4].icell.Ien VPWR 0.18829f
C435 XThC.Tn[12] Iout 0.2243f
C436 XThC.Tn[12] XThR.Tn[9] 0.40738f
C437 XThC.Tn[10] XA.XIR[4].XIC[10].icell.Ien 0.04604f
C438 XA.XIR[4].XIC[14].icell.Ien Iout 0.06801f
C439 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PDM 0.04035f
C440 XThC.Tn[8] XThR.Tn[8] 0.40738f
C441 XA.XIR[8].XIC[12].icell.Ien VPWR 0.18829f
C442 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PDM 0.04035f
C443 XA.XIR[8].XIC[8].icell.Ien Iout 0.06801f
C444 XThC.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.04604f
C445 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.Ien 0.04854f
C446 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.PDM 0.02104f
C447 XA.XIR[2].XIC_15.icell.Ien Vbias 0.19195f
C448 XA.XIR[12].XIC[11].icell.Ien Vbias 0.19161f
C449 XThC.XTBN.Y XThC.Tn[6] 0.49549f
C450 XThC.Tn[3] XThR.Tn[4] 0.40738f
C451 XThR.XTB7.B a_n997_3979# 0.01152f
C452 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.Ien 0.04854f
C453 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PDM 0.04035f
C454 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.Ien 0.04854f
C455 XA.XIR[0].XIC[14].icell.Ien VPWR 0.18783f
C456 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.Ien 0.04854f
C457 XThC.Tn[7] XThR.Tn[10] 0.40738f
C458 XThR.Tn[14] XA.XIR[14].XIC[3].icell.Ien 0.14211f
C459 XA.XIR[10].XIC[1].icell.PDM Vbias 0.03928f
C460 XA.XIR[0].XIC[10].icell.Ien Iout 0.0675f
C461 XThR.Tn[1] XA.XIR[1].XIC[3].icell.Ien 0.14211f
C462 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.PDM 0.02104f
C463 XA.XIR[13].XIC[11].icell.Ien VPWR 0.18829f
C464 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.04035f
C465 a_7651_9569# XThC.Tn[8] 0.1927f
C466 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PDM 0.02601f
C467 XThR.Tn[13] XA.XIR[13].XIC[7].icell.Ien 0.14211f
C468 XA.XIR[7].XIC[13].icell.Ien Iout 0.06801f
C469 XA.XIR[5].XIC[5].icell.Ien Vbias 0.19161f
C470 XThR.Tn[12] XA.XIR[12].XIC_15.icell.Ien 0.13564f
C471 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.Ien 0.04854f
C472 XA.XIR[11].XIC[1].icell.PDM VPWR 0.01171f
C473 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PDM 0.02601f
C474 XThC.Tn[2] XA.XIR[6].XIC[2].icell.Ien 0.04604f
C475 XA.XIR[10].XIC[5].icell.PDM VPWR 0.01171f
C476 XThR.XTB2.Y XThR.Tn[1] 0.17876f
C477 XThC.Tn[8] XA.XIR[3].XIC[8].icell.Ien 0.04604f
C478 XA.XIR[13].XIC[0].icell.Ien Iout 0.06795f
C479 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PDM 0.02602f
C480 XA.XIR[6].XIC[4].icell.Ien VPWR 0.18829f
C481 XThR.Tn[5] Vbias 1.39526f
C482 XThC.Tn[3] XA.XIR[12].XIC[3].icell.Ien 0.04604f
C483 XThR.XTB7.B XThR.Tn[7] 0.07415f
C484 XThR.XTB7.B a_n997_2891# 0.0168f
C485 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PDM 0.02601f
C486 XA.XIR[0].XIC[9].icell.PDM Vbias 0.03945f
C487 XThC.Tn[1] XA.XIR[9].XIC[1].icell.Ien 0.04604f
C488 XA.XIR[12].XIC[11].icell.PDM VPWR 0.01171f
C489 XThC.XTB7.B a_8963_9569# 0.02071f
C490 XThC.XTB7.B data[0] 0.0138f
C491 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.Ien 0.04854f
C492 XThC.Tn[5] XThR.Tn[14] 0.40738f
C493 XThR.Tn[6] XA.XIR[6].XIC[12].icell.Ien 0.14211f
C494 XA.XIR[15].XIC[12].icell.PDM VPWR 0.01512f
C495 XThC.XTB6.A XThC.XTB7.A 0.44014f
C496 XThR.XTB6.A data[4] 0.48493f
C497 XThR.XTB6.A XThR.XTB7.Y 0.01596f
C498 XThR.XTB3.Y XThR.XTB5.Y 0.04438f
C499 XThC.Tn[7] XA.XIR[13].XIC[7].icell.Ien 0.04604f
C500 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.PDM 0.02104f
C501 XA.XIR[0].XIC[13].icell.PDM VPWR 0.01132f
C502 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.Ien 0.04854f
C503 XA.XIR[11].XIC[3].icell.Ien VPWR 0.18829f
C504 XThC.XTB2.Y XThC.Tn[1] 0.18085f
C505 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.PDM 0.02104f
C506 XA.XIR[10].XIC[5].icell.Ien VPWR 0.18829f
C507 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout 0.06446f
C508 XThC.Tn[6] XA.XIR[8].XIC[6].icell.Ien 0.04604f
C509 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PDM 0.04035f
C510 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.Ien 0.04854f
C511 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PDM 0.04035f
C512 XA.XIR[3].XIC[14].icell.Ien VPWR 0.18835f
C513 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PDM 0.02601f
C514 XThR.XTBN.Y a_n997_3979# 0.23021f
C515 XA.XIR[3].XIC[10].icell.Ien Iout 0.06801f
C516 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.Ien 0.04854f
C517 XA.XIR[2].XIC[7].icell.Ien VPWR 0.18829f
C518 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PDM 0.04056f
C519 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.PDM 0.02104f
C520 XA.XIR[2].XIC[3].icell.Ien Iout 0.06801f
C521 XA.XIR[1].XIC[9].icell.Ien VPWR 0.18829f
C522 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PDM 0.02601f
C523 XThR.Tn[8] XA.XIR[8].XIC[4].icell.Ien 0.14211f
C524 XA.XIR[14].XIC_dummy_left.icell.Iout XA.XIR[15].XIC_dummy_left.icell.Iout 0.03665f
C525 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PDM 0.02601f
C526 XA.XIR[1].XIC[5].icell.Ien Iout 0.06801f
C527 XA.XIR[6].XIC[0].icell.PDM Vbias 0.03915f
C528 XA.XIR[2].XIC_dummy_left.icell.Iout XA.XIR[3].XIC_dummy_left.icell.Iout 0.03665f
C529 XA.XIR[15].XIC[13].icell.Ien Vbias 0.15966f
C530 XA.XIR[1].XIC_dummy_right.icell.Iout XA.XIR[2].XIC_dummy_right.icell.Iout 0.04047f
C531 XThC.Tn[9] XA.XIR[5].XIC[9].icell.Ien 0.04604f
C532 XThC.XTB3.Y a_4067_9615# 0.23056f
C533 XThR.XTB1.Y XThR.XTB3.Y 0.04033f
C534 XA.XIR[5].XIC[7].icell.PDM Vbias 0.03928f
C535 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.Ien 0.04854f
C536 XA.XIR[8].XIC[13].icell.Ien Iout 0.06801f
C537 XThC.Tn[7] XThR.Tn[13] 0.40738f
C538 a_4067_9615# XThC.Tn[2] 0.27296f
C539 XA.XIR[13].XIC[1].icell.PDM Vbias 0.03928f
C540 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PDM 0.02601f
C541 XThR.Tn[5] XA.XIR[5].XIC[3].icell.Ien 0.14211f
C542 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PDM 0.0404f
C543 XThC.Tn[13] XA.XIR[12].XIC[13].icell.Ien 0.04604f
C544 XThC.Tn[1] Iout 0.22482f
C545 XA.XIR[12].XIC[6].icell.PDM Vbias 0.03928f
C546 XThC.Tn[1] XThR.Tn[9] 0.40738f
C547 XThC.XTB5.A XThC.XTB6.A 1.80461f
C548 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout 0.06446f
C549 XA.XIR[6].XIC[4].icell.PDM VPWR 0.01171f
C550 XThC.Tn[6] XThR.Tn[8] 0.40738f
C551 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PDM 0.04056f
C552 XThR.XTB7.A a_n1049_6699# 0.02294f
C553 XThR.Tn[1] XA.XIR[1].XIC[8].icell.Ien 0.14211f
C554 XThR.Tn[14] XA.XIR[14].XIC[8].icell.Ien 0.14211f
C555 XA.XIR[0].XIC_15.icell.Ien Iout 0.06774f
C556 XThR.XTB5.Y VPWR 1.0269f
C557 XA.XIR[14].XIC[1].icell.PDM VPWR 0.01171f
C558 XA.XIR[5].XIC[11].icell.PDM VPWR 0.01171f
C559 XThR.XTBN.Y XThR.Tn[7] 0.89994f
C560 XThR.XTBN.Y a_n997_2891# 0.22804f
C561 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PDM 0.02602f
C562 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.Ien 0.04854f
C563 XA.XIR[13].XIC[5].icell.PDM VPWR 0.01171f
C564 XThC.XTB6.Y Vbias 0.01779f
C565 XA.XIR[6].XIC[0].icell.Ien Iout 0.06795f
C566 XA.XIR[12].XIC[10].icell.PDM VPWR 0.01171f
C567 XA.XIR[5].XIC[10].icell.Ien Vbias 0.19161f
C568 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.02601f
C569 XA.XIR[15].XIC_dummy_left.icell.Iout Iout 0.03553f
C570 XThC.XTB3.Y XThC.Tn[3] 0.01335f
C571 XA.XIR[3].XIC[2].icell.PDM Vbias 0.03928f
C572 XA.XIR[8].XIC[4].icell.PDM Vbias 0.03928f
C573 XA.XIR[15].XIC[11].icell.PDM VPWR 0.01512f
C574 XThR.Tn[5] XThR.Tn[6] 0.11432f
C575 XThC.Tn[2] XThC.Tn[3] 0.59596f
C576 XA.XIR[2].XIC[8].icell.PDM Vbias 0.03928f
C577 XThR.XTB4.Y XThR.Tn[7] 0.01797f
C578 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PDM 0.04035f
C579 XA.XIR[0].XIC_dummy_right.icell.Iout Iout 0.01732f
C580 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PDM 0.02601f
C581 XA.XIR[12].XIC[5].icell.Ien Vbias 0.19161f
C582 XA.XIR[6].XIC[9].icell.Ien VPWR 0.18829f
C583 XA.XIR[6].XIC[5].icell.Ien Iout 0.06801f
C584 XThR.Tn[10] a_n997_2891# 0.1927f
C585 XThC.Tn[8] XA.XIR[1].XIC[8].icell.Ien 0.04606f
C586 XA.XIR[15].XIC[11].icell.Ien Vbias 0.15966f
C587 XA.XIR[8].XIC[8].icell.PDM VPWR 0.01171f
C588 XA.XIR[3].XIC[6].icell.PDM VPWR 0.01171f
C589 XA.XIR[14].XIC[3].icell.Ien VPWR 0.18883f
C590 XThC.Tn[9] XThR.Tn[7] 0.40738f
C591 XThC.XTB4.Y Vbias 0.01644f
C592 XA.XIR[2].XIC[12].icell.PDM VPWR 0.01171f
C593 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.PDM 0.02104f
C594 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PDM 0.04035f
C595 XA.XIR[13].XIC[5].icell.Ien VPWR 0.18829f
C596 XThR.XTB1.Y VPWR 1.13148f
C597 XThC.XTB2.Y a_3523_10575# 0.01006f
C598 XThC.XTB7.Y XThC.Tn[11] 0.07422f
C599 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.Ien 0.04854f
C600 XThR.XTB6.Y a_n1319_5611# 0.01283f
C601 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.PDM 0.02104f
C602 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR 0.01691f
C603 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PDM 0.0404f
C604 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PDM 0.02601f
C605 XA.XIR[11].XIC[8].icell.Ien VPWR 0.18829f
C606 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PDM 0.02601f
C607 XA.XIR[11].XIC[4].icell.Ien Iout 0.06801f
C608 XThR.XTB7.Y XThR.Tn[12] 0.07066f
C609 XThC.Tn[12] XA.XIR[7].XIC[12].icell.Ien 0.04604f
C610 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.02804f
C611 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.Ien 0.04854f
C612 XA.XIR[10].XIC[6].icell.Ien Iout 0.06801f
C613 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PDM 0.02601f
C614 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PDM 0.02601f
C615 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PDM 0.04035f
C616 XThR.Tn[4] XThR.Tn[5] 0.12171f
C617 XA.XIR[3].XIC_15.icell.Ien Iout 0.0694f
C618 XThC.Tn[8] XThR.Tn[3] 0.40738f
C619 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PDM 0.04035f
C620 XA.XIR[2].XIC[12].icell.Ien VPWR 0.18829f
C621 XThC.Tn[3] XA.XIR[15].XIC[3].icell.Ien 0.04292f
C622 XA.XIR[2].XIC[8].icell.Ien Iout 0.06801f
C623 XA.XIR[1].XIC[14].icell.Ien VPWR 0.18835f
C624 XThC.Tn[5] VPWR 3.59867f
C625 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PDM 0.04056f
C626 XA.XIR[7].XIC[8].icell.PDM Vbias 0.03928f
C627 XThR.Tn[8] XA.XIR[8].XIC[9].icell.Ien 0.14211f
C628 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PDM 0.02601f
C629 XA.XIR[9].XIC[1].icell.Ien Vbias 0.19161f
C630 XA.XIR[1].XIC[10].icell.Ien Iout 0.06801f
C631 XA.XIR[4].XIC[3].icell.Ien Vbias 0.19161f
C632 XA.XIR[6].XIC_15.icell.PDM Vbias 0.03927f
C633 XA.XIR[15].XIC[6].icell.PDM Vbias 0.03928f
C634 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.PDM 0.02104f
C635 XA.XIR[3].XIC_dummy_left.icell.Iout VPWR 0.11229f
C636 XThR.XTB6.Y XThR.Tn[5] 0.20186f
C637 XThC.Tn[11] XThR.Tn[0] 0.40763f
C638 XThC.Tn[14] XA.XIR[9].XIC[14].icell.Ien 0.04604f
C639 XThC.Tn[13] XThR.Tn[5] 0.40739f
C640 XThC.Tn[4] XA.XIR[11].XIC[4].icell.Ien 0.04604f
C641 XA.XIR[12].XIC[1].icell.Ien VPWR 0.18829f
C642 XThC.Tn[8] XA.XIR[6].XIC[8].icell.Ien 0.04604f
C643 XThR.Tn[5] XA.XIR[5].XIC[8].icell.Ien 0.14211f
C644 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.Ien 0.04854f
C645 XA.XIR[9].XIC[4].icell.PDM Vbias 0.03928f
C646 XThR.XTBN.Y a_n997_1579# 0.23006f
C647 XA.XIR[3].XIC_dummy_right.icell.Iout Iout 0.01732f
C648 XThR.XTB7.Y a_n1049_5317# 0.27822f
C649 XA.XIR[5].XIC[2].icell.Ien VPWR 0.18829f
C650 XThC.XTB2.Y Vbias 0.01484f
C651 XA.XIR[7].XIC[12].icell.PDM VPWR 0.01171f
C652 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout 0.06446f
C653 XThC.Tn[9] XA.XIR[12].XIC[9].icell.Ien 0.04604f
C654 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.PDM 0.02104f
C655 XA.XIR[9].XIC[6].icell.Ien Vbias 0.19161f
C656 XA.XIR[15].XIC[10].icell.PDM VPWR 0.01512f
C657 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PDM 0.02601f
C658 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PDM 0.02601f
C659 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.Ien 0.04854f
C660 XThR.Tn[1] XA.XIR[1].XIC[13].icell.Ien 0.14211f
C661 XA.XIR[1].XIC[9].icell.PDM Vbias 0.03928f
C662 XA.XIR[9].XIC[8].icell.PDM VPWR 0.01171f
C663 XA.XIR[0].XIC[0].icell.PDM VPWR 0.01132f
C664 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.Ien 0.04854f
C665 XA.XIR[7].XIC[2].icell.Ien Vbias 0.19161f
C666 XA.XIR[4].XIC[9].icell.PDM Vbias 0.03928f
C667 XA.XIR[5].XIC_15.icell.Ien Vbias 0.19195f
C668 XThC.Tn[10] XThR.Tn[2] 0.40741f
C669 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12] 0.14211f
C670 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.Ien 0.04854f
C671 XA.XIR[12].XIC_15.icell.PDM Vbias 0.03927f
C672 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PDM 0.04035f
C673 XThR.Tn[11] XThR.Tn[12] 0.1626f
C674 XA.XIR[1].XIC[13].icell.PDM VPWR 0.01171f
C675 XA.XIR[6].XIC[14].icell.Ien VPWR 0.18835f
C676 XThC.Tn[12] XA.XIR[8].XIC[12].icell.Ien 0.04604f
C677 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PDM 0.04035f
C678 XA.XIR[6].XIC[10].icell.Ien Iout 0.06801f
C679 XA.XIR[4].XIC[13].icell.PDM VPWR 0.01171f
C680 XThC.XTB7.A XThC.Tn[6] 0.10502f
C681 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PDM 0.04035f
C682 Vbias Iout 74.00211f
C683 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR 0.01691f
C684 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PDM 0.02601f
C685 XThR.Tn[9] Vbias 1.39532f
C686 XA.XIR[14].XIC[8].icell.Ien VPWR 0.18883f
C687 XThR.XTB5.A XThR.XTBN.A 0.06303f
C688 XThC.Tn[13] XA.XIR[15].XIC[13].icell.Ien 0.04292f
C689 XA.XIR[14].XIC[4].icell.Ien Iout 0.06801f
C690 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.PDM 0.02104f
C691 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PDM 0.04035f
C692 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PDM 0.02601f
C693 XA.XIR[13].XIC[6].icell.Ien Iout 0.06801f
C694 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.PDM 0.02104f
C695 XThC.Tn[6] XA.XIR[2].XIC[6].icell.Ien 0.04605f
C696 XThC.Tn[8] XThR.Tn[11] 0.40738f
C697 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR 0.39005f
C698 XA.XIR[15].XIC[0].icell.Ien Vbias 0.15953f
C699 XA.XIR[11].XIC[9].icell.Ien Iout 0.06801f
C700 XThR.XTBN.Y a_n1049_6699# 0.07601f
C701 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PDM 0.04035f
C702 XThC.Tn[7] XThR.Tn[7] 0.40738f
C703 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.PDM 0.02104f
C704 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.PDM 0.02104f
C705 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PDM 0.04035f
C706 XThC.XTB5.Y XThC.Tn[9] 0.01732f
C707 XA.XIR[10].XIC[3].icell.PDM Vbias 0.03928f
C708 XThC.Tn[4] Vbias 0.84011f
C709 XThC.XTB6.Y XThC.Tn[13] 0.32317f
C710 XThR.XTBN.A data[5] 0.0148f
C711 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PDM 0.04035f
C712 XThC.Tn[4] XA.XIR[14].XIC[4].icell.Ien 0.04604f
C713 XThC.Tn[11] XThR.Tn[1] 0.40744f
C714 XA.XIR[2].XIC[13].icell.Ien Iout 0.06801f
C715 XA.XIR[15].XIC[5].icell.Ien Vbias 0.15966f
C716 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.PDM 0.02104f
C717 XThC.XTB6.A data[1] 0.37233f
C718 XThR.Tn[8] XA.XIR[8].XIC[14].icell.Ien 0.144f
C719 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.Ien 0.04854f
C720 XThR.XTB4.Y a_n1049_6699# 0.23756f
C721 XA.XIR[10].XIC_dummy_left.icell.Iout XA.XIR[11].XIC_dummy_left.icell.Iout 0.03665f
C722 XThR.XTB6.A XThR.XTB3.Y 0.03869f
C723 XThR.XTB2.Y XThR.XTB7.A 0.2319f
C724 XA.XIR[11].XIC[3].icell.PDM VPWR 0.01171f
C725 XA.XIR[1].XIC_15.icell.Ien Iout 0.0694f
C726 XA.XIR[4].XIC[8].icell.Ien Vbias 0.19161f
C727 XThC.Tn[11] XThR.Tn[12] 0.40738f
C728 XThC.Tn[1] XA.XIR[3].XIC[1].icell.Ien 0.04604f
C729 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.Ien 0.04854f
C730 XA.XIR[10].XIC[7].icell.PDM VPWR 0.01171f
C731 XThR.XTB7.B XThR.Tn[8] 0.05091f
C732 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.PDM 0.02104f
C733 XThC.XTBN.Y XThC.Tn[9] 0.39932f
C734 XA.XIR[8].XIC[2].icell.Ien Vbias 0.19161f
C735 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PDM 0.02601f
C736 XThC.Tn[6] XThR.Tn[3] 0.40738f
C737 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.Ien 0.04854f
C738 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR 0.08547f
C739 XThR.Tn[5] XA.XIR[5].XIC[13].icell.Ien 0.14211f
C740 XA.XIR[0].XIC[11].icell.PDM Vbias 0.03945f
C741 XA.XIR[5].XIC[7].icell.Ien VPWR 0.18829f
C742 XThR.XTB7.A a_n1049_5611# 0.01824f
C743 XA.XIR[5].XIC[3].icell.Ien Iout 0.06801f
C744 XThC.Tn[0] XThR.Tn[0] 0.41303f
C745 XA.XIR[9].XIC[11].icell.Ien Vbias 0.19161f
C746 XThC.Tn[10] XThR.Tn[10] 0.40738f
C747 XThC.Tn[2] XThR.Tn[5] 0.40738f
C748 XA.XIR[12].XIC[14].icell.PDM Vbias 0.03928f
C749 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PDM 0.02601f
C750 XA.XIR[0].XIC[4].icell.Ien Vbias 0.19213f
C751 XA.XIR[1].XIC_dummy_right.icell.Iout Iout 0.01732f
C752 XThC.Tn[9] XThC.Tn[10] 0.0671f
C753 XThR.Tn[13] a_n997_1579# 0.19413f
C754 XA.XIR[15].XIC_15.icell.PDM Vbias 0.03927f
C755 XA.XIR[12].XIC[2].icell.Ien VPWR 0.18829f
C756 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PDM 0.04035f
C757 XA.XIR[0].XIC_15.icell.PDM VPWR 0.07389f
C758 XThC.XTB7.Y VPWR 1.07721f
C759 XA.XIR[7].XIC[7].icell.Ien Vbias 0.19161f
C760 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.PDM 0.02104f
C761 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.PDM 0.02104f
C762 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.PDM 0.02104f
C763 XThR.Tn[4] XA.XIR[4].XIC[3].icell.Ien 0.14211f
C764 XThC.XTBN.A XThC.XTB6.Y 0.06405f
C765 XThR.XTBN.A XThR.Tn[9] 0.12398f
C766 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.PDM 0.02104f
C767 XThR.Tn[6] Iout 1.12758f
C768 XA.XIR[11].XIC[14].icell.Ien Iout 0.06801f
C769 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.Ien 0.04854f
C770 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR 0.01604f
C771 XA.XIR[6].XIC_15.icell.Ien Iout 0.0694f
C772 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.02602f
C773 XThR.XTB6.A VPWR 0.68638f
C774 XThC.Tn[8] XThR.Tn[14] 0.40738f
C775 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.PDM 0.02104f
C776 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PDM 0.04035f
C777 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.Ien 0.04854f
C778 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Iout 0.01728f
C779 a_6243_9615# Vbias 0.01011f
C780 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR 0.39002f
C781 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PDM 0.02601f
C782 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.Ien 0.04854f
C783 XA.XIR[6].XIC[2].icell.PDM Vbias 0.03928f
C784 XA.XIR[14].XIC[9].icell.Ien Iout 0.06801f
C785 XThC.Tn[9] XA.XIR[15].XIC[9].icell.Ien 0.04292f
C786 XThR.XTB1.Y a_n1049_8581# 0.21263f
C787 XA.XIR[5].XIC[9].icell.PDM Vbias 0.03928f
C788 XThR.Tn[3] XA.XIR[3].XIC[6].icell.Ien 0.14211f
C789 XThC.Tn[5] XA.XIR[0].XIC[5].icell.Ien 0.04659f
C790 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.PDM 0.02104f
C791 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.Ien 0.04854f
C792 XThR.Tn[0] VPWR 8.08835f
C793 XA.XIR[13].XIC[3].icell.PDM Vbias 0.03928f
C794 XThC.XTB4.Y XThC.XTBN.A 0.03415f
C795 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PDM 0.04035f
C796 XA.XIR[12].XIC[8].icell.PDM Vbias 0.03928f
C797 XThR.XTB7.B XThR.XTB2.Y 0.22599f
C798 XThR.XTB7.B a_n997_3755# 0.01174f
C799 XA.XIR[6].XIC_dummy_right.icell.Iout Iout 0.01732f
C800 XThC.Tn[4] XThR.Tn[6] 0.40738f
C801 XA.XIR[5].XIC_dummy_right.icell.Iout XA.XIR[6].XIC_dummy_right.icell.Iout 0.04047f
C802 XThR.XTBN.Y XThR.Tn[8] 0.4783f
C803 XA.XIR[6].XIC[6].icell.PDM VPWR 0.01171f
C804 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.Ien 0.04854f
C805 XA.XIR[5].XIC[13].icell.PDM VPWR 0.01171f
C806 XA.XIR[14].XIC[3].icell.PDM VPWR 0.01171f
C807 XThC.Tn[7] XA.XIR[4].XIC[7].icell.Ien 0.04604f
C808 XThC.Tn[6] XThR.Tn[11] 0.40738f
C809 XA.XIR[3].XIC[4].icell.Ien Vbias 0.19161f
C810 XA.XIR[10].XIC[13].icell.Ien Vbias 0.19161f
C811 XA.XIR[13].XIC[7].icell.PDM VPWR 0.01171f
C812 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.PDM 0.02104f
C813 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.PDM 0.02104f
C814 XThR.Tn[4] Iout 1.12761f
C815 XThC.XTB3.Y XThC.XTB6.Y 0.04428f
C816 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.Ien 0.04854f
C817 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.Ien 0.04854f
C818 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PDM 0.02601f
C819 XA.XIR[9].XIC[3].icell.Ien VPWR 0.18829f
C820 XA.XIR[3].XIC[4].icell.PDM Vbias 0.03928f
C821 XA.XIR[8].XIC[6].icell.PDM Vbias 0.03928f
C822 XA.XIR[12].XIC[13].icell.PDM Vbias 0.03928f
C823 XA.XIR[4].XIC[13].icell.Ien Vbias 0.19161f
C824 XThR.XTB4.Y XThR.Tn[8] 0.01306f
C825 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.Ien 0.04854f
C826 XThC.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.04606f
C827 XA.XIR[11].XIC[12].icell.Ien Iout 0.06801f
C828 XThC.Tn[10] XThR.Tn[13] 0.40738f
C829 XA.XIR[2].XIC[10].icell.PDM Vbias 0.03928f
C830 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.02601f
C831 XA.XIR[8].XIC[7].icell.Ien Vbias 0.19161f
C832 XThC.Tn[0] XA.XIR[4].XIC[0].icell.Ien 0.04604f
C833 XThC.Tn[0] XThR.Tn[1] 0.40748f
C834 XA.XIR[15].XIC[14].icell.PDM Vbias 0.03928f
C835 XA.XIR[1].XIC[0].icell.PDM VPWR 0.01171f
C836 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PDM 0.02602f
C837 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PDM 0.04035f
C838 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.02601f
C839 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.PDM 0.02104f
C840 XThR.XTB6.Y XThR.Tn[9] 0.0246f
C841 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.Ien 0.04854f
C842 XThR.XTB7.A XThR.Tn[3] 0.0306f
C843 XThC.Tn[13] Iout 0.22423f
C844 XThC.Tn[13] XThR.Tn[9] 0.40739f
C845 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.PDM 0.02104f
C846 XThC.Tn[0] XThR.Tn[12] 0.40738f
C847 XThC.Tn[9] XThR.Tn[8] 0.40738f
C848 XA.XIR[4].XIC[0].icell.PDM VPWR 0.01171f
C849 XA.XIR[5].XIC[12].icell.Ien VPWR 0.18829f
C850 XThC.XTB6.A VPWR 0.68179f
C851 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.PDM 0.02104f
C852 XA.XIR[5].XIC[8].icell.Ien Iout 0.06801f
C853 XThC.XTB7.B XThC.XTB7.Y 0.33493f
C854 XA.XIR[8].XIC[10].icell.PDM VPWR 0.01171f
C855 XA.XIR[3].XIC[8].icell.PDM VPWR 0.01171f
C856 XA.XIR[4].XIC_15.icell.PUM VPWR 0.01655f
C857 XA.XIR[10].XIC_dummy_left.icell.Iout Iout 0.03553f
C858 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Iout 0.01779f
C859 XThR.XTB7.A XThR.XTB7.Y 0.37429f
C860 XA.XIR[2].XIC[14].icell.PDM VPWR 0.0118f
C861 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.PDM 0.02104f
C862 XThR.XTB7.A data[4] 0.8689f
C863 XThC.XTBN.A a_7875_9569# 0.01939f
C864 XA.XIR[0].XIC[9].icell.Ien Vbias 0.19213f
C865 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PDM 0.04035f
C866 XThC.XTBN.Y XThC.Tn[7] 0.85979f
C867 XThC.Tn[4] XThR.Tn[4] 0.40738f
C868 XThC.XTB3.Y XThC.XTB4.Y 2.13136f
C869 XThC.XTB2.Y XThC.XTBN.A 0.04716f
C870 XA.XIR[12].XIC[7].icell.Ien VPWR 0.18829f
C871 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.PDM 0.02104f
C872 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR 0.08209f
C873 XA.XIR[7].XIC_dummy_right.icell.Iout XA.XIR[8].XIC_dummy_right.icell.Iout 0.04047f
C874 XA.XIR[12].XIC[3].icell.Ien Iout 0.06801f
C875 XThC.Tn[5] XA.XIR[3].XIC[5].icell.Ien 0.04604f
C876 XA.XIR[7].XIC[12].icell.Ien Vbias 0.19161f
C877 XA.XIR[14].XIC[14].icell.Ien Iout 0.06801f
C878 XThC.Tn[12] XA.XIR[2].XIC[12].icell.Ien 0.04605f
C879 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR 0.01669f
C880 XThR.Tn[4] XA.XIR[4].XIC[8].icell.Ien 0.14211f
C881 XThR.Tn[11] XA.XIR[11].XIC[13].icell.Ien 0.14211f
C882 XA.XIR[10].XIC[11].icell.Ien Vbias 0.19161f
C883 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.PDM 0.02104f
C884 XA.XIR[3].XIC[1].icell.Ien Vbias 0.19161f
C885 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PDM 0.04035f
C886 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR 0.38995f
C887 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PDM 0.04035f
C888 XThC.XTB1.Y XThC.XTB6.Y 0.05752f
C889 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.PDM 0.02104f
C890 XThR.XTBN.Y a_n997_3755# 0.229f
C891 XThR.XTBN.Y XThR.XTB2.Y 0.2075f
C892 XA.XIR[1].XIC[0].icell.Ien VPWR 0.18829f
C893 XThR.Tn[2] XA.XIR[2].XIC[1].icell.Ien 0.14211f
C894 XA.XIR[7].XIC[10].icell.PDM Vbias 0.03928f
C895 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.Ien 0.04854f
C896 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.Ien 0.04854f
C897 XA.XIR[11].XIC[10].icell.Ien Iout 0.06801f
C898 XThR.Tn[1] VPWR 8.09331f
C899 XA.XIR[4].XIC[0].icell.Ien VPWR 0.18829f
C900 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PDM 0.02601f
C901 XA.XIR[15].XIC[8].icell.PDM Vbias 0.03928f
C902 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.Ien 0.04854f
C903 XThR.Tn[12] XA.XIR[12].XIC[6].icell.Ien 0.14211f
C904 XThC.XTBN.Y a_3773_9615# 0.08456f
C905 XThR.Tn[3] XA.XIR[3].XIC[11].icell.Ien 0.14211f
C906 XThR.Tn[12] VPWR 8.99609f
C907 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.PDM 0.02104f
C908 XA.XIR[13].XIC_dummy_left.icell.Iout XA.XIR[14].XIC_dummy_left.icell.Iout 0.03665f
C909 XThR.XTBN.Y a_n1049_5611# 0.0768f
C910 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.Ien 0.04854f
C911 XA.XIR[9].XIC[6].icell.PDM Vbias 0.03928f
C912 XThR.XTB2.Y XThR.XTB4.Y 0.04006f
C913 XThC.Tn[6] XThR.Tn[14] 0.40738f
C914 XA.XIR[13].XIC[13].icell.Ien Vbias 0.19161f
C915 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.Ien 0.04854f
C916 XA.XIR[15].XIC[2].icell.Ien VPWR 0.31713f
C917 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.PDM 0.02104f
C918 XA.XIR[7].XIC[14].icell.PDM VPWR 0.0118f
C919 XA.XIR[11].XIC[0].icell.Ien Iout 0.06795f
C920 XThR.Tn[2] XA.XIR[2].XIC[6].icell.Ien 0.14211f
C921 XA.XIR[12].XIC[12].icell.PDM Vbias 0.03928f
C922 XThC.Tn[3] XA.XIR[10].XIC[3].icell.Ien 0.04604f
C923 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.PDM 0.02104f
C924 XA.XIR[4].XIC[5].icell.Ien VPWR 0.18829f
C925 XThC.XTB2.Y XThC.XTB3.Y 2.04808f
C926 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.Ien 0.04854f
C927 XThC.XTB1.Y XThC.XTB4.Y 0.05121f
C928 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.PDM 0.02104f
C929 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PDM 0.02601f
C930 XA.XIR[15].XIC[13].icell.PDM Vbias 0.03928f
C931 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR 0.08221f
C932 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.PDM 0.02104f
C933 XA.XIR[3].XIC[9].icell.Ien Vbias 0.19161f
C934 XA.XIR[14].XIC[12].icell.Ien Iout 0.06801f
C935 XA.XIR[1].XIC[11].icell.PDM Vbias 0.03928f
C936 XA.XIR[9].XIC[10].icell.PDM VPWR 0.01171f
C937 XThC.Tn[8] VPWR 4.5473f
C938 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PDM 0.02602f
C939 XThC.Tn[6] XA.XIR[5].XIC[6].icell.Ien 0.04604f
C940 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR 0.08221f
C941 XA.XIR[0].XIC[2].icell.PDM VPWR 0.01132f
C942 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PDM 0.02601f
C943 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.Ien 0.04854f
C944 XA.XIR[4].XIC[11].icell.PDM Vbias 0.03928f
C945 XA.XIR[2].XIC[2].icell.Ien Vbias 0.19161f
C946 XThR.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.14211f
C947 XA.XIR[9].XIC[8].icell.Ien VPWR 0.18829f
C948 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.Ien 0.04854f
C949 XA.XIR[1].XIC[4].icell.Ien Vbias 0.19173f
C950 XThR.XTB7.B data[4] 0.01382f
C951 XThR.XTB7.B XThR.XTB7.Y 0.33493f
C952 XThR.Tn[9] XA.XIR[9].XIC[4].icell.Ien 0.14211f
C953 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.Ien 0.04854f
C954 XA.XIR[9].XIC[4].icell.Ien Iout 0.06801f
C955 XThC.XTB6.A XThC.XTB7.B 1.47641f
C956 XThC.Tn[2] XA.XIR[7].XIC[2].icell.Ien 0.04604f
C957 XThR.XTB5.Y a_n1319_6405# 0.01188f
C958 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.PDM 0.02104f
C959 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PDM 0.04035f
C960 XA.XIR[8].XIC[12].icell.Ien Vbias 0.19161f
C961 a_n1049_5317# VPWR 0.72036f
C962 XA.XIR[13].XIC_dummy_left.icell.Iout Iout 0.03553f
C963 XA.XIR[1].XIC_15.icell.PDM VPWR 0.07527f
C964 XA.XIR[4].XIC_15.icell.PDM VPWR 0.07527f
C965 XA.XIR[7].XIC[4].icell.Ien VPWR 0.18829f
C966 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.PDM 0.02104f
C967 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.Ien 0.04854f
C968 XThR.Tn[2] XThR.Tn[3] 0.15335f
C969 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR 0.08209f
C970 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.PDM 0.02104f
C971 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout 0.06446f
C972 XA.XIR[5].XIC[13].icell.Ien Iout 0.06801f
C973 XThR.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.14251f
C974 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PDM 0.04056f
C975 XA.XIR[0].XIC[14].icell.Ien Vbias 0.19213f
C976 XThC.Tn[2] Iout 0.22439f
C977 XThC.Tn[2] XThR.Tn[9] 0.40738f
C978 XA.XIR[13].XIC[11].icell.Ien Vbias 0.19161f
C979 XThR.XTBN.Y a_n997_715# 0.21503f
C980 XA.XIR[11].XIC_15.icell.Ien Iout 0.0694f
C981 XThC.Tn[4] XA.XIR[9].XIC[4].icell.Ien 0.04604f
C982 XThR.Tn[7] XA.XIR[7].XIC[1].icell.Ien 0.14211f
C983 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.Ien 0.04854f
C984 VPWR data[7] 0.212f
C985 XA.XIR[12].XIC[8].icell.Ien Iout 0.06801f
C986 XThC.Tn[7] XThR.Tn[8] 0.40738f
C987 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.PDM 0.02104f
C988 XThC.XTB1.Y XThC.XTB2.Y 2.14864f
C989 XThC.Tn[11] XA.XIR[0].XIC[11].icell.Ien 0.04662f
C990 XThR.Tn[4] XA.XIR[4].XIC[13].icell.Ien 0.14211f
C991 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PDM 0.04035f
C992 XA.XIR[11].XIC[1].icell.PDM Vbias 0.03928f
C993 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR 0.01499f
C994 XThR.Tn[0] XA.XIR[0].XIC[5].icell.Ien 0.14211f
C995 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.Ien 0.04854f
C996 XThR.Tn[10] XA.XIR[10].XIC[4].icell.Ien 0.14211f
C997 XThR.XTB7.B a_n997_2667# 0.02071f
C998 XThC.Tn[5] XA.XIR[1].XIC[5].icell.Ien 0.04606f
C999 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PDM 0.04035f
C1000 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PDM 0.02601f
C1001 XA.XIR[14].XIC[10].icell.Ien Iout 0.06801f
C1002 XThC.Tn[13] XA.XIR[10].XIC[13].icell.Ien 0.04604f
C1003 XA.XIR[10].XIC[5].icell.PDM Vbias 0.03928f
C1004 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.PDM 0.02104f
C1005 XA.XIR[5].XIC[0].icell.PDM VPWR 0.01171f
C1006 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PDM 0.04035f
C1007 XThC.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.04604f
C1008 XThR.Tn[7] XA.XIR[7].XIC[6].icell.Ien 0.14211f
C1009 XA.XIR[6].XIC[4].icell.Ien Vbias 0.19161f
C1010 a_n1049_6405# VPWR 0.72095f
C1011 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.Ien 0.04854f
C1012 XA.XIR[8].XIC_dummy_left.icell.Ien XThR.Tn[8] 0.0125f
C1013 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.Ien 0.04854f
C1014 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PDM 0.02601f
C1015 XThC.Tn[13] XA.XIR[4].XIC[13].icell.Ien 0.04604f
C1016 XA.XIR[11].XIC_dummy_right.icell.Iout Iout 0.01732f
C1017 XA.XIR[12].XIC[11].icell.PDM Vbias 0.03928f
C1018 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.PDM 0.02104f
C1019 XA.XIR[11].XIC[5].icell.PDM VPWR 0.01171f
C1020 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.Ien 0.04854f
C1021 XA.XIR[4].XIC[1].icell.Ien Iout 0.06801f
C1022 XA.XIR[10].XIC[9].icell.PDM VPWR 0.01171f
C1023 XA.XIR[15].XIC[12].icell.PDM Vbias 0.03928f
C1024 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.Ien 0.04854f
C1025 XThC.Tn[3] XA.XIR[13].XIC[3].icell.Ien 0.04604f
C1026 XThC.Tn[1] XA.XIR[12].XIC[1].icell.Ien 0.04604f
C1027 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.PDM 0.02104f
C1028 XThR.XTBN.Y XThR.Tn[3] 0.62501f
C1029 XA.XIR[11].XIC_dummy_left.icell.Ien XThR.Tn[11] 0.01244f
C1030 a_n1049_8581# XThR.Tn[0] 0.2685f
C1031 XThR.XTB7.B XThR.Tn[11] 0.03888f
C1032 XThC.Tn[10] XThR.Tn[7] 0.40738f
C1033 XA.XIR[0].XIC[13].icell.PDM Vbias 0.03945f
C1034 XA.XIR[11].XIC[3].icell.Ien Vbias 0.19161f
C1035 XA.XIR[15].XIC[7].icell.Ien VPWR 0.31713f
C1036 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.Ien 0.04854f
C1037 XThC.XTB7.B XThC.Tn[8] 0.05151f
C1038 XThC.Tn[2] XA.XIR[8].XIC[2].icell.Ien 0.04604f
C1039 XThR.Tn[2] XA.XIR[2].XIC[11].icell.Ien 0.14211f
C1040 XThC.Tn[0] XA.XIR[2].XIC[0].icell.Ien 0.04605f
C1041 XThR.XTBN.Y XThR.XTB7.Y 0.50018f
C1042 XA.XIR[15].XIC[3].icell.Ien Iout 0.07192f
C1043 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR 0.38902f
C1044 XA.XIR[10].XIC[5].icell.Ien Vbias 0.19161f
C1045 XThC.XTB7.Y XThC.Tn[12] 0.07091f
C1046 XA.XIR[4].XIC[10].icell.Ien VPWR 0.18829f
C1047 XA.XIR[0].XIC[1].icell.Ien VPWR 0.18776f
C1048 XA.XIR[4].XIC[6].icell.Ien Iout 0.06801f
C1049 XA.XIR[2].XIC[1].icell.PDM VPWR 0.01171f
C1050 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.PDM 0.02104f
C1051 XA.XIR[8].XIC[4].icell.Ien VPWR 0.18829f
C1052 XThR.XTB4.Y XThR.Tn[3] 0.1895f
C1053 XA.XIR[3].XIC[14].icell.Ien Vbias 0.19161f
C1054 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.Ien 0.04854f
C1055 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.PDM 0.02104f
C1056 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PDM 0.04035f
C1057 XA.XIR[2].XIC[7].icell.Ien Vbias 0.19161f
C1058 XThC.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.04604f
C1059 XA.XIR[7].XIC[0].icell.Ien Iout 0.06795f
C1060 XA.XIR[9].XIC[13].icell.Ien VPWR 0.18829f
C1061 XThR.XTB4.Y XThR.XTB7.Y 0.03475f
C1062 XA.XIR[1].XIC[9].icell.Ien Vbias 0.19173f
C1063 XThC.Tn[11] XA.XIR[3].XIC[11].icell.Ien 0.04604f
C1064 XA.XIR[9].XIC[9].icell.Ien Iout 0.06801f
C1065 XThR.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.14211f
C1066 XA.XIR[0].XIC[6].icell.Ien VPWR 0.1878f
C1067 XThC.Tn[9] XThR.Tn[3] 0.40738f
C1068 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.Ien 0.04854f
C1069 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1070 XThC.Tn[6] XA.XIR[12].XIC[6].icell.Ien 0.04604f
C1071 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1072 XThR.XTB7.Y XThR.Tn[10] 0.07406f
C1073 XA.XIR[0].XIC[2].icell.Ien Iout 0.0675f
C1074 XThC.Tn[6] VPWR 3.63495f
C1075 XThR.Tn[5] XA.XIR[5].XIC[0].icell.Ien 0.1423f
C1076 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.Ien 0.04854f
C1077 XA.XIR[7].XIC[9].icell.Ien VPWR 0.18829f
C1078 XThR.Tn[14] XA.XIR[14].XIC[13].icell.Ien 0.14211f
C1079 XThC.Tn[12] XThR.Tn[0] 0.40763f
C1080 XA.XIR[7].XIC[5].icell.Ien Iout 0.06801f
C1081 XA.XIR[14].XIC_15.icell.Ien Iout 0.0694f
C1082 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PDM 0.04035f
C1083 XThC.Tn[14] XThR.Tn[5] 0.40742f
C1084 XThR.XTBN.Y a_n997_2667# 0.22784f
C1085 XA.XIR[9].XIC_dummy_left.icell.Iout XA.XIR[10].XIC_dummy_left.icell.Iout 0.03665f
C1086 XA.XIR[6].XIC[4].icell.PDM Vbias 0.03928f
C1087 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.PDM 0.02104f
C1088 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1089 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.PDM 0.02104f
C1090 XThR.Tn[8] a_n997_3979# 0.1927f
C1091 XA.XIR[14].XIC[1].icell.PDM Vbias 0.03928f
C1092 XA.XIR[5].XIC[11].icell.PDM Vbias 0.03928f
C1093 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.Ien 0.04854f
C1094 XA.XIR[2].XIC[0].icell.Ien VPWR 0.18829f
C1095 XThC.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.04604f
C1096 XA.XIR[13].XIC[5].icell.PDM Vbias 0.03928f
C1097 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PDM 0.02601f
C1098 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PDM 0.04035f
C1099 XThR.Tn[11] XA.XIR[11].XIC[5].icell.Ien 0.14211f
C1100 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PDM 0.02602f
C1101 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Ien 0.01557f
C1102 XA.XIR[12].XIC[10].icell.PDM Vbias 0.03928f
C1103 XA.XIR[10].XIC[1].icell.Ien VPWR 0.18829f
C1104 XA.XIR[7].XIC[1].icell.PDM VPWR 0.01171f
C1105 XThC.Tn[11] XA.XIR[14].XIC[11].icell.Ien 0.04604f
C1106 XThR.XTB4.Y a_n997_2667# 0.07199f
C1107 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PDM 0.02601f
C1108 XA.XIR[6].XIC[8].icell.PDM VPWR 0.01171f
C1109 XThR.Tn[0] XA.XIR[0].XIC[10].icell.Ien 0.14211f
C1110 XThR.Tn[10] XA.XIR[10].XIC[9].icell.Ien 0.14211f
C1111 XA.XIR[14].XIC_dummy_right.icell.Iout Iout 0.01732f
C1112 XA.XIR[15].XIC[11].icell.PDM Vbias 0.03928f
C1113 XA.XIR[14].XIC[5].icell.PDM VPWR 0.01171f
C1114 XThR.Tn[6] XA.XIR[6].XIC[4].icell.Ien 0.14211f
C1115 XA.XIR[5].XIC_15.icell.PDM VPWR 0.07527f
C1116 XThC.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.04604f
C1117 XThR.XTBN.Y XThR.Tn[11] 0.52268f
C1118 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.Ien 0.04854f
C1119 XA.XIR[13].XIC[9].icell.PDM VPWR 0.01171f
C1120 XThC.Tn[11] XThR.Tn[2] 0.40741f
C1121 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.Ien 0.04854f
C1122 XA.XIR[6].XIC[9].icell.Ien Vbias 0.19161f
C1123 XThR.Tn[7] XA.XIR[7].XIC[11].icell.Ien 0.14211f
C1124 XThC.XTB7.Y a_10915_9569# 0.06874f
C1125 XThR.XTB7.A XThR.XTB3.Y 0.57441f
C1126 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1127 XThC.Tn[12] XA.XIR[5].XIC[12].icell.Ien 0.04604f
C1128 XA.XIR[8].XIC[8].icell.PDM Vbias 0.03928f
C1129 XA.XIR[3].XIC[6].icell.PDM Vbias 0.03928f
C1130 XA.XIR[14].XIC[3].icell.Ien Vbias 0.19161f
C1131 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout 0.06446f
C1132 XA.XIR[11].XIC[13].icell.Ien VPWR 0.18829f
C1133 XThR.Tn[7] XThR.Tn[8] 0.12208f
C1134 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.PDM 0.02104f
C1135 XA.XIR[2].XIC[12].icell.PDM Vbias 0.03928f
C1136 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.Ien 0.04854f
C1137 XA.XIR[13].XIC[5].icell.Ien Vbias 0.19161f
C1138 XA.XIR[3].XIC[6].icell.Ien VPWR 0.18829f
C1139 XThR.XTB4.Y XThR.Tn[11] 0.3042f
C1140 XA.XIR[1].XIC[2].icell.PDM VPWR 0.01171f
C1141 XThR.Tn[14] XA.XIR[14].XIC[11].icell.Ien 0.14211f
C1142 XThC.Tn[8] XA.XIR[7].XIC[8].icell.Ien 0.04604f
C1143 XA.XIR[3].XIC[2].icell.Ien Iout 0.06801f
C1144 XA.XIR[4].XIC[2].icell.PDM VPWR 0.01171f
C1145 XA.XIR[11].XIC[8].icell.Ien Vbias 0.19161f
C1146 XThR.Tn[10] XThR.Tn[11] 0.10691f
C1147 XA.XIR[15].XIC[8].icell.Ien Iout 0.07192f
C1148 XA.XIR[3].XIC[10].icell.PDM VPWR 0.01171f
C1149 XA.XIR[4].XIC_15.icell.Ien VPWR 0.26829f
C1150 XThC.XTB5.Y XThC.XTBN.Y 0.162f
C1151 XA.XIR[8].XIC[12].icell.PDM VPWR 0.01171f
C1152 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout 0.06446f
C1153 XThC.Tn[9] XThR.Tn[11] 0.40738f
C1154 XThC.XTBN.A a_8963_9569# 0.01679f
C1155 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1156 XA.XIR[4].XIC[11].icell.Ien Iout 0.06801f
C1157 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PDM 0.04035f
C1158 XThC.XTBN.A data[0] 0.02545f
C1159 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PDM 0.04035f
C1160 XA.XIR[8].XIC[9].icell.Ien VPWR 0.18829f
C1161 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.Ien 0.04854f
C1162 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PDM 0.02601f
C1163 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.Ien 0.04854f
C1164 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.PDM 0.02104f
C1165 XA.XIR[8].XIC[5].icell.Ien Iout 0.06801f
C1166 XThR.XTB7.Y XThR.Tn[13] 0.10781f
C1167 XThC.XTB7.B XThC.Tn[6] 0.04318f
C1168 XA.XIR[2].XIC[12].icell.Ien Vbias 0.19161f
C1169 XThC.XTB5.Y XThC.Tn[10] 0.01755f
C1170 XA.XIR[1].XIC[14].icell.Ien Vbias 0.19173f
C1171 XThC.Tn[5] Vbias 0.82298f
C1172 XThC.Tn[10] XA.XIR[9].XIC[10].icell.Ien 0.04604f
C1173 XA.XIR[9].XIC[14].icell.Ien Iout 0.06801f
C1174 XThR.Tn[9] XA.XIR[9].XIC[14].icell.Ien 0.144f
C1175 XA.XIR[0].XIC[11].icell.Ien VPWR 0.18882f
C1176 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.Ien 0.04854f
C1177 XA.XIR[4].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1178 XThR.Tn[12] XA.XIR[12].XIC_dummy_left.icell.Iout 0.03385f
C1179 XThC.Tn[12] XThR.Tn[1] 0.40744f
C1180 XA.XIR[0].XIC[7].icell.Ien Iout 0.0675f
C1181 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PDM 0.04056f
C1182 XA.XIR[12].XIC[1].icell.Ien Vbias 0.19161f
C1183 XA.XIR[6].XIC_dummy_left.icell.Iout XA.XIR[7].XIC_dummy_left.icell.Iout 0.03665f
C1184 XThC.Tn[11] XA.XIR[1].XIC[11].icell.Ien 0.04606f
C1185 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PDM 0.0404f
C1186 XThR.XTB5.Y XThR.XTBN.A 0.10854f
C1187 XThC.Tn[12] XThR.Tn[12] 0.40738f
C1188 XA.XIR[7].XIC[14].icell.Ien VPWR 0.18835f
C1189 XThR.XTB7.A VPWR 0.88595f
C1190 XThR.Tn[13] XA.XIR[13].XIC[4].icell.Ien 0.14211f
C1191 XThR.Tn[10] XA.XIR[10].XIC[14].icell.Ien 0.144f
C1192 XA.XIR[7].XIC[10].icell.Ien Iout 0.06801f
C1193 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PDM 0.02602f
C1194 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1195 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Iout 0.03842f
C1196 XA.XIR[7].XIC[12].icell.PDM Vbias 0.03928f
C1197 XA.XIR[11].XIC[11].icell.Ien VPWR 0.18829f
C1198 XA.XIR[5].XIC[2].icell.Ien Vbias 0.19161f
C1199 XThC.XTBN.Y XThC.Tn[10] 0.4511f
C1200 XThC.Tn[7] XThR.Tn[3] 0.40738f
C1201 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PDM 0.02601f
C1202 XA.XIR[15].XIC[10].icell.PDM Vbias 0.03928f
C1203 XA.XIR[13].XIC[1].icell.Ien VPWR 0.18829f
C1204 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.PDM 0.02104f
C1205 XThC.XTBN.Y a_4861_9615# 0.07601f
C1206 XA.XIR[8].XIC[0].icell.Ien Iout 0.06795f
C1207 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PDM 0.0279f
C1208 XThC.Tn[1] XThR.Tn[0] 0.40762f
C1209 XThC.Tn[11] XThR.Tn[10] 0.40738f
C1210 XThC.Tn[3] XThR.Tn[5] 0.40738f
C1211 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.Ien 0.04854f
C1212 XA.XIR[9].XIC[8].icell.PDM Vbias 0.03928f
C1213 a_10051_9569# Vbias 0.0105f
C1214 XThC.XTB5.Y a_5155_10571# 0.01188f
C1215 XThR.XTB7.B XThR.XTB3.Y 0.23315f
C1216 XThC.Tn[9] XA.XIR[13].XIC[9].icell.Ien 0.04604f
C1217 XThR.XTBN.Y XThR.Tn[14] 0.47807f
C1218 XA.XIR[0].XIC[0].icell.PDM Vbias 0.03932f
C1219 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.Ien 0.04854f
C1220 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1221 XThC.XTB3.Y data[0] 0.03253f
C1222 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PDM 0.02601f
C1223 XThR.Tn[0] XA.XIR[0].XIC_15.icell.Ien 0.13564f
C1224 XThC.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.04604f
C1225 XThR.Tn[6] XA.XIR[6].XIC[9].icell.Ien 0.14211f
C1226 XA.XIR[1].XIC[13].icell.PDM Vbias 0.03928f
C1227 XA.XIR[14].XIC[13].icell.Ien VPWR 0.18883f
C1228 XThC.Tn[6] XA.XIR[15].XIC[6].icell.Ien 0.04292f
C1229 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.PDM 0.02104f
C1230 XA.XIR[6].XIC[14].icell.Ien Vbias 0.19161f
C1231 XA.XIR[9].XIC[12].icell.PDM VPWR 0.01171f
C1232 XThR.XTB1.Y XThR.XTBN.A 0.12307f
C1233 XA.XIR[0].XIC[4].icell.PDM VPWR 0.01136f
C1234 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout 0.06446f
C1235 XA.XIR[4].XIC[13].icell.PDM Vbias 0.03928f
C1236 XA.XIR[1].XIC[1].icell.Ien VPWR 0.18829f
C1237 XThR.XTB3.Y XThR.Tn[2] 0.18254f
C1238 XA.XIR[10].XIC[2].icell.Ien VPWR 0.18829f
C1239 XA.XIR[14].XIC[8].icell.Ien Vbias 0.19161f
C1240 XThC.Tn[7] XA.XIR[11].XIC[7].icell.Ien 0.04604f
C1241 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.Ien 0.04854f
C1242 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PDM 0.04035f
C1243 XThC.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.04605f
C1244 XThC.Tn[11] XA.XIR[6].XIC[11].icell.Ien 0.04604f
C1245 XThC.Tn[0] XThR.Tn[2] 0.40744f
C1246 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PDM 0.04035f
C1247 XThR.XTB5.Y XThR.Tn[4] 0.19957f
C1248 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PDM 0.04035f
C1249 XA.XIR[3].XIC[11].icell.Ien VPWR 0.18829f
C1250 XThC.Tn[9] XThR.Tn[14] 0.40738f
C1251 XThR.Tn[10] XA.XIR[10].XIC[12].icell.Ien 0.14211f
C1252 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PDM 0.02601f
C1253 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1254 XA.XIR[3].XIC[7].icell.Ien Iout 0.06801f
C1255 XA.XIR[2].XIC[4].icell.Ien VPWR 0.18829f
C1256 XThR.Tn[1] a_n1049_7787# 0.26879f
C1257 XA.XIR[1].XIC[6].icell.Ien VPWR 0.18829f
C1258 XThR.XTB5.Y XThR.XTB6.Y 2.12831f
C1259 XA.XIR[1].XIC[2].icell.Ien Iout 0.06801f
C1260 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.PDM 0.02104f
C1261 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.Ien 0.04854f
C1262 XA.XIR[8].XIC[14].icell.Ien VPWR 0.18835f
C1263 XA.XIR[8].XIC[10].icell.Ien Iout 0.06801f
C1264 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR 0.38914f
C1265 XThC.Tn[5] XThR.Tn[6] 0.40738f
C1266 XThR.Tn[7] XA.XIR[7].XIC_dummy_left.icell.Iout 0.0402f
C1267 XThR.XTB7.B VPWR 1.67447f
C1268 XThC.XTB1.Y data[0] 0.06453f
C1269 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.PDM 0.02104f
C1270 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PDM 0.0404f
C1271 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.PDM 0.02104f
C1272 XThC.Tn[7] XThR.Tn[11] 0.40738f
C1273 XA.XIR[11].XIC[3].icell.PDM Vbias 0.03928f
C1274 XA.XIR[14].XIC[11].icell.Ien VPWR 0.18883f
C1275 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PDM 0.04035f
C1276 XA.XIR[0].XIC[12].icell.Ien Iout 0.0675f
C1277 XA.XIR[10].XIC[7].icell.PDM Vbias 0.03928f
C1278 XThR.Tn[14] XA.XIR[14].XIC[5].icell.Ien 0.14211f
C1279 XA.XIR[5].XIC[2].icell.PDM VPWR 0.01171f
C1280 XThR.Tn[1] XA.XIR[1].XIC[5].icell.Ien 0.14211f
C1281 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PDM 0.02601f
C1282 XThR.XTBN.Y XThR.XTB3.Y 0.17246f
C1283 XA.XIR[6].XIC[1].icell.Ien VPWR 0.18829f
C1284 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PDM 0.04035f
C1285 XThC.Tn[10] XA.XIR[12].XIC[10].icell.Ien 0.04604f
C1286 XThR.Tn[13] XA.XIR[13].XIC[9].icell.Ien 0.14211f
C1287 XA.XIR[12].XIC[1].icell.PDM VPWR 0.01171f
C1288 XA.XIR[7].XIC_15.icell.Ien Iout 0.0694f
C1289 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.PDM 0.02104f
C1290 XThC.Tn[11] XThR.Tn[13] 0.40738f
C1291 XA.XIR[5].XIC[7].icell.Ien Vbias 0.19161f
C1292 XThR.Tn[2] VPWR 8.04926f
C1293 XA.XIR[5].XIC[0].icell.Ien Iout 0.06795f
C1294 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.PDM 0.02104f
C1295 XThC.Tn[1] XThR.Tn[1] 0.40744f
C1296 XA.XIR[11].XIC[7].icell.PDM VPWR 0.01171f
C1297 XThR.XTB1.Y XThR.XTB6.Y 0.05751f
C1298 XA.XIR[4].XIC_dummy_left.icell.Iout Iout 0.03553f
C1299 XThR.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.14211f
C1300 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.PDM 0.02104f
C1301 XThC.Tn[14] Iout 0.22441f
C1302 XThC.Tn[14] XThR.Tn[9] 0.40742f
C1303 XThC.Tn[1] XThR.Tn[12] 0.40738f
C1304 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PDM 0.02601f
C1305 XThC.Tn[10] XThR.Tn[8] 0.40738f
C1306 XThR.XTB3.Y XThR.XTB4.Y 2.13136f
C1307 XA.XIR[12].XIC[2].icell.Ien Vbias 0.19161f
C1308 XA.XIR[6].XIC[6].icell.Ien VPWR 0.18829f
C1309 XA.XIR[0].XIC_15.icell.PDM Vbias 0.03947f
C1310 XA.XIR[6].XIC[2].icell.Ien Iout 0.06801f
C1311 XThC.XTB7.Y Vbias 0.01962f
C1312 XThC.XTBN.Y a_7651_9569# 0.23021f
C1313 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.PDM 0.02104f
C1314 XThR.XTB3.Y XThR.Tn[10] 0.29462f
C1315 XThC.Tn[5] XThR.Tn[4] 0.40738f
C1316 XA.XIR[7].XIC_dummy_right.icell.Iout Iout 0.01732f
C1317 XA.XIR[0].XIC_dummy_left.icell.Iout VPWR 0.1175f
C1318 XThC.XTB4.Y XThC.Tn[3] 0.1917f
C1319 XThC.Tn[0] XThR.Tn[10] 0.40734f
C1320 XThR.Tn[6] XA.XIR[6].XIC[14].icell.Ien 0.144f
C1321 XA.XIR[2].XIC[3].icell.PDM VPWR 0.01171f
C1322 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14] 0.14211f
C1323 XA.XIR[13].XIC[2].icell.Ien VPWR 0.18829f
C1324 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.Ien 0.04854f
C1325 XThC.Tn[7] XA.XIR[14].XIC[7].icell.Ien 0.04604f
C1326 XThR.Tn[13] XThR.Tn[14] 0.20347f
C1327 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PDM 0.04035f
C1328 XA.XIR[11].XIC[5].icell.Ien VPWR 0.18829f
C1329 XThR.Tn[8] XA.XIR[8].XIC[1].icell.Ien 0.14211f
C1330 XA.XIR[10].XIC[7].icell.Ien VPWR 0.18829f
C1331 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.PDM 0.02104f
C1332 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.PDM 0.02104f
C1333 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1334 XThR.XTB7.Y XThR.Tn[7] 0.0835f
C1335 XA.XIR[10].XIC[3].icell.Ien Iout 0.06801f
C1336 XThC.XTB2.Y a_4067_9615# 0.02133f
C1337 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Iout 0.01728f
C1338 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PDM 0.02601f
C1339 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.PDM 0.02104f
C1340 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PDM 0.04035f
C1341 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.PDM 0.02104f
C1342 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1343 XThR.XTBN.Y VPWR 4.54335f
C1344 XA.XIR[3].XIC[12].icell.Ien Iout 0.06801f
C1345 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PDM 0.0404f
C1346 XA.XIR[2].XIC[9].icell.Ien VPWR 0.18829f
C1347 XThR.Tn[0] Vbias 1.40808f
C1348 XA.XIR[2].XIC[5].icell.Ien Iout 0.06801f
C1349 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.PDM 0.02104f
C1350 XA.XIR[1].XIC[11].icell.Ien VPWR 0.18829f
C1351 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PDM 0.04035f
C1352 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.Ien 0.04854f
C1353 XThR.Tn[8] XA.XIR[8].XIC[6].icell.Ien 0.14211f
C1354 XA.XIR[1].XIC[7].icell.Ien Iout 0.06801f
C1355 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.Ien 0.04854f
C1356 XThC.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.04604f
C1357 XA.XIR[6].XIC[6].icell.PDM Vbias 0.03928f
C1358 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PDM 0.02601f
C1359 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.PDM 0.02104f
C1360 XThC.Tn[7] XThR.Tn[14] 0.40738f
C1361 XA.XIR[14].XIC[3].icell.PDM Vbias 0.03928f
C1362 XThR.Tn[13] XA.XIR[13].XIC[14].icell.Ien 0.144f
C1363 XA.XIR[5].XIC[13].icell.PDM Vbias 0.03928f
C1364 a_10051_9569# XThC.Tn[13] 0.1927f
C1365 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PDM 0.02601f
C1366 XA.XIR[8].XIC_15.icell.Ien Iout 0.0694f
C1367 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.PDM 0.02104f
C1368 XThR.XTB4.Y VPWR 0.92827f
C1369 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.Ien 0.04854f
C1370 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PDM 0.04056f
C1371 XA.XIR[13].XIC[7].icell.PDM Vbias 0.03928f
C1372 XThR.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.14211f
C1373 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PDM 0.04035f
C1374 XThR.Tn[10] XA.XIR[10].XIC_15.icell.Ien 0.13564f
C1375 XA.XIR[7].XIC[3].icell.PDM VPWR 0.01171f
C1376 XThR.Tn[10] VPWR 8.95184f
C1377 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Ien 0.01557f
C1378 XA.XIR[9].XIC[3].icell.Ien Vbias 0.19161f
C1379 XA.XIR[6].XIC[10].icell.PDM VPWR 0.01171f
C1380 XA.XIR[15].XIC[1].icell.PDM VPWR 0.01512f
C1381 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.Ien 0.04854f
C1382 XThC.Tn[9] VPWR 4.54443f
C1383 XThR.XTB5.A a_n1335_4229# 0.01243f
C1384 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PDM 0.02602f
C1385 XThR.Tn[1] XA.XIR[1].XIC[10].icell.Ien 0.14211f
C1386 XA.XIR[14].XIC[7].icell.PDM VPWR 0.01171f
C1387 XA.XIR[1].XIC[0].icell.PDM Vbias 0.03915f
C1388 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PDM 0.02601f
C1389 XA.XIR[8].XIC_dummy_right.icell.Iout Iout 0.01732f
C1390 XA.XIR[4].XIC[0].icell.PDM Vbias 0.03915f
C1391 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.Ien 0.04854f
C1392 XA.XIR[5].XIC[12].icell.Ien Vbias 0.19161f
C1393 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.Ien 0.04854f
C1394 XA.XIR[1].XIC_dummy_left.icell.Iout XA.XIR[2].XIC_dummy_left.icell.Iout 0.03665f
C1395 data[5] data[6] 0.01513f
C1396 XA.XIR[3].XIC[8].icell.PDM Vbias 0.03928f
C1397 XA.XIR[8].XIC[10].icell.PDM Vbias 0.03928f
C1398 XThC.XTB7.A XThC.XTB5.Y 0.11935f
C1399 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.Ien 0.04854f
C1400 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.PDM 0.02104f
C1401 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PDM 0.02601f
C1402 XA.XIR[2].XIC[14].icell.PDM Vbias 0.03928f
C1403 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.Ien 0.04854f
C1404 XThC.Tn[0] XA.XIR[14].XIC[0].icell.Ien 0.04604f
C1405 XA.XIR[1].XIC[4].icell.PDM VPWR 0.01171f
C1406 XThC.Tn[0] XThR.Tn[13] 0.40741f
C1407 XA.XIR[6].XIC[11].icell.Ien VPWR 0.18829f
C1408 XA.XIR[12].XIC[7].icell.Ien Vbias 0.19161f
C1409 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.PDM 0.02104f
C1410 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.Ien 0.04854f
C1411 XThC.Tn[8] XA.XIR[2].XIC[8].icell.Ien 0.04605f
C1412 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.Ien 0.04854f
C1413 XA.XIR[4].XIC[4].icell.PDM VPWR 0.01171f
C1414 XA.XIR[6].XIC[7].icell.Ien Iout 0.06801f
C1415 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PDM 0.04042f
C1416 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.Ien 0.04854f
C1417 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.Ien 0.04854f
C1418 XThC.Tn[3] Iout 0.22443f
C1419 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.PDM 0.02104f
C1420 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout 0.06446f
C1421 XThC.Tn[3] XThR.Tn[9] 0.40738f
C1422 XA.XIR[3].XIC[12].icell.PDM VPWR 0.01171f
C1423 XA.XIR[8].XIC[14].icell.PDM VPWR 0.0118f
C1424 XA.XIR[14].XIC[5].icell.Ien VPWR 0.18883f
C1425 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.Ien 0.04854f
C1426 XThC.Tn[1] XA.XIR[0].XIC[1].icell.Ien 0.04659f
C1427 XThR.Tn[13] XA.XIR[13].XIC[12].icell.Ien 0.14211f
C1428 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.02602f
C1429 XThC.XTB7.A XThC.XTBN.Y 0.59539f
C1430 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PDM 0.04035f
C1431 XA.XIR[13].XIC[7].icell.Ien VPWR 0.18829f
C1432 XThR.XTB6.A XThR.XTBN.A 0.0512f
C1433 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PDM 0.04035f
C1434 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1435 XA.XIR[13].XIC[3].icell.Ien Iout 0.06801f
C1436 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PDM 0.02601f
C1437 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1438 XThR.XTB7.Y a_n997_1579# 0.013f
C1439 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.PDM 0.02104f
C1440 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PDM 0.02601f
C1441 a_n997_1803# VPWR 0.01991f
C1442 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PDM 0.02792f
C1443 XA.XIR[1].XIC[0].icell.Ien Vbias 0.1916f
C1444 XA.XIR[11].XIC[6].icell.Ien Iout 0.06801f
C1445 XThC.Tn[10] XA.XIR[15].XIC[10].icell.Ien 0.04292f
C1446 XA.XIR[9].XIC_dummy_left.icell.Ien XThR.Tn[9] 0.01244f
C1447 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PDM 0.0404f
C1448 XA.XIR[4].XIC[0].icell.Ien Vbias 0.19149f
C1449 XA.XIR[10].XIC[8].icell.Ien Iout 0.06801f
C1450 XThR.Tn[1] Vbias 1.39552f
C1451 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PDM 0.02601f
C1452 XThC.XTB7.A a_4861_9615# 0.02294f
C1453 XThC.Tn[3] XThC.Tn[4] 0.45992f
C1454 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PDM 0.02601f
C1455 XThR.Tn[12] Vbias 1.39531f
C1456 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PDM 0.0404f
C1457 XA.XIR[2].XIC[14].icell.Ien VPWR 0.18835f
C1458 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.PDM 0.02104f
C1459 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.02601f
C1460 XThC.XTB5.A XThC.XTB5.Y 0.0538f
C1461 XA.XIR[2].XIC[10].icell.Ien Iout 0.06801f
C1462 XA.XIR[15].XIC[2].icell.Ien Vbias 0.15966f
C1463 XA.XIR[7].XIC[14].icell.PDM Vbias 0.03928f
C1464 XThR.Tn[8] XA.XIR[8].XIC[11].icell.Ien 0.14211f
C1465 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.Ien 0.04854f
C1466 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.Ien 0.04854f
C1467 XA.XIR[14].XIC[0].icell.Ien VPWR 0.18883f
C1468 XA.XIR[1].XIC[12].icell.Ien Iout 0.06801f
C1469 XA.XIR[4].XIC[5].icell.Ien Vbias 0.19161f
C1470 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.Ien 0.04854f
C1471 XThR.Tn[13] VPWR 9.0331f
C1472 XThC.Tn[11] XThR.Tn[7] 0.40738f
C1473 XThC.XTBN.Y a_5949_9615# 0.07703f
C1474 XThC.Tn[2] XA.XIR[5].XIC[2].icell.Ien 0.04604f
C1475 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.PDM 0.02104f
C1476 XThC.XTB7.B XThC.Tn[9] 0.05542f
C1477 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.PDM 0.02104f
C1478 XThC.XTB7.Y XThC.Tn[13] 0.10846f
C1479 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.PDM 0.02104f
C1480 XThR.Tn[5] XA.XIR[5].XIC[10].icell.Ien 0.14211f
C1481 XThC.Tn[8] Vbias 0.79784f
C1482 XA.XIR[9].XIC[10].icell.PDM Vbias 0.03928f
C1483 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.Ien 0.04854f
C1484 XA.XIR[0].XIC[2].icell.PDM Vbias 0.03945f
C1485 XThR.Tn[13] XA.XIR[13].XIC[10].icell.Ien 0.14211f
C1486 XThC.Tn[1] XA.XIR[10].XIC[1].icell.Ien 0.04604f
C1487 XA.XIR[5].XIC[4].icell.Ien VPWR 0.18829f
C1488 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PDM 0.02601f
C1489 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.PDM 0.02104f
C1490 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PDM 0.02601f
C1491 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.PDM 0.02104f
C1492 XA.XIR[9].XIC[8].icell.Ien Vbias 0.19161f
C1493 XThR.Tn[3] a_n1049_6699# 0.27008f
C1494 XThR.Tn[1] XA.XIR[1].XIC_15.icell.Ien 0.13564f
C1495 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.PDM 0.02104f
C1496 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.02601f
C1497 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.PDM 0.02104f
C1498 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.PDM 0.02104f
C1499 XA.XIR[1].XIC_15.icell.PDM Vbias 0.03927f
C1500 XA.XIR[9].XIC[14].icell.PDM VPWR 0.0118f
C1501 XThR.XTB6.A XThR.XTB6.Y 0.10153f
C1502 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.PDM 0.02104f
C1503 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.Ien 0.04854f
C1504 XA.XIR[0].XIC[6].icell.PDM VPWR 0.01138f
C1505 XThC.Tn[10] XThR.Tn[3] 0.40738f
C1506 XA.XIR[4].XIC_15.icell.PDM Vbias 0.03927f
C1507 XA.XIR[7].XIC[4].icell.Ien Vbias 0.19161f
C1508 XA.XIR[1].XIC_dummy_left.icell.Iout VPWR 0.11048f
C1509 XThC.Tn[7] VPWR 3.9785f
C1510 XA.XIR[12].XIC[13].icell.Ien Iout 0.06801f
C1511 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.Ien 0.04854f
C1512 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PDM 0.04035f
C1513 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PDM 0.0404f
C1514 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PDM 0.04035f
C1515 XThC.Tn[13] XThR.Tn[0] 0.40764f
C1516 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.PDM 0.02104f
C1517 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.PDM 0.02104f
C1518 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1519 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1520 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PDM 0.02601f
C1521 XA.XIR[6].XIC[12].icell.Ien Iout 0.06801f
C1522 XThC.Tn[6] XA.XIR[10].XIC[6].icell.Ien 0.04604f
C1523 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.PDM 0.02104f
C1524 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout 0.06446f
C1525 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PDM 0.02803f
C1526 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Ien 0.01263f
C1527 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.Ien 0.04854f
C1528 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR 0.38999f
C1529 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PDM 0.02601f
C1530 XA.XIR[14].XIC[6].icell.Ien Iout 0.06801f
C1531 XThC.XTBN.A XThC.XTB7.Y 1.11562f
C1532 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.04035f
C1533 XA.XIR[5].XIC[0].icell.PDM Vbias 0.03915f
C1534 XA.XIR[13].XIC[8].icell.Ien Iout 0.06801f
C1535 XThR.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.14211f
C1536 XThC.Tn[9] XA.XIR[4].XIC[9].icell.Ien 0.04604f
C1537 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PDM 0.02601f
C1538 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.Ien 0.04854f
C1539 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.PDM 0.02104f
C1540 XThR.XTBN.A XThR.Tn[12] 0.22096f
C1541 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.PDM 0.02104f
C1542 XThC.Tn[5] XA.XIR[7].XIC[5].icell.Ien 0.04604f
C1543 a_3773_9615# VPWR 0.70508f
C1544 XA.XIR[11].XIC[5].icell.PDM Vbias 0.03928f
C1545 XThC.Tn[12] XThR.Tn[2] 0.40741f
C1546 XThR.XTB2.Y a_n997_3755# 0.06476f
C1547 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.Ien 0.04854f
C1548 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PDM 0.04035f
C1549 XA.XIR[10].XIC[9].icell.PDM Vbias 0.03928f
C1550 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.PDM 0.02104f
C1551 XA.XIR[5].XIC[4].icell.PDM VPWR 0.01171f
C1552 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.PDM 0.02104f
C1553 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout 0.06446f
C1554 XThC.XTB4.Y a_5155_9615# 0.01546f
C1555 XThR.XTBN.Y a_n1049_8581# 0.0607f
C1556 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.PDM 0.02104f
C1557 XThR.Tn[13] XA.XIR[13].XIC_15.icell.Ien 0.13564f
C1558 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PDM 0.04056f
C1559 XA.XIR[6].XIC_dummy_left.icell.Iout VPWR 0.11008f
C1560 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.Ien 0.04854f
C1561 XA.XIR[12].XIC[3].icell.PDM VPWR 0.01171f
C1562 XA.XIR[2].XIC_15.icell.Ien Iout 0.0694f
C1563 XA.XIR[15].XIC[7].icell.Ien Vbias 0.15966f
C1564 XA.XIR[12].XIC[11].icell.Ien Iout 0.06801f
C1565 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.PDM 0.02104f
C1566 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.Ien 0.04854f
C1567 XA.XIR[11].XIC[9].icell.PDM VPWR 0.01171f
C1568 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PDM 0.02601f
C1569 XA.XIR[4].XIC[10].icell.Ien Vbias 0.19161f
C1570 XThC.Tn[1] XA.XIR[13].XIC[1].icell.Ien 0.04604f
C1571 XA.XIR[0].XIC[1].icell.Ien Vbias 0.19213f
C1572 XA.XIR[2].XIC[1].icell.PDM Vbias 0.03928f
C1573 XThC.Tn[8] XThR.Tn[6] 0.40738f
C1574 XThC.Tn[7] XA.XIR[9].XIC[7].icell.Ien 0.04604f
C1575 XA.XIR[8].XIC[4].icell.Ien Vbias 0.19161f
C1576 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PDM 0.04035f
C1577 XThC.Tn[14] XA.XIR[0].XIC[14].icell.Ien 0.04662f
C1578 XThR.Tn[5] XA.XIR[5].XIC_15.icell.Ien 0.13564f
C1579 XThR.XTB3.Y a_n997_2891# 0.07285f
C1580 XThC.Tn[10] XThR.Tn[11] 0.40738f
C1581 XA.XIR[5].XIC[9].icell.Ien VPWR 0.18829f
C1582 XThC.XTBN.Y a_8739_9569# 0.22804f
C1583 XThC.Tn[0] XThR.Tn[7] 0.40736f
C1584 XA.XIR[9].XIC[13].icell.Ien Vbias 0.19161f
C1585 XA.XIR[5].XIC[5].icell.Ien Iout 0.06801f
C1586 XA.XIR[2].XIC_dummy_right.icell.Iout Iout 0.01732f
C1587 XThC.XTB3.Y XThC.XTB7.Y 0.03772f
C1588 XThR.Tn[4] XA.XIR[4].XIC[0].icell.Ien 0.1423f
C1589 XThC.XTB4.Y XThC.XTB6.Y 0.04273f
C1590 XA.XIR[8].XIC[1].icell.PDM VPWR 0.01171f
C1591 XThC.Tn[2] XA.XIR[12].XIC[2].icell.Ien 0.04604f
C1592 a_n1049_5317# XThR.Tn[6] 0.26047f
C1593 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10] 0.14211f
C1594 XThR.Tn[3] XA.XIR[3].XIC[0].icell.Ien 0.14251f
C1595 XA.XIR[2].XIC[5].icell.PDM VPWR 0.01171f
C1596 XA.XIR[0].XIC[6].icell.Ien Vbias 0.19213f
C1597 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout 0.06446f
C1598 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.PDM 0.02104f
C1599 XThC.XTB7.B XThC.Tn[7] 0.07854f
C1600 XThC.XTB5.Y XThC.Tn[11] 0.02112f
C1601 XA.XIR[12].XIC[4].icell.Ien VPWR 0.18829f
C1602 XThC.Tn[6] Vbias 0.81928f
C1603 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout 0.06446f
C1604 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.Ien 0.04854f
C1605 XThR.Tn[5] Iout 1.12761f
C1606 XThR.XTB7.Y XThR.Tn[8] 0.07806f
C1607 a_8739_9569# XThC.Tn[10] 0.21014f
C1608 XThR.Tn[8] data[4] 0.01643f
C1609 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PDM 0.04035f
C1610 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.PDM 0.02104f
C1611 a_n997_3979# VPWR 0.01662f
C1612 XA.XIR[7].XIC[9].icell.Ien Vbias 0.19161f
C1613 XThC.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.04606f
C1614 XA.XIR[9].XIC_15.icell.PUM VPWR 0.01655f
C1615 XThC.Tn[13] XThR.Tn[1] 0.40745f
C1616 XThR.Tn[8] XA.XIR[8].XIC_dummy_left.icell.Iout 0.03962f
C1617 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1618 XThR.XTBN.A data[7] 0.07741f
C1619 XThC.Tn[6] XA.XIR[13].XIC[6].icell.Ien 0.04604f
C1620 XThR.Tn[4] XA.XIR[4].XIC[5].icell.Ien 0.14211f
C1621 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.Ien 0.04854f
C1622 XThR.XTB6.Y XThR.Tn[12] 0.02431f
C1623 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.Ien 0.04854f
C1624 XThC.Tn[13] XThR.Tn[12] 0.40739f
C1625 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PDM 0.04035f
C1626 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PDM 0.04035f
C1627 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.PDM 0.02104f
C1628 XThC.XTB6.A XThC.XTBN.A 0.0513f
C1629 XA.XIR[2].XIC[0].icell.Ien Vbias 0.19149f
C1630 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PDM 0.02602f
C1631 XThC.Tn[5] XA.XIR[8].XIC[5].icell.Ien 0.04604f
C1632 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PDM 0.04035f
C1633 XThC.XTBN.Y XThC.Tn[11] 0.40412f
C1634 XThC.Tn[8] XThR.Tn[4] 0.40738f
C1635 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR 0.38939f
C1636 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PDM 0.02601f
C1637 XA.XIR[7].XIC[1].icell.PDM Vbias 0.03928f
C1638 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.04035f
C1639 XA.XIR[10].XIC[1].icell.Ien Vbias 0.19161f
C1640 XThC.Tn[2] XThR.Tn[0] 0.40765f
C1641 XThC.Tn[12] XThR.Tn[10] 0.40738f
C1642 XA.XIR[6].XIC[8].icell.PDM Vbias 0.03928f
C1643 XThC.Tn[4] XThR.Tn[5] 0.40738f
C1644 XThR.Tn[12] XA.XIR[12].XIC[3].icell.Ien 0.14211f
C1645 XA.XIR[14].XIC[5].icell.PDM Vbias 0.03928f
C1646 XA.XIR[5].XIC_15.icell.PDM Vbias 0.03927f
C1647 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.Ien 0.04854f
C1648 XThR.Tn[3] XA.XIR[3].XIC[8].icell.Ien 0.14211f
C1649 XThC.Tn[10] XThC.Tn[11] 0.07237f
C1650 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PDM 0.02601f
C1651 XThR.Tn[7] VPWR 8.3986f
C1652 XA.XIR[13].XIC[9].icell.PDM Vbias 0.03928f
C1653 a_n997_2891# VPWR 0.01347f
C1654 XThC.Tn[8] XA.XIR[5].XIC[8].icell.Ien 0.04604f
C1655 XThC.XTB2.Y XThC.XTB6.Y 0.04959f
C1656 XThC.XTB1.Y XThC.XTB7.Y 0.05222f
C1657 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PDM 0.04035f
C1658 XThC.Tn[14] XA.XIR[3].XIC[14].icell.Ien 0.04604f
C1659 XA.XIR[7].XIC[5].icell.PDM VPWR 0.01171f
C1660 XThR.Tn[2] XA.XIR[2].XIC[3].icell.Ien 0.14211f
C1661 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout 0.06446f
C1662 XThR.XTB6.Y a_n1049_5317# 0.01199f
C1663 XA.XIR[15].XIC[3].icell.PDM VPWR 0.01512f
C1664 XA.XIR[4].XIC[2].icell.Ien VPWR 0.18829f
C1665 XA.XIR[6].XIC[12].icell.PDM VPWR 0.01171f
C1666 XA.XIR[3].XIC_dummy_right.icell.Iout XA.XIR[4].XIC_dummy_right.icell.Iout 0.04047f
C1667 XA.XIR[11].XIC[13].icell.Ien Vbias 0.19161f
C1668 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.Ien 0.04854f
C1669 XThC.Tn[0] XA.XIR[9].XIC[0].icell.Ien 0.04604f
C1670 XA.XIR[14].XIC[9].icell.PDM VPWR 0.01171f
C1671 XA.XIR[15].XIC[13].icell.Ien Iout 0.07192f
C1672 XThC.Tn[1] XA.XIR[6].XIC[1].icell.Ien 0.04604f
C1673 XA.XIR[3].XIC[6].icell.Ien Vbias 0.19161f
C1674 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.Ien 0.04854f
C1675 XA.XIR[1].XIC[2].icell.PDM Vbias 0.03928f
C1676 XA.XIR[9].XIC[1].icell.PDM VPWR 0.01171f
C1677 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PDM 0.02601f
C1678 XThC.Tn[1] XThR.Tn[2] 0.40741f
C1679 XA.XIR[4].XIC[2].icell.PDM Vbias 0.03928f
C1680 XA.XIR[9].XIC[5].icell.Ien VPWR 0.18829f
C1681 XA.XIR[8].XIC[12].icell.PDM Vbias 0.03928f
C1682 XA.XIR[3].XIC[10].icell.PDM Vbias 0.03928f
C1683 XA.XIR[4].XIC_15.icell.Ien Vbias 0.19195f
C1684 XThR.XTB5.A data[5] 0.11096f
C1685 XThC.Tn[10] XThR.Tn[14] 0.40738f
C1686 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PDM 0.02601f
C1687 XThR.XTBN.Y a_n1049_7787# 0.08456f
C1688 XThC.XTB6.A XThC.XTB3.Y 0.03869f
C1689 XThC.XTB2.Y XThC.XTB4.Y 0.04006f
C1690 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.Ien 0.04854f
C1691 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PDM 0.0404f
C1692 XA.XIR[8].XIC[9].icell.Ien Vbias 0.19161f
C1693 XThR.XTB2.Y XThR.XTB7.Y 0.0437f
C1694 XA.XIR[1].XIC[6].icell.PDM VPWR 0.01171f
C1695 XA.XIR[5].XIC_dummy_left.icell.Iout XA.XIR[6].XIC_dummy_left.icell.Iout 0.03665f
C1696 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PDM 0.02601f
C1697 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11] 0.14211f
C1698 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1699 a_5155_9615# XThC.Tn[4] 0.27224f
C1700 a_n1049_6405# XThR.Tn[4] 0.26564f
C1701 XA.XIR[5].XIC[14].icell.Ien VPWR 0.18835f
C1702 XA.XIR[4].XIC[6].icell.PDM VPWR 0.01171f
C1703 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PDM 0.04035f
C1704 XA.XIR[11].XIC_dummy_left.icell.Iout Iout 0.03553f
C1705 XA.XIR[5].XIC[10].icell.Ien Iout 0.06801f
C1706 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1707 XA.XIR[3].XIC[14].icell.PDM VPWR 0.0118f
C1708 XThC.Tn[6] XThR.Tn[6] 0.40738f
C1709 XThC.XTBN.A XThC.Tn[8] 0.13691f
C1710 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.PDM 0.02104f
C1711 XA.XIR[0].XIC[11].icell.Ien Vbias 0.19213f
C1712 XA.XIR[12].XIC_15.icell.PUM VPWR 0.01655f
C1713 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PDM 0.04035f
C1714 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PDM 0.04035f
C1715 XA.XIR[12].XIC[9].icell.Ien VPWR 0.18829f
C1716 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.Ien 0.04854f
C1717 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1718 XA.XIR[12].XIC[5].icell.Ien Iout 0.06801f
C1719 XA.XIR[7].XIC[14].icell.Ien Vbias 0.19161f
C1720 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PDM 0.02602f
C1721 XA.XIR[9].XIC[0].icell.Ien VPWR 0.18829f
C1722 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Iout 0.01828f
C1723 XA.XIR[11].XIC[11].icell.Ien Vbias 0.19161f
C1724 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PDM 0.04035f
C1725 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PDM 0.02601f
C1726 XThR.Tn[4] XA.XIR[4].XIC[10].icell.Ien 0.14211f
C1727 XA.XIR[15].XIC[11].icell.Ien Iout 0.07192f
C1728 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PDM 0.02601f
C1729 XThR.Tn[0] XA.XIR[0].XIC[2].icell.Ien 0.14211f
C1730 XA.XIR[13].XIC[1].icell.Ien Vbias 0.19161f
C1731 XThC.XTB7.A a_5949_9615# 0.01824f
C1732 XThC.Tn[11] XA.XIR[7].XIC[11].icell.Ien 0.04604f
C1733 XThC.Tn[12] XThR.Tn[13] 0.40738f
C1734 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PDM 0.04035f
C1735 XThC.Tn[2] XThR.Tn[1] 0.40744f
C1736 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.Ien 0.04854f
C1737 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1738 XThR.Tn[7] XA.XIR[7].XIC[3].icell.Ien 0.14211f
C1739 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PDM 0.02601f
C1740 XThC.XTB2.Y a_7875_9569# 0.06476f
C1741 XThC.XTB1.Y XThC.XTB6.A 0.01609f
C1742 XThC.Tn[2] XThR.Tn[12] 0.40738f
C1743 XThC.XTB5.A XThC.XTB7.A 0.07824f
C1744 a_n997_1579# VPWR 0.02417f
C1745 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout 0.06446f
C1746 XThC.Tn[11] XThR.Tn[8] 0.40738f
C1747 XThC.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.04604f
C1748 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.PDM 0.02104f
C1749 XThR.Tn[12] XA.XIR[12].XIC[8].icell.Ien 0.14211f
C1750 XThC.XTBN.Y XThC.Tn[0] 0.45269f
C1751 XA.XIR[10].XIC[0].icell.PDM VPWR 0.01171f
C1752 XA.XIR[7].XIC_dummy_left.icell.Iout XA.XIR[8].XIC_dummy_left.icell.Iout 0.03665f
C1753 XThC.Tn[2] XA.XIR[15].XIC[2].icell.Ien 0.04292f
C1754 XThR.Tn[3] XA.XIR[3].XIC[13].icell.Ien 0.14211f
C1755 XThC.Tn[6] XThR.Tn[4] 0.40738f
C1756 XA.XIR[14].XIC[13].icell.Ien Vbias 0.19161f
C1757 XA.XIR[9].XIC[12].icell.PDM Vbias 0.03928f
C1758 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.Ien 0.04854f
C1759 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.Ien 0.04854f
C1760 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout 0.06446f
C1761 XThC.Tn[13] XA.XIR[9].XIC[13].icell.Ien 0.04604f
C1762 XA.XIR[15].XIC[4].icell.Ien VPWR 0.31713f
C1763 XA.XIR[0].XIC[4].icell.PDM Vbias 0.03945f
C1764 XThC.Tn[1] XThR.Tn[10] 0.40738f
C1765 XThC.Tn[3] XA.XIR[11].XIC[3].icell.Ien 0.04604f
C1766 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PDM 0.02601f
C1767 XThR.Tn[2] XA.XIR[2].XIC[8].icell.Ien 0.14211f
C1768 XA.XIR[1].XIC[1].icell.Ien Vbias 0.19173f
C1769 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PDM 0.02601f
C1770 XA.XIR[10].XIC[2].icell.Ien Vbias 0.19161f
C1771 XA.XIR[4].XIC[7].icell.Ien VPWR 0.18829f
C1772 XA.XIR[9].XIC[1].icell.Ien Iout 0.06801f
C1773 XThR.Tn[9] XA.XIR[9].XIC[1].icell.Ien 0.14211f
C1774 XThR.XTB7.Y a_n997_715# 0.06874f
C1775 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PDM 0.02803f
C1776 XA.XIR[4].XIC[3].icell.Ien Iout 0.06801f
C1777 XThC.Tn[14] XA.XIR[1].XIC[14].icell.Ien 0.04606f
C1778 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PDM 0.02601f
C1779 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PDM 0.02601f
C1780 XThC.Tn[8] XA.XIR[12].XIC[8].icell.Ien 0.04604f
C1781 XA.XIR[3].XIC[11].icell.Ien Vbias 0.19161f
C1782 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1783 XA.XIR[3].XIC_dummy_left.icell.Iout XA.XIR[4].XIC_dummy_left.icell.Iout 0.03665f
C1784 XA.XIR[7].XIC[1].icell.Ien VPWR 0.18829f
C1785 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13] 0.14211f
C1786 XA.XIR[0].XIC[8].icell.PDM VPWR 0.01451f
C1787 XThC.XTB5.Y VPWR 1.01219f
C1788 XA.XIR[2].XIC[4].icell.Ien Vbias 0.19161f
C1789 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PDM 0.02601f
C1790 XA.XIR[9].XIC[10].icell.Ien VPWR 0.18829f
C1791 XA.XIR[1].XIC[6].icell.Ien Vbias 0.19173f
C1792 XA.XIR[9].XIC[6].icell.Ien Iout 0.06801f
C1793 XA.XIR[14].XIC_dummy_left.icell.Iout Iout 0.03553f
C1794 XA.XIR[12].XIC[14].icell.Ien VPWR 0.18835f
C1795 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.Ien 0.04854f
C1796 XThR.Tn[9] XA.XIR[9].XIC[6].icell.Ien 0.14211f
C1797 XA.XIR[0].XIC[3].icell.Ien VPWR 0.18776f
C1798 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PDM 0.04035f
C1799 XA.XIR[8].XIC[14].icell.Ien Vbias 0.19161f
C1800 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PDM 0.04035f
C1801 XA.XIR[7].XIC[6].icell.Ien VPWR 0.18829f
C1802 XThC.XTBN.Y VPWR 4.12335f
C1803 XA.XIR[7].XIC[2].icell.Ien Iout 0.06801f
C1804 XA.XIR[5].XIC_15.icell.Ien Iout 0.0694f
C1805 XThC.XTB6.Y a_6243_9615# 0.01199f
C1806 XThC.Tn[11] XA.XIR[8].XIC[11].icell.Ien 0.04604f
C1807 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.PDM 0.02104f
C1808 XThR.XTB7.A XThR.XTBN.A 0.19736f
C1809 a_n1049_6699# VPWR 0.72162f
C1810 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.PDM 0.02104f
C1811 XA.XIR[14].XIC[11].icell.Ien Vbias 0.19161f
C1812 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1813 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PDM 0.02601f
C1814 XA.XIR[5].XIC[2].icell.PDM Vbias 0.03928f
C1815 XThR.XTB7.A XThR.Tn[6] 0.1056f
C1816 XThC.XTB1.Y XThC.Tn[8] 0.29214f
C1817 XA.XIR[6].XIC[1].icell.Ien Vbias 0.19161f
C1818 XThR.Tn[11] XA.XIR[11].XIC[2].icell.Ien 0.14211f
C1819 XThC.Tn[10] VPWR 4.54895f
C1820 XA.XIR[12].XIC[1].icell.PDM Vbias 0.03928f
C1821 XThC.Tn[14] XA.XIR[6].XIC[14].icell.Ien 0.04604f
C1822 XThC.Tn[5] XA.XIR[2].XIC[5].icell.Ien 0.04605f
C1823 XThR.Tn[2] Vbias 1.39527f
C1824 XThR.Tn[4] XA.XIR[4].XIC_15.icell.Ien 0.13564f
C1825 a_4861_9615# VPWR 0.70519f
C1826 XThC.Tn[13] XA.XIR[11].XIC[13].icell.Ien 0.04604f
C1827 XThR.Tn[9] Iout 1.12762f
C1828 XA.XIR[11].XIC[7].icell.PDM Vbias 0.03928f
C1829 XA.XIR[5].XIC_dummy_right.icell.Iout Iout 0.01732f
C1830 XThR.Tn[0] XA.XIR[0].XIC[7].icell.Ien 0.14211f
C1831 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PDM 0.04035f
C1832 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1833 XThR.Tn[10] XA.XIR[10].XIC[6].icell.Ien 0.14211f
C1834 XA.XIR[5].XIC[6].icell.PDM VPWR 0.01171f
C1835 XThC.Tn[10] XA.XIR[13].XIC[10].icell.Ien 0.04604f
C1836 XA.XIR[13].XIC[0].icell.PDM VPWR 0.01171f
C1837 XThR.Tn[7] XA.XIR[7].XIC[8].icell.Ien 0.14211f
C1838 XA.XIR[6].XIC[6].icell.Ien Vbias 0.19161f
C1839 XThC.XTB5.Y a_9827_9569# 0.06458f
C1840 XA.XIR[12].XIC[5].icell.PDM VPWR 0.01171f
C1841 XA.XIR[12].XIC[12].icell.Ien VPWR 0.18829f
C1842 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.PDM 0.02104f
C1843 XA.XIR[15].XIC[0].icell.Ien Iout 0.07185f
C1844 XThC.Tn[3] XA.XIR[14].XIC[3].icell.Ien 0.04604f
C1845 XThC.Tn[1] XThR.Tn[13] 0.40738f
C1846 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PDM 0.02601f
C1847 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.Ien 0.04854f
C1848 XA.XIR[2].XIC[3].icell.PDM Vbias 0.03928f
C1849 XA.XIR[8].XIC[1].icell.Ien VPWR 0.18829f
C1850 XA.XIR[13].XIC[2].icell.Ien Vbias 0.19161f
C1851 XA.XIR[3].XIC[3].icell.Ien VPWR 0.18829f
C1852 XA.XIR[15].XIC_15.icell.PUM VPWR 0.01655f
C1853 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PDM 0.04035f
C1854 XThC.Tn[4] Iout 0.22518f
C1855 XThC.Tn[4] XThR.Tn[9] 0.40738f
C1856 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PDM 0.02601f
C1857 XThC.Tn[0] XThR.Tn[8] 0.40736f
C1858 XThC.Tn[0] XA.XIR[3].XIC[0].icell.Ien 0.04604f
C1859 XThR.XTB7.A XThR.Tn[4] 0.02736f
C1860 XA.XIR[15].XIC[9].icell.Ien VPWR 0.31713f
C1861 XA.XIR[11].XIC[5].icell.Ien Vbias 0.19161f
C1862 XThC.XTBN.Y a_9827_9569# 0.22873f
C1863 XThR.Tn[2] XA.XIR[2].XIC[13].icell.Ien 0.14211f
C1864 XThR.XTB7.A a_n1049_7493# 0.0127f
C1865 XA.XIR[15].XIC[5].icell.Ien Iout 0.07192f
C1866 XA.XIR[4].XIC[12].icell.Ien VPWR 0.18829f
C1867 XA.XIR[8].XIC[3].icell.PDM VPWR 0.01171f
C1868 XA.XIR[3].XIC[1].icell.PDM VPWR 0.01171f
C1869 XA.XIR[10].XIC[7].icell.Ien Vbias 0.19161f
C1870 XThC.XTB5.Y XThC.XTB7.B 0.30234f
C1871 data[1] data[2] 0.01393f
C1872 XA.XIR[4].XIC[8].icell.Ien Iout 0.06801f
C1873 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14] 0.14211f
C1874 XA.XIR[2].XIC[7].icell.PDM VPWR 0.01171f
C1875 XA.XIR[8].XIC[6].icell.Ien VPWR 0.18829f
C1876 XThR.XTB7.A XThR.XTB6.Y 0.19112f
C1877 XA.XIR[8].XIC[2].icell.Ien Iout 0.06801f
C1878 XA.XIR[2].XIC[9].icell.Ien Vbias 0.19161f
C1879 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PDM 0.04035f
C1880 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.Ien 0.04854f
C1881 XA.XIR[9].XIC_15.icell.Ien VPWR 0.26829f
C1882 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.PDM 0.02104f
C1883 XA.XIR[1].XIC[11].icell.Ien Vbias 0.19173f
C1884 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.PDM 0.02104f
C1885 XThR.XTB7.B XThR.XTBN.A 0.35142f
C1886 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1887 XThR.XTB7.Y XThR.Tn[11] 0.07412f
C1888 XA.XIR[9].XIC[11].icell.Ien Iout 0.06801f
C1889 XThC.XTB7.B XThC.XTBN.Y 0.38751f
C1890 XThR.Tn[9] XA.XIR[9].XIC[11].icell.Ien 0.14211f
C1891 XA.XIR[0].XIC[8].icell.Ien VPWR 0.18959f
C1892 XThR.XTB7.B XThR.Tn[6] 0.04822f
C1893 XA.XIR[0].XIC[4].icell.Ien Iout 0.0675f
C1894 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PDM 0.04035f
C1895 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.PDM 0.02104f
C1896 XA.XIR[12].XIC[10].icell.Ien VPWR 0.18829f
C1897 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PDM 0.04035f
C1898 XA.XIR[7].XIC[11].icell.Ien VPWR 0.18829f
C1899 XThC.Tn[12] XThR.Tn[7] 0.40738f
C1900 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.Ien 0.04854f
C1901 XA.XIR[7].XIC[7].icell.Ien Iout 0.06801f
C1902 XA.XIR[7].XIC[3].icell.PDM Vbias 0.03928f
C1903 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PDM 0.04035f
C1904 XThR.Tn[10] Vbias 1.39532f
C1905 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PDM 0.02601f
C1906 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.Ien 0.04854f
C1907 XThC.XTB7.B XThC.Tn[10] 0.0672f
C1908 XA.XIR[9].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1909 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.Ien 0.04854f
C1910 XThC.XTB7.Y XThC.Tn[14] 0.4237f
C1911 XA.XIR[15].XIC[1].icell.PDM Vbias 0.03928f
C1912 XA.XIR[6].XIC[10].icell.PDM Vbias 0.03928f
C1913 XThR.Tn[6] XA.XIR[6].XIC[1].icell.Ien 0.14211f
C1914 XThC.Tn[9] Vbias 0.79809f
C1915 XThR.Tn[8] VPWR 8.93422f
C1916 XA.XIR[3].XIC[0].icell.Ien VPWR 0.18829f
C1917 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PDM 0.02601f
C1918 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.PDM 0.02104f
C1919 XThC.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.04604f
C1920 XA.XIR[14].XIC[7].icell.PDM Vbias 0.03928f
C1921 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1922 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.PDM 0.02104f
C1923 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.PDM 0.02104f
C1924 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PDM 0.02601f
C1925 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.Ien 0.04854f
C1926 XA.XIR[11].XIC[1].icell.Ien VPWR 0.18829f
C1927 XThC.Tn[8] XA.XIR[15].XIC[8].icell.Ien 0.04292f
C1928 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PDM 0.04035f
C1929 XThR.Tn[11] XA.XIR[11].XIC[7].icell.Ien 0.14211f
C1930 XThC.Tn[4] XA.XIR[0].XIC[4].icell.Ien 0.04658f
C1931 XA.XIR[7].XIC[7].icell.PDM VPWR 0.01171f
C1932 XThC.XTB7.A data[1] 0.06544f
C1933 a_3773_9615# XThC.Tn[1] 0.26251f
C1934 XThR.XTB2.Y XThR.XTB3.Y 2.04808f
C1935 XThR.Tn[14] a_n997_715# 0.1927f
C1936 XThR.Tn[0] XA.XIR[0].XIC[12].icell.Ien 0.14211f
C1937 XA.XIR[15].XIC[5].icell.PDM VPWR 0.01512f
C1938 XA.XIR[6].XIC[14].icell.PDM VPWR 0.0118f
C1939 XThR.Tn[11] a_n997_2667# 0.19413f
C1940 XThC.Tn[9] XA.XIR[11].XIC[9].icell.Ien 0.04604f
C1941 XThR.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.14211f
C1942 XThC.Tn[11] XThR.Tn[3] 0.40738f
C1943 XA.XIR[9].XIC_dummy_right.icell.Iout XA.XIR[10].XIC_dummy_right.icell.Iout 0.04047f
C1944 XA.XIR[15].XIC[14].icell.Ien VPWR 0.31908f
C1945 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Ien 0.01569f
C1946 XA.XIR[1].XIC[4].icell.PDM Vbias 0.03928f
C1947 XA.XIR[6].XIC[11].icell.Ien Vbias 0.19161f
C1948 XThR.Tn[7] XA.XIR[7].XIC[13].icell.Ien 0.14211f
C1949 XA.XIR[9].XIC[3].icell.PDM VPWR 0.01171f
C1950 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.Ien 0.04854f
C1951 XA.XIR[4].XIC[4].icell.PDM Vbias 0.03928f
C1952 XThC.Tn[6] XA.XIR[4].XIC[6].icell.Ien 0.04604f
C1953 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.Ien 0.04854f
C1954 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PDM 0.02602f
C1955 XA.XIR[3].XIC[12].icell.PDM Vbias 0.03928f
C1956 XThC.Tn[14] XThR.Tn[0] 0.40766f
C1957 XA.XIR[8].XIC[14].icell.PDM Vbias 0.03928f
C1958 XThC.XTB4.Y a_8963_9569# 0.07199f
C1959 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.PDM 0.02104f
C1960 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.PDM 0.02104f
C1961 XA.XIR[14].XIC[5].icell.Ien Vbias 0.19161f
C1962 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.Ien 0.04854f
C1963 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.PDM 0.02104f
C1964 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PDM 0.02601f
C1965 XA.XIR[13].XIC[7].icell.Ien Vbias 0.19161f
C1966 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PDM 0.04035f
C1967 XThR.XTB7.B XThR.XTB6.Y 0.30244f
C1968 XA.XIR[3].XIC[8].icell.Ien VPWR 0.18829f
C1969 XA.XIR[1].XIC[8].icell.PDM VPWR 0.01171f
C1970 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.PDM 0.02104f
C1971 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.Ien 0.04854f
C1972 XA.XIR[3].XIC[4].icell.Ien Iout 0.06801f
C1973 XA.XIR[10].XIC[13].icell.Ien Iout 0.06801f
C1974 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.Ien 0.04854f
C1975 XA.XIR[4].XIC[8].icell.PDM VPWR 0.01171f
C1976 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout 0.06446f
C1977 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PDM 0.04035f
C1978 XThR.XTBN.Y XThR.XTBN.A 0.77119f
C1979 XA.XIR[1].XIC[3].icell.Ien VPWR 0.18829f
C1980 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.PDM 0.02104f
C1981 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1982 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PDM 0.02601f
C1983 XThC.XTB7.Y a_6243_10571# 0.01283f
C1984 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.Ien 0.04854f
C1985 a_n1049_7493# XThR.Tn[2] 0.26564f
C1986 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.Ien 0.04854f
C1987 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.Ien 0.04854f
C1988 XA.XIR[4].XIC[13].icell.Ien Iout 0.06801f
C1989 XThR.XTBN.Y XThR.Tn[6] 0.59897f
C1990 XA.XIR[12].XIC_15.icell.Ien VPWR 0.26829f
C1991 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PDM 0.04035f
C1992 XA.XIR[8].XIC[11].icell.Ien VPWR 0.18829f
C1993 XThR.XTB7.Y XThR.Tn[14] 0.4222f
C1994 XA.XIR[8].XIC[7].icell.Ien Iout 0.06801f
C1995 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.PDM 0.02104f
C1996 XThC.XTB5.A data[1] 0.11102f
C1997 XThC.Tn[13] XThR.Tn[2] 0.40742f
C1998 XA.XIR[2].XIC[14].icell.Ien Vbias 0.19161f
C1999 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.Ien 0.04854f
C2000 XThR.XTB2.Y VPWR 0.98845f
C2001 a_n997_3755# VPWR 0.0133f
C2002 XThR.XTB4.Y XThR.XTBN.A 0.03415f
C2003 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PDM 0.04035f
C2004 XA.XIR[14].XIC[0].icell.Ien Vbias 0.19149f
C2005 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PDM 0.02601f
C2006 XThC.Tn[4] XA.XIR[3].XIC[4].icell.Ien 0.04604f
C2007 XA.XIR[0].XIC[13].icell.Ien VPWR 0.18776f
C2008 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout 0.06446f
C2009 XA.XIR[15].XIC[12].icell.Ien VPWR 0.31713f
C2010 XThR.XTB5.Y XThR.Tn[5] 0.01094f
C2011 VPWR data[2] 0.21031f
C2012 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PDM 0.02601f
C2013 XThR.XTBN.A XThR.Tn[10] 0.12147f
C2014 XThR.Tn[13] Vbias 1.39532f
C2015 XThR.Tn[14] XA.XIR[14].XIC[2].icell.Ien 0.14211f
C2016 XThC.Tn[11] XA.XIR[2].XIC[11].icell.Ien 0.04605f
C2017 XThR.Tn[1] XA.XIR[1].XIC[2].icell.Ien 0.14211f
C2018 XA.XIR[0].XIC[9].icell.Ien Iout 0.0675f
C2019 XA.XIR[12].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2020 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PDM 0.02601f
C2021 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PDM 0.04035f
C2022 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PDM 0.02602f
C2023 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2024 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PDM 0.02601f
C2025 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.PDM 0.02104f
C2026 XThR.Tn[13] XA.XIR[13].XIC[6].icell.Ien 0.14211f
C2027 a_n1049_5611# VPWR 0.71817f
C2028 XA.XIR[7].XIC[12].icell.Ien Iout 0.06801f
C2029 XThC.Tn[9] XThR.Tn[6] 0.40738f
C2030 XA.XIR[5].XIC[4].icell.Ien Vbias 0.19161f
C2031 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.Ien 0.04854f
C2032 XA.XIR[14].XIC[1].icell.Ien VPWR 0.18883f
C2033 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.Ien 0.04854f
C2034 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.Ien 0.04854f
C2035 XA.XIR[10].XIC[2].icell.PDM VPWR 0.01171f
C2036 XA.XIR[10].XIC[11].icell.Ien Iout 0.06801f
C2037 XThC.Tn[11] XThR.Tn[11] 0.40738f
C2038 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.PDM 0.02104f
C2039 XA.XIR[3].XIC[1].icell.Ien Iout 0.06801f
C2040 XThR.XTBN.Y XThR.Tn[4] 0.6035f
C2041 XThC.Tn[9] XA.XIR[14].XIC[9].icell.Ien 0.04604f
C2042 XThC.Tn[1] XThR.Tn[7] 0.40738f
C2043 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.PDM 0.02104f
C2044 XA.XIR[6].XIC[3].icell.Ien VPWR 0.18829f
C2045 XA.XIR[9].XIC[14].icell.PDM Vbias 0.03928f
C2046 XThR.XTBN.Y a_n1049_7493# 0.08456f
C2047 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.Ien 0.04854f
C2048 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.PDM 0.02104f
C2049 XA.XIR[0].XIC[6].icell.PDM Vbias 0.03945f
C2050 XThC.XTB7.B a_7651_9569# 0.01152f
C2051 XThC.XTB5.Y XThC.Tn[12] 0.32158f
C2052 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.PDM 0.02104f
C2053 XA.XIR[9].XIC_dummy_left.icell.Iout Iout 0.03553f
C2054 XThC.Tn[7] Vbias 0.82088f
C2055 XThR.Tn[9] XA.XIR[9].XIC_dummy_left.icell.Iout 0.03386f
C2056 XThR.XTBN.Y XThR.XTB6.Y 0.1894f
C2057 XThR.Tn[6] XA.XIR[6].XIC[11].icell.Ien 0.14211f
C2058 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.PDM 0.02104f
C2059 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.PDM 0.02104f
C2060 XThC.Tn[2] XA.XIR[10].XIC[2].icell.Ien 0.04604f
C2061 XThC.Tn[14] XThR.Tn[1] 0.40747f
C2062 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PDM 0.02601f
C2063 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout 0.06446f
C2064 XA.XIR[2].XIC[1].icell.Ien VPWR 0.18829f
C2065 XThR.XTB3.Y XThR.Tn[3] 0.01287f
C2066 XA.XIR[7].XIC_dummy_left.icell.Iout VPWR 0.10954f
C2067 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.Ien 0.04854f
C2068 XA.XIR[0].XIC[10].icell.PDM VPWR 0.01132f
C2069 XA.XIR[11].XIC[2].icell.Ien VPWR 0.18829f
C2070 XThC.Tn[14] XThR.Tn[12] 0.40742f
C2071 XA.XIR[15].XIC[10].icell.Ien VPWR 0.31713f
C2072 XA.XIR[13].XIC[13].icell.Ien Iout 0.06801f
C2073 XThC.XTB7.A VPWR 0.87269f
C2074 XA.XIR[10].XIC[4].icell.Ien VPWR 0.18829f
C2075 XThC.Tn[0] XThR.Tn[3] 0.40742f
C2076 XThC.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.04604f
C2077 XThR.XTBN.A a_n997_1803# 0.09118f
C2078 XThC.XTBN.Y XThC.Tn[12] 0.46758f
C2079 XThR.XTB3.Y data[4] 0.03253f
C2080 XThR.XTB4.Y XThR.XTB6.Y 0.04273f
C2081 XThC.Tn[9] XThR.Tn[4] 0.40738f
C2082 XThR.XTB3.Y XThR.XTB7.Y 0.03772f
C2083 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PDM 0.04035f
C2084 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PDM 0.02601f
C2085 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PDM 0.04035f
C2086 XA.XIR[3].XIC[13].icell.Ien VPWR 0.18829f
C2087 XA.XIR[3].XIC[9].icell.Ien Iout 0.06801f
C2088 XThR.XTB6.Y XThR.Tn[10] 0.02461f
C2089 XA.XIR[2].XIC[6].icell.Ien VPWR 0.18829f
C2090 XThC.Tn[3] XThR.Tn[0] 0.40763f
C2091 XThC.Tn[13] XThR.Tn[10] 0.40739f
C2092 XThC.Tn[5] XThR.Tn[5] 0.40738f
C2093 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.PDM 0.02104f
C2094 a_n997_715# VPWR 0.02818f
C2095 XA.XIR[2].XIC[2].icell.Ien Iout 0.06801f
C2096 XA.XIR[1].XIC[8].icell.Ien VPWR 0.18829f
C2097 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2098 XThR.Tn[8] XA.XIR[8].XIC[3].icell.Ien 0.14211f
C2099 XThR.Tn[10] XA.XIR[10].XIC_dummy_left.icell.Iout 0.03385f
C2100 a_3773_9615# Vbias 0.01444f
C2101 XA.XIR[1].XIC[4].icell.Ien Iout 0.06801f
C2102 XA.XIR[5].XIC[4].icell.PDM Vbias 0.03928f
C2103 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PDM 0.02601f
C2104 XA.XIR[8].XIC[12].icell.Ien Iout 0.06801f
C2105 XThC.XTB7.B data[2] 0.07481f
C2106 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.PDM 0.02104f
C2107 XThR.Tn[5] XA.XIR[5].XIC[2].icell.Ien 0.14211f
C2108 XA.XIR[12].XIC[3].icell.PDM Vbias 0.03928f
C2109 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PDM 0.02601f
C2110 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.PDM 0.02104f
C2111 XThC.Tn[3] XA.XIR[9].XIC[3].icell.Ien 0.04604f
C2112 XA.XIR[11].XIC[9].icell.PDM Vbias 0.03928f
C2113 a_5949_9615# VPWR 0.7053f
C2114 XThC.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.04604f
C2115 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.Ien 0.04854f
C2116 XA.XIR[6].XIC[1].icell.PDM VPWR 0.01171f
C2117 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PDM 0.04035f
C2118 XThC.Tn[10] XA.XIR[0].XIC[10].icell.Ien 0.04662f
C2119 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.PDM 0.02104f
C2120 XThR.Tn[14] XA.XIR[14].XIC[7].icell.Ien 0.14211f
C2121 XA.XIR[0].XIC[14].icell.Ien Iout 0.0675f
C2122 XThR.Tn[1] XA.XIR[1].XIC[7].icell.Ien 0.14211f
C2123 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.PDM 0.02104f
C2124 XA.XIR[5].XIC[8].icell.PDM VPWR 0.01171f
C2125 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.PDM 0.02104f
C2126 XThC.Tn[2] XThR.Tn[2] 0.40741f
C2127 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.PDM 0.02104f
C2128 XA.XIR[13].XIC[2].icell.PDM VPWR 0.01171f
C2129 XThC.Tn[4] XA.XIR[1].XIC[4].icell.Ien 0.04607f
C2130 XA.XIR[13].XIC[11].icell.Ien Iout 0.06801f
C2131 XThC.Tn[11] XThR.Tn[14] 0.40738f
C2132 XThR.Tn[3] VPWR 8.06517f
C2133 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.PDM 0.02104f
C2134 XThC.XTB5.A VPWR 0.82807f
C2135 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout 0.06446f
C2136 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.Ien 0.04854f
C2137 XA.XIR[12].XIC[7].icell.PDM VPWR 0.01171f
C2138 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.Ien 0.04854f
C2139 XA.XIR[5].XIC[9].icell.Ien Vbias 0.19161f
C2140 XA.XIR[12].XIC_dummy_right.icell.Iout XA.XIR[13].XIC_dummy_right.icell.Iout 0.04047f
C2141 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.Ien 0.04854f
C2142 XA.XIR[8].XIC[1].icell.PDM Vbias 0.03928f
C2143 VPWR data[4] 0.5303f
C2144 XThR.XTB7.Y VPWR 1.14768f
C2145 XA.XIR[2].XIC[5].icell.PDM Vbias 0.03928f
C2146 XThC.Tn[12] XA.XIR[4].XIC[12].icell.Ien 0.04604f
C2147 XThR.XTB5.A XThR.XTB5.Y 0.0538f
C2148 XA.XIR[8].XIC_dummy_left.icell.Iout VPWR 0.11f
C2149 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.Ien 0.04854f
C2150 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PDM 0.04035f
C2151 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.Ien 0.04854f
C2152 XA.XIR[15].XIC_15.icell.Ien VPWR 0.37868f
C2153 XA.XIR[12].XIC[4].icell.Ien Vbias 0.19161f
C2154 XA.XIR[6].XIC[8].icell.Ien VPWR 0.18829f
C2155 XThC.Tn[7] XThR.Tn[6] 0.40738f
C2156 XThC.XTBN.A XThC.Tn[9] 0.12399f
C2157 XThC.Tn[0] XA.XIR[12].XIC[0].icell.Ien 0.04604f
C2158 XA.XIR[6].XIC[4].icell.Ien Iout 0.06801f
C2159 XThC.Tn[2] XA.XIR[13].XIC[2].icell.Ien 0.04604f
C2160 XThC.XTBN.Y a_10915_9569# 0.21503f
C2161 XA.XIR[3].XIC[3].icell.PDM VPWR 0.01171f
C2162 XThC.Tn[0] XThR.Tn[11] 0.4074f
C2163 XA.XIR[14].XIC[2].icell.Ien VPWR 0.18883f
C2164 XA.XIR[8].XIC[5].icell.PDM VPWR 0.01171f
C2165 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.Ien 0.04854f
C2166 XA.XIR[2].XIC[9].icell.PDM VPWR 0.01171f
C2167 XThC.XTB7.A XThC.XTB7.B 0.35844f
C2168 XA.XIR[13].XIC[4].icell.Ien VPWR 0.18829f
C2169 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.PDM 0.02104f
C2170 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PDM 0.02601f
C2171 XThC.Tn[1] XA.XIR[7].XIC[1].icell.Ien 0.04604f
C2172 XA.XIR[10].XIC_15.icell.PUM VPWR 0.01655f
C2173 XA.XIR[15].XIC_dummy_right.icell.Iout VPWR 0.21463f
C2174 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.Ien 0.04854f
C2175 XA.XIR[11].XIC[7].icell.Ien VPWR 0.18829f
C2176 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.PDM 0.02104f
C2177 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PDM 0.04035f
C2178 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.PDM 0.02104f
C2179 XThC.XTB6.Y XThC.Tn[5] 0.20249f
C2180 XThR.XTB6.Y XThR.Tn[13] 0.32265f
C2181 XA.XIR[11].XIC[3].icell.Ien Iout 0.06801f
C2182 XA.XIR[10].XIC[9].icell.Ien VPWR 0.18829f
C2183 XThC.Tn[13] XThR.Tn[13] 0.40739f
C2184 XThC.Tn[3] XThR.Tn[1] 0.40744f
C2185 XA.XIR[10].XIC[5].icell.Ien Iout 0.06801f
C2186 a_n997_2667# VPWR 0.01642f
C2187 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.Ien 0.04854f
C2188 XThC.Tn[4] XA.XIR[6].XIC[4].icell.Ien 0.04604f
C2189 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2190 XThR.XTB5.A XThR.XTB1.Y 0.1098f
C2191 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PDM 0.04035f
C2192 XThC.Tn[3] XThR.Tn[12] 0.40738f
C2193 XThC.Tn[10] XA.XIR[3].XIC[10].icell.Ien 0.04604f
C2194 XThC.Tn[12] XThR.Tn[8] 0.40738f
C2195 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR 0.38522f
C2196 XA.XIR[3].XIC[14].icell.Ien Iout 0.06801f
C2197 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PDM 0.04035f
C2198 XThR.Tn[7] Vbias 1.39526f
C2199 XA.XIR[2].XIC[11].icell.Ien VPWR 0.18829f
C2200 XThC.Tn[5] XA.XIR[12].XIC[5].icell.Ien 0.04604f
C2201 XThC.XTBN.Y XThC.Tn[1] 0.49539f
C2202 XA.XIR[2].XIC[7].icell.Ien Iout 0.06801f
C2203 XA.XIR[1].XIC[13].icell.Ien VPWR 0.18829f
C2204 XThR.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.14211f
C2205 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PDM 0.04035f
C2206 XA.XIR[7].XIC[5].icell.PDM Vbias 0.03928f
C2207 XThC.Tn[7] XThR.Tn[4] 0.40738f
C2208 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.Ien 0.04854f
C2209 XA.XIR[1].XIC[9].icell.Ien Iout 0.06801f
C2210 XA.XIR[15].XIC[3].icell.PDM Vbias 0.03928f
C2211 XA.XIR[4].XIC[2].icell.Ien Vbias 0.19161f
C2212 XA.XIR[6].XIC[12].icell.PDM Vbias 0.03928f
C2213 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Iout 0.03777f
C2214 VPWR bias[1] 1.33312f
C2215 XThC.Tn[2] XThR.Tn[10] 0.40738f
C2216 XA.XIR[14].XIC[9].icell.PDM Vbias 0.03928f
C2217 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.Ien 0.04854f
C2218 XA.XIR[12].XIC[0].icell.Ien VPWR 0.18829f
C2219 XThC.XTB6.Y a_10051_9569# 0.07626f
C2220 XThR.Tn[11] VPWR 9.00382f
C2221 XThR.Tn[5] XA.XIR[5].XIC[7].icell.Ien 0.14211f
C2222 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PDM 0.04035f
C2223 XA.XIR[9].XIC[1].icell.PDM Vbias 0.03928f
C2224 XA.XIR[7].XIC[9].icell.PDM VPWR 0.01171f
C2225 XThC.XTB5.A XThC.XTB7.B 0.30355f
C2226 XA.XIR[9].XIC[5].icell.Ien Vbias 0.19161f
C2227 XA.XIR[15].XIC[7].icell.PDM VPWR 0.01512f
C2228 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2229 XThR.Tn[1] XA.XIR[1].XIC[12].icell.Ien 0.14211f
C2230 XA.XIR[1].XIC[6].icell.PDM Vbias 0.03928f
C2231 XThR.XTB5.Y XThR.Tn[9] 0.01732f
C2232 XA.XIR[9].XIC[5].icell.PDM VPWR 0.01171f
C2233 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.Ien 0.04854f
C2234 XA.XIR[4].XIC[6].icell.PDM Vbias 0.03928f
C2235 XA.XIR[5].XIC[14].icell.Ien Vbias 0.19161f
C2236 XThC.Tn[8] XA.XIR[10].XIC[8].icell.Ien 0.04604f
C2237 XA.XIR[3].XIC[14].icell.PDM Vbias 0.03928f
C2238 XThR.XTBN.A a_n997_3979# 0.02087f
C2239 XThC.Tn[1] XA.XIR[8].XIC[1].icell.Ien 0.04604f
C2240 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.Ien 0.04854f
C2241 XThC.Tn[0] XThR.Tn[14] 0.40739f
C2242 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.PDM 0.02104f
C2243 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.Ien 0.04854f
C2244 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.04035f
C2245 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PDM 0.02601f
C2246 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.PDM 0.02104f
C2247 XA.XIR[1].XIC[10].icell.PDM VPWR 0.01171f
C2248 XThC.Tn[11] XA.XIR[5].XIC[11].icell.Ien 0.04604f
C2249 XA.XIR[12].XIC[9].icell.Ien Vbias 0.19161f
C2250 XA.XIR[6].XIC[13].icell.Ien VPWR 0.18829f
C2251 XA.XIR[10].XIC[14].icell.Ien VPWR 0.18835f
C2252 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2253 XA.XIR[4].XIC[10].icell.PDM VPWR 0.01171f
C2254 XA.XIR[6].XIC[9].icell.Ien Iout 0.06801f
C2255 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PDM 0.02601f
C2256 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PDM 0.04035f
C2257 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PDM 0.02602f
C2258 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PDM 0.02601f
C2259 XA.XIR[13].XIC_15.icell.PUM VPWR 0.01655f
C2260 XA.XIR[9].XIC[0].icell.Ien Vbias 0.19149f
C2261 XA.XIR[14].XIC[7].icell.Ien VPWR 0.18883f
C2262 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2263 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PDM 0.04035f
C2264 XA.XIR[14].XIC[3].icell.Ien Iout 0.06801f
C2265 XA.XIR[13].XIC[9].icell.Ien VPWR 0.18829f
C2266 XThC.Tn[12] XA.XIR[15].XIC[12].icell.Ien 0.04292f
C2267 XThC.Tn[11] VPWR 4.57828f
C2268 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.Ien 0.04854f
C2269 XA.XIR[13].XIC[5].icell.Ien Iout 0.06801f
C2270 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2271 XThC.XTBN.A XThC.Tn[7] 0.01451f
C2272 XThR.Tn[12] XA.XIR[12].XIC[13].icell.Ien 0.14211f
C2273 XThR.Tn[13] XA.XIR[13].XIC_dummy_left.icell.Iout 0.03385f
C2274 XA.XIR[11].XIC[8].icell.Ien Iout 0.06801f
C2275 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PDM 0.04035f
C2276 XThR.XTBN.A XThR.Tn[7] 0.01439f
C2277 XThR.XTBN.A a_n997_2891# 0.01719f
C2278 XA.XIR[10].XIC[0].icell.PDM Vbias 0.03915f
C2279 XThR.Tn[6] XThR.Tn[7] 0.11401f
C2280 XThC.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.04604f
C2281 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PDM 0.04056f
C2282 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PDM 0.04035f
C2283 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.Ien 0.04854f
C2284 XThC.Tn[2] XThR.Tn[13] 0.40738f
C2285 data[6] data[7] 0.04128f
C2286 XA.XIR[5].XIC[1].icell.Ien VPWR 0.18829f
C2287 XA.XIR[2].XIC[12].icell.Ien Iout 0.06801f
C2288 XA.XIR[15].XIC[4].icell.Ien Vbias 0.15966f
C2289 XThR.Tn[8] XA.XIR[8].XIC[13].icell.Ien 0.14211f
C2290 XThR.Tn[14] VPWR 9.25423f
C2291 XThC.Tn[10] XA.XIR[1].XIC[10].icell.Ien 0.04606f
C2292 XA.XIR[11].XIC[0].icell.PDM VPWR 0.01171f
C2293 XA.XIR[1].XIC[14].icell.Ien Iout 0.06801f
C2294 XThC.Tn[5] Iout 0.22432f
C2295 XThC.Tn[5] XThR.Tn[9] 0.40738f
C2296 XA.XIR[4].XIC[7].icell.Ien Vbias 0.19161f
C2297 XThC.Tn[1] XThR.Tn[8] 0.40738f
C2298 XThR.XTB2.Y a_n1335_8107# 0.01006f
C2299 XA.XIR[10].XIC[4].icell.PDM VPWR 0.01171f
C2300 XA.XIR[10].XIC[12].icell.Ien VPWR 0.18829f
C2301 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.Ien 0.04854f
C2302 XA.XIR[3].XIC_dummy_left.icell.Iout Iout 0.03553f
C2303 bias[1] bias[0] 0.56718f
C2304 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PDM 0.02601f
C2305 XThC.Tn[1] XA.XIR[11].XIC[1].icell.Ien 0.04604f
C2306 XA.XIR[12].XIC[1].icell.Ien Iout 0.06801f
C2307 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.Ien 0.04854f
C2308 VPWR data[1] 0.44103f
C2309 XThR.Tn[5] XA.XIR[5].XIC[12].icell.Ien 0.14211f
C2310 XThC.XTB6.Y XThC.XTB7.Y 2.05133f
C2311 XA.XIR[0].XIC[8].icell.PDM Vbias 0.03945f
C2312 XA.XIR[7].XIC[1].icell.Ien Vbias 0.19161f
C2313 XA.XIR[5].XIC[6].icell.Ien VPWR 0.18829f
C2314 XThC.XTB5.Y Vbias 0.01606f
C2315 XThC.XTB7.B a_8739_9569# 0.0168f
C2316 XA.XIR[9].XIC[10].icell.Ien Vbias 0.19161f
C2317 XA.XIR[5].XIC[2].icell.Ien Iout 0.06801f
C2318 XThC.Tn[14] XA.XIR[7].XIC[14].icell.Ien 0.04604f
C2319 XA.XIR[12].XIC[14].icell.Ien Vbias 0.19161f
C2320 XThC.Tn[8] XA.XIR[13].XIC[8].icell.Ien 0.04604f
C2321 XA.XIR[0].XIC[3].icell.Ien Vbias 0.19213f
C2322 XThR.Tn[12] XA.XIR[12].XIC[11].icell.Ien 0.14211f
C2323 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR 0.3367f
C2324 XThC.Tn[4] XThC.Tn[5] 0.31867f
C2325 XThR.XTB2.Y a_n1049_7787# 0.2342f
C2326 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PDM 0.02601f
C2327 XA.XIR[2].XIC_dummy_left.icell.Iout VPWR 0.10954f
C2328 XA.XIR[0].XIC[12].icell.PDM VPWR 0.01451f
C2329 XA.XIR[7].XIC[6].icell.Ien Vbias 0.19161f
C2330 XA.XIR[13].XIC[14].icell.Ien VPWR 0.18835f
C2331 XThC.XTBN.Y Vbias 0.22975f
C2332 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PDM 0.02602f
C2333 XThC.Tn[5] XA.XIR[15].XIC[5].icell.Ien 0.04292f
C2334 XThR.Tn[4] XA.XIR[4].XIC[2].icell.Ien 0.14211f
C2335 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.Ien 0.04854f
C2336 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PDM 0.04035f
C2337 XThC.XTB4.Y XThC.XTB7.Y 0.03475f
C2338 XThR.XTB6.Y XThR.Tn[7] 0.01462f
C2339 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.Ien 0.04854f
C2340 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PDM 0.04035f
C2341 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR 0.0824f
C2342 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.PDM 0.02104f
C2343 XThC.Tn[13] XThR.Tn[7] 0.40739f
C2344 XThC.Tn[6] XA.XIR[11].XIC[6].icell.Ien 0.04604f
C2345 XThC.XTB7.B XThC.Tn[11] 0.03651f
C2346 XThC.Tn[10] XA.XIR[6].XIC[10].icell.Ien 0.04604f
C2347 XA.XIR[6].XIC[14].icell.Ien Iout 0.06801f
C2348 XThC.Tn[10] Vbias 0.81591f
C2349 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.PDM 0.02104f
C2350 XA.XIR[10].XIC[10].icell.Ien VPWR 0.18829f
C2351 XA.XIR[14].XIC[8].icell.Ien Iout 0.06801f
C2352 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.PDM 0.02104f
C2353 XA.XIR[5].XIC[6].icell.PDM Vbias 0.03928f
C2354 XThR.Tn[3] XA.XIR[3].XIC[5].icell.Ien 0.14211f
C2355 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PDM 0.0404f
C2356 a_3773_9615# XThC.Tn[2] 0.01043f
C2357 XA.XIR[13].XIC[0].icell.PDM Vbias 0.03915f
C2358 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.Ien 0.04854f
C2359 XThR.XTB3.Y VPWR 1.07975f
C2360 XA.XIR[12].XIC[5].icell.PDM Vbias 0.03928f
C2361 XThC.Tn[12] XThR.Tn[3] 0.40738f
C2362 XThR.XTB5.A XThR.XTB6.A 1.80461f
C2363 XA.XIR[12].XIC[12].icell.Ien Vbias 0.19161f
C2364 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2365 XThC.Tn[0] VPWR 3.67891f
C2366 XA.XIR[6].XIC[3].icell.PDM VPWR 0.01171f
C2367 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PDM 0.0404f
C2368 XA.XIR[14].XIC[0].icell.PDM VPWR 0.01171f
C2369 XA.XIR[5].XIC[10].icell.PDM VPWR 0.01171f
C2370 XA.XIR[8].XIC[1].icell.Ien Vbias 0.19161f
C2371 XThC.Tn[8] XThR.Tn[5] 0.40738f
C2372 XA.XIR[3].XIC[3].icell.Ien Vbias 0.19161f
C2373 XA.XIR[13].XIC[4].icell.PDM VPWR 0.01171f
C2374 XA.XIR[13].XIC[12].icell.Ien VPWR 0.18829f
C2375 XThC.Tn[14] XA.XIR[8].XIC[14].icell.Ien 0.04604f
C2376 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.02601f
C2377 XA.XIR[15].XIC[9].icell.Ien Vbias 0.15966f
C2378 XA.XIR[12].XIC[9].icell.PDM VPWR 0.01171f
C2379 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.PDM 0.02104f
C2380 XThC.Tn[1] XA.XIR[14].XIC[1].icell.Ien 0.04604f
C2381 XThC.XTB6.A XThC.XTB6.Y 0.10153f
C2382 XThC.XTB2.Y XThC.XTB7.Y 0.0437f
C2383 XA.XIR[9].XIC[2].icell.Ien VPWR 0.18829f
C2384 XA.XIR[4].XIC[12].icell.Ien Vbias 0.19161f
C2385 XA.XIR[3].XIC[1].icell.PDM Vbias 0.03928f
C2386 XA.XIR[8].XIC[3].icell.PDM Vbias 0.03928f
C2387 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.Ien 0.04854f
C2388 XThR.XTB6.A data[5] 0.37233f
C2389 XA.XIR[2].XIC[7].icell.PDM Vbias 0.03928f
C2390 XA.XIR[8].XIC[6].icell.Ien Vbias 0.19161f
C2391 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PDM 0.04035f
C2392 XA.XIR[5].XIC[11].icell.Ien VPWR 0.18829f
C2393 XA.XIR[9].XIC_15.icell.Ien Vbias 0.19195f
C2394 XA.XIR[5].XIC[7].icell.Ien Iout 0.06801f
C2395 XA.XIR[8].XIC[7].icell.PDM VPWR 0.01171f
C2396 XA.XIR[3].XIC[5].icell.PDM VPWR 0.01171f
C2397 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.PDM 0.02104f
C2398 XA.XIR[2].XIC[11].icell.PDM VPWR 0.01171f
C2399 XA.XIR[0].XIC[8].icell.Ien Vbias 0.19213f
C2400 XThC.Tn[14] XThR.Tn[2] 0.40744f
C2401 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.PDM 0.02104f
C2402 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PDM 0.04035f
C2403 XThC.XTB6.A XThC.XTB4.Y 0.04137f
C2404 XA.XIR[12].XIC[6].icell.Ien VPWR 0.18829f
C2405 XThC.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.04605f
C2406 XA.XIR[12].XIC[10].icell.Ien Vbias 0.19161f
C2407 XThR.XTB6.Y a_n997_1579# 0.07626f
C2408 XA.XIR[10].XIC_15.icell.Ien VPWR 0.26829f
C2409 XA.XIR[12].XIC[2].icell.Ien Iout 0.06801f
C2410 XA.XIR[7].XIC[11].icell.Ien Vbias 0.19161f
C2411 XThC.Tn[6] XA.XIR[14].XIC[6].icell.Ien 0.04604f
C2412 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.PDM 0.02104f
C2413 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.PDM 0.02104f
C2414 XThR.Tn[4] XA.XIR[4].XIC[7].icell.Ien 0.14211f
C2415 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.Ien 0.04854f
C2416 XA.XIR[3].XIC[0].icell.Ien Vbias 0.19149f
C2417 XA.XIR[13].XIC[10].icell.Ien VPWR 0.18829f
C2418 XThR.Tn[8] Vbias 1.39526f
C2419 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PDM 0.04035f
C2420 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Iout 0.02485f
C2421 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PDM 0.04035f
C2422 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.PDM 0.02104f
C2423 XThC.Tn[10] XThR.Tn[6] 0.40738f
C2424 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PDM 0.04035f
C2425 XA.XIR[11].XIC[1].icell.Ien Vbias 0.19161f
C2426 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.PDM 0.02104f
C2427 XThC.Tn[12] XThR.Tn[11] 0.40738f
C2428 XA.XIR[10].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2429 XA.XIR[7].XIC[7].icell.PDM Vbias 0.03928f
C2430 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PDM 0.0404f
C2431 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.Ien 0.04854f
C2432 XA.XIR[6].XIC[14].icell.PDM Vbias 0.03928f
C2433 XThC.Tn[2] XThR.Tn[7] 0.40738f
C2434 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PDM 0.04056f
C2435 XA.XIR[15].XIC[5].icell.PDM Vbias 0.03928f
C2436 XThR.Tn[12] XA.XIR[12].XIC[5].icell.Ien 0.14211f
C2437 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2438 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.PDM 0.02104f
C2439 XThR.Tn[3] XA.XIR[3].XIC[10].icell.Ien 0.14211f
C2440 XA.XIR[15].XIC[14].icell.Ien Vbias 0.15966f
C2441 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.PDM 0.02104f
C2442 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.Ien 0.04854f
C2443 XThC.XTB6.Y XThC.Tn[8] 0.02463f
C2444 XThC.Tn[2] XA.XIR[4].XIC[2].icell.Ien 0.04604f
C2445 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PDM 0.04056f
C2446 XA.XIR[9].XIC[3].icell.PDM Vbias 0.03928f
C2447 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.Ien 0.04854f
C2448 XThR.Tn[0] Iout 1.12768f
C2449 XA.XIR[7].XIC[11].icell.PDM VPWR 0.01171f
C2450 XThR.XTB7.Y a_n1319_5317# 0.01283f
C2451 XThR.Tn[2] XA.XIR[2].XIC[5].icell.Ien 0.14211f
C2452 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PDM 0.02601f
C2453 XA.XIR[15].XIC[9].icell.PDM VPWR 0.01512f
C2454 XA.XIR[4].XIC[4].icell.Ien VPWR 0.18829f
C2455 XThC.XTB2.Y XThC.XTB6.A 0.18237f
C2456 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PDM 0.02602f
C2457 XA.XIR[3].XIC[8].icell.Ien Vbias 0.19161f
C2458 XA.XIR[1].XIC[8].icell.PDM Vbias 0.03928f
C2459 XThC.Tn[1] XThR.Tn[3] 0.40738f
C2460 XA.XIR[9].XIC[7].icell.PDM VPWR 0.01171f
C2461 XThC.Tn[10] XThR.Tn[4] 0.40738f
C2462 XThC.XTBN.Y XThC.Tn[13] 0.41509f
C2463 XA.XIR[4].XIC[8].icell.PDM Vbias 0.03928f
C2464 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.Ien 0.04854f
C2465 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.Ien 0.04854f
C2466 XA.XIR[9].XIC[7].icell.Ien VPWR 0.18829f
C2467 XA.XIR[1].XIC[3].icell.Ien Vbias 0.19173f
C2468 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.PDM 0.02104f
C2469 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.Ien 0.04854f
C2470 XThC.XTB4.Y XThC.Tn[8] 0.01307f
C2471 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.PDM 0.02104f
C2472 XA.XIR[9].XIC[3].icell.Ien Iout 0.06801f
C2473 XThR.Tn[9] XA.XIR[9].XIC[3].icell.Ien 0.14211f
C2474 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.PDM 0.02104f
C2475 XA.XIR[12].XIC_15.icell.Ien Vbias 0.19195f
C2476 XThC.Tn[14] XThR.Tn[10] 0.40742f
C2477 XThC.Tn[4] XThR.Tn[0] 0.40763f
C2478 XThC.Tn[6] XThR.Tn[5] 0.40738f
C2479 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PDM 0.02601f
C2480 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PDM 0.04035f
C2481 XA.XIR[8].XIC[11].icell.Ien Vbias 0.19161f
C2482 XA.XIR[1].XIC[12].icell.PDM VPWR 0.01171f
C2483 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.PDM 0.02104f
C2484 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.Ien 0.04854f
C2485 XThC.Tn[7] XA.XIR[0].XIC[7].icell.Ien 0.04658f
C2486 XThC.Tn[11] XThC.Tn[12] 0.12311f
C2487 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.Ien 0.04854f
C2488 XA.XIR[4].XIC[12].icell.PDM VPWR 0.01171f
C2489 XA.XIR[7].XIC[3].icell.Ien VPWR 0.18829f
C2490 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PDM 0.04035f
C2491 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.Ien 0.04854f
C2492 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.Ien 0.04854f
C2493 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.PDM 0.02104f
C2494 XThC.XTB7.B VPWR 1.33508f
C2495 XA.XIR[5].XIC[12].icell.Ien Iout 0.06801f
C2496 XA.XIR[13].XIC_15.icell.Ien VPWR 0.26829f
C2497 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.Ien 0.04854f
C2498 XA.XIR[15].XIC[12].icell.Ien Vbias 0.15966f
C2499 XA.XIR[0].XIC[13].icell.Ien Vbias 0.19213f
C2500 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.Ien 0.04854f
C2501 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PDM 0.04035f
C2502 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PDM 0.04035f
C2503 XThC.XTBN.A XThC.XTB5.Y 0.10854f
C2504 XThC.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.04657f
C2505 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.PDM 0.02104f
C2506 XThR.Tn[7] XA.XIR[7].XIC[0].icell.Ien 0.14211f
C2507 XA.XIR[12].XIC[7].icell.Ien Iout 0.06801f
C2508 XThR.XTBN.A XThR.Tn[8] 0.1369f
C2509 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PDM 0.02601f
C2510 VPWR bias[0] 2.10172f
C2511 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PDM 0.04035f
C2512 XThC.Tn[3] XThR.Tn[2] 0.40741f
C2513 XA.XIR[14].XIC[1].icell.Ien Vbias 0.19161f
C2514 XThR.Tn[4] XA.XIR[4].XIC[12].icell.Ien 0.14211f
C2515 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.0404f
C2516 XThR.Tn[0] XA.XIR[0].XIC[4].icell.Ien 0.14211f
C2517 XA.XIR[0].XIC_15.icell.PUM VPWR 0.01577f
C2518 XThC.XTB7.Y a_6243_9615# 0.27822f
C2519 XA.XIR[13].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2520 XThC.Tn[12] XThR.Tn[14] 0.40738f
C2521 XThR.Tn[10] XA.XIR[10].XIC[3].icell.Ien 0.14211f
C2522 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PDM 0.0404f
C2523 XA.XIR[10].XIC[2].icell.PDM Vbias 0.03928f
C2524 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PDM 0.02601f
C2525 XThC.XTBN.A XThC.XTBN.Y 0.77125f
C2526 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PDM 0.04035f
C2527 XThC.Tn[12] XA.XIR[10].XIC[12].icell.Ien 0.04604f
C2528 XA.XIR[6].XIC[3].icell.Ien Vbias 0.19161f
C2529 XThR.XTB7.B data[6] 0.07481f
C2530 XThR.Tn[7] XA.XIR[7].XIC[5].icell.Ien 0.14211f
C2531 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.PDM 0.02104f
C2532 XA.XIR[15].XIC[1].icell.Ien VPWR 0.31713f
C2533 XA.XIR[5].XIC_dummy_left.icell.Iout VPWR 0.11011f
C2534 XThC.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.04604f
C2535 XA.XIR[1].XIC[0].icell.Ien Iout 0.06795f
C2536 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.Ien 0.04854f
C2537 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.Ien 0.04854f
C2538 XA.XIR[11].XIC[2].icell.PDM VPWR 0.01171f
C2539 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.Ien 0.04854f
C2540 XA.XIR[4].XIC[0].icell.Ien Iout 0.06795f
C2541 XA.XIR[10].XIC[6].icell.PDM VPWR 0.01171f
C2542 XThR.Tn[1] Iout 1.12765f
C2543 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PDM 0.02602f
C2544 XThR.Tn[3] XA.XIR[3].XIC_15.icell.Ien 0.13564f
C2545 XThC.XTBN.A XThC.Tn[10] 0.12208f
C2546 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.PDM 0.02104f
C2547 XThR.Tn[12] Iout 1.12762f
C2548 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PDM 0.02601f
C2549 XThC.Tn[1] XThR.Tn[11] 0.40738f
C2550 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout 0.06446f
C2551 XA.XIR[2].XIC[1].icell.Ien Vbias 0.19161f
C2552 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.Ien 0.04854f
C2553 XA.XIR[0].XIC[10].icell.PDM Vbias 0.03945f
C2554 XA.XIR[15].XIC[6].icell.Ien VPWR 0.31713f
C2555 XA.XIR[11].XIC[2].icell.Ien Vbias 0.19161f
C2556 XThC.Tn[7] XA.XIR[3].XIC[7].icell.Ien 0.04604f
C2557 XA.XIR[15].XIC[10].icell.Ien Vbias 0.15966f
C2558 XThR.Tn[2] XA.XIR[2].XIC[10].icell.Ien 0.14211f
C2559 XA.XIR[15].XIC[2].icell.Ien Iout 0.07192f
C2560 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PDM 0.0279f
C2561 XThC.XTB7.A Vbias 0.0148f
C2562 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.PDM 0.02104f
C2563 XThC.XTB3.Y XThC.XTB5.Y 0.04438f
C2564 XA.XIR[4].XIC[9].icell.Ien VPWR 0.18829f
C2565 XA.XIR[10].XIC[4].icell.Ien Vbias 0.19161f
C2566 XThC.Tn[14] XA.XIR[2].XIC[14].icell.Ien 0.04605f
C2567 XA.XIR[0].XIC[0].icell.Ien VPWR 0.18776f
C2568 XA.XIR[4].XIC[5].icell.Ien Iout 0.06801f
C2569 XThC.Tn[0] XA.XIR[10].XIC[0].icell.Ien 0.04604f
C2570 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.PDM 0.02104f
C2571 XA.XIR[8].XIC[3].icell.Ien VPWR 0.18829f
C2572 XThC.XTB6.Y XThC.Tn[6] 0.01038f
C2573 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.Ien 0.04854f
C2574 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.Ien 0.04854f
C2575 XA.XIR[3].XIC[13].icell.Ien Vbias 0.19161f
C2576 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.PDM 0.02104f
C2577 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PDM 0.02601f
C2578 XThC.Tn[14] XThR.Tn[13] 0.40742f
C2579 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PDM 0.02601f
C2580 XThC.Tn[4] XThR.Tn[1] 0.40744f
C2581 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.Ien 0.04854f
C2582 XA.XIR[0].XIC[14].icell.PDM VPWR 0.01141f
C2583 XA.XIR[2].XIC[6].icell.Ien Vbias 0.19161f
C2584 XThC.Tn[8] Iout 0.22393f
C2585 XThC.Tn[8] XThR.Tn[9] 0.40738f
C2586 XA.XIR[9].XIC[12].icell.Ien VPWR 0.18829f
C2587 XThR.XTB6.Y XThR.Tn[8] 0.02461f
C2588 XA.XIR[1].XIC[8].icell.Ien Vbias 0.19173f
C2589 XThC.Tn[4] XThR.Tn[12] 0.40738f
C2590 XA.XIR[9].XIC[8].icell.Ien Iout 0.06801f
C2591 XThC.Tn[13] XThR.Tn[8] 0.40739f
C2592 XThR.Tn[9] XA.XIR[9].XIC[8].icell.Ien 0.14211f
C2593 XThC.XTB3.Y XThC.XTBN.Y 0.17246f
C2594 XA.XIR[0].XIC[5].icell.Ien VPWR 0.18797f
C2595 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.04035f
C2596 XThR.XTBN.A a_n997_3755# 0.01939f
C2597 XThR.XTB2.Y XThR.XTBN.A 0.04716f
C2598 XA.XIR[3].XIC_15.icell.PUM VPWR 0.01655f
C2599 XThC.XTBN.Y XThC.Tn[2] 0.49723f
C2600 XThR.XTB7.A XThR.Tn[5] 0.02751f
C2601 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2602 XA.XIR[7].XIC[8].icell.Ien VPWR 0.18829f
C2603 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.PDM 0.02104f
C2604 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.Ien 0.04854f
C2605 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.Ien 0.04854f
C2606 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PDM 0.02601f
C2607 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PDM 0.0404f
C2608 XA.XIR[7].XIC[4].icell.Ien Iout 0.06801f
C2609 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PDM 0.04035f
C2610 XThC.Tn[3] XThR.Tn[10] 0.40738f
C2611 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PDM 0.02601f
C2612 XThC.XTB3.Y XThC.Tn[10] 0.29566f
C2613 XA.XIR[6].XIC[1].icell.PDM Vbias 0.03928f
C2614 XThC.Tn[5] XA.XIR[10].XIC[5].icell.Ien 0.04604f
C2615 XA.XIR[5].XIC[8].icell.PDM Vbias 0.03928f
C2616 XA.XIR[13].XIC[2].icell.PDM Vbias 0.03928f
C2617 a_n1049_8581# VPWR 0.71708f
C2618 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.PDM 0.02104f
C2619 XThR.Tn[3] Vbias 1.39527f
C2620 XThR.Tn[11] XA.XIR[11].XIC[4].icell.Ien 0.14211f
C2621 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PDM 0.04035f
C2622 XThC.XTB1.Y XThC.XTB5.Y 0.05054f
C2623 XA.XIR[12].XIC[7].icell.PDM Vbias 0.03928f
C2624 XThC.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.04604f
C2625 XA.XIR[10].XIC[0].icell.Ien VPWR 0.18829f
C2626 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout 0.06446f
C2627 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.PDM 0.02104f
C2628 XThC.Tn[8] XA.XIR[4].XIC[8].icell.Ien 0.04604f
C2629 XThR.XTB1.Y XThR.XTB5.Y 0.05054f
C2630 XA.XIR[6].XIC[5].icell.PDM VPWR 0.01171f
C2631 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.Ien 0.04854f
C2632 XThR.Tn[0] XA.XIR[0].XIC[9].icell.Ien 0.14211f
C2633 XThC.Tn[10] XA.XIR[14].XIC[10].icell.Ien 0.04604f
C2634 XThR.Tn[10] XA.XIR[10].XIC[8].icell.Ien 0.14211f
C2635 XThR.Tn[6] XA.XIR[6].XIC[3].icell.Ien 0.14211f
C2636 XA.XIR[5].XIC[12].icell.PDM VPWR 0.01171f
C2637 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.PDM 0.02104f
C2638 XA.XIR[14].XIC[2].icell.PDM VPWR 0.01171f
C2639 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.PDM 0.02104f
C2640 XThC.Tn[4] XA.XIR[7].XIC[4].icell.Ien 0.04604f
C2641 XA.XIR[15].XIC_15.icell.Ien Vbias 0.15966f
C2642 XA.XIR[13].XIC[6].icell.PDM VPWR 0.01171f
C2643 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.PDM 0.02104f
C2644 XA.XIR[6].XIC[8].icell.Ien Vbias 0.19161f
C2645 XThR.Tn[7] XA.XIR[7].XIC[10].icell.Ien 0.14211f
C2646 XThC.Tn[1] XA.XIR[5].XIC[1].icell.Ien 0.04604f
C2647 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.Ien 0.04854f
C2648 XThC.Tn[1] XThR.Tn[14] 0.40738f
C2649 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PDM 0.02601f
C2650 XThC.XTB1.Y XThC.XTBN.Y 0.1979f
C2651 XA.XIR[12].XIC_dummy_left.icell.Ien XThR.Tn[12] 0.01244f
C2652 XA.XIR[8].XIC[5].icell.PDM Vbias 0.03928f
C2653 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.PDM 0.02104f
C2654 XA.XIR[3].XIC[3].icell.PDM Vbias 0.03928f
C2655 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PDM 0.02803f
C2656 XThR.XTB2.Y a_n1049_7493# 0.02133f
C2657 XA.XIR[14].XIC[2].icell.Ien Vbias 0.19161f
C2658 XA.XIR[2].XIC[9].icell.PDM Vbias 0.03928f
C2659 XA.XIR[13].XIC[4].icell.Ien Vbias 0.19161f
C2660 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.PDM 0.02104f
C2661 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Iout 0.01728f
C2662 XA.XIR[3].XIC[5].icell.Ien VPWR 0.18829f
C2663 XA.XIR[12].XIC_dummy_left.icell.Iout VPWR 0.10997f
C2664 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.04035f
C2665 XThC.Tn[0] XA.XIR[13].XIC[0].icell.Ien 0.04604f
C2666 XThR.XTB2.Y XThR.XTB6.Y 0.04959f
C2667 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PDM 0.02601f
C2668 XA.XIR[11].XIC[7].icell.Ien Vbias 0.19161f
C2669 XThC.Tn[6] XA.XIR[9].XIC[6].icell.Ien 0.04604f
C2670 XThR.Tn[2] XA.XIR[2].XIC_15.icell.Ien 0.13564f
C2671 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.PDM 0.02104f
C2672 XThC.Tn[12] VPWR 4.5561f
C2673 XA.XIR[15].XIC[7].icell.Ien Iout 0.07192f
C2674 XThC.Tn[13] XA.XIR[0].XIC[13].icell.Ien 0.04662f
C2675 XA.XIR[4].XIC[14].icell.Ien VPWR 0.18835f
C2676 XA.XIR[8].XIC[9].icell.PDM VPWR 0.01171f
C2677 XA.XIR[3].XIC[7].icell.PDM VPWR 0.01171f
C2678 XA.XIR[10].XIC[9].icell.Ien Vbias 0.19161f
C2679 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Iout 0.0203f
C2680 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.Ien 0.04854f
C2681 XThC.XTBN.A a_7651_9569# 0.02087f
C2682 XA.XIR[4].XIC[10].icell.Ien Iout 0.06801f
C2683 XA.XIR[2].XIC[13].icell.PDM VPWR 0.01171f
C2684 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PDM 0.04035f
C2685 XThC.Tn[7] XA.XIR[1].XIC[7].icell.Ien 0.04606f
C2686 XA.XIR[8].XIC[8].icell.Ien VPWR 0.18829f
C2687 XA.XIR[0].XIC[1].icell.Ien Iout 0.0675f
C2688 XThR.XTB6.Y a_n1049_5611# 0.26831f
C2689 XA.XIR[8].XIC[4].icell.Ien Iout 0.06801f
C2690 XA.XIR[10].XIC_15.icell.PDM VPWR 0.07527f
C2691 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.Ien 0.04854f
C2692 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.Ien 0.04854f
C2693 XA.XIR[2].XIC[11].icell.Ien Vbias 0.19161f
C2694 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.PDM 0.02104f
C2695 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR 0.39107f
C2696 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PDM 0.04035f
C2697 XA.XIR[1].XIC[13].icell.Ien Vbias 0.19173f
C2698 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2699 XA.XIR[9].XIC[13].icell.Ien Iout 0.06801f
C2700 XA.XIR[0].XIC[10].icell.Ien VPWR 0.18776f
C2701 XThR.Tn[9] XA.XIR[9].XIC[13].icell.Ien 0.14211f
C2702 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.Ien 0.04854f
C2703 XThC.Tn[3] XThR.Tn[13] 0.40738f
C2704 bias[1] Vbias 0.05009f
C2705 XA.XIR[0].XIC[6].icell.Ien Iout 0.0675f
C2706 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PDM 0.04035f
C2707 XThC.Tn[5] XA.XIR[13].XIC[5].icell.Ien 0.04604f
C2708 XA.XIR[12].XIC[0].icell.Ien Vbias 0.19149f
C2709 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PDM 0.04035f
C2710 XA.XIR[7].XIC[13].icell.Ien VPWR 0.18829f
C2711 XThC.Tn[6] Iout 0.22423f
C2712 XThR.Tn[11] Vbias 1.39532f
C2713 XThC.Tn[6] XThR.Tn[9] 0.40738f
C2714 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PDM 0.02601f
C2715 XThR.Tn[13] XA.XIR[13].XIC[3].icell.Ien 0.14211f
C2716 XThC.Tn[2] XThR.Tn[8] 0.40738f
C2717 XA.XIR[7].XIC[9].icell.PDM Vbias 0.03928f
C2718 XA.XIR[7].XIC[9].icell.Ien Iout 0.06801f
C2719 XA.XIR[1].XIC_15.icell.PUM VPWR 0.01655f
C2720 XThC.Tn[4] XA.XIR[8].XIC[4].icell.Ien 0.04604f
C2721 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.Ien 0.04854f
C2722 XA.XIR[15].XIC[7].icell.PDM Vbias 0.03928f
C2723 XA.XIR[13].XIC[0].icell.Ien VPWR 0.18829f
C2724 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.Ien 0.04854f
C2725 XThC.XTBN.Y a_2979_9615# 0.0607f
C2726 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.Ien 0.04854f
C2727 XThR.XTB7.Y XThR.XTBN.A 1.11559f
C2728 XThR.XTBN.A data[4] 0.02581f
C2729 XThR.Tn[11] XA.XIR[11].XIC[9].icell.Ien 0.14211f
C2730 XA.XIR[2].XIC[0].icell.Ien Iout 0.06795f
C2731 XA.XIR[9].XIC[5].icell.PDM Vbias 0.03928f
C2732 XThR.XTB5.A XThR.XTB7.A 0.07862f
C2733 data[2] data[3] 0.04128f
C2734 XA.XIR[7].XIC[13].icell.PDM VPWR 0.01171f
C2735 XThR.XTB7.Y XThR.Tn[6] 0.21438f
C2736 a_9827_9569# XThC.Tn[12] 0.20217f
C2737 XThC.Tn[0] XThC.Tn[1] 0.88262f
C2738 XThC.XTB6.A data[0] 0.48493f
C2739 XThC.Tn[7] XA.XIR[6].XIC[7].icell.Ien 0.04604f
C2740 XA.XIR[10].XIC[1].icell.Ien Iout 0.06801f
C2741 XThR.Tn[0] XA.XIR[0].XIC[14].icell.Ien 0.144f
C2742 XThC.Tn[13] XA.XIR[3].XIC[13].icell.Ien 0.04604f
C2743 XThR.Tn[6] XA.XIR[6].XIC[8].icell.Ien 0.14211f
C2744 a_n1049_7787# VPWR 0.72173f
C2745 XA.XIR[1].XIC[10].icell.PDM Vbias 0.03928f
C2746 XA.XIR[6].XIC[13].icell.Ien Vbias 0.19161f
C2747 XThR.Tn[7] XA.XIR[7].XIC_15.icell.Ien 0.13564f
C2748 XA.XIR[9].XIC[9].icell.PDM VPWR 0.01171f
C2749 XA.XIR[10].XIC[14].icell.Ien Vbias 0.19161f
C2750 XA.XIR[0].XIC[1].icell.PDM VPWR 0.01132f
C2751 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PDM 0.02602f
C2752 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.Ien 0.04854f
C2753 XA.XIR[4].XIC[10].icell.PDM Vbias 0.03928f
C2754 XThC.Tn[0] XA.XIR[6].XIC[0].icell.Ien 0.04604f
C2755 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.Ien 0.04854f
C2756 XThC.Tn[14] XThR.Tn[7] 0.40742f
C2757 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PDM 0.02601f
C2758 XThC.XTB5.A a_7331_10587# 0.01243f
C2759 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.Ien 0.04854f
C2760 XA.XIR[14].XIC[7].icell.Ien Vbias 0.19161f
C2761 XThR.XTB7.A data[5] 0.06538f
C2762 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.Ien 0.04854f
C2763 XA.XIR[13].XIC[9].icell.Ien Vbias 0.19161f
C2764 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PDM 0.04035f
C2765 XThR.XTBN.Y XThR.Tn[5] 0.59911f
C2766 XThC.Tn[11] Vbias 0.82596f
C2767 XA.XIR[11].XIC[13].icell.Ien Iout 0.06801f
C2768 XA.XIR[1].XIC[14].icell.PDM VPWR 0.0118f
C2769 XA.XIR[3].XIC[10].icell.Ien VPWR 0.18829f
C2770 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout 0.06446f
C2771 XA.XIR[6].XIC_15.icell.PUM VPWR 0.01655f
C2772 XA.XIR[10].XIC[14].icell.PDM VPWR 0.0118f
C2773 XThR.XTBN.A a_n997_2667# 0.01679f
C2774 XThR.Tn[3] XThR.Tn[4] 0.1175f
C2775 XA.XIR[3].XIC[6].icell.Ien Iout 0.06801f
C2776 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PDM 0.02601f
C2777 XA.XIR[4].XIC[14].icell.PDM VPWR 0.0118f
C2778 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR 0.01493f
C2779 XA.XIR[2].XIC[3].icell.Ien VPWR 0.18829f
C2780 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PDM 0.04035f
C2781 XA.XIR[1].XIC[5].icell.Ien VPWR 0.18829f
C2782 XA.XIR[13].XIC_15.icell.PDM VPWR 0.07527f
C2783 XA.XIR[4].XIC_15.icell.Ien Iout 0.0694f
C2784 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PDM 0.0404f
C2785 XA.XIR[8].XIC[13].icell.Ien VPWR 0.18829f
C2786 XThC.Tn[13] XThR.Tn[3] 0.40739f
C2787 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.Ien 0.04854f
C2788 XThC.XTB7.A XThC.XTBN.A 0.197f
C2789 XA.XIR[8].XIC[9].icell.Ien Iout 0.06801f
C2790 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PDM 0.02602f
C2791 XThC.Tn[1] VPWR 3.60376f
C2792 XThC.XTB1.Y a_7651_9569# 0.06353f
C2793 XA.XIR[5].XIC[1].icell.Ien Vbias 0.19161f
C2794 XThR.XTB6.Y XThR.XTB7.Y 2.05133f
C2795 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PDM 0.02601f
C2796 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PDM 0.04035f
C2797 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.Ien 0.04854f
C2798 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PDM 0.02601f
C2799 XThR.Tn[14] Vbias 1.39537f
C2800 XThC.Tn[9] XThR.Tn[5] 0.40738f
C2801 XThR.XTBN.A XThR.Tn[11] 0.11968f
C2802 XA.XIR[0].XIC_15.icell.Ien VPWR 0.26622f
C2803 XA.XIR[11].XIC[0].icell.PDM Vbias 0.03915f
C2804 XThC.Tn[14] XA.XIR[5].XIC[14].icell.Ien 0.04604f
C2805 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.04035f
C2806 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PDM 0.02801f
C2807 XA.XIR[10].XIC[4].icell.PDM Vbias 0.03928f
C2808 XThR.Tn[14] XA.XIR[14].XIC[4].icell.Ien 0.14211f
C2809 XThR.Tn[1] XA.XIR[1].XIC[4].icell.Ien 0.14211f
C2810 XThR.Tn[11] XA.XIR[11].XIC[14].icell.Ien 0.144f
C2811 XA.XIR[0].XIC[11].icell.Ien Iout 0.0675f
C2812 XA.XIR[10].XIC[12].icell.Ien Vbias 0.19161f
C2813 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PDM 0.02601f
C2814 XA.XIR[4].XIC_dummy_right.icell.Iout Iout 0.01732f
C2815 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout 0.06446f
C2816 XA.XIR[4].XIC_dummy_right.icell.Iout XA.XIR[5].XIC_dummy_right.icell.Iout 0.04047f
C2817 XA.XIR[6].XIC[0].icell.Ien VPWR 0.18829f
C2818 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PDM 0.04035f
C2819 XThC.Tn[8] data[0] 0.01744f
C2820 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.Ien 0.04854f
C2821 XThR.XTB5.A XThR.XTB7.B 0.30355f
C2822 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PDM 0.02601f
C2823 XA.XIR[15].XIC_dummy_left.icell.Iout VPWR 0.24997f
C2824 XThR.Tn[13] XA.XIR[13].XIC[8].icell.Ien 0.14211f
C2825 XThC.Tn[10] XA.XIR[7].XIC[10].icell.Ien 0.04604f
C2826 a_6243_9615# XThC.Tn[6] 0.26385f
C2827 XA.XIR[7].XIC[14].icell.Ien Iout 0.06801f
C2828 XA.XIR[5].XIC[6].icell.Ien Vbias 0.19161f
C2829 XA.XIR[11].XIC[4].icell.PDM VPWR 0.01171f
C2830 XA.XIR[11].XIC[11].icell.Ien Iout 0.06801f
C2831 XA.XIR[10].XIC[8].icell.PDM VPWR 0.01171f
C2832 XA.XIR[0].XIC_dummy_right.icell.Iout VPWR 0.12361f
C2833 XA.XIR[13].XIC[1].icell.Ien Iout 0.06801f
C2834 XA.XIR[11].XIC_dummy_right.icell.Iout XA.XIR[12].XIC_dummy_right.icell.Iout 0.04047f
C2835 XThR.XTB6.A XThR.XTB5.Y 0.01866f
C2836 XA.XIR[6].XIC[5].icell.Ien VPWR 0.18829f
C2837 XA.XIR[0].XIC[12].icell.PDM Vbias 0.03945f
C2838 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PDM 0.02602f
C2839 XA.XIR[13].XIC[14].icell.Ien Vbias 0.19161f
C2840 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PDM 0.02601f
C2841 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PDM 0.02601f
C2842 XThC.Tn[12] XA.XIR[9].XIC[12].icell.Ien 0.04604f
C2843 XA.XIR[2].XIC[0].icell.PDM VPWR 0.01171f
C2844 XThR.Tn[6] XA.XIR[6].XIC[13].icell.Ien 0.14211f
C2845 XThC.XTB7.A XThC.XTB3.Y 0.57441f
C2846 XThC.XTB5.A XThC.XTBN.A 0.06305f
C2847 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PDM 0.02601f
C2848 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PDM 0.02601f
C2849 XThC.Tn[2] XA.XIR[11].XIC[2].icell.Ien 0.04604f
C2850 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR 0.01669f
C2851 XA.XIR[10].XIC[13].icell.PDM VPWR 0.01171f
C2852 XThC.XTB7.A XThC.Tn[2] 0.1255f
C2853 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.Ien 0.04854f
C2854 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR 0.08055f
C2855 XA.XIR[14].XIC[13].icell.Ien Iout 0.06801f
C2856 XA.XIR[11].XIC[4].icell.Ien VPWR 0.18829f
C2857 XThC.Tn[13] XA.XIR[1].XIC[13].icell.Ien 0.04606f
C2858 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PDM 0.04042f
C2859 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PDM 0.02601f
C2860 XA.XIR[13].XIC[14].icell.PDM VPWR 0.0118f
C2861 XA.XIR[10].XIC[6].icell.Ien VPWR 0.18829f
C2862 XThC.Tn[11] XThR.Tn[6] 0.40738f
C2863 XThR.Tn[11] XA.XIR[11].XIC[12].icell.Ien 0.14211f
C2864 XA.XIR[10].XIC[10].icell.Ien Vbias 0.19161f
C2865 XA.XIR[1].XIC[1].icell.Ien Iout 0.06801f
C2866 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.Ien 0.04854f
C2867 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.Ien 0.04854f
C2868 XA.XIR[10].XIC[2].icell.Ien Iout 0.06801f
C2869 XThR.XTB6.Y XThR.Tn[11] 0.02465f
C2870 XA.XIR[3].XIC_15.icell.Ien VPWR 0.26829f
C2871 XThC.Tn[13] XThR.Tn[11] 0.40739f
C2872 XA.XIR[3].XIC[11].icell.Ien Iout 0.06801f
C2873 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR 0.39039f
C2874 XThR.XTB1.Y XThR.XTB6.A 0.01609f
C2875 XA.XIR[2].XIC[8].icell.Ien VPWR 0.18829f
C2876 XThC.Tn[3] XThR.Tn[7] 0.40738f
C2877 XA.XIR[1].XIC[10].icell.Ien VPWR 0.18829f
C2878 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR 0.38912f
C2879 XA.XIR[2].XIC[4].icell.Ien Iout 0.06801f
C2880 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Iout 0.01758f
C2881 XThR.Tn[8] XA.XIR[8].XIC[5].icell.Ien 0.14211f
C2882 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PDM 0.04035f
C2883 XThC.Tn[0] Vbias 0.27573f
C2884 XThC.XTB6.Y XThC.Tn[9] 0.0246f
C2885 XA.XIR[1].XIC[6].icell.Ien Iout 0.06801f
C2886 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PDM 0.02601f
C2887 XA.XIR[6].XIC[3].icell.PDM Vbias 0.03928f
C2888 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.PDM 0.02104f
C2889 XThR.XTB1.Y XThR.Tn[0] 0.1837f
C2890 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PDM 0.02803f
C2891 XThC.Tn[10] XA.XIR[8].XIC[10].icell.Ien 0.04604f
C2892 XA.XIR[5].XIC[10].icell.PDM Vbias 0.03928f
C2893 XA.XIR[14].XIC[0].icell.PDM Vbias 0.03915f
C2894 XA.XIR[8].XIC[14].icell.Ien Iout 0.06801f
C2895 XThC.Tn[14] XA.XIR[12].XIC[14].icell.Ien 0.04604f
C2896 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PDM 0.02601f
C2897 XA.XIR[13].XIC[4].icell.PDM Vbias 0.03928f
C2898 XA.XIR[3].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2899 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.Ien 0.04854f
C2900 XA.XIR[13].XIC[12].icell.Ien Vbias 0.19161f
C2901 XThR.Tn[5] XA.XIR[5].XIC[4].icell.Ien 0.14211f
C2902 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.04035f
C2903 XA.XIR[12].XIC[9].icell.PDM Vbias 0.03928f
C2904 XThR.XTB7.B XThR.Tn[9] 0.0565f
C2905 XA.XIR[7].XIC[0].icell.PDM VPWR 0.01171f
C2906 XThC.XTB1.Y XThC.XTB7.A 0.48957f
C2907 XThC.XTB5.A XThC.XTB3.Y 0.01156f
C2908 XA.XIR[9].XIC[2].icell.Ien Vbias 0.19161f
C2909 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PDM 0.02601f
C2910 XA.XIR[6].XIC[7].icell.PDM VPWR 0.01171f
C2911 XThC.Tn[2] XThR.Tn[3] 0.40738f
C2912 XThR.Tn[14] XA.XIR[14].XIC[9].icell.Ien 0.14211f
C2913 XA.XIR[14].XIC[4].icell.PDM VPWR 0.01171f
C2914 XThC.XTBN.Y XThC.Tn[14] 0.42645f
C2915 XThR.Tn[1] XA.XIR[1].XIC[9].icell.Ien 0.14211f
C2916 XA.XIR[5].XIC[14].icell.PDM VPWR 0.0118f
C2917 XThC.Tn[13] XA.XIR[6].XIC[13].icell.Ien 0.04604f
C2918 XThC.Tn[11] XThR.Tn[4] 0.40738f
C2919 XThC.Tn[4] XA.XIR[2].XIC[4].icell.Ien 0.04605f
C2920 XA.XIR[14].XIC[11].icell.Ien Iout 0.06801f
C2921 XThR.XTB5.A XThR.XTB4.Y 0.02767f
C2922 XA.XIR[13].XIC[8].icell.PDM VPWR 0.01171f
C2923 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.PDM 0.02104f
C2924 XThC.XTB4.Y XThC.Tn[9] 0.01318f
C2925 XThC.Tn[1] XA.XIR[15].XIC[1].icell.Ien 0.04292f
C2926 XThC.XTB7.Y a_10051_9569# 0.013f
C2927 XA.XIR[6].XIC[1].icell.Ien Iout 0.06801f
C2928 XThR.Tn[11] XA.XIR[11].XIC[10].icell.Ien 0.14211f
C2929 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.PDM 0.02104f
C2930 XThC.Tn[5] XThR.Tn[0] 0.40765f
C2931 XA.XIR[5].XIC[11].icell.Ien Vbias 0.19161f
C2932 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8] 0.14211f
C2933 XThC.Tn[7] XThR.Tn[5] 0.40738f
C2934 XA.XIR[8].XIC[7].icell.PDM Vbias 0.03928f
C2935 XThR.Tn[2] Iout 1.12764f
C2936 XA.XIR[3].XIC[5].icell.PDM Vbias 0.03928f
C2937 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2938 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.Ien 0.04854f
C2939 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PDM 0.02601f
C2940 XA.XIR[2].XIC[11].icell.PDM Vbias 0.03928f
C2941 XA.XIR[10].XIC[12].icell.PDM VPWR 0.01171f
C2942 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PDM 0.02601f
C2943 XA.XIR[1].XIC[1].icell.PDM VPWR 0.01171f
C2944 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.Ien 0.04854f
C2945 XThC.Tn[2] XA.XIR[14].XIC[2].icell.Ien 0.04604f
C2946 XA.XIR[6].XIC[10].icell.Ien VPWR 0.18829f
C2947 XA.XIR[12].XIC[6].icell.Ien Vbias 0.19161f
C2948 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11] 0.14211f
C2949 XA.XIR[10].XIC_15.icell.Ien Vbias 0.19195f
C2950 XA.XIR[6].XIC[6].icell.Ien Iout 0.06801f
C2951 VPWR Vbias 98.23621f
C2952 XA.XIR[13].XIC[13].icell.PDM VPWR 0.01171f
C2953 XA.XIR[4].XIC[1].icell.PDM VPWR 0.01171f
C2954 XA.XIR[3].XIC[9].icell.PDM VPWR 0.01171f
C2955 XA.XIR[14].XIC[4].icell.Ien VPWR 0.18883f
C2956 XA.XIR[8].XIC[11].icell.PDM VPWR 0.01171f
C2957 XThR.XTB5.Y XThR.Tn[12] 0.32095f
C2958 XThC.XTBN.A a_8739_9569# 0.01719f
C2959 XA.XIR[2].XIC_15.icell.PDM VPWR 0.07527f
C2960 XA.XIR[13].XIC[6].icell.Ien VPWR 0.18829f
C2961 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PDM 0.0404f
C2962 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PDM 0.04035f
C2963 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.PDM 0.02104f
C2964 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout 0.06446f
C2965 XA.XIR[0].XIC_dummy_left.icell.Iout Iout 0.03553f
C2966 XA.XIR[13].XIC[10].icell.Ien Vbias 0.19161f
C2967 XA.XIR[11].XIC_15.icell.PUM VPWR 0.01655f
C2968 XA.XIR[13].XIC[2].icell.Ien Iout 0.06801f
C2969 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2970 XThC.Tn[4] XThR.Tn[2] 0.40741f
C2971 XThC.XTB5.A XThC.XTB1.Y 0.1098f
C2972 XA.XIR[11].XIC[9].icell.Ien VPWR 0.18829f
C2973 XThC.Tn[13] XThR.Tn[14] 0.40739f
C2974 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2975 XA.XIR[11].XIC[5].icell.Ien Iout 0.06801f
C2976 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.PDM 0.02104f
C2977 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.PDM 0.02104f
C2978 XThR.XTB3.Y XThR.XTBN.A 0.03907f
C2979 XA.XIR[10].XIC[7].icell.Ien Iout 0.06801f
C2980 a_7875_9569# XThC.Tn[9] 0.19271f
C2981 XThC.XTB2.Y XThC.Tn[9] 0.292f
C2982 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PDM 0.0404f
C2983 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.PDM 0.02104f
C2984 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Iout 0.01728f
C2985 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.Ien 0.04854f
C2986 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PDM 0.04035f
C2987 XA.XIR[2].XIC[13].icell.Ien VPWR 0.18829f
C2988 XThR.XTBN.Y XThR.Tn[9] 0.48067f
C2989 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PDM 0.02601f
C2990 XThC.Tn[0] XThR.Tn[6] 0.40736f
C2991 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2992 XA.XIR[2].XIC[9].icell.Ien Iout 0.06801f
C2993 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.PDM 0.02104f
C2994 XA.XIR[1].XIC_15.icell.Ien VPWR 0.26829f
C2995 XThR.Tn[8] XA.XIR[8].XIC[10].icell.Ien 0.14211f
C2996 XThC.XTBN.A XThC.Tn[11] 0.11997f
C2997 XThR.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.144f
C2998 XA.XIR[7].XIC[11].icell.PDM Vbias 0.03928f
C2999 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.Ien 0.04854f
C3000 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PDM 0.02602f
C3001 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.PDM 0.02104f
C3002 XA.XIR[1].XIC[11].icell.Ien Iout 0.06801f
C3003 XA.XIR[15].XIC[9].icell.PDM Vbias 0.03928f
C3004 XThC.Tn[2] XThR.Tn[11] 0.40738f
C3005 XA.XIR[4].XIC[4].icell.Ien Vbias 0.19161f
C3006 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR 0.35555f
C3007 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PDM 0.02601f
C3008 XThC.XTBN.Y a_4067_9615# 0.08456f
C3009 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.PDM 0.02104f
C3010 XThR.Tn[11] XA.XIR[11].XIC_15.icell.Ien 0.13564f
C3011 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.Ien 0.04854f
C3012 XA.XIR[9].XIC[7].icell.PDM Vbias 0.03928f
C3013 XThR.Tn[5] XA.XIR[5].XIC[9].icell.Ien 0.14211f
C3014 XThR.XTB4.Y XThR.Tn[9] 0.01318f
C3015 XA.XIR[7].XIC_15.icell.PDM VPWR 0.07527f
C3016 XA.XIR[5].XIC[3].icell.Ien VPWR 0.18829f
C3017 XThC.XTB3.Y a_8739_9569# 0.07285f
C3018 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.Ien 0.04854f
C3019 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PDM 0.02601f
C3020 XA.XIR[9].XIC[7].icell.Ien Vbias 0.19161f
C3021 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.Ien 0.04854f
C3022 XThC.XTB6.Y XThC.Tn[7] 0.01474f
C3023 XThR.Tn[10] Iout 1.12758f
C3024 XThR.Tn[9] XThR.Tn[10] 0.12586f
C3025 XA.XIR[1].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3026 XThC.Tn[3] XA.XIR[0].XIC[3].icell.Ien 0.04658f
C3027 XThC.Tn[5] XThR.Tn[1] 0.40744f
C3028 XThR.Tn[1] XA.XIR[1].XIC[14].icell.Ien 0.144f
C3029 XA.XIR[10].XIC[11].icell.PDM VPWR 0.01171f
C3030 XThC.Tn[9] Iout 0.22393f
C3031 XThC.Tn[9] XThR.Tn[9] 0.40738f
C3032 XA.XIR[1].XIC[12].icell.PDM Vbias 0.03928f
C3033 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.Ien 0.04854f
C3034 XA.XIR[9].XIC[11].icell.PDM VPWR 0.01171f
C3035 XA.XIR[13].XIC[12].icell.PDM VPWR 0.01171f
C3036 XThC.Tn[5] XThR.Tn[12] 0.40738f
C3037 XThC.Tn[8] XA.XIR[11].XIC[8].icell.Ien 0.04604f
C3038 XThC.Tn[14] XThR.Tn[8] 0.40742f
C3039 XA.XIR[0].XIC[3].icell.PDM VPWR 0.01132f
C3040 XA.XIR[4].XIC[12].icell.PDM Vbias 0.03928f
C3041 XA.XIR[7].XIC[3].icell.Ien Vbias 0.19161f
C3042 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.Ien 0.04854f
C3043 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.Ien 0.04854f
C3044 XThC.XTB6.Y a_5949_10571# 0.01283f
C3045 XThR.XTB3.Y a_n1049_7493# 0.23056f
C3046 XThC.XTBN.Y XThC.Tn[3] 0.49586f
C3047 XThC.XTB7.B Vbias 0.12116f
C3048 XA.XIR[13].XIC_15.icell.Ien Vbias 0.19195f
C3049 XThC.Tn[0] XThR.Tn[4] 0.40739f
C3050 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.Ien 0.04854f
C3051 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.PDM 0.02104f
C3052 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.Ien 0.04854f
C3053 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.02601f
C3054 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.PDM 0.02104f
C3055 XThR.XTBN.A VPWR 0.90694f
C3056 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PDM 0.02601f
C3057 XThC.XTBN.A data[1] 0.01444f
C3058 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12] 0.14211f
C3059 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.PDM 0.02104f
C3060 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PDM 0.04035f
C3061 XThC.Tn[5] XA.XIR[4].XIC[5].icell.Ien 0.04604f
C3062 XThR.XTB5.Y a_n1049_6405# 0.24821f
C3063 XA.XIR[11].XIC[14].icell.Ien VPWR 0.18835f
C3064 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PDM 0.04042f
C3065 XThR.Tn[6] VPWR 7.9997f
C3066 XThR.XTB3.Y XThR.XTB6.Y 0.04428f
C3067 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3068 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.PDM 0.02104f
C3069 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PDM 0.02601f
C3070 XThC.XTB4.Y XThC.Tn[7] 0.01805f
C3071 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Ien 0.01532f
C3072 XA.XIR[6].XIC_15.icell.Ien VPWR 0.26829f
C3073 XThC.Tn[4] XThR.Tn[10] 0.40738f
C3074 XThR.Tn[14] XA.XIR[14].XIC[12].icell.Ien 0.14211f
C3075 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.Ien 0.04854f
C3076 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PDM 0.02601f
C3077 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3078 XA.XIR[14].XIC_15.icell.PUM VPWR 0.01655f
C3079 XA.XIR[6].XIC[11].icell.Ien Iout 0.06801f
C3080 XThC.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.04292f
C3081 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.PDM 0.02104f
C3082 XA.XIR[14].XIC[9].icell.Ien VPWR 0.18883f
C3083 Vbias bias[0] 0.21039f
C3084 bias[1] bias[2] 0.16429f
C3085 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.Ien 0.04854f
C3086 a_4861_9615# XThC.Tn[3] 0.26251f
C3087 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.Ien 0.04854f
C3088 XA.XIR[14].XIC[5].icell.Ien Iout 0.06801f
C3089 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR 0.38902f
C3090 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3091 XA.XIR[13].XIC[7].icell.Ien Iout 0.06801f
C3092 XThR.Tn[3] XA.XIR[3].XIC[2].icell.Ien 0.14211f
C3093 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0222f
C3094 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.PDM 0.02104f
C3095 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.Ien 0.04854f
C3096 XA.XIR[6].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3097 XA.XIR[15].XIC[1].icell.Ien Vbias 0.15966f
C3098 XA.XIR[14].XIC_dummy_right.icell.Iout XA.XIR[15].XIC_dummy_right.icell.Iout 0.04047f
C3099 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PDM 0.04035f
C3100 XA.XIR[11].XIC[2].icell.PDM Vbias 0.03928f
C3101 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PDM 0.02602f
C3102 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PDM 0.04035f
C3103 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.PDM 0.02104f
C3104 XA.XIR[10].XIC[6].icell.PDM Vbias 0.03928f
C3105 XA.XIR[5].XIC[1].icell.PDM VPWR 0.01171f
C3106 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.02601f
C3107 XThC.Tn[2] XThR.Tn[14] 0.40738f
C3108 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PDM 0.04035f
C3109 XThC.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.04604f
C3110 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.02601f
C3111 XThR.Tn[4] VPWR 8.03623f
C3112 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.PDM 0.02104f
C3113 XA.XIR[12].XIC[0].icell.PDM VPWR 0.01171f
C3114 XThC.Tn[10] XA.XIR[2].XIC[10].icell.Ien 0.04605f
C3115 XA.XIR[15].XIC[6].icell.Ien Vbias 0.15966f
C3116 XA.XIR[2].XIC[14].icell.Ien Iout 0.06801f
C3117 a_n1049_7493# VPWR 0.72084f
C3118 XThR.Tn[8] XA.XIR[8].XIC_15.icell.Ien 0.13564f
C3119 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.Ien 0.04854f
C3120 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.Ien 0.04854f
C3121 XA.XIR[11].XIC[6].icell.PDM VPWR 0.01171f
C3122 XA.XIR[11].XIC[12].icell.Ien VPWR 0.18829f
C3123 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.PDM 0.02104f
C3124 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PDM 0.02601f
C3125 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.Ien 0.04854f
C3126 XA.XIR[4].XIC[9].icell.Ien Vbias 0.19161f
C3127 XA.XIR[14].XIC[0].icell.Ien Iout 0.06795f
C3128 XA.XIR[0].XIC[0].icell.Ien Vbias 0.19209f
C3129 XA.XIR[10].XIC[10].icell.PDM VPWR 0.01171f
C3130 XThR.Tn[14] XA.XIR[14].XIC[10].icell.Ien 0.14211f
C3131 XThR.Tn[13] Iout 1.12765f
C3132 XThR.XTB6.Y VPWR 1.05512f
C3133 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.PDM 0.02104f
C3134 XA.XIR[8].XIC[3].icell.Ien Vbias 0.19161f
C3135 XThC.Tn[13] VPWR 4.60106f
C3136 XThR.Tn[5] XA.XIR[5].XIC[14].icell.Ien 0.144f
C3137 XA.XIR[13].XIC[11].icell.PDM VPWR 0.01171f
C3138 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.PDM 0.02104f
C3139 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.Ien 0.04854f
C3140 XA.XIR[0].XIC[14].icell.PDM Vbias 0.03945f
C3141 XA.XIR[5].XIC[8].icell.Ien VPWR 0.18829f
C3142 XA.XIR[8].XIC_dummy_right.icell.Iout XA.XIR[9].XIC_dummy_right.icell.Iout 0.04047f
C3143 XA.XIR[10].XIC_dummy_left.icell.Iout VPWR 0.11161f
C3144 XThC.Tn[8] XA.XIR[14].XIC[8].icell.Ien 0.04604f
C3145 XA.XIR[9].XIC[12].icell.Ien Vbias 0.19161f
C3146 XThC.Tn[0] XA.XIR[11].XIC[0].icell.Ien 0.04604f
C3147 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.PDM 0.02104f
C3148 XA.XIR[5].XIC[4].icell.Ien Iout 0.06801f
C3149 XThC.XTB6.A XThC.XTB7.Y 0.01596f
C3150 XA.XIR[0].XIC[5].icell.Ien Vbias 0.19213f
C3151 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PDM 0.02601f
C3152 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.PDM 0.02104f
C3153 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.PDM 0.02104f
C3154 XA.XIR[2].XIC[2].icell.PDM VPWR 0.01171f
C3155 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PDM 0.02601f
C3156 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.PDM 0.02104f
C3157 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PDM 0.02601f
C3158 XA.XIR[12].XIC[3].icell.Ien VPWR 0.18829f
C3159 XA.XIR[14].XIC[14].icell.Ien VPWR 0.1889f
C3160 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PDM 0.02803f
C3161 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.Ien 0.04854f
C3162 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PDM 0.04035f
C3163 XA.XIR[7].XIC[8].icell.Ien Vbias 0.19161f
C3164 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PDM 0.02601f
C3165 XThC.Tn[4] XThR.Tn[13] 0.40738f
C3166 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PDM 0.02601f
C3167 XThR.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.14211f
C3168 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.PDM 0.02104f
C3169 XA.XIR[1].XIC_dummy_left.icell.Iout Iout 0.03553f
C3170 XThC.XTB2.Y a_3773_9615# 0.2342f
C3171 XThC.Tn[7] Iout 0.22453f
C3172 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.PDM 0.02104f
C3173 XThC.Tn[7] XThR.Tn[9] 0.40738f
C3174 XThC.Tn[3] XThR.Tn[8] 0.40738f
C3175 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.0404f
C3176 XThC.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.04604f
C3177 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.Ien 0.04854f
C3178 XThR.Tn[10] XA.XIR[10].XIC[13].icell.Ien 0.14211f
C3179 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.PDM 0.02104f
C3180 XA.XIR[11].XIC[10].icell.Ien VPWR 0.18829f
C3181 XA.XIR[10].XIC[0].icell.Ien Vbias 0.19149f
C3182 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PDM 0.04035f
C3183 XA.XIR[6].XIC[5].icell.PDM Vbias 0.03928f
C3184 VPWR data[3] 0.20846f
C3185 XThC.XTBN.A VPWR 0.88815f
C3186 XThR.Tn[12] XA.XIR[12].XIC[2].icell.Ien 0.14211f
C3187 XA.XIR[14].XIC[2].icell.PDM Vbias 0.03928f
C3188 XThR.Tn[3] XA.XIR[3].XIC[7].icell.Ien 0.14211f
C3189 XA.XIR[5].XIC[12].icell.PDM Vbias 0.03928f
C3190 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.PDM 0.02104f
C3191 XA.XIR[13].XIC[6].icell.PDM Vbias 0.03928f
C3192 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.PDM 0.02104f
C3193 XA.XIR[11].XIC[0].icell.Ien VPWR 0.18829f
C3194 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PDM 0.04035f
C3195 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PDM 0.02601f
C3196 XThC.Tn[5] XThC.Tn[6] 0.14629f
C3197 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3198 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.PDM 0.02104f
C3199 XA.XIR[7].XIC[2].icell.PDM VPWR 0.01171f
C3200 XThR.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.14211f
C3201 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3202 XThR.Tn[14] XA.XIR[14].XIC_15.icell.Ien 0.13564f
C3203 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.PDM 0.02104f
C3204 XA.XIR[6].XIC[9].icell.PDM VPWR 0.01171f
C3205 XA.XIR[15].XIC[0].icell.PDM VPWR 0.01512f
C3206 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.Ien 0.04854f
C3207 XA.XIR[14].XIC[6].icell.PDM VPWR 0.01171f
C3208 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3209 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.PDM 0.02104f
C3210 XA.XIR[14].XIC[12].icell.Ien VPWR 0.18883f
C3211 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.PDM 0.02104f
C3212 XA.XIR[3].XIC[5].icell.Ien Vbias 0.19161f
C3213 XThC.Tn[2] XA.XIR[9].XIC[2].icell.Ien 0.04604f
C3214 XA.XIR[13].XIC[10].icell.PDM VPWR 0.01171f
C3215 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.PDM 0.02104f
C3216 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PDM 0.02601f
C3217 XThC.Tn[9] XA.XIR[0].XIC[9].icell.Ien 0.04656f
C3218 XA.XIR[6].XIC_dummy_left.icell.Iout Iout 0.03553f
C3219 XThC.XTB7.Y XThC.Tn[8] 0.07809f
C3220 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.Ien 0.04854f
C3221 XA.XIR[9].XIC[4].icell.Ien VPWR 0.18829f
C3222 XThR.Tn[0] XThR.Tn[1] 0.27134f
C3223 XThC.Tn[12] Vbias 0.8219f
C3224 XA.XIR[3].XIC[7].icell.PDM Vbias 0.03928f
C3225 XThC.Tn[3] XA.XIR[1].XIC[3].icell.Ien 0.04607f
C3226 XA.XIR[8].XIC[9].icell.PDM Vbias 0.03928f
C3227 XA.XIR[4].XIC[14].icell.Ien Vbias 0.19161f
C3228 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.Ien 0.04854f
C3229 XA.XIR[13].XIC_dummy_left.icell.Iout VPWR 0.11047f
C3230 XA.XIR[2].XIC[13].icell.PDM Vbias 0.03928f
C3231 XThR.Tn[10] XA.XIR[10].XIC[11].icell.Ien 0.14211f
C3232 XThR.XTB7.A XThR.XTB5.Y 0.11935f
C3233 XA.XIR[8].XIC[8].icell.Ien Vbias 0.19161f
C3234 XA.XIR[1].XIC[3].icell.PDM VPWR 0.01171f
C3235 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PDM 0.02601f
C3236 XA.XIR[10].XIC_15.icell.PDM Vbias 0.03927f
C3237 XThC.Tn[11] XA.XIR[4].XIC[11].icell.Ien 0.04604f
C3238 XA.XIR[5].XIC[13].icell.Ien VPWR 0.18829f
C3239 XA.XIR[4].XIC[3].icell.PDM VPWR 0.01171f
C3240 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Iout 0.01728f
C3241 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.PDM 0.02104f
C3242 XA.XIR[5].XIC[9].icell.Ien Iout 0.06801f
C3243 XA.XIR[3].XIC[11].icell.PDM VPWR 0.01171f
C3244 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Iout 0.01728f
C3245 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3246 XThC.XTB3.Y VPWR 1.07064f
C3247 XThC.XTB1.Y XThC.Tn[0] 0.1842f
C3248 XA.XIR[8].XIC[13].icell.PDM VPWR 0.01171f
C3249 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.02601f
C3250 XThC.Tn[14] XThR.Tn[3] 0.40742f
C3251 XThC.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.04604f
C3252 XThC.Tn[2] VPWR 3.64821f
C3253 XA.XIR[0].XIC[10].icell.Ien Vbias 0.19213f
C3254 XThC.XTBN.A a_9827_9569# 0.09118f
C3255 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PDM 0.04035f
C3256 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PDM 0.04035f
C3257 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.PDM 0.02104f
C3258 XA.XIR[11].XIC_15.icell.PDM VPWR 0.07527f
C3259 XA.XIR[11].XIC_15.icell.Ien VPWR 0.26829f
C3260 XA.XIR[12].XIC[8].icell.Ien VPWR 0.18829f
C3261 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3262 XThC.Tn[8] XThR.Tn[0] 0.40759f
C3263 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.Ien 0.04854f
C3264 XA.XIR[12].XIC[4].icell.Ien Iout 0.06801f
C3265 XThC.Tn[10] XThR.Tn[5] 0.40738f
C3266 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.PDM 0.02104f
C3267 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.Ien 0.04854f
C3268 XA.XIR[7].XIC[13].icell.Ien Vbias 0.19161f
C3269 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.Ien 0.04854f
C3270 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.PDM 0.02104f
C3271 XThR.Tn[4] XA.XIR[4].XIC[9].icell.Ien 0.14211f
C3272 XA.XIR[14].XIC[10].icell.Ien VPWR 0.18883f
C3273 XThC.Tn[0] XA.XIR[7].XIC[0].icell.Ien 0.04604f
C3274 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.Ien 0.04854f
C3275 XThC.XTB5.Y a_5155_9615# 0.24821f
C3276 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.Ien 0.04854f
C3277 XA.XIR[13].XIC[0].icell.Ien Vbias 0.19149f
C3278 XThC.XTB7.A a_4067_9615# 0.0127f
C3279 XThR.XTB1.Y XThR.XTB7.A 0.48957f
C3280 XThC.XTBN.A XThC.XTB7.B 0.35142f
C3281 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PDM 0.04056f
C3282 XA.XIR[11].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3283 XA.XIR[7].XIC_15.icell.PUM VPWR 0.01655f
C3284 XThR.Tn[7] XA.XIR[7].XIC[2].icell.Ien 0.14211f
C3285 XThC.Tn[3] XA.XIR[6].XIC[3].icell.Ien 0.04604f
C3286 XA.XIR[7].XIC[13].icell.PDM Vbias 0.03928f
C3287 XThC.Tn[9] XA.XIR[3].XIC[9].icell.Ien 0.04604f
C3288 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR 0.08252f
C3289 XA.XIR[4].XIC[1].icell.Ien VPWR 0.18829f
C3290 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.Ien 0.04854f
C3291 XThC.Tn[4] XA.XIR[12].XIC[4].icell.Ien 0.04604f
C3292 XThR.Tn[12] XA.XIR[12].XIC[7].icell.Ien 0.14211f
C3293 XThC.XTBN.Y a_5155_9615# 0.07602f
C3294 XThR.Tn[3] XA.XIR[3].XIC[12].icell.Ien 0.14211f
C3295 XThC.XTB1.Y VPWR 1.11809f
C3296 XA.XIR[9].XIC[9].icell.PDM Vbias 0.03928f
C3297 a_10915_9569# Vbias 0.01451f
C3298 XThC.XTB5.Y XThC.XTB6.Y 2.12831f
C3299 XA.XIR[0].XIC[1].icell.PDM Vbias 0.03945f
C3300 XA.XIR[15].XIC[3].icell.Ien VPWR 0.31713f
C3301 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PDM 0.02601f
C3302 XThR.Tn[7] Iout 1.1276f
C3303 XA.XIR[10].XIC_dummy_right.icell.Iout XA.XIR[11].XIC_dummy_right.icell.Iout 0.04047f
C3304 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PDM 0.02601f
C3305 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.02601f
C3306 XThR.Tn[2] XA.XIR[2].XIC[7].icell.Ien 0.14211f
C3307 XA.XIR[4].XIC[6].icell.Ien VPWR 0.18829f
C3308 XThC.XTB7.A XThC.Tn[3] 0.0337f
C3309 XThR.Tn[1] XA.XIR[1].XIC[0].icell.Ien 0.14251f
C3310 XA.XIR[14].XIC_dummy_left.icell.Ien XThR.Tn[14] 0.01244f
C3311 XA.XIR[4].XIC[2].icell.Ien Iout 0.06801f
C3312 XThR.XTB7.B XThR.XTB5.Y 0.30227f
C3313 VPWR bias[2] 1.20331f
C3314 a_2979_9615# XThC.Tn[0] 0.27729f
C3315 XA.XIR[3].XIC[10].icell.Ien Vbias 0.19161f
C3316 XA.XIR[1].XIC[14].icell.PDM Vbias 0.03928f
C3317 XA.XIR[10].XIC[14].icell.PDM Vbias 0.03928f
C3318 XThC.Tn[12] XThR.Tn[6] 0.40738f
C3319 XA.XIR[9].XIC[13].icell.PDM VPWR 0.01171f
C3320 XA.XIR[7].XIC[0].icell.Ien VPWR 0.18829f
C3321 XThC.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.04604f
C3322 XA.XIR[0].XIC[5].icell.PDM VPWR 0.01261f
C3323 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.PDM 0.02104f
C3324 XA.XIR[2].XIC[3].icell.Ien Vbias 0.19161f
C3325 XA.XIR[4].XIC[14].icell.PDM Vbias 0.03928f
C3326 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.Ien 0.04854f
C3327 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.PDM 0.02104f
C3328 XThC.XTB6.Y XThC.XTBN.Y 0.18947f
C3329 XA.XIR[9].XIC[9].icell.Ien VPWR 0.18829f
C3330 XA.XIR[13].XIC_15.icell.PDM Vbias 0.03927f
C3331 XA.XIR[1].XIC[5].icell.Ien Vbias 0.19173f
C3332 XThC.Tn[14] XThR.Tn[11] 0.40742f
C3333 XA.XIR[9].XIC[5].icell.Ien Iout 0.06801f
C3334 XThR.Tn[9] XA.XIR[9].XIC[5].icell.Ien 0.14211f
C3335 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PDM 0.04035f
C3336 XThC.XTB4.Y XThC.XTB5.Y 2.06459f
C3337 XA.XIR[0].XIC[2].icell.Ien VPWR 0.18776f
C3338 XThC.XTB3.Y XThC.XTB7.B 0.23315f
C3339 XThC.Tn[4] XThR.Tn[7] 0.40738f
C3340 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.Ien 0.04854f
C3341 XA.XIR[11].XIC[14].icell.PDM VPWR 0.0118f
C3342 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PDM 0.04035f
C3343 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PDM 0.04035f
C3344 XA.XIR[8].XIC[13].icell.Ien Vbias 0.19161f
C3345 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.02602f
C3346 XThC.XTB7.Y XThC.Tn[6] 0.2182f
C3347 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.PDM 0.02104f
C3348 XThC.Tn[1] Vbias 0.83728f
C3349 XA.XIR[14].XIC_15.icell.PDM VPWR 0.07527f
C3350 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PDM 0.02601f
C3351 XA.XIR[14].XIC_15.icell.Ien VPWR 0.26861f
C3352 XA.XIR[7].XIC[5].icell.Ien VPWR 0.18829f
C3353 XThC.XTB6.Y XThC.Tn[10] 0.02478f
C3354 XThC.Tn[10] XA.XIR[5].XIC[10].icell.Ien 0.04604f
C3355 XA.XIR[5].XIC[14].icell.Ien Iout 0.06801f
C3356 XThC.Tn[8] XThR.Tn[1] 0.40744f
C3357 XThR.Tn[0] XA.XIR[0].XIC[1].icell.Ien 0.14211f
C3358 XA.XIR[0].XIC_15.icell.Ien Vbias 0.19241f
C3359 XThR.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.14211f
C3360 XA.XIR[8].XIC_15.icell.PUM VPWR 0.01655f
C3361 XThR.XTB7.B XThR.XTB1.Y 1.61695f
C3362 XThC.XTB4.Y XThC.XTBN.Y 0.15636f
C3363 XThC.Tn[8] XThR.Tn[12] 0.40738f
C3364 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PDM 0.02601f
C3365 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.Ien 0.04854f
C3366 XA.XIR[6].XIC[0].icell.Ien Vbias 0.19149f
C3367 XA.XIR[12].XIC[9].icell.Ien Iout 0.06801f
C3368 XThC.Tn[3] XThR.Tn[3] 0.40738f
C3369 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.PDM 0.02104f
C3370 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PDM 0.04056f
C3371 XA.XIR[14].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3372 XThC.Tn[12] XThR.Tn[4] 0.40738f
C3373 XThR.Tn[4] XA.XIR[4].XIC[14].icell.Ien 0.144f
C3374 XThC.Tn[14] XA.XIR[10].XIC[14].icell.Ien 0.04604f
C3375 a_2979_9615# VPWR 0.70527f
C3376 XA.XIR[9].XIC[0].icell.Ien Iout 0.06795f
C3377 XA.XIR[11].XIC[4].icell.PDM Vbias 0.03928f
C3378 XThR.Tn[0] XA.XIR[0].XIC[6].icell.Ien 0.14211f
C3379 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9] 0.14211f
C3380 XThR.Tn[10] XA.XIR[10].XIC[5].icell.Ien 0.14211f
C3381 XThC.XTB4.Y XThC.Tn[10] 0.01405f
C3382 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PDM 0.04035f
C3383 XA.XIR[10].XIC[8].icell.PDM Vbias 0.03928f
C3384 XThC.Tn[12] XA.XIR[11].XIC[12].icell.Ien 0.04604f
C3385 XA.XIR[5].XIC[3].icell.PDM VPWR 0.01171f
C3386 XThC.Tn[6] XThR.Tn[0] 0.40767f
C3387 XThC.XTB4.Y a_4861_9615# 0.23756f
C3388 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PDM 0.02601f
C3389 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PDM 0.0404f
C3390 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.Ien 0.04854f
C3391 XA.XIR[6].XIC[5].icell.Ien Vbias 0.19161f
C3392 XThR.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.14211f
C3393 XThC.Tn[12] XThC.Tn[13] 0.17915f
C3394 XA.XIR[12].XIC[2].icell.PDM VPWR 0.01171f
C3395 XThC.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.04604f
C3396 XThC.XTB1.Y XThC.XTB7.B 1.61695f
C3397 XThC.XTB2.Y XThC.XTB5.Y 0.0451f
C3398 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PDM 0.02601f
C3399 XA.XIR[11].XIC[8].icell.PDM VPWR 0.01171f
C3400 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PDM 0.02602f
C3401 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.02601f
C3402 XThR.XTBN.Y XThR.XTB5.Y 0.16186f
C3403 XA.XIR[2].XIC[0].icell.PDM Vbias 0.03915f
C3404 XThC.Tn[9] XA.XIR[1].XIC[9].icell.Ien 0.04606f
C3405 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PDM 0.04042f
C3406 XA.XIR[3].XIC[2].icell.Ien VPWR 0.18829f
C3407 XA.XIR[10].XIC[13].icell.PDM Vbias 0.03928f
C3408 XThC.Tn[0] XA.XIR[8].XIC[0].icell.Ien 0.04604f
C3409 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.PDM 0.02104f
C3410 XA.XIR[15].XIC[8].icell.Ien VPWR 0.31713f
C3411 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PDM 0.02601f
C3412 XA.XIR[11].XIC[4].icell.Ien Vbias 0.19161f
C3413 XA.XIR[13].XIC[14].icell.PDM Vbias 0.03928f
C3414 XThC.XTBN.Y a_7875_9569# 0.229f
C3415 XThR.Tn[2] XA.XIR[2].XIC[12].icell.Ien 0.14211f
C3416 XThR.Tn[13] XA.XIR[13].XIC[11].icell.Ien 0.14211f
C3417 XA.XIR[15].XIC[4].icell.Ien Iout 0.07192f
C3418 XA.XIR[4].XIC[11].icell.Ien VPWR 0.18829f
C3419 XA.XIR[8].XIC[0].icell.PDM VPWR 0.01171f
C3420 XA.XIR[10].XIC[6].icell.Ien Vbias 0.19161f
C3421 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.PDM 0.02104f
C3422 XThC.XTB2.Y XThC.XTBN.Y 0.2075f
C3423 XThC.Tn[5] XThR.Tn[2] 0.40741f
C3424 XThR.XTB4.Y XThR.XTB5.Y 2.06459f
C3425 XA.XIR[4].XIC[7].icell.Ien Iout 0.06801f
C3426 XA.XIR[2].XIC[4].icell.PDM VPWR 0.01171f
C3427 XA.XIR[11].XIC[13].icell.PDM VPWR 0.01171f
C3428 XThC.Tn[14] XThR.Tn[14] 0.40742f
C3429 XA.XIR[8].XIC[5].icell.Ien VPWR 0.18829f
C3430 XA.XIR[3].XIC_15.icell.Ien Vbias 0.19195f
C3431 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Iout 0.01728f
C3432 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.Ien 0.04854f
C3433 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.Ien 0.04854f
C3434 XThC.Tn[13] XA.XIR[7].XIC[13].icell.Ien 0.04604f
C3435 XThR.XTB5.Y XThR.Tn[10] 0.01742f
C3436 XA.XIR[14].XIC[14].icell.PDM VPWR 0.0118f
C3437 XA.XIR[2].XIC[8].icell.Ien Vbias 0.19161f
C3438 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PDM 0.04035f
C3439 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout 0.06446f
C3440 XA.XIR[7].XIC[1].icell.Ien Iout 0.06801f
C3441 XA.XIR[9].XIC[14].icell.Ien VPWR 0.18835f
C3442 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.PDM 0.02104f
C3443 XA.XIR[1].XIC[10].icell.Ien Vbias 0.19173f
C3444 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PDM 0.02601f
C3445 XA.XIR[9].XIC[10].icell.Ien Iout 0.06801f
C3446 XThR.XTB1.Y XThR.XTBN.Y 0.20262f
C3447 XThR.Tn[9] XA.XIR[9].XIC[10].icell.Ien 0.14211f
C3448 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.Ien 0.04854f
C3449 XA.XIR[0].XIC[7].icell.Ien VPWR 0.18776f
C3450 XThC.Tn[1] XThR.Tn[6] 0.40738f
C3451 XA.XIR[12].XIC[14].icell.Ien Iout 0.06801f
C3452 XA.XIR[0].XIC[3].icell.Ien Iout 0.0675f
C3453 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PDM 0.04035f
C3454 XThC.Tn[4] XA.XIR[15].XIC[4].icell.Ien 0.04292f
C3455 XThC.XTBN.A XThC.Tn[12] 0.22871f
C3456 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3457 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.PDM 0.02104f
C3458 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.04035f
C3459 XThR.Tn[5] a_n1049_5611# 0.27042f
C3460 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PDM 0.02601f
C3461 XA.XIR[7].XIC[10].icell.Ien VPWR 0.18829f
C3462 XThC.Tn[3] XThR.Tn[11] 0.40738f
C3463 XA.XIR[0].XIC_dummy_right.icell.Iout XA.XIR[1].XIC_dummy_right.icell.Iout 0.04047f
C3464 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR 0.38902f
C3465 XA.XIR[7].XIC[6].icell.Ien Iout 0.06801f
C3466 XThC.Tn[5] XA.XIR[11].XIC[5].icell.Ien 0.04604f
C3467 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PDM 0.04035f
C3468 XA.XIR[7].XIC[0].icell.PDM Vbias 0.03915f
C3469 XThC.Tn[9] XA.XIR[6].XIC[9].icell.Ien 0.04604f
C3470 XThR.XTB1.Y XThR.XTB4.Y 0.05121f
C3471 XA.XIR[6].XIC[7].icell.PDM Vbias 0.03928f
C3472 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.PDM 0.02104f
C3473 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.Ien 0.04854f
C3474 XThR.Tn[6] XA.XIR[6].XIC[0].icell.Ien 0.14211f
C3475 XA.XIR[8].XIC[0].icell.Ien VPWR 0.18829f
C3476 XThC.Tn[14] XA.XIR[13].XIC[14].icell.Ien 0.04604f
C3477 XA.XIR[5].XIC[14].icell.PDM Vbias 0.03928f
C3478 XA.XIR[14].XIC[4].icell.PDM Vbias 0.03928f
C3479 XThC.XTB5.Y XThC.Tn[4] 0.20108f
C3480 XThC.Tn[12] XA.XIR[14].XIC[12].icell.Ien 0.04604f
C3481 XA.XIR[13].XIC[8].icell.PDM Vbias 0.03928f
C3482 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.Ien 0.04854f
C3483 XThR.Tn[11] XA.XIR[11].XIC[6].icell.Ien 0.14211f
C3484 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PDM 0.04035f
C3485 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PDM 0.02601f
C3486 XA.XIR[7].XIC[4].icell.PDM VPWR 0.01171f
C3487 XThC.Tn[6] XThR.Tn[1] 0.40744f
C3488 XThC.Tn[10] Iout 0.22426f
C3489 XThR.XTB6.A XThR.XTB7.A 0.44014f
C3490 XA.XIR[12].XIC_dummy_left.icell.Iout XA.XIR[13].XIC_dummy_left.icell.Iout 0.03665f
C3491 XThC.Tn[10] XThR.Tn[9] 0.40738f
C3492 XA.XIR[15].XIC[2].icell.PDM VPWR 0.01512f
C3493 XThR.Tn[0] XA.XIR[0].XIC[11].icell.Ien 0.14211f
C3494 XA.XIR[6].XIC[11].icell.PDM VPWR 0.01171f
C3495 XThC.Tn[6] XThR.Tn[12] 0.40738f
C3496 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PDM 0.02601f
C3497 XThR.Tn[6] XA.XIR[6].XIC[5].icell.Ien 0.14211f
C3498 XA.XIR[14].XIC[8].icell.PDM VPWR 0.01171f
C3499 XThR.XTB5.Y a_n997_1803# 0.06458f
C3500 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.Ien 0.04854f
C3501 XA.XIR[10].XIC[12].icell.PDM Vbias 0.03928f
C3502 XA.XIR[13].XIC_dummy_right.icell.Iout XA.XIR[14].XIC_dummy_right.icell.Iout 0.04047f
C3503 XA.XIR[1].XIC[1].icell.PDM Vbias 0.03928f
C3504 XA.XIR[6].XIC[10].icell.Ien Vbias 0.19161f
C3505 XThC.XTBN.Y XThC.Tn[4] 0.49752f
C3506 XThC.Tn[1] XThR.Tn[4] 0.40738f
C3507 XThR.Tn[7] XA.XIR[7].XIC[12].icell.Ien 0.14211f
C3508 XA.XIR[9].XIC[0].icell.PDM VPWR 0.01171f
C3509 XA.XIR[4].XIC[1].icell.PDM Vbias 0.03928f
C3510 XA.XIR[13].XIC[13].icell.PDM Vbias 0.03928f
C3511 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3512 XA.XIR[12].XIC[12].icell.Ien Iout 0.06801f
C3513 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PDM 0.02601f
C3514 XA.XIR[3].XIC[9].icell.PDM Vbias 0.03928f
C3515 XA.XIR[14].XIC[4].icell.Ien Vbias 0.19161f
C3516 XA.XIR[8].XIC[11].icell.PDM Vbias 0.03928f
C3517 XThC.Tn[13] XA.XIR[8].XIC[13].icell.Ien 0.04604f
C3518 XThC.Tn[5] XThR.Tn[10] 0.40738f
C3519 XThC.Tn[0] XA.XIR[5].XIC[0].icell.Ien 0.04604f
C3520 XA.XIR[11].XIC[12].icell.PDM VPWR 0.01171f
C3521 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.Ien 0.04854f
C3522 XA.XIR[2].XIC_15.icell.PDM Vbias 0.03927f
C3523 XA.XIR[13].XIC[6].icell.Ien Vbias 0.19161f
C3524 XA.XIR[3].XIC[7].icell.Ien VPWR 0.18829f
C3525 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.Ien 0.04854f
C3526 XA.XIR[1].XIC[5].icell.PDM VPWR 0.01171f
C3527 XA.XIR[8].XIC[1].icell.Ien Iout 0.06801f
C3528 XA.XIR[14].XIC[13].icell.PDM VPWR 0.01171f
C3529 XA.XIR[3].XIC[3].icell.Ien Iout 0.06801f
C3530 XA.XIR[4].XIC[5].icell.PDM VPWR 0.01171f
C3531 XA.XIR[11].XIC[9].icell.Ien Vbias 0.19161f
C3532 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PDM 0.04035f
C3533 XA.XIR[15].XIC[9].icell.Ien Iout 0.07192f
C3534 XA.XIR[3].XIC[13].icell.PDM VPWR 0.01171f
C3535 XA.XIR[1].XIC[2].icell.Ien VPWR 0.18829f
C3536 XA.XIR[8].XIC_15.icell.PDM VPWR 0.07527f
C3537 XThC.Tn[7] XA.XIR[2].XIC[7].icell.Ien 0.04605f
C3538 XA.XIR[4].XIC[12].icell.Ien Iout 0.06801f
C3539 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PDM 0.04035f
C3540 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.PDM 0.02104f
C3541 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PDM 0.04035f
C3542 XA.XIR[8].XIC[10].icell.Ien VPWR 0.18829f
C3543 XA.XIR[8].XIC[6].icell.Ien Iout 0.06801f
C3544 XA.XIR[2].XIC[13].icell.Ien Vbias 0.19161f
C3545 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR 0.01604f
C3546 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3547 XA.XIR[1].XIC_15.icell.Ien Vbias 0.19206f
C3548 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PDM 0.04035f
C3549 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.PDM 0.02104f
C3550 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.PDM 0.02104f
C3551 XThC.Tn[3] XThR.Tn[14] 0.40738f
C3552 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PDM 0.02601f
C3553 XA.XIR[9].XIC_15.icell.Ien Iout 0.0694f
C3554 XThR.Tn[9] XA.XIR[9].XIC_15.icell.Ien 0.13564f
C3555 XA.XIR[0].XIC[12].icell.Ien VPWR 0.1902f
C3556 XThC.Tn[5] XA.XIR[14].XIC[5].icell.Ien 0.04604f
C3557 XThC.XTB7.A a_5155_9615# 0.02287f
C3558 XA.XIR[0].XIC[8].icell.Ien Iout 0.0675f
C3559 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.PDM 0.02104f
C3560 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.PDM 0.02104f
C3561 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PDM 0.04039f
C3562 XA.XIR[7].XIC_15.icell.Ien VPWR 0.26829f
C3563 XA.XIR[2].XIC_15.icell.PUM VPWR 0.01655f
C3564 XA.XIR[12].XIC[10].icell.Ien Iout 0.06801f
C3565 XThR.Tn[13] XA.XIR[13].XIC[5].icell.Ien 0.14211f
C3566 XA.XIR[5].XIC[0].icell.Ien VPWR 0.18829f
C3567 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.PDM 0.02104f
C3568 XThR.XTB5.A XThR.XTB2.Y 0.02203f
C3569 XA.XIR[5].XIC[3].icell.Ien Vbias 0.19161f
C3570 XA.XIR[7].XIC[11].icell.Ien Iout 0.06801f
C3571 XThR.XTB7.B XThR.XTB6.A 1.47641f
C3572 XA.XIR[7].XIC_15.icell.PDM Vbias 0.03927f
C3573 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.Ien 0.04854f
C3574 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.PDM 0.02104f
C3575 XA.XIR[4].XIC_dummy_left.icell.Iout VPWR 0.10954f
C3576 XThC.Tn[14] VPWR 4.55561f
C3577 XThC.XTBN.Y a_6243_9615# 0.07767f
C3578 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PDM 0.02601f
C3579 XA.XIR[9].XIC_dummy_right.icell.Iout Iout 0.01732f
C3580 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.PDM 0.02104f
C3581 XA.XIR[10].XIC[11].icell.PDM Vbias 0.03928f
C3582 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout 0.06446f
C3583 XA.XIR[3].XIC[0].icell.Ien Iout 0.06795f
C3584 XThR.Tn[8] Iout 1.12761f
C3585 XThR.Tn[8] XThR.Tn[9] 0.10569f
C3586 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.Ien 0.04854f
C3587 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3588 XA.XIR[6].XIC[2].icell.Ien VPWR 0.18829f
C3589 XA.XIR[9].XIC[11].icell.PDM Vbias 0.03928f
C3590 XA.XIR[13].XIC[12].icell.PDM Vbias 0.03928f
C3591 XA.XIR[0].XIC[3].icell.PDM Vbias 0.03945f
C3592 XA.XIR[11].XIC[1].icell.Ien Iout 0.06801f
C3593 XThC.XTB7.A XThC.XTB6.Y 0.19112f
C3594 XA.XIR[7].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3595 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Ien 0.01546f
C3596 XA.XIR[10].XIC_dummy_left.icell.Ien XThR.Tn[10] 0.01244f
C3597 XA.XIR[11].XIC[11].icell.PDM VPWR 0.01171f
C3598 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Ien 0.01597f
C3599 XThR.Tn[6] XA.XIR[6].XIC[10].icell.Ien 0.14211f
C3600 XThR.XTB2.Y data[5] 0.017f
C3601 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.PDM 0.02104f
C3602 XA.XIR[11].XIC[14].icell.Ien Vbias 0.19161f
C3603 XThC.Tn[5] XThR.Tn[13] 0.40738f
C3604 XThR.Tn[6] Vbias 1.39526f
C3605 XA.XIR[14].XIC[12].icell.PDM VPWR 0.01171f
C3606 XA.XIR[6].XIC_15.icell.Ien Vbias 0.19195f
C3607 XA.XIR[15].XIC[14].icell.Ien Iout 0.07192f
C3608 XA.XIR[9].XIC_15.icell.PDM VPWR 0.07527f
C3609 XA.XIR[0].XIC[7].icell.PDM VPWR 0.01132f
C3610 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.Ien 0.04854f
C3611 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.Ien 0.04854f
C3612 XA.XIR[10].XIC[3].icell.Ien VPWR 0.18829f
C3613 XThC.Tn[4] XThR.Tn[8] 0.40738f
C3614 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.PDM 0.02104f
C3615 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.Ien 0.04854f
C3616 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.PDM 0.02104f
C3617 XA.XIR[14].XIC[9].icell.Ien Vbias 0.19161f
C3618 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PDM 0.04035f
C3619 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PDM 0.04056f
C3620 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PDM 0.04035f
C3621 XThC.XTB7.A XThC.XTB4.Y 0.14536f
C3622 XA.XIR[3].XIC[12].icell.Ien VPWR 0.18829f
C3623 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.PDM 0.02104f
C3624 XA.XIR[3].XIC[8].icell.Ien Iout 0.06801f
C3625 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.Ien 0.04854f
C3626 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.Ien 0.04854f
C3627 XA.XIR[2].XIC[5].icell.Ien VPWR 0.18829f
C3628 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.PDM 0.02104f
C3629 XThC.XTB6.Y a_5949_9615# 0.26831f
C3630 XA.XIR[1].XIC[7].icell.Ien VPWR 0.18829f
C3631 XThC.Tn[6] XA.XIR[0].XIC[6].icell.Ien 0.04659f
C3632 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.Ien 0.04854f
C3633 XThR.Tn[8] XA.XIR[8].XIC[2].icell.Ien 0.14211f
C3634 XThC.Tn[1] XThC.Tn[2] 0.71417f
C3635 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.03838f
C3636 XA.XIR[1].XIC[3].icell.Ien Iout 0.06801f
C3637 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PDM 0.02601f
C3638 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.Ien 0.04854f
C3639 XThR.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.14211f
C3640 XA.XIR[8].XIC_15.icell.Ien VPWR 0.26829f
C3641 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PDM 0.02602f
C3642 XA.XIR[12].XIC_15.icell.Ien Iout 0.0694f
C3643 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PDM 0.02601f
C3644 XA.XIR[5].XIC[1].icell.PDM Vbias 0.03928f
C3645 XThR.XTB7.A a_n1049_5317# 0.02018f
C3646 XA.XIR[8].XIC[11].icell.Ien Iout 0.06801f
C3647 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.PDM 0.02104f
C3648 XThR.Tn[4] Vbias 1.39526f
C3649 XThR.XTBN.Y XThR.XTB6.A 0.03867f
C3650 XA.XIR[12].XIC[0].icell.PDM Vbias 0.03915f
C3651 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.PDM 0.02104f
C3652 a_4067_9615# VPWR 0.70663f
C3653 XA.XIR[11].XIC[6].icell.PDM Vbias 0.03928f
C3654 XThR.XTB2.Y XThR.Tn[9] 0.292f
C3655 a_n997_3755# XThR.Tn[9] 0.19352f
C3656 XA.XIR[11].XIC[12].icell.Ien Vbias 0.19161f
C3657 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PDM 0.04035f
C3658 XA.XIR[15].XIC[12].icell.Ien Iout 0.07192f
C3659 XThC.XTB7.Y XThC.Tn[9] 0.07413f
C3660 XThR.Tn[14] XA.XIR[14].XIC[6].icell.Ien 0.14211f
C3661 XA.XIR[10].XIC[10].icell.PDM Vbias 0.03928f
C3662 XA.XIR[0].XIC[13].icell.Ien Iout 0.0675f
C3663 XThR.Tn[1] XA.XIR[1].XIC[6].icell.Ien 0.14211f
C3664 XThC.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.04604f
C3665 XA.XIR[5].XIC[5].icell.PDM VPWR 0.01171f
C3666 XThR.XTBN.Y XThR.Tn[0] 0.55717f
C3667 XA.XIR[8].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3668 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PDM 0.02601f
C3669 XA.XIR[12].XIC_dummy_right.icell.Iout Iout 0.01732f
C3670 XThC.Tn[13] Vbias 0.82511f
C3671 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.PDM 0.02104f
C3672 XA.XIR[13].XIC[11].icell.PDM Vbias 0.03928f
C3673 XThR.XTB6.A XThR.XTB4.Y 0.04137f
C3674 XA.XIR[12].XIC[4].icell.PDM VPWR 0.01171f
C3675 XA.XIR[5].XIC[8].icell.Ien Vbias 0.19161f
C3676 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.Ien 0.04854f
C3677 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.Ien 0.04854f
C3678 XThC.Tn[1] XA.XIR[4].XIC[1].icell.Ien 0.04604f
C3679 XA.XIR[11].XIC[10].icell.PDM VPWR 0.01171f
C3680 XThC.XTB2.Y XThC.XTB7.A 0.2319f
C3681 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.PDM 0.02104f
C3682 XThC.XTB5.A XThC.XTB4.Y 0.02767f
C3683 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.Ien 0.04854f
C3684 XA.XIR[14].XIC[1].icell.Ien Iout 0.06801f
C3685 XA.XIR[2].XIC[2].icell.PDM Vbias 0.03928f
C3686 XA.XIR[14].XIC[11].icell.PDM VPWR 0.01171f
C3687 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PDM 0.04035f
C3688 XA.XIR[12].XIC[3].icell.Ien Vbias 0.19161f
C3689 XA.XIR[6].XIC[7].icell.Ien VPWR 0.18829f
C3690 XThC.XTB1.Y XThC.Tn[1] 0.01068f
C3691 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.Ien 0.04854f
C3692 XA.XIR[14].XIC[14].icell.Ien Vbias 0.19161f
C3693 XThR.XTB7.A a_n1049_6405# 0.02287f
C3694 XThC.Tn[3] VPWR 3.60513f
C3695 XA.XIR[6].XIC[3].icell.Ien Iout 0.06801f
C3696 XThC.XTBN.Y a_8963_9569# 0.22784f
C3697 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PDM 0.02601f
C3698 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.PDM 0.02104f
C3699 XA.XIR[8].XIC[2].icell.PDM VPWR 0.01171f
C3700 XA.XIR[3].XIC[0].icell.PDM VPWR 0.01171f
C3701 XA.XIR[4].XIC_dummy_left.icell.Iout XA.XIR[5].XIC_dummy_left.icell.Iout 0.03665f
C3702 XThR.XTB5.A data[4] 0.14415f
C3703 XThC.Tn[9] XThR.Tn[0] 0.40759f
C3704 XThR.Tn[6] XA.XIR[6].XIC_15.icell.Ien 0.13564f
C3705 XThC.Tn[11] XThR.Tn[5] 0.40738f
C3706 XThR.Tn[1] XThR.Tn[2] 0.15279f
C3707 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.PDM 0.02104f
C3708 XThC.Tn[6] XA.XIR[3].XIC[6].icell.Ien 0.04604f
C3709 XA.XIR[2].XIC[6].icell.PDM VPWR 0.01171f
C3710 XA.XIR[13].XIC[3].icell.Ien VPWR 0.18829f
C3711 XThR.XTB1.Y a_n997_3979# 0.06353f
C3712 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.PDM 0.02104f
C3713 XThC.Tn[13] XA.XIR[2].XIC[13].icell.Ien 0.04605f
C3714 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.Ien 0.04854f
C3715 XA.XIR[11].XIC[6].icell.Ien VPWR 0.18829f
C3716 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR 0.38914f
C3717 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PDM 0.04035f
C3718 XA.XIR[2].XIC[1].icell.Ien Iout 0.06801f
C3719 XA.XIR[11].XIC[10].icell.Ien Vbias 0.19161f
C3720 XA.XIR[7].XIC_dummy_left.icell.Iout Iout 0.03553f
C3721 XA.XIR[11].XIC[2].icell.Ien Iout 0.06801f
C3722 XA.XIR[10].XIC[8].icell.Ien VPWR 0.18829f
C3723 XA.XIR[15].XIC[10].icell.Ien Iout 0.07192f
C3724 XA.XIR[10].XIC[4].icell.Ien Iout 0.06801f
C3725 XThC.XTBN.A Vbias 0.01693f
C3726 XThR.XTB7.B a_n1049_5317# 0.01743f
C3727 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PDM 0.04035f
C3728 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PDM 0.02602f
C3729 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.PDM 0.02104f
C3730 data[5] data[4] 0.64735f
C3731 XA.XIR[3].XIC[13].icell.Ien Iout 0.06801f
C3732 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.Ien 0.04854f
C3733 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PDM 0.04035f
C3734 VPWR data[6] 0.21221f
C3735 XThR.Tn[5] XA.XIR[5].XIC[1].icell.Ien 0.14211f
C3736 XThR.Tn[11] XA.XIR[11].XIC_dummy_left.icell.Iout 0.03385f
C3737 XA.XIR[2].XIC[10].icell.Ien VPWR 0.18829f
C3738 XA.XIR[11].XIC[0].icell.Ien Vbias 0.19149f
C3739 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.PDM 0.02104f
C3740 XThC.XTB5.A XThC.XTB2.Y 0.02203f
C3741 XThC.Tn[8] XThR.Tn[2] 0.40741f
C3742 XA.XIR[2].XIC[6].icell.Ien Iout 0.06801f
C3743 XThR.Tn[8] XA.XIR[8].XIC[7].icell.Ien 0.14211f
C3744 XA.XIR[1].XIC[12].icell.Ien VPWR 0.18829f
C3745 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PDM 0.04035f
C3746 XA.XIR[7].XIC[2].icell.PDM Vbias 0.03928f
C3747 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.Ien 0.04854f
C3748 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.Ien 0.04854f
C3749 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PDM 0.02792f
C3750 XA.XIR[1].XIC[8].icell.Ien Iout 0.06801f
C3751 XA.XIR[15].XIC[0].icell.PDM Vbias 0.03915f
C3752 XA.XIR[6].XIC[9].icell.PDM Vbias 0.03928f
C3753 XA.XIR[14].XIC[6].icell.PDM Vbias 0.03928f
C3754 XA.XIR[14].XIC[12].icell.Ien Vbias 0.19161f
C3755 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.PDM 0.02104f
C3756 XA.XIR[13].XIC[10].icell.PDM Vbias 0.03928f
C3757 XThC.XTB7.A XThC.Tn[4] 0.02779f
C3758 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PDM 0.02601f
C3759 XThC.Tn[4] XA.XIR[10].XIC[4].icell.Ien 0.04604f
C3760 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.PDM 0.02104f
C3761 XThR.Tn[5] XA.XIR[5].XIC[6].icell.Ien 0.14211f
C3762 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PDM 0.04035f
C3763 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3764 XThR.XTB6.Y XThR.XTBN.A 0.06405f
C3765 XThR.XTBN.Y XThR.Tn[1] 0.61094f
C3766 XA.XIR[7].XIC[6].icell.PDM VPWR 0.01171f
C3767 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.PDM 0.02104f
C3768 XA.XIR[9].XIC[4].icell.Ien Vbias 0.19161f
C3769 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.Ien 0.04854f
C3770 XA.XIR[15].XIC[4].icell.PDM VPWR 0.01512f
C3771 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.Ien 0.04854f
C3772 XA.XIR[6].XIC[13].icell.PDM VPWR 0.01171f
C3773 XThC.Tn[13] XThR.Tn[6] 0.40739f
C3774 XThC.Tn[7] XA.XIR[5].XIC[7].icell.Ien 0.04604f
C3775 XThR.XTBN.Y XThR.Tn[12] 0.50762f
C3776 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.PDM 0.02104f
C3777 XThR.Tn[1] XA.XIR[1].XIC[11].icell.Ien 0.14211f
C3778 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.PDM 0.02104f
C3779 XA.XIR[14].XIC[10].icell.PDM VPWR 0.01171f
C3780 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PDM 0.02601f
C3781 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.PDM 0.02104f
C3782 XA.XIR[13].XIC_dummy_left.icell.Ien XThR.Tn[13] 0.01244f
C3783 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.PDM 0.02104f
C3784 XA.XIR[1].XIC[3].icell.PDM Vbias 0.03928f
C3785 XA.XIR[9].XIC[2].icell.PDM VPWR 0.01171f
C3786 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.Ien 0.04854f
C3787 XA.XIR[5].XIC[13].icell.Ien Vbias 0.19161f
C3788 XThR.Tn[3] Iout 1.12764f
C3789 XA.XIR[4].XIC[3].icell.PDM Vbias 0.03928f
C3790 XThC.Tn[5] XThR.Tn[7] 0.40738f
C3791 XThC.Tn[3] XA.XIR[7].XIC[3].icell.Ien 0.04604f
C3792 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.PDM 0.02104f
C3793 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3794 XA.XIR[12].XIC[13].icell.Ien VPWR 0.18829f
C3795 XThC.XTB3.Y Vbias 0.01224f
C3796 XA.XIR[3].XIC[11].icell.PDM Vbias 0.03928f
C3797 XA.XIR[8].XIC[13].icell.PDM Vbias 0.03928f
C3798 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PDM 0.02601f
C3799 XThC.XTB7.Y XThC.Tn[7] 0.08399f
C3800 XThC.Tn[2] Vbias 0.83223f
C3801 XThC.XTB6.Y XThC.Tn[11] 0.02473f
C3802 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PDM 0.04035f
C3803 XThR.XTB7.Y XThR.Tn[9] 0.07413f
C3804 XA.XIR[11].XIC_15.icell.PDM Vbias 0.03927f
C3805 XA.XIR[1].XIC[7].icell.PDM VPWR 0.01171f
C3806 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Iout 0.01728f
C3807 XA.XIR[8].XIC_dummy_left.icell.Iout Iout 0.03553f
C3808 XA.XIR[11].XIC_15.icell.Ien Vbias 0.19195f
C3809 XA.XIR[12].XIC[8].icell.Ien Vbias 0.19161f
C3810 XA.XIR[6].XIC[12].icell.Ien VPWR 0.18829f
C3811 XThC.Tn[9] XThR.Tn[1] 0.40744f
C3812 XA.XIR[15].XIC_15.icell.Ien Iout 0.0733f
C3813 XA.XIR[6].XIC[8].icell.Ien Iout 0.06801f
C3814 XA.XIR[4].XIC[7].icell.PDM VPWR 0.01171f
C3815 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.PDM 0.02104f
C3816 XA.XIR[5].XIC_15.icell.PUM VPWR 0.01655f
C3817 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PDM 0.04035f
C3818 XThC.Tn[9] XThR.Tn[12] 0.40738f
C3819 XA.XIR[3].XIC_15.icell.PDM VPWR 0.07527f
C3820 XA.XIR[14].XIC[6].icell.Ien VPWR 0.18883f
C3821 XA.XIR[14].XIC[10].icell.Ien Vbias 0.19161f
C3822 XThR.XTBN.Y a_n1049_5317# 0.07731f
C3823 XThC.Tn[5] XA.XIR[9].XIC[5].icell.Ien 0.04604f
C3824 XA.XIR[14].XIC[2].icell.Ien Iout 0.06801f
C3825 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PDM 0.04035f
C3826 XA.XIR[13].XIC[8].icell.Ien VPWR 0.18829f
C3827 XThC.Tn[4] XThR.Tn[3] 0.40738f
C3828 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout 0.06446f
C3829 XThC.Tn[12] XA.XIR[0].XIC[12].icell.Ien 0.04662f
C3830 XA.XIR[13].XIC[4].icell.Ien Iout 0.06801f
C3831 XThC.Tn[13] XThR.Tn[4] 0.40739f
C3832 XThC.Tn[11] XA.XIR[15].XIC[11].icell.Ien 0.04292f
C3833 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.Ien 0.04854f
C3834 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.PDM 0.02104f
C3835 XThC.Tn[6] XA.XIR[1].XIC[6].icell.Ien 0.04606f
C3836 XThC.XTB4.Y XThC.Tn[11] 0.30457f
C3837 XA.XIR[15].XIC_dummy_right.icell.Iout Iout 0.01732f
C3838 XThC.Tn[8] XThR.Tn[10] 0.40738f
C3839 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.01728f
C3840 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.Ien 0.04854f
C3841 XA.XIR[11].XIC[7].icell.Ien Iout 0.06801f
C3842 XThC.Tn[0] XThR.Tn[5] 0.40739f
C3843 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PDM 0.04035f
C3844 XThC.Tn[7] XThR.Tn[0] 0.40759f
C3845 XA.XIR[4].XIC[1].icell.Ien Vbias 0.19161f
C3846 XA.XIR[10].XIC[9].icell.Ien Iout 0.06801f
C3847 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.Ien 0.04854f
C3848 XThC.Tn[8] XThC.Tn[9] 0.0619f
C3849 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.Ien 0.04854f
C3850 XThC.XTB7.A a_6243_9615# 0.02018f
C3851 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3852 XThC.Tn[14] XA.XIR[4].XIC[14].icell.Ien 0.04604f
C3853 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PDM 0.04035f
C3854 XA.XIR[2].XIC_15.icell.Ien VPWR 0.26829f
C3855 XA.XIR[12].XIC[11].icell.Ien VPWR 0.18829f
C3856 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.Ien 0.04854f
C3857 XThC.XTB1.Y Vbias 0.01576f
C3858 XA.XIR[2].XIC[11].icell.Ien Iout 0.06801f
C3859 XA.XIR[15].XIC[3].icell.Ien Vbias 0.15966f
C3860 XThR.Tn[8] XA.XIR[8].XIC[12].icell.Ien 0.14211f
C3861 XThC.Tn[4] XA.XIR[13].XIC[4].icell.Ien 0.04604f
C3862 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PDM 0.02601f
C3863 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.Ien 0.04854f
C3864 XA.XIR[1].XIC[13].icell.Ien Iout 0.06801f
C3865 XA.XIR[4].XIC[6].icell.Ien Vbias 0.19161f
C3866 XA.XIR[10].XIC[1].icell.PDM VPWR 0.01171f
C3867 Vbias bias[2] 0.06133f
C3868 XThC.Tn[3] XA.XIR[8].XIC[3].icell.Ien 0.04604f
C3869 XThR.XTBN.Y a_n1049_6405# 0.07602f
C3870 XThR.Tn[12] a_n997_1803# 0.18719f
C3871 XA.XIR[12].XIC[0].icell.Ien Iout 0.06795f
C3872 XA.XIR[9].XIC[13].icell.PDM Vbias 0.03928f
C3873 XThR.Tn[5] XA.XIR[5].XIC[11].icell.Ien 0.14211f
C3874 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PDM 0.02601f
C3875 XThC.Tn[6] XThR.Tn[2] 0.40741f
C3876 XA.XIR[7].XIC[0].icell.Ien Vbias 0.19149f
C3877 XA.XIR[0].XIC[5].icell.PDM Vbias 0.03945f
C3878 XThR.Tn[11] Iout 1.12764f
C3879 XA.XIR[5].XIC[5].icell.Ien VPWR 0.18829f
C3880 XA.XIR[2].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3881 XA.XIR[9].XIC[9].icell.Ien Vbias 0.19161f
C3882 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.Ien 0.04854f
C3883 XA.XIR[0].XIC[2].icell.Ien Vbias 0.19213f
C3884 XThC.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.04604f
C3885 XA.XIR[11].XIC[14].icell.PDM Vbias 0.03928f
C3886 XThR.XTB4.Y a_n1049_6405# 0.01546f
C3887 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PDM 0.02601f
C3888 XThR.Tn[5] VPWR 8.03417f
C3889 XThC.Tn[12] XA.XIR[3].XIC[12].icell.Ien 0.04604f
C3890 XA.XIR[0].XIC[9].icell.PDM VPWR 0.01451f
C3891 XThR.Tn[2] XA.XIR[2].XIC[0].icell.Ien 0.14251f
C3892 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.Ien 0.04854f
C3893 XA.XIR[14].XIC_15.icell.PDM Vbias 0.03927f
C3894 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.PDM 0.02104f
C3895 XA.XIR[14].XIC_15.icell.Ien Vbias 0.19195f
C3896 XA.XIR[7].XIC[5].icell.Ien Vbias 0.19161f
C3897 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.PDM 0.02104f
C3898 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PDM 0.02601f
C3899 XThC.Tn[2] XThR.Tn[6] 0.40738f
C3900 XThC.Tn[7] XA.XIR[12].XIC[7].icell.Ien 0.04604f
C3901 XThR.Tn[12] XThR.Tn[13] 0.11103f
C3902 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.Ien 0.04854f
C3903 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.Ien 0.04854f
C3904 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PDM 0.04035f
C3905 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PDM 0.04035f
C3906 XThC.Tn[4] XThR.Tn[11] 0.40738f
C3907 XA.XIR[6].XIC[13].icell.Ien Iout 0.06801f
C3908 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.02601f
C3909 XA.XIR[10].XIC[14].icell.Ien Iout 0.06801f
C3910 XThC.XTB5.Y XThC.Tn[5] 0.01168f
C3911 a_10915_9569# XThC.Tn[14] 0.20879f
C3912 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR 0.38998f
C3913 a_2979_9615# Vbias 0.01381f
C3914 XThC.Tn[8] XThR.Tn[13] 0.40738f
C3915 XA.XIR[14].XIC[7].icell.Ien Iout 0.06801f
C3916 XThR.Tn[14] XA.XIR[14].XIC_dummy_left.icell.Iout 0.03385f
C3917 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Iout 0.03842f
C3918 XA.XIR[13].XIC[9].icell.Ien Iout 0.06801f
C3919 XThR.Tn[3] XA.XIR[3].XIC[4].icell.Ien 0.14211f
C3920 XA.XIR[5].XIC[3].icell.PDM Vbias 0.03928f
C3921 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.Ien 0.04854f
C3922 XThC.Tn[7] XThR.Tn[1] 0.40744f
C3923 XThC.Tn[11] XThR.Tn[9] 0.40738f
C3924 XThC.Tn[11] Iout 0.22485f
C3925 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout 0.06446f
C3926 XThC.XTB2.Y data[1] 0.017f
C3927 XThC.Tn[7] XThR.Tn[12] 0.40738f
C3928 XA.XIR[12].XIC[2].icell.PDM Vbias 0.03928f
C3929 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PDM 0.02602f
C3930 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PDM 0.02601f
C3931 a_5155_9615# VPWR 0.7051f
C3932 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PDM 0.04056f
C3933 XA.XIR[11].XIC[8].icell.PDM Vbias 0.03928f
C3934 XA.XIR[6].XIC[0].icell.PDM VPWR 0.01171f
C3935 XThC.XTBN.Y XThC.Tn[5] 0.49425f
C3936 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PDM 0.02601f
C3937 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PDM 0.04035f
C3938 XThC.Tn[2] XThR.Tn[4] 0.40738f
C3939 XA.XIR[15].XIC[13].icell.Ien VPWR 0.31713f
C3940 XA.XIR[5].XIC[7].icell.PDM VPWR 0.01171f
C3941 XA.XIR[3].XIC[2].icell.Ien Vbias 0.19161f
C3942 XA.XIR[13].XIC[1].icell.PDM VPWR 0.01171f
C3943 XThC.Tn[13] XA.XIR[5].XIC[13].icell.Ien 0.04604f
C3944 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.Ien 0.04854f
C3945 XThC.Tn[6] XThR.Tn[10] 0.40738f
C3946 XThR.XTB5.A XThR.XTB3.Y 0.01152f
C3947 XThR.XTB7.B XThR.XTB7.A 0.35833f
C3948 XA.XIR[12].XIC[6].icell.PDM VPWR 0.01171f
C3949 XThC.XTBN.A data[3] 0.07741f
C3950 data[7] VGND 0.49949f
C3951 data[6] VGND 0.47974f
C3952 data[4] VGND 0.59317f
C3953 data[5] VGND 1.17814f
C3954 Iout VGND 0.32108p
C3955 bias[2] VGND 0.8011f
C3956 bias[0] VGND 2.64942f
C3957 Vbias VGND 0.17035p
C3958 bias[1] VGND 0.72457f
C3959 data[3] VGND 0.49926f
C3960 data[2] VGND 0.48064f
C3961 data[0] VGND 0.59269f
C3962 data[1] VGND 1.17844f
C3963 VPWR VGND 0.37297p
C3964 a_n997_715# VGND 0.5638f
C3965 XA.XIR[15].XIC_dummy_right.icell.Iout VGND 0.7524f
C3966 XA.XIR[15].XIC_dummy_right.icell.SM VGND 0.01013f
C3967 XA.XIR[15].XIC_dummy_right.icell.Ien VGND 0.64532f
C3968 XA.XIR[15].XIC_15.icell.Ien VGND 0.44493f
C3969 XA.XIR[15].XIC[14].icell.Ien VGND 0.4451f
C3970 XA.XIR[15].XIC[13].icell.Ien VGND 0.44506f
C3971 XA.XIR[15].XIC[12].icell.Ien VGND 0.44506f
C3972 XA.XIR[15].XIC[11].icell.Ien VGND 0.44506f
C3973 XA.XIR[15].XIC[10].icell.Ien VGND 0.44506f
C3974 XA.XIR[15].XIC[9].icell.Ien VGND 0.44506f
C3975 XA.XIR[15].XIC[8].icell.Ien VGND 0.44506f
C3976 XA.XIR[15].XIC[7].icell.Ien VGND 0.44506f
C3977 XA.XIR[15].XIC[6].icell.Ien VGND 0.44506f
C3978 XA.XIR[15].XIC[5].icell.Ien VGND 0.44506f
C3979 XA.XIR[15].XIC[4].icell.Ien VGND 0.44506f
C3980 XA.XIR[15].XIC[3].icell.Ien VGND 0.44506f
C3981 XA.XIR[15].XIC[2].icell.Ien VGND 0.44506f
C3982 XA.XIR[15].XIC_dummy_left.icell.Iout VGND 0.70682f
C3983 XA.XIR[15].XIC[1].icell.Ien VGND 0.44506f
C3984 XA.XIR[15].XIC[0].icell.Ien VGND 0.44521f
C3985 XA.XIR[15].XIC_dummy_left.icell.SM VGND 0.01033f
C3986 XA.XIR[15].XIC_dummy_left.icell.Ien VGND 0.6116f
C3987 XA.XIR[15].XIC_dummy_right.icell.PDM VGND 0.23278f
C3988 XA.XIR[15].XIC_15.icell.PDM VGND 0.18786f
C3989 XA.XIR[15].XIC[14].icell.PDM VGND 0.18744f
C3990 XA.XIR[15].XIC[13].icell.PDM VGND 0.18744f
C3991 XA.XIR[15].XIC[12].icell.PDM VGND 0.18744f
C3992 XA.XIR[15].XIC[11].icell.PDM VGND 0.18744f
C3993 XA.XIR[15].XIC[10].icell.PDM VGND 0.18744f
C3994 XA.XIR[15].XIC[9].icell.PDM VGND 0.18744f
C3995 XA.XIR[15].XIC[8].icell.PDM VGND 0.18744f
C3996 XA.XIR[15].XIC[7].icell.PDM VGND 0.18744f
C3997 XA.XIR[15].XIC[6].icell.PDM VGND 0.18744f
C3998 XA.XIR[15].XIC[5].icell.PDM VGND 0.18744f
C3999 XA.XIR[15].XIC[4].icell.PDM VGND 0.18744f
C4000 XA.XIR[15].XIC[3].icell.PDM VGND 0.18744f
C4001 XA.XIR[15].XIC[2].icell.PDM VGND 0.18744f
C4002 XA.XIR[15].XIC[1].icell.PDM VGND 0.18744f
C4003 XA.XIR[15].XIC[0].icell.PDM VGND 0.1876f
C4004 XA.XIR[15].XIC_dummy_left.icell.PDM VGND 0.22703f
C4005 XA.XIR[14].XIC_dummy_right.icell.Iout VGND 0.85788f
C4006 XA.XIR[14].XIC_dummy_right.icell.SM VGND 0.01013f
C4007 XA.XIR[14].XIC_dummy_right.icell.Ien VGND 0.60818f
C4008 XA.XIR[14].XIC_15.icell.Ien VGND 0.37264f
C4009 XA.XIR[14].XIC[14].icell.Ien VGND 0.37333f
C4010 XA.XIR[14].XIC[13].icell.Ien VGND 0.3733f
C4011 XA.XIR[14].XIC[12].icell.Ien VGND 0.3733f
C4012 XA.XIR[14].XIC[11].icell.Ien VGND 0.3733f
C4013 XA.XIR[14].XIC[10].icell.Ien VGND 0.3733f
C4014 XA.XIR[14].XIC[9].icell.Ien VGND 0.3733f
C4015 XA.XIR[14].XIC[8].icell.Ien VGND 0.3733f
C4016 XA.XIR[14].XIC[7].icell.Ien VGND 0.3733f
C4017 XA.XIR[14].XIC[6].icell.Ien VGND 0.3733f
C4018 XA.XIR[14].XIC[5].icell.Ien VGND 0.3733f
C4019 XA.XIR[14].XIC[4].icell.Ien VGND 0.3733f
C4020 XA.XIR[14].XIC[3].icell.Ien VGND 0.3733f
C4021 XA.XIR[14].XIC[2].icell.Ien VGND 0.3733f
C4022 XA.XIR[14].XIC_dummy_left.icell.Iout VGND 0.8066f
C4023 XThR.Tn[14] VGND 13.06755f
C4024 XA.XIR[14].XIC[1].icell.Ien VGND 0.3733f
C4025 a_n997_1579# VGND 0.54776f
C4026 XA.XIR[14].XIC[0].icell.Ien VGND 0.37345f
C4027 XA.XIR[14].XIC_dummy_left.icell.SM VGND 0.01033f
C4028 XA.XIR[14].XIC_dummy_left.icell.Ien VGND 0.57576f
C4029 a_n997_1803# VGND 0.53619f
C4030 XA.XIR[14].XIC_dummy_right.icell.PDM VGND 0.23384f
C4031 XA.XIR[14].XIC_15.icell.PDM VGND 0.18862f
C4032 XA.XIR[14].XIC[14].icell.PDM VGND 0.1882f
C4033 XA.XIR[14].XIC[13].icell.PDM VGND 0.1882f
C4034 XA.XIR[14].XIC[12].icell.PDM VGND 0.1882f
C4035 XA.XIR[14].XIC[11].icell.PDM VGND 0.1882f
C4036 XA.XIR[14].XIC[10].icell.PDM VGND 0.1882f
C4037 XA.XIR[14].XIC[9].icell.PDM VGND 0.1882f
C4038 XA.XIR[14].XIC[8].icell.PDM VGND 0.1882f
C4039 XA.XIR[14].XIC[7].icell.PDM VGND 0.1882f
C4040 XA.XIR[14].XIC[6].icell.PDM VGND 0.1882f
C4041 XA.XIR[14].XIC[5].icell.PDM VGND 0.1882f
C4042 XA.XIR[14].XIC[4].icell.PDM VGND 0.1882f
C4043 XA.XIR[14].XIC[3].icell.PDM VGND 0.1882f
C4044 XA.XIR[14].XIC[2].icell.PDM VGND 0.1882f
C4045 XA.XIR[14].XIC[1].icell.PDM VGND 0.1882f
C4046 XA.XIR[14].XIC[0].icell.PDM VGND 0.18836f
C4047 XA.XIR[14].XIC_dummy_left.icell.PDM VGND 0.22809f
C4048 XA.XIR[13].XIC_dummy_right.icell.Iout VGND 0.85788f
C4049 XA.XIR[13].XIC_dummy_right.icell.SM VGND 0.01013f
C4050 XA.XIR[13].XIC_dummy_right.icell.Ien VGND 0.60818f
C4051 XA.XIR[13].XIC_15.icell.Ien VGND 0.37264f
C4052 XA.XIR[13].XIC[14].icell.Ien VGND 0.37333f
C4053 XA.XIR[13].XIC[13].icell.Ien VGND 0.3733f
C4054 XA.XIR[13].XIC[12].icell.Ien VGND 0.3733f
C4055 XA.XIR[13].XIC[11].icell.Ien VGND 0.3733f
C4056 XA.XIR[13].XIC[10].icell.Ien VGND 0.3733f
C4057 XA.XIR[13].XIC[9].icell.Ien VGND 0.3733f
C4058 XA.XIR[13].XIC[8].icell.Ien VGND 0.3733f
C4059 XA.XIR[13].XIC[7].icell.Ien VGND 0.3733f
C4060 XA.XIR[13].XIC[6].icell.Ien VGND 0.3733f
C4061 XA.XIR[13].XIC[5].icell.Ien VGND 0.3733f
C4062 XA.XIR[13].XIC[4].icell.Ien VGND 0.3733f
C4063 XA.XIR[13].XIC[3].icell.Ien VGND 0.3733f
C4064 XA.XIR[13].XIC[2].icell.Ien VGND 0.3733f
C4065 XA.XIR[13].XIC_dummy_left.icell.Iout VGND 0.80664f
C4066 XThR.Tn[13] VGND 12.91167f
C4067 XA.XIR[13].XIC[1].icell.Ien VGND 0.3733f
C4068 XA.XIR[13].XIC[0].icell.Ien VGND 0.37345f
C4069 XA.XIR[13].XIC_dummy_left.icell.SM VGND 0.01033f
C4070 XA.XIR[13].XIC_dummy_left.icell.Ien VGND 0.57422f
C4071 XA.XIR[13].XIC_dummy_right.icell.PDM VGND 0.23384f
C4072 XA.XIR[13].XIC_15.icell.PDM VGND 0.18862f
C4073 XA.XIR[13].XIC[14].icell.PDM VGND 0.1882f
C4074 XA.XIR[13].XIC[13].icell.PDM VGND 0.1882f
C4075 XA.XIR[13].XIC[12].icell.PDM VGND 0.1882f
C4076 XA.XIR[13].XIC[11].icell.PDM VGND 0.1882f
C4077 XA.XIR[13].XIC[10].icell.PDM VGND 0.1882f
C4078 XA.XIR[13].XIC[9].icell.PDM VGND 0.1882f
C4079 XA.XIR[13].XIC[8].icell.PDM VGND 0.1882f
C4080 XA.XIR[13].XIC[7].icell.PDM VGND 0.1882f
C4081 XA.XIR[13].XIC[6].icell.PDM VGND 0.1882f
C4082 XA.XIR[13].XIC[5].icell.PDM VGND 0.1882f
C4083 XA.XIR[13].XIC[4].icell.PDM VGND 0.1882f
C4084 XA.XIR[13].XIC[3].icell.PDM VGND 0.1882f
C4085 XA.XIR[13].XIC[2].icell.PDM VGND 0.1882f
C4086 XA.XIR[13].XIC[1].icell.PDM VGND 0.1882f
C4087 XA.XIR[13].XIC[0].icell.PDM VGND 0.18836f
C4088 XA.XIR[13].XIC_dummy_left.icell.PDM VGND 0.22809f
C4089 XA.XIR[12].XIC_dummy_right.icell.Iout VGND 0.85788f
C4090 XA.XIR[12].XIC_dummy_right.icell.SM VGND 0.01013f
C4091 XA.XIR[12].XIC_dummy_right.icell.Ien VGND 0.60818f
C4092 XA.XIR[12].XIC_15.icell.Ien VGND 0.37264f
C4093 XA.XIR[12].XIC[14].icell.Ien VGND 0.37333f
C4094 XA.XIR[12].XIC[13].icell.Ien VGND 0.3733f
C4095 XA.XIR[12].XIC[12].icell.Ien VGND 0.3733f
C4096 XA.XIR[12].XIC[11].icell.Ien VGND 0.3733f
C4097 XA.XIR[12].XIC[10].icell.Ien VGND 0.3733f
C4098 XA.XIR[12].XIC[9].icell.Ien VGND 0.3733f
C4099 XA.XIR[12].XIC[8].icell.Ien VGND 0.3733f
C4100 XA.XIR[12].XIC[7].icell.Ien VGND 0.3733f
C4101 XA.XIR[12].XIC[6].icell.Ien VGND 0.3733f
C4102 XA.XIR[12].XIC[5].icell.Ien VGND 0.3733f
C4103 XA.XIR[12].XIC[4].icell.Ien VGND 0.3733f
C4104 XA.XIR[12].XIC[3].icell.Ien VGND 0.3733f
C4105 XA.XIR[12].XIC[2].icell.Ien VGND 0.3733f
C4106 XA.XIR[12].XIC_dummy_left.icell.Iout VGND 0.80529f
C4107 XThR.Tn[12] VGND 12.80173f
C4108 XA.XIR[12].XIC[1].icell.Ien VGND 0.3733f
C4109 XA.XIR[12].XIC[0].icell.Ien VGND 0.37345f
C4110 XA.XIR[12].XIC_dummy_left.icell.SM VGND 0.01033f
C4111 XA.XIR[12].XIC_dummy_left.icell.Ien VGND 0.5728f
C4112 a_n997_2667# VGND 0.5457f
C4113 XA.XIR[12].XIC_dummy_right.icell.PDM VGND 0.23384f
C4114 XA.XIR[12].XIC_15.icell.PDM VGND 0.18862f
C4115 XA.XIR[12].XIC[14].icell.PDM VGND 0.1882f
C4116 XA.XIR[12].XIC[13].icell.PDM VGND 0.1882f
C4117 XA.XIR[12].XIC[12].icell.PDM VGND 0.1882f
C4118 XA.XIR[12].XIC[11].icell.PDM VGND 0.1882f
C4119 XA.XIR[12].XIC[10].icell.PDM VGND 0.1882f
C4120 XA.XIR[12].XIC[9].icell.PDM VGND 0.1882f
C4121 XA.XIR[12].XIC[8].icell.PDM VGND 0.1882f
C4122 XA.XIR[12].XIC[7].icell.PDM VGND 0.1882f
C4123 XA.XIR[12].XIC[6].icell.PDM VGND 0.1882f
C4124 XA.XIR[12].XIC[5].icell.PDM VGND 0.1882f
C4125 XA.XIR[12].XIC[4].icell.PDM VGND 0.1882f
C4126 XA.XIR[12].XIC[3].icell.PDM VGND 0.1882f
C4127 XA.XIR[12].XIC[2].icell.PDM VGND 0.1882f
C4128 XA.XIR[12].XIC[1].icell.PDM VGND 0.1882f
C4129 XA.XIR[12].XIC[0].icell.PDM VGND 0.18836f
C4130 XA.XIR[12].XIC_dummy_left.icell.PDM VGND 0.22809f
C4131 XA.XIR[11].XIC_dummy_right.icell.Iout VGND 0.85788f
C4132 XA.XIR[11].XIC_dummy_right.icell.SM VGND 0.01013f
C4133 XA.XIR[11].XIC_dummy_right.icell.Ien VGND 0.60818f
C4134 XA.XIR[11].XIC_15.icell.Ien VGND 0.37264f
C4135 XA.XIR[11].XIC[14].icell.Ien VGND 0.37333f
C4136 XA.XIR[11].XIC[13].icell.Ien VGND 0.3733f
C4137 XA.XIR[11].XIC[12].icell.Ien VGND 0.3733f
C4138 XA.XIR[11].XIC[11].icell.Ien VGND 0.3733f
C4139 XA.XIR[11].XIC[10].icell.Ien VGND 0.3733f
C4140 XA.XIR[11].XIC[9].icell.Ien VGND 0.3733f
C4141 XA.XIR[11].XIC[8].icell.Ien VGND 0.3733f
C4142 XA.XIR[11].XIC[7].icell.Ien VGND 0.3733f
C4143 XA.XIR[11].XIC[6].icell.Ien VGND 0.3733f
C4144 XA.XIR[11].XIC[5].icell.Ien VGND 0.3733f
C4145 XA.XIR[11].XIC[4].icell.Ien VGND 0.3733f
C4146 XA.XIR[11].XIC[3].icell.Ien VGND 0.3733f
C4147 XA.XIR[11].XIC[2].icell.Ien VGND 0.3733f
C4148 XA.XIR[11].XIC_dummy_left.icell.Iout VGND 0.80765f
C4149 XThR.Tn[11] VGND 12.86402f
C4150 XA.XIR[11].XIC[1].icell.Ien VGND 0.3733f
C4151 a_n997_2891# VGND 0.54795f
C4152 XA.XIR[11].XIC[0].icell.Ien VGND 0.37345f
C4153 XA.XIR[11].XIC_dummy_left.icell.SM VGND 0.01033f
C4154 XA.XIR[11].XIC_dummy_left.icell.Ien VGND 0.57294f
C4155 XA.XIR[11].XIC_dummy_right.icell.PDM VGND 0.23384f
C4156 XA.XIR[11].XIC_15.icell.PDM VGND 0.18862f
C4157 XA.XIR[11].XIC[14].icell.PDM VGND 0.1882f
C4158 XA.XIR[11].XIC[13].icell.PDM VGND 0.1882f
C4159 XA.XIR[11].XIC[12].icell.PDM VGND 0.1882f
C4160 XA.XIR[11].XIC[11].icell.PDM VGND 0.1882f
C4161 XA.XIR[11].XIC[10].icell.PDM VGND 0.1882f
C4162 XA.XIR[11].XIC[9].icell.PDM VGND 0.1882f
C4163 XA.XIR[11].XIC[8].icell.PDM VGND 0.1882f
C4164 XA.XIR[11].XIC[7].icell.PDM VGND 0.1882f
C4165 XA.XIR[11].XIC[6].icell.PDM VGND 0.1882f
C4166 XA.XIR[11].XIC[5].icell.PDM VGND 0.1882f
C4167 XA.XIR[11].XIC[4].icell.PDM VGND 0.1882f
C4168 XA.XIR[11].XIC[3].icell.PDM VGND 0.1882f
C4169 XA.XIR[11].XIC[2].icell.PDM VGND 0.1882f
C4170 XA.XIR[11].XIC[1].icell.PDM VGND 0.1882f
C4171 XA.XIR[11].XIC[0].icell.PDM VGND 0.18836f
C4172 XA.XIR[11].XIC_dummy_left.icell.PDM VGND 0.22809f
C4173 XA.XIR[10].XIC_dummy_right.icell.Iout VGND 0.85788f
C4174 XA.XIR[10].XIC_dummy_right.icell.SM VGND 0.01013f
C4175 XA.XIR[10].XIC_dummy_right.icell.Ien VGND 0.60818f
C4176 XA.XIR[10].XIC_15.icell.Ien VGND 0.37264f
C4177 XA.XIR[10].XIC[14].icell.Ien VGND 0.37333f
C4178 XA.XIR[10].XIC[13].icell.Ien VGND 0.3733f
C4179 XA.XIR[10].XIC[12].icell.Ien VGND 0.3733f
C4180 XA.XIR[10].XIC[11].icell.Ien VGND 0.3733f
C4181 XA.XIR[10].XIC[10].icell.Ien VGND 0.3733f
C4182 XA.XIR[10].XIC[9].icell.Ien VGND 0.3733f
C4183 XA.XIR[10].XIC[8].icell.Ien VGND 0.3733f
C4184 XA.XIR[10].XIC[7].icell.Ien VGND 0.3733f
C4185 XA.XIR[10].XIC[6].icell.Ien VGND 0.3733f
C4186 XA.XIR[10].XIC[5].icell.Ien VGND 0.3733f
C4187 XA.XIR[10].XIC[4].icell.Ien VGND 0.3733f
C4188 XA.XIR[10].XIC[3].icell.Ien VGND 0.3733f
C4189 XA.XIR[10].XIC[2].icell.Ien VGND 0.3733f
C4190 XA.XIR[10].XIC_dummy_left.icell.Iout VGND 0.80648f
C4191 XThR.Tn[10] VGND 12.83941f
C4192 XA.XIR[10].XIC[1].icell.Ien VGND 0.3733f
C4193 XA.XIR[10].XIC[0].icell.Ien VGND 0.37345f
C4194 XA.XIR[10].XIC_dummy_left.icell.SM VGND 0.01033f
C4195 XA.XIR[10].XIC_dummy_left.icell.Ien VGND 0.57422f
C4196 XA.XIR[10].XIC_dummy_right.icell.PDM VGND 0.23384f
C4197 XA.XIR[10].XIC_15.icell.PDM VGND 0.18862f
C4198 XA.XIR[10].XIC[14].icell.PDM VGND 0.1882f
C4199 XA.XIR[10].XIC[13].icell.PDM VGND 0.1882f
C4200 XA.XIR[10].XIC[12].icell.PDM VGND 0.1882f
C4201 XA.XIR[10].XIC[11].icell.PDM VGND 0.1882f
C4202 XA.XIR[10].XIC[10].icell.PDM VGND 0.1882f
C4203 XA.XIR[10].XIC[9].icell.PDM VGND 0.1882f
C4204 XA.XIR[10].XIC[8].icell.PDM VGND 0.1882f
C4205 XA.XIR[10].XIC[7].icell.PDM VGND 0.1882f
C4206 XA.XIR[10].XIC[6].icell.PDM VGND 0.1882f
C4207 XA.XIR[10].XIC[5].icell.PDM VGND 0.1882f
C4208 XA.XIR[10].XIC[4].icell.PDM VGND 0.1882f
C4209 XA.XIR[10].XIC[3].icell.PDM VGND 0.1882f
C4210 XA.XIR[10].XIC[2].icell.PDM VGND 0.1882f
C4211 XA.XIR[10].XIC[1].icell.PDM VGND 0.1882f
C4212 XA.XIR[10].XIC[0].icell.PDM VGND 0.18836f
C4213 XA.XIR[10].XIC_dummy_left.icell.PDM VGND 0.22809f
C4214 XA.XIR[9].XIC_dummy_right.icell.Iout VGND 0.85788f
C4215 XA.XIR[9].XIC_dummy_right.icell.SM VGND 0.01013f
C4216 XA.XIR[9].XIC_dummy_right.icell.Ien VGND 0.60818f
C4217 XA.XIR[9].XIC_15.icell.Ien VGND 0.37264f
C4218 XA.XIR[9].XIC[14].icell.Ien VGND 0.37333f
C4219 XA.XIR[9].XIC[13].icell.Ien VGND 0.3733f
C4220 XA.XIR[9].XIC[12].icell.Ien VGND 0.3733f
C4221 XA.XIR[9].XIC[11].icell.Ien VGND 0.3733f
C4222 XA.XIR[9].XIC[10].icell.Ien VGND 0.3733f
C4223 XA.XIR[9].XIC[9].icell.Ien VGND 0.3733f
C4224 XA.XIR[9].XIC[8].icell.Ien VGND 0.3733f
C4225 XA.XIR[9].XIC[7].icell.Ien VGND 0.3733f
C4226 XA.XIR[9].XIC[6].icell.Ien VGND 0.3733f
C4227 XA.XIR[9].XIC[5].icell.Ien VGND 0.3733f
C4228 XA.XIR[9].XIC[4].icell.Ien VGND 0.3733f
C4229 XA.XIR[9].XIC[3].icell.Ien VGND 0.3733f
C4230 XA.XIR[9].XIC[2].icell.Ien VGND 0.3733f
C4231 XA.XIR[9].XIC_dummy_left.icell.Iout VGND 0.80834f
C4232 XA.XIR[9].XIC[1].icell.Ien VGND 0.3733f
C4233 XThR.Tn[9] VGND 12.8472f
C4234 a_n997_3755# VGND 0.54861f
C4235 XA.XIR[9].XIC[0].icell.Ien VGND 0.37345f
C4236 XA.XIR[9].XIC_dummy_left.icell.SM VGND 0.01033f
C4237 XA.XIR[9].XIC_dummy_left.icell.Ien VGND 0.5732f
C4238 a_n997_3979# VGND 0.54721f
C4239 XA.XIR[9].XIC_dummy_right.icell.PDM VGND 0.23384f
C4240 XA.XIR[9].XIC_15.icell.PDM VGND 0.18862f
C4241 XA.XIR[9].XIC[14].icell.PDM VGND 0.1882f
C4242 XA.XIR[9].XIC[13].icell.PDM VGND 0.1882f
C4243 XA.XIR[9].XIC[12].icell.PDM VGND 0.1882f
C4244 XA.XIR[9].XIC[11].icell.PDM VGND 0.1882f
C4245 XA.XIR[9].XIC[10].icell.PDM VGND 0.1882f
C4246 XA.XIR[9].XIC[9].icell.PDM VGND 0.1882f
C4247 XA.XIR[9].XIC[8].icell.PDM VGND 0.1882f
C4248 XA.XIR[9].XIC[7].icell.PDM VGND 0.1882f
C4249 XA.XIR[9].XIC[6].icell.PDM VGND 0.1882f
C4250 XA.XIR[9].XIC[5].icell.PDM VGND 0.1882f
C4251 XA.XIR[9].XIC[4].icell.PDM VGND 0.1882f
C4252 XA.XIR[9].XIC[3].icell.PDM VGND 0.1882f
C4253 XA.XIR[9].XIC[2].icell.PDM VGND 0.1882f
C4254 XA.XIR[9].XIC[1].icell.PDM VGND 0.1882f
C4255 XA.XIR[9].XIC[0].icell.PDM VGND 0.18836f
C4256 XA.XIR[9].XIC_dummy_left.icell.PDM VGND 0.22809f
C4257 XA.XIR[8].XIC_dummy_right.icell.Iout VGND 0.85788f
C4258 XA.XIR[8].XIC_dummy_right.icell.SM VGND 0.01013f
C4259 XA.XIR[8].XIC_dummy_right.icell.Ien VGND 0.60818f
C4260 XA.XIR[8].XIC_15.icell.Ien VGND 0.37264f
C4261 XA.XIR[8].XIC[14].icell.Ien VGND 0.37333f
C4262 XA.XIR[8].XIC[13].icell.Ien VGND 0.3733f
C4263 XA.XIR[8].XIC[12].icell.Ien VGND 0.3733f
C4264 XA.XIR[8].XIC[11].icell.Ien VGND 0.3733f
C4265 XA.XIR[8].XIC[10].icell.Ien VGND 0.3733f
C4266 XA.XIR[8].XIC[9].icell.Ien VGND 0.3733f
C4267 XA.XIR[8].XIC[8].icell.Ien VGND 0.3733f
C4268 XA.XIR[8].XIC[7].icell.Ien VGND 0.3733f
C4269 XA.XIR[8].XIC[6].icell.Ien VGND 0.3733f
C4270 XA.XIR[8].XIC[5].icell.Ien VGND 0.3733f
C4271 XA.XIR[8].XIC[4].icell.Ien VGND 0.3733f
C4272 XA.XIR[8].XIC[3].icell.Ien VGND 0.3733f
C4273 XA.XIR[8].XIC[2].icell.Ien VGND 0.3733f
C4274 XA.XIR[8].XIC_dummy_left.icell.Iout VGND 0.80566f
C4275 XA.XIR[8].XIC[1].icell.Ien VGND 0.3733f
C4276 XThR.Tn[8] VGND 12.78722f
C4277 XA.XIR[8].XIC[0].icell.Ien VGND 0.37345f
C4278 XA.XIR[8].XIC_dummy_left.icell.SM VGND 0.01033f
C4279 XA.XIR[8].XIC_dummy_left.icell.Ien VGND 0.57308f
C4280 XA.XIR[8].XIC_dummy_right.icell.PDM VGND 0.23384f
C4281 XA.XIR[8].XIC_15.icell.PDM VGND 0.18862f
C4282 XA.XIR[8].XIC[14].icell.PDM VGND 0.1882f
C4283 XA.XIR[8].XIC[13].icell.PDM VGND 0.1882f
C4284 XA.XIR[8].XIC[12].icell.PDM VGND 0.1882f
C4285 XA.XIR[8].XIC[11].icell.PDM VGND 0.1882f
C4286 XA.XIR[8].XIC[10].icell.PDM VGND 0.1882f
C4287 XA.XIR[8].XIC[9].icell.PDM VGND 0.1882f
C4288 XA.XIR[8].XIC[8].icell.PDM VGND 0.1882f
C4289 XA.XIR[8].XIC[7].icell.PDM VGND 0.1882f
C4290 XA.XIR[8].XIC[6].icell.PDM VGND 0.1882f
C4291 XA.XIR[8].XIC[5].icell.PDM VGND 0.1882f
C4292 XA.XIR[8].XIC[4].icell.PDM VGND 0.1882f
C4293 XA.XIR[8].XIC[3].icell.PDM VGND 0.1882f
C4294 XA.XIR[8].XIC[2].icell.PDM VGND 0.1882f
C4295 XA.XIR[8].XIC[1].icell.PDM VGND 0.1882f
C4296 XA.XIR[8].XIC[0].icell.PDM VGND 0.18836f
C4297 XA.XIR[8].XIC_dummy_left.icell.PDM VGND 0.22809f
C4298 XA.XIR[7].XIC_dummy_right.icell.Iout VGND 0.85788f
C4299 XA.XIR[7].XIC_dummy_right.icell.SM VGND 0.01013f
C4300 XA.XIR[7].XIC_dummy_right.icell.Ien VGND 0.60818f
C4301 XA.XIR[7].XIC_15.icell.Ien VGND 0.37264f
C4302 XA.XIR[7].XIC[14].icell.Ien VGND 0.37333f
C4303 XA.XIR[7].XIC[13].icell.Ien VGND 0.3733f
C4304 XA.XIR[7].XIC[12].icell.Ien VGND 0.3733f
C4305 XA.XIR[7].XIC[11].icell.Ien VGND 0.3733f
C4306 XA.XIR[7].XIC[10].icell.Ien VGND 0.3733f
C4307 XA.XIR[7].XIC[9].icell.Ien VGND 0.3733f
C4308 XA.XIR[7].XIC[8].icell.Ien VGND 0.3733f
C4309 XA.XIR[7].XIC[7].icell.Ien VGND 0.3733f
C4310 XA.XIR[7].XIC[6].icell.Ien VGND 0.3733f
C4311 XA.XIR[7].XIC[5].icell.Ien VGND 0.3733f
C4312 XA.XIR[7].XIC[4].icell.Ien VGND 0.3733f
C4313 XA.XIR[7].XIC[3].icell.Ien VGND 0.3733f
C4314 XA.XIR[7].XIC[2].icell.Ien VGND 0.3733f
C4315 XA.XIR[7].XIC_dummy_left.icell.Iout VGND 0.80598f
C4316 XA.XIR[7].XIC[1].icell.Ien VGND 0.3733f
C4317 XA.XIR[7].XIC[0].icell.Ien VGND 0.37345f
C4318 XA.XIR[7].XIC_dummy_left.icell.SM VGND 0.01033f
C4319 XThR.Tn[7] VGND 13.23029f
C4320 XThR.XTBN.A VGND 1.22814f
C4321 XA.XIR[7].XIC_dummy_left.icell.Ien VGND 0.57576f
C4322 XA.XIR[7].XIC_dummy_right.icell.PDM VGND 0.23384f
C4323 XA.XIR[7].XIC_15.icell.PDM VGND 0.18862f
C4324 XA.XIR[7].XIC[14].icell.PDM VGND 0.1882f
C4325 XA.XIR[7].XIC[13].icell.PDM VGND 0.1882f
C4326 XA.XIR[7].XIC[12].icell.PDM VGND 0.1882f
C4327 XA.XIR[7].XIC[11].icell.PDM VGND 0.1882f
C4328 XA.XIR[7].XIC[10].icell.PDM VGND 0.1882f
C4329 XA.XIR[7].XIC[9].icell.PDM VGND 0.1882f
C4330 XA.XIR[7].XIC[8].icell.PDM VGND 0.1882f
C4331 XA.XIR[7].XIC[7].icell.PDM VGND 0.1882f
C4332 XA.XIR[7].XIC[6].icell.PDM VGND 0.1882f
C4333 XA.XIR[7].XIC[5].icell.PDM VGND 0.1882f
C4334 XA.XIR[7].XIC[4].icell.PDM VGND 0.1882f
C4335 XA.XIR[7].XIC[3].icell.PDM VGND 0.1882f
C4336 XA.XIR[7].XIC[2].icell.PDM VGND 0.1882f
C4337 XA.XIR[7].XIC[1].icell.PDM VGND 0.1882f
C4338 XA.XIR[7].XIC[0].icell.PDM VGND 0.18836f
C4339 XA.XIR[7].XIC_dummy_left.icell.PDM VGND 0.22809f
C4340 XA.XIR[6].XIC_dummy_right.icell.Iout VGND 0.85788f
C4341 XA.XIR[6].XIC_dummy_right.icell.SM VGND 0.01013f
C4342 XA.XIR[6].XIC_dummy_right.icell.Ien VGND 0.60818f
C4343 XA.XIR[6].XIC_15.icell.Ien VGND 0.37264f
C4344 XA.XIR[6].XIC[14].icell.Ien VGND 0.37333f
C4345 XA.XIR[6].XIC[13].icell.Ien VGND 0.3733f
C4346 XA.XIR[6].XIC[12].icell.Ien VGND 0.3733f
C4347 XA.XIR[6].XIC[11].icell.Ien VGND 0.3733f
C4348 XA.XIR[6].XIC[10].icell.Ien VGND 0.3733f
C4349 XA.XIR[6].XIC[9].icell.Ien VGND 0.3733f
C4350 XA.XIR[6].XIC[8].icell.Ien VGND 0.3733f
C4351 XA.XIR[6].XIC[7].icell.Ien VGND 0.3733f
C4352 XA.XIR[6].XIC[6].icell.Ien VGND 0.3733f
C4353 XA.XIR[6].XIC[5].icell.Ien VGND 0.3733f
C4354 XA.XIR[6].XIC[4].icell.Ien VGND 0.3733f
C4355 XA.XIR[6].XIC[3].icell.Ien VGND 0.3733f
C4356 XA.XIR[6].XIC[2].icell.Ien VGND 0.3733f
C4357 XA.XIR[6].XIC_dummy_left.icell.Iout VGND 0.80693f
C4358 XA.XIR[6].XIC[1].icell.Ien VGND 0.3733f
C4359 XA.XIR[6].XIC[0].icell.Ien VGND 0.37345f
C4360 XA.XIR[6].XIC_dummy_left.icell.SM VGND 0.01033f
C4361 XA.XIR[6].XIC_dummy_left.icell.Ien VGND 0.57422f
C4362 XThR.Tn[6] VGND 12.9018f
C4363 a_n1049_5317# VGND 0.02283f
C4364 XThR.XTB7.Y VGND 1.36132f
C4365 XA.XIR[6].XIC_dummy_right.icell.PDM VGND 0.23384f
C4366 XA.XIR[6].XIC_15.icell.PDM VGND 0.18862f
C4367 XA.XIR[6].XIC[14].icell.PDM VGND 0.1882f
C4368 XA.XIR[6].XIC[13].icell.PDM VGND 0.1882f
C4369 XA.XIR[6].XIC[12].icell.PDM VGND 0.1882f
C4370 XA.XIR[6].XIC[11].icell.PDM VGND 0.1882f
C4371 XA.XIR[6].XIC[10].icell.PDM VGND 0.1882f
C4372 XA.XIR[6].XIC[9].icell.PDM VGND 0.1882f
C4373 XA.XIR[6].XIC[8].icell.PDM VGND 0.1882f
C4374 XA.XIR[6].XIC[7].icell.PDM VGND 0.1882f
C4375 XA.XIR[6].XIC[6].icell.PDM VGND 0.1882f
C4376 XA.XIR[6].XIC[5].icell.PDM VGND 0.1882f
C4377 XA.XIR[6].XIC[4].icell.PDM VGND 0.1882f
C4378 XA.XIR[6].XIC[3].icell.PDM VGND 0.1882f
C4379 XA.XIR[6].XIC[2].icell.PDM VGND 0.1882f
C4380 XA.XIR[6].XIC[1].icell.PDM VGND 0.1882f
C4381 XA.XIR[6].XIC[0].icell.PDM VGND 0.18836f
C4382 XA.XIR[6].XIC_dummy_left.icell.PDM VGND 0.22809f
C4383 XA.XIR[5].XIC_dummy_right.icell.Iout VGND 0.85788f
C4384 XA.XIR[5].XIC_dummy_right.icell.SM VGND 0.01013f
C4385 XA.XIR[5].XIC_dummy_right.icell.Ien VGND 0.60818f
C4386 XA.XIR[5].XIC_15.icell.Ien VGND 0.37264f
C4387 XA.XIR[5].XIC[14].icell.Ien VGND 0.37333f
C4388 XA.XIR[5].XIC[13].icell.Ien VGND 0.3733f
C4389 XA.XIR[5].XIC[12].icell.Ien VGND 0.3733f
C4390 XA.XIR[5].XIC[11].icell.Ien VGND 0.3733f
C4391 XA.XIR[5].XIC[10].icell.Ien VGND 0.3733f
C4392 XA.XIR[5].XIC[9].icell.Ien VGND 0.3733f
C4393 XA.XIR[5].XIC[8].icell.Ien VGND 0.3733f
C4394 XA.XIR[5].XIC[7].icell.Ien VGND 0.3733f
C4395 XA.XIR[5].XIC[6].icell.Ien VGND 0.3733f
C4396 XA.XIR[5].XIC[5].icell.Ien VGND 0.3733f
C4397 XA.XIR[5].XIC[4].icell.Ien VGND 0.3733f
C4398 XA.XIR[5].XIC[3].icell.Ien VGND 0.3733f
C4399 XA.XIR[5].XIC[2].icell.Ien VGND 0.3733f
C4400 XA.XIR[5].XIC_dummy_left.icell.Iout VGND 0.80562f
C4401 XA.XIR[5].XIC[1].icell.Ien VGND 0.3733f
C4402 a_n1049_5611# VGND 0.02888f
C4403 XA.XIR[5].XIC[0].icell.Ien VGND 0.37345f
C4404 XA.XIR[5].XIC_dummy_left.icell.SM VGND 0.01033f
C4405 XA.XIR[5].XIC_dummy_left.icell.Ien VGND 0.57288f
C4406 XThR.Tn[5] VGND 12.89248f
C4407 XThR.XTB6.Y VGND 1.38212f
C4408 XA.XIR[5].XIC_dummy_right.icell.PDM VGND 0.23384f
C4409 XA.XIR[5].XIC_15.icell.PDM VGND 0.18862f
C4410 XA.XIR[5].XIC[14].icell.PDM VGND 0.1882f
C4411 XA.XIR[5].XIC[13].icell.PDM VGND 0.1882f
C4412 XA.XIR[5].XIC[12].icell.PDM VGND 0.1882f
C4413 XA.XIR[5].XIC[11].icell.PDM VGND 0.1882f
C4414 XA.XIR[5].XIC[10].icell.PDM VGND 0.1882f
C4415 XA.XIR[5].XIC[9].icell.PDM VGND 0.1882f
C4416 XA.XIR[5].XIC[8].icell.PDM VGND 0.1882f
C4417 XA.XIR[5].XIC[7].icell.PDM VGND 0.1882f
C4418 XA.XIR[5].XIC[6].icell.PDM VGND 0.1882f
C4419 XA.XIR[5].XIC[5].icell.PDM VGND 0.1882f
C4420 XA.XIR[5].XIC[4].icell.PDM VGND 0.1882f
C4421 XA.XIR[5].XIC[3].icell.PDM VGND 0.1882f
C4422 XA.XIR[5].XIC[2].icell.PDM VGND 0.1882f
C4423 XA.XIR[5].XIC[1].icell.PDM VGND 0.1882f
C4424 XA.XIR[5].XIC[0].icell.PDM VGND 0.18836f
C4425 XA.XIR[5].XIC_dummy_left.icell.PDM VGND 0.22809f
C4426 XA.XIR[4].XIC_dummy_right.icell.Iout VGND 0.85788f
C4427 XA.XIR[4].XIC_dummy_right.icell.SM VGND 0.01013f
C4428 XA.XIR[4].XIC_dummy_right.icell.Ien VGND 0.60818f
C4429 XA.XIR[4].XIC_15.icell.Ien VGND 0.37264f
C4430 XA.XIR[4].XIC[14].icell.Ien VGND 0.37333f
C4431 XA.XIR[4].XIC[13].icell.Ien VGND 0.3733f
C4432 XA.XIR[4].XIC[12].icell.Ien VGND 0.3733f
C4433 XA.XIR[4].XIC[11].icell.Ien VGND 0.3733f
C4434 XA.XIR[4].XIC[10].icell.Ien VGND 0.3733f
C4435 XA.XIR[4].XIC[9].icell.Ien VGND 0.3733f
C4436 XA.XIR[4].XIC[8].icell.Ien VGND 0.3733f
C4437 XA.XIR[4].XIC[7].icell.Ien VGND 0.3733f
C4438 XA.XIR[4].XIC[6].icell.Ien VGND 0.3733f
C4439 XA.XIR[4].XIC[5].icell.Ien VGND 0.3733f
C4440 XA.XIR[4].XIC[4].icell.Ien VGND 0.3733f
C4441 XA.XIR[4].XIC[3].icell.Ien VGND 0.3733f
C4442 XA.XIR[4].XIC[2].icell.Ien VGND 0.3733f
C4443 XA.XIR[4].XIC_dummy_left.icell.Iout VGND 0.80734f
C4444 XA.XIR[4].XIC[1].icell.Ien VGND 0.3733f
C4445 XA.XIR[4].XIC[0].icell.Ien VGND 0.37345f
C4446 XA.XIR[4].XIC_dummy_left.icell.SM VGND 0.01033f
C4447 XA.XIR[4].XIC_dummy_left.icell.Ien VGND 0.57333f
C4448 XA.XIR[4].XIC_dummy_right.icell.PDM VGND 0.23384f
C4449 XA.XIR[4].XIC_15.icell.PDM VGND 0.18862f
C4450 XA.XIR[4].XIC[14].icell.PDM VGND 0.1882f
C4451 XA.XIR[4].XIC[13].icell.PDM VGND 0.1882f
C4452 XA.XIR[4].XIC[12].icell.PDM VGND 0.1882f
C4453 XA.XIR[4].XIC[11].icell.PDM VGND 0.1882f
C4454 XA.XIR[4].XIC[10].icell.PDM VGND 0.1882f
C4455 XA.XIR[4].XIC[9].icell.PDM VGND 0.1882f
C4456 XA.XIR[4].XIC[8].icell.PDM VGND 0.1882f
C4457 XA.XIR[4].XIC[7].icell.PDM VGND 0.1882f
C4458 XA.XIR[4].XIC[6].icell.PDM VGND 0.1882f
C4459 XA.XIR[4].XIC[5].icell.PDM VGND 0.1882f
C4460 XA.XIR[4].XIC[4].icell.PDM VGND 0.1882f
C4461 XA.XIR[4].XIC[3].icell.PDM VGND 0.1882f
C4462 XA.XIR[4].XIC[2].icell.PDM VGND 0.1882f
C4463 XA.XIR[4].XIC[1].icell.PDM VGND 0.1882f
C4464 XA.XIR[4].XIC[0].icell.PDM VGND 0.18836f
C4465 XA.XIR[4].XIC_dummy_left.icell.PDM VGND 0.22809f
C4466 XThR.Tn[4] VGND 12.95212f
C4467 a_n1049_6405# VGND 0.02935f
C4468 XA.XIR[3].XIC_dummy_right.icell.Iout VGND 0.85788f
C4469 XA.XIR[3].XIC_dummy_right.icell.SM VGND 0.01013f
C4470 XA.XIR[3].XIC_dummy_right.icell.Ien VGND 0.60818f
C4471 XA.XIR[3].XIC_15.icell.Ien VGND 0.37264f
C4472 XA.XIR[3].XIC[14].icell.Ien VGND 0.37333f
C4473 XA.XIR[3].XIC[13].icell.Ien VGND 0.3733f
C4474 XA.XIR[3].XIC[12].icell.Ien VGND 0.3733f
C4475 XA.XIR[3].XIC[11].icell.Ien VGND 0.3733f
C4476 XA.XIR[3].XIC[10].icell.Ien VGND 0.3733f
C4477 XA.XIR[3].XIC[9].icell.Ien VGND 0.3733f
C4478 XA.XIR[3].XIC[8].icell.Ien VGND 0.3733f
C4479 XA.XIR[3].XIC[7].icell.Ien VGND 0.3733f
C4480 XA.XIR[3].XIC[6].icell.Ien VGND 0.3733f
C4481 XA.XIR[3].XIC[5].icell.Ien VGND 0.3733f
C4482 XA.XIR[3].XIC[4].icell.Ien VGND 0.3733f
C4483 XA.XIR[3].XIC[3].icell.Ien VGND 0.3733f
C4484 XA.XIR[3].XIC[2].icell.Ien VGND 0.3733f
C4485 XThR.XTB5.Y VGND 1.32753f
C4486 XA.XIR[3].XIC_dummy_left.icell.Iout VGND 0.80575f
C4487 XA.XIR[3].XIC[1].icell.Ien VGND 0.3733f
C4488 XA.XIR[3].XIC[0].icell.Ien VGND 0.37345f
C4489 XA.XIR[3].XIC_dummy_left.icell.SM VGND 0.01033f
C4490 XA.XIR[3].XIC_dummy_left.icell.Ien VGND 0.57422f
C4491 a_n1049_6699# VGND 0.02979f
C4492 XA.XIR[3].XIC_dummy_right.icell.PDM VGND 0.23384f
C4493 XA.XIR[3].XIC_15.icell.PDM VGND 0.18862f
C4494 XA.XIR[3].XIC[14].icell.PDM VGND 0.1882f
C4495 XA.XIR[3].XIC[13].icell.PDM VGND 0.1882f
C4496 XA.XIR[3].XIC[12].icell.PDM VGND 0.1882f
C4497 XA.XIR[3].XIC[11].icell.PDM VGND 0.1882f
C4498 XA.XIR[3].XIC[10].icell.PDM VGND 0.1882f
C4499 XA.XIR[3].XIC[9].icell.PDM VGND 0.1882f
C4500 XA.XIR[3].XIC[8].icell.PDM VGND 0.1882f
C4501 XA.XIR[3].XIC[7].icell.PDM VGND 0.1882f
C4502 XA.XIR[3].XIC[6].icell.PDM VGND 0.1882f
C4503 XA.XIR[3].XIC[5].icell.PDM VGND 0.1882f
C4504 XA.XIR[3].XIC[4].icell.PDM VGND 0.1882f
C4505 XA.XIR[3].XIC[3].icell.PDM VGND 0.1882f
C4506 XA.XIR[3].XIC[2].icell.PDM VGND 0.1882f
C4507 XA.XIR[3].XIC[1].icell.PDM VGND 0.1882f
C4508 XA.XIR[3].XIC[0].icell.PDM VGND 0.18836f
C4509 XA.XIR[3].XIC_dummy_left.icell.PDM VGND 0.22809f
C4510 XA.XIR[2].XIC_dummy_right.icell.Iout VGND 0.85788f
C4511 XA.XIR[2].XIC_dummy_right.icell.SM VGND 0.01013f
C4512 XA.XIR[2].XIC_dummy_right.icell.Ien VGND 0.60818f
C4513 XA.XIR[2].XIC_15.icell.Ien VGND 0.37264f
C4514 XA.XIR[2].XIC[14].icell.Ien VGND 0.37333f
C4515 XA.XIR[2].XIC[13].icell.Ien VGND 0.3733f
C4516 XA.XIR[2].XIC[12].icell.Ien VGND 0.3733f
C4517 XA.XIR[2].XIC[11].icell.Ien VGND 0.3733f
C4518 XA.XIR[2].XIC[10].icell.Ien VGND 0.3733f
C4519 XA.XIR[2].XIC[9].icell.Ien VGND 0.3733f
C4520 XA.XIR[2].XIC[8].icell.Ien VGND 0.3733f
C4521 XA.XIR[2].XIC[7].icell.Ien VGND 0.3733f
C4522 XA.XIR[2].XIC[6].icell.Ien VGND 0.3733f
C4523 XA.XIR[2].XIC[5].icell.Ien VGND 0.3733f
C4524 XA.XIR[2].XIC[4].icell.Ien VGND 0.3733f
C4525 XA.XIR[2].XIC[3].icell.Ien VGND 0.3733f
C4526 XA.XIR[2].XIC[2].icell.Ien VGND 0.3733f
C4527 XA.XIR[2].XIC_dummy_left.icell.Iout VGND 0.80789f
C4528 XA.XIR[2].XIC[1].icell.Ien VGND 0.3733f
C4529 XThR.Tn[3] VGND 12.94485f
C4530 XThR.XTB4.Y VGND 1.48815f
C4531 XA.XIR[2].XIC[0].icell.Ien VGND 0.37345f
C4532 XA.XIR[2].XIC_dummy_left.icell.SM VGND 0.01033f
C4533 XA.XIR[2].XIC_dummy_left.icell.Ien VGND 0.57556f
C4534 XA.XIR[2].XIC_dummy_right.icell.PDM VGND 0.23384f
C4535 XA.XIR[2].XIC_15.icell.PDM VGND 0.18862f
C4536 XA.XIR[2].XIC[14].icell.PDM VGND 0.1882f
C4537 XA.XIR[2].XIC[13].icell.PDM VGND 0.1882f
C4538 XA.XIR[2].XIC[12].icell.PDM VGND 0.1882f
C4539 XA.XIR[2].XIC[11].icell.PDM VGND 0.1882f
C4540 XA.XIR[2].XIC[10].icell.PDM VGND 0.1882f
C4541 XA.XIR[2].XIC[9].icell.PDM VGND 0.1882f
C4542 XA.XIR[2].XIC[8].icell.PDM VGND 0.1882f
C4543 XA.XIR[2].XIC[7].icell.PDM VGND 0.1882f
C4544 XA.XIR[2].XIC[6].icell.PDM VGND 0.1882f
C4545 XA.XIR[2].XIC[5].icell.PDM VGND 0.1882f
C4546 XA.XIR[2].XIC[4].icell.PDM VGND 0.1882f
C4547 XA.XIR[2].XIC[3].icell.PDM VGND 0.1882f
C4548 XA.XIR[2].XIC[2].icell.PDM VGND 0.1882f
C4549 XA.XIR[2].XIC[1].icell.PDM VGND 0.1882f
C4550 XA.XIR[2].XIC[0].icell.PDM VGND 0.18836f
C4551 XA.XIR[2].XIC_dummy_left.icell.PDM VGND 0.22809f
C4552 XA.XIR[1].XIC_dummy_right.icell.Iout VGND 0.85788f
C4553 XA.XIR[1].XIC_dummy_right.icell.SM VGND 0.01013f
C4554 XA.XIR[1].XIC_dummy_right.icell.Ien VGND 0.60818f
C4555 XA.XIR[1].XIC_15.icell.Ien VGND 0.37264f
C4556 XA.XIR[1].XIC[14].icell.Ien VGND 0.37333f
C4557 XA.XIR[1].XIC[13].icell.Ien VGND 0.3733f
C4558 XA.XIR[1].XIC[12].icell.Ien VGND 0.3733f
C4559 XA.XIR[1].XIC[11].icell.Ien VGND 0.3733f
C4560 XA.XIR[1].XIC[10].icell.Ien VGND 0.3733f
C4561 XA.XIR[1].XIC[9].icell.Ien VGND 0.3733f
C4562 XA.XIR[1].XIC[8].icell.Ien VGND 0.3733f
C4563 XA.XIR[1].XIC[7].icell.Ien VGND 0.3733f
C4564 XA.XIR[1].XIC[6].icell.Ien VGND 0.3733f
C4565 XA.XIR[1].XIC[5].icell.Ien VGND 0.3733f
C4566 XA.XIR[1].XIC[4].icell.Ien VGND 0.3733f
C4567 XA.XIR[1].XIC[3].icell.Ien VGND 0.3733f
C4568 XA.XIR[1].XIC[2].icell.Ien VGND 0.3733f
C4569 XA.XIR[1].XIC_dummy_left.icell.Iout VGND 0.80575f
C4570 XA.XIR[1].XIC[1].icell.Ien VGND 0.3733f
C4571 XThR.Tn[2] VGND 12.94933f
C4572 a_n1049_7493# VGND 0.02484f
C4573 XThR.XTB3.Y VGND 1.24035f
C4574 XThR.XTB7.A VGND 1.95537f
C4575 XA.XIR[1].XIC[0].icell.Ien VGND 0.37345f
C4576 XA.XIR[1].XIC_dummy_left.icell.SM VGND 0.01033f
C4577 XA.XIR[1].XIC_dummy_left.icell.Ien VGND 0.57376f
C4578 XA.XIR[1].XIC_dummy_right.icell.PDM VGND 0.23384f
C4579 XA.XIR[1].XIC_15.icell.PDM VGND 0.18862f
C4580 XA.XIR[1].XIC[14].icell.PDM VGND 0.1882f
C4581 XA.XIR[1].XIC[13].icell.PDM VGND 0.1882f
C4582 XA.XIR[1].XIC[12].icell.PDM VGND 0.1882f
C4583 XA.XIR[1].XIC[11].icell.PDM VGND 0.1882f
C4584 XA.XIR[1].XIC[10].icell.PDM VGND 0.1882f
C4585 XA.XIR[1].XIC[9].icell.PDM VGND 0.1882f
C4586 XA.XIR[1].XIC[8].icell.PDM VGND 0.1882f
C4587 XA.XIR[1].XIC[7].icell.PDM VGND 0.1882f
C4588 XA.XIR[1].XIC[6].icell.PDM VGND 0.1882f
C4589 XA.XIR[1].XIC[5].icell.PDM VGND 0.1882f
C4590 XA.XIR[1].XIC[4].icell.PDM VGND 0.1882f
C4591 XA.XIR[1].XIC[3].icell.PDM VGND 0.1882f
C4592 XA.XIR[1].XIC[2].icell.PDM VGND 0.1882f
C4593 XA.XIR[1].XIC[1].icell.PDM VGND 0.1882f
C4594 XA.XIR[1].XIC[0].icell.PDM VGND 0.18836f
C4595 XA.XIR[1].XIC_dummy_left.icell.PDM VGND 0.22809f
C4596 a_n1049_7787# VGND 0.03397f
C4597 XA.XIR[0].XIC_dummy_right.icell.Iout VGND 0.87403f
C4598 XA.XIR[0].XIC_dummy_right.icell.SM VGND 0.01013f
C4599 XA.XIR[0].XIC_dummy_right.icell.Ien VGND 0.61797f
C4600 XA.XIR[0].XIC_15.icell.Ien VGND 0.37874f
C4601 XA.XIR[0].XIC[14].icell.Ien VGND 0.39158f
C4602 XA.XIR[0].XIC[13].icell.Ien VGND 0.39155f
C4603 XA.XIR[0].XIC[12].icell.Ien VGND 0.38822f
C4604 XA.XIR[0].XIC[11].icell.Ien VGND 0.3889f
C4605 XA.XIR[0].XIC[10].icell.Ien VGND 0.39022f
C4606 XA.XIR[0].XIC[9].icell.Ien VGND 0.3885f
C4607 XA.XIR[0].XIC[8].icell.Ien VGND 0.38898f
C4608 XA.XIR[0].XIC[7].icell.Ien VGND 0.38927f
C4609 XA.XIR[0].XIC[6].icell.Ien VGND 0.38927f
C4610 XA.XIR[0].XIC[5].icell.Ien VGND 0.38822f
C4611 XA.XIR[0].XIC[4].icell.Ien VGND 0.38827f
C4612 XA.XIR[0].XIC[3].icell.Ien VGND 0.38951f
C4613 XA.XIR[0].XIC[2].icell.Ien VGND 0.39155f
C4614 XA.XIR[0].XIC_dummy_left.icell.Iout VGND 0.83191f
C4615 XA.XIR[0].XIC[1].icell.Ien VGND 0.39155f
C4616 XA.XIR[0].XIC[0].icell.Ien VGND 0.39086f
C4617 XA.XIR[0].XIC_dummy_left.icell.SM VGND 0.01033f
C4618 XThR.Tn[1] VGND 12.98843f
C4619 XThR.XTB2.Y VGND 1.47619f
C4620 XThR.XTB6.A VGND 0.95635f
C4621 XA.XIR[0].XIC_dummy_left.icell.Ien VGND 0.58431f
C4622 XA.XIR[0].XIC_dummy_right.icell.PDM VGND 0.251f
C4623 XA.XIR[0].XIC_15.icell.PDM VGND 0.20773f
C4624 XA.XIR[0].XIC[14].icell.PDM VGND 0.24601f
C4625 XA.XIR[0].XIC[13].icell.PDM VGND 0.24585f
C4626 XA.XIR[0].XIC[12].icell.PDM VGND 0.24146f
C4627 XA.XIR[0].XIC[11].icell.PDM VGND 0.24184f
C4628 XA.XIR[0].XIC[10].icell.PDM VGND 0.24174f
C4629 XA.XIR[0].XIC[9].icell.PDM VGND 0.24147f
C4630 XA.XIR[0].XIC[8].icell.PDM VGND 0.24147f
C4631 XA.XIR[0].XIC[7].icell.PDM VGND 0.2442f
C4632 XA.XIR[0].XIC[6].icell.PDM VGND 0.24156f
C4633 XA.XIR[0].XIC[5].icell.PDM VGND 0.24321f
C4634 XA.XIR[0].XIC[4].icell.PDM VGND 0.24159f
C4635 XA.XIR[0].XIC[3].icell.PDM VGND 0.24451f
C4636 XA.XIR[0].XIC[2].icell.PDM VGND 0.2458f
C4637 XA.XIR[0].XIC[1].icell.PDM VGND 0.2458f
C4638 XA.XIR[0].XIC[0].icell.PDM VGND 0.2446f
C4639 XA.XIR[0].XIC_dummy_left.icell.PDM VGND 0.24577f
C4640 XThR.Tn[0] VGND 13.29619f
C4641 a_n1049_8581# VGND 0.04333f
C4642 XThR.XTBN.Y VGND 7.77803f
C4643 XThR.XTB1.Y VGND 1.45322f
C4644 XThR.XTB7.B VGND 2.61063f
C4645 XThR.XTB5.A VGND 1.75777f
C4646 XThC.Tn[14] VGND 5.52615f
C4647 XThC.Tn[13] VGND 5.16689f
C4648 XThC.Tn[12] VGND 5.1562f
C4649 XThC.Tn[11] VGND 5.52379f
C4650 XThC.Tn[10] VGND 5.0515f
C4651 XThC.Tn[9] VGND 5.34336f
C4652 XThC.Tn[8] VGND 4.89287f
C4653 a_10915_9569# VGND 0.55912f
C4654 a_10051_9569# VGND 0.55747f
C4655 a_9827_9569# VGND 0.54584f
C4656 a_8963_9569# VGND 0.55439f
C4657 a_8739_9569# VGND 0.553f
C4658 a_7875_9569# VGND 0.55432f
C4659 a_7651_9569# VGND 0.55717f
C4660 XThC.Tn[7] VGND 5.47379f
C4661 XThC.Tn[6] VGND 5.48958f
C4662 XThC.Tn[5] VGND 5.60438f
C4663 XThC.Tn[4] VGND 5.55465f
C4664 XThC.Tn[3] VGND 5.88113f
C4665 XThC.Tn[2] VGND 5.58437f
C4666 XThC.Tn[1] VGND 5.71923f
C4667 XThC.Tn[0] VGND 6.86777f
C4668 a_6243_9615# VGND 0.03028f
C4669 a_5949_9615# VGND 0.03456f
C4670 a_5155_9615# VGND 0.03624f
C4671 a_4861_9615# VGND 0.03647f
C4672 a_4067_9615# VGND 0.03118f
C4673 a_3773_9615# VGND 0.03896f
C4674 a_2979_9615# VGND 0.04122f
C4675 XThC.XTBN.Y VGND 8.71711f
C4676 XThC.XTB7.Y VGND 1.35988f
C4677 XThC.XTB6.Y VGND 1.3794f
C4678 XThC.XTB7.B VGND 2.83799f
C4679 XThC.XTB5.Y VGND 1.32558f
C4680 XThC.XTBN.A VGND 1.2246f
C4681 XThC.XTB4.Y VGND 1.6934f
C4682 XThC.XTB3.Y VGND 1.96717f
C4683 XThC.XTB7.A VGND 1.94951f
C4684 XThC.XTB6.A VGND 0.95452f
C4685 XThC.XTB2.Y VGND 1.4752f
C4686 XThC.XTB1.Y VGND 1.77643f
C4687 XThC.XTB5.A VGND 1.75974f
C4688 bias[0].t0 VGND 0.94587f
C4689 XThR.Tn[13].t2 VGND 0.01241f
C4690 XThR.Tn[13].t0 VGND 0.01241f
C4691 XThR.Tn[13].n0 VGND 0.02481f
C4692 XThR.Tn[13].t3 VGND 0.01241f
C4693 XThR.Tn[13].t1 VGND 0.01241f
C4694 XThR.Tn[13].n1 VGND 0.03094f
C4695 XThR.Tn[13].n2 VGND 0.06242f
C4696 XThR.Tn[13].t9 VGND 0.01909f
C4697 XThR.Tn[13].t11 VGND 0.01909f
C4698 XThR.Tn[13].n3 VGND 0.05796f
C4699 XThR.Tn[13].t10 VGND 0.01909f
C4700 XThR.Tn[13].t8 VGND 0.01909f
C4701 XThR.Tn[13].n4 VGND 0.04243f
C4702 XThR.Tn[13].n5 VGND 0.19293f
C4703 XThR.Tn[13].t6 VGND 0.01909f
C4704 XThR.Tn[13].t4 VGND 0.01909f
C4705 XThR.Tn[13].n6 VGND 0.04124f
C4706 XThR.Tn[13].t7 VGND 0.01909f
C4707 XThR.Tn[13].t5 VGND 0.01909f
C4708 XThR.Tn[13].n7 VGND 0.06277f
C4709 XThR.Tn[13].n8 VGND 0.17429f
C4710 XThR.Tn[13].n9 VGND 0.02334f
C4711 XThR.Tn[13].t72 VGND 0.01492f
C4712 XThR.Tn[13].t64 VGND 0.01633f
C4713 XThR.Tn[13].n10 VGND 0.03989f
C4714 XThR.Tn[13].n11 VGND 0.07663f
C4715 XThR.Tn[13].t28 VGND 0.01492f
C4716 XThR.Tn[13].t21 VGND 0.01633f
C4717 XThR.Tn[13].n12 VGND 0.03989f
C4718 XThR.Tn[13].t44 VGND 0.01487f
C4719 XThR.Tn[13].t12 VGND 0.01628f
C4720 XThR.Tn[13].n13 VGND 0.0415f
C4721 XThR.Tn[13].n14 VGND 0.02916f
C4722 XThR.Tn[13].n16 VGND 0.09357f
C4723 XThR.Tn[13].t65 VGND 0.01492f
C4724 XThR.Tn[13].t57 VGND 0.01633f
C4725 XThR.Tn[13].n17 VGND 0.03989f
C4726 XThR.Tn[13].t19 VGND 0.01487f
C4727 XThR.Tn[13].t52 VGND 0.01628f
C4728 XThR.Tn[13].n18 VGND 0.0415f
C4729 XThR.Tn[13].n19 VGND 0.02916f
C4730 XThR.Tn[13].n21 VGND 0.09357f
C4731 XThR.Tn[13].t22 VGND 0.01492f
C4732 XThR.Tn[13].t14 VGND 0.01633f
C4733 XThR.Tn[13].n22 VGND 0.03989f
C4734 XThR.Tn[13].t34 VGND 0.01487f
C4735 XThR.Tn[13].t70 VGND 0.01628f
C4736 XThR.Tn[13].n23 VGND 0.0415f
C4737 XThR.Tn[13].n24 VGND 0.02916f
C4738 XThR.Tn[13].n26 VGND 0.09357f
C4739 XThR.Tn[13].t49 VGND 0.01492f
C4740 XThR.Tn[13].t39 VGND 0.01633f
C4741 XThR.Tn[13].n27 VGND 0.03989f
C4742 XThR.Tn[13].t66 VGND 0.01487f
C4743 XThR.Tn[13].t35 VGND 0.01628f
C4744 XThR.Tn[13].n28 VGND 0.0415f
C4745 XThR.Tn[13].n29 VGND 0.02916f
C4746 XThR.Tn[13].n31 VGND 0.09357f
C4747 XThR.Tn[13].t24 VGND 0.01492f
C4748 XThR.Tn[13].t16 VGND 0.01633f
C4749 XThR.Tn[13].n32 VGND 0.03989f
C4750 XThR.Tn[13].t37 VGND 0.01487f
C4751 XThR.Tn[13].t71 VGND 0.01628f
C4752 XThR.Tn[13].n33 VGND 0.0415f
C4753 XThR.Tn[13].n34 VGND 0.02916f
C4754 XThR.Tn[13].n36 VGND 0.09357f
C4755 XThR.Tn[13].t60 VGND 0.01492f
C4756 XThR.Tn[13].t30 VGND 0.01633f
C4757 XThR.Tn[13].n37 VGND 0.03989f
C4758 XThR.Tn[13].t13 VGND 0.01487f
C4759 XThR.Tn[13].t26 VGND 0.01628f
C4760 XThR.Tn[13].n38 VGND 0.0415f
C4761 XThR.Tn[13].n39 VGND 0.02916f
C4762 XThR.Tn[13].n41 VGND 0.09357f
C4763 XThR.Tn[13].t29 VGND 0.01492f
C4764 XThR.Tn[13].t25 VGND 0.01633f
C4765 XThR.Tn[13].n42 VGND 0.03989f
C4766 XThR.Tn[13].t43 VGND 0.01487f
C4767 XThR.Tn[13].t18 VGND 0.01628f
C4768 XThR.Tn[13].n43 VGND 0.0415f
C4769 XThR.Tn[13].n44 VGND 0.02916f
C4770 XThR.Tn[13].n46 VGND 0.09357f
C4771 XThR.Tn[13].t32 VGND 0.01492f
C4772 XThR.Tn[13].t38 VGND 0.01633f
C4773 XThR.Tn[13].n47 VGND 0.03989f
C4774 XThR.Tn[13].t48 VGND 0.01487f
C4775 XThR.Tn[13].t33 VGND 0.01628f
C4776 XThR.Tn[13].n48 VGND 0.0415f
C4777 XThR.Tn[13].n49 VGND 0.02916f
C4778 XThR.Tn[13].n51 VGND 0.09357f
C4779 XThR.Tn[13].t51 VGND 0.01492f
C4780 XThR.Tn[13].t59 VGND 0.01633f
C4781 XThR.Tn[13].n52 VGND 0.03989f
C4782 XThR.Tn[13].t68 VGND 0.01487f
C4783 XThR.Tn[13].t53 VGND 0.01628f
C4784 XThR.Tn[13].n53 VGND 0.0415f
C4785 XThR.Tn[13].n54 VGND 0.02916f
C4786 XThR.Tn[13].n56 VGND 0.09357f
C4787 XThR.Tn[13].t41 VGND 0.01492f
C4788 XThR.Tn[13].t17 VGND 0.01633f
C4789 XThR.Tn[13].n57 VGND 0.03989f
C4790 XThR.Tn[13].t58 VGND 0.01487f
C4791 XThR.Tn[13].t73 VGND 0.01628f
C4792 XThR.Tn[13].n58 VGND 0.0415f
C4793 XThR.Tn[13].n59 VGND 0.02916f
C4794 XThR.Tn[13].n61 VGND 0.09357f
C4795 XThR.Tn[13].t63 VGND 0.01492f
C4796 XThR.Tn[13].t55 VGND 0.01633f
C4797 XThR.Tn[13].n62 VGND 0.03989f
C4798 XThR.Tn[13].t15 VGND 0.01487f
C4799 XThR.Tn[13].t45 VGND 0.01628f
C4800 XThR.Tn[13].n63 VGND 0.0415f
C4801 XThR.Tn[13].n64 VGND 0.02916f
C4802 XThR.Tn[13].n66 VGND 0.09357f
C4803 XThR.Tn[13].t31 VGND 0.01492f
C4804 XThR.Tn[13].t27 VGND 0.01633f
C4805 XThR.Tn[13].n67 VGND 0.03989f
C4806 XThR.Tn[13].t46 VGND 0.01487f
C4807 XThR.Tn[13].t20 VGND 0.01628f
C4808 XThR.Tn[13].n68 VGND 0.0415f
C4809 XThR.Tn[13].n69 VGND 0.02916f
C4810 XThR.Tn[13].n71 VGND 0.09357f
C4811 XThR.Tn[13].t50 VGND 0.01492f
C4812 XThR.Tn[13].t40 VGND 0.01633f
C4813 XThR.Tn[13].n72 VGND 0.03989f
C4814 XThR.Tn[13].t67 VGND 0.01487f
C4815 XThR.Tn[13].t36 VGND 0.01628f
C4816 XThR.Tn[13].n73 VGND 0.0415f
C4817 XThR.Tn[13].n74 VGND 0.02916f
C4818 XThR.Tn[13].n76 VGND 0.09357f
C4819 XThR.Tn[13].t69 VGND 0.01492f
C4820 XThR.Tn[13].t62 VGND 0.01633f
C4821 XThR.Tn[13].n77 VGND 0.03989f
C4822 XThR.Tn[13].t23 VGND 0.01487f
C4823 XThR.Tn[13].t54 VGND 0.01628f
C4824 XThR.Tn[13].n78 VGND 0.0415f
C4825 XThR.Tn[13].n79 VGND 0.02916f
C4826 XThR.Tn[13].n81 VGND 0.09357f
C4827 XThR.Tn[13].t42 VGND 0.01492f
C4828 XThR.Tn[13].t56 VGND 0.01633f
C4829 XThR.Tn[13].n82 VGND 0.03989f
C4830 XThR.Tn[13].t61 VGND 0.01487f
C4831 XThR.Tn[13].t47 VGND 0.01628f
C4832 XThR.Tn[13].n83 VGND 0.0415f
C4833 XThR.Tn[13].n84 VGND 0.02916f
C4834 XThR.Tn[13].n86 VGND 0.09357f
C4835 XThR.Tn[13].n87 VGND 0.08503f
C4836 XThR.Tn[13].n88 VGND 0.33338f
C4837 XThC.XTB3.Y.t1 VGND 0.06296f
C4838 XThC.XTB3.Y.n0 VGND 0.04069f
C4839 XThC.XTB3.Y.n1 VGND 0.05192f
C4840 XThC.XTB3.Y.t2 VGND 0.03159f
C4841 XThC.XTB3.Y.t0 VGND 0.03159f
C4842 XThC.XTB3.Y.n2 VGND 0.06782f
C4843 XThC.XTB3.Y.t10 VGND 0.04914f
C4844 XThC.XTB3.Y.t17 VGND 0.02896f
C4845 XThC.XTB3.Y.n3 VGND 0.05852f
C4846 XThC.XTB3.Y.t14 VGND 0.04914f
C4847 XThC.XTB3.Y.t5 VGND 0.02896f
C4848 XThC.XTB3.Y.n4 VGND 0.03012f
C4849 XThC.XTB3.Y.t15 VGND 0.04914f
C4850 XThC.XTB3.Y.t6 VGND 0.02896f
C4851 XThC.XTB3.Y.n5 VGND 0.06469f
C4852 XThC.XTB3.Y.t3 VGND 0.04914f
C4853 XThC.XTB3.Y.t9 VGND 0.02896f
C4854 XThC.XTB3.Y.n6 VGND 0.06006f
C4855 XThC.XTB3.Y.n7 VGND 0.03654f
C4856 XThC.XTB3.Y.n8 VGND 0.06049f
C4857 XThC.XTB3.Y.n9 VGND 0.0234f
C4858 XThC.XTB3.Y.n10 VGND 0.02857f
C4859 XThC.XTB3.Y.n11 VGND 0.06469f
C4860 XThC.XTB3.Y.n12 VGND 0.03243f
C4861 XThC.XTB3.Y.n13 VGND 0.05514f
C4862 XThC.XTB3.Y.t16 VGND 0.04914f
C4863 XThC.XTB3.Y.t7 VGND 0.02896f
C4864 XThC.XTB3.Y.n14 VGND 0.06624f
C4865 XThC.XTB3.Y.t4 VGND 0.04914f
C4866 XThC.XTB3.Y.t13 VGND 0.02896f
C4867 XThC.XTB3.Y.t12 VGND 0.04914f
C4868 XThC.XTB3.Y.t18 VGND 0.02896f
C4869 XThC.XTB3.Y.t11 VGND 0.04914f
C4870 XThC.XTB3.Y.t8 VGND 0.02896f
C4871 XThC.XTB3.Y.n15 VGND 0.08245f
C4872 XThC.XTB3.Y.n16 VGND 0.08709f
C4873 XThC.XTB3.Y.n17 VGND 0.03356f
C4874 XThC.XTB3.Y.n18 VGND 0.07087f
C4875 XThC.XTB3.Y.n19 VGND 0.03243f
C4876 XThC.XTB3.Y.n20 VGND 0.02691f
C4877 XThC.XTB3.Y.n21 VGND 1.39635f
C4878 XThC.XTB3.Y.n22 VGND 0.14933f
C4879 XThR.Tn[8].t10 VGND 0.01919f
C4880 XThR.Tn[8].t8 VGND 0.01919f
C4881 XThR.Tn[8].n0 VGND 0.05828f
C4882 XThR.Tn[8].t11 VGND 0.01919f
C4883 XThR.Tn[8].t9 VGND 0.01919f
C4884 XThR.Tn[8].n1 VGND 0.04267f
C4885 XThR.Tn[8].n2 VGND 0.19401f
C4886 XThR.Tn[8].t6 VGND 0.01919f
C4887 XThR.Tn[8].t4 VGND 0.01919f
C4888 XThR.Tn[8].n3 VGND 0.04147f
C4889 XThR.Tn[8].t7 VGND 0.01919f
C4890 XThR.Tn[8].t5 VGND 0.01919f
C4891 XThR.Tn[8].n4 VGND 0.06312f
C4892 XThR.Tn[8].n5 VGND 0.17526f
C4893 XThR.Tn[8].t39 VGND 0.015f
C4894 XThR.Tn[8].t33 VGND 0.01643f
C4895 XThR.Tn[8].n7 VGND 0.04011f
C4896 XThR.Tn[8].n8 VGND 0.07706f
C4897 XThR.Tn[8].t59 VGND 0.015f
C4898 XThR.Tn[8].t49 VGND 0.01643f
C4899 XThR.Tn[8].n9 VGND 0.04011f
C4900 XThR.Tn[8].t13 VGND 0.01495f
C4901 XThR.Tn[8].t45 VGND 0.01637f
C4902 XThR.Tn[8].n10 VGND 0.04174f
C4903 XThR.Tn[8].n11 VGND 0.02932f
C4904 XThR.Tn[8].n13 VGND 0.09409f
C4905 XThR.Tn[8].t34 VGND 0.015f
C4906 XThR.Tn[8].t26 VGND 0.01643f
C4907 XThR.Tn[8].n14 VGND 0.04011f
C4908 XThR.Tn[8].t53 VGND 0.01495f
C4909 XThR.Tn[8].t22 VGND 0.01637f
C4910 XThR.Tn[8].n15 VGND 0.04174f
C4911 XThR.Tn[8].n16 VGND 0.02932f
C4912 XThR.Tn[8].n18 VGND 0.09409f
C4913 XThR.Tn[8].t50 VGND 0.015f
C4914 XThR.Tn[8].t43 VGND 0.01643f
C4915 XThR.Tn[8].n19 VGND 0.04011f
C4916 XThR.Tn[8].t65 VGND 0.01495f
C4917 XThR.Tn[8].t40 VGND 0.01637f
C4918 XThR.Tn[8].n20 VGND 0.04174f
C4919 XThR.Tn[8].n21 VGND 0.02932f
C4920 XThR.Tn[8].n23 VGND 0.09409f
C4921 XThR.Tn[8].t12 VGND 0.015f
C4922 XThR.Tn[8].t70 VGND 0.01643f
C4923 XThR.Tn[8].n24 VGND 0.04011f
C4924 XThR.Tn[8].t36 VGND 0.01495f
C4925 XThR.Tn[8].t66 VGND 0.01637f
C4926 XThR.Tn[8].n25 VGND 0.04174f
C4927 XThR.Tn[8].n26 VGND 0.02932f
C4928 XThR.Tn[8].n28 VGND 0.09409f
C4929 XThR.Tn[8].t52 VGND 0.015f
C4930 XThR.Tn[8].t44 VGND 0.01643f
C4931 XThR.Tn[8].n29 VGND 0.04011f
C4932 XThR.Tn[8].t68 VGND 0.01495f
C4933 XThR.Tn[8].t41 VGND 0.01637f
C4934 XThR.Tn[8].n30 VGND 0.04174f
C4935 XThR.Tn[8].n31 VGND 0.02932f
C4936 XThR.Tn[8].n33 VGND 0.09409f
C4937 XThR.Tn[8].t28 VGND 0.015f
C4938 XThR.Tn[8].t61 VGND 0.01643f
C4939 XThR.Tn[8].n34 VGND 0.04011f
C4940 XThR.Tn[8].t47 VGND 0.01495f
C4941 XThR.Tn[8].t58 VGND 0.01637f
C4942 XThR.Tn[8].n35 VGND 0.04174f
C4943 XThR.Tn[8].n36 VGND 0.02932f
C4944 XThR.Tn[8].n38 VGND 0.09409f
C4945 XThR.Tn[8].t60 VGND 0.015f
C4946 XThR.Tn[8].t56 VGND 0.01643f
C4947 XThR.Tn[8].n39 VGND 0.04011f
C4948 XThR.Tn[8].t14 VGND 0.01495f
C4949 XThR.Tn[8].t51 VGND 0.01637f
C4950 XThR.Tn[8].n40 VGND 0.04174f
C4951 XThR.Tn[8].n41 VGND 0.02932f
C4952 XThR.Tn[8].n43 VGND 0.09409f
C4953 XThR.Tn[8].t63 VGND 0.015f
C4954 XThR.Tn[8].t69 VGND 0.01643f
C4955 XThR.Tn[8].n44 VGND 0.04011f
C4956 XThR.Tn[8].t20 VGND 0.01495f
C4957 XThR.Tn[8].t64 VGND 0.01637f
C4958 XThR.Tn[8].n45 VGND 0.04174f
C4959 XThR.Tn[8].n46 VGND 0.02932f
C4960 XThR.Tn[8].n48 VGND 0.09409f
C4961 XThR.Tn[8].t17 VGND 0.015f
C4962 XThR.Tn[8].t27 VGND 0.01643f
C4963 XThR.Tn[8].n49 VGND 0.04011f
C4964 XThR.Tn[8].t38 VGND 0.01495f
C4965 XThR.Tn[8].t24 VGND 0.01637f
C4966 XThR.Tn[8].n50 VGND 0.04174f
C4967 XThR.Tn[8].n51 VGND 0.02932f
C4968 XThR.Tn[8].n53 VGND 0.09409f
C4969 XThR.Tn[8].t72 VGND 0.015f
C4970 XThR.Tn[8].t46 VGND 0.01643f
C4971 XThR.Tn[8].n54 VGND 0.04011f
C4972 XThR.Tn[8].t31 VGND 0.01495f
C4973 XThR.Tn[8].t42 VGND 0.01637f
C4974 XThR.Tn[8].n55 VGND 0.04174f
C4975 XThR.Tn[8].n56 VGND 0.02932f
C4976 XThR.Tn[8].n58 VGND 0.09409f
C4977 XThR.Tn[8].t30 VGND 0.015f
C4978 XThR.Tn[8].t21 VGND 0.01643f
C4979 XThR.Tn[8].n59 VGND 0.04011f
C4980 XThR.Tn[8].t48 VGND 0.01495f
C4981 XThR.Tn[8].t16 VGND 0.01637f
C4982 XThR.Tn[8].n60 VGND 0.04174f
C4983 XThR.Tn[8].n61 VGND 0.02932f
C4984 XThR.Tn[8].n63 VGND 0.09409f
C4985 XThR.Tn[8].t62 VGND 0.015f
C4986 XThR.Tn[8].t57 VGND 0.01643f
C4987 XThR.Tn[8].n64 VGND 0.04011f
C4988 XThR.Tn[8].t18 VGND 0.01495f
C4989 XThR.Tn[8].t54 VGND 0.01637f
C4990 XThR.Tn[8].n65 VGND 0.04174f
C4991 XThR.Tn[8].n66 VGND 0.02932f
C4992 XThR.Tn[8].n68 VGND 0.09409f
C4993 XThR.Tn[8].t15 VGND 0.015f
C4994 XThR.Tn[8].t71 VGND 0.01643f
C4995 XThR.Tn[8].n69 VGND 0.04011f
C4996 XThR.Tn[8].t37 VGND 0.01495f
C4997 XThR.Tn[8].t67 VGND 0.01637f
C4998 XThR.Tn[8].n70 VGND 0.04174f
C4999 XThR.Tn[8].n71 VGND 0.02932f
C5000 XThR.Tn[8].n73 VGND 0.09409f
C5001 XThR.Tn[8].t35 VGND 0.015f
C5002 XThR.Tn[8].t29 VGND 0.01643f
C5003 XThR.Tn[8].n74 VGND 0.04011f
C5004 XThR.Tn[8].t55 VGND 0.01495f
C5005 XThR.Tn[8].t25 VGND 0.01637f
C5006 XThR.Tn[8].n75 VGND 0.04174f
C5007 XThR.Tn[8].n76 VGND 0.02932f
C5008 XThR.Tn[8].n78 VGND 0.09409f
C5009 XThR.Tn[8].t73 VGND 0.015f
C5010 XThR.Tn[8].t23 VGND 0.01643f
C5011 XThR.Tn[8].n79 VGND 0.04011f
C5012 XThR.Tn[8].t32 VGND 0.01495f
C5013 XThR.Tn[8].t19 VGND 0.01637f
C5014 XThR.Tn[8].n80 VGND 0.04174f
C5015 XThR.Tn[8].n81 VGND 0.02932f
C5016 XThR.Tn[8].n83 VGND 0.09409f
C5017 XThR.Tn[8].n84 VGND 0.08551f
C5018 XThR.Tn[8].n85 VGND 0.26201f
C5019 XThR.Tn[8].t0 VGND 0.01248f
C5020 XThR.Tn[8].t2 VGND 0.01248f
C5021 XThR.Tn[8].n86 VGND 0.02495f
C5022 XThR.Tn[8].t1 VGND 0.01248f
C5023 XThR.Tn[8].t3 VGND 0.01248f
C5024 XThR.Tn[8].n87 VGND 0.03112f
C5025 XThR.Tn[8].n88 VGND 0.05754f
C5026 XThR.Tn[0].t6 VGND 0.01769f
C5027 XThR.Tn[0].t7 VGND 0.01769f
C5028 XThR.Tn[0].n0 VGND 0.03571f
C5029 XThR.Tn[0].t5 VGND 0.01769f
C5030 XThR.Tn[0].t4 VGND 0.01769f
C5031 XThR.Tn[0].n1 VGND 0.04178f
C5032 XThR.Tn[0].n2 VGND 0.12532f
C5033 XThR.Tn[0].t9 VGND 0.0115f
C5034 XThR.Tn[0].t10 VGND 0.0115f
C5035 XThR.Tn[0].n3 VGND 0.02618f
C5036 XThR.Tn[0].t8 VGND 0.0115f
C5037 XThR.Tn[0].t11 VGND 0.0115f
C5038 XThR.Tn[0].n4 VGND 0.02618f
C5039 XThR.Tn[0].t1 VGND 0.0115f
C5040 XThR.Tn[0].t2 VGND 0.0115f
C5041 XThR.Tn[0].n5 VGND 0.04363f
C5042 XThR.Tn[0].t0 VGND 0.0115f
C5043 XThR.Tn[0].t3 VGND 0.0115f
C5044 XThR.Tn[0].n6 VGND 0.02618f
C5045 XThR.Tn[0].n7 VGND 0.12469f
C5046 XThR.Tn[0].n8 VGND 0.07708f
C5047 XThR.Tn[0].n9 VGND 0.08699f
C5048 XThR.Tn[0].t48 VGND 0.01383f
C5049 XThR.Tn[0].t40 VGND 0.01514f
C5050 XThR.Tn[0].n10 VGND 0.03697f
C5051 XThR.Tn[0].n11 VGND 0.07101f
C5052 XThR.Tn[0].t67 VGND 0.01383f
C5053 XThR.Tn[0].t58 VGND 0.01514f
C5054 XThR.Tn[0].n12 VGND 0.03697f
C5055 XThR.Tn[0].t24 VGND 0.01378f
C5056 XThR.Tn[0].t50 VGND 0.01509f
C5057 XThR.Tn[0].n13 VGND 0.03846f
C5058 XThR.Tn[0].n14 VGND 0.02702f
C5059 XThR.Tn[0].n16 VGND 0.08671f
C5060 XThR.Tn[0].t41 VGND 0.01383f
C5061 XThR.Tn[0].t33 VGND 0.01514f
C5062 XThR.Tn[0].n17 VGND 0.03697f
C5063 XThR.Tn[0].t61 VGND 0.01378f
C5064 XThR.Tn[0].t26 VGND 0.01509f
C5065 XThR.Tn[0].n18 VGND 0.03846f
C5066 XThR.Tn[0].n19 VGND 0.02702f
C5067 XThR.Tn[0].n21 VGND 0.08671f
C5068 XThR.Tn[0].t59 VGND 0.01383f
C5069 XThR.Tn[0].t51 VGND 0.01514f
C5070 XThR.Tn[0].n22 VGND 0.03697f
C5071 XThR.Tn[0].t12 VGND 0.01378f
C5072 XThR.Tn[0].t44 VGND 0.01509f
C5073 XThR.Tn[0].n23 VGND 0.03846f
C5074 XThR.Tn[0].n24 VGND 0.02702f
C5075 XThR.Tn[0].n26 VGND 0.08671f
C5076 XThR.Tn[0].t21 VGND 0.01383f
C5077 XThR.Tn[0].t15 VGND 0.01514f
C5078 XThR.Tn[0].n27 VGND 0.03697f
C5079 XThR.Tn[0].t43 VGND 0.01378f
C5080 XThR.Tn[0].t72 VGND 0.01509f
C5081 XThR.Tn[0].n28 VGND 0.03846f
C5082 XThR.Tn[0].n29 VGND 0.02702f
C5083 XThR.Tn[0].n31 VGND 0.08671f
C5084 XThR.Tn[0].t60 VGND 0.01383f
C5085 XThR.Tn[0].t52 VGND 0.01514f
C5086 XThR.Tn[0].n32 VGND 0.03697f
C5087 XThR.Tn[0].t13 VGND 0.01378f
C5088 XThR.Tn[0].t46 VGND 0.01509f
C5089 XThR.Tn[0].n33 VGND 0.03846f
C5090 XThR.Tn[0].n34 VGND 0.02702f
C5091 XThR.Tn[0].n36 VGND 0.08671f
C5092 XThR.Tn[0].t35 VGND 0.01383f
C5093 XThR.Tn[0].t68 VGND 0.01514f
C5094 XThR.Tn[0].n37 VGND 0.03697f
C5095 XThR.Tn[0].t54 VGND 0.01378f
C5096 XThR.Tn[0].t64 VGND 0.01509f
C5097 XThR.Tn[0].n38 VGND 0.03846f
C5098 XThR.Tn[0].n39 VGND 0.02702f
C5099 XThR.Tn[0].n41 VGND 0.08671f
C5100 XThR.Tn[0].t66 VGND 0.01383f
C5101 XThR.Tn[0].t63 VGND 0.01514f
C5102 XThR.Tn[0].n42 VGND 0.03697f
C5103 XThR.Tn[0].t23 VGND 0.01378f
C5104 XThR.Tn[0].t55 VGND 0.01509f
C5105 XThR.Tn[0].n43 VGND 0.03846f
C5106 XThR.Tn[0].n44 VGND 0.02702f
C5107 XThR.Tn[0].n46 VGND 0.08671f
C5108 XThR.Tn[0].t70 VGND 0.01383f
C5109 XThR.Tn[0].t14 VGND 0.01514f
C5110 XThR.Tn[0].n47 VGND 0.03697f
C5111 XThR.Tn[0].t28 VGND 0.01378f
C5112 XThR.Tn[0].t71 VGND 0.01509f
C5113 XThR.Tn[0].n48 VGND 0.03846f
C5114 XThR.Tn[0].n49 VGND 0.02702f
C5115 XThR.Tn[0].n51 VGND 0.08671f
C5116 XThR.Tn[0].t25 VGND 0.01383f
C5117 XThR.Tn[0].t34 VGND 0.01514f
C5118 XThR.Tn[0].n52 VGND 0.03697f
C5119 XThR.Tn[0].t47 VGND 0.01378f
C5120 XThR.Tn[0].t29 VGND 0.01509f
C5121 XThR.Tn[0].n53 VGND 0.03846f
C5122 XThR.Tn[0].n54 VGND 0.02702f
C5123 XThR.Tn[0].n56 VGND 0.08671f
C5124 XThR.Tn[0].t17 VGND 0.01383f
C5125 XThR.Tn[0].t53 VGND 0.01514f
C5126 XThR.Tn[0].n57 VGND 0.03697f
C5127 XThR.Tn[0].t38 VGND 0.01378f
C5128 XThR.Tn[0].t49 VGND 0.01509f
C5129 XThR.Tn[0].n58 VGND 0.03846f
C5130 XThR.Tn[0].n59 VGND 0.02702f
C5131 XThR.Tn[0].n61 VGND 0.08671f
C5132 XThR.Tn[0].t37 VGND 0.01383f
C5133 XThR.Tn[0].t31 VGND 0.01514f
C5134 XThR.Tn[0].n62 VGND 0.03697f
C5135 XThR.Tn[0].t56 VGND 0.01378f
C5136 XThR.Tn[0].t19 VGND 0.01509f
C5137 XThR.Tn[0].n63 VGND 0.03846f
C5138 XThR.Tn[0].n64 VGND 0.02702f
C5139 XThR.Tn[0].n66 VGND 0.08671f
C5140 XThR.Tn[0].t69 VGND 0.01383f
C5141 XThR.Tn[0].t65 VGND 0.01514f
C5142 XThR.Tn[0].n67 VGND 0.03697f
C5143 XThR.Tn[0].t27 VGND 0.01378f
C5144 XThR.Tn[0].t57 VGND 0.01509f
C5145 XThR.Tn[0].n68 VGND 0.03846f
C5146 XThR.Tn[0].n69 VGND 0.02702f
C5147 XThR.Tn[0].n71 VGND 0.08671f
C5148 XThR.Tn[0].t22 VGND 0.01383f
C5149 XThR.Tn[0].t16 VGND 0.01514f
C5150 XThR.Tn[0].n72 VGND 0.03697f
C5151 XThR.Tn[0].t45 VGND 0.01378f
C5152 XThR.Tn[0].t73 VGND 0.01509f
C5153 XThR.Tn[0].n73 VGND 0.03846f
C5154 XThR.Tn[0].n74 VGND 0.02702f
C5155 XThR.Tn[0].n76 VGND 0.08671f
C5156 XThR.Tn[0].t42 VGND 0.01383f
C5157 XThR.Tn[0].t36 VGND 0.01514f
C5158 XThR.Tn[0].n77 VGND 0.03697f
C5159 XThR.Tn[0].t62 VGND 0.01378f
C5160 XThR.Tn[0].t30 VGND 0.01509f
C5161 XThR.Tn[0].n78 VGND 0.03846f
C5162 XThR.Tn[0].n79 VGND 0.02702f
C5163 XThR.Tn[0].n81 VGND 0.08671f
C5164 XThR.Tn[0].t18 VGND 0.01383f
C5165 XThR.Tn[0].t32 VGND 0.01514f
C5166 XThR.Tn[0].n82 VGND 0.03697f
C5167 XThR.Tn[0].t39 VGND 0.01378f
C5168 XThR.Tn[0].t20 VGND 0.01509f
C5169 XThR.Tn[0].n83 VGND 0.03846f
C5170 XThR.Tn[0].n84 VGND 0.02702f
C5171 XThR.Tn[0].n86 VGND 0.08671f
C5172 XThR.Tn[0].n87 VGND 0.0788f
C5173 XThR.Tn[0].n88 VGND 0.22563f
C5174 XThR.Tn[7].t2 VGND 0.0118f
C5175 XThR.Tn[7].t1 VGND 0.0118f
C5176 XThR.Tn[7].n0 VGND 0.02606f
C5177 XThR.Tn[7].t3 VGND 0.0118f
C5178 XThR.Tn[7].t0 VGND 0.0118f
C5179 XThR.Tn[7].n1 VGND 0.03641f
C5180 XThR.Tn[7].n2 VGND 0.13363f
C5181 XThR.Tn[7].t6 VGND 0.01815f
C5182 XThR.Tn[7].t7 VGND 0.01815f
C5183 XThR.Tn[7].n3 VGND 0.05527f
C5184 XThR.Tn[7].t5 VGND 0.01815f
C5185 XThR.Tn[7].t4 VGND 0.01815f
C5186 XThR.Tn[7].n4 VGND 0.04021f
C5187 XThR.Tn[7].n5 VGND 0.17693f
C5188 XThR.Tn[7].n6 VGND 0.02205f
C5189 XThR.Tn[7].t53 VGND 0.01419f
C5190 XThR.Tn[7].t45 VGND 0.01553f
C5191 XThR.Tn[7].n7 VGND 0.03793f
C5192 XThR.Tn[7].n8 VGND 0.07287f
C5193 XThR.Tn[7].t8 VGND 0.01419f
C5194 XThR.Tn[7].t60 VGND 0.01553f
C5195 XThR.Tn[7].n9 VGND 0.03793f
C5196 XThR.Tn[7].t26 VGND 0.01414f
C5197 XThR.Tn[7].t38 VGND 0.01548f
C5198 XThR.Tn[7].n10 VGND 0.03947f
C5199 XThR.Tn[7].n11 VGND 0.02773f
C5200 XThR.Tn[7].n13 VGND 0.08897f
C5201 XThR.Tn[7].t47 VGND 0.01419f
C5202 XThR.Tn[7].t37 VGND 0.01553f
C5203 XThR.Tn[7].n14 VGND 0.03793f
C5204 XThR.Tn[7].t66 VGND 0.01414f
C5205 XThR.Tn[7].t15 VGND 0.01548f
C5206 XThR.Tn[7].n15 VGND 0.03947f
C5207 XThR.Tn[7].n16 VGND 0.02773f
C5208 XThR.Tn[7].n18 VGND 0.08897f
C5209 XThR.Tn[7].t62 VGND 0.01419f
C5210 XThR.Tn[7].t55 VGND 0.01553f
C5211 XThR.Tn[7].n19 VGND 0.03793f
C5212 XThR.Tn[7].t18 VGND 0.01414f
C5213 XThR.Tn[7].t32 VGND 0.01548f
C5214 XThR.Tn[7].n20 VGND 0.03947f
C5215 XThR.Tn[7].n21 VGND 0.02773f
C5216 XThR.Tn[7].n23 VGND 0.08897f
C5217 XThR.Tn[7].t25 VGND 0.01419f
C5218 XThR.Tn[7].t21 VGND 0.01553f
C5219 XThR.Tn[7].n24 VGND 0.03793f
C5220 XThR.Tn[7].t50 VGND 0.01414f
C5221 XThR.Tn[7].t63 VGND 0.01548f
C5222 XThR.Tn[7].n25 VGND 0.03947f
C5223 XThR.Tn[7].n26 VGND 0.02773f
C5224 XThR.Tn[7].n28 VGND 0.08897f
C5225 XThR.Tn[7].t65 VGND 0.01419f
C5226 XThR.Tn[7].t56 VGND 0.01553f
C5227 XThR.Tn[7].n29 VGND 0.03793f
C5228 XThR.Tn[7].t19 VGND 0.01414f
C5229 XThR.Tn[7].t34 VGND 0.01548f
C5230 XThR.Tn[7].n30 VGND 0.03947f
C5231 XThR.Tn[7].n31 VGND 0.02773f
C5232 XThR.Tn[7].n33 VGND 0.08897f
C5233 XThR.Tn[7].t40 VGND 0.01419f
C5234 XThR.Tn[7].t11 VGND 0.01553f
C5235 XThR.Tn[7].n34 VGND 0.03793f
C5236 XThR.Tn[7].t58 VGND 0.01414f
C5237 XThR.Tn[7].t54 VGND 0.01548f
C5238 XThR.Tn[7].n35 VGND 0.03947f
C5239 XThR.Tn[7].n36 VGND 0.02773f
C5240 XThR.Tn[7].n38 VGND 0.08897f
C5241 XThR.Tn[7].t9 VGND 0.01419f
C5242 XThR.Tn[7].t68 VGND 0.01553f
C5243 XThR.Tn[7].n39 VGND 0.03793f
C5244 XThR.Tn[7].t27 VGND 0.01414f
C5245 XThR.Tn[7].t46 VGND 0.01548f
C5246 XThR.Tn[7].n40 VGND 0.03947f
C5247 XThR.Tn[7].n41 VGND 0.02773f
C5248 XThR.Tn[7].n43 VGND 0.08897f
C5249 XThR.Tn[7].t14 VGND 0.01419f
C5250 XThR.Tn[7].t20 VGND 0.01553f
C5251 XThR.Tn[7].n44 VGND 0.03793f
C5252 XThR.Tn[7].t31 VGND 0.01414f
C5253 XThR.Tn[7].t61 VGND 0.01548f
C5254 XThR.Tn[7].n45 VGND 0.03947f
C5255 XThR.Tn[7].n46 VGND 0.02773f
C5256 XThR.Tn[7].n48 VGND 0.08897f
C5257 XThR.Tn[7].t29 VGND 0.01419f
C5258 XThR.Tn[7].t39 VGND 0.01553f
C5259 XThR.Tn[7].n49 VGND 0.03793f
C5260 XThR.Tn[7].t52 VGND 0.01414f
C5261 XThR.Tn[7].t16 VGND 0.01548f
C5262 XThR.Tn[7].n50 VGND 0.03947f
C5263 XThR.Tn[7].n51 VGND 0.02773f
C5264 XThR.Tn[7].n53 VGND 0.08897f
C5265 XThR.Tn[7].t23 VGND 0.01419f
C5266 XThR.Tn[7].t57 VGND 0.01553f
C5267 XThR.Tn[7].n54 VGND 0.03793f
C5268 XThR.Tn[7].t43 VGND 0.01414f
C5269 XThR.Tn[7].t36 VGND 0.01548f
C5270 XThR.Tn[7].n55 VGND 0.03947f
C5271 XThR.Tn[7].n56 VGND 0.02773f
C5272 XThR.Tn[7].n58 VGND 0.08897f
C5273 XThR.Tn[7].t42 VGND 0.01419f
C5274 XThR.Tn[7].t33 VGND 0.01553f
C5275 XThR.Tn[7].n59 VGND 0.03793f
C5276 XThR.Tn[7].t59 VGND 0.01414f
C5277 XThR.Tn[7].t10 VGND 0.01548f
C5278 XThR.Tn[7].n60 VGND 0.03947f
C5279 XThR.Tn[7].n61 VGND 0.02773f
C5280 XThR.Tn[7].n63 VGND 0.08897f
C5281 XThR.Tn[7].t12 VGND 0.01419f
C5282 XThR.Tn[7].t69 VGND 0.01553f
C5283 XThR.Tn[7].n64 VGND 0.03793f
C5284 XThR.Tn[7].t30 VGND 0.01414f
C5285 XThR.Tn[7].t48 VGND 0.01548f
C5286 XThR.Tn[7].n65 VGND 0.03947f
C5287 XThR.Tn[7].n66 VGND 0.02773f
C5288 XThR.Tn[7].n68 VGND 0.08897f
C5289 XThR.Tn[7].t28 VGND 0.01419f
C5290 XThR.Tn[7].t22 VGND 0.01553f
C5291 XThR.Tn[7].n69 VGND 0.03793f
C5292 XThR.Tn[7].t51 VGND 0.01414f
C5293 XThR.Tn[7].t64 VGND 0.01548f
C5294 XThR.Tn[7].n70 VGND 0.03947f
C5295 XThR.Tn[7].n71 VGND 0.02773f
C5296 XThR.Tn[7].n73 VGND 0.08897f
C5297 XThR.Tn[7].t49 VGND 0.01419f
C5298 XThR.Tn[7].t41 VGND 0.01553f
C5299 XThR.Tn[7].n74 VGND 0.03793f
C5300 XThR.Tn[7].t67 VGND 0.01414f
C5301 XThR.Tn[7].t17 VGND 0.01548f
C5302 XThR.Tn[7].n75 VGND 0.03947f
C5303 XThR.Tn[7].n76 VGND 0.02773f
C5304 XThR.Tn[7].n78 VGND 0.08897f
C5305 XThR.Tn[7].t24 VGND 0.01419f
C5306 XThR.Tn[7].t35 VGND 0.01553f
C5307 XThR.Tn[7].n79 VGND 0.03793f
C5308 XThR.Tn[7].t44 VGND 0.01414f
C5309 XThR.Tn[7].t13 VGND 0.01548f
C5310 XThR.Tn[7].n80 VGND 0.03947f
C5311 XThR.Tn[7].n81 VGND 0.02773f
C5312 XThR.Tn[7].n83 VGND 0.08897f
C5313 XThR.Tn[7].n84 VGND 0.08086f
C5314 XThR.Tn[7].n85 VGND 0.32824f
C5315 XThR.Tn[11].t2 VGND 0.01248f
C5316 XThR.Tn[11].t0 VGND 0.01248f
C5317 XThR.Tn[11].n0 VGND 0.02496f
C5318 XThR.Tn[11].t3 VGND 0.01248f
C5319 XThR.Tn[11].t1 VGND 0.01248f
C5320 XThR.Tn[11].n1 VGND 0.03112f
C5321 XThR.Tn[11].n2 VGND 0.06279f
C5322 XThR.Tn[11].t8 VGND 0.0192f
C5323 XThR.Tn[11].t10 VGND 0.0192f
C5324 XThR.Tn[11].n3 VGND 0.05829f
C5325 XThR.Tn[11].t9 VGND 0.0192f
C5326 XThR.Tn[11].t11 VGND 0.0192f
C5327 XThR.Tn[11].n4 VGND 0.04268f
C5328 XThR.Tn[11].n5 VGND 0.19406f
C5329 XThR.Tn[11].t4 VGND 0.0192f
C5330 XThR.Tn[11].t6 VGND 0.0192f
C5331 XThR.Tn[11].n6 VGND 0.04148f
C5332 XThR.Tn[11].t5 VGND 0.0192f
C5333 XThR.Tn[11].t7 VGND 0.0192f
C5334 XThR.Tn[11].n7 VGND 0.06313f
C5335 XThR.Tn[11].n8 VGND 0.1753f
C5336 XThR.Tn[11].n9 VGND 0.02347f
C5337 XThR.Tn[11].t56 VGND 0.015f
C5338 XThR.Tn[11].t48 VGND 0.01643f
C5339 XThR.Tn[11].n10 VGND 0.04012f
C5340 XThR.Tn[11].n11 VGND 0.07707f
C5341 XThR.Tn[11].t12 VGND 0.015f
C5342 XThR.Tn[11].t67 VGND 0.01643f
C5343 XThR.Tn[11].n12 VGND 0.04012f
C5344 XThR.Tn[11].t27 VGND 0.01496f
C5345 XThR.Tn[11].t58 VGND 0.01638f
C5346 XThR.Tn[11].n13 VGND 0.04174f
C5347 XThR.Tn[11].n14 VGND 0.02933f
C5348 XThR.Tn[11].n16 VGND 0.09411f
C5349 XThR.Tn[11].t49 VGND 0.015f
C5350 XThR.Tn[11].t41 VGND 0.01643f
C5351 XThR.Tn[11].n17 VGND 0.04012f
C5352 XThR.Tn[11].t65 VGND 0.01496f
C5353 XThR.Tn[11].t36 VGND 0.01638f
C5354 XThR.Tn[11].n18 VGND 0.04174f
C5355 XThR.Tn[11].n19 VGND 0.02933f
C5356 XThR.Tn[11].n21 VGND 0.09411f
C5357 XThR.Tn[11].t68 VGND 0.015f
C5358 XThR.Tn[11].t60 VGND 0.01643f
C5359 XThR.Tn[11].n22 VGND 0.04012f
C5360 XThR.Tn[11].t18 VGND 0.01496f
C5361 XThR.Tn[11].t54 VGND 0.01638f
C5362 XThR.Tn[11].n23 VGND 0.04174f
C5363 XThR.Tn[11].n24 VGND 0.02933f
C5364 XThR.Tn[11].n26 VGND 0.09411f
C5365 XThR.Tn[11].t33 VGND 0.015f
C5366 XThR.Tn[11].t23 VGND 0.01643f
C5367 XThR.Tn[11].n27 VGND 0.04012f
C5368 XThR.Tn[11].t50 VGND 0.01496f
C5369 XThR.Tn[11].t19 VGND 0.01638f
C5370 XThR.Tn[11].n28 VGND 0.04174f
C5371 XThR.Tn[11].n29 VGND 0.02933f
C5372 XThR.Tn[11].n31 VGND 0.09411f
C5373 XThR.Tn[11].t70 VGND 0.015f
C5374 XThR.Tn[11].t62 VGND 0.01643f
C5375 XThR.Tn[11].n32 VGND 0.04012f
C5376 XThR.Tn[11].t21 VGND 0.01496f
C5377 XThR.Tn[11].t55 VGND 0.01638f
C5378 XThR.Tn[11].n33 VGND 0.04174f
C5379 XThR.Tn[11].n34 VGND 0.02933f
C5380 XThR.Tn[11].n36 VGND 0.09411f
C5381 XThR.Tn[11].t44 VGND 0.015f
C5382 XThR.Tn[11].t14 VGND 0.01643f
C5383 XThR.Tn[11].n37 VGND 0.04012f
C5384 XThR.Tn[11].t59 VGND 0.01496f
C5385 XThR.Tn[11].t72 VGND 0.01638f
C5386 XThR.Tn[11].n38 VGND 0.04174f
C5387 XThR.Tn[11].n39 VGND 0.02933f
C5388 XThR.Tn[11].n41 VGND 0.09411f
C5389 XThR.Tn[11].t13 VGND 0.015f
C5390 XThR.Tn[11].t71 VGND 0.01643f
C5391 XThR.Tn[11].n42 VGND 0.04012f
C5392 XThR.Tn[11].t28 VGND 0.01496f
C5393 XThR.Tn[11].t64 VGND 0.01638f
C5394 XThR.Tn[11].n43 VGND 0.04174f
C5395 XThR.Tn[11].n44 VGND 0.02933f
C5396 XThR.Tn[11].n46 VGND 0.09411f
C5397 XThR.Tn[11].t16 VGND 0.015f
C5398 XThR.Tn[11].t22 VGND 0.01643f
C5399 XThR.Tn[11].n47 VGND 0.04012f
C5400 XThR.Tn[11].t32 VGND 0.01496f
C5401 XThR.Tn[11].t17 VGND 0.01638f
C5402 XThR.Tn[11].n48 VGND 0.04174f
C5403 XThR.Tn[11].n49 VGND 0.02933f
C5404 XThR.Tn[11].n51 VGND 0.09411f
C5405 XThR.Tn[11].t35 VGND 0.015f
C5406 XThR.Tn[11].t43 VGND 0.01643f
C5407 XThR.Tn[11].n52 VGND 0.04012f
C5408 XThR.Tn[11].t52 VGND 0.01496f
C5409 XThR.Tn[11].t37 VGND 0.01638f
C5410 XThR.Tn[11].n53 VGND 0.04174f
C5411 XThR.Tn[11].n54 VGND 0.02933f
C5412 XThR.Tn[11].n56 VGND 0.09411f
C5413 XThR.Tn[11].t25 VGND 0.015f
C5414 XThR.Tn[11].t63 VGND 0.01643f
C5415 XThR.Tn[11].n57 VGND 0.04012f
C5416 XThR.Tn[11].t42 VGND 0.01496f
C5417 XThR.Tn[11].t57 VGND 0.01638f
C5418 XThR.Tn[11].n58 VGND 0.04174f
C5419 XThR.Tn[11].n59 VGND 0.02933f
C5420 XThR.Tn[11].n61 VGND 0.09411f
C5421 XThR.Tn[11].t47 VGND 0.015f
C5422 XThR.Tn[11].t39 VGND 0.01643f
C5423 XThR.Tn[11].n62 VGND 0.04012f
C5424 XThR.Tn[11].t61 VGND 0.01496f
C5425 XThR.Tn[11].t29 VGND 0.01638f
C5426 XThR.Tn[11].n63 VGND 0.04174f
C5427 XThR.Tn[11].n64 VGND 0.02933f
C5428 XThR.Tn[11].n66 VGND 0.09411f
C5429 XThR.Tn[11].t15 VGND 0.015f
C5430 XThR.Tn[11].t73 VGND 0.01643f
C5431 XThR.Tn[11].n67 VGND 0.04012f
C5432 XThR.Tn[11].t30 VGND 0.01496f
C5433 XThR.Tn[11].t66 VGND 0.01638f
C5434 XThR.Tn[11].n68 VGND 0.04174f
C5435 XThR.Tn[11].n69 VGND 0.02933f
C5436 XThR.Tn[11].n71 VGND 0.09411f
C5437 XThR.Tn[11].t34 VGND 0.015f
C5438 XThR.Tn[11].t24 VGND 0.01643f
C5439 XThR.Tn[11].n72 VGND 0.04012f
C5440 XThR.Tn[11].t51 VGND 0.01496f
C5441 XThR.Tn[11].t20 VGND 0.01638f
C5442 XThR.Tn[11].n73 VGND 0.04174f
C5443 XThR.Tn[11].n74 VGND 0.02933f
C5444 XThR.Tn[11].n76 VGND 0.09411f
C5445 XThR.Tn[11].t53 VGND 0.015f
C5446 XThR.Tn[11].t46 VGND 0.01643f
C5447 XThR.Tn[11].n77 VGND 0.04012f
C5448 XThR.Tn[11].t69 VGND 0.01496f
C5449 XThR.Tn[11].t38 VGND 0.01638f
C5450 XThR.Tn[11].n78 VGND 0.04174f
C5451 XThR.Tn[11].n79 VGND 0.02933f
C5452 XThR.Tn[11].n81 VGND 0.09411f
C5453 XThR.Tn[11].t26 VGND 0.015f
C5454 XThR.Tn[11].t40 VGND 0.01643f
C5455 XThR.Tn[11].n82 VGND 0.04012f
C5456 XThR.Tn[11].t45 VGND 0.01496f
C5457 XThR.Tn[11].t31 VGND 0.01638f
C5458 XThR.Tn[11].n83 VGND 0.04174f
C5459 XThR.Tn[11].n84 VGND 0.02933f
C5460 XThR.Tn[11].n86 VGND 0.09411f
C5461 XThR.Tn[11].n87 VGND 0.08553f
C5462 XThR.Tn[11].n88 VGND 0.30653f
C5463 XThR.Tn[4].t5 VGND 0.01806f
C5464 XThR.Tn[4].t6 VGND 0.01806f
C5465 XThR.Tn[4].n0 VGND 0.03645f
C5466 XThR.Tn[4].t4 VGND 0.01806f
C5467 XThR.Tn[4].t7 VGND 0.01806f
C5468 XThR.Tn[4].n1 VGND 0.04265f
C5469 XThR.Tn[4].n2 VGND 0.12794f
C5470 XThR.Tn[4].t11 VGND 0.01174f
C5471 XThR.Tn[4].t8 VGND 0.01174f
C5472 XThR.Tn[4].n3 VGND 0.02673f
C5473 XThR.Tn[4].t10 VGND 0.01174f
C5474 XThR.Tn[4].t9 VGND 0.01174f
C5475 XThR.Tn[4].n4 VGND 0.02673f
C5476 XThR.Tn[4].t0 VGND 0.01174f
C5477 XThR.Tn[4].t1 VGND 0.01174f
C5478 XThR.Tn[4].n5 VGND 0.04454f
C5479 XThR.Tn[4].t3 VGND 0.01174f
C5480 XThR.Tn[4].t2 VGND 0.01174f
C5481 XThR.Tn[4].n6 VGND 0.02673f
C5482 XThR.Tn[4].n7 VGND 0.1273f
C5483 XThR.Tn[4].n8 VGND 0.0787f
C5484 XThR.Tn[4].n9 VGND 0.08881f
C5485 XThR.Tn[4].t44 VGND 0.01411f
C5486 XThR.Tn[4].t38 VGND 0.01545f
C5487 XThR.Tn[4].n10 VGND 0.03774f
C5488 XThR.Tn[4].n11 VGND 0.0725f
C5489 XThR.Tn[4].t65 VGND 0.01411f
C5490 XThR.Tn[4].t54 VGND 0.01545f
C5491 XThR.Tn[4].n12 VGND 0.03774f
C5492 XThR.Tn[4].t19 VGND 0.01407f
C5493 XThR.Tn[4].t50 VGND 0.01541f
C5494 XThR.Tn[4].n13 VGND 0.03927f
C5495 XThR.Tn[4].n14 VGND 0.02759f
C5496 XThR.Tn[4].n16 VGND 0.08853f
C5497 XThR.Tn[4].t39 VGND 0.01411f
C5498 XThR.Tn[4].t31 VGND 0.01545f
C5499 XThR.Tn[4].n17 VGND 0.03774f
C5500 XThR.Tn[4].t58 VGND 0.01407f
C5501 XThR.Tn[4].t27 VGND 0.01541f
C5502 XThR.Tn[4].n18 VGND 0.03927f
C5503 XThR.Tn[4].n19 VGND 0.02759f
C5504 XThR.Tn[4].n21 VGND 0.08853f
C5505 XThR.Tn[4].t55 VGND 0.01411f
C5506 XThR.Tn[4].t48 VGND 0.01545f
C5507 XThR.Tn[4].n22 VGND 0.03774f
C5508 XThR.Tn[4].t70 VGND 0.01407f
C5509 XThR.Tn[4].t45 VGND 0.01541f
C5510 XThR.Tn[4].n23 VGND 0.03927f
C5511 XThR.Tn[4].n24 VGND 0.02759f
C5512 XThR.Tn[4].n26 VGND 0.08853f
C5513 XThR.Tn[4].t17 VGND 0.01411f
C5514 XThR.Tn[4].t13 VGND 0.01545f
C5515 XThR.Tn[4].n27 VGND 0.03774f
C5516 XThR.Tn[4].t41 VGND 0.01407f
C5517 XThR.Tn[4].t71 VGND 0.01541f
C5518 XThR.Tn[4].n28 VGND 0.03927f
C5519 XThR.Tn[4].n29 VGND 0.02759f
C5520 XThR.Tn[4].n31 VGND 0.08853f
C5521 XThR.Tn[4].t57 VGND 0.01411f
C5522 XThR.Tn[4].t49 VGND 0.01545f
C5523 XThR.Tn[4].n32 VGND 0.03774f
C5524 XThR.Tn[4].t73 VGND 0.01407f
C5525 XThR.Tn[4].t46 VGND 0.01541f
C5526 XThR.Tn[4].n33 VGND 0.03927f
C5527 XThR.Tn[4].n34 VGND 0.02759f
C5528 XThR.Tn[4].n36 VGND 0.08853f
C5529 XThR.Tn[4].t33 VGND 0.01411f
C5530 XThR.Tn[4].t66 VGND 0.01545f
C5531 XThR.Tn[4].n37 VGND 0.03774f
C5532 XThR.Tn[4].t52 VGND 0.01407f
C5533 XThR.Tn[4].t63 VGND 0.01541f
C5534 XThR.Tn[4].n38 VGND 0.03927f
C5535 XThR.Tn[4].n39 VGND 0.02759f
C5536 XThR.Tn[4].n41 VGND 0.08853f
C5537 XThR.Tn[4].t64 VGND 0.01411f
C5538 XThR.Tn[4].t61 VGND 0.01545f
C5539 XThR.Tn[4].n42 VGND 0.03774f
C5540 XThR.Tn[4].t18 VGND 0.01407f
C5541 XThR.Tn[4].t56 VGND 0.01541f
C5542 XThR.Tn[4].n43 VGND 0.03927f
C5543 XThR.Tn[4].n44 VGND 0.02759f
C5544 XThR.Tn[4].n46 VGND 0.08853f
C5545 XThR.Tn[4].t68 VGND 0.01411f
C5546 XThR.Tn[4].t12 VGND 0.01545f
C5547 XThR.Tn[4].n47 VGND 0.03774f
C5548 XThR.Tn[4].t25 VGND 0.01407f
C5549 XThR.Tn[4].t69 VGND 0.01541f
C5550 XThR.Tn[4].n48 VGND 0.03927f
C5551 XThR.Tn[4].n49 VGND 0.02759f
C5552 XThR.Tn[4].n51 VGND 0.08853f
C5553 XThR.Tn[4].t22 VGND 0.01411f
C5554 XThR.Tn[4].t32 VGND 0.01545f
C5555 XThR.Tn[4].n52 VGND 0.03774f
C5556 XThR.Tn[4].t43 VGND 0.01407f
C5557 XThR.Tn[4].t29 VGND 0.01541f
C5558 XThR.Tn[4].n53 VGND 0.03927f
C5559 XThR.Tn[4].n54 VGND 0.02759f
C5560 XThR.Tn[4].n56 VGND 0.08853f
C5561 XThR.Tn[4].t15 VGND 0.01411f
C5562 XThR.Tn[4].t51 VGND 0.01545f
C5563 XThR.Tn[4].n57 VGND 0.03774f
C5564 XThR.Tn[4].t36 VGND 0.01407f
C5565 XThR.Tn[4].t47 VGND 0.01541f
C5566 XThR.Tn[4].n58 VGND 0.03927f
C5567 XThR.Tn[4].n59 VGND 0.02759f
C5568 XThR.Tn[4].n61 VGND 0.08853f
C5569 XThR.Tn[4].t35 VGND 0.01411f
C5570 XThR.Tn[4].t26 VGND 0.01545f
C5571 XThR.Tn[4].n62 VGND 0.03774f
C5572 XThR.Tn[4].t53 VGND 0.01407f
C5573 XThR.Tn[4].t21 VGND 0.01541f
C5574 XThR.Tn[4].n63 VGND 0.03927f
C5575 XThR.Tn[4].n64 VGND 0.02759f
C5576 XThR.Tn[4].n66 VGND 0.08853f
C5577 XThR.Tn[4].t67 VGND 0.01411f
C5578 XThR.Tn[4].t62 VGND 0.01545f
C5579 XThR.Tn[4].n67 VGND 0.03774f
C5580 XThR.Tn[4].t23 VGND 0.01407f
C5581 XThR.Tn[4].t59 VGND 0.01541f
C5582 XThR.Tn[4].n68 VGND 0.03927f
C5583 XThR.Tn[4].n69 VGND 0.02759f
C5584 XThR.Tn[4].n71 VGND 0.08853f
C5585 XThR.Tn[4].t20 VGND 0.01411f
C5586 XThR.Tn[4].t14 VGND 0.01545f
C5587 XThR.Tn[4].n72 VGND 0.03774f
C5588 XThR.Tn[4].t42 VGND 0.01407f
C5589 XThR.Tn[4].t72 VGND 0.01541f
C5590 XThR.Tn[4].n73 VGND 0.03927f
C5591 XThR.Tn[4].n74 VGND 0.02759f
C5592 XThR.Tn[4].n76 VGND 0.08853f
C5593 XThR.Tn[4].t40 VGND 0.01411f
C5594 XThR.Tn[4].t34 VGND 0.01545f
C5595 XThR.Tn[4].n77 VGND 0.03774f
C5596 XThR.Tn[4].t60 VGND 0.01407f
C5597 XThR.Tn[4].t30 VGND 0.01541f
C5598 XThR.Tn[4].n78 VGND 0.03927f
C5599 XThR.Tn[4].n79 VGND 0.02759f
C5600 XThR.Tn[4].n81 VGND 0.08853f
C5601 XThR.Tn[4].t16 VGND 0.01411f
C5602 XThR.Tn[4].t28 VGND 0.01545f
C5603 XThR.Tn[4].n82 VGND 0.03774f
C5604 XThR.Tn[4].t37 VGND 0.01407f
C5605 XThR.Tn[4].t24 VGND 0.01541f
C5606 XThR.Tn[4].n83 VGND 0.03927f
C5607 XThR.Tn[4].n84 VGND 0.02759f
C5608 XThR.Tn[4].n86 VGND 0.08853f
C5609 XThR.Tn[4].n87 VGND 0.08045f
C5610 XThR.Tn[4].n88 VGND 0.15199f
C5611 XThC.Tn[7].t4 VGND 0.01305f
C5612 XThC.Tn[7].t7 VGND 0.01305f
C5613 XThC.Tn[7].n0 VGND 0.0281f
C5614 XThC.Tn[7].t6 VGND 0.01305f
C5615 XThC.Tn[7].t5 VGND 0.01305f
C5616 XThC.Tn[7].n1 VGND 0.04266f
C5617 XThC.Tn[7].n2 VGND 0.12542f
C5618 XThC.Tn[7].t8 VGND 0.01034f
C5619 XThC.Tn[7].t11 VGND 0.01129f
C5620 XThC.Tn[7].n3 VGND 0.02522f
C5621 XThC.Tn[7].n4 VGND 0.01441f
C5622 XThC.Tn[7].n5 VGND 0.01753f
C5623 XThC.Tn[7].t25 VGND 0.01034f
C5624 XThC.Tn[7].t30 VGND 0.01129f
C5625 XThC.Tn[7].n6 VGND 0.02522f
C5626 XThC.Tn[7].n7 VGND 0.01441f
C5627 XThC.Tn[7].n8 VGND 0.08328f
C5628 XThC.Tn[7].t27 VGND 0.01034f
C5629 XThC.Tn[7].t34 VGND 0.01129f
C5630 XThC.Tn[7].n9 VGND 0.02522f
C5631 XThC.Tn[7].n10 VGND 0.01441f
C5632 XThC.Tn[7].n11 VGND 0.08328f
C5633 XThC.Tn[7].t29 VGND 0.01034f
C5634 XThC.Tn[7].t35 VGND 0.01129f
C5635 XThC.Tn[7].n12 VGND 0.02522f
C5636 XThC.Tn[7].n13 VGND 0.01441f
C5637 XThC.Tn[7].n14 VGND 0.08328f
C5638 XThC.Tn[7].t18 VGND 0.01034f
C5639 XThC.Tn[7].t22 VGND 0.01129f
C5640 XThC.Tn[7].n15 VGND 0.02522f
C5641 XThC.Tn[7].n16 VGND 0.01441f
C5642 XThC.Tn[7].n17 VGND 0.08328f
C5643 XThC.Tn[7].t20 VGND 0.01034f
C5644 XThC.Tn[7].t23 VGND 0.01129f
C5645 XThC.Tn[7].n18 VGND 0.02522f
C5646 XThC.Tn[7].n19 VGND 0.01441f
C5647 XThC.Tn[7].n20 VGND 0.08328f
C5648 XThC.Tn[7].t33 VGND 0.01034f
C5649 XThC.Tn[7].t39 VGND 0.01129f
C5650 XThC.Tn[7].n21 VGND 0.02522f
C5651 XThC.Tn[7].n22 VGND 0.01441f
C5652 XThC.Tn[7].n23 VGND 0.08328f
C5653 XThC.Tn[7].t10 VGND 0.01034f
C5654 XThC.Tn[7].t14 VGND 0.01129f
C5655 XThC.Tn[7].n24 VGND 0.02522f
C5656 XThC.Tn[7].n25 VGND 0.01441f
C5657 XThC.Tn[7].n26 VGND 0.08328f
C5658 XThC.Tn[7].t12 VGND 0.01034f
C5659 XThC.Tn[7].t16 VGND 0.01129f
C5660 XThC.Tn[7].n27 VGND 0.02522f
C5661 XThC.Tn[7].n28 VGND 0.01441f
C5662 XThC.Tn[7].n29 VGND 0.08328f
C5663 XThC.Tn[7].t31 VGND 0.01034f
C5664 XThC.Tn[7].t36 VGND 0.01129f
C5665 XThC.Tn[7].n30 VGND 0.02522f
C5666 XThC.Tn[7].n31 VGND 0.01441f
C5667 XThC.Tn[7].n32 VGND 0.08328f
C5668 XThC.Tn[7].t32 VGND 0.01034f
C5669 XThC.Tn[7].t38 VGND 0.01129f
C5670 XThC.Tn[7].n33 VGND 0.02522f
C5671 XThC.Tn[7].n34 VGND 0.01441f
C5672 XThC.Tn[7].n35 VGND 0.08328f
C5673 XThC.Tn[7].t13 VGND 0.01034f
C5674 XThC.Tn[7].t17 VGND 0.01129f
C5675 XThC.Tn[7].n36 VGND 0.02522f
C5676 XThC.Tn[7].n37 VGND 0.01441f
C5677 XThC.Tn[7].n38 VGND 0.08328f
C5678 XThC.Tn[7].t21 VGND 0.01034f
C5679 XThC.Tn[7].t26 VGND 0.01129f
C5680 XThC.Tn[7].n39 VGND 0.02522f
C5681 XThC.Tn[7].n40 VGND 0.01441f
C5682 XThC.Tn[7].n41 VGND 0.08328f
C5683 XThC.Tn[7].t24 VGND 0.01034f
C5684 XThC.Tn[7].t28 VGND 0.01129f
C5685 XThC.Tn[7].n42 VGND 0.02522f
C5686 XThC.Tn[7].n43 VGND 0.01441f
C5687 XThC.Tn[7].n44 VGND 0.08328f
C5688 XThC.Tn[7].t37 VGND 0.01034f
C5689 XThC.Tn[7].t9 VGND 0.01129f
C5690 XThC.Tn[7].n45 VGND 0.02522f
C5691 XThC.Tn[7].n46 VGND 0.01441f
C5692 XThC.Tn[7].n47 VGND 0.08328f
C5693 XThC.Tn[7].t15 VGND 0.01034f
C5694 XThC.Tn[7].t19 VGND 0.01129f
C5695 XThC.Tn[7].n48 VGND 0.02522f
C5696 XThC.Tn[7].n49 VGND 0.01441f
C5697 XThC.Tn[7].n50 VGND 0.08328f
C5698 XThC.Tn[7].n51 VGND 0.52699f
C5699 XThC.Tn[7].n52 VGND 0.03388f
C5700 XThC.Tn[7].n53 VGND 0.02617f
C5701 XThC.Tn[7].n54 VGND 0.01873f
C5702 XThC.Tn[7].n55 VGND 0.09263f
C5703 XThC.Tn[7].n56 VGND 0.01561f
C5704 XThR.Tn[1].t4 VGND 0.01794f
C5705 XThR.Tn[1].t5 VGND 0.01794f
C5706 XThR.Tn[1].n0 VGND 0.03622f
C5707 XThR.Tn[1].t7 VGND 0.01794f
C5708 XThR.Tn[1].t6 VGND 0.01794f
C5709 XThR.Tn[1].n1 VGND 0.04238f
C5710 XThR.Tn[1].n2 VGND 0.11863f
C5711 XThR.Tn[1].t11 VGND 0.01166f
C5712 XThR.Tn[1].t8 VGND 0.01166f
C5713 XThR.Tn[1].n3 VGND 0.02656f
C5714 XThR.Tn[1].t10 VGND 0.01166f
C5715 XThR.Tn[1].t9 VGND 0.01166f
C5716 XThR.Tn[1].n4 VGND 0.02656f
C5717 XThR.Tn[1].t2 VGND 0.01166f
C5718 XThR.Tn[1].t1 VGND 0.01166f
C5719 XThR.Tn[1].n5 VGND 0.02656f
C5720 XThR.Tn[1].t3 VGND 0.01166f
C5721 XThR.Tn[1].t0 VGND 0.01166f
C5722 XThR.Tn[1].n6 VGND 0.04425f
C5723 XThR.Tn[1].n7 VGND 0.12648f
C5724 XThR.Tn[1].n8 VGND 0.07819f
C5725 XThR.Tn[1].n9 VGND 0.08824f
C5726 XThR.Tn[1].t24 VGND 0.01402f
C5727 XThR.Tn[1].t18 VGND 0.01536f
C5728 XThR.Tn[1].n10 VGND 0.0375f
C5729 XThR.Tn[1].n11 VGND 0.07203f
C5730 XThR.Tn[1].t44 VGND 0.01402f
C5731 XThR.Tn[1].t34 VGND 0.01536f
C5732 XThR.Tn[1].n12 VGND 0.0375f
C5733 XThR.Tn[1].t61 VGND 0.01398f
C5734 XThR.Tn[1].t30 VGND 0.01531f
C5735 XThR.Tn[1].n13 VGND 0.03901f
C5736 XThR.Tn[1].n14 VGND 0.02741f
C5737 XThR.Tn[1].n16 VGND 0.08795f
C5738 XThR.Tn[1].t19 VGND 0.01402f
C5739 XThR.Tn[1].t73 VGND 0.01536f
C5740 XThR.Tn[1].n17 VGND 0.0375f
C5741 XThR.Tn[1].t38 VGND 0.01398f
C5742 XThR.Tn[1].t69 VGND 0.01531f
C5743 XThR.Tn[1].n18 VGND 0.03901f
C5744 XThR.Tn[1].n19 VGND 0.02741f
C5745 XThR.Tn[1].n21 VGND 0.08795f
C5746 XThR.Tn[1].t35 VGND 0.01402f
C5747 XThR.Tn[1].t28 VGND 0.01536f
C5748 XThR.Tn[1].n22 VGND 0.0375f
C5749 XThR.Tn[1].t50 VGND 0.01398f
C5750 XThR.Tn[1].t25 VGND 0.01531f
C5751 XThR.Tn[1].n23 VGND 0.03901f
C5752 XThR.Tn[1].n24 VGND 0.02741f
C5753 XThR.Tn[1].n26 VGND 0.08795f
C5754 XThR.Tn[1].t59 VGND 0.01402f
C5755 XThR.Tn[1].t55 VGND 0.01536f
C5756 XThR.Tn[1].n27 VGND 0.0375f
C5757 XThR.Tn[1].t21 VGND 0.01398f
C5758 XThR.Tn[1].t51 VGND 0.01531f
C5759 XThR.Tn[1].n28 VGND 0.03901f
C5760 XThR.Tn[1].n29 VGND 0.02741f
C5761 XThR.Tn[1].n31 VGND 0.08795f
C5762 XThR.Tn[1].t37 VGND 0.01402f
C5763 XThR.Tn[1].t29 VGND 0.01536f
C5764 XThR.Tn[1].n32 VGND 0.0375f
C5765 XThR.Tn[1].t53 VGND 0.01398f
C5766 XThR.Tn[1].t26 VGND 0.01531f
C5767 XThR.Tn[1].n33 VGND 0.03901f
C5768 XThR.Tn[1].n34 VGND 0.02741f
C5769 XThR.Tn[1].n36 VGND 0.08795f
C5770 XThR.Tn[1].t13 VGND 0.01402f
C5771 XThR.Tn[1].t46 VGND 0.01536f
C5772 XThR.Tn[1].n37 VGND 0.0375f
C5773 XThR.Tn[1].t32 VGND 0.01398f
C5774 XThR.Tn[1].t43 VGND 0.01531f
C5775 XThR.Tn[1].n38 VGND 0.03901f
C5776 XThR.Tn[1].n39 VGND 0.02741f
C5777 XThR.Tn[1].n41 VGND 0.08795f
C5778 XThR.Tn[1].t45 VGND 0.01402f
C5779 XThR.Tn[1].t41 VGND 0.01536f
C5780 XThR.Tn[1].n42 VGND 0.0375f
C5781 XThR.Tn[1].t60 VGND 0.01398f
C5782 XThR.Tn[1].t36 VGND 0.01531f
C5783 XThR.Tn[1].n43 VGND 0.03901f
C5784 XThR.Tn[1].n44 VGND 0.02741f
C5785 XThR.Tn[1].n46 VGND 0.08795f
C5786 XThR.Tn[1].t48 VGND 0.01402f
C5787 XThR.Tn[1].t54 VGND 0.01536f
C5788 XThR.Tn[1].n47 VGND 0.0375f
C5789 XThR.Tn[1].t67 VGND 0.01398f
C5790 XThR.Tn[1].t49 VGND 0.01531f
C5791 XThR.Tn[1].n48 VGND 0.03901f
C5792 XThR.Tn[1].n49 VGND 0.02741f
C5793 XThR.Tn[1].n51 VGND 0.08795f
C5794 XThR.Tn[1].t64 VGND 0.01402f
C5795 XThR.Tn[1].t12 VGND 0.01536f
C5796 XThR.Tn[1].n52 VGND 0.0375f
C5797 XThR.Tn[1].t23 VGND 0.01398f
C5798 XThR.Tn[1].t71 VGND 0.01531f
C5799 XThR.Tn[1].n53 VGND 0.03901f
C5800 XThR.Tn[1].n54 VGND 0.02741f
C5801 XThR.Tn[1].n56 VGND 0.08795f
C5802 XThR.Tn[1].t57 VGND 0.01402f
C5803 XThR.Tn[1].t31 VGND 0.01536f
C5804 XThR.Tn[1].n57 VGND 0.0375f
C5805 XThR.Tn[1].t16 VGND 0.01398f
C5806 XThR.Tn[1].t27 VGND 0.01531f
C5807 XThR.Tn[1].n58 VGND 0.03901f
C5808 XThR.Tn[1].n59 VGND 0.02741f
C5809 XThR.Tn[1].n61 VGND 0.08795f
C5810 XThR.Tn[1].t15 VGND 0.01402f
C5811 XThR.Tn[1].t68 VGND 0.01536f
C5812 XThR.Tn[1].n62 VGND 0.0375f
C5813 XThR.Tn[1].t33 VGND 0.01398f
C5814 XThR.Tn[1].t63 VGND 0.01531f
C5815 XThR.Tn[1].n63 VGND 0.03901f
C5816 XThR.Tn[1].n64 VGND 0.02741f
C5817 XThR.Tn[1].n66 VGND 0.08795f
C5818 XThR.Tn[1].t47 VGND 0.01402f
C5819 XThR.Tn[1].t42 VGND 0.01536f
C5820 XThR.Tn[1].n67 VGND 0.0375f
C5821 XThR.Tn[1].t65 VGND 0.01398f
C5822 XThR.Tn[1].t39 VGND 0.01531f
C5823 XThR.Tn[1].n68 VGND 0.03901f
C5824 XThR.Tn[1].n69 VGND 0.02741f
C5825 XThR.Tn[1].n71 VGND 0.08795f
C5826 XThR.Tn[1].t62 VGND 0.01402f
C5827 XThR.Tn[1].t56 VGND 0.01536f
C5828 XThR.Tn[1].n72 VGND 0.0375f
C5829 XThR.Tn[1].t22 VGND 0.01398f
C5830 XThR.Tn[1].t52 VGND 0.01531f
C5831 XThR.Tn[1].n73 VGND 0.03901f
C5832 XThR.Tn[1].n74 VGND 0.02741f
C5833 XThR.Tn[1].n76 VGND 0.08795f
C5834 XThR.Tn[1].t20 VGND 0.01402f
C5835 XThR.Tn[1].t14 VGND 0.01536f
C5836 XThR.Tn[1].n77 VGND 0.0375f
C5837 XThR.Tn[1].t40 VGND 0.01398f
C5838 XThR.Tn[1].t72 VGND 0.01531f
C5839 XThR.Tn[1].n78 VGND 0.03901f
C5840 XThR.Tn[1].n79 VGND 0.02741f
C5841 XThR.Tn[1].n81 VGND 0.08795f
C5842 XThR.Tn[1].t58 VGND 0.01402f
C5843 XThR.Tn[1].t70 VGND 0.01536f
C5844 XThR.Tn[1].n82 VGND 0.0375f
C5845 XThR.Tn[1].t17 VGND 0.01398f
C5846 XThR.Tn[1].t66 VGND 0.01531f
C5847 XThR.Tn[1].n83 VGND 0.03901f
C5848 XThR.Tn[1].n84 VGND 0.02741f
C5849 XThR.Tn[1].n86 VGND 0.08795f
C5850 XThR.Tn[1].n87 VGND 0.07993f
C5851 XThR.Tn[1].n88 VGND 0.23008f
C5852 XThR.Tn[1].n89 VGND 0.03755f
C5853 XThC.Tn[8].n0 VGND 0.02379f
C5854 XThC.Tn[8].n1 VGND 0.01907f
C5855 XThC.Tn[8].n2 VGND 0.04799f
C5856 XThC.Tn[8].t5 VGND 0.01467f
C5857 XThC.Tn[8].t6 VGND 0.01467f
C5858 XThC.Tn[8].n3 VGND 0.0317f
C5859 XThC.Tn[8].t4 VGND 0.01467f
C5860 XThC.Tn[8].t7 VGND 0.01467f
C5861 XThC.Tn[8].n4 VGND 0.04825f
C5862 XThC.Tn[8].n5 VGND 0.13407f
C5863 XThC.Tn[8].t8 VGND 0.01467f
C5864 XThC.Tn[8].t11 VGND 0.01467f
C5865 XThC.Tn[8].n6 VGND 0.04455f
C5866 XThC.Tn[8].t10 VGND 0.01467f
C5867 XThC.Tn[8].t9 VGND 0.01467f
C5868 XThC.Tn[8].n7 VGND 0.03262f
C5869 XThC.Tn[8].n8 VGND 0.14517f
C5870 XThC.Tn[8].n9 VGND 0.02108f
C5871 XThC.Tn[8].t43 VGND 0.01163f
C5872 XThC.Tn[8].t41 VGND 0.0127f
C5873 XThC.Tn[8].n10 VGND 0.02837f
C5874 XThC.Tn[8].n11 VGND 0.01621f
C5875 XThC.Tn[8].n12 VGND 0.01972f
C5876 XThC.Tn[8].t29 VGND 0.01163f
C5877 XThC.Tn[8].t26 VGND 0.0127f
C5878 XThC.Tn[8].n13 VGND 0.02837f
C5879 XThC.Tn[8].n14 VGND 0.01621f
C5880 XThC.Tn[8].n15 VGND 0.09367f
C5881 XThC.Tn[8].t34 VGND 0.01163f
C5882 XThC.Tn[8].t28 VGND 0.0127f
C5883 XThC.Tn[8].n16 VGND 0.02837f
C5884 XThC.Tn[8].n17 VGND 0.01621f
C5885 XThC.Tn[8].n18 VGND 0.09367f
C5886 XThC.Tn[8].t35 VGND 0.01163f
C5887 XThC.Tn[8].t30 VGND 0.0127f
C5888 XThC.Tn[8].n19 VGND 0.02837f
C5889 XThC.Tn[8].n20 VGND 0.01621f
C5890 XThC.Tn[8].n21 VGND 0.09367f
C5891 XThC.Tn[8].t22 VGND 0.01163f
C5892 XThC.Tn[8].t19 VGND 0.0127f
C5893 XThC.Tn[8].n22 VGND 0.02837f
C5894 XThC.Tn[8].n23 VGND 0.01621f
C5895 XThC.Tn[8].n24 VGND 0.09367f
C5896 XThC.Tn[8].t23 VGND 0.01163f
C5897 XThC.Tn[8].t20 VGND 0.0127f
C5898 XThC.Tn[8].n25 VGND 0.02837f
C5899 XThC.Tn[8].n26 VGND 0.01621f
C5900 XThC.Tn[8].n27 VGND 0.09367f
C5901 XThC.Tn[8].t39 VGND 0.01163f
C5902 XThC.Tn[8].t33 VGND 0.0127f
C5903 XThC.Tn[8].n28 VGND 0.02837f
C5904 XThC.Tn[8].n29 VGND 0.01621f
C5905 XThC.Tn[8].n30 VGND 0.09367f
C5906 XThC.Tn[8].t14 VGND 0.01163f
C5907 XThC.Tn[8].t42 VGND 0.0127f
C5908 XThC.Tn[8].n31 VGND 0.02837f
C5909 XThC.Tn[8].n32 VGND 0.01621f
C5910 XThC.Tn[8].n33 VGND 0.09367f
C5911 XThC.Tn[8].t16 VGND 0.01163f
C5912 XThC.Tn[8].t12 VGND 0.0127f
C5913 XThC.Tn[8].n34 VGND 0.02837f
C5914 XThC.Tn[8].n35 VGND 0.01621f
C5915 XThC.Tn[8].n36 VGND 0.09367f
C5916 XThC.Tn[8].t36 VGND 0.01163f
C5917 XThC.Tn[8].t31 VGND 0.0127f
C5918 XThC.Tn[8].n37 VGND 0.02837f
C5919 XThC.Tn[8].n38 VGND 0.01621f
C5920 XThC.Tn[8].n39 VGND 0.09367f
C5921 XThC.Tn[8].t38 VGND 0.01163f
C5922 XThC.Tn[8].t32 VGND 0.0127f
C5923 XThC.Tn[8].n40 VGND 0.02837f
C5924 XThC.Tn[8].n41 VGND 0.01621f
C5925 XThC.Tn[8].n42 VGND 0.09367f
C5926 XThC.Tn[8].t17 VGND 0.01163f
C5927 XThC.Tn[8].t13 VGND 0.0127f
C5928 XThC.Tn[8].n43 VGND 0.02837f
C5929 XThC.Tn[8].n44 VGND 0.01621f
C5930 XThC.Tn[8].n45 VGND 0.09367f
C5931 XThC.Tn[8].t25 VGND 0.01163f
C5932 XThC.Tn[8].t21 VGND 0.0127f
C5933 XThC.Tn[8].n46 VGND 0.02837f
C5934 XThC.Tn[8].n47 VGND 0.01621f
C5935 XThC.Tn[8].n48 VGND 0.09367f
C5936 XThC.Tn[8].t27 VGND 0.01163f
C5937 XThC.Tn[8].t24 VGND 0.0127f
C5938 XThC.Tn[8].n49 VGND 0.02837f
C5939 XThC.Tn[8].n50 VGND 0.01621f
C5940 XThC.Tn[8].n51 VGND 0.09367f
C5941 XThC.Tn[8].t40 VGND 0.01163f
C5942 XThC.Tn[8].t37 VGND 0.0127f
C5943 XThC.Tn[8].n52 VGND 0.02837f
C5944 XThC.Tn[8].n53 VGND 0.01621f
C5945 XThC.Tn[8].n54 VGND 0.09367f
C5946 XThC.Tn[8].t18 VGND 0.01163f
C5947 XThC.Tn[8].t15 VGND 0.0127f
C5948 XThC.Tn[8].n55 VGND 0.02837f
C5949 XThC.Tn[8].n56 VGND 0.01621f
C5950 XThC.Tn[8].n57 VGND 0.09367f
C5951 XThC.Tn[8].n58 VGND 0.04332f
C5952 XThC.Tn[8].n59 VGND 0.41007f
C5953 XThC.Tn[8].n60 VGND 0.03291f
C5954 XThC.XTB1.Y.t1 VGND 0.03224f
C5955 XThC.XTB1.Y.n0 VGND 0.02084f
C5956 XThC.XTB1.Y.n1 VGND 0.02659f
C5957 XThC.XTB1.Y.t0 VGND 0.01618f
C5958 XThC.XTB1.Y.t2 VGND 0.01618f
C5959 XThC.XTB1.Y.n2 VGND 0.03473f
C5960 XThC.XTB1.Y.t17 VGND 0.02517f
C5961 XThC.XTB1.Y.t5 VGND 0.01483f
C5962 XThC.XTB1.Y.n3 VGND 0.02997f
C5963 XThC.XTB1.Y.t6 VGND 0.02517f
C5964 XThC.XTB1.Y.t12 VGND 0.01483f
C5965 XThC.XTB1.Y.n4 VGND 0.01542f
C5966 XThC.XTB1.Y.t8 VGND 0.02517f
C5967 XThC.XTB1.Y.t13 VGND 0.01483f
C5968 XThC.XTB1.Y.n5 VGND 0.03313f
C5969 XThC.XTB1.Y.t11 VGND 0.02517f
C5970 XThC.XTB1.Y.t16 VGND 0.01483f
C5971 XThC.XTB1.Y.n6 VGND 0.03076f
C5972 XThC.XTB1.Y.n7 VGND 0.01871f
C5973 XThC.XTB1.Y.n8 VGND 0.03098f
C5974 XThC.XTB1.Y.n9 VGND 0.01198f
C5975 XThC.XTB1.Y.n10 VGND 0.01463f
C5976 XThC.XTB1.Y.n11 VGND 0.03313f
C5977 XThC.XTB1.Y.n12 VGND 0.01661f
C5978 XThC.XTB1.Y.n13 VGND 0.02824f
C5979 XThC.XTB1.Y.t18 VGND 0.02517f
C5980 XThC.XTB1.Y.t9 VGND 0.01483f
C5981 XThC.XTB1.Y.n14 VGND 0.03392f
C5982 XThC.XTB1.Y.t7 VGND 0.02517f
C5983 XThC.XTB1.Y.t15 VGND 0.01483f
C5984 XThC.XTB1.Y.t14 VGND 0.02517f
C5985 XThC.XTB1.Y.t3 VGND 0.01483f
C5986 XThC.XTB1.Y.t10 VGND 0.02517f
C5987 XThC.XTB1.Y.t4 VGND 0.01483f
C5988 XThC.XTB1.Y.n15 VGND 0.04223f
C5989 XThC.XTB1.Y.n16 VGND 0.0446f
C5990 XThC.XTB1.Y.n17 VGND 0.01719f
C5991 XThC.XTB1.Y.n18 VGND 0.0363f
C5992 XThC.XTB1.Y.n19 VGND 0.01661f
C5993 XThC.XTB1.Y.n20 VGND 0.01378f
C5994 XThC.XTB1.Y.n21 VGND 0.77148f
C5995 XThC.XTB1.Y.n22 VGND 0.07634f
C5996 XThC.Tn[14].n0 VGND 0.02301f
C5997 XThC.Tn[14].n1 VGND 0.01845f
C5998 XThC.Tn[14].n2 VGND 0.04642f
C5999 XThC.Tn[14].t4 VGND 0.01419f
C6000 XThC.Tn[14].t5 VGND 0.01419f
C6001 XThC.Tn[14].n3 VGND 0.03067f
C6002 XThC.Tn[14].t7 VGND 0.01419f
C6003 XThC.Tn[14].t6 VGND 0.01419f
C6004 XThC.Tn[14].n4 VGND 0.04667f
C6005 XThC.Tn[14].n5 VGND 0.12968f
C6006 XThC.Tn[14].t11 VGND 0.01419f
C6007 XThC.Tn[14].t10 VGND 0.01419f
C6008 XThC.Tn[14].n6 VGND 0.04309f
C6009 XThC.Tn[14].t9 VGND 0.01419f
C6010 XThC.Tn[14].t8 VGND 0.01419f
C6011 XThC.Tn[14].n7 VGND 0.03155f
C6012 XThC.Tn[14].n8 VGND 0.14042f
C6013 XThC.Tn[14].n9 VGND 0.02039f
C6014 XThC.Tn[14].t43 VGND 0.01125f
C6015 XThC.Tn[14].t38 VGND 0.01229f
C6016 XThC.Tn[14].n10 VGND 0.02744f
C6017 XThC.Tn[14].n11 VGND 0.01568f
C6018 XThC.Tn[14].n12 VGND 0.01907f
C6019 XThC.Tn[14].t29 VGND 0.01125f
C6020 XThC.Tn[14].t22 VGND 0.01229f
C6021 XThC.Tn[14].n13 VGND 0.02744f
C6022 XThC.Tn[14].n14 VGND 0.01568f
C6023 XThC.Tn[14].n15 VGND 0.09061f
C6024 XThC.Tn[14].t32 VGND 0.01125f
C6025 XThC.Tn[14].t25 VGND 0.01229f
C6026 XThC.Tn[14].n16 VGND 0.02744f
C6027 XThC.Tn[14].n17 VGND 0.01568f
C6028 XThC.Tn[14].n18 VGND 0.09061f
C6029 XThC.Tn[14].t34 VGND 0.01125f
C6030 XThC.Tn[14].t26 VGND 0.01229f
C6031 XThC.Tn[14].n19 VGND 0.02744f
C6032 XThC.Tn[14].n20 VGND 0.01568f
C6033 XThC.Tn[14].n21 VGND 0.09061f
C6034 XThC.Tn[14].t20 VGND 0.01125f
C6035 XThC.Tn[14].t14 VGND 0.01229f
C6036 XThC.Tn[14].n22 VGND 0.02744f
C6037 XThC.Tn[14].n23 VGND 0.01568f
C6038 XThC.Tn[14].n24 VGND 0.09061f
C6039 XThC.Tn[14].t23 VGND 0.01125f
C6040 XThC.Tn[14].t17 VGND 0.01229f
C6041 XThC.Tn[14].n25 VGND 0.02744f
C6042 XThC.Tn[14].n26 VGND 0.01568f
C6043 XThC.Tn[14].n27 VGND 0.09061f
C6044 XThC.Tn[14].t37 VGND 0.01125f
C6045 XThC.Tn[14].t31 VGND 0.01229f
C6046 XThC.Tn[14].n28 VGND 0.02744f
C6047 XThC.Tn[14].n29 VGND 0.01568f
C6048 XThC.Tn[14].n30 VGND 0.09061f
C6049 XThC.Tn[14].t13 VGND 0.01125f
C6050 XThC.Tn[14].t39 VGND 0.01229f
C6051 XThC.Tn[14].n31 VGND 0.02744f
C6052 XThC.Tn[14].n32 VGND 0.01568f
C6053 XThC.Tn[14].n33 VGND 0.09061f
C6054 XThC.Tn[14].t15 VGND 0.01125f
C6055 XThC.Tn[14].t41 VGND 0.01229f
C6056 XThC.Tn[14].n34 VGND 0.02744f
C6057 XThC.Tn[14].n35 VGND 0.01568f
C6058 XThC.Tn[14].n36 VGND 0.09061f
C6059 XThC.Tn[14].t35 VGND 0.01125f
C6060 XThC.Tn[14].t27 VGND 0.01229f
C6061 XThC.Tn[14].n37 VGND 0.02744f
C6062 XThC.Tn[14].n38 VGND 0.01568f
C6063 XThC.Tn[14].n39 VGND 0.09061f
C6064 XThC.Tn[14].t36 VGND 0.01125f
C6065 XThC.Tn[14].t30 VGND 0.01229f
C6066 XThC.Tn[14].n40 VGND 0.02744f
C6067 XThC.Tn[14].n41 VGND 0.01568f
C6068 XThC.Tn[14].n42 VGND 0.09061f
C6069 XThC.Tn[14].t16 VGND 0.01125f
C6070 XThC.Tn[14].t42 VGND 0.01229f
C6071 XThC.Tn[14].n43 VGND 0.02744f
C6072 XThC.Tn[14].n44 VGND 0.01568f
C6073 XThC.Tn[14].n45 VGND 0.09061f
C6074 XThC.Tn[14].t24 VGND 0.01125f
C6075 XThC.Tn[14].t19 VGND 0.01229f
C6076 XThC.Tn[14].n46 VGND 0.02744f
C6077 XThC.Tn[14].n47 VGND 0.01568f
C6078 XThC.Tn[14].n48 VGND 0.09061f
C6079 XThC.Tn[14].t28 VGND 0.01125f
C6080 XThC.Tn[14].t21 VGND 0.01229f
C6081 XThC.Tn[14].n49 VGND 0.02744f
C6082 XThC.Tn[14].n50 VGND 0.01568f
C6083 XThC.Tn[14].n51 VGND 0.09061f
C6084 XThC.Tn[14].t40 VGND 0.01125f
C6085 XThC.Tn[14].t33 VGND 0.01229f
C6086 XThC.Tn[14].n52 VGND 0.02744f
C6087 XThC.Tn[14].n53 VGND 0.01568f
C6088 XThC.Tn[14].n54 VGND 0.09061f
C6089 XThC.Tn[14].t18 VGND 0.01125f
C6090 XThC.Tn[14].t12 VGND 0.01229f
C6091 XThC.Tn[14].n55 VGND 0.02744f
C6092 XThC.Tn[14].n56 VGND 0.01568f
C6093 XThC.Tn[14].n57 VGND 0.09061f
C6094 XThC.Tn[14].n58 VGND 0.54091f
C6095 XThC.Tn[14].n59 VGND 0.03454f
C6096 XThR.Tn[10].t10 VGND 0.01941f
C6097 XThR.Tn[10].t8 VGND 0.01941f
C6098 XThR.Tn[10].n0 VGND 0.05892f
C6099 XThR.Tn[10].t11 VGND 0.01941f
C6100 XThR.Tn[10].t9 VGND 0.01941f
C6101 XThR.Tn[10].n1 VGND 0.04314f
C6102 XThR.Tn[10].n2 VGND 0.19615f
C6103 XThR.Tn[10].t6 VGND 0.01941f
C6104 XThR.Tn[10].t4 VGND 0.01941f
C6105 XThR.Tn[10].n3 VGND 0.04193f
C6106 XThR.Tn[10].t7 VGND 0.01941f
C6107 XThR.Tn[10].t5 VGND 0.01941f
C6108 XThR.Tn[10].n4 VGND 0.06382f
C6109 XThR.Tn[10].n5 VGND 0.1772f
C6110 XThR.Tn[10].t54 VGND 0.01517f
C6111 XThR.Tn[10].t47 VGND 0.01661f
C6112 XThR.Tn[10].n7 VGND 0.04056f
C6113 XThR.Tn[10].n8 VGND 0.07791f
C6114 XThR.Tn[10].t13 VGND 0.01517f
C6115 XThR.Tn[10].t63 VGND 0.01661f
C6116 XThR.Tn[10].n9 VGND 0.04056f
C6117 XThR.Tn[10].t50 VGND 0.01512f
C6118 XThR.Tn[10].t60 VGND 0.01655f
C6119 XThR.Tn[10].n10 VGND 0.0422f
C6120 XThR.Tn[10].n11 VGND 0.02964f
C6121 XThR.Tn[10].n13 VGND 0.09513f
C6122 XThR.Tn[10].t48 VGND 0.01517f
C6123 XThR.Tn[10].t41 VGND 0.01661f
C6124 XThR.Tn[10].n14 VGND 0.04056f
C6125 XThR.Tn[10].t23 VGND 0.01512f
C6126 XThR.Tn[10].t36 VGND 0.01655f
C6127 XThR.Tn[10].n15 VGND 0.0422f
C6128 XThR.Tn[10].n16 VGND 0.02964f
C6129 XThR.Tn[10].n18 VGND 0.09513f
C6130 XThR.Tn[10].t65 VGND 0.01517f
C6131 XThR.Tn[10].t58 VGND 0.01661f
C6132 XThR.Tn[10].n19 VGND 0.04056f
C6133 XThR.Tn[10].t40 VGND 0.01512f
C6134 XThR.Tn[10].t55 VGND 0.01655f
C6135 XThR.Tn[10].n20 VGND 0.0422f
C6136 XThR.Tn[10].n21 VGND 0.02964f
C6137 XThR.Tn[10].n23 VGND 0.09513f
C6138 XThR.Tn[10].t30 VGND 0.01517f
C6139 XThR.Tn[10].t26 VGND 0.01661f
C6140 XThR.Tn[10].n24 VGND 0.04056f
C6141 XThR.Tn[10].t70 VGND 0.01512f
C6142 XThR.Tn[10].t21 VGND 0.01655f
C6143 XThR.Tn[10].n25 VGND 0.0422f
C6144 XThR.Tn[10].n26 VGND 0.02964f
C6145 XThR.Tn[10].n28 VGND 0.09513f
C6146 XThR.Tn[10].t67 VGND 0.01517f
C6147 XThR.Tn[10].t59 VGND 0.01661f
C6148 XThR.Tn[10].n29 VGND 0.04056f
C6149 XThR.Tn[10].t42 VGND 0.01512f
C6150 XThR.Tn[10].t56 VGND 0.01655f
C6151 XThR.Tn[10].n30 VGND 0.0422f
C6152 XThR.Tn[10].n31 VGND 0.02964f
C6153 XThR.Tn[10].n33 VGND 0.09513f
C6154 XThR.Tn[10].t44 VGND 0.01517f
C6155 XThR.Tn[10].t15 VGND 0.01661f
C6156 XThR.Tn[10].n34 VGND 0.04056f
C6157 XThR.Tn[10].t18 VGND 0.01512f
C6158 XThR.Tn[10].t12 VGND 0.01655f
C6159 XThR.Tn[10].n35 VGND 0.0422f
C6160 XThR.Tn[10].n36 VGND 0.02964f
C6161 XThR.Tn[10].n38 VGND 0.09513f
C6162 XThR.Tn[10].t14 VGND 0.01517f
C6163 XThR.Tn[10].t69 VGND 0.01661f
C6164 XThR.Tn[10].n39 VGND 0.04056f
C6165 XThR.Tn[10].t51 VGND 0.01512f
C6166 XThR.Tn[10].t66 VGND 0.01655f
C6167 XThR.Tn[10].n40 VGND 0.0422f
C6168 XThR.Tn[10].n41 VGND 0.02964f
C6169 XThR.Tn[10].n43 VGND 0.09513f
C6170 XThR.Tn[10].t17 VGND 0.01517f
C6171 XThR.Tn[10].t24 VGND 0.01661f
C6172 XThR.Tn[10].n44 VGND 0.04056f
C6173 XThR.Tn[10].t53 VGND 0.01512f
C6174 XThR.Tn[10].t20 VGND 0.01655f
C6175 XThR.Tn[10].n45 VGND 0.0422f
C6176 XThR.Tn[10].n46 VGND 0.02964f
C6177 XThR.Tn[10].n48 VGND 0.09513f
C6178 XThR.Tn[10].t33 VGND 0.01517f
C6179 XThR.Tn[10].t43 VGND 0.01661f
C6180 XThR.Tn[10].n49 VGND 0.04056f
C6181 XThR.Tn[10].t73 VGND 0.01512f
C6182 XThR.Tn[10].t38 VGND 0.01655f
C6183 XThR.Tn[10].n50 VGND 0.0422f
C6184 XThR.Tn[10].n51 VGND 0.02964f
C6185 XThR.Tn[10].n53 VGND 0.09513f
C6186 XThR.Tn[10].t28 VGND 0.01517f
C6187 XThR.Tn[10].t61 VGND 0.01661f
C6188 XThR.Tn[10].n54 VGND 0.04056f
C6189 XThR.Tn[10].t62 VGND 0.01512f
C6190 XThR.Tn[10].t57 VGND 0.01655f
C6191 XThR.Tn[10].n55 VGND 0.0422f
C6192 XThR.Tn[10].n56 VGND 0.02964f
C6193 XThR.Tn[10].n58 VGND 0.09513f
C6194 XThR.Tn[10].t46 VGND 0.01517f
C6195 XThR.Tn[10].t35 VGND 0.01661f
C6196 XThR.Tn[10].n59 VGND 0.04056f
C6197 XThR.Tn[10].t19 VGND 0.01512f
C6198 XThR.Tn[10].t32 VGND 0.01655f
C6199 XThR.Tn[10].n60 VGND 0.0422f
C6200 XThR.Tn[10].n61 VGND 0.02964f
C6201 XThR.Tn[10].n63 VGND 0.09513f
C6202 XThR.Tn[10].t16 VGND 0.01517f
C6203 XThR.Tn[10].t72 VGND 0.01661f
C6204 XThR.Tn[10].n64 VGND 0.04056f
C6205 XThR.Tn[10].t52 VGND 0.01512f
C6206 XThR.Tn[10].t68 VGND 0.01655f
C6207 XThR.Tn[10].n65 VGND 0.0422f
C6208 XThR.Tn[10].n66 VGND 0.02964f
C6209 XThR.Tn[10].n68 VGND 0.09513f
C6210 XThR.Tn[10].t31 VGND 0.01517f
C6211 XThR.Tn[10].t27 VGND 0.01661f
C6212 XThR.Tn[10].n69 VGND 0.04056f
C6213 XThR.Tn[10].t71 VGND 0.01512f
C6214 XThR.Tn[10].t22 VGND 0.01655f
C6215 XThR.Tn[10].n70 VGND 0.0422f
C6216 XThR.Tn[10].n71 VGND 0.02964f
C6217 XThR.Tn[10].n73 VGND 0.09513f
C6218 XThR.Tn[10].t49 VGND 0.01517f
C6219 XThR.Tn[10].t45 VGND 0.01661f
C6220 XThR.Tn[10].n74 VGND 0.04056f
C6221 XThR.Tn[10].t25 VGND 0.01512f
C6222 XThR.Tn[10].t39 VGND 0.01655f
C6223 XThR.Tn[10].n75 VGND 0.0422f
C6224 XThR.Tn[10].n76 VGND 0.02964f
C6225 XThR.Tn[10].n78 VGND 0.09513f
C6226 XThR.Tn[10].t29 VGND 0.01517f
C6227 XThR.Tn[10].t37 VGND 0.01661f
C6228 XThR.Tn[10].n79 VGND 0.04056f
C6229 XThR.Tn[10].t64 VGND 0.01512f
C6230 XThR.Tn[10].t34 VGND 0.01655f
C6231 XThR.Tn[10].n80 VGND 0.0422f
C6232 XThR.Tn[10].n81 VGND 0.02964f
C6233 XThR.Tn[10].n83 VGND 0.09513f
C6234 XThR.Tn[10].n84 VGND 0.08645f
C6235 XThR.Tn[10].n85 VGND 0.26614f
C6236 XThR.Tn[10].t0 VGND 0.01261f
C6237 XThR.Tn[10].t2 VGND 0.01261f
C6238 XThR.Tn[10].n86 VGND 0.02523f
C6239 XThR.Tn[10].t1 VGND 0.01261f
C6240 XThR.Tn[10].t3 VGND 0.01261f
C6241 XThR.Tn[10].n87 VGND 0.03146f
C6242 XThR.Tn[10].n88 VGND 0.05817f
C6243 XThC.Tn[3].t1 VGND 0.01185f
C6244 XThC.Tn[3].t0 VGND 0.01185f
C6245 XThC.Tn[3].n0 VGND 0.02391f
C6246 XThC.Tn[3].t3 VGND 0.01185f
C6247 XThC.Tn[3].t2 VGND 0.01185f
C6248 XThC.Tn[3].n1 VGND 0.02797f
C6249 XThC.Tn[3].n2 VGND 0.08391f
C6250 XThC.Tn[3].n3 VGND 0.02921f
C6251 XThC.Tn[3].n4 VGND 0.01753f
C6252 XThC.Tn[3].n5 VGND 0.0835f
C6253 XThC.Tn[3].n6 VGND 0.01753f
C6254 XThC.Tn[3].n7 VGND 0.05162f
C6255 XThC.Tn[3].n8 VGND 0.01753f
C6256 XThC.Tn[3].n9 VGND 0.05825f
C6257 XThC.Tn[3].t42 VGND 0.01025f
C6258 XThC.Tn[3].n10 VGND 0.0229f
C6259 XThC.Tn[3].n11 VGND 0.01309f
C6260 XThC.Tn[3].n12 VGND 0.01592f
C6261 XThC.Tn[3].t27 VGND 0.01025f
C6262 XThC.Tn[3].n13 VGND 0.0229f
C6263 XThC.Tn[3].n14 VGND 0.01309f
C6264 XThC.Tn[3].n15 VGND 0.07562f
C6265 XThC.Tn[3].t29 VGND 0.01025f
C6266 XThC.Tn[3].n16 VGND 0.0229f
C6267 XThC.Tn[3].n17 VGND 0.01309f
C6268 XThC.Tn[3].n18 VGND 0.07562f
C6269 XThC.Tn[3].t31 VGND 0.01025f
C6270 XThC.Tn[3].n19 VGND 0.0229f
C6271 XThC.Tn[3].n20 VGND 0.01309f
C6272 XThC.Tn[3].n21 VGND 0.07562f
C6273 XThC.Tn[3].t20 VGND 0.01025f
C6274 XThC.Tn[3].n22 VGND 0.0229f
C6275 XThC.Tn[3].n23 VGND 0.01309f
C6276 XThC.Tn[3].n24 VGND 0.07562f
C6277 XThC.Tn[3].t21 VGND 0.01025f
C6278 XThC.Tn[3].n25 VGND 0.0229f
C6279 XThC.Tn[3].n26 VGND 0.01309f
C6280 XThC.Tn[3].n27 VGND 0.07562f
C6281 XThC.Tn[3].t34 VGND 0.01025f
C6282 XThC.Tn[3].n28 VGND 0.0229f
C6283 XThC.Tn[3].n29 VGND 0.01309f
C6284 XThC.Tn[3].n30 VGND 0.07562f
C6285 XThC.Tn[3].t43 VGND 0.01025f
C6286 XThC.Tn[3].n31 VGND 0.0229f
C6287 XThC.Tn[3].n32 VGND 0.01309f
C6288 XThC.Tn[3].n33 VGND 0.07562f
C6289 XThC.Tn[3].t13 VGND 0.01025f
C6290 XThC.Tn[3].n34 VGND 0.0229f
C6291 XThC.Tn[3].n35 VGND 0.01309f
C6292 XThC.Tn[3].n36 VGND 0.07562f
C6293 XThC.Tn[3].t32 VGND 0.01025f
C6294 XThC.Tn[3].n37 VGND 0.0229f
C6295 XThC.Tn[3].n38 VGND 0.01309f
C6296 XThC.Tn[3].n39 VGND 0.07562f
C6297 XThC.Tn[3].t33 VGND 0.01025f
C6298 XThC.Tn[3].n40 VGND 0.0229f
C6299 XThC.Tn[3].n41 VGND 0.01309f
C6300 XThC.Tn[3].n42 VGND 0.07562f
C6301 XThC.Tn[3].t14 VGND 0.01025f
C6302 XThC.Tn[3].n43 VGND 0.0229f
C6303 XThC.Tn[3].n44 VGND 0.01309f
C6304 XThC.Tn[3].n45 VGND 0.07562f
C6305 XThC.Tn[3].t22 VGND 0.01025f
C6306 XThC.Tn[3].n46 VGND 0.0229f
C6307 XThC.Tn[3].n47 VGND 0.01309f
C6308 XThC.Tn[3].n48 VGND 0.07562f
C6309 XThC.Tn[3].t25 VGND 0.01025f
C6310 XThC.Tn[3].n49 VGND 0.0229f
C6311 XThC.Tn[3].n50 VGND 0.01309f
C6312 XThC.Tn[3].n51 VGND 0.07562f
C6313 XThC.Tn[3].t38 VGND 0.01025f
C6314 XThC.Tn[3].n52 VGND 0.0229f
C6315 XThC.Tn[3].n53 VGND 0.01309f
C6316 XThC.Tn[3].n54 VGND 0.07562f
C6317 XThC.Tn[3].t16 VGND 0.01025f
C6318 XThC.Tn[3].n55 VGND 0.0229f
C6319 XThC.Tn[3].n56 VGND 0.01309f
C6320 XThC.Tn[3].n57 VGND 0.07562f
C6321 XThC.Tn[3].n58 VGND 0.03994f
C6322 XThC.Tn[1].t7 VGND 0.0116f
C6323 XThC.Tn[1].t6 VGND 0.0116f
C6324 XThC.Tn[1].n0 VGND 0.02342f
C6325 XThC.Tn[1].t5 VGND 0.0116f
C6326 XThC.Tn[1].t4 VGND 0.0116f
C6327 XThC.Tn[1].n1 VGND 0.02741f
C6328 XThC.Tn[1].n2 VGND 0.08221f
C6329 XThC.Tn[1].n3 VGND 0.01718f
C6330 XThC.Tn[1].n4 VGND 0.01718f
C6331 XThC.Tn[1].n5 VGND 0.01718f
C6332 XThC.Tn[1].n6 VGND 0.02862f
C6333 XThC.Tn[1].n7 VGND 0.0818f
C6334 XThC.Tn[1].n8 VGND 0.05057f
C6335 XThC.Tn[1].n9 VGND 0.05707f
C6336 XThC.Tn[1].t29 VGND 0.01005f
C6337 XThC.Tn[1].n10 VGND 0.02244f
C6338 XThC.Tn[1].n11 VGND 0.01282f
C6339 XThC.Tn[1].n12 VGND 0.01559f
C6340 XThC.Tn[1].t14 VGND 0.01005f
C6341 XThC.Tn[1].n13 VGND 0.02244f
C6342 XThC.Tn[1].n14 VGND 0.01282f
C6343 XThC.Tn[1].n15 VGND 0.07408f
C6344 XThC.Tn[1].t16 VGND 0.01005f
C6345 XThC.Tn[1].n16 VGND 0.02244f
C6346 XThC.Tn[1].n17 VGND 0.01282f
C6347 XThC.Tn[1].n18 VGND 0.07408f
C6348 XThC.Tn[1].t18 VGND 0.01005f
C6349 XThC.Tn[1].n19 VGND 0.02244f
C6350 XThC.Tn[1].n20 VGND 0.01282f
C6351 XThC.Tn[1].n21 VGND 0.07408f
C6352 XThC.Tn[1].t39 VGND 0.01005f
C6353 XThC.Tn[1].n22 VGND 0.02244f
C6354 XThC.Tn[1].n23 VGND 0.01282f
C6355 XThC.Tn[1].n24 VGND 0.07408f
C6356 XThC.Tn[1].t40 VGND 0.01005f
C6357 XThC.Tn[1].n25 VGND 0.02244f
C6358 XThC.Tn[1].n26 VGND 0.01282f
C6359 XThC.Tn[1].n27 VGND 0.07408f
C6360 XThC.Tn[1].t21 VGND 0.01005f
C6361 XThC.Tn[1].n28 VGND 0.02244f
C6362 XThC.Tn[1].n29 VGND 0.01282f
C6363 XThC.Tn[1].n30 VGND 0.07408f
C6364 XThC.Tn[1].t30 VGND 0.01005f
C6365 XThC.Tn[1].n31 VGND 0.02244f
C6366 XThC.Tn[1].n32 VGND 0.01282f
C6367 XThC.Tn[1].n33 VGND 0.07408f
C6368 XThC.Tn[1].t32 VGND 0.01005f
C6369 XThC.Tn[1].n34 VGND 0.02244f
C6370 XThC.Tn[1].n35 VGND 0.01282f
C6371 XThC.Tn[1].n36 VGND 0.07408f
C6372 XThC.Tn[1].t19 VGND 0.01005f
C6373 XThC.Tn[1].n37 VGND 0.02244f
C6374 XThC.Tn[1].n38 VGND 0.01282f
C6375 XThC.Tn[1].n39 VGND 0.07408f
C6376 XThC.Tn[1].t20 VGND 0.01005f
C6377 XThC.Tn[1].n40 VGND 0.02244f
C6378 XThC.Tn[1].n41 VGND 0.01282f
C6379 XThC.Tn[1].n42 VGND 0.07408f
C6380 XThC.Tn[1].t33 VGND 0.01005f
C6381 XThC.Tn[1].n43 VGND 0.02244f
C6382 XThC.Tn[1].n44 VGND 0.01282f
C6383 XThC.Tn[1].n45 VGND 0.07408f
C6384 XThC.Tn[1].t41 VGND 0.01005f
C6385 XThC.Tn[1].n46 VGND 0.02244f
C6386 XThC.Tn[1].n47 VGND 0.01282f
C6387 XThC.Tn[1].n48 VGND 0.07408f
C6388 XThC.Tn[1].t12 VGND 0.01005f
C6389 XThC.Tn[1].n49 VGND 0.02244f
C6390 XThC.Tn[1].n50 VGND 0.01282f
C6391 XThC.Tn[1].n51 VGND 0.07408f
C6392 XThC.Tn[1].t25 VGND 0.01005f
C6393 XThC.Tn[1].n52 VGND 0.02244f
C6394 XThC.Tn[1].n53 VGND 0.01282f
C6395 XThC.Tn[1].n54 VGND 0.07408f
C6396 XThC.Tn[1].t35 VGND 0.01005f
C6397 XThC.Tn[1].n55 VGND 0.02244f
C6398 XThC.Tn[1].n56 VGND 0.01282f
C6399 XThC.Tn[1].n57 VGND 0.07408f
C6400 XThC.Tn[1].n58 VGND 0.27353f
C6401 XThC.Tn[1].n59 VGND 0.0276f
C6402 Vbias.t260 VGND 0.17882f
C6403 Vbias.n0 VGND 0.19466f
C6404 Vbias.t79 VGND 0.17882f
C6405 Vbias.n1 VGND 0.19501f
C6406 Vbias.n2 VGND 0.12932f
C6407 Vbias.t174 VGND 0.17882f
C6408 Vbias.n3 VGND 0.19501f
C6409 Vbias.n4 VGND 0.12932f
C6410 Vbias.t182 VGND 0.17882f
C6411 Vbias.n5 VGND 0.19501f
C6412 Vbias.n6 VGND 0.12932f
C6413 Vbias.t15 VGND 0.17882f
C6414 Vbias.n7 VGND 0.19501f
C6415 Vbias.n8 VGND 0.12932f
C6416 Vbias.t101 VGND 0.17882f
C6417 Vbias.n9 VGND 0.19501f
C6418 Vbias.n10 VGND 0.12932f
C6419 Vbias.t184 VGND 0.17882f
C6420 Vbias.n11 VGND 0.19501f
C6421 Vbias.n12 VGND 0.12932f
C6422 Vbias.t19 VGND 0.17882f
C6423 Vbias.n13 VGND 0.19501f
C6424 Vbias.n14 VGND 0.12932f
C6425 Vbias.t39 VGND 0.17882f
C6426 Vbias.n15 VGND 0.19501f
C6427 Vbias.n16 VGND 0.12932f
C6428 Vbias.t111 VGND 0.17882f
C6429 Vbias.n17 VGND 0.19501f
C6430 Vbias.n18 VGND 0.12932f
C6431 Vbias.t202 VGND 0.17882f
C6432 Vbias.n19 VGND 0.19501f
C6433 Vbias.n20 VGND 0.12932f
C6434 Vbias.t223 VGND 0.17882f
C6435 Vbias.n21 VGND 0.19501f
C6436 Vbias.n22 VGND 0.12932f
C6437 Vbias.t114 VGND 0.17882f
C6438 Vbias.n23 VGND 0.19501f
C6439 Vbias.n24 VGND 0.12932f
C6440 Vbias.t142 VGND 0.17882f
C6441 Vbias.n25 VGND 0.19501f
C6442 Vbias.n26 VGND 0.12932f
C6443 Vbias.t151 VGND 0.17882f
C6444 Vbias.n27 VGND 0.19501f
C6445 Vbias.n28 VGND 0.12932f
C6446 Vbias.t61 VGND 0.17882f
C6447 Vbias.n29 VGND 0.19501f
C6448 Vbias.n30 VGND 0.12932f
C6449 Vbias.n31 VGND 0.54269f
C6450 Vbias.t140 VGND 0.17882f
C6451 Vbias.n32 VGND 0.19466f
C6452 Vbias.t216 VGND 0.17882f
C6453 Vbias.n33 VGND 0.19501f
C6454 Vbias.n34 VGND 0.12932f
C6455 Vbias.t59 VGND 0.17882f
C6456 Vbias.n35 VGND 0.19501f
C6457 Vbias.n36 VGND 0.12932f
C6458 Vbias.t67 VGND 0.17882f
C6459 Vbias.n37 VGND 0.19501f
C6460 Vbias.n38 VGND 0.12932f
C6461 Vbias.t152 VGND 0.17882f
C6462 Vbias.n39 VGND 0.19501f
C6463 Vbias.n40 VGND 0.12932f
C6464 Vbias.t245 VGND 0.17882f
C6465 Vbias.n41 VGND 0.19501f
C6466 Vbias.n42 VGND 0.12932f
C6467 Vbias.t72 VGND 0.17882f
C6468 Vbias.n43 VGND 0.19501f
C6469 Vbias.n44 VGND 0.12932f
C6470 Vbias.t158 VGND 0.17882f
C6471 Vbias.n45 VGND 0.19501f
C6472 Vbias.n46 VGND 0.12932f
C6473 Vbias.t178 VGND 0.17882f
C6474 Vbias.n47 VGND 0.19501f
C6475 Vbias.n48 VGND 0.12932f
C6476 Vbias.t254 VGND 0.17882f
C6477 Vbias.n49 VGND 0.19501f
C6478 Vbias.n50 VGND 0.12932f
C6479 Vbias.t84 VGND 0.17882f
C6480 Vbias.n51 VGND 0.19501f
C6481 Vbias.n52 VGND 0.12932f
C6482 Vbias.t106 VGND 0.17882f
C6483 Vbias.n53 VGND 0.19501f
C6484 Vbias.n54 VGND 0.12932f
C6485 Vbias.t259 VGND 0.17882f
C6486 Vbias.n55 VGND 0.19501f
C6487 Vbias.n56 VGND 0.12932f
C6488 Vbias.t26 VGND 0.17882f
C6489 Vbias.n57 VGND 0.19501f
C6490 Vbias.n58 VGND 0.12932f
C6491 Vbias.t35 VGND 0.17882f
C6492 Vbias.n59 VGND 0.19501f
C6493 Vbias.n60 VGND 0.12932f
C6494 Vbias.t194 VGND 0.17882f
C6495 Vbias.n61 VGND 0.19501f
C6496 Vbias.n62 VGND 0.12932f
C6497 Vbias.n63 VGND 0.55831f
C6498 Vbias.t215 VGND 0.17882f
C6499 Vbias.n64 VGND 0.19466f
C6500 Vbias.t31 VGND 0.17882f
C6501 Vbias.n65 VGND 0.19501f
C6502 Vbias.n66 VGND 0.12932f
C6503 Vbias.t132 VGND 0.17882f
C6504 Vbias.n67 VGND 0.19501f
C6505 Vbias.n68 VGND 0.12932f
C6506 Vbias.t139 VGND 0.17882f
C6507 Vbias.n69 VGND 0.19501f
C6508 Vbias.n70 VGND 0.12932f
C6509 Vbias.t224 VGND 0.17882f
C6510 Vbias.n71 VGND 0.19501f
C6511 Vbias.n72 VGND 0.12932f
C6512 Vbias.t58 VGND 0.17882f
C6513 Vbias.n73 VGND 0.19501f
C6514 Vbias.n74 VGND 0.12932f
C6515 Vbias.t145 VGND 0.17882f
C6516 Vbias.n75 VGND 0.19501f
C6517 Vbias.n76 VGND 0.12932f
C6518 Vbias.t230 VGND 0.17882f
C6519 Vbias.n77 VGND 0.19501f
C6520 Vbias.n78 VGND 0.12932f
C6521 Vbias.t253 VGND 0.17882f
C6522 Vbias.n79 VGND 0.19501f
C6523 Vbias.n80 VGND 0.12932f
C6524 Vbias.t71 VGND 0.17882f
C6525 Vbias.n81 VGND 0.19501f
C6526 Vbias.n82 VGND 0.12932f
C6527 Vbias.t157 VGND 0.17882f
C6528 Vbias.n83 VGND 0.19501f
C6529 Vbias.n84 VGND 0.12932f
C6530 Vbias.t177 VGND 0.17882f
C6531 Vbias.n85 VGND 0.19501f
C6532 Vbias.n86 VGND 0.12932f
C6533 Vbias.t77 VGND 0.17882f
C6534 Vbias.n87 VGND 0.19501f
C6535 Vbias.n88 VGND 0.12932f
C6536 Vbias.t97 VGND 0.17882f
C6537 Vbias.n89 VGND 0.19501f
C6538 Vbias.n90 VGND 0.12932f
C6539 Vbias.t104 VGND 0.17882f
C6540 Vbias.n91 VGND 0.19501f
C6541 Vbias.n92 VGND 0.12932f
C6542 Vbias.t13 VGND 0.17882f
C6543 Vbias.n93 VGND 0.19501f
C6544 Vbias.n94 VGND 0.12932f
C6545 Vbias.n95 VGND 0.55831f
C6546 Vbias.t30 VGND 0.17882f
C6547 Vbias.n96 VGND 0.19466f
C6548 Vbias.t100 VGND 0.17882f
C6549 Vbias.n97 VGND 0.19501f
C6550 Vbias.n98 VGND 0.12932f
C6551 Vbias.t203 VGND 0.17882f
C6552 Vbias.n99 VGND 0.19501f
C6553 Vbias.n100 VGND 0.12932f
C6554 Vbias.t214 VGND 0.17882f
C6555 Vbias.n101 VGND 0.19501f
C6556 Vbias.n102 VGND 0.12932f
C6557 Vbias.t38 VGND 0.17882f
C6558 Vbias.n103 VGND 0.19501f
C6559 Vbias.n104 VGND 0.12932f
C6560 Vbias.t131 VGND 0.17882f
C6561 Vbias.n105 VGND 0.19501f
C6562 Vbias.n106 VGND 0.12932f
C6563 Vbias.t218 VGND 0.17882f
C6564 Vbias.n107 VGND 0.19501f
C6565 Vbias.n108 VGND 0.12932f
C6566 Vbias.t42 VGND 0.17882f
C6567 Vbias.n109 VGND 0.19501f
C6568 Vbias.n110 VGND 0.12932f
C6569 Vbias.t70 VGND 0.17882f
C6570 Vbias.n111 VGND 0.19501f
C6571 Vbias.n112 VGND 0.12932f
C6572 Vbias.t143 VGND 0.17882f
C6573 Vbias.n113 VGND 0.19501f
C6574 Vbias.n114 VGND 0.12932f
C6575 Vbias.t228 VGND 0.17882f
C6576 Vbias.n115 VGND 0.19501f
C6577 Vbias.n116 VGND 0.12932f
C6578 Vbias.t252 VGND 0.17882f
C6579 Vbias.n117 VGND 0.19501f
C6580 Vbias.n118 VGND 0.12932f
C6581 Vbias.t148 VGND 0.17882f
C6582 Vbias.n119 VGND 0.19501f
C6583 Vbias.n120 VGND 0.12932f
C6584 Vbias.t170 VGND 0.17882f
C6585 Vbias.n121 VGND 0.19501f
C6586 Vbias.n122 VGND 0.12932f
C6587 Vbias.t175 VGND 0.17882f
C6588 Vbias.n123 VGND 0.19501f
C6589 Vbias.n124 VGND 0.12932f
C6590 Vbias.t86 VGND 0.17882f
C6591 Vbias.n125 VGND 0.19501f
C6592 Vbias.n126 VGND 0.12932f
C6593 Vbias.n127 VGND 0.55831f
C6594 Vbias.t186 VGND 0.17882f
C6595 Vbias.n128 VGND 0.19466f
C6596 Vbias.t6 VGND 0.17882f
C6597 Vbias.n129 VGND 0.19501f
C6598 Vbias.n130 VGND 0.12932f
C6599 Vbias.t103 VGND 0.17882f
C6600 Vbias.n131 VGND 0.19501f
C6601 Vbias.n132 VGND 0.12932f
C6602 Vbias.t115 VGND 0.17882f
C6603 Vbias.n133 VGND 0.19501f
C6604 Vbias.n134 VGND 0.12932f
C6605 Vbias.t206 VGND 0.17882f
C6606 Vbias.n135 VGND 0.19501f
C6607 Vbias.n136 VGND 0.12932f
C6608 Vbias.t34 VGND 0.17882f
C6609 Vbias.n137 VGND 0.19501f
C6610 Vbias.n138 VGND 0.12932f
C6611 Vbias.t116 VGND 0.17882f
C6612 Vbias.n139 VGND 0.19501f
C6613 Vbias.n140 VGND 0.12932f
C6614 Vbias.t209 VGND 0.17882f
C6615 Vbias.n141 VGND 0.19501f
C6616 Vbias.n142 VGND 0.12932f
C6617 Vbias.t231 VGND 0.17882f
C6618 Vbias.n143 VGND 0.19501f
C6619 Vbias.n144 VGND 0.12932f
C6620 Vbias.t43 VGND 0.17882f
C6621 Vbias.n145 VGND 0.19501f
C6622 Vbias.n146 VGND 0.12932f
C6623 Vbias.t134 VGND 0.17882f
C6624 Vbias.n147 VGND 0.19501f
C6625 Vbias.n148 VGND 0.12932f
C6626 Vbias.t159 VGND 0.17882f
C6627 Vbias.n149 VGND 0.19501f
C6628 Vbias.n150 VGND 0.12932f
C6629 Vbias.t47 VGND 0.17882f
C6630 Vbias.n151 VGND 0.19501f
C6631 Vbias.n152 VGND 0.12932f
C6632 Vbias.t78 VGND 0.17882f
C6633 Vbias.n153 VGND 0.19501f
C6634 Vbias.n154 VGND 0.12932f
C6635 Vbias.t85 VGND 0.17882f
C6636 Vbias.n155 VGND 0.19501f
C6637 Vbias.n156 VGND 0.12932f
C6638 Vbias.t249 VGND 0.17882f
C6639 Vbias.n157 VGND 0.19501f
C6640 Vbias.n158 VGND 0.12932f
C6641 Vbias.n159 VGND 0.55831f
C6642 Vbias.t55 VGND 0.17882f
C6643 Vbias.n160 VGND 0.19466f
C6644 Vbias.t128 VGND 0.17882f
C6645 Vbias.n161 VGND 0.19501f
C6646 Vbias.n162 VGND 0.12932f
C6647 Vbias.t226 VGND 0.17882f
C6648 Vbias.n163 VGND 0.19501f
C6649 Vbias.n164 VGND 0.12932f
C6650 Vbias.t241 VGND 0.17882f
C6651 Vbias.n165 VGND 0.19501f
C6652 Vbias.n166 VGND 0.12932f
C6653 Vbias.t66 VGND 0.17882f
C6654 Vbias.n167 VGND 0.19501f
C6655 Vbias.n168 VGND 0.12932f
C6656 Vbias.t155 VGND 0.17882f
C6657 Vbias.n169 VGND 0.19501f
C6658 Vbias.n170 VGND 0.12932f
C6659 Vbias.t244 VGND 0.17882f
C6660 Vbias.n171 VGND 0.19501f
C6661 Vbias.n172 VGND 0.12932f
C6662 Vbias.t74 VGND 0.17882f
C6663 Vbias.n173 VGND 0.19501f
C6664 Vbias.n174 VGND 0.12932f
C6665 Vbias.t94 VGND 0.17882f
C6666 Vbias.n175 VGND 0.19501f
C6667 Vbias.n176 VGND 0.12932f
C6668 Vbias.t167 VGND 0.17882f
C6669 Vbias.n177 VGND 0.19501f
C6670 Vbias.n178 VGND 0.12932f
C6671 Vbias.t256 VGND 0.17882f
C6672 Vbias.n179 VGND 0.19501f
C6673 Vbias.n180 VGND 0.12932f
C6674 Vbias.t22 VGND 0.17882f
C6675 Vbias.n181 VGND 0.19501f
C6676 Vbias.n182 VGND 0.12932f
C6677 Vbias.t172 VGND 0.17882f
C6678 Vbias.n183 VGND 0.19501f
C6679 Vbias.n184 VGND 0.12932f
C6680 Vbias.t191 VGND 0.17882f
C6681 Vbias.n185 VGND 0.19501f
C6682 Vbias.n186 VGND 0.12932f
C6683 Vbias.t207 VGND 0.17882f
C6684 Vbias.n187 VGND 0.19501f
C6685 Vbias.n188 VGND 0.12932f
C6686 Vbias.t109 VGND 0.17882f
C6687 Vbias.n189 VGND 0.19501f
C6688 Vbias.n190 VGND 0.12932f
C6689 Vbias.n191 VGND 0.55831f
C6690 Vbias.t189 VGND 0.17882f
C6691 Vbias.n192 VGND 0.19466f
C6692 Vbias.t10 VGND 0.17882f
C6693 Vbias.n193 VGND 0.19501f
C6694 Vbias.n194 VGND 0.12932f
C6695 Vbias.t108 VGND 0.17882f
C6696 Vbias.n195 VGND 0.19501f
C6697 Vbias.n196 VGND 0.12932f
C6698 Vbias.t117 VGND 0.17882f
C6699 Vbias.n197 VGND 0.19501f
C6700 Vbias.n198 VGND 0.12932f
C6701 Vbias.t208 VGND 0.17882f
C6702 Vbias.n199 VGND 0.19501f
C6703 Vbias.n200 VGND 0.12932f
C6704 Vbias.t36 VGND 0.17882f
C6705 Vbias.n201 VGND 0.19501f
C6706 Vbias.n202 VGND 0.12932f
C6707 Vbias.t120 VGND 0.17882f
C6708 Vbias.n203 VGND 0.19501f
C6709 Vbias.n204 VGND 0.12932f
C6710 Vbias.t212 VGND 0.17882f
C6711 Vbias.n205 VGND 0.19501f
C6712 Vbias.n206 VGND 0.12932f
C6713 Vbias.t234 VGND 0.17882f
C6714 Vbias.n207 VGND 0.19501f
C6715 Vbias.n208 VGND 0.12932f
C6716 Vbias.t46 VGND 0.17882f
C6717 Vbias.n209 VGND 0.19501f
C6718 Vbias.n210 VGND 0.12932f
C6719 Vbias.t136 VGND 0.17882f
C6720 Vbias.n211 VGND 0.19501f
C6721 Vbias.n212 VGND 0.12932f
C6722 Vbias.t162 VGND 0.17882f
C6723 Vbias.n213 VGND 0.19501f
C6724 Vbias.n214 VGND 0.12932f
C6725 Vbias.t51 VGND 0.17882f
C6726 Vbias.n215 VGND 0.19501f
C6727 Vbias.n216 VGND 0.12932f
C6728 Vbias.t80 VGND 0.17882f
C6729 Vbias.n217 VGND 0.19501f
C6730 Vbias.n218 VGND 0.12932f
C6731 Vbias.t89 VGND 0.17882f
C6732 Vbias.n219 VGND 0.19501f
C6733 Vbias.n220 VGND 0.12932f
C6734 Vbias.t250 VGND 0.17882f
C6735 Vbias.n221 VGND 0.19501f
C6736 Vbias.n222 VGND 0.12932f
C6737 Vbias.n223 VGND 0.55831f
C6738 Vbias.t9 VGND 0.17882f
C6739 Vbias.n224 VGND 0.19466f
C6740 Vbias.t83 VGND 0.17882f
C6741 Vbias.n225 VGND 0.19501f
C6742 Vbias.n226 VGND 0.12932f
C6743 Vbias.t180 VGND 0.17882f
C6744 Vbias.n227 VGND 0.19501f
C6745 Vbias.n228 VGND 0.12932f
C6746 Vbias.t188 VGND 0.17882f
C6747 Vbias.n229 VGND 0.19501f
C6748 Vbias.n230 VGND 0.12932f
C6749 Vbias.t23 VGND 0.17882f
C6750 Vbias.n231 VGND 0.19501f
C6751 Vbias.n232 VGND 0.12932f
C6752 Vbias.t107 VGND 0.17882f
C6753 Vbias.n233 VGND 0.19501f
C6754 Vbias.n234 VGND 0.12932f
C6755 Vbias.t192 VGND 0.17882f
C6756 Vbias.n235 VGND 0.19501f
C6757 Vbias.n236 VGND 0.12932f
C6758 Vbias.t28 VGND 0.17882f
C6759 Vbias.n237 VGND 0.19501f
C6760 Vbias.n238 VGND 0.12932f
C6761 Vbias.t45 VGND 0.17882f
C6762 Vbias.n239 VGND 0.19501f
C6763 Vbias.n240 VGND 0.12932f
C6764 Vbias.t119 VGND 0.17882f
C6765 Vbias.n241 VGND 0.19501f
C6766 Vbias.n242 VGND 0.12932f
C6767 Vbias.t211 VGND 0.17882f
C6768 Vbias.n243 VGND 0.19501f
C6769 Vbias.n244 VGND 0.12932f
C6770 Vbias.t233 VGND 0.17882f
C6771 Vbias.n245 VGND 0.19501f
C6772 Vbias.n246 VGND 0.12932f
C6773 Vbias.t123 VGND 0.17882f
C6774 Vbias.n247 VGND 0.19501f
C6775 Vbias.n248 VGND 0.12932f
C6776 Vbias.t149 VGND 0.17882f
C6777 Vbias.n249 VGND 0.19501f
C6778 Vbias.n250 VGND 0.12932f
C6779 Vbias.t161 VGND 0.17882f
C6780 Vbias.n251 VGND 0.19501f
C6781 Vbias.n252 VGND 0.12932f
C6782 Vbias.t64 VGND 0.17882f
C6783 Vbias.n253 VGND 0.19501f
C6784 Vbias.n254 VGND 0.12932f
C6785 Vbias.n255 VGND 0.55831f
C6786 Vbias.t82 VGND 0.17882f
C6787 Vbias.n256 VGND 0.19466f
C6788 Vbias.t154 VGND 0.17882f
C6789 Vbias.n257 VGND 0.19501f
C6790 Vbias.n258 VGND 0.12932f
C6791 Vbias.t257 VGND 0.17882f
C6792 Vbias.n259 VGND 0.19501f
C6793 Vbias.n260 VGND 0.12932f
C6794 Vbias.t8 VGND 0.17882f
C6795 Vbias.n261 VGND 0.19501f
C6796 Vbias.n262 VGND 0.12932f
C6797 Vbias.t93 VGND 0.17882f
C6798 Vbias.n263 VGND 0.19501f
C6799 Vbias.n264 VGND 0.12932f
C6800 Vbias.t179 VGND 0.17882f
C6801 Vbias.n265 VGND 0.19501f
C6802 Vbias.n266 VGND 0.12932f
C6803 Vbias.t11 VGND 0.17882f
C6804 Vbias.n267 VGND 0.19501f
C6805 Vbias.n268 VGND 0.12932f
C6806 Vbias.t98 VGND 0.17882f
C6807 Vbias.n269 VGND 0.19501f
C6808 Vbias.n270 VGND 0.12932f
C6809 Vbias.t118 VGND 0.17882f
C6810 Vbias.n271 VGND 0.19501f
C6811 Vbias.n272 VGND 0.12932f
C6812 Vbias.t190 VGND 0.17882f
C6813 Vbias.n273 VGND 0.19501f
C6814 Vbias.n274 VGND 0.12932f
C6815 Vbias.t27 VGND 0.17882f
C6816 Vbias.n275 VGND 0.19501f
C6817 Vbias.n276 VGND 0.12932f
C6818 Vbias.t44 VGND 0.17882f
C6819 Vbias.n277 VGND 0.19501f
C6820 Vbias.n278 VGND 0.12932f
C6821 Vbias.t197 VGND 0.17882f
C6822 Vbias.n279 VGND 0.19501f
C6823 Vbias.n280 VGND 0.12932f
C6824 Vbias.t220 VGND 0.17882f
C6825 Vbias.n281 VGND 0.19501f
C6826 Vbias.n282 VGND 0.12932f
C6827 Vbias.t232 VGND 0.17882f
C6828 Vbias.n283 VGND 0.19501f
C6829 Vbias.n284 VGND 0.12932f
C6830 Vbias.t137 VGND 0.17882f
C6831 Vbias.n285 VGND 0.19501f
C6832 Vbias.n286 VGND 0.12932f
C6833 Vbias.n287 VGND 0.55831f
C6834 Vbias.t49 VGND 0.17882f
C6835 Vbias.n288 VGND 0.19466f
C6836 Vbias.t122 VGND 0.17882f
C6837 Vbias.n289 VGND 0.19501f
C6838 Vbias.n290 VGND 0.12932f
C6839 Vbias.t222 VGND 0.17882f
C6840 Vbias.n291 VGND 0.19501f
C6841 Vbias.n292 VGND 0.12932f
C6842 Vbias.t235 VGND 0.17882f
C6843 Vbias.n293 VGND 0.19501f
C6844 Vbias.n294 VGND 0.12932f
C6845 Vbias.t63 VGND 0.17882f
C6846 Vbias.n295 VGND 0.19501f
C6847 Vbias.n296 VGND 0.12932f
C6848 Vbias.t150 VGND 0.17882f
C6849 Vbias.n297 VGND 0.19501f
C6850 Vbias.n298 VGND 0.12932f
C6851 Vbias.t237 VGND 0.17882f
C6852 Vbias.n299 VGND 0.19501f
C6853 Vbias.n300 VGND 0.12932f
C6854 Vbias.t68 VGND 0.17882f
C6855 Vbias.n301 VGND 0.19501f
C6856 Vbias.n302 VGND 0.12932f
C6857 Vbias.t91 VGND 0.17882f
C6858 Vbias.n303 VGND 0.19501f
C6859 Vbias.n304 VGND 0.12932f
C6860 Vbias.t164 VGND 0.17882f
C6861 Vbias.n305 VGND 0.19501f
C6862 Vbias.n306 VGND 0.12932f
C6863 Vbias.t251 VGND 0.17882f
C6864 Vbias.n307 VGND 0.19501f
C6865 Vbias.n308 VGND 0.12932f
C6866 Vbias.t21 VGND 0.17882f
C6867 Vbias.n309 VGND 0.19501f
C6868 Vbias.n310 VGND 0.12932f
C6869 Vbias.t168 VGND 0.17882f
C6870 Vbias.n311 VGND 0.19501f
C6871 Vbias.n312 VGND 0.12932f
C6872 Vbias.t187 VGND 0.17882f
C6873 Vbias.n313 VGND 0.19501f
C6874 Vbias.n314 VGND 0.12932f
C6875 Vbias.t204 VGND 0.17882f
C6876 Vbias.n315 VGND 0.19501f
C6877 Vbias.n316 VGND 0.12932f
C6878 Vbias.t105 VGND 0.17882f
C6879 Vbias.n317 VGND 0.19501f
C6880 Vbias.n318 VGND 0.12932f
C6881 Vbias.n319 VGND 0.55831f
C6882 Vbias.t121 VGND 0.17882f
C6883 Vbias.n320 VGND 0.19466f
C6884 Vbias.t195 VGND 0.17882f
C6885 Vbias.n321 VGND 0.19501f
C6886 Vbias.n322 VGND 0.12932f
C6887 Vbias.t37 VGND 0.17882f
C6888 Vbias.n323 VGND 0.19501f
C6889 Vbias.n324 VGND 0.12932f
C6890 Vbias.t48 VGND 0.17882f
C6891 Vbias.n325 VGND 0.19501f
C6892 Vbias.n326 VGND 0.12932f
C6893 Vbias.t135 VGND 0.17882f
C6894 Vbias.n327 VGND 0.19501f
C6895 Vbias.n328 VGND 0.12932f
C6896 Vbias.t221 VGND 0.17882f
C6897 Vbias.n329 VGND 0.19501f
C6898 Vbias.n330 VGND 0.12932f
C6899 Vbias.t50 VGND 0.17882f
C6900 Vbias.n331 VGND 0.19501f
C6901 Vbias.n332 VGND 0.12932f
C6902 Vbias.t138 VGND 0.17882f
C6903 Vbias.n333 VGND 0.19501f
C6904 Vbias.n334 VGND 0.12932f
C6905 Vbias.t163 VGND 0.17882f
C6906 Vbias.n335 VGND 0.19501f
C6907 Vbias.n336 VGND 0.12932f
C6908 Vbias.t236 VGND 0.17882f
C6909 Vbias.n337 VGND 0.19501f
C6910 Vbias.n338 VGND 0.12932f
C6911 Vbias.t65 VGND 0.17882f
C6912 Vbias.n339 VGND 0.19501f
C6913 Vbias.n340 VGND 0.12932f
C6914 Vbias.t90 VGND 0.17882f
C6915 Vbias.n341 VGND 0.19501f
C6916 Vbias.n342 VGND 0.12932f
C6917 Vbias.t243 VGND 0.17882f
C6918 Vbias.n343 VGND 0.19501f
C6919 Vbias.n344 VGND 0.12932f
C6920 Vbias.t7 VGND 0.17882f
C6921 Vbias.n345 VGND 0.19501f
C6922 Vbias.n346 VGND 0.12932f
C6923 Vbias.t20 VGND 0.17882f
C6924 Vbias.n347 VGND 0.19501f
C6925 Vbias.n348 VGND 0.12932f
C6926 Vbias.t176 VGND 0.17882f
C6927 Vbias.n349 VGND 0.19501f
C6928 Vbias.n350 VGND 0.12932f
C6929 Vbias.n351 VGND 0.55831f
C6930 Vbias.t198 VGND 0.17882f
C6931 Vbias.n352 VGND 0.19466f
C6932 Vbias.t17 VGND 0.17882f
C6933 Vbias.n353 VGND 0.19501f
C6934 Vbias.n354 VGND 0.12932f
C6935 Vbias.t113 VGND 0.17882f
C6936 Vbias.n355 VGND 0.19501f
C6937 Vbias.n356 VGND 0.12932f
C6938 Vbias.t124 VGND 0.17882f
C6939 Vbias.n357 VGND 0.19501f
C6940 Vbias.n358 VGND 0.12932f
C6941 Vbias.t213 VGND 0.17882f
C6942 Vbias.n359 VGND 0.19501f
C6943 Vbias.n360 VGND 0.12932f
C6944 Vbias.t40 VGND 0.17882f
C6945 Vbias.n361 VGND 0.19501f
C6946 Vbias.n362 VGND 0.12932f
C6947 Vbias.t127 VGND 0.17882f
C6948 Vbias.n363 VGND 0.19501f
C6949 Vbias.n364 VGND 0.12932f
C6950 Vbias.t219 VGND 0.17882f
C6951 Vbias.n365 VGND 0.19501f
C6952 Vbias.n366 VGND 0.12932f
C6953 Vbias.t240 VGND 0.17882f
C6954 Vbias.n367 VGND 0.19501f
C6955 Vbias.n368 VGND 0.12932f
C6956 Vbias.t54 VGND 0.17882f
C6957 Vbias.n369 VGND 0.19501f
C6958 Vbias.n370 VGND 0.12932f
C6959 Vbias.t144 VGND 0.17882f
C6960 Vbias.n371 VGND 0.19501f
C6961 Vbias.n372 VGND 0.12932f
C6962 Vbias.t166 VGND 0.17882f
C6963 Vbias.n373 VGND 0.19501f
C6964 Vbias.n374 VGND 0.12932f
C6965 Vbias.t62 VGND 0.17882f
C6966 Vbias.n375 VGND 0.19501f
C6967 Vbias.n376 VGND 0.12932f
C6968 Vbias.t81 VGND 0.17882f
C6969 Vbias.n377 VGND 0.19501f
C6970 Vbias.n378 VGND 0.12932f
C6971 Vbias.t92 VGND 0.17882f
C6972 Vbias.n379 VGND 0.19501f
C6973 Vbias.n380 VGND 0.12932f
C6974 Vbias.t255 VGND 0.17882f
C6975 Vbias.n381 VGND 0.19501f
C6976 Vbias.n382 VGND 0.12932f
C6977 Vbias.n383 VGND 0.55831f
C6978 Vbias.t16 VGND 0.17882f
C6979 Vbias.n384 VGND 0.19466f
C6980 Vbias.t88 VGND 0.17882f
C6981 Vbias.n385 VGND 0.19501f
C6982 Vbias.n386 VGND 0.12932f
C6983 Vbias.t185 VGND 0.17882f
C6984 Vbias.n387 VGND 0.19501f
C6985 Vbias.n388 VGND 0.12932f
C6986 Vbias.t196 VGND 0.17882f
C6987 Vbias.n389 VGND 0.19501f
C6988 Vbias.n390 VGND 0.12932f
C6989 Vbias.t29 VGND 0.17882f
C6990 Vbias.n391 VGND 0.19501f
C6991 Vbias.n392 VGND 0.12932f
C6992 Vbias.t112 VGND 0.17882f
C6993 Vbias.n393 VGND 0.19501f
C6994 Vbias.n394 VGND 0.12932f
C6995 Vbias.t200 VGND 0.17882f
C6996 Vbias.n395 VGND 0.19501f
C6997 Vbias.n396 VGND 0.12932f
C6998 Vbias.t33 VGND 0.17882f
C6999 Vbias.n397 VGND 0.19501f
C7000 Vbias.n398 VGND 0.12932f
C7001 Vbias.t53 VGND 0.17882f
C7002 Vbias.n399 VGND 0.19501f
C7003 Vbias.n400 VGND 0.12932f
C7004 Vbias.t126 VGND 0.17882f
C7005 Vbias.n401 VGND 0.19501f
C7006 Vbias.n402 VGND 0.12932f
C7007 Vbias.t217 VGND 0.17882f
C7008 Vbias.n403 VGND 0.19501f
C7009 Vbias.n404 VGND 0.12932f
C7010 Vbias.t239 VGND 0.17882f
C7011 Vbias.n405 VGND 0.19501f
C7012 Vbias.n406 VGND 0.12932f
C7013 Vbias.t133 VGND 0.17882f
C7014 Vbias.n407 VGND 0.19501f
C7015 Vbias.n408 VGND 0.12932f
C7016 Vbias.t153 VGND 0.17882f
C7017 Vbias.n409 VGND 0.19501f
C7018 Vbias.n410 VGND 0.12932f
C7019 Vbias.t165 VGND 0.17882f
C7020 Vbias.n411 VGND 0.19501f
C7021 Vbias.n412 VGND 0.12932f
C7022 Vbias.t73 VGND 0.17882f
C7023 Vbias.n413 VGND 0.19501f
C7024 Vbias.n414 VGND 0.12932f
C7025 Vbias.n415 VGND 0.55831f
C7026 Vbias.t87 VGND 0.17882f
C7027 Vbias.n416 VGND 0.19466f
C7028 Vbias.t160 VGND 0.17882f
C7029 Vbias.n417 VGND 0.19501f
C7030 Vbias.n418 VGND 0.12932f
C7031 Vbias.t261 VGND 0.17882f
C7032 Vbias.n419 VGND 0.19501f
C7033 Vbias.n420 VGND 0.12932f
C7034 Vbias.t14 VGND 0.17882f
C7035 Vbias.n421 VGND 0.19501f
C7036 Vbias.n422 VGND 0.12932f
C7037 Vbias.t99 VGND 0.17882f
C7038 Vbias.n423 VGND 0.19501f
C7039 Vbias.n424 VGND 0.12932f
C7040 Vbias.t183 VGND 0.17882f
C7041 Vbias.n425 VGND 0.19501f
C7042 Vbias.n426 VGND 0.12932f
C7043 Vbias.t18 VGND 0.17882f
C7044 Vbias.n427 VGND 0.19501f
C7045 Vbias.n428 VGND 0.12932f
C7046 Vbias.t102 VGND 0.17882f
C7047 Vbias.n429 VGND 0.19501f
C7048 Vbias.n430 VGND 0.12932f
C7049 Vbias.t125 VGND 0.17882f
C7050 Vbias.n431 VGND 0.19501f
C7051 Vbias.n432 VGND 0.12932f
C7052 Vbias.t199 VGND 0.17882f
C7053 Vbias.n433 VGND 0.19501f
C7054 Vbias.n434 VGND 0.12932f
C7055 Vbias.t32 VGND 0.17882f
C7056 Vbias.n435 VGND 0.19501f
C7057 Vbias.n436 VGND 0.12932f
C7058 Vbias.t52 VGND 0.17882f
C7059 Vbias.n437 VGND 0.19501f
C7060 Vbias.n438 VGND 0.12932f
C7061 Vbias.t205 VGND 0.17882f
C7062 Vbias.n439 VGND 0.19501f
C7063 Vbias.n440 VGND 0.12932f
C7064 Vbias.t225 VGND 0.17882f
C7065 Vbias.n441 VGND 0.19501f
C7066 Vbias.n442 VGND 0.12932f
C7067 Vbias.t238 VGND 0.17882f
C7068 Vbias.n443 VGND 0.19501f
C7069 Vbias.n444 VGND 0.12932f
C7070 Vbias.t146 VGND 0.17882f
C7071 Vbias.n445 VGND 0.19501f
C7072 Vbias.n446 VGND 0.12932f
C7073 Vbias.n447 VGND 0.55831f
C7074 Vbias.t57 VGND 0.17882f
C7075 Vbias.n448 VGND 0.19466f
C7076 Vbias.t130 VGND 0.17882f
C7077 Vbias.n449 VGND 0.19501f
C7078 Vbias.n450 VGND 0.12932f
C7079 Vbias.t229 VGND 0.17882f
C7080 Vbias.n451 VGND 0.19501f
C7081 Vbias.n452 VGND 0.12932f
C7082 Vbias.t242 VGND 0.17882f
C7083 Vbias.n453 VGND 0.19501f
C7084 Vbias.n454 VGND 0.12932f
C7085 Vbias.t69 VGND 0.17882f
C7086 Vbias.n455 VGND 0.19501f
C7087 Vbias.n456 VGND 0.12932f
C7088 Vbias.t156 VGND 0.17882f
C7089 Vbias.n457 VGND 0.19501f
C7090 Vbias.n458 VGND 0.12932f
C7091 Vbias.t247 VGND 0.17882f
C7092 Vbias.n459 VGND 0.19501f
C7093 Vbias.n460 VGND 0.12932f
C7094 Vbias.t76 VGND 0.17882f
C7095 Vbias.n461 VGND 0.19501f
C7096 Vbias.n462 VGND 0.12932f
C7097 Vbias.t96 VGND 0.17882f
C7098 Vbias.n463 VGND 0.19501f
C7099 Vbias.n464 VGND 0.12932f
C7100 Vbias.t171 VGND 0.17882f
C7101 Vbias.n465 VGND 0.19501f
C7102 Vbias.n466 VGND 0.12932f
C7103 Vbias.t258 VGND 0.17882f
C7104 Vbias.n467 VGND 0.19501f
C7105 Vbias.n468 VGND 0.12932f
C7106 Vbias.t25 VGND 0.17882f
C7107 Vbias.n469 VGND 0.19501f
C7108 Vbias.n470 VGND 0.12932f
C7109 Vbias.t173 VGND 0.17882f
C7110 Vbias.n471 VGND 0.19501f
C7111 Vbias.n472 VGND 0.12932f
C7112 Vbias.t193 VGND 0.17882f
C7113 Vbias.n473 VGND 0.19501f
C7114 Vbias.n474 VGND 0.12932f
C7115 Vbias.t210 VGND 0.17882f
C7116 Vbias.n475 VGND 0.19501f
C7117 Vbias.n476 VGND 0.12932f
C7118 Vbias.t110 VGND 0.17882f
C7119 Vbias.n477 VGND 0.19501f
C7120 Vbias.n478 VGND 0.12932f
C7121 Vbias.n479 VGND 0.55831f
C7122 Vbias.t129 VGND 0.17882f
C7123 Vbias.n480 VGND 0.19466f
C7124 Vbias.t201 VGND 0.17882f
C7125 Vbias.n481 VGND 0.19501f
C7126 Vbias.n482 VGND 0.12932f
C7127 Vbias.t41 VGND 0.17882f
C7128 Vbias.n483 VGND 0.19501f
C7129 Vbias.n484 VGND 0.12932f
C7130 Vbias.t56 VGND 0.17882f
C7131 Vbias.n485 VGND 0.19501f
C7132 Vbias.n486 VGND 0.12932f
C7133 Vbias.t141 VGND 0.17882f
C7134 Vbias.n487 VGND 0.19501f
C7135 Vbias.n488 VGND 0.12932f
C7136 Vbias.t227 VGND 0.17882f
C7137 Vbias.n489 VGND 0.19501f
C7138 Vbias.n490 VGND 0.12932f
C7139 Vbias.t60 VGND 0.17882f
C7140 Vbias.n491 VGND 0.19501f
C7141 Vbias.n492 VGND 0.12932f
C7142 Vbias.t147 VGND 0.17882f
C7143 Vbias.n493 VGND 0.19501f
C7144 Vbias.n494 VGND 0.12932f
C7145 Vbias.t169 VGND 0.17882f
C7146 Vbias.n495 VGND 0.19501f
C7147 Vbias.n496 VGND 0.12932f
C7148 Vbias.t246 VGND 0.17882f
C7149 Vbias.n497 VGND 0.19501f
C7150 Vbias.n498 VGND 0.12932f
C7151 Vbias.t75 VGND 0.17882f
C7152 Vbias.n499 VGND 0.19501f
C7153 Vbias.n500 VGND 0.12932f
C7154 Vbias.t95 VGND 0.17882f
C7155 Vbias.n501 VGND 0.19501f
C7156 Vbias.n502 VGND 0.12932f
C7157 Vbias.t248 VGND 0.17882f
C7158 Vbias.n503 VGND 0.19501f
C7159 Vbias.n504 VGND 0.12932f
C7160 Vbias.t12 VGND 0.17882f
C7161 Vbias.n505 VGND 0.19501f
C7162 Vbias.n506 VGND 0.12932f
C7163 Vbias.t24 VGND 0.17882f
C7164 Vbias.n507 VGND 0.19501f
C7165 Vbias.n508 VGND 0.12932f
C7166 Vbias.t181 VGND 0.17882f
C7167 Vbias.n509 VGND 0.19501f
C7168 Vbias.n510 VGND 0.12932f
C7169 Vbias.n511 VGND 0.64934f
C7170 Vbias.t3 VGND 0.03654f
C7171 Vbias.t4 VGND 0.03654f
C7172 Vbias.n512 VGND 0.24617f
C7173 Vbias.t5 VGND 0.03654f
C7174 Vbias.t0 VGND 0.03654f
C7175 Vbias.n513 VGND 0.24617f
C7176 Vbias.n514 VGND 0.74304f
C7177 Vbias.t2 VGND 0.17043f
C7178 Vbias.t1 VGND 0.67015f
C7179 Vbias.n515 VGND 1.2407f
C7180 Vbias.n516 VGND 0.47721f
C7181 Vbias.n517 VGND 1.11739f
C7182 XThC.Tn[2].t4 VGND 0.01169f
C7183 XThC.Tn[2].t3 VGND 0.01169f
C7184 XThC.Tn[2].n0 VGND 0.02361f
C7185 XThC.Tn[2].t2 VGND 0.01169f
C7186 XThC.Tn[2].t1 VGND 0.01169f
C7187 XThC.Tn[2].n1 VGND 0.02762f
C7188 XThC.Tn[2].n2 VGND 0.07732f
C7189 XThC.Tn[2].n3 VGND 0.01731f
C7190 XThC.Tn[2].n4 VGND 0.01731f
C7191 XThC.Tn[2].n5 VGND 0.02884f
C7192 XThC.Tn[2].n6 VGND 0.01731f
C7193 XThC.Tn[2].n7 VGND 0.08243f
C7194 XThC.Tn[2].n8 VGND 0.05096f
C7195 XThC.Tn[2].n9 VGND 0.05751f
C7196 XThC.Tn[2].t18 VGND 0.01012f
C7197 XThC.Tn[2].n10 VGND 0.02261f
C7198 XThC.Tn[2].n11 VGND 0.01292f
C7199 XThC.Tn[2].n12 VGND 0.01571f
C7200 XThC.Tn[2].t35 VGND 0.01012f
C7201 XThC.Tn[2].n13 VGND 0.02261f
C7202 XThC.Tn[2].n14 VGND 0.01292f
C7203 XThC.Tn[2].n15 VGND 0.07465f
C7204 XThC.Tn[2].t37 VGND 0.01012f
C7205 XThC.Tn[2].n16 VGND 0.02261f
C7206 XThC.Tn[2].n17 VGND 0.01292f
C7207 XThC.Tn[2].n18 VGND 0.07465f
C7208 XThC.Tn[2].t39 VGND 0.01012f
C7209 XThC.Tn[2].n19 VGND 0.02261f
C7210 XThC.Tn[2].n20 VGND 0.01292f
C7211 XThC.Tn[2].n21 VGND 0.07465f
C7212 XThC.Tn[2].t28 VGND 0.01012f
C7213 XThC.Tn[2].n22 VGND 0.02261f
C7214 XThC.Tn[2].n23 VGND 0.01292f
C7215 XThC.Tn[2].n24 VGND 0.07465f
C7216 XThC.Tn[2].t29 VGND 0.01012f
C7217 XThC.Tn[2].n25 VGND 0.02261f
C7218 XThC.Tn[2].n26 VGND 0.01292f
C7219 XThC.Tn[2].n27 VGND 0.07465f
C7220 XThC.Tn[2].t42 VGND 0.01012f
C7221 XThC.Tn[2].n28 VGND 0.02261f
C7222 XThC.Tn[2].n29 VGND 0.01292f
C7223 XThC.Tn[2].n30 VGND 0.07465f
C7224 XThC.Tn[2].t19 VGND 0.01012f
C7225 XThC.Tn[2].n31 VGND 0.02261f
C7226 XThC.Tn[2].n32 VGND 0.01292f
C7227 XThC.Tn[2].n33 VGND 0.07465f
C7228 XThC.Tn[2].t21 VGND 0.01012f
C7229 XThC.Tn[2].n34 VGND 0.02261f
C7230 XThC.Tn[2].n35 VGND 0.01292f
C7231 XThC.Tn[2].n36 VGND 0.07465f
C7232 XThC.Tn[2].t40 VGND 0.01012f
C7233 XThC.Tn[2].n37 VGND 0.02261f
C7234 XThC.Tn[2].n38 VGND 0.01292f
C7235 XThC.Tn[2].n39 VGND 0.07465f
C7236 XThC.Tn[2].t41 VGND 0.01012f
C7237 XThC.Tn[2].n40 VGND 0.02261f
C7238 XThC.Tn[2].n41 VGND 0.01292f
C7239 XThC.Tn[2].n42 VGND 0.07465f
C7240 XThC.Tn[2].t22 VGND 0.01012f
C7241 XThC.Tn[2].n43 VGND 0.02261f
C7242 XThC.Tn[2].n44 VGND 0.01292f
C7243 XThC.Tn[2].n45 VGND 0.07465f
C7244 XThC.Tn[2].t30 VGND 0.01012f
C7245 XThC.Tn[2].n46 VGND 0.02261f
C7246 XThC.Tn[2].n47 VGND 0.01292f
C7247 XThC.Tn[2].n48 VGND 0.07465f
C7248 XThC.Tn[2].t33 VGND 0.01012f
C7249 XThC.Tn[2].n49 VGND 0.02261f
C7250 XThC.Tn[2].n50 VGND 0.01292f
C7251 XThC.Tn[2].n51 VGND 0.07465f
C7252 XThC.Tn[2].t14 VGND 0.01012f
C7253 XThC.Tn[2].n52 VGND 0.02261f
C7254 XThC.Tn[2].n53 VGND 0.01292f
C7255 XThC.Tn[2].n54 VGND 0.07465f
C7256 XThC.Tn[2].t24 VGND 0.01012f
C7257 XThC.Tn[2].n55 VGND 0.02261f
C7258 XThC.Tn[2].n56 VGND 0.01292f
C7259 XThC.Tn[2].n57 VGND 0.07465f
C7260 XThC.Tn[2].n58 VGND 0.27153f
C7261 XThC.Tn[2].n59 VGND 0.0441f
C7262 XThC.Tn[2].n60 VGND 0.02447f
C7263 XThC.Tn[4].t5 VGND 0.01194f
C7264 XThC.Tn[4].t4 VGND 0.01194f
C7265 XThC.Tn[4].n0 VGND 0.02411f
C7266 XThC.Tn[4].t7 VGND 0.01194f
C7267 XThC.Tn[4].t6 VGND 0.01194f
C7268 XThC.Tn[4].n1 VGND 0.02821f
C7269 XThC.Tn[4].n2 VGND 0.07897f
C7270 XThC.Tn[4].n3 VGND 0.01768f
C7271 XThC.Tn[4].n4 VGND 0.01768f
C7272 XThC.Tn[4].n5 VGND 0.01768f
C7273 XThC.Tn[4].n6 VGND 0.02946f
C7274 XThC.Tn[4].n7 VGND 0.0842f
C7275 XThC.Tn[4].n8 VGND 0.05205f
C7276 XThC.Tn[4].n9 VGND 0.05874f
C7277 XThC.Tn[4].t26 VGND 0.01034f
C7278 XThC.Tn[4].n10 VGND 0.02309f
C7279 XThC.Tn[4].n11 VGND 0.0132f
C7280 XThC.Tn[4].n12 VGND 0.01605f
C7281 XThC.Tn[4].t43 VGND 0.01034f
C7282 XThC.Tn[4].n13 VGND 0.02309f
C7283 XThC.Tn[4].n14 VGND 0.0132f
C7284 XThC.Tn[4].n15 VGND 0.07625f
C7285 XThC.Tn[4].t13 VGND 0.01034f
C7286 XThC.Tn[4].n16 VGND 0.02309f
C7287 XThC.Tn[4].n17 VGND 0.0132f
C7288 XThC.Tn[4].n18 VGND 0.07625f
C7289 XThC.Tn[4].t15 VGND 0.01034f
C7290 XThC.Tn[4].n19 VGND 0.02309f
C7291 XThC.Tn[4].n20 VGND 0.0132f
C7292 XThC.Tn[4].n21 VGND 0.07625f
C7293 XThC.Tn[4].t36 VGND 0.01034f
C7294 XThC.Tn[4].n22 VGND 0.02309f
C7295 XThC.Tn[4].n23 VGND 0.0132f
C7296 XThC.Tn[4].n24 VGND 0.07625f
C7297 XThC.Tn[4].t37 VGND 0.01034f
C7298 XThC.Tn[4].n25 VGND 0.02309f
C7299 XThC.Tn[4].n26 VGND 0.0132f
C7300 XThC.Tn[4].n27 VGND 0.07625f
C7301 XThC.Tn[4].t18 VGND 0.01034f
C7302 XThC.Tn[4].n28 VGND 0.02309f
C7303 XThC.Tn[4].n29 VGND 0.0132f
C7304 XThC.Tn[4].n30 VGND 0.07625f
C7305 XThC.Tn[4].t27 VGND 0.01034f
C7306 XThC.Tn[4].n31 VGND 0.02309f
C7307 XThC.Tn[4].n32 VGND 0.0132f
C7308 XThC.Tn[4].n33 VGND 0.07625f
C7309 XThC.Tn[4].t29 VGND 0.01034f
C7310 XThC.Tn[4].n34 VGND 0.02309f
C7311 XThC.Tn[4].n35 VGND 0.0132f
C7312 XThC.Tn[4].n36 VGND 0.07625f
C7313 XThC.Tn[4].t16 VGND 0.01034f
C7314 XThC.Tn[4].n37 VGND 0.02309f
C7315 XThC.Tn[4].n38 VGND 0.0132f
C7316 XThC.Tn[4].n39 VGND 0.07625f
C7317 XThC.Tn[4].t17 VGND 0.01034f
C7318 XThC.Tn[4].n40 VGND 0.02309f
C7319 XThC.Tn[4].n41 VGND 0.0132f
C7320 XThC.Tn[4].n42 VGND 0.07625f
C7321 XThC.Tn[4].t30 VGND 0.01034f
C7322 XThC.Tn[4].n43 VGND 0.02309f
C7323 XThC.Tn[4].n44 VGND 0.0132f
C7324 XThC.Tn[4].n45 VGND 0.07625f
C7325 XThC.Tn[4].t38 VGND 0.01034f
C7326 XThC.Tn[4].n46 VGND 0.02309f
C7327 XThC.Tn[4].n47 VGND 0.0132f
C7328 XThC.Tn[4].n48 VGND 0.07625f
C7329 XThC.Tn[4].t41 VGND 0.01034f
C7330 XThC.Tn[4].n49 VGND 0.02309f
C7331 XThC.Tn[4].n50 VGND 0.0132f
C7332 XThC.Tn[4].n51 VGND 0.07625f
C7333 XThC.Tn[4].t22 VGND 0.01034f
C7334 XThC.Tn[4].n52 VGND 0.02309f
C7335 XThC.Tn[4].n53 VGND 0.0132f
C7336 XThC.Tn[4].n54 VGND 0.07625f
C7337 XThC.Tn[4].t32 VGND 0.01034f
C7338 XThC.Tn[4].n55 VGND 0.02309f
C7339 XThC.Tn[4].n56 VGND 0.0132f
C7340 XThC.Tn[4].n57 VGND 0.07625f
C7341 XThC.Tn[4].n58 VGND 0.23757f
C7342 XThC.Tn[4].n59 VGND 0.04514f
C7343 XThC.Tn[4].n60 VGND 0.025f
C7344 XThR.Tn[5].t10 VGND 0.01808f
C7345 XThR.Tn[5].t11 VGND 0.01808f
C7346 XThR.Tn[5].n0 VGND 0.03649f
C7347 XThR.Tn[5].t9 VGND 0.01808f
C7348 XThR.Tn[5].t8 VGND 0.01808f
C7349 XThR.Tn[5].n1 VGND 0.04269f
C7350 XThR.Tn[5].n2 VGND 0.11952f
C7351 XThR.Tn[5].t7 VGND 0.01175f
C7352 XThR.Tn[5].t4 VGND 0.01175f
C7353 XThR.Tn[5].n3 VGND 0.02676f
C7354 XThR.Tn[5].t6 VGND 0.01175f
C7355 XThR.Tn[5].t5 VGND 0.01175f
C7356 XThR.Tn[5].n4 VGND 0.02676f
C7357 XThR.Tn[5].t0 VGND 0.01175f
C7358 XThR.Tn[5].t1 VGND 0.01175f
C7359 XThR.Tn[5].n5 VGND 0.04459f
C7360 XThR.Tn[5].t3 VGND 0.01175f
C7361 XThR.Tn[5].t2 VGND 0.01175f
C7362 XThR.Tn[5].n6 VGND 0.02676f
C7363 XThR.Tn[5].n7 VGND 0.12743f
C7364 XThR.Tn[5].n8 VGND 0.07877f
C7365 XThR.Tn[5].n9 VGND 0.0889f
C7366 XThR.Tn[5].t17 VGND 0.01413f
C7367 XThR.Tn[5].t72 VGND 0.01547f
C7368 XThR.Tn[5].n10 VGND 0.03778f
C7369 XThR.Tn[5].n11 VGND 0.07257f
C7370 XThR.Tn[5].t39 VGND 0.01413f
C7371 XThR.Tn[5].t26 VGND 0.01547f
C7372 XThR.Tn[5].n12 VGND 0.03778f
C7373 XThR.Tn[5].t13 VGND 0.01408f
C7374 XThR.Tn[5].t23 VGND 0.01542f
C7375 XThR.Tn[5].n13 VGND 0.03931f
C7376 XThR.Tn[5].n14 VGND 0.02761f
C7377 XThR.Tn[5].n16 VGND 0.08862f
C7378 XThR.Tn[5].t73 VGND 0.01413f
C7379 XThR.Tn[5].t66 VGND 0.01547f
C7380 XThR.Tn[5].n17 VGND 0.03778f
C7381 XThR.Tn[5].t48 VGND 0.01408f
C7382 XThR.Tn[5].t61 VGND 0.01542f
C7383 XThR.Tn[5].n18 VGND 0.03931f
C7384 XThR.Tn[5].n19 VGND 0.02761f
C7385 XThR.Tn[5].n21 VGND 0.08862f
C7386 XThR.Tn[5].t28 VGND 0.01413f
C7387 XThR.Tn[5].t21 VGND 0.01547f
C7388 XThR.Tn[5].n22 VGND 0.03778f
C7389 XThR.Tn[5].t65 VGND 0.01408f
C7390 XThR.Tn[5].t18 VGND 0.01542f
C7391 XThR.Tn[5].n23 VGND 0.03931f
C7392 XThR.Tn[5].n24 VGND 0.02761f
C7393 XThR.Tn[5].n26 VGND 0.08862f
C7394 XThR.Tn[5].t55 VGND 0.01413f
C7395 XThR.Tn[5].t51 VGND 0.01547f
C7396 XThR.Tn[5].n27 VGND 0.03778f
C7397 XThR.Tn[5].t33 VGND 0.01408f
C7398 XThR.Tn[5].t46 VGND 0.01542f
C7399 XThR.Tn[5].n28 VGND 0.03931f
C7400 XThR.Tn[5].n29 VGND 0.02761f
C7401 XThR.Tn[5].n31 VGND 0.08862f
C7402 XThR.Tn[5].t30 VGND 0.01413f
C7403 XThR.Tn[5].t22 VGND 0.01547f
C7404 XThR.Tn[5].n32 VGND 0.03778f
C7405 XThR.Tn[5].t67 VGND 0.01408f
C7406 XThR.Tn[5].t19 VGND 0.01542f
C7407 XThR.Tn[5].n33 VGND 0.03931f
C7408 XThR.Tn[5].n34 VGND 0.02761f
C7409 XThR.Tn[5].n36 VGND 0.08862f
C7410 XThR.Tn[5].t69 VGND 0.01413f
C7411 XThR.Tn[5].t40 VGND 0.01547f
C7412 XThR.Tn[5].n37 VGND 0.03778f
C7413 XThR.Tn[5].t43 VGND 0.01408f
C7414 XThR.Tn[5].t37 VGND 0.01542f
C7415 XThR.Tn[5].n38 VGND 0.03931f
C7416 XThR.Tn[5].n39 VGND 0.02761f
C7417 XThR.Tn[5].n41 VGND 0.08862f
C7418 XThR.Tn[5].t38 VGND 0.01413f
C7419 XThR.Tn[5].t32 VGND 0.01547f
C7420 XThR.Tn[5].n42 VGND 0.03778f
C7421 XThR.Tn[5].t14 VGND 0.01408f
C7422 XThR.Tn[5].t29 VGND 0.01542f
C7423 XThR.Tn[5].n43 VGND 0.03931f
C7424 XThR.Tn[5].n44 VGND 0.02761f
C7425 XThR.Tn[5].n46 VGND 0.08862f
C7426 XThR.Tn[5].t42 VGND 0.01413f
C7427 XThR.Tn[5].t49 VGND 0.01547f
C7428 XThR.Tn[5].n47 VGND 0.03778f
C7429 XThR.Tn[5].t16 VGND 0.01408f
C7430 XThR.Tn[5].t45 VGND 0.01542f
C7431 XThR.Tn[5].n48 VGND 0.03931f
C7432 XThR.Tn[5].n49 VGND 0.02761f
C7433 XThR.Tn[5].n51 VGND 0.08862f
C7434 XThR.Tn[5].t58 VGND 0.01413f
C7435 XThR.Tn[5].t68 VGND 0.01547f
C7436 XThR.Tn[5].n52 VGND 0.03778f
C7437 XThR.Tn[5].t36 VGND 0.01408f
C7438 XThR.Tn[5].t63 VGND 0.01542f
C7439 XThR.Tn[5].n53 VGND 0.03931f
C7440 XThR.Tn[5].n54 VGND 0.02761f
C7441 XThR.Tn[5].n56 VGND 0.08862f
C7442 XThR.Tn[5].t53 VGND 0.01413f
C7443 XThR.Tn[5].t24 VGND 0.01547f
C7444 XThR.Tn[5].n57 VGND 0.03778f
C7445 XThR.Tn[5].t25 VGND 0.01408f
C7446 XThR.Tn[5].t20 VGND 0.01542f
C7447 XThR.Tn[5].n58 VGND 0.03931f
C7448 XThR.Tn[5].n59 VGND 0.02761f
C7449 XThR.Tn[5].n61 VGND 0.08862f
C7450 XThR.Tn[5].t71 VGND 0.01413f
C7451 XThR.Tn[5].t60 VGND 0.01547f
C7452 XThR.Tn[5].n62 VGND 0.03778f
C7453 XThR.Tn[5].t44 VGND 0.01408f
C7454 XThR.Tn[5].t57 VGND 0.01542f
C7455 XThR.Tn[5].n63 VGND 0.03931f
C7456 XThR.Tn[5].n64 VGND 0.02761f
C7457 XThR.Tn[5].n66 VGND 0.08862f
C7458 XThR.Tn[5].t41 VGND 0.01413f
C7459 XThR.Tn[5].t35 VGND 0.01547f
C7460 XThR.Tn[5].n67 VGND 0.03778f
C7461 XThR.Tn[5].t15 VGND 0.01408f
C7462 XThR.Tn[5].t31 VGND 0.01542f
C7463 XThR.Tn[5].n68 VGND 0.03931f
C7464 XThR.Tn[5].n69 VGND 0.02761f
C7465 XThR.Tn[5].n71 VGND 0.08862f
C7466 XThR.Tn[5].t56 VGND 0.01413f
C7467 XThR.Tn[5].t52 VGND 0.01547f
C7468 XThR.Tn[5].n72 VGND 0.03778f
C7469 XThR.Tn[5].t34 VGND 0.01408f
C7470 XThR.Tn[5].t47 VGND 0.01542f
C7471 XThR.Tn[5].n73 VGND 0.03931f
C7472 XThR.Tn[5].n74 VGND 0.02761f
C7473 XThR.Tn[5].n76 VGND 0.08862f
C7474 XThR.Tn[5].t12 VGND 0.01413f
C7475 XThR.Tn[5].t70 VGND 0.01547f
C7476 XThR.Tn[5].n77 VGND 0.03778f
C7477 XThR.Tn[5].t50 VGND 0.01408f
C7478 XThR.Tn[5].t64 VGND 0.01542f
C7479 XThR.Tn[5].n78 VGND 0.03931f
C7480 XThR.Tn[5].n79 VGND 0.02761f
C7481 XThR.Tn[5].n81 VGND 0.08862f
C7482 XThR.Tn[5].t54 VGND 0.01413f
C7483 XThR.Tn[5].t62 VGND 0.01547f
C7484 XThR.Tn[5].n82 VGND 0.03778f
C7485 XThR.Tn[5].t27 VGND 0.01408f
C7486 XThR.Tn[5].t59 VGND 0.01542f
C7487 XThR.Tn[5].n83 VGND 0.03931f
C7488 XThR.Tn[5].n84 VGND 0.02761f
C7489 XThR.Tn[5].n86 VGND 0.08862f
C7490 XThR.Tn[5].n87 VGND 0.08053f
C7491 XThR.Tn[5].n88 VGND 0.15597f
C7492 XThR.Tn[5].n89 VGND 0.03783f
C7493 XThR.Tn[3].t5 VGND 0.01821f
C7494 XThR.Tn[3].t6 VGND 0.01821f
C7495 XThR.Tn[3].n0 VGND 0.03675f
C7496 XThR.Tn[3].t4 VGND 0.01821f
C7497 XThR.Tn[3].t7 VGND 0.01821f
C7498 XThR.Tn[3].n1 VGND 0.043f
C7499 XThR.Tn[3].n2 VGND 0.12037f
C7500 XThR.Tn[3].t11 VGND 0.01183f
C7501 XThR.Tn[3].t8 VGND 0.01183f
C7502 XThR.Tn[3].n3 VGND 0.02695f
C7503 XThR.Tn[3].t10 VGND 0.01183f
C7504 XThR.Tn[3].t9 VGND 0.01183f
C7505 XThR.Tn[3].n4 VGND 0.02695f
C7506 XThR.Tn[3].t0 VGND 0.01183f
C7507 XThR.Tn[3].t1 VGND 0.01183f
C7508 XThR.Tn[3].n5 VGND 0.0449f
C7509 XThR.Tn[3].t3 VGND 0.01183f
C7510 XThR.Tn[3].t2 VGND 0.01183f
C7511 XThR.Tn[3].n6 VGND 0.02695f
C7512 XThR.Tn[3].n7 VGND 0.12834f
C7513 XThR.Tn[3].n8 VGND 0.07933f
C7514 XThR.Tn[3].n9 VGND 0.08953f
C7515 XThR.Tn[3].t64 VGND 0.01423f
C7516 XThR.Tn[3].t57 VGND 0.01558f
C7517 XThR.Tn[3].n10 VGND 0.03805f
C7518 XThR.Tn[3].n11 VGND 0.07309f
C7519 XThR.Tn[3].t18 VGND 0.01423f
C7520 XThR.Tn[3].t70 VGND 0.01558f
C7521 XThR.Tn[3].n12 VGND 0.03805f
C7522 XThR.Tn[3].t24 VGND 0.01418f
C7523 XThR.Tn[3].t55 VGND 0.01553f
C7524 XThR.Tn[3].n13 VGND 0.03959f
C7525 XThR.Tn[3].n14 VGND 0.02781f
C7526 XThR.Tn[3].n16 VGND 0.08925f
C7527 XThR.Tn[3].t59 VGND 0.01423f
C7528 XThR.Tn[3].t49 VGND 0.01558f
C7529 XThR.Tn[3].n17 VGND 0.03805f
C7530 XThR.Tn[3].t62 VGND 0.01418f
C7531 XThR.Tn[3].t29 VGND 0.01553f
C7532 XThR.Tn[3].n18 VGND 0.03959f
C7533 XThR.Tn[3].n19 VGND 0.02781f
C7534 XThR.Tn[3].n21 VGND 0.08925f
C7535 XThR.Tn[3].t71 VGND 0.01423f
C7536 XThR.Tn[3].t67 VGND 0.01558f
C7537 XThR.Tn[3].n22 VGND 0.03805f
C7538 XThR.Tn[3].t12 VGND 0.01418f
C7539 XThR.Tn[3].t47 VGND 0.01553f
C7540 XThR.Tn[3].n23 VGND 0.03959f
C7541 XThR.Tn[3].n24 VGND 0.02781f
C7542 XThR.Tn[3].n26 VGND 0.08925f
C7543 XThR.Tn[3].t39 VGND 0.01423f
C7544 XThR.Tn[3].t33 VGND 0.01558f
C7545 XThR.Tn[3].n27 VGND 0.03805f
C7546 XThR.Tn[3].t42 VGND 0.01418f
C7547 XThR.Tn[3].t13 VGND 0.01553f
C7548 XThR.Tn[3].n28 VGND 0.03959f
C7549 XThR.Tn[3].n29 VGND 0.02781f
C7550 XThR.Tn[3].n31 VGND 0.08925f
C7551 XThR.Tn[3].t72 VGND 0.01423f
C7552 XThR.Tn[3].t68 VGND 0.01558f
C7553 XThR.Tn[3].n32 VGND 0.03805f
C7554 XThR.Tn[3].t16 VGND 0.01418f
C7555 XThR.Tn[3].t48 VGND 0.01553f
C7556 XThR.Tn[3].n33 VGND 0.03959f
C7557 XThR.Tn[3].n34 VGND 0.02781f
C7558 XThR.Tn[3].n36 VGND 0.08925f
C7559 XThR.Tn[3].t52 VGND 0.01423f
C7560 XThR.Tn[3].t20 VGND 0.01558f
C7561 XThR.Tn[3].n37 VGND 0.03805f
C7562 XThR.Tn[3].t56 VGND 0.01418f
C7563 XThR.Tn[3].t66 VGND 0.01553f
C7564 XThR.Tn[3].n38 VGND 0.03959f
C7565 XThR.Tn[3].n39 VGND 0.02781f
C7566 XThR.Tn[3].n41 VGND 0.08925f
C7567 XThR.Tn[3].t19 VGND 0.01423f
C7568 XThR.Tn[3].t14 VGND 0.01558f
C7569 XThR.Tn[3].n42 VGND 0.03805f
C7570 XThR.Tn[3].t23 VGND 0.01418f
C7571 XThR.Tn[3].t61 VGND 0.01553f
C7572 XThR.Tn[3].n43 VGND 0.03959f
C7573 XThR.Tn[3].n44 VGND 0.02781f
C7574 XThR.Tn[3].n46 VGND 0.08925f
C7575 XThR.Tn[3].t22 VGND 0.01423f
C7576 XThR.Tn[3].t31 VGND 0.01558f
C7577 XThR.Tn[3].n47 VGND 0.03805f
C7578 XThR.Tn[3].t28 VGND 0.01418f
C7579 XThR.Tn[3].t73 VGND 0.01553f
C7580 XThR.Tn[3].n48 VGND 0.03959f
C7581 XThR.Tn[3].n49 VGND 0.02781f
C7582 XThR.Tn[3].n51 VGND 0.08925f
C7583 XThR.Tn[3].t41 VGND 0.01423f
C7584 XThR.Tn[3].t51 VGND 0.01558f
C7585 XThR.Tn[3].n52 VGND 0.03805f
C7586 XThR.Tn[3].t45 VGND 0.01418f
C7587 XThR.Tn[3].t30 VGND 0.01553f
C7588 XThR.Tn[3].n53 VGND 0.03959f
C7589 XThR.Tn[3].n54 VGND 0.02781f
C7590 XThR.Tn[3].n56 VGND 0.08925f
C7591 XThR.Tn[3].t35 VGND 0.01423f
C7592 XThR.Tn[3].t69 VGND 0.01558f
C7593 XThR.Tn[3].n57 VGND 0.03805f
C7594 XThR.Tn[3].t37 VGND 0.01418f
C7595 XThR.Tn[3].t50 VGND 0.01553f
C7596 XThR.Tn[3].n58 VGND 0.03959f
C7597 XThR.Tn[3].n59 VGND 0.02781f
C7598 XThR.Tn[3].n61 VGND 0.08925f
C7599 XThR.Tn[3].t54 VGND 0.01423f
C7600 XThR.Tn[3].t44 VGND 0.01558f
C7601 XThR.Tn[3].n62 VGND 0.03805f
C7602 XThR.Tn[3].t58 VGND 0.01418f
C7603 XThR.Tn[3].t25 VGND 0.01553f
C7604 XThR.Tn[3].n63 VGND 0.03959f
C7605 XThR.Tn[3].n64 VGND 0.02781f
C7606 XThR.Tn[3].n66 VGND 0.08925f
C7607 XThR.Tn[3].t21 VGND 0.01423f
C7608 XThR.Tn[3].t17 VGND 0.01558f
C7609 XThR.Tn[3].n67 VGND 0.03805f
C7610 XThR.Tn[3].t26 VGND 0.01418f
C7611 XThR.Tn[3].t63 VGND 0.01553f
C7612 XThR.Tn[3].n68 VGND 0.03959f
C7613 XThR.Tn[3].n69 VGND 0.02781f
C7614 XThR.Tn[3].n71 VGND 0.08925f
C7615 XThR.Tn[3].t40 VGND 0.01423f
C7616 XThR.Tn[3].t34 VGND 0.01558f
C7617 XThR.Tn[3].n72 VGND 0.03805f
C7618 XThR.Tn[3].t43 VGND 0.01418f
C7619 XThR.Tn[3].t15 VGND 0.01553f
C7620 XThR.Tn[3].n73 VGND 0.03959f
C7621 XThR.Tn[3].n74 VGND 0.02781f
C7622 XThR.Tn[3].n76 VGND 0.08925f
C7623 XThR.Tn[3].t60 VGND 0.01423f
C7624 XThR.Tn[3].t53 VGND 0.01558f
C7625 XThR.Tn[3].n77 VGND 0.03805f
C7626 XThR.Tn[3].t65 VGND 0.01418f
C7627 XThR.Tn[3].t32 VGND 0.01553f
C7628 XThR.Tn[3].n78 VGND 0.03959f
C7629 XThR.Tn[3].n79 VGND 0.02781f
C7630 XThR.Tn[3].n81 VGND 0.08925f
C7631 XThR.Tn[3].t36 VGND 0.01423f
C7632 XThR.Tn[3].t46 VGND 0.01558f
C7633 XThR.Tn[3].n82 VGND 0.03805f
C7634 XThR.Tn[3].t38 VGND 0.01418f
C7635 XThR.Tn[3].t27 VGND 0.01553f
C7636 XThR.Tn[3].n83 VGND 0.03959f
C7637 XThR.Tn[3].n84 VGND 0.02781f
C7638 XThR.Tn[3].n86 VGND 0.08925f
C7639 XThR.Tn[3].n87 VGND 0.0811f
C7640 XThR.Tn[3].n88 VGND 0.17963f
C7641 XThR.Tn[3].n89 VGND 0.0381f
C7642 XThC.XTB4.Y.t1 VGND 0.12238f
C7643 XThC.XTB4.Y.n0 VGND 0.16166f
C7644 XThC.XTB4.Y.t4 VGND 0.02956f
C7645 XThC.XTB4.Y.t13 VGND 0.05016f
C7646 XThC.XTB4.Y.n1 VGND 0.05972f
C7647 XThC.XTB4.Y.t7 VGND 0.02956f
C7648 XThC.XTB4.Y.t17 VGND 0.05016f
C7649 XThC.XTB4.Y.n2 VGND 0.03074f
C7650 XThC.XTB4.Y.t10 VGND 0.02956f
C7651 XThC.XTB4.Y.t2 VGND 0.05016f
C7652 XThC.XTB4.Y.n3 VGND 0.06603f
C7653 XThC.XTB4.Y.t14 VGND 0.02956f
C7654 XThC.XTB4.Y.t3 VGND 0.05016f
C7655 XThC.XTB4.Y.n4 VGND 0.0613f
C7656 XThC.XTB4.Y.n5 VGND 0.03729f
C7657 XThC.XTB4.Y.n6 VGND 0.06174f
C7658 XThC.XTB4.Y.n7 VGND 0.02389f
C7659 XThC.XTB4.Y.n8 VGND 0.02916f
C7660 XThC.XTB4.Y.n9 VGND 0.06603f
C7661 XThC.XTB4.Y.n10 VGND 0.0331f
C7662 XThC.XTB4.Y.n11 VGND 0.06459f
C7663 XThC.XTB4.Y.t5 VGND 0.02956f
C7664 XThC.XTB4.Y.t16 VGND 0.05016f
C7665 XThC.XTB4.Y.n12 VGND 0.06761f
C7666 XThC.XTB4.Y.t9 VGND 0.02956f
C7667 XThC.XTB4.Y.t6 VGND 0.05016f
C7668 XThC.XTB4.Y.t15 VGND 0.02956f
C7669 XThC.XTB4.Y.t12 VGND 0.05016f
C7670 XThC.XTB4.Y.t11 VGND 0.02956f
C7671 XThC.XTB4.Y.t8 VGND 0.05016f
C7672 XThC.XTB4.Y.n13 VGND 0.08416f
C7673 XThC.XTB4.Y.n14 VGND 0.08889f
C7674 XThC.XTB4.Y.n15 VGND 0.03426f
C7675 XThC.XTB4.Y.n16 VGND 0.07234f
C7676 XThC.XTB4.Y.n17 VGND 0.0331f
C7677 XThC.XTB4.Y.n18 VGND 0.02701f
C7678 XThC.XTB4.Y.n19 VGND 0.63971f
C7679 XThC.XTB4.Y.n20 VGND 1.29767f
C7680 XThC.XTB4.Y.n21 VGND 0.08408f
C7681 XThC.XTB4.Y.t0 VGND 0.06491f
C7682 XThC.XTB4.Y.n22 VGND 0.04329f
C7683 XThC.Tn[0].n0 VGND 0.02911f
C7684 XThC.Tn[0].n1 VGND 0.01747f
C7685 XThC.Tn[0].n2 VGND 0.0832f
C7686 XThC.Tn[0].n3 VGND 0.01747f
C7687 XThC.Tn[0].n4 VGND 0.05143f
C7688 XThC.Tn[0].n5 VGND 0.01747f
C7689 XThC.Tn[0].n6 VGND 0.05805f
C7690 XThC.Tn[0].t22 VGND 0.01022f
C7691 XThC.Tn[0].n7 VGND 0.02282f
C7692 XThC.Tn[0].n8 VGND 0.01304f
C7693 XThC.Tn[0].n9 VGND 0.01586f
C7694 XThC.Tn[0].t41 VGND 0.01022f
C7695 XThC.Tn[0].n10 VGND 0.02282f
C7696 XThC.Tn[0].n11 VGND 0.01304f
C7697 XThC.Tn[0].n12 VGND 0.07535f
C7698 XThC.Tn[0].t12 VGND 0.01022f
C7699 XThC.Tn[0].n13 VGND 0.02282f
C7700 XThC.Tn[0].n14 VGND 0.01304f
C7701 XThC.Tn[0].n15 VGND 0.07535f
C7702 XThC.Tn[0].t13 VGND 0.01022f
C7703 XThC.Tn[0].n16 VGND 0.02282f
C7704 XThC.Tn[0].n17 VGND 0.01304f
C7705 XThC.Tn[0].n18 VGND 0.07535f
C7706 XThC.Tn[0].t32 VGND 0.01022f
C7707 XThC.Tn[0].n19 VGND 0.02282f
C7708 XThC.Tn[0].n20 VGND 0.01304f
C7709 XThC.Tn[0].n21 VGND 0.07535f
C7710 XThC.Tn[0].t34 VGND 0.01022f
C7711 XThC.Tn[0].n22 VGND 0.02282f
C7712 XThC.Tn[0].n23 VGND 0.01304f
C7713 XThC.Tn[0].n24 VGND 0.07535f
C7714 XThC.Tn[0].t17 VGND 0.01022f
C7715 XThC.Tn[0].n25 VGND 0.02282f
C7716 XThC.Tn[0].n26 VGND 0.01304f
C7717 XThC.Tn[0].n27 VGND 0.07535f
C7718 XThC.Tn[0].t25 VGND 0.01022f
C7719 XThC.Tn[0].n28 VGND 0.02282f
C7720 XThC.Tn[0].n29 VGND 0.01304f
C7721 XThC.Tn[0].n30 VGND 0.07535f
C7722 XThC.Tn[0].t26 VGND 0.01022f
C7723 XThC.Tn[0].n31 VGND 0.02282f
C7724 XThC.Tn[0].n32 VGND 0.01304f
C7725 XThC.Tn[0].n33 VGND 0.07535f
C7726 XThC.Tn[0].t15 VGND 0.01022f
C7727 XThC.Tn[0].n34 VGND 0.02282f
C7728 XThC.Tn[0].n35 VGND 0.01304f
C7729 XThC.Tn[0].n36 VGND 0.07535f
C7730 XThC.Tn[0].t16 VGND 0.01022f
C7731 XThC.Tn[0].n37 VGND 0.02282f
C7732 XThC.Tn[0].n38 VGND 0.01304f
C7733 XThC.Tn[0].n39 VGND 0.07535f
C7734 XThC.Tn[0].t27 VGND 0.01022f
C7735 XThC.Tn[0].n40 VGND 0.02282f
C7736 XThC.Tn[0].n41 VGND 0.01304f
C7737 XThC.Tn[0].n42 VGND 0.07535f
C7738 XThC.Tn[0].t36 VGND 0.01022f
C7739 XThC.Tn[0].n43 VGND 0.02282f
C7740 XThC.Tn[0].n44 VGND 0.01304f
C7741 XThC.Tn[0].n45 VGND 0.07535f
C7742 XThC.Tn[0].t38 VGND 0.01022f
C7743 XThC.Tn[0].n46 VGND 0.02282f
C7744 XThC.Tn[0].n47 VGND 0.01304f
C7745 XThC.Tn[0].n48 VGND 0.07535f
C7746 XThC.Tn[0].t19 VGND 0.01022f
C7747 XThC.Tn[0].n49 VGND 0.02282f
C7748 XThC.Tn[0].n50 VGND 0.01304f
C7749 XThC.Tn[0].n51 VGND 0.07535f
C7750 XThC.Tn[0].t29 VGND 0.01022f
C7751 XThC.Tn[0].n52 VGND 0.02282f
C7752 XThC.Tn[0].n53 VGND 0.01304f
C7753 XThC.Tn[0].n54 VGND 0.07535f
C7754 XThC.Tn[0].n55 VGND 0.13474f
C7755 XThC.Tn[0].n56 VGND 0.03416f
C7756 XThC.Tn[0].t1 VGND 0.0118f
C7757 XThC.Tn[0].t0 VGND 0.0118f
C7758 XThC.Tn[0].n57 VGND 0.02383f
C7759 XThC.Tn[0].t3 VGND 0.0118f
C7760 XThC.Tn[0].t2 VGND 0.0118f
C7761 XThC.Tn[0].n58 VGND 0.02788f
C7762 XThC.Tn[0].n59 VGND 0.07804f
C7763 XThC.Tn[0].n60 VGND 0.0247f
C7764 XThC.Tn[13].t6 VGND 0.01445f
C7765 XThC.Tn[13].t5 VGND 0.01445f
C7766 XThC.Tn[13].n0 VGND 0.03122f
C7767 XThC.Tn[13].t4 VGND 0.01445f
C7768 XThC.Tn[13].t7 VGND 0.01445f
C7769 XThC.Tn[13].n1 VGND 0.04921f
C7770 XThC.Tn[13].n2 VGND 0.13032f
C7771 XThC.Tn[13].t9 VGND 0.01445f
C7772 XThC.Tn[13].t8 VGND 0.01445f
C7773 XThC.Tn[13].n3 VGND 0.04387f
C7774 XThC.Tn[13].t11 VGND 0.01445f
C7775 XThC.Tn[13].t10 VGND 0.01445f
C7776 XThC.Tn[13].n4 VGND 0.03212f
C7777 XThC.Tn[13].n5 VGND 0.14294f
C7778 XThC.Tn[13].t29 VGND 0.01145f
C7779 XThC.Tn[13].t27 VGND 0.01251f
C7780 XThC.Tn[13].n7 VGND 0.02793f
C7781 XThC.Tn[13].n8 VGND 0.01596f
C7782 XThC.Tn[13].n9 VGND 0.01941f
C7783 XThC.Tn[13].t15 VGND 0.01145f
C7784 XThC.Tn[13].t12 VGND 0.01251f
C7785 XThC.Tn[13].n10 VGND 0.02793f
C7786 XThC.Tn[13].n11 VGND 0.01596f
C7787 XThC.Tn[13].n12 VGND 0.09223f
C7788 XThC.Tn[13].t20 VGND 0.01145f
C7789 XThC.Tn[13].t14 VGND 0.01251f
C7790 XThC.Tn[13].n13 VGND 0.02793f
C7791 XThC.Tn[13].n14 VGND 0.01596f
C7792 XThC.Tn[13].n15 VGND 0.09223f
C7793 XThC.Tn[13].t21 VGND 0.01145f
C7794 XThC.Tn[13].t16 VGND 0.01251f
C7795 XThC.Tn[13].n16 VGND 0.02793f
C7796 XThC.Tn[13].n17 VGND 0.01596f
C7797 XThC.Tn[13].n18 VGND 0.09223f
C7798 XThC.Tn[13].t40 VGND 0.01145f
C7799 XThC.Tn[13].t37 VGND 0.01251f
C7800 XThC.Tn[13].n19 VGND 0.02793f
C7801 XThC.Tn[13].n20 VGND 0.01596f
C7802 XThC.Tn[13].n21 VGND 0.09223f
C7803 XThC.Tn[13].t41 VGND 0.01145f
C7804 XThC.Tn[13].t38 VGND 0.01251f
C7805 XThC.Tn[13].n22 VGND 0.02793f
C7806 XThC.Tn[13].n23 VGND 0.01596f
C7807 XThC.Tn[13].n24 VGND 0.09223f
C7808 XThC.Tn[13].t25 VGND 0.01145f
C7809 XThC.Tn[13].t19 VGND 0.01251f
C7810 XThC.Tn[13].n25 VGND 0.02793f
C7811 XThC.Tn[13].n26 VGND 0.01596f
C7812 XThC.Tn[13].n27 VGND 0.09223f
C7813 XThC.Tn[13].t32 VGND 0.01145f
C7814 XThC.Tn[13].t28 VGND 0.01251f
C7815 XThC.Tn[13].n28 VGND 0.02793f
C7816 XThC.Tn[13].n29 VGND 0.01596f
C7817 XThC.Tn[13].n30 VGND 0.09223f
C7818 XThC.Tn[13].t34 VGND 0.01145f
C7819 XThC.Tn[13].t30 VGND 0.01251f
C7820 XThC.Tn[13].n31 VGND 0.02793f
C7821 XThC.Tn[13].n32 VGND 0.01596f
C7822 XThC.Tn[13].n33 VGND 0.09223f
C7823 XThC.Tn[13].t22 VGND 0.01145f
C7824 XThC.Tn[13].t17 VGND 0.01251f
C7825 XThC.Tn[13].n34 VGND 0.02793f
C7826 XThC.Tn[13].n35 VGND 0.01596f
C7827 XThC.Tn[13].n36 VGND 0.09223f
C7828 XThC.Tn[13].t24 VGND 0.01145f
C7829 XThC.Tn[13].t18 VGND 0.01251f
C7830 XThC.Tn[13].n37 VGND 0.02793f
C7831 XThC.Tn[13].n38 VGND 0.01596f
C7832 XThC.Tn[13].n39 VGND 0.09223f
C7833 XThC.Tn[13].t35 VGND 0.01145f
C7834 XThC.Tn[13].t31 VGND 0.01251f
C7835 XThC.Tn[13].n40 VGND 0.02793f
C7836 XThC.Tn[13].n41 VGND 0.01596f
C7837 XThC.Tn[13].n42 VGND 0.09223f
C7838 XThC.Tn[13].t43 VGND 0.01145f
C7839 XThC.Tn[13].t39 VGND 0.01251f
C7840 XThC.Tn[13].n43 VGND 0.02793f
C7841 XThC.Tn[13].n44 VGND 0.01596f
C7842 XThC.Tn[13].n45 VGND 0.09223f
C7843 XThC.Tn[13].t13 VGND 0.01145f
C7844 XThC.Tn[13].t42 VGND 0.01251f
C7845 XThC.Tn[13].n46 VGND 0.02793f
C7846 XThC.Tn[13].n47 VGND 0.01596f
C7847 XThC.Tn[13].n48 VGND 0.09223f
C7848 XThC.Tn[13].t26 VGND 0.01145f
C7849 XThC.Tn[13].t23 VGND 0.01251f
C7850 XThC.Tn[13].n49 VGND 0.02793f
C7851 XThC.Tn[13].n50 VGND 0.01596f
C7852 XThC.Tn[13].n51 VGND 0.09223f
C7853 XThC.Tn[13].t36 VGND 0.01145f
C7854 XThC.Tn[13].t33 VGND 0.01251f
C7855 XThC.Tn[13].n52 VGND 0.02793f
C7856 XThC.Tn[13].n53 VGND 0.01596f
C7857 XThC.Tn[13].n54 VGND 0.09223f
C7858 XThC.Tn[13].n55 VGND 0.51097f
C7859 XThC.Tn[13].n56 VGND 0.04181f
C7860 XThC.Tn[13].n57 VGND 0.01878f
C7861 XThC.Tn[13].n58 VGND 0.02342f
C7862 XThC.Tn[13].n59 VGND 0.04331f
C7863 XThC.Tn[12].n0 VGND 0.01883f
C7864 XThC.Tn[12].n1 VGND 0.02348f
C7865 XThC.Tn[12].n2 VGND 0.04736f
C7866 XThC.Tn[12].t5 VGND 0.01448f
C7867 XThC.Tn[12].t6 VGND 0.01448f
C7868 XThC.Tn[12].n3 VGND 0.03129f
C7869 XThC.Tn[12].t4 VGND 0.01448f
C7870 XThC.Tn[12].t7 VGND 0.01448f
C7871 XThC.Tn[12].n4 VGND 0.04762f
C7872 XThC.Tn[12].n5 VGND 0.13232f
C7873 XThC.Tn[12].t9 VGND 0.01448f
C7874 XThC.Tn[12].t8 VGND 0.01448f
C7875 XThC.Tn[12].n6 VGND 0.04397f
C7876 XThC.Tn[12].t11 VGND 0.01448f
C7877 XThC.Tn[12].t10 VGND 0.01448f
C7878 XThC.Tn[12].n7 VGND 0.03219f
C7879 XThC.Tn[12].n8 VGND 0.14328f
C7880 XThC.Tn[12].n9 VGND 0.02081f
C7881 XThC.Tn[12].t37 VGND 0.01148f
C7882 XThC.Tn[12].t35 VGND 0.01254f
C7883 XThC.Tn[12].n10 VGND 0.028f
C7884 XThC.Tn[12].n11 VGND 0.016f
C7885 XThC.Tn[12].n12 VGND 0.01946f
C7886 XThC.Tn[12].t23 VGND 0.01148f
C7887 XThC.Tn[12].t20 VGND 0.01254f
C7888 XThC.Tn[12].n13 VGND 0.028f
C7889 XThC.Tn[12].n14 VGND 0.016f
C7890 XThC.Tn[12].n15 VGND 0.09245f
C7891 XThC.Tn[12].t28 VGND 0.01148f
C7892 XThC.Tn[12].t22 VGND 0.01254f
C7893 XThC.Tn[12].n16 VGND 0.028f
C7894 XThC.Tn[12].n17 VGND 0.016f
C7895 XThC.Tn[12].n18 VGND 0.09245f
C7896 XThC.Tn[12].t29 VGND 0.01148f
C7897 XThC.Tn[12].t24 VGND 0.01254f
C7898 XThC.Tn[12].n19 VGND 0.028f
C7899 XThC.Tn[12].n20 VGND 0.016f
C7900 XThC.Tn[12].n21 VGND 0.09245f
C7901 XThC.Tn[12].t16 VGND 0.01148f
C7902 XThC.Tn[12].t13 VGND 0.01254f
C7903 XThC.Tn[12].n22 VGND 0.028f
C7904 XThC.Tn[12].n23 VGND 0.016f
C7905 XThC.Tn[12].n24 VGND 0.09245f
C7906 XThC.Tn[12].t17 VGND 0.01148f
C7907 XThC.Tn[12].t14 VGND 0.01254f
C7908 XThC.Tn[12].n25 VGND 0.028f
C7909 XThC.Tn[12].n26 VGND 0.016f
C7910 XThC.Tn[12].n27 VGND 0.09245f
C7911 XThC.Tn[12].t33 VGND 0.01148f
C7912 XThC.Tn[12].t27 VGND 0.01254f
C7913 XThC.Tn[12].n28 VGND 0.028f
C7914 XThC.Tn[12].n29 VGND 0.016f
C7915 XThC.Tn[12].n30 VGND 0.09245f
C7916 XThC.Tn[12].t40 VGND 0.01148f
C7917 XThC.Tn[12].t36 VGND 0.01254f
C7918 XThC.Tn[12].n31 VGND 0.028f
C7919 XThC.Tn[12].n32 VGND 0.016f
C7920 XThC.Tn[12].n33 VGND 0.09245f
C7921 XThC.Tn[12].t42 VGND 0.01148f
C7922 XThC.Tn[12].t38 VGND 0.01254f
C7923 XThC.Tn[12].n34 VGND 0.028f
C7924 XThC.Tn[12].n35 VGND 0.016f
C7925 XThC.Tn[12].n36 VGND 0.09245f
C7926 XThC.Tn[12].t30 VGND 0.01148f
C7927 XThC.Tn[12].t25 VGND 0.01254f
C7928 XThC.Tn[12].n37 VGND 0.028f
C7929 XThC.Tn[12].n38 VGND 0.016f
C7930 XThC.Tn[12].n39 VGND 0.09245f
C7931 XThC.Tn[12].t32 VGND 0.01148f
C7932 XThC.Tn[12].t26 VGND 0.01254f
C7933 XThC.Tn[12].n40 VGND 0.028f
C7934 XThC.Tn[12].n41 VGND 0.016f
C7935 XThC.Tn[12].n42 VGND 0.09245f
C7936 XThC.Tn[12].t43 VGND 0.01148f
C7937 XThC.Tn[12].t39 VGND 0.01254f
C7938 XThC.Tn[12].n43 VGND 0.028f
C7939 XThC.Tn[12].n44 VGND 0.016f
C7940 XThC.Tn[12].n45 VGND 0.09245f
C7941 XThC.Tn[12].t19 VGND 0.01148f
C7942 XThC.Tn[12].t15 VGND 0.01254f
C7943 XThC.Tn[12].n46 VGND 0.028f
C7944 XThC.Tn[12].n47 VGND 0.016f
C7945 XThC.Tn[12].n48 VGND 0.09245f
C7946 XThC.Tn[12].t21 VGND 0.01148f
C7947 XThC.Tn[12].t18 VGND 0.01254f
C7948 XThC.Tn[12].n49 VGND 0.028f
C7949 XThC.Tn[12].n50 VGND 0.016f
C7950 XThC.Tn[12].n51 VGND 0.09245f
C7951 XThC.Tn[12].t34 VGND 0.01148f
C7952 XThC.Tn[12].t31 VGND 0.01254f
C7953 XThC.Tn[12].n52 VGND 0.028f
C7954 XThC.Tn[12].n53 VGND 0.016f
C7955 XThC.Tn[12].n54 VGND 0.09245f
C7956 XThC.Tn[12].t12 VGND 0.01148f
C7957 XThC.Tn[12].t41 VGND 0.01254f
C7958 XThC.Tn[12].n55 VGND 0.028f
C7959 XThC.Tn[12].n56 VGND 0.016f
C7960 XThC.Tn[12].n57 VGND 0.09245f
C7961 XThC.Tn[12].n58 VGND 0.5067f
C7962 XThC.Tn[12].n59 VGND 0.03519f
C7963 XThC.Tn[11].n0 VGND 0.0239f
C7964 XThC.Tn[11].n1 VGND 0.01917f
C7965 XThC.Tn[11].n2 VGND 0.0442f
C7966 XThC.Tn[11].t20 VGND 0.01169f
C7967 XThC.Tn[11].t18 VGND 0.01277f
C7968 XThC.Tn[11].n3 VGND 0.02851f
C7969 XThC.Tn[11].n4 VGND 0.01629f
C7970 XThC.Tn[11].n5 VGND 0.01981f
C7971 XThC.Tn[11].t38 VGND 0.01169f
C7972 XThC.Tn[11].t35 VGND 0.01277f
C7973 XThC.Tn[11].n6 VGND 0.02851f
C7974 XThC.Tn[11].n7 VGND 0.01629f
C7975 XThC.Tn[11].n8 VGND 0.09412f
C7976 XThC.Tn[11].t43 VGND 0.01169f
C7977 XThC.Tn[11].t37 VGND 0.01277f
C7978 XThC.Tn[11].n9 VGND 0.02851f
C7979 XThC.Tn[11].n10 VGND 0.01629f
C7980 XThC.Tn[11].n11 VGND 0.09412f
C7981 XThC.Tn[11].t12 VGND 0.01169f
C7982 XThC.Tn[11].t39 VGND 0.01277f
C7983 XThC.Tn[11].n12 VGND 0.02851f
C7984 XThC.Tn[11].n13 VGND 0.01629f
C7985 XThC.Tn[11].n14 VGND 0.09412f
C7986 XThC.Tn[11].t31 VGND 0.01169f
C7987 XThC.Tn[11].t28 VGND 0.01277f
C7988 XThC.Tn[11].n15 VGND 0.02851f
C7989 XThC.Tn[11].n16 VGND 0.01629f
C7990 XThC.Tn[11].n17 VGND 0.09412f
C7991 XThC.Tn[11].t32 VGND 0.01169f
C7992 XThC.Tn[11].t29 VGND 0.01277f
C7993 XThC.Tn[11].n18 VGND 0.02851f
C7994 XThC.Tn[11].n19 VGND 0.01629f
C7995 XThC.Tn[11].n20 VGND 0.09412f
C7996 XThC.Tn[11].t16 VGND 0.01169f
C7997 XThC.Tn[11].t42 VGND 0.01277f
C7998 XThC.Tn[11].n21 VGND 0.02851f
C7999 XThC.Tn[11].n22 VGND 0.01629f
C8000 XThC.Tn[11].n23 VGND 0.09412f
C8001 XThC.Tn[11].t23 VGND 0.01169f
C8002 XThC.Tn[11].t19 VGND 0.01277f
C8003 XThC.Tn[11].n24 VGND 0.02851f
C8004 XThC.Tn[11].n25 VGND 0.01629f
C8005 XThC.Tn[11].n26 VGND 0.09412f
C8006 XThC.Tn[11].t25 VGND 0.01169f
C8007 XThC.Tn[11].t21 VGND 0.01277f
C8008 XThC.Tn[11].n27 VGND 0.02851f
C8009 XThC.Tn[11].n28 VGND 0.01629f
C8010 XThC.Tn[11].n29 VGND 0.09412f
C8011 XThC.Tn[11].t13 VGND 0.01169f
C8012 XThC.Tn[11].t40 VGND 0.01277f
C8013 XThC.Tn[11].n30 VGND 0.02851f
C8014 XThC.Tn[11].n31 VGND 0.01629f
C8015 XThC.Tn[11].n32 VGND 0.09412f
C8016 XThC.Tn[11].t15 VGND 0.01169f
C8017 XThC.Tn[11].t41 VGND 0.01277f
C8018 XThC.Tn[11].n33 VGND 0.02851f
C8019 XThC.Tn[11].n34 VGND 0.01629f
C8020 XThC.Tn[11].n35 VGND 0.09412f
C8021 XThC.Tn[11].t26 VGND 0.01169f
C8022 XThC.Tn[11].t22 VGND 0.01277f
C8023 XThC.Tn[11].n36 VGND 0.02851f
C8024 XThC.Tn[11].n37 VGND 0.01629f
C8025 XThC.Tn[11].n38 VGND 0.09412f
C8026 XThC.Tn[11].t34 VGND 0.01169f
C8027 XThC.Tn[11].t30 VGND 0.01277f
C8028 XThC.Tn[11].n39 VGND 0.02851f
C8029 XThC.Tn[11].n40 VGND 0.01629f
C8030 XThC.Tn[11].n41 VGND 0.09412f
C8031 XThC.Tn[11].t36 VGND 0.01169f
C8032 XThC.Tn[11].t33 VGND 0.01277f
C8033 XThC.Tn[11].n42 VGND 0.02851f
C8034 XThC.Tn[11].n43 VGND 0.01629f
C8035 XThC.Tn[11].n44 VGND 0.09412f
C8036 XThC.Tn[11].t17 VGND 0.01169f
C8037 XThC.Tn[11].t14 VGND 0.01277f
C8038 XThC.Tn[11].n45 VGND 0.02851f
C8039 XThC.Tn[11].n46 VGND 0.01629f
C8040 XThC.Tn[11].n47 VGND 0.09412f
C8041 XThC.Tn[11].t27 VGND 0.01169f
C8042 XThC.Tn[11].t24 VGND 0.01277f
C8043 XThC.Tn[11].n48 VGND 0.02851f
C8044 XThC.Tn[11].n49 VGND 0.01629f
C8045 XThC.Tn[11].n50 VGND 0.09412f
C8046 XThC.Tn[11].n51 VGND 0.04302f
C8047 XThC.Tn[11].t8 VGND 0.01474f
C8048 XThC.Tn[11].t5 VGND 0.01474f
C8049 XThC.Tn[11].n52 VGND 0.03186f
C8050 XThC.Tn[11].t0 VGND 0.01474f
C8051 XThC.Tn[11].t11 VGND 0.01474f
C8052 XThC.Tn[11].n53 VGND 0.05022f
C8053 XThC.Tn[11].n54 VGND 0.13299f
C8054 XThC.Tn[11].t1 VGND 0.01474f
C8055 XThC.Tn[11].t4 VGND 0.01474f
C8056 XThC.Tn[11].n56 VGND 0.04477f
C8057 XThC.Tn[11].t3 VGND 0.01474f
C8058 XThC.Tn[11].t2 VGND 0.01474f
C8059 XThC.Tn[11].n57 VGND 0.03278f
C8060 XThC.Tn[11].n58 VGND 0.14588f
C8061 XThC.Tn[9].t4 VGND 0.01469f
C8062 XThC.Tn[9].t7 VGND 0.01469f
C8063 XThC.Tn[9].n0 VGND 0.03174f
C8064 XThC.Tn[9].t6 VGND 0.01469f
C8065 XThC.Tn[9].t5 VGND 0.01469f
C8066 XThC.Tn[9].n1 VGND 0.05003f
C8067 XThC.Tn[9].n2 VGND 0.1325f
C8068 XThC.Tn[9].t9 VGND 0.01469f
C8069 XThC.Tn[9].t8 VGND 0.01469f
C8070 XThC.Tn[9].n3 VGND 0.0446f
C8071 XThC.Tn[9].t11 VGND 0.01469f
C8072 XThC.Tn[9].t10 VGND 0.01469f
C8073 XThC.Tn[9].n4 VGND 0.03266f
C8074 XThC.Tn[9].n5 VGND 0.14534f
C8075 XThC.Tn[9].t26 VGND 0.01164f
C8076 XThC.Tn[9].t12 VGND 0.01272f
C8077 XThC.Tn[9].n7 VGND 0.0284f
C8078 XThC.Tn[9].n8 VGND 0.01623f
C8079 XThC.Tn[9].n9 VGND 0.01974f
C8080 XThC.Tn[9].t13 VGND 0.01164f
C8081 XThC.Tn[9].t30 VGND 0.01272f
C8082 XThC.Tn[9].n10 VGND 0.0284f
C8083 XThC.Tn[9].n11 VGND 0.01623f
C8084 XThC.Tn[9].n12 VGND 0.09378f
C8085 XThC.Tn[9].t15 VGND 0.01164f
C8086 XThC.Tn[9].t34 VGND 0.01272f
C8087 XThC.Tn[9].n13 VGND 0.0284f
C8088 XThC.Tn[9].n14 VGND 0.01623f
C8089 XThC.Tn[9].n15 VGND 0.09378f
C8090 XThC.Tn[9].t17 VGND 0.01164f
C8091 XThC.Tn[9].t35 VGND 0.01272f
C8092 XThC.Tn[9].n16 VGND 0.0284f
C8093 XThC.Tn[9].n17 VGND 0.01623f
C8094 XThC.Tn[9].n18 VGND 0.09378f
C8095 XThC.Tn[9].t39 VGND 0.01164f
C8096 XThC.Tn[9].t24 VGND 0.01272f
C8097 XThC.Tn[9].n19 VGND 0.0284f
C8098 XThC.Tn[9].n20 VGND 0.01623f
C8099 XThC.Tn[9].n21 VGND 0.09378f
C8100 XThC.Tn[9].t40 VGND 0.01164f
C8101 XThC.Tn[9].t25 VGND 0.01272f
C8102 XThC.Tn[9].n22 VGND 0.0284f
C8103 XThC.Tn[9].n23 VGND 0.01623f
C8104 XThC.Tn[9].n24 VGND 0.09378f
C8105 XThC.Tn[9].t22 VGND 0.01164f
C8106 XThC.Tn[9].t38 VGND 0.01272f
C8107 XThC.Tn[9].n25 VGND 0.0284f
C8108 XThC.Tn[9].n26 VGND 0.01623f
C8109 XThC.Tn[9].n27 VGND 0.09378f
C8110 XThC.Tn[9].t28 VGND 0.01164f
C8111 XThC.Tn[9].t14 VGND 0.01272f
C8112 XThC.Tn[9].n28 VGND 0.0284f
C8113 XThC.Tn[9].n29 VGND 0.01623f
C8114 XThC.Tn[9].n30 VGND 0.09378f
C8115 XThC.Tn[9].t31 VGND 0.01164f
C8116 XThC.Tn[9].t16 VGND 0.01272f
C8117 XThC.Tn[9].n31 VGND 0.0284f
C8118 XThC.Tn[9].n32 VGND 0.01623f
C8119 XThC.Tn[9].n33 VGND 0.09378f
C8120 XThC.Tn[9].t19 VGND 0.01164f
C8121 XThC.Tn[9].t36 VGND 0.01272f
C8122 XThC.Tn[9].n34 VGND 0.0284f
C8123 XThC.Tn[9].n35 VGND 0.01623f
C8124 XThC.Tn[9].n36 VGND 0.09378f
C8125 XThC.Tn[9].t21 VGND 0.01164f
C8126 XThC.Tn[9].t37 VGND 0.01272f
C8127 XThC.Tn[9].n37 VGND 0.0284f
C8128 XThC.Tn[9].n38 VGND 0.01623f
C8129 XThC.Tn[9].n39 VGND 0.09378f
C8130 XThC.Tn[9].t32 VGND 0.01164f
C8131 XThC.Tn[9].t18 VGND 0.01272f
C8132 XThC.Tn[9].n40 VGND 0.0284f
C8133 XThC.Tn[9].n41 VGND 0.01623f
C8134 XThC.Tn[9].n42 VGND 0.09378f
C8135 XThC.Tn[9].t42 VGND 0.01164f
C8136 XThC.Tn[9].t27 VGND 0.01272f
C8137 XThC.Tn[9].n43 VGND 0.0284f
C8138 XThC.Tn[9].n44 VGND 0.01623f
C8139 XThC.Tn[9].n45 VGND 0.09378f
C8140 XThC.Tn[9].t43 VGND 0.01164f
C8141 XThC.Tn[9].t29 VGND 0.01272f
C8142 XThC.Tn[9].n46 VGND 0.0284f
C8143 XThC.Tn[9].n47 VGND 0.01623f
C8144 XThC.Tn[9].n48 VGND 0.09378f
C8145 XThC.Tn[9].t23 VGND 0.01164f
C8146 XThC.Tn[9].t41 VGND 0.01272f
C8147 XThC.Tn[9].n49 VGND 0.0284f
C8148 XThC.Tn[9].n50 VGND 0.01623f
C8149 XThC.Tn[9].n51 VGND 0.09378f
C8150 XThC.Tn[9].t33 VGND 0.01164f
C8151 XThC.Tn[9].t20 VGND 0.01272f
C8152 XThC.Tn[9].n52 VGND 0.0284f
C8153 XThC.Tn[9].n53 VGND 0.01623f
C8154 XThC.Tn[9].n54 VGND 0.09378f
C8155 XThC.Tn[9].n55 VGND 0.04286f
C8156 XThC.Tn[9].n56 VGND 0.02381f
C8157 XThC.Tn[9].n57 VGND 0.0191f
C8158 XThC.Tn[9].n58 VGND 0.04403f
C8159 XThC.Tn[5].t7 VGND 0.0121f
C8160 XThC.Tn[5].t6 VGND 0.0121f
C8161 XThC.Tn[5].n0 VGND 0.02443f
C8162 XThC.Tn[5].t5 VGND 0.0121f
C8163 XThC.Tn[5].t4 VGND 0.0121f
C8164 XThC.Tn[5].n1 VGND 0.02858f
C8165 XThC.Tn[5].n2 VGND 0.08573f
C8166 XThC.Tn[5].n3 VGND 0.01791f
C8167 XThC.Tn[5].n4 VGND 0.01791f
C8168 XThC.Tn[5].n5 VGND 0.01791f
C8169 XThC.Tn[5].n6 VGND 0.02985f
C8170 XThC.Tn[5].n7 VGND 0.0853f
C8171 XThC.Tn[5].n8 VGND 0.05273f
C8172 XThC.Tn[5].n9 VGND 0.05951f
C8173 XThC.Tn[5].t33 VGND 0.01048f
C8174 XThC.Tn[5].n10 VGND 0.0234f
C8175 XThC.Tn[5].n11 VGND 0.01337f
C8176 XThC.Tn[5].n12 VGND 0.01626f
C8177 XThC.Tn[5].t19 VGND 0.01048f
C8178 XThC.Tn[5].n13 VGND 0.0234f
C8179 XThC.Tn[5].n14 VGND 0.01337f
C8180 XThC.Tn[5].n15 VGND 0.07725f
C8181 XThC.Tn[5].t23 VGND 0.01048f
C8182 XThC.Tn[5].n16 VGND 0.0234f
C8183 XThC.Tn[5].n17 VGND 0.01337f
C8184 XThC.Tn[5].n18 VGND 0.07725f
C8185 XThC.Tn[5].t24 VGND 0.01048f
C8186 XThC.Tn[5].n19 VGND 0.0234f
C8187 XThC.Tn[5].n20 VGND 0.01337f
C8188 XThC.Tn[5].n21 VGND 0.07725f
C8189 XThC.Tn[5].t13 VGND 0.01048f
C8190 XThC.Tn[5].n22 VGND 0.0234f
C8191 XThC.Tn[5].n23 VGND 0.01337f
C8192 XThC.Tn[5].n24 VGND 0.07725f
C8193 XThC.Tn[5].t14 VGND 0.01048f
C8194 XThC.Tn[5].n25 VGND 0.0234f
C8195 XThC.Tn[5].n26 VGND 0.01337f
C8196 XThC.Tn[5].n27 VGND 0.07725f
C8197 XThC.Tn[5].t27 VGND 0.01048f
C8198 XThC.Tn[5].n28 VGND 0.0234f
C8199 XThC.Tn[5].n29 VGND 0.01337f
C8200 XThC.Tn[5].n30 VGND 0.07725f
C8201 XThC.Tn[5].t35 VGND 0.01048f
C8202 XThC.Tn[5].n31 VGND 0.0234f
C8203 XThC.Tn[5].n32 VGND 0.01337f
C8204 XThC.Tn[5].n33 VGND 0.07725f
C8205 XThC.Tn[5].t37 VGND 0.01048f
C8206 XThC.Tn[5].n34 VGND 0.0234f
C8207 XThC.Tn[5].n35 VGND 0.01337f
C8208 XThC.Tn[5].n36 VGND 0.07725f
C8209 XThC.Tn[5].t25 VGND 0.01048f
C8210 XThC.Tn[5].n37 VGND 0.0234f
C8211 XThC.Tn[5].n38 VGND 0.01337f
C8212 XThC.Tn[5].n39 VGND 0.07725f
C8213 XThC.Tn[5].t26 VGND 0.01048f
C8214 XThC.Tn[5].n40 VGND 0.0234f
C8215 XThC.Tn[5].n41 VGND 0.01337f
C8216 XThC.Tn[5].n42 VGND 0.07725f
C8217 XThC.Tn[5].t39 VGND 0.01048f
C8218 XThC.Tn[5].n43 VGND 0.0234f
C8219 XThC.Tn[5].n44 VGND 0.01337f
C8220 XThC.Tn[5].n45 VGND 0.07725f
C8221 XThC.Tn[5].t16 VGND 0.01048f
C8222 XThC.Tn[5].n46 VGND 0.0234f
C8223 XThC.Tn[5].n47 VGND 0.01337f
C8224 XThC.Tn[5].n48 VGND 0.07725f
C8225 XThC.Tn[5].t18 VGND 0.01048f
C8226 XThC.Tn[5].n49 VGND 0.0234f
C8227 XThC.Tn[5].n50 VGND 0.01337f
C8228 XThC.Tn[5].n51 VGND 0.07725f
C8229 XThC.Tn[5].t30 VGND 0.01048f
C8230 XThC.Tn[5].n52 VGND 0.0234f
C8231 XThC.Tn[5].n53 VGND 0.01337f
C8232 XThC.Tn[5].n54 VGND 0.07725f
C8233 XThC.Tn[5].t41 VGND 0.01048f
C8234 XThC.Tn[5].n55 VGND 0.0234f
C8235 XThC.Tn[5].n56 VGND 0.01337f
C8236 XThC.Tn[5].n57 VGND 0.07725f
C8237 XThC.Tn[5].n58 VGND 0.2186f
C8238 XThC.Tn[5].n59 VGND 0.04035f
C8239 XThR.Tn[9].t0 VGND 0.01255f
C8240 XThR.Tn[9].t2 VGND 0.01255f
C8241 XThR.Tn[9].n0 VGND 0.0251f
C8242 XThR.Tn[9].t1 VGND 0.01255f
C8243 XThR.Tn[9].t3 VGND 0.01255f
C8244 XThR.Tn[9].n1 VGND 0.03131f
C8245 XThR.Tn[9].n2 VGND 0.06315f
C8246 XThR.Tn[9].t10 VGND 0.01931f
C8247 XThR.Tn[9].t8 VGND 0.01931f
C8248 XThR.Tn[9].n3 VGND 0.05863f
C8249 XThR.Tn[9].t11 VGND 0.01931f
C8250 XThR.Tn[9].t9 VGND 0.01931f
C8251 XThR.Tn[9].n4 VGND 0.04293f
C8252 XThR.Tn[9].n5 VGND 0.19519f
C8253 XThR.Tn[9].t6 VGND 0.01931f
C8254 XThR.Tn[9].t4 VGND 0.01931f
C8255 XThR.Tn[9].n6 VGND 0.04172f
C8256 XThR.Tn[9].t7 VGND 0.01931f
C8257 XThR.Tn[9].t5 VGND 0.01931f
C8258 XThR.Tn[9].n7 VGND 0.0635f
C8259 XThR.Tn[9].n8 VGND 0.17633f
C8260 XThR.Tn[9].n9 VGND 0.02361f
C8261 XThR.Tn[9].t17 VGND 0.01509f
C8262 XThR.Tn[9].t71 VGND 0.01653f
C8263 XThR.Tn[9].n10 VGND 0.04036f
C8264 XThR.Tn[9].n11 VGND 0.07752f
C8265 XThR.Tn[9].t35 VGND 0.01509f
C8266 XThR.Tn[9].t28 VGND 0.01653f
C8267 XThR.Tn[9].n12 VGND 0.04036f
C8268 XThR.Tn[9].t50 VGND 0.01504f
C8269 XThR.Tn[9].t19 VGND 0.01647f
C8270 XThR.Tn[9].n13 VGND 0.04199f
C8271 XThR.Tn[9].n14 VGND 0.0295f
C8272 XThR.Tn[9].n16 VGND 0.09466f
C8273 XThR.Tn[9].t72 VGND 0.01509f
C8274 XThR.Tn[9].t64 VGND 0.01653f
C8275 XThR.Tn[9].n17 VGND 0.04036f
C8276 XThR.Tn[9].t26 VGND 0.01504f
C8277 XThR.Tn[9].t59 VGND 0.01647f
C8278 XThR.Tn[9].n18 VGND 0.04199f
C8279 XThR.Tn[9].n19 VGND 0.0295f
C8280 XThR.Tn[9].n21 VGND 0.09466f
C8281 XThR.Tn[9].t29 VGND 0.01509f
C8282 XThR.Tn[9].t21 VGND 0.01653f
C8283 XThR.Tn[9].n22 VGND 0.04036f
C8284 XThR.Tn[9].t41 VGND 0.01504f
C8285 XThR.Tn[9].t15 VGND 0.01647f
C8286 XThR.Tn[9].n23 VGND 0.04199f
C8287 XThR.Tn[9].n24 VGND 0.0295f
C8288 XThR.Tn[9].n26 VGND 0.09466f
C8289 XThR.Tn[9].t56 VGND 0.01509f
C8290 XThR.Tn[9].t46 VGND 0.01653f
C8291 XThR.Tn[9].n27 VGND 0.04036f
C8292 XThR.Tn[9].t73 VGND 0.01504f
C8293 XThR.Tn[9].t42 VGND 0.01647f
C8294 XThR.Tn[9].n28 VGND 0.04199f
C8295 XThR.Tn[9].n29 VGND 0.0295f
C8296 XThR.Tn[9].n31 VGND 0.09466f
C8297 XThR.Tn[9].t31 VGND 0.01509f
C8298 XThR.Tn[9].t23 VGND 0.01653f
C8299 XThR.Tn[9].n32 VGND 0.04036f
C8300 XThR.Tn[9].t44 VGND 0.01504f
C8301 XThR.Tn[9].t16 VGND 0.01647f
C8302 XThR.Tn[9].n33 VGND 0.04199f
C8303 XThR.Tn[9].n34 VGND 0.0295f
C8304 XThR.Tn[9].n36 VGND 0.09466f
C8305 XThR.Tn[9].t67 VGND 0.01509f
C8306 XThR.Tn[9].t37 VGND 0.01653f
C8307 XThR.Tn[9].n37 VGND 0.04036f
C8308 XThR.Tn[9].t20 VGND 0.01504f
C8309 XThR.Tn[9].t33 VGND 0.01647f
C8310 XThR.Tn[9].n38 VGND 0.04199f
C8311 XThR.Tn[9].n39 VGND 0.0295f
C8312 XThR.Tn[9].n41 VGND 0.09466f
C8313 XThR.Tn[9].t36 VGND 0.01509f
C8314 XThR.Tn[9].t32 VGND 0.01653f
C8315 XThR.Tn[9].n42 VGND 0.04036f
C8316 XThR.Tn[9].t51 VGND 0.01504f
C8317 XThR.Tn[9].t25 VGND 0.01647f
C8318 XThR.Tn[9].n43 VGND 0.04199f
C8319 XThR.Tn[9].n44 VGND 0.0295f
C8320 XThR.Tn[9].n46 VGND 0.09466f
C8321 XThR.Tn[9].t39 VGND 0.01509f
C8322 XThR.Tn[9].t45 VGND 0.01653f
C8323 XThR.Tn[9].n47 VGND 0.04036f
C8324 XThR.Tn[9].t55 VGND 0.01504f
C8325 XThR.Tn[9].t40 VGND 0.01647f
C8326 XThR.Tn[9].n48 VGND 0.04199f
C8327 XThR.Tn[9].n49 VGND 0.0295f
C8328 XThR.Tn[9].n51 VGND 0.09466f
C8329 XThR.Tn[9].t58 VGND 0.01509f
C8330 XThR.Tn[9].t66 VGND 0.01653f
C8331 XThR.Tn[9].n52 VGND 0.04036f
C8332 XThR.Tn[9].t13 VGND 0.01504f
C8333 XThR.Tn[9].t60 VGND 0.01647f
C8334 XThR.Tn[9].n53 VGND 0.04199f
C8335 XThR.Tn[9].n54 VGND 0.0295f
C8336 XThR.Tn[9].n56 VGND 0.09466f
C8337 XThR.Tn[9].t48 VGND 0.01509f
C8338 XThR.Tn[9].t24 VGND 0.01653f
C8339 XThR.Tn[9].n57 VGND 0.04036f
C8340 XThR.Tn[9].t65 VGND 0.01504f
C8341 XThR.Tn[9].t18 VGND 0.01647f
C8342 XThR.Tn[9].n58 VGND 0.04199f
C8343 XThR.Tn[9].n59 VGND 0.0295f
C8344 XThR.Tn[9].n61 VGND 0.09466f
C8345 XThR.Tn[9].t70 VGND 0.01509f
C8346 XThR.Tn[9].t62 VGND 0.01653f
C8347 XThR.Tn[9].n62 VGND 0.04036f
C8348 XThR.Tn[9].t22 VGND 0.01504f
C8349 XThR.Tn[9].t52 VGND 0.01647f
C8350 XThR.Tn[9].n63 VGND 0.04199f
C8351 XThR.Tn[9].n64 VGND 0.0295f
C8352 XThR.Tn[9].n66 VGND 0.09466f
C8353 XThR.Tn[9].t38 VGND 0.01509f
C8354 XThR.Tn[9].t34 VGND 0.01653f
C8355 XThR.Tn[9].n67 VGND 0.04036f
C8356 XThR.Tn[9].t53 VGND 0.01504f
C8357 XThR.Tn[9].t27 VGND 0.01647f
C8358 XThR.Tn[9].n68 VGND 0.04199f
C8359 XThR.Tn[9].n69 VGND 0.0295f
C8360 XThR.Tn[9].n71 VGND 0.09466f
C8361 XThR.Tn[9].t57 VGND 0.01509f
C8362 XThR.Tn[9].t47 VGND 0.01653f
C8363 XThR.Tn[9].n72 VGND 0.04036f
C8364 XThR.Tn[9].t12 VGND 0.01504f
C8365 XThR.Tn[9].t43 VGND 0.01647f
C8366 XThR.Tn[9].n73 VGND 0.04199f
C8367 XThR.Tn[9].n74 VGND 0.0295f
C8368 XThR.Tn[9].n76 VGND 0.09466f
C8369 XThR.Tn[9].t14 VGND 0.01509f
C8370 XThR.Tn[9].t69 VGND 0.01653f
C8371 XThR.Tn[9].n77 VGND 0.04036f
C8372 XThR.Tn[9].t30 VGND 0.01504f
C8373 XThR.Tn[9].t61 VGND 0.01647f
C8374 XThR.Tn[9].n78 VGND 0.04199f
C8375 XThR.Tn[9].n79 VGND 0.0295f
C8376 XThR.Tn[9].n81 VGND 0.09466f
C8377 XThR.Tn[9].t49 VGND 0.01509f
C8378 XThR.Tn[9].t63 VGND 0.01653f
C8379 XThR.Tn[9].n82 VGND 0.04036f
C8380 XThR.Tn[9].t68 VGND 0.01504f
C8381 XThR.Tn[9].t54 VGND 0.01647f
C8382 XThR.Tn[9].n83 VGND 0.04199f
C8383 XThR.Tn[9].n84 VGND 0.0295f
C8384 XThR.Tn[9].n86 VGND 0.09466f
C8385 XThR.Tn[9].n87 VGND 0.08603f
C8386 XThR.Tn[9].n88 VGND 0.27907f
C8387 XThC.Tn[6].t7 VGND 0.01221f
C8388 XThC.Tn[6].t6 VGND 0.01221f
C8389 XThC.Tn[6].n0 VGND 0.02464f
C8390 XThC.Tn[6].t5 VGND 0.01221f
C8391 XThC.Tn[6].t4 VGND 0.01221f
C8392 XThC.Tn[6].n1 VGND 0.02883f
C8393 XThC.Tn[6].n2 VGND 0.0807f
C8394 XThC.Tn[6].n3 VGND 0.01807f
C8395 XThC.Tn[6].n4 VGND 0.01807f
C8396 XThC.Tn[6].n5 VGND 0.01807f
C8397 XThC.Tn[6].n6 VGND 0.0301f
C8398 XThC.Tn[6].n7 VGND 0.08604f
C8399 XThC.Tn[6].n8 VGND 0.05319f
C8400 XThC.Tn[6].n9 VGND 0.06003f
C8401 XThC.Tn[6].t26 VGND 0.01057f
C8402 XThC.Tn[6].n10 VGND 0.0236f
C8403 XThC.Tn[6].n11 VGND 0.01349f
C8404 XThC.Tn[6].n12 VGND 0.0164f
C8405 XThC.Tn[6].t13 VGND 0.01057f
C8406 XThC.Tn[6].n13 VGND 0.0236f
C8407 XThC.Tn[6].n14 VGND 0.01349f
C8408 XThC.Tn[6].n15 VGND 0.07792f
C8409 XThC.Tn[6].t17 VGND 0.01057f
C8410 XThC.Tn[6].n16 VGND 0.0236f
C8411 XThC.Tn[6].n17 VGND 0.01349f
C8412 XThC.Tn[6].n18 VGND 0.07792f
C8413 XThC.Tn[6].t18 VGND 0.01057f
C8414 XThC.Tn[6].n19 VGND 0.0236f
C8415 XThC.Tn[6].n20 VGND 0.01349f
C8416 XThC.Tn[6].n21 VGND 0.07792f
C8417 XThC.Tn[6].t37 VGND 0.01057f
C8418 XThC.Tn[6].n22 VGND 0.0236f
C8419 XThC.Tn[6].n23 VGND 0.01349f
C8420 XThC.Tn[6].n24 VGND 0.07792f
C8421 XThC.Tn[6].t38 VGND 0.01057f
C8422 XThC.Tn[6].n25 VGND 0.0236f
C8423 XThC.Tn[6].n26 VGND 0.01349f
C8424 XThC.Tn[6].n27 VGND 0.07792f
C8425 XThC.Tn[6].t22 VGND 0.01057f
C8426 XThC.Tn[6].n28 VGND 0.0236f
C8427 XThC.Tn[6].n29 VGND 0.01349f
C8428 XThC.Tn[6].n30 VGND 0.07792f
C8429 XThC.Tn[6].t29 VGND 0.01057f
C8430 XThC.Tn[6].n31 VGND 0.0236f
C8431 XThC.Tn[6].n32 VGND 0.01349f
C8432 XThC.Tn[6].n33 VGND 0.07792f
C8433 XThC.Tn[6].t31 VGND 0.01057f
C8434 XThC.Tn[6].n34 VGND 0.0236f
C8435 XThC.Tn[6].n35 VGND 0.01349f
C8436 XThC.Tn[6].n36 VGND 0.07792f
C8437 XThC.Tn[6].t19 VGND 0.01057f
C8438 XThC.Tn[6].n37 VGND 0.0236f
C8439 XThC.Tn[6].n38 VGND 0.01349f
C8440 XThC.Tn[6].n39 VGND 0.07792f
C8441 XThC.Tn[6].t21 VGND 0.01057f
C8442 XThC.Tn[6].n40 VGND 0.0236f
C8443 XThC.Tn[6].n41 VGND 0.01349f
C8444 XThC.Tn[6].n42 VGND 0.07792f
C8445 XThC.Tn[6].t32 VGND 0.01057f
C8446 XThC.Tn[6].n43 VGND 0.0236f
C8447 XThC.Tn[6].n44 VGND 0.01349f
C8448 XThC.Tn[6].n45 VGND 0.07792f
C8449 XThC.Tn[6].t41 VGND 0.01057f
C8450 XThC.Tn[6].n46 VGND 0.0236f
C8451 XThC.Tn[6].n47 VGND 0.01349f
C8452 XThC.Tn[6].n48 VGND 0.07792f
C8453 XThC.Tn[6].t43 VGND 0.01057f
C8454 XThC.Tn[6].n49 VGND 0.0236f
C8455 XThC.Tn[6].n50 VGND 0.01349f
C8456 XThC.Tn[6].n51 VGND 0.07792f
C8457 XThC.Tn[6].t24 VGND 0.01057f
C8458 XThC.Tn[6].n52 VGND 0.0236f
C8459 XThC.Tn[6].n53 VGND 0.01349f
C8460 XThC.Tn[6].n54 VGND 0.07792f
C8461 XThC.Tn[6].t34 VGND 0.01057f
C8462 XThC.Tn[6].n55 VGND 0.0236f
C8463 XThC.Tn[6].n56 VGND 0.01349f
C8464 XThC.Tn[6].n57 VGND 0.07792f
C8465 XThC.Tn[6].n58 VGND 0.20284f
C8466 XThC.Tn[6].n59 VGND 0.04609f
C8467 XThC.Tn[6].n60 VGND 0.02554f
C8468 XThC.XTBN.Y.n0 VGND 0.01531f
C8469 XThC.XTBN.Y.t50 VGND 0.01024f
C8470 XThC.XTBN.Y.t18 VGND 0.01024f
C8471 XThC.XTBN.Y.n1 VGND 0.01477f
C8472 XThC.XTBN.Y.t120 VGND 0.01024f
C8473 XThC.XTBN.Y.t114 VGND 0.01024f
C8474 XThC.XTBN.Y.n3 VGND 0.0138f
C8475 XThC.XTBN.Y.n5 VGND 0.01477f
C8476 XThC.XTBN.Y.n10 VGND 0.02164f
C8477 XThC.XTBN.Y.t79 VGND 0.01024f
C8478 XThC.XTBN.Y.t36 VGND 0.01024f
C8479 XThC.XTBN.Y.n13 VGND 0.01477f
C8480 XThC.XTBN.Y.t26 VGND 0.01024f
C8481 XThC.XTBN.Y.t21 VGND 0.01024f
C8482 XThC.XTBN.Y.n15 VGND 0.0138f
C8483 XThC.XTBN.Y.n17 VGND 0.01477f
C8484 XThC.XTBN.Y.n22 VGND 0.02164f
C8485 XThC.XTBN.Y.n25 VGND 0.11789f
C8486 XThC.XTBN.Y.t106 VGND 0.01024f
C8487 XThC.XTBN.Y.t70 VGND 0.01024f
C8488 XThC.XTBN.Y.n26 VGND 0.01477f
C8489 XThC.XTBN.Y.t56 VGND 0.01024f
C8490 XThC.XTBN.Y.t48 VGND 0.01024f
C8491 XThC.XTBN.Y.n28 VGND 0.0138f
C8492 XThC.XTBN.Y.n30 VGND 0.01477f
C8493 XThC.XTBN.Y.n35 VGND 0.02164f
C8494 XThC.XTBN.Y.n38 VGND 0.07443f
C8495 XThC.XTBN.Y.t39 VGND 0.01024f
C8496 XThC.XTBN.Y.t122 VGND 0.01024f
C8497 XThC.XTBN.Y.n39 VGND 0.01477f
C8498 XThC.XTBN.Y.t109 VGND 0.01024f
C8499 XThC.XTBN.Y.t102 VGND 0.01024f
C8500 XThC.XTBN.Y.n41 VGND 0.0138f
C8501 XThC.XTBN.Y.n43 VGND 0.01477f
C8502 XThC.XTBN.Y.n48 VGND 0.02164f
C8503 XThC.XTBN.Y.n51 VGND 0.07443f
C8504 XThC.XTBN.Y.t47 VGND 0.01024f
C8505 XThC.XTBN.Y.t17 VGND 0.01024f
C8506 XThC.XTBN.Y.n52 VGND 0.01477f
C8507 XThC.XTBN.Y.t116 VGND 0.01024f
C8508 XThC.XTBN.Y.t111 VGND 0.01024f
C8509 XThC.XTBN.Y.n54 VGND 0.0138f
C8510 XThC.XTBN.Y.n56 VGND 0.01477f
C8511 XThC.XTBN.Y.n61 VGND 0.02164f
C8512 XThC.XTBN.Y.n64 VGND 0.07443f
C8513 XThC.XTBN.Y.t101 VGND 0.01024f
C8514 XThC.XTBN.Y.t63 VGND 0.01024f
C8515 XThC.XTBN.Y.n65 VGND 0.01477f
C8516 XThC.XTBN.Y.t52 VGND 0.01024f
C8517 XThC.XTBN.Y.t44 VGND 0.01024f
C8518 XThC.XTBN.Y.n67 VGND 0.0138f
C8519 XThC.XTBN.Y.n69 VGND 0.01477f
C8520 XThC.XTBN.Y.n74 VGND 0.02164f
C8521 XThC.XTBN.Y.n77 VGND 0.07443f
C8522 XThC.XTBN.Y.t25 VGND 0.01024f
C8523 XThC.XTBN.Y.t100 VGND 0.01024f
C8524 XThC.XTBN.Y.n78 VGND 0.01477f
C8525 XThC.XTBN.Y.t93 VGND 0.01024f
C8526 XThC.XTBN.Y.t90 VGND 0.01024f
C8527 XThC.XTBN.Y.n80 VGND 0.0138f
C8528 XThC.XTBN.Y.n82 VGND 0.01477f
C8529 XThC.XTBN.Y.n87 VGND 0.02164f
C8530 XThC.XTBN.Y.n90 VGND 0.06646f
C8531 XThC.XTBN.Y.t46 VGND 0.01024f
C8532 XThC.XTBN.Y.t6 VGND 0.01024f
C8533 XThC.XTBN.Y.n92 VGND 0.01243f
C8534 XThC.XTBN.Y.t12 VGND 0.01024f
C8535 XThC.XTBN.Y.n93 VGND 0.01348f
C8536 XThC.XTBN.Y.n95 VGND 0.01252f
C8537 XThC.XTBN.Y.n98 VGND 0.01348f
C8538 XThC.XTBN.Y.t54 VGND 0.01024f
C8539 XThC.XTBN.Y.n99 VGND 0.01227f
C8540 XThC.XTBN.Y.n101 VGND 0.01009f
C8541 XThC.XTBN.Y.t38 VGND 0.01024f
C8542 XThC.XTBN.Y.t113 VGND 0.01024f
C8543 XThC.XTBN.Y.n103 VGND 0.01243f
C8544 XThC.XTBN.Y.t119 VGND 0.01024f
C8545 XThC.XTBN.Y.n104 VGND 0.01348f
C8546 XThC.XTBN.Y.n106 VGND 0.01252f
C8547 XThC.XTBN.Y.n109 VGND 0.01348f
C8548 XThC.XTBN.Y.t42 VGND 0.01024f
C8549 XThC.XTBN.Y.n110 VGND 0.01227f
C8550 XThC.XTBN.Y.n113 VGND 0.11256f
C8551 XThC.XTBN.Y.t30 VGND 0.01024f
C8552 XThC.XTBN.Y.t98 VGND 0.01024f
C8553 XThC.XTBN.Y.n115 VGND 0.01243f
C8554 XThC.XTBN.Y.t103 VGND 0.01024f
C8555 XThC.XTBN.Y.n116 VGND 0.01348f
C8556 XThC.XTBN.Y.n118 VGND 0.01252f
C8557 XThC.XTBN.Y.n121 VGND 0.01348f
C8558 XThC.XTBN.Y.t34 VGND 0.01024f
C8559 XThC.XTBN.Y.n122 VGND 0.01227f
C8560 XThC.XTBN.Y.n125 VGND 0.07521f
C8561 XThC.XTBN.Y.t96 VGND 0.01024f
C8562 XThC.XTBN.Y.t51 VGND 0.01024f
C8563 XThC.XTBN.Y.n127 VGND 0.01243f
C8564 XThC.XTBN.Y.t58 VGND 0.01024f
C8565 XThC.XTBN.Y.n128 VGND 0.01348f
C8566 XThC.XTBN.Y.n130 VGND 0.01252f
C8567 XThC.XTBN.Y.n133 VGND 0.01348f
C8568 XThC.XTBN.Y.t99 VGND 0.01024f
C8569 XThC.XTBN.Y.n134 VGND 0.01227f
C8570 XThC.XTBN.Y.n137 VGND 0.07521f
C8571 XThC.XTBN.Y.t88 VGND 0.01024f
C8572 XThC.XTBN.Y.t37 VGND 0.01024f
C8573 XThC.XTBN.Y.n139 VGND 0.01243f
C8574 XThC.XTBN.Y.t40 VGND 0.01024f
C8575 XThC.XTBN.Y.n140 VGND 0.01348f
C8576 XThC.XTBN.Y.n142 VGND 0.01252f
C8577 XThC.XTBN.Y.n145 VGND 0.01348f
C8578 XThC.XTBN.Y.t91 VGND 0.01024f
C8579 XThC.XTBN.Y.n146 VGND 0.01227f
C8580 XThC.XTBN.Y.n149 VGND 0.07534f
C8581 XThC.XTBN.Y.t7 VGND 0.01024f
C8582 XThC.XTBN.Y.t81 VGND 0.01024f
C8583 XThC.XTBN.Y.n151 VGND 0.01243f
C8584 XThC.XTBN.Y.t86 VGND 0.01024f
C8585 XThC.XTBN.Y.n152 VGND 0.01348f
C8586 XThC.XTBN.Y.n154 VGND 0.01252f
C8587 XThC.XTBN.Y.n157 VGND 0.01348f
C8588 XThC.XTBN.Y.t13 VGND 0.01024f
C8589 XThC.XTBN.Y.n158 VGND 0.01227f
C8590 XThC.XTBN.Y.n161 VGND 0.07521f
C8591 XThC.XTBN.Y.t23 VGND 0.01024f
C8592 XThC.XTBN.Y.t95 VGND 0.01024f
C8593 XThC.XTBN.Y.n163 VGND 0.01243f
C8594 XThC.XTBN.Y.t97 VGND 0.01024f
C8595 XThC.XTBN.Y.n164 VGND 0.01348f
C8596 XThC.XTBN.Y.n166 VGND 0.01252f
C8597 XThC.XTBN.Y.n169 VGND 0.01348f
C8598 XThC.XTBN.Y.t28 VGND 0.01024f
C8599 XThC.XTBN.Y.n170 VGND 0.01227f
C8600 XThC.XTBN.Y.n173 VGND 0.08751f
C8601 XThC.XTBN.Y.n174 VGND 0.11019f
C8602 XThC.XTBN.Y.t75 VGND 0.01024f
C8603 XThC.XTBN.Y.t33 VGND 0.01024f
C8604 XThC.XTBN.Y.n175 VGND 0.01477f
C8605 XThC.XTBN.Y.t27 VGND 0.01024f
C8606 XThC.XTBN.Y.n176 VGND 0.02293f
C8607 XThC.XTBN.Y.n181 VGND 0.01477f
C8608 XThC.XTBN.Y.t9 VGND 0.01024f
C8609 XThC.XTBN.Y.n182 VGND 0.0138f
C8610 XThC.XTBN.Y.n186 VGND 0.11129f
C8611 XThC.XTBN.Y.n187 VGND 0.02169f
C8612 XThC.XTBN.Y.n188 VGND 0.01513f
C8613 XThC.XTBN.Y.n189 VGND 0.0307f
C8614 XThR.Tn[12].t11 VGND 0.01931f
C8615 XThR.Tn[12].t9 VGND 0.01931f
C8616 XThR.Tn[12].n0 VGND 0.05864f
C8617 XThR.Tn[12].t8 VGND 0.01931f
C8618 XThR.Tn[12].t10 VGND 0.01931f
C8619 XThR.Tn[12].n1 VGND 0.04293f
C8620 XThR.Tn[12].n2 VGND 0.1952f
C8621 XThR.Tn[12].t6 VGND 0.01931f
C8622 XThR.Tn[12].t4 VGND 0.01931f
C8623 XThR.Tn[12].n3 VGND 0.04172f
C8624 XThR.Tn[12].t7 VGND 0.01931f
C8625 XThR.Tn[12].t5 VGND 0.01931f
C8626 XThR.Tn[12].n4 VGND 0.06351f
C8627 XThR.Tn[12].n5 VGND 0.17633f
C8628 XThR.Tn[12].t36 VGND 0.01509f
C8629 XThR.Tn[12].t28 VGND 0.01653f
C8630 XThR.Tn[12].n7 VGND 0.04036f
C8631 XThR.Tn[12].n8 VGND 0.07753f
C8632 XThR.Tn[12].t53 VGND 0.01509f
C8633 XThR.Tn[12].t43 VGND 0.01653f
C8634 XThR.Tn[12].n9 VGND 0.04036f
C8635 XThR.Tn[12].t71 VGND 0.01504f
C8636 XThR.Tn[12].t21 VGND 0.01647f
C8637 XThR.Tn[12].n10 VGND 0.04199f
C8638 XThR.Tn[12].n11 VGND 0.0295f
C8639 XThR.Tn[12].n13 VGND 0.09466f
C8640 XThR.Tn[12].t30 VGND 0.01509f
C8641 XThR.Tn[12].t20 VGND 0.01653f
C8642 XThR.Tn[12].n14 VGND 0.04036f
C8643 XThR.Tn[12].t49 VGND 0.01504f
C8644 XThR.Tn[12].t60 VGND 0.01647f
C8645 XThR.Tn[12].n15 VGND 0.04199f
C8646 XThR.Tn[12].n16 VGND 0.0295f
C8647 XThR.Tn[12].n18 VGND 0.09466f
C8648 XThR.Tn[12].t45 VGND 0.01509f
C8649 XThR.Tn[12].t38 VGND 0.01653f
C8650 XThR.Tn[12].n19 VGND 0.04036f
C8651 XThR.Tn[12].t63 VGND 0.01504f
C8652 XThR.Tn[12].t15 VGND 0.01647f
C8653 XThR.Tn[12].n20 VGND 0.04199f
C8654 XThR.Tn[12].n21 VGND 0.0295f
C8655 XThR.Tn[12].n23 VGND 0.09466f
C8656 XThR.Tn[12].t70 VGND 0.01509f
C8657 XThR.Tn[12].t66 VGND 0.01653f
C8658 XThR.Tn[12].n24 VGND 0.04036f
C8659 XThR.Tn[12].t33 VGND 0.01504f
C8660 XThR.Tn[12].t46 VGND 0.01647f
C8661 XThR.Tn[12].n25 VGND 0.04199f
C8662 XThR.Tn[12].n26 VGND 0.0295f
C8663 XThR.Tn[12].n28 VGND 0.09466f
C8664 XThR.Tn[12].t48 VGND 0.01509f
C8665 XThR.Tn[12].t39 VGND 0.01653f
C8666 XThR.Tn[12].n29 VGND 0.04036f
C8667 XThR.Tn[12].t64 VGND 0.01504f
C8668 XThR.Tn[12].t17 VGND 0.01647f
C8669 XThR.Tn[12].n30 VGND 0.04199f
C8670 XThR.Tn[12].n31 VGND 0.0295f
C8671 XThR.Tn[12].n33 VGND 0.09466f
C8672 XThR.Tn[12].t23 VGND 0.01509f
C8673 XThR.Tn[12].t56 VGND 0.01653f
C8674 XThR.Tn[12].n34 VGND 0.04036f
C8675 XThR.Tn[12].t41 VGND 0.01504f
C8676 XThR.Tn[12].t37 VGND 0.01647f
C8677 XThR.Tn[12].n35 VGND 0.04199f
C8678 XThR.Tn[12].n36 VGND 0.0295f
C8679 XThR.Tn[12].n38 VGND 0.09466f
C8680 XThR.Tn[12].t54 VGND 0.01509f
C8681 XThR.Tn[12].t51 VGND 0.01653f
C8682 XThR.Tn[12].n39 VGND 0.04036f
C8683 XThR.Tn[12].t72 VGND 0.01504f
C8684 XThR.Tn[12].t29 VGND 0.01647f
C8685 XThR.Tn[12].n40 VGND 0.04199f
C8686 XThR.Tn[12].n41 VGND 0.0295f
C8687 XThR.Tn[12].n43 VGND 0.09466f
C8688 XThR.Tn[12].t59 VGND 0.01509f
C8689 XThR.Tn[12].t65 VGND 0.01653f
C8690 XThR.Tn[12].n44 VGND 0.04036f
C8691 XThR.Tn[12].t14 VGND 0.01504f
C8692 XThR.Tn[12].t44 VGND 0.01647f
C8693 XThR.Tn[12].n45 VGND 0.04199f
C8694 XThR.Tn[12].n46 VGND 0.0295f
C8695 XThR.Tn[12].n48 VGND 0.09466f
C8696 XThR.Tn[12].t12 VGND 0.01509f
C8697 XThR.Tn[12].t22 VGND 0.01653f
C8698 XThR.Tn[12].n49 VGND 0.04036f
C8699 XThR.Tn[12].t35 VGND 0.01504f
C8700 XThR.Tn[12].t61 VGND 0.01647f
C8701 XThR.Tn[12].n50 VGND 0.04199f
C8702 XThR.Tn[12].n51 VGND 0.0295f
C8703 XThR.Tn[12].n53 VGND 0.09466f
C8704 XThR.Tn[12].t68 VGND 0.01509f
C8705 XThR.Tn[12].t40 VGND 0.01653f
C8706 XThR.Tn[12].n54 VGND 0.04036f
C8707 XThR.Tn[12].t26 VGND 0.01504f
C8708 XThR.Tn[12].t19 VGND 0.01647f
C8709 XThR.Tn[12].n55 VGND 0.04199f
C8710 XThR.Tn[12].n56 VGND 0.0295f
C8711 XThR.Tn[12].n58 VGND 0.09466f
C8712 XThR.Tn[12].t25 VGND 0.01509f
C8713 XThR.Tn[12].t16 VGND 0.01653f
C8714 XThR.Tn[12].n59 VGND 0.04036f
C8715 XThR.Tn[12].t42 VGND 0.01504f
C8716 XThR.Tn[12].t55 VGND 0.01647f
C8717 XThR.Tn[12].n60 VGND 0.04199f
C8718 XThR.Tn[12].n61 VGND 0.0295f
C8719 XThR.Tn[12].n63 VGND 0.09466f
C8720 XThR.Tn[12].t57 VGND 0.01509f
C8721 XThR.Tn[12].t52 VGND 0.01653f
C8722 XThR.Tn[12].n64 VGND 0.04036f
C8723 XThR.Tn[12].t13 VGND 0.01504f
C8724 XThR.Tn[12].t31 VGND 0.01647f
C8725 XThR.Tn[12].n65 VGND 0.04199f
C8726 XThR.Tn[12].n66 VGND 0.0295f
C8727 XThR.Tn[12].n68 VGND 0.09466f
C8728 XThR.Tn[12].t73 VGND 0.01509f
C8729 XThR.Tn[12].t67 VGND 0.01653f
C8730 XThR.Tn[12].n69 VGND 0.04036f
C8731 XThR.Tn[12].t34 VGND 0.01504f
C8732 XThR.Tn[12].t47 VGND 0.01647f
C8733 XThR.Tn[12].n70 VGND 0.04199f
C8734 XThR.Tn[12].n71 VGND 0.0295f
C8735 XThR.Tn[12].n73 VGND 0.09466f
C8736 XThR.Tn[12].t32 VGND 0.01509f
C8737 XThR.Tn[12].t24 VGND 0.01653f
C8738 XThR.Tn[12].n74 VGND 0.04036f
C8739 XThR.Tn[12].t50 VGND 0.01504f
C8740 XThR.Tn[12].t62 VGND 0.01647f
C8741 XThR.Tn[12].n75 VGND 0.04199f
C8742 XThR.Tn[12].n76 VGND 0.0295f
C8743 XThR.Tn[12].n78 VGND 0.09466f
C8744 XThR.Tn[12].t69 VGND 0.01509f
C8745 XThR.Tn[12].t18 VGND 0.01653f
C8746 XThR.Tn[12].n79 VGND 0.04036f
C8747 XThR.Tn[12].t27 VGND 0.01504f
C8748 XThR.Tn[12].t58 VGND 0.01647f
C8749 XThR.Tn[12].n80 VGND 0.04199f
C8750 XThR.Tn[12].n81 VGND 0.0295f
C8751 XThR.Tn[12].n83 VGND 0.09466f
C8752 XThR.Tn[12].n84 VGND 0.08603f
C8753 XThR.Tn[12].n85 VGND 0.29341f
C8754 XThR.Tn[12].t2 VGND 0.01255f
C8755 XThR.Tn[12].t0 VGND 0.01255f
C8756 XThR.Tn[12].n86 VGND 0.0251f
C8757 XThR.Tn[12].t3 VGND 0.01255f
C8758 XThR.Tn[12].t1 VGND 0.01255f
C8759 XThR.Tn[12].n87 VGND 0.03131f
C8760 XThR.Tn[12].n88 VGND 0.05789f
C8761 XThR.Tn[14].t8 VGND 0.0197f
C8762 XThR.Tn[14].t9 VGND 0.0197f
C8763 XThR.Tn[14].n0 VGND 0.0598f
C8764 XThR.Tn[14].t10 VGND 0.0197f
C8765 XThR.Tn[14].t11 VGND 0.0197f
C8766 XThR.Tn[14].n1 VGND 0.04378f
C8767 XThR.Tn[14].n2 VGND 0.19909f
C8768 XThR.Tn[14].t6 VGND 0.0197f
C8769 XThR.Tn[14].t7 VGND 0.0197f
C8770 XThR.Tn[14].n3 VGND 0.04256f
C8771 XThR.Tn[14].t4 VGND 0.0197f
C8772 XThR.Tn[14].t5 VGND 0.0197f
C8773 XThR.Tn[14].n4 VGND 0.06477f
C8774 XThR.Tn[14].n5 VGND 0.17985f
C8775 XThR.Tn[14].t69 VGND 0.01539f
C8776 XThR.Tn[14].t62 VGND 0.01686f
C8777 XThR.Tn[14].n7 VGND 0.04116f
C8778 XThR.Tn[14].n8 VGND 0.07907f
C8779 XThR.Tn[14].t24 VGND 0.01539f
C8780 XThR.Tn[14].t13 VGND 0.01686f
C8781 XThR.Tn[14].n9 VGND 0.04116f
C8782 XThR.Tn[14].t28 VGND 0.01534f
C8783 XThR.Tn[14].t60 VGND 0.0168f
C8784 XThR.Tn[14].n10 VGND 0.04283f
C8785 XThR.Tn[14].n11 VGND 0.03009f
C8786 XThR.Tn[14].n13 VGND 0.09655f
C8787 XThR.Tn[14].t64 VGND 0.01539f
C8788 XThR.Tn[14].t54 VGND 0.01686f
C8789 XThR.Tn[14].n14 VGND 0.04116f
C8790 XThR.Tn[14].t67 VGND 0.01534f
C8791 XThR.Tn[14].t34 VGND 0.0168f
C8792 XThR.Tn[14].n15 VGND 0.04283f
C8793 XThR.Tn[14].n16 VGND 0.03009f
C8794 XThR.Tn[14].n18 VGND 0.09655f
C8795 XThR.Tn[14].t14 VGND 0.01539f
C8796 XThR.Tn[14].t72 VGND 0.01686f
C8797 XThR.Tn[14].n19 VGND 0.04116f
C8798 XThR.Tn[14].t17 VGND 0.01534f
C8799 XThR.Tn[14].t52 VGND 0.0168f
C8800 XThR.Tn[14].n20 VGND 0.04283f
C8801 XThR.Tn[14].n21 VGND 0.03009f
C8802 XThR.Tn[14].n23 VGND 0.09655f
C8803 XThR.Tn[14].t44 VGND 0.01539f
C8804 XThR.Tn[14].t38 VGND 0.01686f
C8805 XThR.Tn[14].n24 VGND 0.04116f
C8806 XThR.Tn[14].t47 VGND 0.01534f
C8807 XThR.Tn[14].t18 VGND 0.0168f
C8808 XThR.Tn[14].n25 VGND 0.04283f
C8809 XThR.Tn[14].n26 VGND 0.03009f
C8810 XThR.Tn[14].n28 VGND 0.09655f
C8811 XThR.Tn[14].t15 VGND 0.01539f
C8812 XThR.Tn[14].t73 VGND 0.01686f
C8813 XThR.Tn[14].n29 VGND 0.04116f
C8814 XThR.Tn[14].t21 VGND 0.01534f
C8815 XThR.Tn[14].t53 VGND 0.0168f
C8816 XThR.Tn[14].n30 VGND 0.04283f
C8817 XThR.Tn[14].n31 VGND 0.03009f
C8818 XThR.Tn[14].n33 VGND 0.09655f
C8819 XThR.Tn[14].t57 VGND 0.01539f
C8820 XThR.Tn[14].t25 VGND 0.01686f
C8821 XThR.Tn[14].n34 VGND 0.04116f
C8822 XThR.Tn[14].t61 VGND 0.01534f
C8823 XThR.Tn[14].t71 VGND 0.0168f
C8824 XThR.Tn[14].n35 VGND 0.04283f
C8825 XThR.Tn[14].n36 VGND 0.03009f
C8826 XThR.Tn[14].n38 VGND 0.09655f
C8827 XThR.Tn[14].t23 VGND 0.01539f
C8828 XThR.Tn[14].t19 VGND 0.01686f
C8829 XThR.Tn[14].n39 VGND 0.04116f
C8830 XThR.Tn[14].t29 VGND 0.01534f
C8831 XThR.Tn[14].t66 VGND 0.0168f
C8832 XThR.Tn[14].n40 VGND 0.04283f
C8833 XThR.Tn[14].n41 VGND 0.03009f
C8834 XThR.Tn[14].n43 VGND 0.09655f
C8835 XThR.Tn[14].t27 VGND 0.01539f
C8836 XThR.Tn[14].t36 VGND 0.01686f
C8837 XThR.Tn[14].n44 VGND 0.04116f
C8838 XThR.Tn[14].t33 VGND 0.01534f
C8839 XThR.Tn[14].t16 VGND 0.0168f
C8840 XThR.Tn[14].n45 VGND 0.04283f
C8841 XThR.Tn[14].n46 VGND 0.03009f
C8842 XThR.Tn[14].n48 VGND 0.09655f
C8843 XThR.Tn[14].t46 VGND 0.01539f
C8844 XThR.Tn[14].t56 VGND 0.01686f
C8845 XThR.Tn[14].n49 VGND 0.04116f
C8846 XThR.Tn[14].t50 VGND 0.01534f
C8847 XThR.Tn[14].t35 VGND 0.0168f
C8848 XThR.Tn[14].n50 VGND 0.04283f
C8849 XThR.Tn[14].n51 VGND 0.03009f
C8850 XThR.Tn[14].n53 VGND 0.09655f
C8851 XThR.Tn[14].t40 VGND 0.01539f
C8852 XThR.Tn[14].t12 VGND 0.01686f
C8853 XThR.Tn[14].n54 VGND 0.04116f
C8854 XThR.Tn[14].t42 VGND 0.01534f
C8855 XThR.Tn[14].t55 VGND 0.0168f
C8856 XThR.Tn[14].n55 VGND 0.04283f
C8857 XThR.Tn[14].n56 VGND 0.03009f
C8858 XThR.Tn[14].n58 VGND 0.09655f
C8859 XThR.Tn[14].t59 VGND 0.01539f
C8860 XThR.Tn[14].t49 VGND 0.01686f
C8861 XThR.Tn[14].n59 VGND 0.04116f
C8862 XThR.Tn[14].t63 VGND 0.01534f
C8863 XThR.Tn[14].t30 VGND 0.0168f
C8864 XThR.Tn[14].n60 VGND 0.04283f
C8865 XThR.Tn[14].n61 VGND 0.03009f
C8866 XThR.Tn[14].n63 VGND 0.09655f
C8867 XThR.Tn[14].t26 VGND 0.01539f
C8868 XThR.Tn[14].t22 VGND 0.01686f
C8869 XThR.Tn[14].n64 VGND 0.04116f
C8870 XThR.Tn[14].t31 VGND 0.01534f
C8871 XThR.Tn[14].t68 VGND 0.0168f
C8872 XThR.Tn[14].n65 VGND 0.04283f
C8873 XThR.Tn[14].n66 VGND 0.03009f
C8874 XThR.Tn[14].n68 VGND 0.09655f
C8875 XThR.Tn[14].t45 VGND 0.01539f
C8876 XThR.Tn[14].t39 VGND 0.01686f
C8877 XThR.Tn[14].n69 VGND 0.04116f
C8878 XThR.Tn[14].t48 VGND 0.01534f
C8879 XThR.Tn[14].t20 VGND 0.0168f
C8880 XThR.Tn[14].n70 VGND 0.04283f
C8881 XThR.Tn[14].n71 VGND 0.03009f
C8882 XThR.Tn[14].n73 VGND 0.09655f
C8883 XThR.Tn[14].t65 VGND 0.01539f
C8884 XThR.Tn[14].t58 VGND 0.01686f
C8885 XThR.Tn[14].n74 VGND 0.04116f
C8886 XThR.Tn[14].t70 VGND 0.01534f
C8887 XThR.Tn[14].t37 VGND 0.0168f
C8888 XThR.Tn[14].n75 VGND 0.04283f
C8889 XThR.Tn[14].n76 VGND 0.03009f
C8890 XThR.Tn[14].n78 VGND 0.09655f
C8891 XThR.Tn[14].t41 VGND 0.01539f
C8892 XThR.Tn[14].t51 VGND 0.01686f
C8893 XThR.Tn[14].n79 VGND 0.04116f
C8894 XThR.Tn[14].t43 VGND 0.01534f
C8895 XThR.Tn[14].t32 VGND 0.0168f
C8896 XThR.Tn[14].n80 VGND 0.04283f
C8897 XThR.Tn[14].n81 VGND 0.03009f
C8898 XThR.Tn[14].n83 VGND 0.09655f
C8899 XThR.Tn[14].n84 VGND 0.08774f
C8900 XThR.Tn[14].n85 VGND 0.35247f
C8901 XThR.Tn[14].t0 VGND 0.0128f
C8902 XThR.Tn[14].t1 VGND 0.0128f
C8903 XThR.Tn[14].n86 VGND 0.02561f
C8904 XThR.Tn[14].t2 VGND 0.0128f
C8905 XThR.Tn[14].t3 VGND 0.0128f
C8906 XThR.Tn[14].n87 VGND 0.03193f
C8907 XThR.Tn[14].n88 VGND 0.05904f
C8908 XThR.Tn[6].t7 VGND 0.01813f
C8909 XThR.Tn[6].t4 VGND 0.01813f
C8910 XThR.Tn[6].n0 VGND 0.0366f
C8911 XThR.Tn[6].t6 VGND 0.01813f
C8912 XThR.Tn[6].t5 VGND 0.01813f
C8913 XThR.Tn[6].n1 VGND 0.04282f
C8914 XThR.Tn[6].n2 VGND 0.12845f
C8915 XThR.Tn[6].t8 VGND 0.01179f
C8916 XThR.Tn[6].t9 VGND 0.01179f
C8917 XThR.Tn[6].n3 VGND 0.02684f
C8918 XThR.Tn[6].t11 VGND 0.01179f
C8919 XThR.Tn[6].t10 VGND 0.01179f
C8920 XThR.Tn[6].n4 VGND 0.02684f
C8921 XThR.Tn[6].t0 VGND 0.01179f
C8922 XThR.Tn[6].t1 VGND 0.01179f
C8923 XThR.Tn[6].n5 VGND 0.04472f
C8924 XThR.Tn[6].t3 VGND 0.01179f
C8925 XThR.Tn[6].t2 VGND 0.01179f
C8926 XThR.Tn[6].n6 VGND 0.02684f
C8927 XThR.Tn[6].n7 VGND 0.12781f
C8928 XThR.Tn[6].n8 VGND 0.07901f
C8929 XThR.Tn[6].n9 VGND 0.08917f
C8930 XThR.Tn[6].t62 VGND 0.01417f
C8931 XThR.Tn[6].t56 VGND 0.01552f
C8932 XThR.Tn[6].n10 VGND 0.03789f
C8933 XThR.Tn[6].n11 VGND 0.07279f
C8934 XThR.Tn[6].t20 VGND 0.01417f
C8935 XThR.Tn[6].t72 VGND 0.01552f
C8936 XThR.Tn[6].n12 VGND 0.03789f
C8937 XThR.Tn[6].t36 VGND 0.01412f
C8938 XThR.Tn[6].t68 VGND 0.01547f
C8939 XThR.Tn[6].n13 VGND 0.03943f
C8940 XThR.Tn[6].n14 VGND 0.0277f
C8941 XThR.Tn[6].n16 VGND 0.08888f
C8942 XThR.Tn[6].t57 VGND 0.01417f
C8943 XThR.Tn[6].t49 VGND 0.01552f
C8944 XThR.Tn[6].n17 VGND 0.03789f
C8945 XThR.Tn[6].t14 VGND 0.01412f
C8946 XThR.Tn[6].t45 VGND 0.01547f
C8947 XThR.Tn[6].n18 VGND 0.03943f
C8948 XThR.Tn[6].n19 VGND 0.0277f
C8949 XThR.Tn[6].n21 VGND 0.08888f
C8950 XThR.Tn[6].t73 VGND 0.01417f
C8951 XThR.Tn[6].t66 VGND 0.01552f
C8952 XThR.Tn[6].n22 VGND 0.03789f
C8953 XThR.Tn[6].t26 VGND 0.01412f
C8954 XThR.Tn[6].t63 VGND 0.01547f
C8955 XThR.Tn[6].n23 VGND 0.03943f
C8956 XThR.Tn[6].n24 VGND 0.0277f
C8957 XThR.Tn[6].n26 VGND 0.08888f
C8958 XThR.Tn[6].t35 VGND 0.01417f
C8959 XThR.Tn[6].t31 VGND 0.01552f
C8960 XThR.Tn[6].n27 VGND 0.03789f
C8961 XThR.Tn[6].t59 VGND 0.01412f
C8962 XThR.Tn[6].t27 VGND 0.01547f
C8963 XThR.Tn[6].n28 VGND 0.03943f
C8964 XThR.Tn[6].n29 VGND 0.0277f
C8965 XThR.Tn[6].n31 VGND 0.08888f
C8966 XThR.Tn[6].t13 VGND 0.01417f
C8967 XThR.Tn[6].t67 VGND 0.01552f
C8968 XThR.Tn[6].n32 VGND 0.03789f
C8969 XThR.Tn[6].t29 VGND 0.01412f
C8970 XThR.Tn[6].t64 VGND 0.01547f
C8971 XThR.Tn[6].n33 VGND 0.03943f
C8972 XThR.Tn[6].n34 VGND 0.0277f
C8973 XThR.Tn[6].n36 VGND 0.08888f
C8974 XThR.Tn[6].t51 VGND 0.01417f
C8975 XThR.Tn[6].t22 VGND 0.01552f
C8976 XThR.Tn[6].n37 VGND 0.03789f
C8977 XThR.Tn[6].t70 VGND 0.01412f
C8978 XThR.Tn[6].t19 VGND 0.01547f
C8979 XThR.Tn[6].n38 VGND 0.03943f
C8980 XThR.Tn[6].n39 VGND 0.0277f
C8981 XThR.Tn[6].n41 VGND 0.08888f
C8982 XThR.Tn[6].t21 VGND 0.01417f
C8983 XThR.Tn[6].t17 VGND 0.01552f
C8984 XThR.Tn[6].n42 VGND 0.03789f
C8985 XThR.Tn[6].t37 VGND 0.01412f
C8986 XThR.Tn[6].t12 VGND 0.01547f
C8987 XThR.Tn[6].n43 VGND 0.03943f
C8988 XThR.Tn[6].n44 VGND 0.0277f
C8989 XThR.Tn[6].n46 VGND 0.08888f
C8990 XThR.Tn[6].t24 VGND 0.01417f
C8991 XThR.Tn[6].t30 VGND 0.01552f
C8992 XThR.Tn[6].n47 VGND 0.03789f
C8993 XThR.Tn[6].t43 VGND 0.01412f
C8994 XThR.Tn[6].t25 VGND 0.01547f
C8995 XThR.Tn[6].n48 VGND 0.03943f
C8996 XThR.Tn[6].n49 VGND 0.0277f
C8997 XThR.Tn[6].n51 VGND 0.08888f
C8998 XThR.Tn[6].t40 VGND 0.01417f
C8999 XThR.Tn[6].t50 VGND 0.01552f
C9000 XThR.Tn[6].n52 VGND 0.03789f
C9001 XThR.Tn[6].t61 VGND 0.01412f
C9002 XThR.Tn[6].t47 VGND 0.01547f
C9003 XThR.Tn[6].n53 VGND 0.03943f
C9004 XThR.Tn[6].n54 VGND 0.0277f
C9005 XThR.Tn[6].n56 VGND 0.08888f
C9006 XThR.Tn[6].t33 VGND 0.01417f
C9007 XThR.Tn[6].t69 VGND 0.01552f
C9008 XThR.Tn[6].n57 VGND 0.03789f
C9009 XThR.Tn[6].t54 VGND 0.01412f
C9010 XThR.Tn[6].t65 VGND 0.01547f
C9011 XThR.Tn[6].n58 VGND 0.03943f
C9012 XThR.Tn[6].n59 VGND 0.0277f
C9013 XThR.Tn[6].n61 VGND 0.08888f
C9014 XThR.Tn[6].t53 VGND 0.01417f
C9015 XThR.Tn[6].t44 VGND 0.01552f
C9016 XThR.Tn[6].n62 VGND 0.03789f
C9017 XThR.Tn[6].t71 VGND 0.01412f
C9018 XThR.Tn[6].t39 VGND 0.01547f
C9019 XThR.Tn[6].n63 VGND 0.03943f
C9020 XThR.Tn[6].n64 VGND 0.0277f
C9021 XThR.Tn[6].n66 VGND 0.08888f
C9022 XThR.Tn[6].t23 VGND 0.01417f
C9023 XThR.Tn[6].t18 VGND 0.01552f
C9024 XThR.Tn[6].n67 VGND 0.03789f
C9025 XThR.Tn[6].t41 VGND 0.01412f
C9026 XThR.Tn[6].t15 VGND 0.01547f
C9027 XThR.Tn[6].n68 VGND 0.03943f
C9028 XThR.Tn[6].n69 VGND 0.0277f
C9029 XThR.Tn[6].n71 VGND 0.08888f
C9030 XThR.Tn[6].t38 VGND 0.01417f
C9031 XThR.Tn[6].t32 VGND 0.01552f
C9032 XThR.Tn[6].n72 VGND 0.03789f
C9033 XThR.Tn[6].t60 VGND 0.01412f
C9034 XThR.Tn[6].t28 VGND 0.01547f
C9035 XThR.Tn[6].n73 VGND 0.03943f
C9036 XThR.Tn[6].n74 VGND 0.0277f
C9037 XThR.Tn[6].n76 VGND 0.08888f
C9038 XThR.Tn[6].t58 VGND 0.01417f
C9039 XThR.Tn[6].t52 VGND 0.01552f
C9040 XThR.Tn[6].n77 VGND 0.03789f
C9041 XThR.Tn[6].t16 VGND 0.01412f
C9042 XThR.Tn[6].t48 VGND 0.01547f
C9043 XThR.Tn[6].n78 VGND 0.03943f
C9044 XThR.Tn[6].n79 VGND 0.0277f
C9045 XThR.Tn[6].n81 VGND 0.08888f
C9046 XThR.Tn[6].t34 VGND 0.01417f
C9047 XThR.Tn[6].t46 VGND 0.01552f
C9048 XThR.Tn[6].n82 VGND 0.03789f
C9049 XThR.Tn[6].t55 VGND 0.01412f
C9050 XThR.Tn[6].t42 VGND 0.01547f
C9051 XThR.Tn[6].n83 VGND 0.03943f
C9052 XThR.Tn[6].n84 VGND 0.0277f
C9053 XThR.Tn[6].n86 VGND 0.08888f
C9054 XThR.Tn[6].n87 VGND 0.08078f
C9055 XThR.Tn[6].n88 VGND 0.13446f
C9056 XThR.XTBN.Y.t60 VGND 0.01124f
C9057 XThR.XTBN.Y.n1 VGND 0.01347f
C9058 XThR.XTBN.Y.t12 VGND 0.01124f
C9059 XThR.XTBN.Y.t81 VGND 0.01124f
C9060 XThR.XTBN.Y.n2 VGND 0.01479f
C9061 XThR.XTBN.Y.t121 VGND 0.01124f
C9062 XThR.XTBN.Y.n3 VGND 0.01365f
C9063 XThR.XTBN.Y.n5 VGND 0.01304f
C9064 XThR.XTBN.Y.n8 VGND 0.01479f
C9065 XThR.XTBN.Y.n10 VGND 0.0122f
C9066 XThR.XTBN.Y.t115 VGND 0.01124f
C9067 XThR.XTBN.Y.n12 VGND 0.01347f
C9068 XThR.XTBN.Y.t65 VGND 0.01124f
C9069 XThR.XTBN.Y.t21 VGND 0.01124f
C9070 XThR.XTBN.Y.n13 VGND 0.01479f
C9071 XThR.XTBN.Y.t57 VGND 0.01124f
C9072 XThR.XTBN.Y.n14 VGND 0.01365f
C9073 XThR.XTBN.Y.n16 VGND 0.01304f
C9074 XThR.XTBN.Y.n19 VGND 0.01479f
C9075 XThR.XTBN.Y.n22 VGND 0.12354f
C9076 XThR.XTBN.Y.t27 VGND 0.01124f
C9077 XThR.XTBN.Y.n24 VGND 0.01347f
C9078 XThR.XTBN.Y.t96 VGND 0.01124f
C9079 XThR.XTBN.Y.t46 VGND 0.01124f
C9080 XThR.XTBN.Y.n25 VGND 0.01479f
C9081 XThR.XTBN.Y.t89 VGND 0.01124f
C9082 XThR.XTBN.Y.n26 VGND 0.01365f
C9083 XThR.XTBN.Y.n28 VGND 0.01304f
C9084 XThR.XTBN.Y.n31 VGND 0.01479f
C9085 XThR.XTBN.Y.n34 VGND 0.08255f
C9086 XThR.XTBN.Y.t80 VGND 0.01124f
C9087 XThR.XTBN.Y.n36 VGND 0.01347f
C9088 XThR.XTBN.Y.t31 VGND 0.01124f
C9089 XThR.XTBN.Y.t102 VGND 0.01124f
C9090 XThR.XTBN.Y.n37 VGND 0.01479f
C9091 XThR.XTBN.Y.t25 VGND 0.01124f
C9092 XThR.XTBN.Y.n38 VGND 0.01365f
C9093 XThR.XTBN.Y.n40 VGND 0.01304f
C9094 XThR.XTBN.Y.n43 VGND 0.01479f
C9095 XThR.XTBN.Y.n46 VGND 0.08255f
C9096 XThR.XTBN.Y.t85 VGND 0.01124f
C9097 XThR.XTBN.Y.n48 VGND 0.01347f
C9098 XThR.XTBN.Y.t33 VGND 0.01124f
C9099 XThR.XTBN.Y.t105 VGND 0.01124f
C9100 XThR.XTBN.Y.n49 VGND 0.01479f
C9101 XThR.XTBN.Y.t26 VGND 0.01124f
C9102 XThR.XTBN.Y.n50 VGND 0.01365f
C9103 XThR.XTBN.Y.n52 VGND 0.01304f
C9104 XThR.XTBN.Y.n55 VGND 0.01479f
C9105 XThR.XTBN.Y.n58 VGND 0.08269f
C9106 XThR.XTBN.Y.t54 VGND 0.01124f
C9107 XThR.XTBN.Y.n60 VGND 0.01347f
C9108 XThR.XTBN.Y.t5 VGND 0.01124f
C9109 XThR.XTBN.Y.t73 VGND 0.01124f
C9110 XThR.XTBN.Y.n61 VGND 0.01479f
C9111 XThR.XTBN.Y.t114 VGND 0.01124f
C9112 XThR.XTBN.Y.n62 VGND 0.01365f
C9113 XThR.XTBN.Y.n64 VGND 0.01304f
C9114 XThR.XTBN.Y.n67 VGND 0.01479f
C9115 XThR.XTBN.Y.n70 VGND 0.08255f
C9116 XThR.XTBN.Y.t49 VGND 0.01124f
C9117 XThR.XTBN.Y.n72 VGND 0.01347f
C9118 XThR.XTBN.Y.t119 VGND 0.01124f
C9119 XThR.XTBN.Y.t69 VGND 0.01124f
C9120 XThR.XTBN.Y.n73 VGND 0.01479f
C9121 XThR.XTBN.Y.t108 VGND 0.01124f
C9122 XThR.XTBN.Y.n74 VGND 0.01365f
C9123 XThR.XTBN.Y.n76 VGND 0.01304f
C9124 XThR.XTBN.Y.n79 VGND 0.01479f
C9125 XThR.XTBN.Y.n82 VGND 0.09424f
C9126 XThR.XTBN.Y.t99 VGND 0.01124f
C9127 XThR.XTBN.Y.t87 VGND 0.01124f
C9128 XThR.XTBN.Y.n83 VGND 0.01621f
C9129 XThR.XTBN.Y.t77 VGND 0.01124f
C9130 XThR.XTBN.Y.t68 VGND 0.01124f
C9131 XThR.XTBN.Y.n84 VGND 0.01515f
C9132 XThR.XTBN.Y.n87 VGND 0.01621f
C9133 XThR.XTBN.Y.n92 VGND 0.02375f
C9134 XThR.XTBN.Y.n93 VGND 0.01318f
C9135 XThR.XTBN.Y.t66 VGND 0.01124f
C9136 XThR.XTBN.Y.t23 VGND 0.01124f
C9137 XThR.XTBN.Y.n94 VGND 0.01621f
C9138 XThR.XTBN.Y.t59 VGND 0.01124f
C9139 XThR.XTBN.Y.t97 VGND 0.01124f
C9140 XThR.XTBN.Y.n95 VGND 0.01515f
C9141 XThR.XTBN.Y.n98 VGND 0.01621f
C9142 XThR.XTBN.Y.n103 VGND 0.02375f
C9143 XThR.XTBN.Y.n105 VGND 0.13142f
C9144 XThR.XTBN.Y.t15 VGND 0.01124f
C9145 XThR.XTBN.Y.t83 VGND 0.01124f
C9146 XThR.XTBN.Y.n106 VGND 0.01621f
C9147 XThR.XTBN.Y.t123 VGND 0.01124f
C9148 XThR.XTBN.Y.t39 VGND 0.01124f
C9149 XThR.XTBN.Y.n107 VGND 0.01515f
C9150 XThR.XTBN.Y.n110 VGND 0.01621f
C9151 XThR.XTBN.Y.n115 VGND 0.02375f
C9152 XThR.XTBN.Y.n117 VGND 0.08248f
C9153 XThR.XTBN.Y.t100 VGND 0.01124f
C9154 XThR.XTBN.Y.t50 VGND 0.01124f
C9155 XThR.XTBN.Y.n118 VGND 0.01621f
C9156 XThR.XTBN.Y.t92 VGND 0.01124f
C9157 XThR.XTBN.Y.t13 VGND 0.01124f
C9158 XThR.XTBN.Y.n119 VGND 0.01515f
C9159 XThR.XTBN.Y.n122 VGND 0.01621f
C9160 XThR.XTBN.Y.n127 VGND 0.02375f
C9161 XThR.XTBN.Y.n129 VGND 0.08248f
C9162 XThR.XTBN.Y.t45 VGND 0.01124f
C9163 XThR.XTBN.Y.t117 VGND 0.01124f
C9164 XThR.XTBN.Y.n130 VGND 0.01621f
C9165 XThR.XTBN.Y.t36 VGND 0.01124f
C9166 XThR.XTBN.Y.t75 VGND 0.01124f
C9167 XThR.XTBN.Y.n131 VGND 0.01515f
C9168 XThR.XTBN.Y.n134 VGND 0.01621f
C9169 XThR.XTBN.Y.n139 VGND 0.02375f
C9170 XThR.XTBN.Y.n141 VGND 0.08248f
C9171 XThR.XTBN.Y.t19 VGND 0.01124f
C9172 XThR.XTBN.Y.t86 VGND 0.01124f
C9173 XThR.XTBN.Y.n142 VGND 0.01621f
C9174 XThR.XTBN.Y.t6 VGND 0.01124f
C9175 XThR.XTBN.Y.t43 VGND 0.01124f
C9176 XThR.XTBN.Y.n143 VGND 0.01515f
C9177 XThR.XTBN.Y.n146 VGND 0.01621f
C9178 XThR.XTBN.Y.n151 VGND 0.02375f
C9179 XThR.XTBN.Y.n153 VGND 0.08248f
C9180 XThR.XTBN.Y.t41 VGND 0.01124f
C9181 XThR.XTBN.Y.t113 VGND 0.01124f
C9182 XThR.XTBN.Y.n154 VGND 0.01621f
C9183 XThR.XTBN.Y.t34 VGND 0.01124f
C9184 XThR.XTBN.Y.t72 VGND 0.01124f
C9185 XThR.XTBN.Y.n155 VGND 0.01515f
C9186 XThR.XTBN.Y.n158 VGND 0.01621f
C9187 XThR.XTBN.Y.n163 VGND 0.02375f
C9188 XThR.XTBN.Y.n165 VGND 0.07589f
C9189 XThR.XTBN.Y.n166 VGND 0.12019f
C9190 XThR.XTBN.Y.t106 VGND 0.01124f
C9191 XThR.XTBN.Y.t63 VGND 0.01124f
C9192 XThR.XTBN.Y.n167 VGND 0.01515f
C9193 XThR.XTBN.Y.n169 VGND 0.01621f
C9194 XThR.XTBN.Y.t56 VGND 0.01124f
C9195 XThR.XTBN.Y.t7 VGND 0.01124f
C9196 XThR.XTBN.Y.n170 VGND 0.02517f
C9197 XThR.XTBN.Y.n174 VGND 0.01621f
C9198 XThR.XTBN.Y.n178 VGND 0.12255f
C9199 XThR.XTBN.Y.n179 VGND 0.02242f
C9200 XThR.XTBN.Y.n180 VGND 0.01587f
C9201 XThR.XTBN.Y.n183 VGND 0.0112f
C9202 XThR.XTBN.Y.n184 VGND 0.022f
C9203 XThC.Tn[10].n0 VGND 0.02345f
C9204 XThC.Tn[10].n1 VGND 0.0188f
C9205 XThC.Tn[10].n2 VGND 0.0473f
C9206 XThC.Tn[10].t38 VGND 0.01146f
C9207 XThC.Tn[10].t36 VGND 0.01252f
C9208 XThC.Tn[10].n3 VGND 0.02796f
C9209 XThC.Tn[10].n4 VGND 0.01598f
C9210 XThC.Tn[10].n5 VGND 0.01943f
C9211 XThC.Tn[10].t24 VGND 0.01146f
C9212 XThC.Tn[10].t21 VGND 0.01252f
C9213 XThC.Tn[10].n6 VGND 0.02796f
C9214 XThC.Tn[10].n7 VGND 0.01598f
C9215 XThC.Tn[10].n8 VGND 0.09232f
C9216 XThC.Tn[10].t29 VGND 0.01146f
C9217 XThC.Tn[10].t23 VGND 0.01252f
C9218 XThC.Tn[10].n9 VGND 0.02796f
C9219 XThC.Tn[10].n10 VGND 0.01598f
C9220 XThC.Tn[10].n11 VGND 0.09232f
C9221 XThC.Tn[10].t30 VGND 0.01146f
C9222 XThC.Tn[10].t25 VGND 0.01252f
C9223 XThC.Tn[10].n12 VGND 0.02796f
C9224 XThC.Tn[10].n13 VGND 0.01598f
C9225 XThC.Tn[10].n14 VGND 0.09232f
C9226 XThC.Tn[10].t17 VGND 0.01146f
C9227 XThC.Tn[10].t14 VGND 0.01252f
C9228 XThC.Tn[10].n15 VGND 0.02796f
C9229 XThC.Tn[10].n16 VGND 0.01598f
C9230 XThC.Tn[10].n17 VGND 0.09232f
C9231 XThC.Tn[10].t18 VGND 0.01146f
C9232 XThC.Tn[10].t15 VGND 0.01252f
C9233 XThC.Tn[10].n18 VGND 0.02796f
C9234 XThC.Tn[10].n19 VGND 0.01598f
C9235 XThC.Tn[10].n20 VGND 0.09232f
C9236 XThC.Tn[10].t34 VGND 0.01146f
C9237 XThC.Tn[10].t28 VGND 0.01252f
C9238 XThC.Tn[10].n21 VGND 0.02796f
C9239 XThC.Tn[10].n22 VGND 0.01598f
C9240 XThC.Tn[10].n23 VGND 0.09232f
C9241 XThC.Tn[10].t41 VGND 0.01146f
C9242 XThC.Tn[10].t37 VGND 0.01252f
C9243 XThC.Tn[10].n24 VGND 0.02796f
C9244 XThC.Tn[10].n25 VGND 0.01598f
C9245 XThC.Tn[10].n26 VGND 0.09232f
C9246 XThC.Tn[10].t43 VGND 0.01146f
C9247 XThC.Tn[10].t39 VGND 0.01252f
C9248 XThC.Tn[10].n27 VGND 0.02796f
C9249 XThC.Tn[10].n28 VGND 0.01598f
C9250 XThC.Tn[10].n29 VGND 0.09232f
C9251 XThC.Tn[10].t31 VGND 0.01146f
C9252 XThC.Tn[10].t26 VGND 0.01252f
C9253 XThC.Tn[10].n30 VGND 0.02796f
C9254 XThC.Tn[10].n31 VGND 0.01598f
C9255 XThC.Tn[10].n32 VGND 0.09232f
C9256 XThC.Tn[10].t33 VGND 0.01146f
C9257 XThC.Tn[10].t27 VGND 0.01252f
C9258 XThC.Tn[10].n33 VGND 0.02796f
C9259 XThC.Tn[10].n34 VGND 0.01598f
C9260 XThC.Tn[10].n35 VGND 0.09232f
C9261 XThC.Tn[10].t12 VGND 0.01146f
C9262 XThC.Tn[10].t40 VGND 0.01252f
C9263 XThC.Tn[10].n36 VGND 0.02796f
C9264 XThC.Tn[10].n37 VGND 0.01598f
C9265 XThC.Tn[10].n38 VGND 0.09232f
C9266 XThC.Tn[10].t20 VGND 0.01146f
C9267 XThC.Tn[10].t16 VGND 0.01252f
C9268 XThC.Tn[10].n39 VGND 0.02796f
C9269 XThC.Tn[10].n40 VGND 0.01598f
C9270 XThC.Tn[10].n41 VGND 0.09232f
C9271 XThC.Tn[10].t22 VGND 0.01146f
C9272 XThC.Tn[10].t19 VGND 0.01252f
C9273 XThC.Tn[10].n42 VGND 0.02796f
C9274 XThC.Tn[10].n43 VGND 0.01598f
C9275 XThC.Tn[10].n44 VGND 0.09232f
C9276 XThC.Tn[10].t35 VGND 0.01146f
C9277 XThC.Tn[10].t32 VGND 0.01252f
C9278 XThC.Tn[10].n45 VGND 0.02796f
C9279 XThC.Tn[10].n46 VGND 0.01598f
C9280 XThC.Tn[10].n47 VGND 0.09232f
C9281 XThC.Tn[10].t13 VGND 0.01146f
C9282 XThC.Tn[10].t42 VGND 0.01252f
C9283 XThC.Tn[10].n48 VGND 0.02796f
C9284 XThC.Tn[10].n49 VGND 0.01598f
C9285 XThC.Tn[10].n50 VGND 0.09232f
C9286 XThC.Tn[10].n51 VGND 0.46113f
C9287 XThC.Tn[10].n52 VGND 0.03515f
C9288 XThC.Tn[10].t2 VGND 0.01446f
C9289 XThC.Tn[10].t1 VGND 0.01446f
C9290 XThC.Tn[10].n53 VGND 0.03125f
C9291 XThC.Tn[10].t5 VGND 0.01446f
C9292 XThC.Tn[10].t9 VGND 0.01446f
C9293 XThC.Tn[10].n54 VGND 0.04756f
C9294 XThC.Tn[10].n55 VGND 0.13215f
C9295 XThC.Tn[10].n56 VGND 0.02078f
C9296 XThC.Tn[10].t7 VGND 0.01446f
C9297 XThC.Tn[10].t8 VGND 0.01446f
C9298 XThC.Tn[10].n57 VGND 0.03215f
C9299 XThC.Tn[10].t0 VGND 0.01446f
C9300 XThC.Tn[10].t4 VGND 0.01446f
C9301 XThC.Tn[10].n58 VGND 0.04391f
C9302 XThC.Tn[10].n59 VGND 0.14309f
C9303 Iout.n0 VGND 0.22972f
C9304 Iout.n1 VGND 1.20114f
C9305 Iout.n2 VGND 0.22972f
C9306 Iout.n3 VGND 0.22972f
C9307 Iout.t234 VGND 0.02212f
C9308 Iout.n4 VGND 0.04919f
C9309 Iout.n5 VGND 0.19431f
C9310 Iout.n6 VGND 0.22972f
C9311 Iout.n7 VGND 1.20114f
C9312 Iout.n8 VGND 0.22972f
C9313 Iout.t75 VGND 0.02212f
C9314 Iout.n9 VGND 0.04919f
C9315 Iout.n10 VGND 0.19431f
C9316 Iout.n11 VGND 0.22972f
C9317 Iout.n12 VGND 1.20114f
C9318 Iout.n13 VGND 0.22972f
C9319 Iout.t32 VGND 0.02212f
C9320 Iout.n14 VGND 0.04919f
C9321 Iout.n15 VGND 0.19431f
C9322 Iout.n16 VGND 0.22972f
C9323 Iout.n17 VGND 1.20114f
C9324 Iout.n18 VGND 0.22972f
C9325 Iout.t10 VGND 0.02212f
C9326 Iout.n19 VGND 0.04919f
C9327 Iout.n20 VGND 0.19431f
C9328 Iout.n21 VGND 0.47625f
C9329 Iout.t79 VGND 0.02212f
C9330 Iout.n22 VGND 0.04919f
C9331 Iout.n23 VGND 0.28657f
C9332 Iout.n24 VGND 0.22972f
C9333 Iout.n25 VGND 0.22972f
C9334 Iout.n26 VGND 0.22972f
C9335 Iout.n27 VGND 0.22972f
C9336 Iout.n28 VGND 0.22972f
C9337 Iout.n29 VGND 0.22972f
C9338 Iout.n30 VGND 0.22972f
C9339 Iout.n31 VGND 0.22972f
C9340 Iout.n32 VGND 0.22972f
C9341 Iout.n33 VGND 0.22972f
C9342 Iout.n34 VGND 0.22972f
C9343 Iout.n35 VGND 0.22972f
C9344 Iout.n36 VGND 0.22972f
C9345 Iout.n37 VGND 0.22972f
C9346 Iout.t44 VGND 0.02212f
C9347 Iout.n38 VGND 0.04919f
C9348 Iout.n39 VGND 0.02502f
C9349 Iout.n40 VGND 0.22972f
C9350 Iout.n41 VGND 0.04584f
C9351 Iout.t184 VGND 0.02212f
C9352 Iout.n42 VGND 0.04919f
C9353 Iout.n43 VGND 0.02502f
C9354 Iout.t201 VGND 0.02212f
C9355 Iout.n44 VGND 0.04919f
C9356 Iout.n45 VGND 0.02502f
C9357 Iout.n46 VGND 0.22972f
C9358 Iout.t94 VGND 0.02212f
C9359 Iout.n47 VGND 0.04919f
C9360 Iout.n48 VGND 0.02502f
C9361 Iout.n49 VGND 0.22972f
C9362 Iout.t200 VGND 0.02212f
C9363 Iout.n50 VGND 0.04919f
C9364 Iout.n51 VGND 0.02502f
C9365 Iout.n52 VGND 0.22972f
C9366 Iout.t120 VGND 0.02212f
C9367 Iout.n53 VGND 0.04919f
C9368 Iout.n54 VGND 0.02502f
C9369 Iout.n55 VGND 0.22972f
C9370 Iout.t69 VGND 0.02212f
C9371 Iout.n56 VGND 0.04919f
C9372 Iout.n57 VGND 0.02502f
C9373 Iout.n58 VGND 0.22972f
C9374 Iout.t24 VGND 0.02212f
C9375 Iout.n59 VGND 0.04919f
C9376 Iout.n60 VGND 0.02502f
C9377 Iout.n61 VGND 0.22972f
C9378 Iout.t92 VGND 0.02212f
C9379 Iout.n62 VGND 0.04919f
C9380 Iout.n63 VGND 0.02502f
C9381 Iout.n64 VGND 0.22972f
C9382 Iout.t61 VGND 0.02212f
C9383 Iout.n65 VGND 0.04919f
C9384 Iout.n66 VGND 0.02502f
C9385 Iout.n67 VGND 0.22972f
C9386 Iout.t85 VGND 0.02212f
C9387 Iout.n68 VGND 0.04919f
C9388 Iout.n69 VGND 0.02502f
C9389 Iout.n70 VGND 0.22972f
C9390 Iout.t112 VGND 0.02212f
C9391 Iout.n71 VGND 0.04919f
C9392 Iout.n72 VGND 0.02502f
C9393 Iout.n73 VGND 0.22972f
C9394 Iout.t136 VGND 0.02212f
C9395 Iout.n74 VGND 0.04919f
C9396 Iout.n75 VGND 0.02502f
C9397 Iout.n76 VGND 0.22972f
C9398 Iout.t110 VGND 0.02212f
C9399 Iout.n77 VGND 0.04919f
C9400 Iout.n78 VGND 0.02502f
C9401 Iout.n79 VGND 0.22972f
C9402 Iout.n80 VGND 0.22972f
C9403 Iout.t131 VGND 0.02212f
C9404 Iout.n81 VGND 0.04919f
C9405 Iout.n82 VGND 0.02502f
C9406 Iout.n83 VGND 0.22972f
C9407 Iout.n84 VGND 0.04584f
C9408 Iout.t50 VGND 0.02212f
C9409 Iout.n85 VGND 0.04919f
C9410 Iout.n86 VGND 0.02502f
C9411 Iout.t52 VGND 0.02212f
C9412 Iout.n87 VGND 0.04919f
C9413 Iout.n88 VGND 0.02502f
C9414 Iout.n89 VGND 0.22972f
C9415 Iout.t20 VGND 0.02212f
C9416 Iout.n90 VGND 0.04919f
C9417 Iout.n91 VGND 0.02502f
C9418 Iout.n92 VGND 0.22972f
C9419 Iout.t173 VGND 0.02212f
C9420 Iout.n93 VGND 0.04919f
C9421 Iout.n94 VGND 0.02502f
C9422 Iout.n95 VGND 0.22972f
C9423 Iout.t253 VGND 0.02212f
C9424 Iout.n96 VGND 0.04919f
C9425 Iout.n97 VGND 0.02502f
C9426 Iout.n98 VGND 0.22972f
C9427 Iout.t132 VGND 0.02212f
C9428 Iout.n99 VGND 0.04919f
C9429 Iout.n100 VGND 0.02502f
C9430 Iout.n101 VGND 0.22972f
C9431 Iout.t93 VGND 0.02212f
C9432 Iout.n102 VGND 0.04919f
C9433 Iout.n103 VGND 0.02502f
C9434 Iout.n104 VGND 0.22972f
C9435 Iout.t203 VGND 0.02212f
C9436 Iout.n105 VGND 0.04919f
C9437 Iout.n106 VGND 0.02502f
C9438 Iout.n107 VGND 0.22972f
C9439 Iout.t211 VGND 0.02212f
C9440 Iout.n108 VGND 0.04919f
C9441 Iout.n109 VGND 0.02502f
C9442 Iout.n110 VGND 0.22972f
C9443 Iout.t250 VGND 0.02212f
C9444 Iout.n111 VGND 0.04919f
C9445 Iout.n112 VGND 0.02502f
C9446 Iout.n113 VGND 0.22972f
C9447 Iout.t175 VGND 0.02212f
C9448 Iout.n114 VGND 0.04919f
C9449 Iout.n115 VGND 0.02502f
C9450 Iout.n116 VGND 0.22972f
C9451 Iout.t34 VGND 0.02212f
C9452 Iout.n117 VGND 0.04919f
C9453 Iout.n118 VGND 0.02502f
C9454 Iout.n119 VGND 0.22972f
C9455 Iout.t6 VGND 0.02212f
C9456 Iout.n120 VGND 0.04919f
C9457 Iout.n121 VGND 0.02502f
C9458 Iout.n122 VGND 0.04584f
C9459 Iout.t168 VGND 0.02212f
C9460 Iout.n123 VGND 0.04919f
C9461 Iout.n124 VGND 0.02502f
C9462 Iout.n125 VGND 0.22972f
C9463 Iout.n126 VGND 0.22972f
C9464 Iout.t101 VGND 0.02212f
C9465 Iout.n127 VGND 0.04919f
C9466 Iout.n128 VGND 0.02502f
C9467 Iout.n129 VGND 0.04584f
C9468 Iout.t225 VGND 0.02212f
C9469 Iout.n130 VGND 0.04919f
C9470 Iout.n131 VGND 0.02502f
C9471 Iout.n132 VGND 0.22972f
C9472 Iout.t84 VGND 0.02212f
C9473 Iout.n133 VGND 0.04919f
C9474 Iout.n134 VGND 0.02502f
C9475 Iout.n135 VGND 0.04584f
C9476 Iout.t214 VGND 0.02212f
C9477 Iout.n136 VGND 0.04919f
C9478 Iout.n137 VGND 0.02502f
C9479 Iout.n138 VGND 0.22972f
C9480 Iout.n139 VGND 0.22972f
C9481 Iout.t185 VGND 0.02212f
C9482 Iout.n140 VGND 0.04919f
C9483 Iout.n141 VGND 0.02502f
C9484 Iout.n142 VGND 0.04584f
C9485 Iout.t0 VGND 0.02212f
C9486 Iout.n143 VGND 0.04919f
C9487 Iout.n144 VGND 0.02502f
C9488 Iout.n145 VGND 0.13561f
C9489 Iout.t125 VGND 0.02212f
C9490 Iout.n146 VGND 0.04919f
C9491 Iout.n147 VGND 0.02502f
C9492 Iout.n148 VGND 0.04584f
C9493 Iout.t7 VGND 0.02212f
C9494 Iout.n149 VGND 0.04919f
C9495 Iout.n150 VGND 0.02502f
C9496 Iout.n151 VGND 0.22972f
C9497 Iout.n152 VGND 0.13561f
C9498 Iout.n153 VGND 0.22972f
C9499 Iout.n154 VGND 0.22972f
C9500 Iout.n155 VGND 0.22972f
C9501 Iout.t40 VGND 0.02212f
C9502 Iout.n156 VGND 0.04919f
C9503 Iout.n157 VGND 0.02502f
C9504 Iout.n158 VGND 0.22972f
C9505 Iout.n159 VGND 0.22972f
C9506 Iout.n160 VGND 0.22972f
C9507 Iout.n161 VGND 0.22972f
C9508 Iout.n162 VGND 0.22972f
C9509 Iout.n163 VGND 0.22972f
C9510 Iout.n164 VGND 0.22972f
C9511 Iout.n165 VGND 0.22972f
C9512 Iout.n166 VGND 0.22972f
C9513 Iout.n167 VGND 0.22972f
C9514 Iout.t189 VGND 0.02212f
C9515 Iout.n168 VGND 0.04919f
C9516 Iout.n169 VGND 0.02502f
C9517 Iout.n170 VGND 0.22972f
C9518 Iout.n171 VGND 0.04584f
C9519 Iout.t91 VGND 0.02212f
C9520 Iout.n172 VGND 0.04919f
C9521 Iout.n173 VGND 0.02502f
C9522 Iout.t248 VGND 0.02212f
C9523 Iout.n174 VGND 0.04919f
C9524 Iout.n175 VGND 0.02502f
C9525 Iout.n176 VGND 0.22972f
C9526 Iout.t12 VGND 0.02212f
C9527 Iout.n177 VGND 0.04919f
C9528 Iout.n178 VGND 0.02502f
C9529 Iout.n179 VGND 0.22972f
C9530 Iout.t13 VGND 0.02212f
C9531 Iout.n180 VGND 0.04919f
C9532 Iout.n181 VGND 0.02502f
C9533 Iout.n182 VGND 0.22972f
C9534 Iout.t230 VGND 0.02212f
C9535 Iout.n183 VGND 0.04919f
C9536 Iout.n184 VGND 0.02502f
C9537 Iout.n185 VGND 0.22972f
C9538 Iout.t29 VGND 0.02212f
C9539 Iout.n186 VGND 0.04919f
C9540 Iout.n187 VGND 0.02502f
C9541 Iout.n188 VGND 0.22972f
C9542 Iout.t118 VGND 0.02212f
C9543 Iout.n189 VGND 0.04919f
C9544 Iout.n190 VGND 0.02502f
C9545 Iout.n191 VGND 0.13561f
C9546 Iout.t167 VGND 0.02212f
C9547 Iout.n192 VGND 0.04919f
C9548 Iout.n193 VGND 0.02502f
C9549 Iout.n194 VGND 0.04584f
C9550 Iout.t197 VGND 0.02212f
C9551 Iout.n195 VGND 0.04919f
C9552 Iout.n196 VGND 0.02502f
C9553 Iout.n197 VGND 0.13561f
C9554 Iout.n198 VGND 0.04584f
C9555 Iout.t233 VGND 0.02212f
C9556 Iout.n199 VGND 0.04919f
C9557 Iout.n200 VGND 0.02502f
C9558 Iout.n201 VGND 0.04584f
C9559 Iout.t18 VGND 0.02212f
C9560 Iout.n202 VGND 0.04919f
C9561 Iout.n203 VGND 0.02502f
C9562 Iout.n204 VGND 0.13561f
C9563 Iout.n205 VGND 0.04584f
C9564 Iout.t193 VGND 0.02212f
C9565 Iout.n206 VGND 0.04919f
C9566 Iout.n207 VGND 0.02502f
C9567 Iout.n208 VGND 0.13561f
C9568 Iout.n209 VGND 0.04584f
C9569 Iout.t89 VGND 0.02212f
C9570 Iout.n210 VGND 0.04919f
C9571 Iout.n211 VGND 0.02502f
C9572 Iout.n212 VGND 0.13561f
C9573 Iout.n213 VGND 0.04584f
C9574 Iout.t78 VGND 0.02212f
C9575 Iout.n214 VGND 0.04919f
C9576 Iout.n215 VGND 0.02502f
C9577 Iout.n216 VGND 0.13561f
C9578 Iout.n217 VGND 0.04584f
C9579 Iout.t161 VGND 0.02212f
C9580 Iout.n218 VGND 0.04919f
C9581 Iout.n219 VGND 0.02502f
C9582 Iout.n220 VGND 0.13561f
C9583 Iout.n221 VGND 0.04584f
C9584 Iout.t181 VGND 0.02212f
C9585 Iout.n222 VGND 0.04919f
C9586 Iout.n223 VGND 0.02502f
C9587 Iout.n224 VGND 0.13561f
C9588 Iout.n225 VGND 0.04584f
C9589 Iout.t48 VGND 0.02212f
C9590 Iout.n226 VGND 0.04919f
C9591 Iout.n227 VGND 0.02502f
C9592 Iout.n228 VGND 0.04584f
C9593 Iout.n229 VGND 0.13561f
C9594 Iout.n230 VGND 0.22972f
C9595 Iout.n231 VGND 0.04584f
C9596 Iout.t133 VGND 0.02212f
C9597 Iout.n232 VGND 0.04919f
C9598 Iout.n233 VGND 0.02502f
C9599 Iout.n234 VGND 0.04584f
C9600 Iout.t126 VGND 0.02212f
C9601 Iout.n235 VGND 0.04919f
C9602 Iout.n236 VGND 0.02502f
C9603 Iout.n237 VGND 0.04584f
C9604 Iout.t3 VGND 0.02212f
C9605 Iout.n238 VGND 0.04919f
C9606 Iout.n239 VGND 0.02502f
C9607 Iout.n240 VGND 0.04584f
C9608 Iout.t2 VGND 0.02212f
C9609 Iout.n241 VGND 0.04919f
C9610 Iout.n242 VGND 0.02502f
C9611 Iout.n243 VGND 0.04584f
C9612 Iout.t255 VGND 0.02212f
C9613 Iout.n244 VGND 0.04919f
C9614 Iout.n245 VGND 0.02502f
C9615 Iout.n246 VGND 0.04584f
C9616 Iout.t8 VGND 0.02212f
C9617 Iout.n247 VGND 0.04919f
C9618 Iout.n248 VGND 0.02502f
C9619 Iout.n249 VGND 0.04584f
C9620 Iout.t245 VGND 0.02212f
C9621 Iout.n250 VGND 0.04919f
C9622 Iout.n251 VGND 0.02502f
C9623 Iout.t212 VGND 0.02212f
C9624 Iout.n252 VGND 0.04919f
C9625 Iout.n253 VGND 0.02502f
C9626 Iout.n254 VGND 0.04584f
C9627 Iout.t21 VGND 0.02212f
C9628 Iout.n255 VGND 0.04919f
C9629 Iout.n256 VGND 0.02502f
C9630 Iout.n257 VGND 0.04584f
C9631 Iout.n258 VGND 0.22972f
C9632 Iout.t227 VGND 0.02212f
C9633 Iout.n259 VGND 0.04919f
C9634 Iout.n260 VGND 0.02502f
C9635 Iout.n261 VGND 0.04584f
C9636 Iout.n262 VGND 0.22972f
C9637 Iout.n263 VGND 0.22972f
C9638 Iout.n264 VGND 0.04584f
C9639 Iout.t229 VGND 0.02212f
C9640 Iout.n265 VGND 0.04919f
C9641 Iout.n266 VGND 0.02502f
C9642 Iout.n267 VGND 0.04584f
C9643 Iout.n268 VGND 0.22972f
C9644 Iout.n269 VGND 0.22972f
C9645 Iout.n270 VGND 0.04584f
C9646 Iout.t81 VGND 0.02212f
C9647 Iout.n271 VGND 0.04919f
C9648 Iout.n272 VGND 0.02502f
C9649 Iout.n273 VGND 0.04584f
C9650 Iout.n274 VGND 0.22972f
C9651 Iout.n275 VGND 0.22972f
C9652 Iout.n276 VGND 0.04584f
C9653 Iout.t247 VGND 0.02212f
C9654 Iout.n277 VGND 0.04919f
C9655 Iout.n278 VGND 0.02502f
C9656 Iout.n279 VGND 0.04584f
C9657 Iout.n280 VGND 0.22972f
C9658 Iout.n281 VGND 0.22972f
C9659 Iout.n282 VGND 0.04584f
C9660 Iout.t198 VGND 0.02212f
C9661 Iout.n283 VGND 0.04919f
C9662 Iout.n284 VGND 0.02502f
C9663 Iout.n285 VGND 0.04584f
C9664 Iout.n286 VGND 0.22972f
C9665 Iout.n287 VGND 0.22972f
C9666 Iout.n288 VGND 0.04584f
C9667 Iout.t149 VGND 0.02212f
C9668 Iout.n289 VGND 0.04919f
C9669 Iout.n290 VGND 0.02502f
C9670 Iout.n291 VGND 0.04584f
C9671 Iout.n292 VGND 0.22972f
C9672 Iout.n293 VGND 0.22972f
C9673 Iout.n294 VGND 0.04584f
C9674 Iout.t177 VGND 0.02212f
C9675 Iout.n295 VGND 0.04919f
C9676 Iout.n296 VGND 0.02502f
C9677 Iout.n297 VGND 0.04584f
C9678 Iout.n298 VGND 0.22972f
C9679 Iout.n299 VGND 0.22972f
C9680 Iout.n300 VGND 0.04584f
C9681 Iout.t67 VGND 0.02212f
C9682 Iout.n301 VGND 0.04919f
C9683 Iout.n302 VGND 0.02502f
C9684 Iout.n303 VGND 0.04584f
C9685 Iout.n304 VGND 0.22972f
C9686 Iout.t208 VGND 0.02212f
C9687 Iout.n305 VGND 0.04919f
C9688 Iout.n306 VGND 0.02502f
C9689 Iout.n307 VGND 0.04584f
C9690 Iout.t218 VGND 0.02212f
C9691 Iout.n308 VGND 0.04919f
C9692 Iout.n309 VGND 0.02502f
C9693 Iout.n310 VGND 0.04584f
C9694 Iout.t244 VGND 0.02212f
C9695 Iout.n311 VGND 0.04919f
C9696 Iout.n312 VGND 0.02502f
C9697 Iout.n313 VGND 0.04584f
C9698 Iout.t199 VGND 0.02212f
C9699 Iout.n314 VGND 0.04919f
C9700 Iout.n315 VGND 0.02502f
C9701 Iout.n316 VGND 0.04584f
C9702 Iout.t145 VGND 0.02212f
C9703 Iout.n317 VGND 0.04919f
C9704 Iout.n318 VGND 0.02502f
C9705 Iout.n319 VGND 0.04584f
C9706 Iout.t113 VGND 0.02212f
C9707 Iout.n320 VGND 0.04919f
C9708 Iout.n321 VGND 0.02502f
C9709 Iout.n322 VGND 0.04584f
C9710 Iout.t121 VGND 0.02212f
C9711 Iout.n323 VGND 0.04919f
C9712 Iout.n324 VGND 0.02502f
C9713 Iout.n325 VGND 0.04584f
C9714 Iout.t73 VGND 0.02212f
C9715 Iout.n326 VGND 0.04919f
C9716 Iout.n327 VGND 0.02502f
C9717 Iout.n328 VGND 0.04584f
C9718 Iout.t49 VGND 0.02212f
C9719 Iout.n329 VGND 0.04919f
C9720 Iout.n330 VGND 0.02502f
C9721 Iout.n331 VGND 0.04584f
C9722 Iout.n332 VGND 0.22972f
C9723 Iout.t74 VGND 0.02212f
C9724 Iout.n333 VGND 0.04919f
C9725 Iout.n334 VGND 0.02502f
C9726 Iout.n335 VGND 0.04584f
C9727 Iout.t223 VGND 0.02212f
C9728 Iout.n336 VGND 0.04919f
C9729 Iout.n337 VGND 0.02502f
C9730 Iout.n338 VGND 0.04584f
C9731 Iout.t59 VGND 0.02212f
C9732 Iout.n339 VGND 0.04919f
C9733 Iout.n340 VGND 0.02502f
C9734 Iout.n341 VGND 0.04584f
C9735 Iout.t155 VGND 0.02212f
C9736 Iout.n342 VGND 0.04919f
C9737 Iout.n343 VGND 0.02502f
C9738 Iout.n344 VGND 0.04584f
C9739 Iout.t207 VGND 0.02212f
C9740 Iout.n345 VGND 0.04919f
C9741 Iout.n346 VGND 0.02502f
C9742 Iout.n347 VGND 0.04584f
C9743 Iout.t172 VGND 0.02212f
C9744 Iout.n348 VGND 0.04919f
C9745 Iout.n349 VGND 0.02502f
C9746 Iout.n350 VGND 0.04584f
C9747 Iout.t194 VGND 0.02212f
C9748 Iout.n351 VGND 0.04919f
C9749 Iout.n352 VGND 0.02502f
C9750 Iout.n353 VGND 0.04584f
C9751 Iout.t102 VGND 0.02212f
C9752 Iout.n354 VGND 0.04919f
C9753 Iout.n355 VGND 0.02502f
C9754 Iout.n356 VGND 0.04584f
C9755 Iout.t138 VGND 0.02212f
C9756 Iout.n357 VGND 0.04919f
C9757 Iout.n358 VGND 0.02502f
C9758 Iout.n359 VGND 0.04584f
C9759 Iout.t210 VGND 0.02212f
C9760 Iout.n360 VGND 0.04919f
C9761 Iout.n361 VGND 0.02502f
C9762 Iout.n362 VGND 0.04584f
C9763 Iout.t147 VGND 0.02212f
C9764 Iout.n363 VGND 0.04919f
C9765 Iout.n364 VGND 0.02502f
C9766 Iout.n365 VGND 0.04584f
C9767 Iout.t25 VGND 0.02212f
C9768 Iout.n366 VGND 0.04919f
C9769 Iout.n367 VGND 0.02502f
C9770 Iout.n368 VGND 0.04584f
C9771 Iout.n369 VGND 0.22972f
C9772 Iout.t209 VGND 0.02212f
C9773 Iout.n370 VGND 0.04919f
C9774 Iout.n371 VGND 0.02502f
C9775 Iout.n372 VGND 0.04584f
C9776 Iout.n373 VGND 0.22972f
C9777 Iout.n374 VGND 0.22972f
C9778 Iout.n375 VGND 0.04584f
C9779 Iout.t157 VGND 0.02212f
C9780 Iout.n376 VGND 0.04919f
C9781 Iout.n377 VGND 0.02502f
C9782 Iout.t54 VGND 0.02212f
C9783 Iout.n378 VGND 0.04919f
C9784 Iout.n379 VGND 0.02502f
C9785 Iout.n380 VGND 0.04584f
C9786 Iout.n381 VGND 0.22972f
C9787 Iout.n382 VGND 0.22972f
C9788 Iout.n383 VGND 0.04584f
C9789 Iout.t104 VGND 0.02212f
C9790 Iout.n384 VGND 0.04919f
C9791 Iout.n385 VGND 0.02502f
C9792 Iout.t27 VGND 0.02212f
C9793 Iout.n386 VGND 0.04919f
C9794 Iout.n387 VGND 0.02502f
C9795 Iout.n388 VGND 0.04584f
C9796 Iout.n389 VGND 0.22972f
C9797 Iout.n390 VGND 0.22972f
C9798 Iout.n391 VGND 0.04584f
C9799 Iout.t226 VGND 0.02212f
C9800 Iout.n392 VGND 0.04919f
C9801 Iout.n393 VGND 0.02502f
C9802 Iout.t46 VGND 0.02212f
C9803 Iout.n394 VGND 0.04919f
C9804 Iout.n395 VGND 0.02502f
C9805 Iout.n396 VGND 0.04584f
C9806 Iout.n397 VGND 0.22972f
C9807 Iout.n398 VGND 0.22972f
C9808 Iout.n399 VGND 0.04584f
C9809 Iout.t182 VGND 0.02212f
C9810 Iout.n400 VGND 0.04919f
C9811 Iout.n401 VGND 0.02502f
C9812 Iout.t190 VGND 0.02212f
C9813 Iout.n402 VGND 0.04919f
C9814 Iout.n403 VGND 0.02502f
C9815 Iout.n404 VGND 0.04584f
C9816 Iout.n405 VGND 0.22972f
C9817 Iout.n406 VGND 0.22972f
C9818 Iout.n407 VGND 0.04584f
C9819 Iout.t228 VGND 0.02212f
C9820 Iout.n408 VGND 0.04919f
C9821 Iout.n409 VGND 0.02502f
C9822 Iout.t169 VGND 0.02212f
C9823 Iout.n410 VGND 0.04919f
C9824 Iout.n411 VGND 0.02502f
C9825 Iout.n412 VGND 0.04584f
C9826 Iout.n413 VGND 0.22972f
C9827 Iout.n414 VGND 0.22972f
C9828 Iout.n415 VGND 0.04584f
C9829 Iout.t90 VGND 0.02212f
C9830 Iout.n416 VGND 0.04919f
C9831 Iout.n417 VGND 0.02502f
C9832 Iout.t128 VGND 0.02212f
C9833 Iout.n418 VGND 0.04919f
C9834 Iout.n419 VGND 0.02502f
C9835 Iout.n420 VGND 0.04584f
C9836 Iout.n421 VGND 0.22972f
C9837 Iout.n422 VGND 0.22972f
C9838 Iout.n423 VGND 0.04584f
C9839 Iout.t88 VGND 0.02212f
C9840 Iout.n424 VGND 0.04919f
C9841 Iout.n425 VGND 0.02502f
C9842 Iout.t162 VGND 0.02212f
C9843 Iout.n426 VGND 0.04919f
C9844 Iout.n427 VGND 0.02502f
C9845 Iout.n428 VGND 0.04584f
C9846 Iout.n429 VGND 0.22972f
C9847 Iout.n430 VGND 0.22972f
C9848 Iout.n431 VGND 0.04584f
C9849 Iout.t134 VGND 0.02212f
C9850 Iout.n432 VGND 0.04919f
C9851 Iout.n433 VGND 0.02502f
C9852 Iout.t232 VGND 0.02212f
C9853 Iout.n434 VGND 0.04919f
C9854 Iout.n435 VGND 0.02502f
C9855 Iout.n436 VGND 0.22972f
C9856 Iout.n437 VGND 0.04584f
C9857 Iout.t156 VGND 0.02212f
C9858 Iout.n438 VGND 0.04919f
C9859 Iout.n439 VGND 0.02502f
C9860 Iout.n440 VGND 0.04584f
C9861 Iout.t42 VGND 0.02212f
C9862 Iout.n441 VGND 0.04919f
C9863 Iout.n442 VGND 0.02502f
C9864 Iout.n443 VGND 0.04584f
C9865 Iout.n444 VGND 0.22972f
C9866 Iout.n445 VGND 0.22972f
C9867 Iout.n446 VGND 0.04584f
C9868 Iout.t249 VGND 0.02212f
C9869 Iout.n447 VGND 0.04919f
C9870 Iout.n448 VGND 0.02502f
C9871 Iout.t158 VGND 0.02212f
C9872 Iout.n449 VGND 0.04919f
C9873 Iout.n450 VGND 0.02502f
C9874 Iout.n451 VGND 0.04584f
C9875 Iout.t37 VGND 0.02212f
C9876 Iout.n452 VGND 0.04919f
C9877 Iout.n453 VGND 0.02502f
C9878 Iout.n454 VGND 0.04584f
C9879 Iout.n455 VGND 0.22972f
C9880 Iout.n456 VGND 0.22972f
C9881 Iout.n457 VGND 0.04584f
C9882 Iout.t191 VGND 0.02212f
C9883 Iout.n458 VGND 0.04919f
C9884 Iout.n459 VGND 0.02502f
C9885 Iout.t108 VGND 0.02212f
C9886 Iout.n460 VGND 0.04919f
C9887 Iout.n461 VGND 0.02502f
C9888 Iout.n462 VGND 0.04584f
C9889 Iout.t216 VGND 0.02212f
C9890 Iout.n463 VGND 0.04919f
C9891 Iout.n464 VGND 0.02502f
C9892 Iout.n465 VGND 0.04584f
C9893 Iout.n466 VGND 0.22972f
C9894 Iout.n467 VGND 0.22972f
C9895 Iout.n468 VGND 0.04584f
C9896 Iout.t178 VGND 0.02212f
C9897 Iout.n469 VGND 0.04919f
C9898 Iout.n470 VGND 0.02502f
C9899 Iout.n471 VGND 0.04584f
C9900 Iout.t43 VGND 0.02212f
C9901 Iout.n472 VGND 0.04919f
C9902 Iout.n473 VGND 0.02502f
C9903 Iout.n474 VGND 0.04584f
C9904 Iout.n475 VGND 0.22972f
C9905 Iout.n476 VGND 0.22972f
C9906 Iout.n477 VGND 0.04584f
C9907 Iout.t17 VGND 0.02212f
C9908 Iout.n478 VGND 0.04919f
C9909 Iout.n479 VGND 0.02502f
C9910 Iout.t171 VGND 0.02212f
C9911 Iout.n480 VGND 0.04919f
C9912 Iout.n481 VGND 0.02502f
C9913 Iout.n482 VGND 0.04584f
C9914 Iout.t195 VGND 0.02212f
C9915 Iout.n483 VGND 0.04919f
C9916 Iout.n484 VGND 0.02502f
C9917 Iout.n485 VGND 0.04584f
C9918 Iout.n486 VGND 0.22972f
C9919 Iout.n487 VGND 0.22972f
C9920 Iout.n488 VGND 0.04584f
C9921 Iout.t170 VGND 0.02212f
C9922 Iout.n489 VGND 0.04919f
C9923 Iout.n490 VGND 0.02502f
C9924 Iout.t135 VGND 0.02212f
C9925 Iout.n491 VGND 0.04919f
C9926 Iout.n492 VGND 0.02502f
C9927 Iout.n493 VGND 0.04584f
C9928 Iout.t188 VGND 0.02212f
C9929 Iout.n494 VGND 0.04919f
C9930 Iout.n495 VGND 0.02502f
C9931 Iout.n496 VGND 0.04584f
C9932 Iout.n497 VGND 0.22972f
C9933 Iout.n498 VGND 0.13561f
C9934 Iout.n499 VGND 0.04584f
C9935 Iout.t148 VGND 0.02212f
C9936 Iout.n500 VGND 0.04919f
C9937 Iout.n501 VGND 0.02502f
C9938 Iout.n502 VGND 0.13561f
C9939 Iout.n503 VGND 0.04584f
C9940 Iout.t127 VGND 0.02212f
C9941 Iout.n504 VGND 0.04919f
C9942 Iout.n505 VGND 0.02502f
C9943 Iout.n506 VGND 0.04584f
C9944 Iout.t159 VGND 0.02212f
C9945 Iout.n507 VGND 0.04919f
C9946 Iout.n508 VGND 0.02502f
C9947 Iout.t142 VGND 0.02212f
C9948 Iout.n509 VGND 0.04919f
C9949 Iout.n510 VGND 0.02502f
C9950 Iout.n511 VGND 0.13561f
C9951 Iout.n512 VGND 0.04584f
C9952 Iout.t23 VGND 0.02212f
C9953 Iout.n513 VGND 0.04919f
C9954 Iout.n514 VGND 0.02502f
C9955 Iout.n515 VGND 0.04584f
C9956 Iout.n516 VGND 0.13561f
C9957 Iout.n517 VGND 0.22972f
C9958 Iout.n518 VGND 0.04584f
C9959 Iout.t139 VGND 0.02212f
C9960 Iout.n519 VGND 0.04919f
C9961 Iout.n520 VGND 0.02502f
C9962 Iout.n521 VGND 0.04584f
C9963 Iout.n522 VGND 0.22972f
C9964 Iout.n523 VGND 0.22972f
C9965 Iout.n524 VGND 0.04584f
C9966 Iout.t246 VGND 0.02212f
C9967 Iout.n525 VGND 0.04919f
C9968 Iout.n526 VGND 0.02502f
C9969 Iout.n527 VGND 0.04584f
C9970 Iout.n528 VGND 0.22972f
C9971 Iout.n529 VGND 0.22972f
C9972 Iout.n530 VGND 0.04584f
C9973 Iout.t22 VGND 0.02212f
C9974 Iout.n531 VGND 0.04919f
C9975 Iout.n532 VGND 0.02502f
C9976 Iout.n533 VGND 0.04584f
C9977 Iout.t163 VGND 0.02212f
C9978 Iout.n534 VGND 0.04919f
C9979 Iout.n535 VGND 0.02502f
C9980 Iout.t80 VGND 0.02212f
C9981 Iout.n536 VGND 0.04919f
C9982 Iout.n537 VGND 0.02502f
C9983 Iout.n538 VGND 0.04584f
C9984 Iout.n539 VGND 0.22972f
C9985 Iout.n540 VGND 0.22972f
C9986 Iout.n541 VGND 0.04584f
C9987 Iout.t28 VGND 0.02212f
C9988 Iout.n542 VGND 0.04919f
C9989 Iout.n543 VGND 0.02502f
C9990 Iout.n544 VGND 0.04584f
C9991 Iout.n545 VGND 0.22972f
C9992 Iout.n546 VGND 0.22972f
C9993 Iout.n547 VGND 0.04584f
C9994 Iout.t72 VGND 0.02212f
C9995 Iout.n548 VGND 0.04919f
C9996 Iout.n549 VGND 0.02502f
C9997 Iout.n550 VGND 0.04584f
C9998 Iout.n551 VGND 0.22972f
C9999 Iout.n552 VGND 0.22972f
C10000 Iout.n553 VGND 0.04584f
C10001 Iout.t51 VGND 0.02212f
C10002 Iout.n554 VGND 0.04919f
C10003 Iout.n555 VGND 0.02502f
C10004 Iout.n556 VGND 0.04584f
C10005 Iout.t116 VGND 0.02212f
C10006 Iout.n557 VGND 0.04919f
C10007 Iout.n558 VGND 0.02502f
C10008 Iout.t196 VGND 0.02212f
C10009 Iout.n559 VGND 0.04919f
C10010 Iout.n560 VGND 0.02502f
C10011 Iout.n561 VGND 0.04584f
C10012 Iout.n562 VGND 0.22972f
C10013 Iout.t114 VGND 0.02212f
C10014 Iout.n563 VGND 0.04919f
C10015 Iout.n564 VGND 0.02502f
C10016 Iout.n565 VGND 0.04584f
C10017 Iout.n566 VGND 0.22972f
C10018 Iout.n567 VGND 0.22972f
C10019 Iout.n568 VGND 0.04584f
C10020 Iout.t237 VGND 0.02212f
C10021 Iout.n569 VGND 0.04919f
C10022 Iout.n570 VGND 0.02502f
C10023 Iout.n571 VGND 0.04584f
C10024 Iout.n572 VGND 0.22972f
C10025 Iout.t68 VGND 0.02212f
C10026 Iout.n573 VGND 0.04919f
C10027 Iout.n574 VGND 0.02502f
C10028 Iout.n575 VGND 0.04584f
C10029 Iout.t45 VGND 0.02212f
C10030 Iout.n576 VGND 0.04919f
C10031 Iout.n577 VGND 0.02502f
C10032 Iout.n578 VGND 0.04584f
C10033 Iout.n579 VGND 0.22972f
C10034 Iout.n580 VGND 0.22972f
C10035 Iout.n581 VGND 0.04584f
C10036 Iout.t123 VGND 0.02212f
C10037 Iout.n582 VGND 0.04919f
C10038 Iout.n583 VGND 0.02502f
C10039 Iout.n584 VGND 0.04584f
C10040 Iout.n585 VGND 0.22972f
C10041 Iout.n586 VGND 0.22972f
C10042 Iout.n587 VGND 0.04584f
C10043 Iout.t231 VGND 0.02212f
C10044 Iout.n588 VGND 0.04919f
C10045 Iout.n589 VGND 0.02502f
C10046 Iout.n590 VGND 0.04584f
C10047 Iout.n591 VGND 0.22972f
C10048 Iout.n592 VGND 0.22972f
C10049 Iout.n593 VGND 0.04584f
C10050 Iout.t117 VGND 0.02212f
C10051 Iout.n594 VGND 0.04919f
C10052 Iout.n595 VGND 0.02502f
C10053 Iout.n596 VGND 0.04584f
C10054 Iout.n597 VGND 0.22972f
C10055 Iout.n598 VGND 0.22972f
C10056 Iout.n599 VGND 0.04584f
C10057 Iout.t70 VGND 0.02212f
C10058 Iout.n600 VGND 0.04919f
C10059 Iout.n601 VGND 0.02502f
C10060 Iout.n602 VGND 0.04584f
C10061 Iout.n603 VGND 0.22972f
C10062 Iout.n604 VGND 0.22972f
C10063 Iout.n605 VGND 0.04584f
C10064 Iout.t205 VGND 0.02212f
C10065 Iout.n606 VGND 0.04919f
C10066 Iout.n607 VGND 0.02502f
C10067 Iout.n608 VGND 0.04584f
C10068 Iout.n609 VGND 0.22972f
C10069 Iout.n610 VGND 0.22972f
C10070 Iout.n611 VGND 0.04584f
C10071 Iout.t57 VGND 0.02212f
C10072 Iout.n612 VGND 0.04919f
C10073 Iout.n613 VGND 0.02502f
C10074 Iout.n614 VGND 0.04584f
C10075 Iout.n615 VGND 0.22972f
C10076 Iout.n616 VGND 0.22972f
C10077 Iout.n617 VGND 0.04584f
C10078 Iout.t64 VGND 0.02212f
C10079 Iout.n618 VGND 0.04919f
C10080 Iout.n619 VGND 0.02502f
C10081 Iout.n620 VGND 0.04584f
C10082 Iout.n621 VGND 0.22972f
C10083 Iout.n622 VGND 0.22972f
C10084 Iout.n623 VGND 0.04584f
C10085 Iout.t152 VGND 0.02212f
C10086 Iout.n624 VGND 0.04919f
C10087 Iout.n625 VGND 0.02502f
C10088 Iout.n626 VGND 0.04584f
C10089 Iout.n627 VGND 0.22972f
C10090 Iout.n628 VGND 0.22972f
C10091 Iout.n629 VGND 0.04584f
C10092 Iout.t9 VGND 0.02212f
C10093 Iout.n630 VGND 0.04919f
C10094 Iout.n631 VGND 0.02502f
C10095 Iout.n632 VGND 0.04584f
C10096 Iout.n633 VGND 0.22972f
C10097 Iout.n634 VGND 0.22972f
C10098 Iout.n635 VGND 0.04584f
C10099 Iout.t140 VGND 0.02212f
C10100 Iout.n636 VGND 0.04919f
C10101 Iout.n637 VGND 0.02502f
C10102 Iout.n638 VGND 0.04584f
C10103 Iout.n639 VGND 0.22972f
C10104 Iout.n640 VGND 0.22972f
C10105 Iout.n641 VGND 0.04584f
C10106 Iout.t180 VGND 0.02212f
C10107 Iout.n642 VGND 0.04919f
C10108 Iout.n643 VGND 0.02502f
C10109 Iout.n644 VGND 0.04584f
C10110 Iout.n645 VGND 0.22972f
C10111 Iout.n646 VGND 0.22972f
C10112 Iout.n647 VGND 0.04584f
C10113 Iout.t220 VGND 0.02212f
C10114 Iout.n648 VGND 0.04919f
C10115 Iout.n649 VGND 0.02502f
C10116 Iout.n650 VGND 0.04584f
C10117 Iout.n651 VGND 0.22972f
C10118 Iout.n652 VGND 0.22972f
C10119 Iout.n653 VGND 0.04584f
C10120 Iout.t221 VGND 0.02212f
C10121 Iout.n654 VGND 0.04919f
C10122 Iout.n655 VGND 0.02502f
C10123 Iout.n656 VGND 0.04584f
C10124 Iout.t96 VGND 0.02212f
C10125 Iout.n657 VGND 0.04919f
C10126 Iout.n658 VGND 0.02502f
C10127 Iout.n659 VGND 0.04584f
C10128 Iout.t41 VGND 0.02212f
C10129 Iout.n660 VGND 0.04919f
C10130 Iout.n661 VGND 0.02502f
C10131 Iout.n662 VGND 0.04584f
C10132 Iout.t58 VGND 0.02212f
C10133 Iout.n663 VGND 0.04919f
C10134 Iout.n664 VGND 0.02502f
C10135 Iout.n665 VGND 0.04584f
C10136 Iout.t86 VGND 0.02212f
C10137 Iout.n666 VGND 0.04919f
C10138 Iout.n667 VGND 0.02502f
C10139 Iout.n668 VGND 0.04584f
C10140 Iout.t164 VGND 0.02212f
C10141 Iout.n669 VGND 0.04919f
C10142 Iout.n670 VGND 0.02502f
C10143 Iout.n671 VGND 0.04584f
C10144 Iout.t186 VGND 0.02212f
C10145 Iout.n672 VGND 0.04919f
C10146 Iout.n673 VGND 0.02502f
C10147 Iout.n674 VGND 0.04584f
C10148 Iout.t47 VGND 0.02212f
C10149 Iout.n675 VGND 0.04919f
C10150 Iout.n676 VGND 0.02502f
C10151 Iout.n677 VGND 0.04584f
C10152 Iout.t143 VGND 0.02212f
C10153 Iout.n678 VGND 0.04919f
C10154 Iout.n679 VGND 0.02502f
C10155 Iout.n680 VGND 0.04584f
C10156 Iout.t39 VGND 0.02212f
C10157 Iout.n681 VGND 0.04919f
C10158 Iout.n682 VGND 0.02502f
C10159 Iout.n683 VGND 0.04584f
C10160 Iout.t31 VGND 0.02212f
C10161 Iout.n684 VGND 0.04919f
C10162 Iout.n685 VGND 0.02502f
C10163 Iout.n686 VGND 0.04584f
C10164 Iout.t105 VGND 0.02212f
C10165 Iout.n687 VGND 0.04919f
C10166 Iout.n688 VGND 0.02502f
C10167 Iout.n689 VGND 0.04584f
C10168 Iout.t242 VGND 0.02212f
C10169 Iout.n690 VGND 0.04919f
C10170 Iout.n691 VGND 0.02502f
C10171 Iout.t183 VGND 0.02212f
C10172 Iout.n692 VGND 0.04919f
C10173 Iout.n693 VGND 0.02502f
C10174 Iout.n694 VGND 0.04584f
C10175 Iout.t82 VGND 0.02212f
C10176 Iout.n695 VGND 0.04919f
C10177 Iout.n696 VGND 0.02502f
C10178 Iout.n697 VGND 0.04584f
C10179 Iout.n698 VGND 0.22972f
C10180 Iout.t222 VGND 0.02212f
C10181 Iout.n699 VGND 0.04919f
C10182 Iout.n700 VGND 0.02502f
C10183 Iout.n701 VGND 0.04584f
C10184 Iout.n702 VGND 0.22972f
C10185 Iout.n703 VGND 0.22972f
C10186 Iout.n704 VGND 0.04584f
C10187 Iout.t154 VGND 0.02212f
C10188 Iout.n705 VGND 0.04919f
C10189 Iout.n706 VGND 0.02502f
C10190 Iout.n707 VGND 0.04584f
C10191 Iout.n708 VGND 0.22972f
C10192 Iout.n709 VGND 0.22972f
C10193 Iout.n710 VGND 0.04584f
C10194 Iout.t109 VGND 0.02212f
C10195 Iout.n711 VGND 0.04919f
C10196 Iout.n712 VGND 0.02502f
C10197 Iout.n713 VGND 0.04584f
C10198 Iout.n714 VGND 0.22972f
C10199 Iout.n715 VGND 0.22972f
C10200 Iout.n716 VGND 0.04584f
C10201 Iout.t146 VGND 0.02212f
C10202 Iout.n717 VGND 0.04919f
C10203 Iout.n718 VGND 0.02502f
C10204 Iout.n719 VGND 0.04584f
C10205 Iout.n720 VGND 0.22972f
C10206 Iout.n721 VGND 0.22972f
C10207 Iout.n722 VGND 0.04584f
C10208 Iout.t100 VGND 0.02212f
C10209 Iout.n723 VGND 0.04919f
C10210 Iout.n724 VGND 0.02502f
C10211 Iout.n725 VGND 0.04584f
C10212 Iout.n726 VGND 0.22972f
C10213 Iout.n727 VGND 0.22972f
C10214 Iout.n728 VGND 0.04584f
C10215 Iout.t217 VGND 0.02212f
C10216 Iout.n729 VGND 0.04919f
C10217 Iout.n730 VGND 0.02502f
C10218 Iout.n731 VGND 0.04584f
C10219 Iout.n732 VGND 0.22972f
C10220 Iout.n733 VGND 0.22972f
C10221 Iout.n734 VGND 0.04584f
C10222 Iout.t97 VGND 0.02212f
C10223 Iout.n735 VGND 0.04919f
C10224 Iout.n736 VGND 0.02502f
C10225 Iout.n737 VGND 0.04584f
C10226 Iout.n738 VGND 0.22972f
C10227 Iout.n739 VGND 0.22972f
C10228 Iout.n740 VGND 0.04584f
C10229 Iout.t103 VGND 0.02212f
C10230 Iout.n741 VGND 0.04919f
C10231 Iout.n742 VGND 0.02502f
C10232 Iout.n743 VGND 0.04584f
C10233 Iout.n744 VGND 0.22972f
C10234 Iout.n745 VGND 0.22972f
C10235 Iout.n746 VGND 0.04584f
C10236 Iout.t236 VGND 0.02212f
C10237 Iout.n747 VGND 0.04919f
C10238 Iout.n748 VGND 0.02502f
C10239 Iout.n749 VGND 0.04584f
C10240 Iout.n750 VGND 0.22972f
C10241 Iout.n751 VGND 0.22972f
C10242 Iout.n752 VGND 0.04584f
C10243 Iout.t151 VGND 0.02212f
C10244 Iout.n753 VGND 0.04919f
C10245 Iout.n754 VGND 0.02502f
C10246 Iout.n755 VGND 0.04584f
C10247 Iout.n756 VGND 0.22972f
C10248 Iout.n757 VGND 0.22972f
C10249 Iout.n758 VGND 0.04584f
C10250 Iout.t137 VGND 0.02212f
C10251 Iout.n759 VGND 0.04919f
C10252 Iout.n760 VGND 0.02502f
C10253 Iout.n761 VGND 0.04584f
C10254 Iout.n762 VGND 0.22972f
C10255 Iout.n763 VGND 0.22972f
C10256 Iout.n764 VGND 0.04584f
C10257 Iout.t252 VGND 0.02212f
C10258 Iout.n765 VGND 0.04919f
C10259 Iout.n766 VGND 0.02502f
C10260 Iout.n767 VGND 0.04584f
C10261 Iout.n768 VGND 0.22972f
C10262 Iout.n769 VGND 0.22972f
C10263 Iout.n770 VGND 0.04584f
C10264 Iout.t35 VGND 0.02212f
C10265 Iout.n771 VGND 0.04919f
C10266 Iout.n772 VGND 0.02502f
C10267 Iout.n773 VGND 0.04584f
C10268 Iout.n774 VGND 0.22972f
C10269 Iout.n775 VGND 0.22972f
C10270 Iout.n776 VGND 0.04584f
C10271 Iout.t60 VGND 0.02212f
C10272 Iout.n777 VGND 0.04919f
C10273 Iout.n778 VGND 0.02502f
C10274 Iout.n779 VGND 0.04584f
C10275 Iout.n780 VGND 0.22972f
C10276 Iout.t87 VGND 0.02212f
C10277 Iout.n781 VGND 0.04919f
C10278 Iout.n782 VGND 0.02502f
C10279 Iout.n783 VGND 0.04584f
C10280 Iout.t26 VGND 0.02212f
C10281 Iout.n784 VGND 0.04919f
C10282 Iout.n785 VGND 0.02502f
C10283 Iout.n786 VGND 0.04584f
C10284 Iout.t4 VGND 0.02212f
C10285 Iout.n787 VGND 0.04919f
C10286 Iout.n788 VGND 0.02502f
C10287 Iout.n789 VGND 0.04584f
C10288 Iout.t83 VGND 0.02212f
C10289 Iout.n790 VGND 0.04919f
C10290 Iout.n791 VGND 0.02502f
C10291 Iout.n792 VGND 0.04584f
C10292 Iout.t77 VGND 0.02212f
C10293 Iout.n793 VGND 0.04919f
C10294 Iout.n794 VGND 0.02502f
C10295 Iout.n795 VGND 0.04584f
C10296 Iout.t187 VGND 0.02212f
C10297 Iout.n796 VGND 0.04919f
C10298 Iout.n797 VGND 0.02502f
C10299 Iout.n798 VGND 0.04584f
C10300 Iout.t192 VGND 0.02212f
C10301 Iout.n799 VGND 0.04919f
C10302 Iout.n800 VGND 0.02502f
C10303 Iout.n801 VGND 0.04584f
C10304 Iout.t243 VGND 0.02212f
C10305 Iout.n802 VGND 0.04919f
C10306 Iout.n803 VGND 0.02502f
C10307 Iout.n804 VGND 0.04584f
C10308 Iout.t160 VGND 0.02212f
C10309 Iout.n805 VGND 0.04919f
C10310 Iout.n806 VGND 0.02502f
C10311 Iout.n807 VGND 0.04584f
C10312 Iout.t239 VGND 0.02212f
C10313 Iout.n808 VGND 0.04919f
C10314 Iout.n809 VGND 0.02502f
C10315 Iout.n810 VGND 0.04584f
C10316 Iout.t202 VGND 0.02212f
C10317 Iout.n811 VGND 0.04919f
C10318 Iout.n812 VGND 0.02502f
C10319 Iout.n813 VGND 0.04584f
C10320 Iout.t119 VGND 0.02212f
C10321 Iout.n814 VGND 0.04919f
C10322 Iout.n815 VGND 0.02502f
C10323 Iout.n816 VGND 0.04584f
C10324 Iout.t19 VGND 0.02212f
C10325 Iout.n817 VGND 0.04919f
C10326 Iout.n818 VGND 0.02502f
C10327 Iout.n819 VGND 0.04584f
C10328 Iout.t63 VGND 0.02212f
C10329 Iout.n820 VGND 0.04919f
C10330 Iout.n821 VGND 0.02502f
C10331 Iout.n822 VGND 0.04584f
C10332 Iout.t166 VGND 0.02212f
C10333 Iout.n823 VGND 0.04919f
C10334 Iout.n824 VGND 0.02502f
C10335 Iout.n825 VGND 0.04584f
C10336 Iout.n826 VGND 0.22972f
C10337 Iout.t141 VGND 0.02212f
C10338 Iout.n827 VGND 0.04919f
C10339 Iout.n828 VGND 0.02502f
C10340 Iout.n829 VGND 0.07841f
C10341 Iout.n830 VGND 0.47625f
C10342 Iout.n831 VGND 0.04584f
C10343 Iout.t241 VGND 0.02212f
C10344 Iout.n832 VGND 0.04919f
C10345 Iout.n833 VGND 0.02502f
C10346 Iout.t30 VGND 0.02212f
C10347 Iout.n834 VGND 0.04919f
C10348 Iout.n835 VGND 0.02502f
C10349 Iout.n836 VGND 0.04584f
C10350 Iout.n837 VGND 0.47625f
C10351 Iout.n838 VGND 0.07841f
C10352 Iout.t11 VGND 0.02212f
C10353 Iout.n839 VGND 0.04919f
C10354 Iout.n840 VGND 0.02502f
C10355 Iout.t129 VGND 0.02212f
C10356 Iout.n841 VGND 0.04919f
C10357 Iout.n842 VGND 0.02502f
C10358 Iout.n843 VGND 0.07841f
C10359 Iout.n844 VGND 0.47625f
C10360 Iout.n845 VGND 0.04584f
C10361 Iout.t144 VGND 0.02212f
C10362 Iout.n846 VGND 0.04919f
C10363 Iout.n847 VGND 0.02502f
C10364 Iout.t215 VGND 0.02212f
C10365 Iout.n848 VGND 0.04919f
C10366 Iout.n849 VGND 0.02502f
C10367 Iout.n850 VGND 0.04584f
C10368 Iout.n851 VGND 0.47625f
C10369 Iout.n852 VGND 0.07841f
C10370 Iout.t66 VGND 0.02212f
C10371 Iout.n853 VGND 0.04919f
C10372 Iout.n854 VGND 0.02502f
C10373 Iout.t130 VGND 0.02212f
C10374 Iout.n855 VGND 0.04919f
C10375 Iout.n856 VGND 0.02502f
C10376 Iout.n857 VGND 0.07841f
C10377 Iout.n858 VGND 0.47625f
C10378 Iout.n859 VGND 0.04584f
C10379 Iout.t153 VGND 0.02212f
C10380 Iout.n860 VGND 0.04919f
C10381 Iout.n861 VGND 0.02502f
C10382 Iout.t251 VGND 0.02212f
C10383 Iout.n862 VGND 0.04919f
C10384 Iout.n863 VGND 0.02502f
C10385 Iout.n864 VGND 0.04584f
C10386 Iout.n865 VGND 0.47625f
C10387 Iout.n866 VGND 0.07841f
C10388 Iout.t219 VGND 0.02212f
C10389 Iout.n867 VGND 0.04919f
C10390 Iout.n868 VGND 0.02502f
C10391 Iout.t176 VGND 0.02212f
C10392 Iout.n869 VGND 0.04919f
C10393 Iout.n870 VGND 0.02502f
C10394 Iout.n871 VGND 0.07841f
C10395 Iout.n872 VGND 0.47625f
C10396 Iout.n873 VGND 0.04584f
C10397 Iout.t55 VGND 0.02212f
C10398 Iout.n874 VGND 0.04919f
C10399 Iout.n875 VGND 0.02502f
C10400 Iout.t204 VGND 0.02212f
C10401 Iout.n876 VGND 0.04919f
C10402 Iout.n877 VGND 0.02502f
C10403 Iout.n878 VGND 0.04584f
C10404 Iout.n879 VGND 0.47625f
C10405 Iout.n880 VGND 0.07841f
C10406 Iout.t56 VGND 0.02212f
C10407 Iout.n881 VGND 0.04919f
C10408 Iout.n882 VGND 0.02502f
C10409 Iout.t150 VGND 0.02212f
C10410 Iout.n883 VGND 0.04919f
C10411 Iout.n884 VGND 0.02502f
C10412 Iout.n885 VGND 0.07841f
C10413 Iout.n886 VGND 0.47625f
C10414 Iout.n887 VGND 0.04584f
C10415 Iout.t71 VGND 0.02212f
C10416 Iout.n888 VGND 0.04919f
C10417 Iout.n889 VGND 0.02502f
C10418 Iout.t165 VGND 0.02212f
C10419 Iout.n890 VGND 0.04919f
C10420 Iout.n891 VGND 0.02502f
C10421 Iout.n892 VGND 0.04584f
C10422 Iout.n893 VGND 0.47625f
C10423 Iout.n894 VGND 0.07841f
C10424 Iout.t76 VGND 0.02212f
C10425 Iout.n895 VGND 0.04919f
C10426 Iout.n896 VGND 0.02502f
C10427 Iout.t14 VGND 0.02212f
C10428 Iout.n897 VGND 0.04919f
C10429 Iout.n898 VGND 0.02502f
C10430 Iout.n899 VGND 0.07841f
C10431 Iout.n900 VGND 0.47625f
C10432 Iout.n901 VGND 0.04584f
C10433 Iout.t65 VGND 0.02212f
C10434 Iout.n902 VGND 0.04919f
C10435 Iout.n903 VGND 0.02502f
C10436 Iout.t206 VGND 0.02212f
C10437 Iout.n904 VGND 0.04919f
C10438 Iout.n905 VGND 0.02502f
C10439 Iout.n906 VGND 0.04584f
C10440 Iout.n907 VGND 0.47625f
C10441 Iout.n908 VGND 0.07841f
C10442 Iout.t254 VGND 0.02212f
C10443 Iout.n909 VGND 0.04919f
C10444 Iout.n910 VGND 0.02502f
C10445 Iout.t62 VGND 0.02212f
C10446 Iout.n911 VGND 0.04919f
C10447 Iout.n912 VGND 0.02502f
C10448 Iout.n913 VGND 0.07841f
C10449 Iout.n914 VGND 0.47625f
C10450 Iout.n915 VGND 0.04584f
C10451 Iout.t213 VGND 0.02212f
C10452 Iout.n916 VGND 0.04919f
C10453 Iout.n917 VGND 0.02502f
C10454 Iout.t99 VGND 0.02212f
C10455 Iout.n918 VGND 0.04919f
C10456 Iout.n919 VGND 0.02502f
C10457 Iout.n920 VGND 0.04584f
C10458 Iout.n921 VGND 0.47625f
C10459 Iout.n922 VGND 0.07841f
C10460 Iout.t33 VGND 0.02212f
C10461 Iout.n923 VGND 0.04919f
C10462 Iout.n924 VGND 0.02502f
C10463 Iout.n925 VGND 0.07841f
C10464 Iout.t115 VGND 0.02212f
C10465 Iout.n926 VGND 0.04919f
C10466 Iout.n927 VGND 0.02502f
C10467 Iout.n928 VGND 0.07841f
C10468 Iout.n929 VGND 0.47625f
C10469 Iout.n930 VGND 0.04584f
C10470 Iout.t179 VGND 0.02212f
C10471 Iout.n931 VGND 0.04919f
C10472 Iout.n932 VGND 0.02502f
C10473 Iout.n933 VGND 0.04584f
C10474 Iout.t224 VGND 0.02212f
C10475 Iout.n934 VGND 0.04919f
C10476 Iout.n935 VGND 0.19431f
C10477 Iout.n936 VGND 2.54526f
C10478 Iout.n937 VGND 1.20114f
C10479 Iout.t235 VGND 0.02212f
C10480 Iout.n938 VGND 0.04919f
C10481 Iout.n939 VGND 0.19431f
C10482 Iout.n940 VGND 0.04584f
C10483 Iout.n941 VGND 0.22972f
C10484 Iout.n942 VGND 0.22972f
C10485 Iout.n943 VGND 0.04584f
C10486 Iout.t5 VGND 0.02212f
C10487 Iout.n944 VGND 0.04919f
C10488 Iout.n945 VGND 0.02502f
C10489 Iout.n946 VGND 0.04584f
C10490 Iout.n947 VGND 0.22972f
C10491 Iout.n948 VGND 0.22972f
C10492 Iout.n949 VGND 0.04584f
C10493 Iout.t238 VGND 0.02212f
C10494 Iout.n950 VGND 0.04919f
C10495 Iout.n951 VGND 0.02502f
C10496 Iout.n952 VGND 0.04584f
C10497 Iout.t15 VGND 0.02212f
C10498 Iout.n953 VGND 0.04919f
C10499 Iout.n954 VGND 0.19431f
C10500 Iout.n955 VGND 1.20114f
C10501 Iout.n956 VGND 1.20114f
C10502 Iout.t95 VGND 0.02212f
C10503 Iout.n957 VGND 0.04919f
C10504 Iout.n958 VGND 0.19431f
C10505 Iout.n959 VGND 0.04584f
C10506 Iout.n960 VGND 0.22972f
C10507 Iout.n961 VGND 0.22972f
C10508 Iout.n962 VGND 0.04584f
C10509 Iout.t36 VGND 0.02212f
C10510 Iout.n963 VGND 0.04919f
C10511 Iout.n964 VGND 0.02502f
C10512 Iout.n965 VGND 0.04584f
C10513 Iout.n966 VGND 0.22972f
C10514 Iout.n967 VGND 0.22972f
C10515 Iout.n968 VGND 0.04584f
C10516 Iout.t122 VGND 0.02212f
C10517 Iout.n969 VGND 0.04919f
C10518 Iout.n970 VGND 0.02502f
C10519 Iout.n971 VGND 0.04584f
C10520 Iout.t1 VGND 0.02212f
C10521 Iout.n972 VGND 0.04919f
C10522 Iout.n973 VGND 0.19431f
C10523 Iout.n974 VGND 1.20114f
C10524 Iout.n975 VGND 1.20114f
C10525 Iout.t107 VGND 0.02212f
C10526 Iout.n976 VGND 0.04919f
C10527 Iout.n977 VGND 0.19431f
C10528 Iout.n978 VGND 0.04584f
C10529 Iout.n979 VGND 0.22972f
C10530 Iout.n980 VGND 0.22972f
C10531 Iout.n981 VGND 0.04584f
C10532 Iout.t240 VGND 0.02212f
C10533 Iout.n982 VGND 0.04919f
C10534 Iout.n983 VGND 0.02502f
C10535 Iout.n984 VGND 0.04584f
C10536 Iout.n985 VGND 0.22972f
C10537 Iout.n986 VGND 0.22972f
C10538 Iout.n987 VGND 0.04584f
C10539 Iout.t111 VGND 0.02212f
C10540 Iout.n988 VGND 0.04919f
C10541 Iout.n989 VGND 0.02502f
C10542 Iout.n990 VGND 0.04584f
C10543 Iout.t38 VGND 0.02212f
C10544 Iout.n991 VGND 0.04919f
C10545 Iout.n992 VGND 0.19431f
C10546 Iout.n993 VGND 1.20114f
C10547 Iout.n994 VGND 1.20114f
C10548 Iout.t53 VGND 0.02212f
C10549 Iout.n995 VGND 0.04919f
C10550 Iout.n996 VGND 0.19431f
C10551 Iout.n997 VGND 0.04584f
C10552 Iout.n998 VGND 0.22972f
C10553 Iout.n999 VGND 0.22972f
C10554 Iout.n1000 VGND 0.04584f
C10555 Iout.t124 VGND 0.02212f
C10556 Iout.n1001 VGND 0.04919f
C10557 Iout.n1002 VGND 0.02502f
C10558 Iout.n1003 VGND 0.04584f
C10559 Iout.n1004 VGND 0.22972f
C10560 Iout.n1005 VGND 0.22972f
C10561 Iout.n1006 VGND 0.04584f
C10562 Iout.t16 VGND 0.02212f
C10563 Iout.n1007 VGND 0.04919f
C10564 Iout.n1008 VGND 0.02502f
C10565 Iout.n1009 VGND 0.04584f
C10566 Iout.t106 VGND 0.02212f
C10567 Iout.n1010 VGND 0.04919f
C10568 Iout.n1011 VGND 0.19431f
C10569 Iout.n1012 VGND 1.20114f
C10570 Iout.n1013 VGND 1.07853f
C10571 Iout.t98 VGND 0.02212f
C10572 Iout.n1014 VGND 0.04919f
C10573 Iout.n1015 VGND 0.19431f
C10574 Iout.n1016 VGND 0.04584f
C10575 Iout.n1017 VGND 0.22972f
C10576 Iout.n1018 VGND 0.13561f
C10577 Iout.n1019 VGND 0.04584f
C10578 Iout.t174 VGND 0.02212f
C10579 Iout.n1020 VGND 0.04919f
C10580 Iout.n1021 VGND 0.19431f
C10581 Iout.n1022 VGND 0.22314f
C10582 VPWR.n0 VGND 0.03466f
C10583 VPWR.t551 VGND 0.21918f
C10584 VPWR.t740 VGND 0.09699f
C10585 VPWR.t955 VGND 0.27964f
C10586 VPWR.t938 VGND 0.10581f
C10587 VPWR.t332 VGND 0.10581f
C10588 VPWR.t329 VGND 0.10581f
C10589 VPWR.t1194 VGND 0.10581f
C10590 VPWR.t985 VGND 0.10581f
C10591 VPWR.t981 VGND 0.10581f
C10592 VPWR.t1117 VGND 0.07432f
C10593 VPWR.n1 VGND 0.13503f
C10594 VPWR.n2 VGND 0.07145f
C10595 VPWR.t741 VGND 0.04227f
C10596 VPWR.t1118 VGND 0.0106f
C10597 VPWR.t982 VGND 0.0106f
C10598 VPWR.n4 VGND 0.02326f
C10599 VPWR.t986 VGND 0.0106f
C10600 VPWR.t1195 VGND 0.0106f
C10601 VPWR.n5 VGND 0.02322f
C10602 VPWR.n6 VGND 0.0477f
C10603 VPWR.n7 VGND 0.13446f
C10604 VPWR.n8 VGND 0.04257f
C10605 VPWR.n9 VGND 0.03127f
C10606 VPWR.n10 VGND 0.05604f
C10607 VPWR.n12 VGND 0.01206f
C10608 VPWR.n13 VGND 0.01413f
C10609 VPWR.n14 VGND 0.02072f
C10610 VPWR.n15 VGND 0.06272f
C10611 VPWR.t552 VGND 0.04226f
C10612 VPWR.n17 VGND 0.05435f
C10613 VPWR.n18 VGND 0.2482f
C10614 VPWR.n19 VGND 0.72374f
C10615 VPWR.n20 VGND 0.23558f
C10616 VPWR.n21 VGND 0.75117f
C10617 VPWR.n22 VGND 0.1027f
C10618 VPWR.n23 VGND 0.02214f
C10619 VPWR.n24 VGND 0.05881f
C10620 VPWR.n25 VGND 0.02214f
C10621 VPWR.n26 VGND 0.11837f
C10622 VPWR.n27 VGND 0.02214f
C10623 VPWR.n28 VGND 0.09431f
C10624 VPWR.n29 VGND 0.02214f
C10625 VPWR.n30 VGND 0.09431f
C10626 VPWR.n31 VGND 0.02214f
C10627 VPWR.n32 VGND 0.09431f
C10628 VPWR.n33 VGND 0.02214f
C10629 VPWR.n34 VGND 0.09431f
C10630 VPWR.n35 VGND 0.02214f
C10631 VPWR.n36 VGND 0.09431f
C10632 VPWR.n37 VGND 0.02214f
C10633 VPWR.n38 VGND 0.09431f
C10634 VPWR.n39 VGND 0.02214f
C10635 VPWR.n40 VGND 0.09431f
C10636 VPWR.n41 VGND 0.02214f
C10637 VPWR.n42 VGND 0.09431f
C10638 VPWR.n43 VGND 0.02214f
C10639 VPWR.n44 VGND 0.09431f
C10640 VPWR.n45 VGND 0.02214f
C10641 VPWR.n46 VGND 0.09431f
C10642 VPWR.n47 VGND 0.02214f
C10643 VPWR.n48 VGND 0.09431f
C10644 VPWR.n49 VGND 0.02214f
C10645 VPWR.n50 VGND 0.09431f
C10646 VPWR.n51 VGND 0.02214f
C10647 VPWR.n52 VGND 0.09431f
C10648 VPWR.n53 VGND 0.02214f
C10649 VPWR.n54 VGND 0.10211f
C10650 VPWR.n55 VGND 0.08525f
C10651 VPWR.t1486 VGND 0.02464f
C10652 VPWR.t1591 VGND 0.02189f
C10653 VPWR.n56 VGND 0.06768f
C10654 VPWR.t1354 VGND 0.06817f
C10655 VPWR.t1361 VGND 0.02464f
C10656 VPWR.t1355 VGND 0.02189f
C10657 VPWR.n57 VGND 0.06768f
C10658 VPWR.n58 VGND 0.02542f
C10659 VPWR.n59 VGND 0.10289f
C10660 VPWR.n60 VGND 0.10289f
C10661 VPWR.n61 VGND 0.02542f
C10662 VPWR.t1342 VGND 0.02464f
C10663 VPWR.t1715 VGND 0.02189f
C10664 VPWR.n62 VGND 0.06768f
C10665 VPWR.t1581 VGND 0.06817f
C10666 VPWR.t1492 VGND 0.02464f
C10667 VPWR.t1582 VGND 0.02189f
C10668 VPWR.n63 VGND 0.06768f
C10669 VPWR.n64 VGND 0.02542f
C10670 VPWR.n65 VGND 0.10289f
C10671 VPWR.n66 VGND 0.10289f
C10672 VPWR.n67 VGND 0.02542f
C10673 VPWR.t1462 VGND 0.02464f
C10674 VPWR.t1454 VGND 0.02189f
C10675 VPWR.n68 VGND 0.06768f
C10676 VPWR.t1435 VGND 0.06817f
C10677 VPWR.t1718 VGND 0.02464f
C10678 VPWR.t1436 VGND 0.02189f
C10679 VPWR.n69 VGND 0.06768f
C10680 VPWR.n70 VGND 0.02542f
C10681 VPWR.n71 VGND 0.10289f
C10682 VPWR.n72 VGND 0.10289f
C10683 VPWR.n73 VGND 0.02542f
C10684 VPWR.t1588 VGND 0.02464f
C10685 VPWR.t1669 VGND 0.02189f
C10686 VPWR.n74 VGND 0.06768f
C10687 VPWR.t1558 VGND 0.06817f
C10688 VPWR.t1572 VGND 0.02464f
C10689 VPWR.t1559 VGND 0.02189f
C10690 VPWR.n75 VGND 0.06768f
C10691 VPWR.n76 VGND 0.02542f
C10692 VPWR.n77 VGND 0.10289f
C10693 VPWR.n78 VGND 0.10289f
C10694 VPWR.n79 VGND 0.02542f
C10695 VPWR.t1412 VGND 0.02464f
C10696 VPWR.t1431 VGND 0.02189f
C10697 VPWR.n80 VGND 0.06768f
C10698 VPWR.t1395 VGND 0.06817f
C10699 VPWR.t1691 VGND 0.02464f
C10700 VPWR.t1396 VGND 0.02189f
C10701 VPWR.n81 VGND 0.06768f
C10702 VPWR.n82 VGND 0.02542f
C10703 VPWR.n83 VGND 0.10289f
C10704 VPWR.n84 VGND 0.10289f
C10705 VPWR.n85 VGND 0.02542f
C10706 VPWR.t1535 VGND 0.02464f
C10707 VPWR.t1672 VGND 0.02189f
C10708 VPWR.n86 VGND 0.06768f
C10709 VPWR.t1516 VGND 0.06817f
C10710 VPWR.t1526 VGND 0.02464f
C10711 VPWR.t1517 VGND 0.02189f
C10712 VPWR.n87 VGND 0.06768f
C10713 VPWR.n88 VGND 0.02542f
C10714 VPWR.n89 VGND 0.10289f
C10715 VPWR.n90 VGND 0.10289f
C10716 VPWR.n91 VGND 0.02542f
C10717 VPWR.t1415 VGND 0.02464f
C10718 VPWR.t1409 VGND 0.02189f
C10719 VPWR.n92 VGND 0.06768f
C10720 VPWR.t1646 VGND 0.06817f
C10721 VPWR.t1650 VGND 0.02464f
C10722 VPWR.t1647 VGND 0.02189f
C10723 VPWR.n93 VGND 0.06768f
C10724 VPWR.n94 VGND 0.02542f
C10725 VPWR.n95 VGND 0.10289f
C10726 VPWR.n96 VGND 0.10289f
C10727 VPWR.n97 VGND 0.02542f
C10728 VPWR.t1538 VGND 0.02464f
C10729 VPWR.t1629 VGND 0.02189f
C10730 VPWR.n98 VGND 0.06768f
C10731 VPWR.t1392 VGND 0.10732f
C10732 VPWR.t1368 VGND 0.05805f
C10733 VPWR.t1499 VGND 0.06817f
C10734 VPWR.t1393 VGND 0.02464f
C10735 VPWR.t1500 VGND 0.02189f
C10736 VPWR.n99 VGND 0.06768f
C10737 VPWR.n100 VGND 0.02213f
C10738 VPWR.n101 VGND 0.02429f
C10739 VPWR.n103 VGND 0.01347f
C10740 VPWR.n104 VGND 0.02213f
C10741 VPWR.n105 VGND 0.02429f
C10742 VPWR.n106 VGND 0.02304f
C10743 VPWR.n107 VGND 0.01456f
C10744 VPWR.n108 VGND 0.02047f
C10745 VPWR.n109 VGND 0.02084f
C10746 VPWR.n110 VGND 0.01313f
C10747 VPWR.n112 VGND 0.01347f
C10748 VPWR.n113 VGND 0.01963f
C10749 VPWR.n114 VGND 0.02213f
C10750 VPWR.n115 VGND 0.02429f
C10751 VPWR.n116 VGND 0.02304f
C10752 VPWR.n117 VGND 0.02731f
C10753 VPWR.n119 VGND 0.02047f
C10754 VPWR.n120 VGND 0.02084f
C10755 VPWR.n121 VGND 0.01313f
C10756 VPWR.n123 VGND 0.01347f
C10757 VPWR.n124 VGND 0.01879f
C10758 VPWR.n125 VGND 0.02213f
C10759 VPWR.n126 VGND 0.02429f
C10760 VPWR.n127 VGND 0.02304f
C10761 VPWR.n128 VGND 0.02731f
C10762 VPWR.n130 VGND 0.02047f
C10763 VPWR.n131 VGND 0.02084f
C10764 VPWR.n132 VGND 0.01313f
C10765 VPWR.n134 VGND 0.01347f
C10766 VPWR.n135 VGND 0.01763f
C10767 VPWR.n136 VGND 0.1565f
C10768 VPWR.n137 VGND 0.02213f
C10769 VPWR.n138 VGND 0.02429f
C10770 VPWR.n139 VGND 0.02304f
C10771 VPWR.n140 VGND 0.02731f
C10772 VPWR.n142 VGND 0.02047f
C10773 VPWR.n143 VGND 0.02084f
C10774 VPWR.n144 VGND 0.01313f
C10775 VPWR.n146 VGND 0.01347f
C10776 VPWR.n147 VGND 0.01763f
C10777 VPWR.n148 VGND 0.13004f
C10778 VPWR.n149 VGND 0.02213f
C10779 VPWR.n150 VGND 0.02429f
C10780 VPWR.n151 VGND 0.02304f
C10781 VPWR.n152 VGND 0.02731f
C10782 VPWR.n154 VGND 0.02047f
C10783 VPWR.n155 VGND 0.02084f
C10784 VPWR.n156 VGND 0.01313f
C10785 VPWR.n158 VGND 0.01347f
C10786 VPWR.n159 VGND 0.01763f
C10787 VPWR.n160 VGND 0.13004f
C10788 VPWR.n161 VGND 0.02213f
C10789 VPWR.n162 VGND 0.02429f
C10790 VPWR.n163 VGND 0.02304f
C10791 VPWR.n164 VGND 0.02731f
C10792 VPWR.n166 VGND 0.02047f
C10793 VPWR.n167 VGND 0.02084f
C10794 VPWR.n168 VGND 0.01313f
C10795 VPWR.n170 VGND 0.01347f
C10796 VPWR.n171 VGND 0.01763f
C10797 VPWR.n172 VGND 0.13004f
C10798 VPWR.n173 VGND 0.02213f
C10799 VPWR.n174 VGND 0.02429f
C10800 VPWR.n175 VGND 0.02304f
C10801 VPWR.n176 VGND 0.02731f
C10802 VPWR.n178 VGND 0.02047f
C10803 VPWR.n179 VGND 0.02084f
C10804 VPWR.n180 VGND 0.01313f
C10805 VPWR.n182 VGND 0.01347f
C10806 VPWR.n183 VGND 0.01763f
C10807 VPWR.n184 VGND 0.13004f
C10808 VPWR.n185 VGND 0.02213f
C10809 VPWR.n186 VGND 0.02429f
C10810 VPWR.n187 VGND 0.02304f
C10811 VPWR.n188 VGND 0.02731f
C10812 VPWR.n190 VGND 0.02047f
C10813 VPWR.n191 VGND 0.02084f
C10814 VPWR.n192 VGND 0.01313f
C10815 VPWR.n194 VGND 0.01347f
C10816 VPWR.n195 VGND 0.01763f
C10817 VPWR.n196 VGND 0.13004f
C10818 VPWR.n197 VGND 0.02213f
C10819 VPWR.n198 VGND 0.02429f
C10820 VPWR.n199 VGND 0.02304f
C10821 VPWR.n200 VGND 0.02731f
C10822 VPWR.n202 VGND 0.02047f
C10823 VPWR.n203 VGND 0.02084f
C10824 VPWR.n204 VGND 0.01313f
C10825 VPWR.n206 VGND 0.01347f
C10826 VPWR.n207 VGND 0.01763f
C10827 VPWR.n208 VGND 0.13004f
C10828 VPWR.n209 VGND 0.02213f
C10829 VPWR.n210 VGND 0.02429f
C10830 VPWR.n211 VGND 0.02304f
C10831 VPWR.n212 VGND 0.02731f
C10832 VPWR.n214 VGND 0.02047f
C10833 VPWR.n215 VGND 0.02084f
C10834 VPWR.n216 VGND 0.01313f
C10835 VPWR.n218 VGND 0.01347f
C10836 VPWR.n219 VGND 0.01763f
C10837 VPWR.n220 VGND 0.13004f
C10838 VPWR.n221 VGND 0.02213f
C10839 VPWR.n222 VGND 0.02429f
C10840 VPWR.n223 VGND 0.02304f
C10841 VPWR.n224 VGND 0.02731f
C10842 VPWR.n226 VGND 0.02047f
C10843 VPWR.n227 VGND 0.02084f
C10844 VPWR.n228 VGND 0.01313f
C10845 VPWR.n230 VGND 0.01347f
C10846 VPWR.n231 VGND 0.01763f
C10847 VPWR.n232 VGND 0.13004f
C10848 VPWR.n233 VGND 0.02213f
C10849 VPWR.n234 VGND 0.02429f
C10850 VPWR.n235 VGND 0.02304f
C10851 VPWR.n236 VGND 0.02731f
C10852 VPWR.n238 VGND 0.02047f
C10853 VPWR.n239 VGND 0.02084f
C10854 VPWR.n240 VGND 0.01313f
C10855 VPWR.n242 VGND 0.01347f
C10856 VPWR.n243 VGND 0.01763f
C10857 VPWR.n244 VGND 0.13004f
C10858 VPWR.n245 VGND 0.02213f
C10859 VPWR.n246 VGND 0.02429f
C10860 VPWR.n247 VGND 0.02304f
C10861 VPWR.n248 VGND 0.02731f
C10862 VPWR.n250 VGND 0.02047f
C10863 VPWR.n251 VGND 0.02084f
C10864 VPWR.n252 VGND 0.01313f
C10865 VPWR.n254 VGND 0.01347f
C10866 VPWR.n255 VGND 0.01763f
C10867 VPWR.n256 VGND 0.13004f
C10868 VPWR.n257 VGND 0.02213f
C10869 VPWR.n258 VGND 0.02429f
C10870 VPWR.n259 VGND 0.02304f
C10871 VPWR.n260 VGND 0.02731f
C10872 VPWR.n262 VGND 0.02047f
C10873 VPWR.n263 VGND 0.02084f
C10874 VPWR.n264 VGND 0.01313f
C10875 VPWR.n266 VGND 0.01347f
C10876 VPWR.n267 VGND 0.01763f
C10877 VPWR.n268 VGND 0.13004f
C10878 VPWR.n269 VGND 0.02213f
C10879 VPWR.n270 VGND 0.02429f
C10880 VPWR.n271 VGND 0.02304f
C10881 VPWR.n272 VGND 0.02731f
C10882 VPWR.n274 VGND 0.02047f
C10883 VPWR.n275 VGND 0.02084f
C10884 VPWR.n276 VGND 0.01313f
C10885 VPWR.n278 VGND 0.01347f
C10886 VPWR.n279 VGND 0.01763f
C10887 VPWR.n280 VGND 0.13004f
C10888 VPWR.n281 VGND 0.17544f
C10889 VPWR.n282 VGND 0.01763f
C10890 VPWR.n283 VGND 0.01313f
C10891 VPWR.n284 VGND 0.02047f
C10892 VPWR.n285 VGND 0.02084f
C10893 VPWR.n287 VGND 0.02304f
C10894 VPWR.n288 VGND 0.02731f
C10895 VPWR.n289 VGND 0.02542f
C10896 VPWR.t1062 VGND 0.02464f
C10897 VPWR.t904 VGND 0.02189f
C10898 VPWR.n290 VGND 0.06768f
C10899 VPWR.t1061 VGND 0.10732f
C10900 VPWR.t676 VGND 0.05805f
C10901 VPWR.t903 VGND 0.06817f
C10902 VPWR.t880 VGND 0.02464f
C10903 VPWR.t1699 VGND 0.02189f
C10904 VPWR.n291 VGND 0.06768f
C10905 VPWR.n292 VGND 0.01329f
C10906 VPWR.n293 VGND 0.05634f
C10907 VPWR.t1698 VGND 0.0986f
C10908 VPWR.t1879 VGND 0.05805f
C10909 VPWR.t879 VGND 0.08842f
C10910 VPWR.t19 VGND 0.02464f
C10911 VPWR.t196 VGND 0.02189f
C10912 VPWR.n294 VGND 0.06768f
C10913 VPWR.n295 VGND 0.01329f
C10914 VPWR.n297 VGND 0.08003f
C10915 VPWR.t195 VGND 0.06817f
C10916 VPWR.t1882 VGND 0.05805f
C10917 VPWR.t18 VGND 0.08842f
C10918 VPWR.t1245 VGND 0.02464f
C10919 VPWR.t1789 VGND 0.02189f
C10920 VPWR.n298 VGND 0.06768f
C10921 VPWR.n299 VGND 0.01329f
C10922 VPWR.n301 VGND 0.08003f
C10923 VPWR.t1788 VGND 0.06817f
C10924 VPWR.t1873 VGND 0.05805f
C10925 VPWR.t1244 VGND 0.08842f
C10926 VPWR.t99 VGND 0.02464f
C10927 VPWR.t970 VGND 0.02189f
C10928 VPWR.n302 VGND 0.06768f
C10929 VPWR.n303 VGND 0.01329f
C10930 VPWR.n305 VGND 0.08003f
C10931 VPWR.t969 VGND 0.06817f
C10932 VPWR.t1874 VGND 0.05805f
C10933 VPWR.t98 VGND 0.08842f
C10934 VPWR.t522 VGND 0.02464f
C10935 VPWR.t1803 VGND 0.02189f
C10936 VPWR.n306 VGND 0.06768f
C10937 VPWR.n307 VGND 0.01329f
C10938 VPWR.n309 VGND 0.08003f
C10939 VPWR.t1802 VGND 0.06817f
C10940 VPWR.t677 VGND 0.05805f
C10941 VPWR.t521 VGND 0.08842f
C10942 VPWR.t358 VGND 0.02464f
C10943 VPWR.t528 VGND 0.02189f
C10944 VPWR.n310 VGND 0.06768f
C10945 VPWR.n311 VGND 0.01329f
C10946 VPWR.n313 VGND 0.08003f
C10947 VPWR.t527 VGND 0.06817f
C10948 VPWR.t678 VGND 0.05805f
C10949 VPWR.t357 VGND 0.08842f
C10950 VPWR.t729 VGND 0.02464f
C10951 VPWR.t368 VGND 0.02189f
C10952 VPWR.n314 VGND 0.06768f
C10953 VPWR.n315 VGND 0.01329f
C10954 VPWR.n317 VGND 0.08003f
C10955 VPWR.t367 VGND 0.06817f
C10956 VPWR.t1877 VGND 0.05805f
C10957 VPWR.t728 VGND 0.08842f
C10958 VPWR.t70 VGND 0.02464f
C10959 VPWR.t1897 VGND 0.02189f
C10960 VPWR.n318 VGND 0.06768f
C10961 VPWR.n319 VGND 0.01329f
C10962 VPWR.n321 VGND 0.08003f
C10963 VPWR.t1896 VGND 0.06817f
C10964 VPWR.t673 VGND 0.05805f
C10965 VPWR.t69 VGND 0.08842f
C10966 VPWR.t1733 VGND 0.02464f
C10967 VPWR.t848 VGND 0.02189f
C10968 VPWR.n322 VGND 0.06768f
C10969 VPWR.n323 VGND 0.01329f
C10970 VPWR.n325 VGND 0.08003f
C10971 VPWR.t847 VGND 0.06817f
C10972 VPWR.t674 VGND 0.05805f
C10973 VPWR.t1732 VGND 0.08842f
C10974 VPWR.t1819 VGND 0.02464f
C10975 VPWR.t1739 VGND 0.02189f
C10976 VPWR.n326 VGND 0.06768f
C10977 VPWR.n327 VGND 0.01329f
C10978 VPWR.n329 VGND 0.08003f
C10979 VPWR.t1738 VGND 0.06817f
C10980 VPWR.t1875 VGND 0.05805f
C10981 VPWR.t1818 VGND 0.08842f
C10982 VPWR.t655 VGND 0.02464f
C10983 VPWR.t1755 VGND 0.02189f
C10984 VPWR.n330 VGND 0.06768f
C10985 VPWR.n331 VGND 0.01329f
C10986 VPWR.n333 VGND 0.08003f
C10987 VPWR.t1754 VGND 0.06817f
C10988 VPWR.t1876 VGND 0.05805f
C10989 VPWR.t654 VGND 0.08842f
C10990 VPWR.t682 VGND 0.02464f
C10991 VPWR.t661 VGND 0.02189f
C10992 VPWR.n334 VGND 0.06768f
C10993 VPWR.n335 VGND 0.01329f
C10994 VPWR.n337 VGND 0.08003f
C10995 VPWR.t660 VGND 0.06817f
C10996 VPWR.t675 VGND 0.05805f
C10997 VPWR.t681 VGND 0.08842f
C10998 VPWR.t802 VGND 0.02464f
C10999 VPWR.t1034 VGND 0.02189f
C11000 VPWR.n338 VGND 0.06768f
C11001 VPWR.n339 VGND 0.01329f
C11002 VPWR.n341 VGND 0.08003f
C11003 VPWR.t1033 VGND 0.06817f
C11004 VPWR.t1880 VGND 0.05805f
C11005 VPWR.t801 VGND 0.08842f
C11006 VPWR.t1231 VGND 0.02464f
C11007 VPWR.t778 VGND 0.02189f
C11008 VPWR.n342 VGND 0.06768f
C11009 VPWR.n343 VGND 0.01329f
C11010 VPWR.n345 VGND 0.08003f
C11011 VPWR.t777 VGND 0.06817f
C11012 VPWR.t1881 VGND 0.05805f
C11013 VPWR.t1230 VGND 0.08842f
C11014 VPWR.t1023 VGND 0.02464f
C11015 VPWR.t1211 VGND 0.02189f
C11016 VPWR.n346 VGND 0.06768f
C11017 VPWR.n347 VGND 0.01329f
C11018 VPWR.n349 VGND 0.08003f
C11019 VPWR.t1210 VGND 0.06817f
C11020 VPWR.t1878 VGND 0.05805f
C11021 VPWR.t1022 VGND 0.08842f
C11022 VPWR.n350 VGND 0.08003f
C11023 VPWR.n352 VGND 0.01329f
C11024 VPWR.n353 VGND 0.10289f
C11025 VPWR.n354 VGND 0.74646f
C11026 VPWR.n355 VGND 0.10289f
C11027 VPWR.t1056 VGND 0.02464f
C11028 VPWR.t894 VGND 0.02189f
C11029 VPWR.n356 VGND 0.06768f
C11030 VPWR.t1055 VGND 0.10732f
C11031 VPWR.t1921 VGND 0.05805f
C11032 VPWR.t893 VGND 0.06817f
C11033 VPWR.t1214 VGND 0.08842f
C11034 VPWR.t900 VGND 0.02464f
C11035 VPWR.t1140 VGND 0.02189f
C11036 VPWR.n357 VGND 0.06768f
C11037 VPWR.n358 VGND 0.10289f
C11038 VPWR.n359 VGND 0.10289f
C11039 VPWR.t1215 VGND 0.02464f
C11040 VPWR.t770 VGND 0.02189f
C11041 VPWR.n360 VGND 0.06768f
C11042 VPWR.t940 VGND 0.05805f
C11043 VPWR.t769 VGND 0.06817f
C11044 VPWR.t632 VGND 0.08842f
C11045 VPWR.t794 VGND 0.02464f
C11046 VPWR.t1046 VGND 0.02189f
C11047 VPWR.n361 VGND 0.06768f
C11048 VPWR.n362 VGND 0.10289f
C11049 VPWR.n363 VGND 0.10289f
C11050 VPWR.t633 VGND 0.02464f
C11051 VPWR.t408 VGND 0.02189f
C11052 VPWR.n364 VGND 0.06768f
C11053 VPWR.t1920 VGND 0.05805f
C11054 VPWR.t407 VGND 0.06817f
C11055 VPWR.t1758 VGND 0.08842f
C11056 VPWR.t402 VGND 0.02464f
C11057 VPWR.t696 VGND 0.02189f
C11058 VPWR.n365 VGND 0.06768f
C11059 VPWR.n366 VGND 0.10289f
C11060 VPWR.n367 VGND 0.10289f
C11061 VPWR.t1759 VGND 0.02464f
C11062 VPWR.t1749 VGND 0.02189f
C11063 VPWR.n368 VGND 0.06768f
C11064 VPWR.t458 VGND 0.05805f
C11065 VPWR.t1748 VGND 0.06817f
C11066 VPWR.t569 VGND 0.08842f
C11067 VPWR.t1743 VGND 0.02464f
C11068 VPWR.t289 VGND 0.02189f
C11069 VPWR.n369 VGND 0.06768f
C11070 VPWR.n370 VGND 0.10289f
C11071 VPWR.n371 VGND 0.10289f
C11072 VPWR.t570 VGND 0.02464f
C11073 VPWR.t1106 VGND 0.02189f
C11074 VPWR.n372 VGND 0.06768f
C11075 VPWR.t1182 VGND 0.05805f
C11076 VPWR.t1105 VGND 0.06817f
C11077 VPWR.t363 VGND 0.08842f
C11078 VPWR.t1901 VGND 0.02464f
C11079 VPWR.t386 VGND 0.02189f
C11080 VPWR.n373 VGND 0.06768f
C11081 VPWR.n374 VGND 0.10289f
C11082 VPWR.n375 VGND 0.10289f
C11083 VPWR.t364 VGND 0.02464f
C11084 VPWR.t219 VGND 0.02189f
C11085 VPWR.n376 VGND 0.06768f
C11086 VPWR.t1923 VGND 0.05805f
C11087 VPWR.t218 VGND 0.06817f
C11088 VPWR.t1798 VGND 0.08842f
C11089 VPWR.t532 VGND 0.02464f
C11090 VPWR.t1158 VGND 0.02189f
C11091 VPWR.n377 VGND 0.06768f
C11092 VPWR.n378 VGND 0.10289f
C11093 VPWR.n379 VGND 0.10289f
C11094 VPWR.t1799 VGND 0.02464f
C11095 VPWR.t540 VGND 0.02189f
C11096 VPWR.n380 VGND 0.06768f
C11097 VPWR.t457 VGND 0.05805f
C11098 VPWR.t539 VGND 0.06817f
C11099 VPWR.t1784 VGND 0.08842f
C11100 VPWR.t1251 VGND 0.02464f
C11101 VPWR.t1025 VGND 0.02189f
C11102 VPWR.n381 VGND 0.06768f
C11103 VPWR.n382 VGND 0.10289f
C11104 VPWR.n383 VGND 0.10289f
C11105 VPWR.t1785 VGND 0.02464f
C11106 VPWR.t208 VGND 0.02189f
C11107 VPWR.n384 VGND 0.06768f
C11108 VPWR.t941 VGND 0.05805f
C11109 VPWR.t207 VGND 0.06817f
C11110 VPWR.t1009 VGND 0.02464f
C11111 VPWR.t1659 VGND 0.02189f
C11112 VPWR.n385 VGND 0.06768f
C11113 VPWR.t872 VGND 0.02464f
C11114 VPWR.t1377 VGND 0.02189f
C11115 VPWR.n386 VGND 0.06768f
C11116 VPWR.t1065 VGND 0.10732f
C11117 VPWR.t1269 VGND 0.05805f
C11118 VPWR.t1018 VGND 0.06817f
C11119 VPWR.t1066 VGND 0.02464f
C11120 VPWR.t1019 VGND 0.02189f
C11121 VPWR.n387 VGND 0.06768f
C11122 VPWR.n388 VGND 0.01329f
C11123 VPWR.n390 VGND 0.08003f
C11124 VPWR.t483 VGND 0.08842f
C11125 VPWR.t1925 VGND 0.05805f
C11126 VPWR.t145 VGND 0.06817f
C11127 VPWR.t484 VGND 0.02464f
C11128 VPWR.t146 VGND 0.02189f
C11129 VPWR.n391 VGND 0.06768f
C11130 VPWR.n392 VGND 0.01329f
C11131 VPWR.n394 VGND 0.08003f
C11132 VPWR.t513 VGND 0.08842f
C11133 VPWR.t1273 VGND 0.05805f
C11134 VPWR.t787 VGND 0.06817f
C11135 VPWR.t514 VGND 0.02464f
C11136 VPWR.t788 VGND 0.02189f
C11137 VPWR.n395 VGND 0.06768f
C11138 VPWR.n396 VGND 0.01329f
C11139 VPWR.n398 VGND 0.08003f
C11140 VPWR.t813 VGND 0.08842f
C11141 VPWR.t1272 VGND 0.05805f
C11142 VPWR.t636 VGND 0.06817f
C11143 VPWR.t814 VGND 0.02464f
C11144 VPWR.t637 VGND 0.02189f
C11145 VPWR.n399 VGND 0.06768f
C11146 VPWR.n400 VGND 0.01329f
C11147 VPWR.n402 VGND 0.08003f
C11148 VPWR.t1334 VGND 0.08842f
C11149 VPWR.t949 VGND 0.05805f
C11150 VPWR.t722 VGND 0.06817f
C11151 VPWR.t1335 VGND 0.02464f
C11152 VPWR.t723 VGND 0.02189f
C11153 VPWR.n403 VGND 0.06768f
C11154 VPWR.n404 VGND 0.01329f
C11155 VPWR.n406 VGND 0.08003f
C11156 VPWR.t1204 VGND 0.08842f
C11157 VPWR.t1278 VGND 0.05805f
C11158 VPWR.t1814 VGND 0.06817f
C11159 VPWR.t1205 VGND 0.02464f
C11160 VPWR.t1815 VGND 0.02189f
C11161 VPWR.n407 VGND 0.06768f
C11162 VPWR.n408 VGND 0.01329f
C11163 VPWR.n410 VGND 0.08003f
C11164 VPWR.t61 VGND 0.08842f
C11165 VPWR.t1277 VGND 0.05805f
C11166 VPWR.t1871 VGND 0.06817f
C11167 VPWR.t62 VGND 0.02464f
C11168 VPWR.t1872 VGND 0.02189f
C11169 VPWR.n411 VGND 0.06768f
C11170 VPWR.n412 VGND 0.01329f
C11171 VPWR.n414 VGND 0.08003f
C11172 VPWR.t1865 VGND 0.08842f
C11173 VPWR.t948 VGND 0.05805f
C11174 VPWR.t575 VGND 0.06817f
C11175 VPWR.t1866 VGND 0.02464f
C11176 VPWR.t576 VGND 0.02189f
C11177 VPWR.n415 VGND 0.06768f
C11178 VPWR.n416 VGND 0.01329f
C11179 VPWR.n418 VGND 0.08003f
C11180 VPWR.t599 VGND 0.08842f
C11181 VPWR.t947 VGND 0.05805f
C11182 VPWR.t724 VGND 0.06817f
C11183 VPWR.t600 VGND 0.02464f
C11184 VPWR.t725 VGND 0.02189f
C11185 VPWR.n419 VGND 0.06768f
C11186 VPWR.n420 VGND 0.01329f
C11187 VPWR.n422 VGND 0.08003f
C11188 VPWR.t1222 VGND 0.08842f
C11189 VPWR.t951 VGND 0.05805f
C11190 VPWR.t346 VGND 0.06817f
C11191 VPWR.t1223 VGND 0.02464f
C11192 VPWR.t347 VGND 0.02189f
C11193 VPWR.n423 VGND 0.06768f
C11194 VPWR.n424 VGND 0.01329f
C11195 VPWR.n426 VGND 0.08003f
C11196 VPWR.t340 VGND 0.08842f
C11197 VPWR.t1271 VGND 0.05805f
C11198 VPWR.t1826 VGND 0.06817f
C11199 VPWR.t341 VGND 0.02464f
C11200 VPWR.t1827 VGND 0.02189f
C11201 VPWR.n427 VGND 0.06768f
C11202 VPWR.n428 VGND 0.01329f
C11203 VPWR.n430 VGND 0.08003f
C11204 VPWR.t1841 VGND 0.08842f
C11205 VPWR.t1270 VGND 0.05805f
C11206 VPWR.t1810 VGND 0.06817f
C11207 VPWR.t1842 VGND 0.02464f
C11208 VPWR.t1811 VGND 0.02189f
C11209 VPWR.n431 VGND 0.06768f
C11210 VPWR.n432 VGND 0.01329f
C11211 VPWR.n434 VGND 0.08003f
C11212 VPWR.t923 VGND 0.08842f
C11213 VPWR.t1276 VGND 0.05805f
C11214 VPWR.t944 VGND 0.06817f
C11215 VPWR.t924 VGND 0.02464f
C11216 VPWR.t945 VGND 0.02189f
C11217 VPWR.n435 VGND 0.06768f
C11218 VPWR.n436 VGND 0.01329f
C11219 VPWR.n438 VGND 0.08003f
C11220 VPWR.t1293 VGND 0.08842f
C11221 VPWR.t1275 VGND 0.05805f
C11222 VPWR.t14 VGND 0.06817f
C11223 VPWR.t1294 VGND 0.02464f
C11224 VPWR.t15 VGND 0.02189f
C11225 VPWR.n439 VGND 0.06768f
C11226 VPWR.n440 VGND 0.01329f
C11227 VPWR.n442 VGND 0.08003f
C11228 VPWR.t8 VGND 0.08842f
C11229 VPWR.t1274 VGND 0.05805f
C11230 VPWR.t1012 VGND 0.06817f
C11231 VPWR.t9 VGND 0.02464f
C11232 VPWR.t1013 VGND 0.02189f
C11233 VPWR.n443 VGND 0.06768f
C11234 VPWR.n444 VGND 0.01329f
C11235 VPWR.n446 VGND 0.08003f
C11236 VPWR.t871 VGND 0.08842f
C11237 VPWR.t946 VGND 0.05805f
C11238 VPWR.t1376 VGND 0.0986f
C11239 VPWR.n447 VGND 0.05634f
C11240 VPWR.n448 VGND 0.01329f
C11241 VPWR.n449 VGND 0.10289f
C11242 VPWR.n450 VGND 0.75117f
C11243 VPWR.n451 VGND 0.10289f
C11244 VPWR.t182 VGND 0.02464f
C11245 VPWR.t1489 VGND 0.02189f
C11246 VPWR.n452 VGND 0.06768f
C11247 VPWR.t873 VGND 0.06817f
C11248 VPWR.t884 VGND 0.02464f
C11249 VPWR.t874 VGND 0.02189f
C11250 VPWR.n453 VGND 0.06768f
C11251 VPWR.n454 VGND 0.10289f
C11252 VPWR.n455 VGND 0.10289f
C11253 VPWR.t546 VGND 0.02464f
C11254 VPWR.t892 VGND 0.02189f
C11255 VPWR.n456 VGND 0.06768f
C11256 VPWR.t1238 VGND 0.06817f
C11257 VPWR.t1781 VGND 0.02464f
C11258 VPWR.t1239 VGND 0.02189f
C11259 VPWR.n457 VGND 0.06768f
C11260 VPWR.n458 VGND 0.10289f
C11261 VPWR.n459 VGND 0.10289f
C11262 VPWR.t1915 VGND 0.02464f
C11263 VPWR.t95 VGND 0.02189f
C11264 VPWR.n460 VGND 0.06768f
C11265 VPWR.t1918 VGND 0.06817f
C11266 VPWR.t432 VGND 0.02464f
C11267 VPWR.t1919 VGND 0.02189f
C11268 VPWR.n461 VGND 0.06768f
C11269 VPWR.n462 VGND 0.10289f
C11270 VPWR.n463 VGND 0.10289f
C11271 VPWR.t580 VGND 0.02464f
C11272 VPWR.t440 VGND 0.02189f
C11273 VPWR.n464 VGND 0.06768f
C11274 VPWR.t853 VGND 0.06817f
C11275 VPWR.t737 VGND 0.02464f
C11276 VPWR.t854 VGND 0.02189f
C11277 VPWR.n465 VGND 0.06768f
C11278 VPWR.n466 VGND 0.10289f
C11279 VPWR.n467 VGND 0.10289f
C11280 VPWR.t1257 VGND 0.02464f
C11281 VPWR.t604 VGND 0.02189f
C11282 VPWR.n468 VGND 0.06768f
C11283 VPWR.t1260 VGND 0.06817f
C11284 VPWR.t1177 VGND 0.02464f
C11285 VPWR.t1261 VGND 0.02189f
C11286 VPWR.n469 VGND 0.06768f
C11287 VPWR.n470 VGND 0.10289f
C11288 VPWR.n471 VGND 0.10289f
C11289 VPWR.t1122 VGND 0.02464f
C11290 VPWR.t1162 VGND 0.02189f
C11291 VPWR.n472 VGND 0.06768f
C11292 VPWR.t1125 VGND 0.06817f
C11293 VPWR.t154 VGND 0.02464f
C11294 VPWR.t1126 VGND 0.02189f
C11295 VPWR.n473 VGND 0.06768f
C11296 VPWR.n474 VGND 0.10289f
C11297 VPWR.n475 VGND 0.10289f
C11298 VPWR.t828 VGND 0.02464f
C11299 VPWR.t1337 VGND 0.02189f
C11300 VPWR.n476 VGND 0.06768f
C11301 VPWR.t805 VGND 0.06817f
C11302 VPWR.t1130 VGND 0.02464f
C11303 VPWR.t806 VGND 0.02189f
C11304 VPWR.n477 VGND 0.06768f
C11305 VPWR.n478 VGND 0.10289f
C11306 VPWR.n479 VGND 0.10289f
C11307 VPWR.t958 VGND 0.02464f
C11308 VPWR.t1134 VGND 0.02189f
C11309 VPWR.n480 VGND 0.06768f
C11310 VPWR.t1074 VGND 0.10732f
C11311 VPWR.t1268 VGND 0.05805f
C11312 VPWR.t1726 VGND 0.06817f
C11313 VPWR.t1075 VGND 0.02464f
C11314 VPWR.t1727 VGND 0.02189f
C11315 VPWR.n481 VGND 0.06768f
C11316 VPWR.t1064 VGND 0.02464f
C11317 VPWR.t902 VGND 0.02189f
C11318 VPWR.n482 VGND 0.06768f
C11319 VPWR.t1063 VGND 0.10732f
C11320 VPWR.t86 VGND 0.05805f
C11321 VPWR.t901 VGND 0.06817f
C11322 VPWR.t878 VGND 0.02464f
C11323 VPWR.t1707 VGND 0.02189f
C11324 VPWR.n483 VGND 0.06768f
C11325 VPWR.n484 VGND 0.01329f
C11326 VPWR.n485 VGND 0.05634f
C11327 VPWR.t1706 VGND 0.0986f
C11328 VPWR.t672 VGND 0.05805f
C11329 VPWR.t877 VGND 0.08842f
C11330 VPWR.t17 VGND 0.02464f
C11331 VPWR.t1015 VGND 0.02189f
C11332 VPWR.n486 VGND 0.06768f
C11333 VPWR.n487 VGND 0.01329f
C11334 VPWR.n489 VGND 0.08003f
C11335 VPWR.t1014 VGND 0.06817f
C11336 VPWR.t79 VGND 0.05805f
C11337 VPWR.t16 VGND 0.08842f
C11338 VPWR.t1241 VGND 0.02464f
C11339 VPWR.t1787 VGND 0.02189f
C11340 VPWR.n490 VGND 0.06768f
C11341 VPWR.n491 VGND 0.01329f
C11342 VPWR.n493 VGND 0.08003f
C11343 VPWR.t1786 VGND 0.06817f
C11344 VPWR.t1848 VGND 0.05805f
C11345 VPWR.t1240 VGND 0.08842f
C11346 VPWR.t97 VGND 0.02464f
C11347 VPWR.t966 VGND 0.02189f
C11348 VPWR.n494 VGND 0.06768f
C11349 VPWR.n495 VGND 0.01329f
C11350 VPWR.n497 VGND 0.08003f
C11351 VPWR.t965 VGND 0.06817f
C11352 VPWR.t1849 VGND 0.05805f
C11353 VPWR.t96 VGND 0.08842f
C11354 VPWR.t1829 VGND 0.02464f
C11355 VPWR.t1801 VGND 0.02189f
C11356 VPWR.n498 VGND 0.06768f
C11357 VPWR.n499 VGND 0.01329f
C11358 VPWR.n501 VGND 0.08003f
C11359 VPWR.t1800 VGND 0.06817f
C11360 VPWR.t75 VGND 0.05805f
C11361 VPWR.t1828 VGND 0.08842f
C11362 VPWR.t356 VGND 0.02464f
C11363 VPWR.t524 VGND 0.02189f
C11364 VPWR.n502 VGND 0.06768f
C11365 VPWR.n503 VGND 0.01329f
C11366 VPWR.n505 VGND 0.08003f
C11367 VPWR.t523 VGND 0.06817f
C11368 VPWR.t76 VGND 0.05805f
C11369 VPWR.t355 VGND 0.08842f
C11370 VPWR.t727 VGND 0.02464f
C11371 VPWR.t366 VGND 0.02189f
C11372 VPWR.n506 VGND 0.06768f
C11373 VPWR.n507 VGND 0.01329f
C11374 VPWR.n509 VGND 0.08003f
C11375 VPWR.t365 VGND 0.06817f
C11376 VPWR.t670 VGND 0.05805f
C11377 VPWR.t726 VGND 0.08842f
C11378 VPWR.t66 VGND 0.02464f
C11379 VPWR.t731 VGND 0.02189f
C11380 VPWR.n510 VGND 0.06768f
C11381 VPWR.n511 VGND 0.01329f
C11382 VPWR.n513 VGND 0.08003f
C11383 VPWR.t730 VGND 0.06817f
C11384 VPWR.t83 VGND 0.05805f
C11385 VPWR.t65 VGND 0.08842f
C11386 VPWR.t1731 VGND 0.02464f
C11387 VPWR.t844 VGND 0.02189f
C11388 VPWR.n514 VGND 0.06768f
C11389 VPWR.n515 VGND 0.01329f
C11390 VPWR.n517 VGND 0.08003f
C11391 VPWR.t843 VGND 0.06817f
C11392 VPWR.t84 VGND 0.05805f
C11393 VPWR.t1730 VGND 0.08842f
C11394 VPWR.t1817 VGND 0.02464f
C11395 VPWR.t1735 VGND 0.02189f
C11396 VPWR.n518 VGND 0.06768f
C11397 VPWR.n519 VGND 0.01329f
C11398 VPWR.n521 VGND 0.08003f
C11399 VPWR.t1734 VGND 0.06817f
C11400 VPWR.t1850 VGND 0.05805f
C11401 VPWR.t1816 VGND 0.08842f
C11402 VPWR.t113 VGND 0.02464f
C11403 VPWR.t1751 VGND 0.02189f
C11404 VPWR.n522 VGND 0.06768f
C11405 VPWR.n523 VGND 0.01329f
C11406 VPWR.n525 VGND 0.08003f
C11407 VPWR.t1750 VGND 0.06817f
C11408 VPWR.t1851 VGND 0.05805f
C11409 VPWR.t112 VGND 0.08842f
C11410 VPWR.t680 VGND 0.02464f
C11411 VPWR.t657 VGND 0.02189f
C11412 VPWR.n526 VGND 0.06768f
C11413 VPWR.n527 VGND 0.01329f
C11414 VPWR.n529 VGND 0.08003f
C11415 VPWR.t656 VGND 0.06817f
C11416 VPWR.t85 VGND 0.05805f
C11417 VPWR.t679 VGND 0.08842f
C11418 VPWR.t804 VGND 0.02464f
C11419 VPWR.t1032 VGND 0.02189f
C11420 VPWR.n530 VGND 0.06768f
C11421 VPWR.n531 VGND 0.01329f
C11422 VPWR.n533 VGND 0.08003f
C11423 VPWR.t1031 VGND 0.06817f
C11424 VPWR.t77 VGND 0.05805f
C11425 VPWR.t803 VGND 0.08842f
C11426 VPWR.t1229 VGND 0.02464f
C11427 VPWR.t780 VGND 0.02189f
C11428 VPWR.n534 VGND 0.06768f
C11429 VPWR.n535 VGND 0.01329f
C11430 VPWR.n537 VGND 0.08003f
C11431 VPWR.t779 VGND 0.06817f
C11432 VPWR.t78 VGND 0.05805f
C11433 VPWR.t1228 VGND 0.08842f
C11434 VPWR.t1021 VGND 0.02464f
C11435 VPWR.t1207 VGND 0.02189f
C11436 VPWR.n538 VGND 0.06768f
C11437 VPWR.n539 VGND 0.01329f
C11438 VPWR.n541 VGND 0.08003f
C11439 VPWR.t1206 VGND 0.06817f
C11440 VPWR.t671 VGND 0.05805f
C11441 VPWR.t1020 VGND 0.08842f
C11442 VPWR.n542 VGND 0.08003f
C11443 VPWR.n544 VGND 0.01329f
C11444 VPWR.n545 VGND 0.10289f
C11445 VPWR.n546 VGND 0.74646f
C11446 VPWR.n547 VGND 0.10289f
C11447 VPWR.t1050 VGND 0.02464f
C11448 VPWR.t619 VGND 0.02189f
C11449 VPWR.n548 VGND 0.06768f
C11450 VPWR.t1049 VGND 0.10732f
C11451 VPWR.t1001 VGND 0.05805f
C11452 VPWR.t618 VGND 0.06817f
C11453 VPWR.t259 VGND 0.08842f
C11454 VPWR.t1911 VGND 0.02464f
C11455 VPWR.t268 VGND 0.02189f
C11456 VPWR.n549 VGND 0.06768f
C11457 VPWR.n550 VGND 0.10289f
C11458 VPWR.n551 VGND 0.10289f
C11459 VPWR.t260 VGND 0.02464f
C11460 VPWR.t820 VGND 0.02189f
C11461 VPWR.n552 VGND 0.06768f
C11462 VPWR.t1776 VGND 0.05805f
C11463 VPWR.t819 VGND 0.06817f
C11464 VPWR.t1041 VGND 0.08842f
C11465 VPWR.t782 VGND 0.02464f
C11466 VPWR.t376 VGND 0.02189f
C11467 VPWR.n553 VGND 0.06768f
C11468 VPWR.n554 VGND 0.10289f
C11469 VPWR.n555 VGND 0.10289f
C11470 VPWR.t1042 VGND 0.02464f
C11471 VPWR.t1187 VGND 0.02189f
C11472 VPWR.n556 VGND 0.06768f
C11473 VPWR.t1000 VGND 0.05805f
C11474 VPWR.t1186 VGND 0.06817f
C11475 VPWR.t557 VGND 0.08842f
C11476 VPWR.t1321 VGND 0.02464f
C11477 VPWR.t1171 VGND 0.02189f
C11478 VPWR.n557 VGND 0.06768f
C11479 VPWR.n558 VGND 0.10289f
C11480 VPWR.n559 VGND 0.10289f
C11481 VPWR.t558 VGND 0.02464f
C11482 VPWR.t500 VGND 0.02189f
C11483 VPWR.n560 VGND 0.06768f
C11484 VPWR.t861 VGND 0.05805f
C11485 VPWR.t499 VGND 0.06817f
C11486 VPWR.t849 VGND 0.08842f
C11487 VPWR.t492 VGND 0.02464f
C11488 VPWR.t7 VGND 0.02189f
C11489 VPWR.n561 VGND 0.06768f
C11490 VPWR.n562 VGND 0.10289f
C11491 VPWR.n563 VGND 0.10289f
C11492 VPWR.t850 VGND 0.02464f
C11493 VPWR.t109 VGND 0.02189f
C11494 VPWR.n564 VGND 0.06768f
C11495 VPWR.t866 VGND 0.05805f
C11496 VPWR.t108 VGND 0.06817f
C11497 VPWR.t587 VGND 0.08842f
C11498 VPWR.t520 VGND 0.02464f
C11499 VPWR.t428 VGND 0.02189f
C11500 VPWR.n565 VGND 0.06768f
C11501 VPWR.n566 VGND 0.10289f
C11502 VPWR.n567 VGND 0.10289f
C11503 VPWR.t588 VGND 0.02464f
C11504 VPWR.t715 VGND 0.02189f
C11505 VPWR.n568 VGND 0.06768f
C11506 VPWR.t1774 VGND 0.05805f
C11507 VPWR.t714 VGND 0.06817f
C11508 VPWR.t1141 VGND 0.08842f
C11509 VPWR.t707 VGND 0.02464f
C11510 VPWR.t1150 VGND 0.02189f
C11511 VPWR.n569 VGND 0.06768f
C11512 VPWR.n570 VGND 0.10289f
C11513 VPWR.n571 VGND 0.10289f
C11514 VPWR.t1142 VGND 0.02464f
C11515 VPWR.t1286 VGND 0.02189f
C11516 VPWR.n572 VGND 0.06768f
C11517 VPWR.t860 VGND 0.05805f
C11518 VPWR.t1285 VGND 0.06817f
C11519 VPWR.t477 VGND 0.08842f
C11520 VPWR.t972 VGND 0.02464f
C11521 VPWR.t42 VGND 0.02189f
C11522 VPWR.n573 VGND 0.06768f
C11523 VPWR.n574 VGND 0.10289f
C11524 VPWR.n575 VGND 0.10289f
C11525 VPWR.t478 VGND 0.02464f
C11526 VPWR.t162 VGND 0.02189f
C11527 VPWR.n576 VGND 0.06768f
C11528 VPWR.t1777 VGND 0.05805f
C11529 VPWR.t161 VGND 0.06817f
C11530 VPWR.t204 VGND 0.02464f
C11531 VPWR.t1556 VGND 0.02189f
C11532 VPWR.n577 VGND 0.06768f
C11533 VPWR.t1005 VGND 0.02464f
C11534 VPWR.t1664 VGND 0.02189f
C11535 VPWR.n578 VGND 0.06768f
C11536 VPWR.t1057 VGND 0.10732f
C11537 VPWR.t352 VGND 0.05805f
C11538 VPWR.t907 VGND 0.06817f
C11539 VPWR.t1058 VGND 0.02464f
C11540 VPWR.t908 VGND 0.02189f
C11541 VPWR.n579 VGND 0.06768f
C11542 VPWR.n580 VGND 0.01329f
C11543 VPWR.n582 VGND 0.08003f
C11544 VPWR.t897 VGND 0.08842f
C11545 VPWR.t424 VGND 0.05805f
C11546 VPWR.t1137 VGND 0.06817f
C11547 VPWR.t898 VGND 0.02464f
C11548 VPWR.t1138 VGND 0.02189f
C11549 VPWR.n583 VGND 0.06768f
C11550 VPWR.n584 VGND 0.01329f
C11551 VPWR.n586 VGND 0.08003f
C11552 VPWR.t1212 VGND 0.08842f
C11553 VPWR.t328 VGND 0.05805f
C11554 VPWR.t771 VGND 0.06817f
C11555 VPWR.t1213 VGND 0.02464f
C11556 VPWR.t772 VGND 0.02189f
C11557 VPWR.n587 VGND 0.06768f
C11558 VPWR.n588 VGND 0.01329f
C11559 VPWR.n590 VGND 0.08003f
C11560 VPWR.t795 VGND 0.08842f
C11561 VPWR.t327 VGND 0.05805f
C11562 VPWR.t1043 VGND 0.06817f
C11563 VPWR.t796 VGND 0.02464f
C11564 VPWR.t1044 VGND 0.02189f
C11565 VPWR.n591 VGND 0.06768f
C11566 VPWR.n592 VGND 0.01329f
C11567 VPWR.n594 VGND 0.08003f
C11568 VPWR.t685 VGND 0.08842f
C11569 VPWR.t351 VGND 0.05805f
C11570 VPWR.t405 VGND 0.06817f
C11571 VPWR.t686 VGND 0.02464f
C11572 VPWR.t406 VGND 0.02189f
C11573 VPWR.n595 VGND 0.06768f
C11574 VPWR.n596 VGND 0.01329f
C11575 VPWR.n598 VGND 0.08003f
C11576 VPWR.t399 VGND 0.08842f
C11577 VPWR.t422 VGND 0.05805f
C11578 VPWR.t1762 VGND 0.06817f
C11579 VPWR.t400 VGND 0.02464f
C11580 VPWR.t1763 VGND 0.02189f
C11581 VPWR.n599 VGND 0.06768f
C11582 VPWR.n600 VGND 0.01329f
C11583 VPWR.n602 VGND 0.08003f
C11584 VPWR.t1756 VGND 0.08842f
C11585 VPWR.t421 VGND 0.05805f
C11586 VPWR.t1746 VGND 0.06817f
C11587 VPWR.t1757 VGND 0.02464f
C11588 VPWR.t1747 VGND 0.02189f
C11589 VPWR.n603 VGND 0.06768f
C11590 VPWR.n604 VGND 0.01329f
C11591 VPWR.n606 VGND 0.08003f
C11592 VPWR.t1740 VGND 0.08842f
C11593 VPWR.t350 VGND 0.05805f
C11594 VPWR.t286 VGND 0.06817f
C11595 VPWR.t1741 VGND 0.02464f
C11596 VPWR.t287 VGND 0.02189f
C11597 VPWR.n607 VGND 0.06768f
C11598 VPWR.n608 VGND 0.01329f
C11599 VPWR.n610 VGND 0.08003f
C11600 VPWR.t73 VGND 0.08842f
C11601 VPWR.t349 VGND 0.05805f
C11602 VPWR.t1904 VGND 0.06817f
C11603 VPWR.t74 VGND 0.02464f
C11604 VPWR.t1905 VGND 0.02189f
C11605 VPWR.n611 VGND 0.06768f
C11606 VPWR.n612 VGND 0.01329f
C11607 VPWR.n614 VGND 0.08003f
C11608 VPWR.t1898 VGND 0.08842f
C11609 VPWR.t423 VGND 0.05805f
C11610 VPWR.t383 VGND 0.06817f
C11611 VPWR.t1899 VGND 0.02464f
C11612 VPWR.t384 VGND 0.02189f
C11613 VPWR.n615 VGND 0.06768f
C11614 VPWR.n616 VGND 0.01329f
C11615 VPWR.n618 VGND 0.08003f
C11616 VPWR.t361 VGND 0.08842f
C11617 VPWR.t354 VGND 0.05805f
C11618 VPWR.t216 VGND 0.06817f
C11619 VPWR.t362 VGND 0.02464f
C11620 VPWR.t217 VGND 0.02189f
C11621 VPWR.n619 VGND 0.06768f
C11622 VPWR.n620 VGND 0.01329f
C11623 VPWR.n622 VGND 0.08003f
C11624 VPWR.t529 VGND 0.08842f
C11625 VPWR.t353 VGND 0.05805f
C11626 VPWR.t1155 VGND 0.06817f
C11627 VPWR.t530 VGND 0.02464f
C11628 VPWR.t1156 VGND 0.02189f
C11629 VPWR.n623 VGND 0.06768f
C11630 VPWR.n624 VGND 0.01329f
C11631 VPWR.n626 VGND 0.08003f
C11632 VPWR.t1796 VGND 0.08842f
C11633 VPWR.t420 VGND 0.05805f
C11634 VPWR.t537 VGND 0.06817f
C11635 VPWR.t1797 VGND 0.02464f
C11636 VPWR.t538 VGND 0.02189f
C11637 VPWR.n627 VGND 0.06768f
C11638 VPWR.n628 VGND 0.01329f
C11639 VPWR.n630 VGND 0.08003f
C11640 VPWR.t1248 VGND 0.08842f
C11641 VPWR.t419 VGND 0.05805f
C11642 VPWR.t1792 VGND 0.06817f
C11643 VPWR.t1249 VGND 0.02464f
C11644 VPWR.t1793 VGND 0.02189f
C11645 VPWR.n631 VGND 0.06768f
C11646 VPWR.n632 VGND 0.01329f
C11647 VPWR.n634 VGND 0.08003f
C11648 VPWR.t33 VGND 0.08842f
C11649 VPWR.t418 VGND 0.05805f
C11650 VPWR.t205 VGND 0.06817f
C11651 VPWR.t34 VGND 0.02464f
C11652 VPWR.t206 VGND 0.02189f
C11653 VPWR.n635 VGND 0.06768f
C11654 VPWR.n636 VGND 0.01329f
C11655 VPWR.n638 VGND 0.08003f
C11656 VPWR.t1004 VGND 0.08842f
C11657 VPWR.t348 VGND 0.05805f
C11658 VPWR.t1663 VGND 0.0986f
C11659 VPWR.n639 VGND 0.05634f
C11660 VPWR.n640 VGND 0.01329f
C11661 VPWR.n641 VGND 0.10289f
C11662 VPWR.n642 VGND 0.75117f
C11663 VPWR.n643 VGND 0.10289f
C11664 VPWR.t166 VGND 0.02464f
C11665 VPWR.t1390 VGND 0.02189f
C11666 VPWR.n644 VGND 0.06768f
C11667 VPWR.t1006 VGND 0.06817f
C11668 VPWR.t23 VGND 0.02464f
C11669 VPWR.t1007 VGND 0.02189f
C11670 VPWR.n645 VGND 0.06768f
C11671 VPWR.n646 VGND 0.10289f
C11672 VPWR.n647 VGND 0.10289f
C11673 VPWR.t1290 VGND 0.02464f
C11674 VPWR.t11 VGND 0.02189f
C11675 VPWR.n648 VGND 0.06768f
C11676 VPWR.t1252 VGND 0.06817f
C11677 VPWR.t920 VGND 0.02464f
C11678 VPWR.t1253 VGND 0.02189f
C11679 VPWR.n649 VGND 0.06768f
C11680 VPWR.n650 VGND 0.10289f
C11681 VPWR.n651 VGND 0.10289f
C11682 VPWR.t1838 VGND 0.02464f
C11683 VPWR.t1807 VGND 0.02189f
C11684 VPWR.n652 VGND 0.06768f
C11685 VPWR.t1843 VGND 0.06817f
C11686 VPWR.t337 VGND 0.02464f
C11687 VPWR.t1844 VGND 0.02189f
C11688 VPWR.n653 VGND 0.06768f
C11689 VPWR.n654 VGND 0.10289f
C11690 VPWR.n655 VGND 0.10289f
C11691 VPWR.t1219 VGND 0.02464f
C11692 VPWR.t343 VGND 0.02189f
C11693 VPWR.n656 VGND 0.06768f
C11694 VPWR.t1224 VGND 0.06817f
C11695 VPWR.t596 VGND 0.02464f
C11696 VPWR.t1225 VGND 0.02189f
C11697 VPWR.n657 VGND 0.06768f
C11698 VPWR.n658 VGND 0.10289f
C11699 VPWR.n659 VGND 0.10289f
C11700 VPWR.t1862 VGND 0.02464f
C11701 VPWR.t572 VGND 0.02189f
C11702 VPWR.n660 VGND 0.06768f
C11703 VPWR.t1867 VGND 0.06817f
C11704 VPWR.t58 VGND 0.02464f
C11705 VPWR.t1868 VGND 0.02189f
C11706 VPWR.n661 VGND 0.06768f
C11707 VPWR.n662 VGND 0.10289f
C11708 VPWR.n663 VGND 0.10289f
C11709 VPWR.t140 VGND 0.02464f
C11710 VPWR.t64 VGND 0.02189f
C11711 VPWR.n664 VGND 0.06768f
C11712 VPWR.t718 VGND 0.06817f
C11713 VPWR.t380 VGND 0.02464f
C11714 VPWR.t719 VGND 0.02189f
C11715 VPWR.n665 VGND 0.06768f
C11716 VPWR.n666 VGND 0.10289f
C11717 VPWR.n667 VGND 0.10289f
C11718 VPWR.t818 VGND 0.02464f
C11719 VPWR.t688 VGND 0.02189f
C11720 VPWR.n668 VGND 0.06768f
C11721 VPWR.t791 VGND 0.06817f
C11722 VPWR.t510 VGND 0.02464f
C11723 VPWR.t792 VGND 0.02189f
C11724 VPWR.n669 VGND 0.06768f
C11725 VPWR.n670 VGND 0.10289f
C11726 VPWR.n671 VGND 0.10289f
C11727 VPWR.t480 VGND 0.02464f
C11728 VPWR.t142 VGND 0.02189f
C11729 VPWR.n672 VGND 0.06768f
C11730 VPWR.t1069 VGND 0.10732f
C11731 VPWR.t568 VGND 0.05805f
C11732 VPWR.t1295 VGND 0.06817f
C11733 VPWR.t1070 VGND 0.02464f
C11734 VPWR.t1296 VGND 0.02189f
C11735 VPWR.n673 VGND 0.06768f
C11736 VPWR.t1077 VGND 0.02464f
C11737 VPWR.t962 VGND 0.02189f
C11738 VPWR.n674 VGND 0.06768f
C11739 VPWR.t1076 VGND 0.10732f
C11740 VPWR.t1169 VGND 0.05805f
C11741 VPWR.t961 VGND 0.06817f
C11742 VPWR.t180 VGND 0.02464f
C11743 VPWR.t1497 VGND 0.02189f
C11744 VPWR.n675 VGND 0.06768f
C11745 VPWR.n676 VGND 0.01329f
C11746 VPWR.n677 VGND 0.05634f
C11747 VPWR.t1496 VGND 0.0986f
C11748 VPWR.t177 VGND 0.05805f
C11749 VPWR.t179 VGND 0.08842f
C11750 VPWR.t882 VGND 0.02464f
C11751 VPWR.t870 VGND 0.02189f
C11752 VPWR.n678 VGND 0.06768f
C11753 VPWR.n679 VGND 0.01329f
C11754 VPWR.n681 VGND 0.08003f
C11755 VPWR.t869 VGND 0.06817f
C11756 VPWR.t1314 VGND 0.05805f
C11757 VPWR.t881 VGND 0.08842f
C11758 VPWR.t544 VGND 0.02464f
C11759 VPWR.t888 VGND 0.02189f
C11760 VPWR.n682 VGND 0.06768f
C11761 VPWR.n683 VGND 0.01329f
C11762 VPWR.n685 VGND 0.08003f
C11763 VPWR.t887 VGND 0.06817f
C11764 VPWR.t1315 VGND 0.05805f
C11765 VPWR.t543 VGND 0.08842f
C11766 VPWR.t1779 VGND 0.02464f
C11767 VPWR.t1237 VGND 0.02189f
C11768 VPWR.n686 VGND 0.06768f
C11769 VPWR.n687 VGND 0.01329f
C11770 VPWR.n689 VGND 0.08003f
C11771 VPWR.t1236 VGND 0.06817f
C11772 VPWR.t689 VGND 0.05805f
C11773 VPWR.t1778 VGND 0.08842f
C11774 VPWR.t1913 VGND 0.02464f
C11775 VPWR.t91 VGND 0.02189f
C11776 VPWR.n690 VGND 0.06768f
C11777 VPWR.n691 VGND 0.01329f
C11778 VPWR.n693 VGND 0.08003f
C11779 VPWR.t90 VGND 0.06817f
C11780 VPWR.t547 VGND 0.05805f
C11781 VPWR.t1912 VGND 0.08842f
C11782 VPWR.t430 VGND 0.02464f
C11783 VPWR.t1917 VGND 0.02189f
C11784 VPWR.n694 VGND 0.06768f
C11785 VPWR.n695 VGND 0.01329f
C11786 VPWR.n697 VGND 0.08003f
C11787 VPWR.t1916 VGND 0.06817f
C11788 VPWR.t548 VGND 0.05805f
C11789 VPWR.t429 VGND 0.08842f
C11790 VPWR.t578 VGND 0.02464f
C11791 VPWR.t436 VGND 0.02189f
C11792 VPWR.n698 VGND 0.06768f
C11793 VPWR.n699 VGND 0.01329f
C11794 VPWR.n701 VGND 0.08003f
C11795 VPWR.t435 VGND 0.06817f
C11796 VPWR.t692 VGND 0.05805f
C11797 VPWR.t577 VGND 0.08842f
C11798 VPWR.t735 VGND 0.02464f
C11799 VPWR.t582 VGND 0.02189f
C11800 VPWR.n702 VGND 0.06768f
C11801 VPWR.n703 VGND 0.01329f
C11802 VPWR.n705 VGND 0.08003f
C11803 VPWR.t581 VGND 0.06817f
C11804 VPWR.t178 VGND 0.05805f
C11805 VPWR.t734 VGND 0.08842f
C11806 VPWR.t1255 VGND 0.02464f
C11807 VPWR.t602 VGND 0.02189f
C11808 VPWR.n706 VGND 0.06768f
C11809 VPWR.n707 VGND 0.01329f
C11810 VPWR.n709 VGND 0.08003f
C11811 VPWR.t601 VGND 0.06817f
C11812 VPWR.t1167 VGND 0.05805f
C11813 VPWR.t1254 VGND 0.08842f
C11814 VPWR.t1175 VGND 0.02464f
C11815 VPWR.t1259 VGND 0.02189f
C11816 VPWR.n710 VGND 0.06768f
C11817 VPWR.n711 VGND 0.01329f
C11818 VPWR.n713 VGND 0.08003f
C11819 VPWR.t1258 VGND 0.06817f
C11820 VPWR.t690 VGND 0.05805f
C11821 VPWR.t1174 VGND 0.08842f
C11822 VPWR.t1191 VGND 0.02464f
C11823 VPWR.t1179 VGND 0.02189f
C11824 VPWR.n714 VGND 0.06768f
C11825 VPWR.n715 VGND 0.01329f
C11826 VPWR.n717 VGND 0.08003f
C11827 VPWR.t1178 VGND 0.06817f
C11828 VPWR.t691 VGND 0.05805f
C11829 VPWR.t1190 VGND 0.08842f
C11830 VPWR.t152 VGND 0.02464f
C11831 VPWR.t1124 VGND 0.02189f
C11832 VPWR.n718 VGND 0.06768f
C11833 VPWR.n719 VGND 0.01329f
C11834 VPWR.n721 VGND 0.08003f
C11835 VPWR.t1123 VGND 0.06817f
C11836 VPWR.t1168 VGND 0.05805f
C11837 VPWR.t151 VGND 0.08842f
C11838 VPWR.t830 VGND 0.02464f
C11839 VPWR.t1333 VGND 0.02189f
C11840 VPWR.n722 VGND 0.06768f
C11841 VPWR.n723 VGND 0.01329f
C11842 VPWR.n725 VGND 0.08003f
C11843 VPWR.t1332 VGND 0.06817f
C11844 VPWR.t549 VGND 0.05805f
C11845 VPWR.t829 VGND 0.08842f
C11846 VPWR.t768 VGND 0.02464f
C11847 VPWR.t810 VGND 0.02189f
C11848 VPWR.n726 VGND 0.06768f
C11849 VPWR.n727 VGND 0.01329f
C11850 VPWR.n729 VGND 0.08003f
C11851 VPWR.t809 VGND 0.06817f
C11852 VPWR.t1313 VGND 0.05805f
C11853 VPWR.t767 VGND 0.08842f
C11854 VPWR.t621 VGND 0.02464f
C11855 VPWR.t1132 VGND 0.02189f
C11856 VPWR.n730 VGND 0.06768f
C11857 VPWR.n731 VGND 0.01329f
C11858 VPWR.n733 VGND 0.08003f
C11859 VPWR.t1131 VGND 0.06817f
C11860 VPWR.t176 VGND 0.05805f
C11861 VPWR.t620 VGND 0.08842f
C11862 VPWR.n734 VGND 0.08003f
C11863 VPWR.n736 VGND 0.01329f
C11864 VPWR.n737 VGND 0.10289f
C11865 VPWR.n738 VGND 0.74646f
C11866 VPWR.n739 VGND 0.10289f
C11867 VPWR.t1073 VGND 0.02464f
C11868 VPWR.t1729 VGND 0.02189f
C11869 VPWR.n740 VGND 0.06768f
C11870 VPWR.t1072 VGND 0.10732f
C11871 VPWR.t30 VGND 0.05805f
C11872 VPWR.t1728 VGND 0.06817f
C11873 VPWR.t1135 VGND 0.08842f
C11874 VPWR.t1725 VGND 0.02464f
C11875 VPWR.t508 VGND 0.02189f
C11876 VPWR.n741 VGND 0.06768f
C11877 VPWR.n742 VGND 0.10289f
C11878 VPWR.n743 VGND 0.10289f
C11879 VPWR.t1136 VGND 0.02464f
C11880 VPWR.t800 VGND 0.02189f
C11881 VPWR.n744 VGND 0.06768f
C11882 VPWR.t1300 VGND 0.05805f
C11883 VPWR.t799 VGND 0.06817f
C11884 VPWR.t369 VGND 0.08842f
C11885 VPWR.t824 VGND 0.02464f
C11886 VPWR.t1339 VGND 0.02189f
C11887 VPWR.n745 VGND 0.06768f
C11888 VPWR.n746 VGND 0.10289f
C11889 VPWR.n747 VGND 0.10289f
C11890 VPWR.t370 VGND 0.02464f
C11891 VPWR.t138 VGND 0.02189f
C11892 VPWR.n748 VGND 0.06768f
C11893 VPWR.t29 VGND 0.05805f
C11894 VPWR.t137 VGND 0.06817f
C11895 VPWR.t1163 VGND 0.08842f
C11896 VPWR.t1128 VGND 0.02464f
C11897 VPWR.t1166 VGND 0.02189f
C11898 VPWR.n749 VGND 0.06768f
C11899 VPWR.n750 VGND 0.10289f
C11900 VPWR.n751 VGND 0.10289f
C11901 VPWR.t1164 VGND 0.02464f
C11902 VPWR.t1860 VGND 0.02189f
C11903 VPWR.n752 VGND 0.06768f
C11904 VPWR.t1262 VGND 0.05805f
C11905 VPWR.t1859 VGND 0.06817f
C11906 VPWR.t0 VGND 0.08842f
C11907 VPWR.t1858 VGND 0.02464f
C11908 VPWR.t68 VGND 0.02189f
C11909 VPWR.n753 VGND 0.06768f
C11910 VPWR.n754 VGND 0.10289f
C11911 VPWR.n755 VGND 0.10289f
C11912 VPWR.t1 VGND 0.02464f
C11913 VPWR.t858 VGND 0.02189f
C11914 VPWR.n756 VGND 0.06768f
C11915 VPWR.t27 VGND 0.05805f
C11916 VPWR.t857 VGND 0.06817f
C11917 VPWR.t437 VGND 0.08842f
C11918 VPWR.t856 VGND 0.02464f
C11919 VPWR.t335 VGND 0.02189f
C11920 VPWR.n757 VGND 0.06768f
C11921 VPWR.n758 VGND 0.10289f
C11922 VPWR.n759 VGND 0.10289f
C11923 VPWR.t438 VGND 0.02464f
C11924 VPWR.t1116 VGND 0.02189f
C11925 VPWR.n760 VGND 0.06768f
C11926 VPWR.t1298 VGND 0.05805f
C11927 VPWR.t1115 VGND 0.06817f
C11928 VPWR.t92 VGND 0.08842f
C11929 VPWR.t1114 VGND 0.02464f
C11930 VPWR.t1079 VGND 0.02189f
C11931 VPWR.n761 VGND 0.06768f
C11932 VPWR.n762 VGND 0.10289f
C11933 VPWR.n763 VGND 0.10289f
C11934 VPWR.t93 VGND 0.02464f
C11935 VPWR.t1243 VGND 0.02189f
C11936 VPWR.n764 VGND 0.06768f
C11937 VPWR.t1303 VGND 0.05805f
C11938 VPWR.t1242 VGND 0.06817f
C11939 VPWR.t889 VGND 0.08842f
C11940 VPWR.t1280 VGND 0.02464f
C11941 VPWR.t21 VGND 0.02189f
C11942 VPWR.n765 VGND 0.06768f
C11943 VPWR.n766 VGND 0.10289f
C11944 VPWR.n767 VGND 0.10289f
C11945 VPWR.t890 VGND 0.02464f
C11946 VPWR.t876 VGND 0.02189f
C11947 VPWR.n768 VGND 0.06768f
C11948 VPWR.t1301 VGND 0.05805f
C11949 VPWR.t875 VGND 0.06817f
C11950 VPWR.t184 VGND 0.02464f
C11951 VPWR.t1457 VGND 0.02189f
C11952 VPWR.n769 VGND 0.06768f
C11953 VPWR.t200 VGND 0.02464f
C11954 VPWR.t1562 VGND 0.02189f
C11955 VPWR.n770 VGND 0.06768f
C11956 VPWR.t1051 VGND 0.10732f
C11957 VPWR.t1310 VGND 0.05805f
C11958 VPWR.t616 VGND 0.06817f
C11959 VPWR.t1052 VGND 0.02464f
C11960 VPWR.t617 VGND 0.02189f
C11961 VPWR.n771 VGND 0.06768f
C11962 VPWR.n772 VGND 0.01329f
C11963 VPWR.n774 VGND 0.08003f
C11964 VPWR.t1908 VGND 0.08842f
C11965 VPWR.t1305 VGND 0.05805f
C11966 VPWR.t263 VGND 0.06817f
C11967 VPWR.t1909 VGND 0.02464f
C11968 VPWR.t264 VGND 0.02189f
C11969 VPWR.n775 VGND 0.06768f
C11970 VPWR.n776 VGND 0.01329f
C11971 VPWR.n778 VGND 0.08003f
C11972 VPWR.t257 VGND 0.08842f
C11973 VPWR.t170 VGND 0.05805f
C11974 VPWR.t807 VGND 0.06817f
C11975 VPWR.t258 VGND 0.02464f
C11976 VPWR.t808 VGND 0.02189f
C11977 VPWR.n779 VGND 0.06768f
C11978 VPWR.n780 VGND 0.01329f
C11979 VPWR.n782 VGND 0.08003f
C11980 VPWR.t783 VGND 0.08842f
C11981 VPWR.t169 VGND 0.05805f
C11982 VPWR.t373 VGND 0.06817f
C11983 VPWR.t784 VGND 0.02464f
C11984 VPWR.t374 VGND 0.02189f
C11985 VPWR.n783 VGND 0.06768f
C11986 VPWR.n784 VGND 0.01329f
C11987 VPWR.n786 VGND 0.08003f
C11988 VPWR.t1037 VGND 0.08842f
C11989 VPWR.t1309 VGND 0.05805f
C11990 VPWR.t1324 VGND 0.06817f
C11991 VPWR.t1038 VGND 0.02464f
C11992 VPWR.t1325 VGND 0.02189f
C11993 VPWR.n787 VGND 0.06768f
C11994 VPWR.n788 VGND 0.01329f
C11995 VPWR.n790 VGND 0.08003f
C11996 VPWR.t1318 VGND 0.08842f
C11997 VPWR.t175 VGND 0.05805f
C11998 VPWR.t561 VGND 0.06817f
C11999 VPWR.t1319 VGND 0.02464f
C12000 VPWR.t562 VGND 0.02189f
C12001 VPWR.n791 VGND 0.06768f
C12002 VPWR.n792 VGND 0.01329f
C12003 VPWR.n794 VGND 0.08003f
C12004 VPWR.t555 VGND 0.08842f
C12005 VPWR.t174 VGND 0.05805f
C12006 VPWR.t495 VGND 0.06817f
C12007 VPWR.t556 VGND 0.02464f
C12008 VPWR.t496 VGND 0.02189f
C12009 VPWR.n795 VGND 0.06768f
C12010 VPWR.n796 VGND 0.01329f
C12011 VPWR.n798 VGND 0.08003f
C12012 VPWR.t489 VGND 0.08842f
C12013 VPWR.t1308 VGND 0.05805f
C12014 VPWR.t4 VGND 0.06817f
C12015 VPWR.t490 VGND 0.02464f
C12016 VPWR.t5 VGND 0.02189f
C12017 VPWR.n799 VGND 0.06768f
C12018 VPWR.n800 VGND 0.01329f
C12019 VPWR.n802 VGND 0.08003f
C12020 VPWR.t845 VGND 0.08842f
C12021 VPWR.t1307 VGND 0.05805f
C12022 VPWR.t104 VGND 0.06817f
C12023 VPWR.t846 VGND 0.02464f
C12024 VPWR.t105 VGND 0.02189f
C12025 VPWR.n803 VGND 0.06768f
C12026 VPWR.n804 VGND 0.01329f
C12027 VPWR.n806 VGND 0.08003f
C12028 VPWR.t517 VGND 0.08842f
C12029 VPWR.t1304 VGND 0.05805f
C12030 VPWR.t425 VGND 0.06817f
C12031 VPWR.t518 VGND 0.02464f
C12032 VPWR.t426 VGND 0.02189f
C12033 VPWR.n807 VGND 0.06768f
C12034 VPWR.n808 VGND 0.01329f
C12035 VPWR.n810 VGND 0.08003f
C12036 VPWR.t585 VGND 0.08842f
C12037 VPWR.t168 VGND 0.05805f
C12038 VPWR.t710 VGND 0.06817f
C12039 VPWR.t586 VGND 0.02464f
C12040 VPWR.t711 VGND 0.02189f
C12041 VPWR.n811 VGND 0.06768f
C12042 VPWR.n812 VGND 0.01329f
C12043 VPWR.n814 VGND 0.08003f
C12044 VPWR.t704 VGND 0.08842f
C12045 VPWR.t167 VGND 0.05805f
C12046 VPWR.t1147 VGND 0.06817f
C12047 VPWR.t705 VGND 0.02464f
C12048 VPWR.t1148 VGND 0.02189f
C12049 VPWR.n815 VGND 0.06768f
C12050 VPWR.n816 VGND 0.01329f
C12051 VPWR.n818 VGND 0.08003f
C12052 VPWR.t1153 VGND 0.08842f
C12053 VPWR.t173 VGND 0.05805f
C12054 VPWR.t1283 VGND 0.06817f
C12055 VPWR.t1154 VGND 0.02464f
C12056 VPWR.t1284 VGND 0.02189f
C12057 VPWR.n819 VGND 0.06768f
C12058 VPWR.n820 VGND 0.01329f
C12059 VPWR.n822 VGND 0.08003f
C12060 VPWR.t967 VGND 0.08842f
C12061 VPWR.t172 VGND 0.05805f
C12062 VPWR.t39 VGND 0.06817f
C12063 VPWR.t968 VGND 0.02464f
C12064 VPWR.t40 VGND 0.02189f
C12065 VPWR.n823 VGND 0.06768f
C12066 VPWR.n824 VGND 0.01329f
C12067 VPWR.n826 VGND 0.08003f
C12068 VPWR.t1890 VGND 0.08842f
C12069 VPWR.t171 VGND 0.05805f
C12070 VPWR.t187 VGND 0.06817f
C12071 VPWR.t1891 VGND 0.02464f
C12072 VPWR.t188 VGND 0.02189f
C12073 VPWR.n827 VGND 0.06768f
C12074 VPWR.n828 VGND 0.01329f
C12075 VPWR.n830 VGND 0.08003f
C12076 VPWR.t199 VGND 0.08842f
C12077 VPWR.t1306 VGND 0.05805f
C12078 VPWR.t1561 VGND 0.0986f
C12079 VPWR.n831 VGND 0.05634f
C12080 VPWR.n832 VGND 0.01329f
C12081 VPWR.n833 VGND 0.10289f
C12082 VPWR.n834 VGND 0.75117f
C12083 VPWR.n835 VGND 0.10289f
C12084 VPWR.t868 VGND 0.02464f
C12085 VPWR.t1385 VGND 0.02189f
C12086 VPWR.n836 VGND 0.06768f
C12087 VPWR.t1010 VGND 0.06817f
C12088 VPWR.t25 VGND 0.02464f
C12089 VPWR.t1011 VGND 0.02189f
C12090 VPWR.n837 VGND 0.06768f
C12091 VPWR.n838 VGND 0.10289f
C12092 VPWR.n839 VGND 0.10289f
C12093 VPWR.t1292 VGND 0.02464f
C12094 VPWR.t13 VGND 0.02189f
C12095 VPWR.n840 VGND 0.06768f
C12096 VPWR.t942 VGND 0.06817f
C12097 VPWR.t922 VGND 0.02464f
C12098 VPWR.t943 VGND 0.02189f
C12099 VPWR.n841 VGND 0.06768f
C12100 VPWR.n842 VGND 0.10289f
C12101 VPWR.n843 VGND 0.10289f
C12102 VPWR.t1840 VGND 0.02464f
C12103 VPWR.t1809 VGND 0.02189f
C12104 VPWR.n844 VGND 0.06768f
C12105 VPWR.t1824 VGND 0.06817f
C12106 VPWR.t339 VGND 0.02464f
C12107 VPWR.t1825 VGND 0.02189f
C12108 VPWR.n845 VGND 0.06768f
C12109 VPWR.n846 VGND 0.10289f
C12110 VPWR.n847 VGND 0.10289f
C12111 VPWR.t1221 VGND 0.02464f
C12112 VPWR.t345 VGND 0.02189f
C12113 VPWR.n848 VGND 0.06768f
C12114 VPWR.t1226 VGND 0.06817f
C12115 VPWR.t598 VGND 0.02464f
C12116 VPWR.t1227 VGND 0.02189f
C12117 VPWR.n849 VGND 0.06768f
C12118 VPWR.n850 VGND 0.10289f
C12119 VPWR.n851 VGND 0.10289f
C12120 VPWR.t1864 VGND 0.02464f
C12121 VPWR.t574 VGND 0.02189f
C12122 VPWR.n852 VGND 0.06768f
C12123 VPWR.t1869 VGND 0.06817f
C12124 VPWR.t60 VGND 0.02464f
C12125 VPWR.t1870 VGND 0.02189f
C12126 VPWR.n853 VGND 0.06768f
C12127 VPWR.n854 VGND 0.10289f
C12128 VPWR.n855 VGND 0.10289f
C12129 VPWR.t1203 VGND 0.02464f
C12130 VPWR.t1813 VGND 0.02189f
C12131 VPWR.n856 VGND 0.06768f
C12132 VPWR.t720 VGND 0.06817f
C12133 VPWR.t1331 VGND 0.02464f
C12134 VPWR.t721 VGND 0.02189f
C12135 VPWR.n857 VGND 0.06768f
C12136 VPWR.n858 VGND 0.10289f
C12137 VPWR.n859 VGND 0.10289f
C12138 VPWR.t816 VGND 0.02464f
C12139 VPWR.t635 VGND 0.02189f
C12140 VPWR.n860 VGND 0.06768f
C12141 VPWR.t789 VGND 0.06817f
C12142 VPWR.t512 VGND 0.02464f
C12143 VPWR.t790 VGND 0.02189f
C12144 VPWR.n861 VGND 0.06768f
C12145 VPWR.n862 VGND 0.10289f
C12146 VPWR.n863 VGND 0.10289f
C12147 VPWR.t482 VGND 0.02464f
C12148 VPWR.t144 VGND 0.02189f
C12149 VPWR.n864 VGND 0.06768f
C12150 VPWR.t1067 VGND 0.10732f
C12151 VPWR.t667 VGND 0.05805f
C12152 VPWR.t1016 VGND 0.06817f
C12153 VPWR.t1068 VGND 0.02464f
C12154 VPWR.t1017 VGND 0.02189f
C12155 VPWR.n865 VGND 0.06768f
C12156 VPWR.t1054 VGND 0.02464f
C12157 VPWR.t615 VGND 0.02189f
C12158 VPWR.n866 VGND 0.06768f
C12159 VPWR.t1053 VGND 0.10732f
C12160 VPWR.t997 VGND 0.05805f
C12161 VPWR.t614 VGND 0.06817f
C12162 VPWR.t198 VGND 0.02464f
C12163 VPWR.t1569 VGND 0.02189f
C12164 VPWR.n867 VGND 0.06768f
C12165 VPWR.n868 VGND 0.01329f
C12166 VPWR.n869 VGND 0.05634f
C12167 VPWR.t1568 VGND 0.0986f
C12168 VPWR.t1886 VGND 0.05805f
C12169 VPWR.t197 VGND 0.08842f
C12170 VPWR.t1889 VGND 0.02464f
C12171 VPWR.t186 VGND 0.02189f
C12172 VPWR.n870 VGND 0.06768f
C12173 VPWR.n871 VGND 0.01329f
C12174 VPWR.n873 VGND 0.08003f
C12175 VPWR.t185 VGND 0.06817f
C12176 VPWR.t608 VGND 0.05805f
C12177 VPWR.t1888 VGND 0.08842f
C12178 VPWR.t964 VGND 0.02464f
C12179 VPWR.t38 VGND 0.02189f
C12180 VPWR.n874 VGND 0.06768f
C12181 VPWR.n875 VGND 0.01329f
C12182 VPWR.n877 VGND 0.08003f
C12183 VPWR.t37 VGND 0.06817f
C12184 VPWR.t609 VGND 0.05805f
C12185 VPWR.t963 VGND 0.08842f
C12186 VPWR.t1152 VGND 0.02464f
C12187 VPWR.t1282 VGND 0.02189f
C12188 VPWR.n878 VGND 0.06768f
C12189 VPWR.n879 VGND 0.01329f
C12190 VPWR.n881 VGND 0.08003f
C12191 VPWR.t1281 VGND 0.06817f
C12192 VPWR.t610 VGND 0.05805f
C12193 VPWR.t1151 VGND 0.08842f
C12194 VPWR.t703 VGND 0.02464f
C12195 VPWR.t1146 VGND 0.02189f
C12196 VPWR.n882 VGND 0.06768f
C12197 VPWR.n883 VGND 0.01329f
C12198 VPWR.n885 VGND 0.08003f
C12199 VPWR.t1145 VGND 0.06817f
C12200 VPWR.t1856 VGND 0.05805f
C12201 VPWR.t702 VGND 0.08842f
C12202 VPWR.t584 VGND 0.02464f
C12203 VPWR.t709 VGND 0.02189f
C12204 VPWR.n886 VGND 0.06768f
C12205 VPWR.n887 VGND 0.01329f
C12206 VPWR.n889 VGND 0.08003f
C12207 VPWR.t708 VGND 0.06817f
C12208 VPWR.t605 VGND 0.05805f
C12209 VPWR.t583 VGND 0.08842f
C12210 VPWR.t516 VGND 0.02464f
C12211 VPWR.t592 VGND 0.02189f
C12212 VPWR.n890 VGND 0.06768f
C12213 VPWR.n891 VGND 0.01329f
C12214 VPWR.n893 VGND 0.08003f
C12215 VPWR.t591 VGND 0.06817f
C12216 VPWR.t1884 VGND 0.05805f
C12217 VPWR.t515 VGND 0.08842f
C12218 VPWR.t842 VGND 0.02464f
C12219 VPWR.t103 VGND 0.02189f
C12220 VPWR.n894 VGND 0.06768f
C12221 VPWR.n895 VGND 0.01329f
C12222 VPWR.n897 VGND 0.08003f
C12223 VPWR.t102 VGND 0.06817f
C12224 VPWR.t1887 VGND 0.05805f
C12225 VPWR.t841 VGND 0.08842f
C12226 VPWR.t488 VGND 0.02464f
C12227 VPWR.t3 VGND 0.02189f
C12228 VPWR.n898 VGND 0.06768f
C12229 VPWR.n899 VGND 0.01329f
C12230 VPWR.n901 VGND 0.08003f
C12231 VPWR.t2 VGND 0.06817f
C12232 VPWR.t995 VGND 0.05805f
C12233 VPWR.t487 VGND 0.08842f
C12234 VPWR.t554 VGND 0.02464f
C12235 VPWR.t494 VGND 0.02189f
C12236 VPWR.n902 VGND 0.06768f
C12237 VPWR.n903 VGND 0.01329f
C12238 VPWR.n905 VGND 0.08003f
C12239 VPWR.t493 VGND 0.06817f
C12240 VPWR.t611 VGND 0.05805f
C12241 VPWR.t553 VGND 0.08842f
C12242 VPWR.t1317 VGND 0.02464f
C12243 VPWR.t560 VGND 0.02189f
C12244 VPWR.n906 VGND 0.06768f
C12245 VPWR.n907 VGND 0.01329f
C12246 VPWR.n909 VGND 0.08003f
C12247 VPWR.t559 VGND 0.06817f
C12248 VPWR.t1883 VGND 0.05805f
C12249 VPWR.t1316 VGND 0.08842f
C12250 VPWR.t1036 VGND 0.02464f
C12251 VPWR.t1323 VGND 0.02189f
C12252 VPWR.n910 VGND 0.06768f
C12253 VPWR.n911 VGND 0.01329f
C12254 VPWR.n913 VGND 0.08003f
C12255 VPWR.t1322 VGND 0.06817f
C12256 VPWR.t996 VGND 0.05805f
C12257 VPWR.t1035 VGND 0.08842f
C12258 VPWR.t786 VGND 0.02464f
C12259 VPWR.t372 VGND 0.02189f
C12260 VPWR.n914 VGND 0.06768f
C12261 VPWR.n915 VGND 0.01329f
C12262 VPWR.n917 VGND 0.08003f
C12263 VPWR.t371 VGND 0.06817f
C12264 VPWR.t606 VGND 0.05805f
C12265 VPWR.t785 VGND 0.08842f
C12266 VPWR.t256 VGND 0.02464f
C12267 VPWR.t822 VGND 0.02189f
C12268 VPWR.n918 VGND 0.06768f
C12269 VPWR.n919 VGND 0.01329f
C12270 VPWR.n921 VGND 0.08003f
C12271 VPWR.t821 VGND 0.06817f
C12272 VPWR.t607 VGND 0.05805f
C12273 VPWR.t255 VGND 0.08842f
C12274 VPWR.t1907 VGND 0.02464f
C12275 VPWR.t262 VGND 0.02189f
C12276 VPWR.n922 VGND 0.06768f
C12277 VPWR.n923 VGND 0.01329f
C12278 VPWR.n925 VGND 0.08003f
C12279 VPWR.t261 VGND 0.06817f
C12280 VPWR.t1885 VGND 0.05805f
C12281 VPWR.t1906 VGND 0.08842f
C12282 VPWR.n926 VGND 0.08003f
C12283 VPWR.n928 VGND 0.01329f
C12284 VPWR.n929 VGND 0.10289f
C12285 VPWR.n930 VGND 0.74646f
C12286 VPWR.n931 VGND 0.10289f
C12287 VPWR.t1060 VGND 0.02464f
C12288 VPWR.t906 VGND 0.02189f
C12289 VPWR.n932 VGND 0.06768f
C12290 VPWR.t1059 VGND 0.10732f
C12291 VPWR.t626 VGND 0.05805f
C12292 VPWR.t905 VGND 0.06817f
C12293 VPWR.t1208 VGND 0.08842f
C12294 VPWR.t910 VGND 0.02464f
C12295 VPWR.t1217 VGND 0.02189f
C12296 VPWR.n933 VGND 0.06768f
C12297 VPWR.n934 VGND 0.10289f
C12298 VPWR.n935 VGND 0.10289f
C12299 VPWR.t1209 VGND 0.02464f
C12300 VPWR.t774 VGND 0.02189f
C12301 VPWR.n936 VGND 0.06768f
C12302 VPWR.t1772 VGND 0.05805f
C12303 VPWR.t773 VGND 0.06817f
C12304 VPWR.t683 VGND 0.08842f
C12305 VPWR.t798 VGND 0.02464f
C12306 VPWR.t1040 VGND 0.02189f
C12307 VPWR.n937 VGND 0.06768f
C12308 VPWR.n938 VGND 0.10289f
C12309 VPWR.n939 VGND 0.10289f
C12310 VPWR.t684 VGND 0.02464f
C12311 VPWR.t404 VGND 0.02189f
C12312 VPWR.n940 VGND 0.06768f
C12313 VPWR.t625 VGND 0.05805f
C12314 VPWR.t403 VGND 0.06817f
C12315 VPWR.t1752 VGND 0.08842f
C12316 VPWR.t659 VGND 0.02464f
C12317 VPWR.t1761 VGND 0.02189f
C12318 VPWR.n941 VGND 0.06768f
C12319 VPWR.n942 VGND 0.10289f
C12320 VPWR.n943 VGND 0.10289f
C12321 VPWR.t1753 VGND 0.02464f
C12322 VPWR.t1745 VGND 0.02189f
C12323 VPWR.n944 VGND 0.06768f
C12324 VPWR.t977 VGND 0.05805f
C12325 VPWR.t1744 VGND 0.06817f
C12326 VPWR.t71 VGND 0.08842f
C12327 VPWR.t1737 VGND 0.02464f
C12328 VPWR.t852 VGND 0.02189f
C12329 VPWR.n945 VGND 0.06768f
C12330 VPWR.n946 VGND 0.10289f
C12331 VPWR.n947 VGND 0.10289f
C12332 VPWR.t72 VGND 0.02464f
C12333 VPWR.t1903 VGND 0.02189f
C12334 VPWR.n948 VGND 0.06768f
C12335 VPWR.t623 VGND 0.05805f
C12336 VPWR.t1902 VGND 0.06817f
C12337 VPWR.t359 VGND 0.08842f
C12338 VPWR.t1895 VGND 0.02464f
C12339 VPWR.t382 VGND 0.02189f
C12340 VPWR.n949 VGND 0.06768f
C12341 VPWR.n950 VGND 0.10289f
C12342 VPWR.n951 VGND 0.10289f
C12343 VPWR.t360 VGND 0.02464f
C12344 VPWR.t534 VGND 0.02189f
C12345 VPWR.n952 VGND 0.06768f
C12346 VPWR.t1770 VGND 0.05805f
C12347 VPWR.t533 VGND 0.06817f
C12348 VPWR.t1794 VGND 0.08842f
C12349 VPWR.t526 VGND 0.02464f
C12350 VPWR.t1805 VGND 0.02189f
C12351 VPWR.n953 VGND 0.06768f
C12352 VPWR.n954 VGND 0.10289f
C12353 VPWR.n955 VGND 0.10289f
C12354 VPWR.t1795 VGND 0.02464f
C12355 VPWR.t974 VGND 0.02189f
C12356 VPWR.n956 VGND 0.06768f
C12357 VPWR.t976 VGND 0.05805f
C12358 VPWR.t973 VGND 0.06817f
C12359 VPWR.t31 VGND 0.08842f
C12360 VPWR.t1247 VGND 0.02464f
C12361 VPWR.t1791 VGND 0.02189f
C12362 VPWR.n957 VGND 0.06768f
C12363 VPWR.n958 VGND 0.10289f
C12364 VPWR.n959 VGND 0.10289f
C12365 VPWR.t32 VGND 0.02464f
C12366 VPWR.t202 VGND 0.02189f
C12367 VPWR.n960 VGND 0.06768f
C12368 VPWR.t998 VGND 0.05805f
C12369 VPWR.t201 VGND 0.06817f
C12370 VPWR.t1003 VGND 0.02464f
C12371 VPWR.t1677 VGND 0.02189f
C12372 VPWR.n961 VGND 0.06768f
C12373 VPWR.t210 VGND 0.02464f
C12374 VPWR.t1529 VGND 0.02189f
C12375 VPWR.n962 VGND 0.06768f
C12376 VPWR.t1047 VGND 0.10732f
C12377 VPWR.t1836 VGND 0.05805f
C12378 VPWR.t959 VGND 0.06817f
C12379 VPWR.t1048 VGND 0.02464f
C12380 VPWR.t960 VGND 0.02189f
C12381 VPWR.n963 VGND 0.06768f
C12382 VPWR.n964 VGND 0.01329f
C12383 VPWR.n966 VGND 0.08003f
C12384 VPWR.t612 VGND 0.08842f
C12385 VPWR.t701 VGND 0.05805f
C12386 VPWR.t765 VGND 0.06817f
C12387 VPWR.t613 VGND 0.02464f
C12388 VPWR.t766 VGND 0.02189f
C12389 VPWR.n967 VGND 0.06768f
C12390 VPWR.n968 VGND 0.01329f
C12391 VPWR.n970 VGND 0.08003f
C12392 VPWR.t265 VGND 0.08842f
C12393 VPWR.t304 VGND 0.05805f
C12394 VPWR.t811 VGND 0.06817f
C12395 VPWR.t266 VGND 0.02464f
C12396 VPWR.t812 VGND 0.02189f
C12397 VPWR.n971 VGND 0.06768f
C12398 VPWR.n972 VGND 0.01329f
C12399 VPWR.n974 VGND 0.08003f
C12400 VPWR.t775 VGND 0.08842f
C12401 VPWR.t89 VGND 0.05805f
C12402 VPWR.t377 VGND 0.06817f
C12403 VPWR.t776 VGND 0.02464f
C12404 VPWR.t378 VGND 0.02189f
C12405 VPWR.n975 VGND 0.06768f
C12406 VPWR.n976 VGND 0.01329f
C12407 VPWR.n978 VGND 0.08003f
C12408 VPWR.t147 VGND 0.08842f
C12409 VPWR.t1112 VGND 0.05805f
C12410 VPWR.t1188 VGND 0.06817f
C12411 VPWR.t148 VGND 0.02464f
C12412 VPWR.t1189 VGND 0.02189f
C12413 VPWR.n979 VGND 0.06768f
C12414 VPWR.n980 VGND 0.01329f
C12415 VPWR.n982 VGND 0.08003f
C12416 VPWR.t1184 VGND 0.08842f
C12417 VPWR.t699 VGND 0.05805f
C12418 VPWR.t1172 VGND 0.06817f
C12419 VPWR.t1185 VGND 0.02464f
C12420 VPWR.t1173 VGND 0.02189f
C12421 VPWR.n983 VGND 0.06768f
C12422 VPWR.n984 VGND 0.01329f
C12423 VPWR.n986 VGND 0.08003f
C12424 VPWR.t563 VGND 0.08842f
C12425 VPWR.t308 VGND 0.05805f
C12426 VPWR.t441 VGND 0.06817f
C12427 VPWR.t564 VGND 0.02464f
C12428 VPWR.t442 VGND 0.02189f
C12429 VPWR.n987 VGND 0.06768f
C12430 VPWR.n988 VGND 0.01329f
C12431 VPWR.n990 VGND 0.08003f
C12432 VPWR.t497 VGND 0.08842f
C12433 VPWR.t1111 VGND 0.05805f
C12434 VPWR.t593 VGND 0.06817f
C12435 VPWR.t498 VGND 0.02464f
C12436 VPWR.t594 VGND 0.02189f
C12437 VPWR.n991 VGND 0.06768f
C12438 VPWR.n992 VGND 0.01329f
C12439 VPWR.n994 VGND 0.08003f
C12440 VPWR.t284 VGND 0.08842f
C12441 VPWR.t1110 VGND 0.05805f
C12442 VPWR.t110 VGND 0.06817f
C12443 VPWR.t285 VGND 0.02464f
C12444 VPWR.t111 VGND 0.02189f
C12445 VPWR.n995 VGND 0.06768f
C12446 VPWR.n996 VGND 0.01329f
C12447 VPWR.n998 VGND 0.08003f
C12448 VPWR.t106 VGND 0.08842f
C12449 VPWR.t700 VGND 0.05805f
C12450 VPWR.t433 VGND 0.06817f
C12451 VPWR.t107 VGND 0.02464f
C12452 VPWR.t434 VGND 0.02189f
C12453 VPWR.n999 VGND 0.06768f
C12454 VPWR.n1000 VGND 0.01329f
C12455 VPWR.n1002 VGND 0.08003f
C12456 VPWR.t589 VGND 0.08842f
C12457 VPWR.t88 VGND 0.05805f
C12458 VPWR.t716 VGND 0.06817f
C12459 VPWR.t590 VGND 0.02464f
C12460 VPWR.t717 VGND 0.02189f
C12461 VPWR.n1003 VGND 0.06768f
C12462 VPWR.n1004 VGND 0.01329f
C12463 VPWR.n1006 VGND 0.08003f
C12464 VPWR.t712 VGND 0.08842f
C12465 VPWR.t87 VGND 0.05805f
C12466 VPWR.t1782 VGND 0.06817f
C12467 VPWR.t713 VGND 0.02464f
C12468 VPWR.t1783 VGND 0.02189f
C12469 VPWR.n1007 VGND 0.06768f
C12470 VPWR.n1008 VGND 0.01329f
C12471 VPWR.n1010 VGND 0.08003f
C12472 VPWR.t1143 VGND 0.08842f
C12473 VPWR.t307 VGND 0.05805f
C12474 VPWR.t1287 VGND 0.06817f
C12475 VPWR.t1144 VGND 0.02464f
C12476 VPWR.t1288 VGND 0.02189f
C12477 VPWR.n1011 VGND 0.06768f
C12478 VPWR.n1012 VGND 0.01329f
C12479 VPWR.n1014 VGND 0.08003f
C12480 VPWR.t535 VGND 0.08842f
C12481 VPWR.t306 VGND 0.05805f
C12482 VPWR.t885 VGND 0.06817f
C12483 VPWR.t536 VGND 0.02464f
C12484 VPWR.t886 VGND 0.02189f
C12485 VPWR.n1015 VGND 0.06768f
C12486 VPWR.n1016 VGND 0.01329f
C12487 VPWR.n1018 VGND 0.08003f
C12488 VPWR.t35 VGND 0.08842f
C12489 VPWR.t305 VGND 0.05805f
C12490 VPWR.t163 VGND 0.06817f
C12491 VPWR.t36 VGND 0.02464f
C12492 VPWR.t164 VGND 0.02189f
C12493 VPWR.n1019 VGND 0.06768f
C12494 VPWR.n1020 VGND 0.01329f
C12495 VPWR.n1022 VGND 0.08003f
C12496 VPWR.t209 VGND 0.08842f
C12497 VPWR.t1109 VGND 0.05805f
C12498 VPWR.t1528 VGND 0.0986f
C12499 VPWR.n1023 VGND 0.05634f
C12500 VPWR.n1024 VGND 0.01329f
C12501 VPWR.n1025 VGND 0.10289f
C12502 VPWR.n1026 VGND 4.32396f
C12503 VPWR.n1027 VGND 0.04856f
C12504 VPWR.n1028 VGND -0.0138f
C12505 VPWR.n1029 VGND 0.0225f
C12506 VPWR.t1532 VGND 0.01981f
C12507 VPWR.n1031 VGND 0.04233f
C12508 VPWR.t1640 VGND 0.02189f
C12509 VPWR.n1032 VGND 0.0347f
C12510 VPWR.t211 VGND 0.06817f
C12511 VPWR.n1033 VGND 0.0225f
C12512 VPWR.t1424 VGND 0.01981f
C12513 VPWR.n1035 VGND 0.04233f
C12514 VPWR.t212 VGND 0.02189f
C12515 VPWR.n1036 VGND 0.0347f
C12516 VPWR.n1037 VGND -0.0138f
C12517 VPWR.n1038 VGND 0.04856f
C12518 VPWR.n1039 VGND 0.02048f
C12519 VPWR.n1040 VGND 0.01403f
C12520 VPWR.n1041 VGND 0.04617f
C12521 VPWR.n1042 VGND 0.07207f
C12522 VPWR.n1043 VGND 0.04023f
C12523 VPWR.n1044 VGND 0.04856f
C12524 VPWR.n1045 VGND -0.0138f
C12525 VPWR.n1046 VGND 0.0225f
C12526 VPWR.t1510 VGND 0.01981f
C12527 VPWR.n1048 VGND 0.04233f
C12528 VPWR.t1160 VGND 0.02189f
C12529 VPWR.n1049 VGND 0.0347f
C12530 VPWR.t1159 VGND 0.06817f
C12531 VPWR.t1373 VGND 0.08842f
C12532 VPWR.n1050 VGND 0.0225f
C12533 VPWR.t1551 VGND 0.01981f
C12534 VPWR.n1052 VGND 0.04233f
C12535 VPWR.t542 VGND 0.02189f
C12536 VPWR.n1053 VGND 0.0347f
C12537 VPWR.n1055 VGND 0.14325f
C12538 VPWR.n1056 VGND 0.06176f
C12539 VPWR.n1057 VGND 0.02542f
C12540 VPWR.t1604 VGND 0.02464f
C12541 VPWR.t1596 VGND 0.02189f
C12542 VPWR.n1058 VGND 0.06768f
C12543 VPWR.t1595 VGND 0.06817f
C12544 VPWR.t1351 VGND 0.08842f
C12545 VPWR.t1632 VGND 0.02464f
C12546 VPWR.t1624 VGND 0.02189f
C12547 VPWR.n1059 VGND 0.06768f
C12548 VPWR.t1352 VGND 0.02464f
C12549 VPWR.t1475 VGND 0.02189f
C12550 VPWR.n1061 VGND 0.06768f
C12551 VPWR.t1347 VGND 0.05805f
C12552 VPWR.t1474 VGND 0.0986f
C12553 VPWR.n1062 VGND 0.05631f
C12554 VPWR.n1063 VGND 0.01256f
C12555 VPWR.n1064 VGND 0.02213f
C12556 VPWR.n1065 VGND 0.02429f
C12557 VPWR.n1067 VGND 0.01347f
C12558 VPWR.n1068 VGND 0.13004f
C12559 VPWR.n1069 VGND 0.02213f
C12560 VPWR.n1070 VGND 0.02429f
C12561 VPWR.n1071 VGND 0.01268f
C12562 VPWR.n1074 VGND 0.01268f
C12563 VPWR.n1076 VGND 0.02047f
C12564 VPWR.n1077 VGND 0.02084f
C12565 VPWR.n1078 VGND 0.01347f
C12566 VPWR.n1079 VGND 0.13004f
C12567 VPWR.n1080 VGND 0.02213f
C12568 VPWR.n1081 VGND 0.02429f
C12569 VPWR.n1082 VGND 0.01268f
C12570 VPWR.n1084 VGND 0.01268f
C12571 VPWR.n1086 VGND 0.02047f
C12572 VPWR.n1087 VGND 0.02084f
C12573 VPWR.n1088 VGND 0.01347f
C12574 VPWR.n1089 VGND 0.13004f
C12575 VPWR.n1090 VGND 0.02213f
C12576 VPWR.n1091 VGND 0.02429f
C12577 VPWR.n1092 VGND 0.01268f
C12578 VPWR.n1094 VGND 0.01268f
C12579 VPWR.n1096 VGND 0.02047f
C12580 VPWR.n1097 VGND 0.02084f
C12581 VPWR.n1098 VGND 0.01347f
C12582 VPWR.n1099 VGND 0.13004f
C12583 VPWR.n1100 VGND 0.02213f
C12584 VPWR.n1101 VGND 0.02429f
C12585 VPWR.n1102 VGND 0.01268f
C12586 VPWR.n1104 VGND 0.01268f
C12587 VPWR.n1106 VGND 0.02047f
C12588 VPWR.n1107 VGND 0.02084f
C12589 VPWR.n1108 VGND 0.01347f
C12590 VPWR.n1109 VGND 0.01963f
C12591 VPWR.n1110 VGND 0.02213f
C12592 VPWR.n1111 VGND 0.02429f
C12593 VPWR.n1112 VGND 0.01347f
C12594 VPWR.n1114 VGND 0.02304f
C12595 VPWR.n1115 VGND 0.01456f
C12596 VPWR.n1116 VGND 0.02047f
C12597 VPWR.n1117 VGND 0.02084f
C12598 VPWR.n1118 VGND 0.01313f
C12599 VPWR.n1119 VGND 0.02213f
C12600 VPWR.n1120 VGND 0.02429f
C12601 VPWR.t1653 VGND 0.02464f
C12602 VPWR.t1371 VGND 0.02189f
C12603 VPWR.n1122 VGND 0.06768f
C12604 VPWR.t1652 VGND 0.10732f
C12605 VPWR.t1642 VGND 0.05805f
C12606 VPWR.t1370 VGND 0.06817f
C12607 VPWR.t1522 VGND 0.08842f
C12608 VPWR.t1421 VGND 0.02464f
C12609 VPWR.t1507 VGND 0.02189f
C12610 VPWR.n1123 VGND 0.06768f
C12611 VPWR.n1125 VGND 0.02304f
C12612 VPWR.n1126 VGND 0.02731f
C12613 VPWR.n1127 VGND 0.02542f
C12614 VPWR.n1128 VGND 0.10289f
C12615 VPWR.n1130 VGND 0.01329f
C12616 VPWR.n1131 VGND 0.04856f
C12617 VPWR.n1132 VGND 0.04023f
C12618 VPWR.n1133 VGND 0.02048f
C12619 VPWR.n1134 VGND 0.01403f
C12620 VPWR.n1135 VGND 0.04617f
C12621 VPWR.n1136 VGND 0.07207f
C12622 VPWR.n1137 VGND 0.04856f
C12623 VPWR.n1138 VGND 0.04856f
C12624 VPWR.n1139 VGND 0.04856f
C12625 VPWR.n1140 VGND 0.04856f
C12626 VPWR.n1141 VGND 0.04856f
C12627 VPWR.n1142 VGND 0.04856f
C12628 VPWR.n1143 VGND 0.04023f
C12629 VPWR.n1145 VGND -0.0138f
C12630 VPWR.n1146 VGND 0.0225f
C12631 VPWR.t1637 VGND 0.01981f
C12632 VPWR.n1148 VGND 0.04233f
C12633 VPWR.t388 VGND 0.02189f
C12634 VPWR.n1149 VGND 0.0347f
C12635 VPWR.t387 VGND 0.06817f
C12636 VPWR.t1382 VGND 0.05805f
C12637 VPWR.t1509 VGND 0.08842f
C12638 VPWR.n1150 VGND 0.0225f
C12639 VPWR.t1380 VGND 0.01981f
C12640 VPWR.n1152 VGND 0.04233f
C12641 VPWR.t221 VGND 0.02189f
C12642 VPWR.n1153 VGND 0.0347f
C12643 VPWR.n1156 VGND 0.0225f
C12644 VPWR.t1621 VGND 0.01981f
C12645 VPWR.n1158 VGND 0.04233f
C12646 VPWR.t1108 VGND 0.02189f
C12647 VPWR.n1159 VGND 0.0347f
C12648 VPWR.t732 VGND 0.06817f
C12649 VPWR.n1160 VGND 0.0225f
C12650 VPWR.t1480 VGND 0.01981f
C12651 VPWR.n1162 VGND 0.04233f
C12652 VPWR.t733 VGND 0.02189f
C12653 VPWR.n1163 VGND 0.0347f
C12654 VPWR.n1166 VGND 0.0225f
C12655 VPWR.t1358 VGND 0.01981f
C12656 VPWR.n1168 VGND 0.04233f
C12657 VPWR.t486 VGND 0.02189f
C12658 VPWR.n1169 VGND 0.0347f
C12659 VPWR.t697 VGND 0.06817f
C12660 VPWR.n1170 VGND 0.0225f
C12661 VPWR.t1607 VGND 0.01981f
C12662 VPWR.n1172 VGND 0.04233f
C12663 VPWR.t698 VGND 0.02189f
C12664 VPWR.n1173 VGND 0.0347f
C12665 VPWR.n1176 VGND 0.02304f
C12666 VPWR.n1177 VGND 0.02731f
C12667 VPWR.n1178 VGND 0.02542f
C12668 VPWR.t1406 VGND 0.02464f
C12669 VPWR.t1401 VGND 0.02189f
C12670 VPWR.n1179 VGND 0.06768f
C12671 VPWR.t1512 VGND 0.05805f
C12672 VPWR.t1519 VGND 0.06817f
C12673 VPWR.t1523 VGND 0.02464f
C12674 VPWR.t1520 VGND 0.02189f
C12675 VPWR.n1180 VGND 0.06768f
C12676 VPWR.n1182 VGND 0.08003f
C12677 VPWR.t1687 VGND 0.08842f
C12678 VPWR.t1553 VGND 0.05805f
C12679 VPWR.t1679 VGND 0.06817f
C12680 VPWR.t1688 VGND 0.02464f
C12681 VPWR.t1680 VGND 0.02189f
C12682 VPWR.n1183 VGND 0.06768f
C12683 VPWR.n1185 VGND 0.08003f
C12684 VPWR.t1405 VGND 0.08842f
C12685 VPWR.t1661 VGND 0.05805f
C12686 VPWR.t1400 VGND 0.06817f
C12687 VPWR.t1477 VGND 0.05805f
C12688 VPWR.t1603 VGND 0.08842f
C12689 VPWR.t1366 VGND 0.02464f
C12690 VPWR.t1467 VGND 0.02189f
C12691 VPWR.n1186 VGND 0.06768f
C12692 VPWR.n1188 VGND 0.08003f
C12693 VPWR.t1466 VGND 0.06817f
C12694 VPWR.t1451 VGND 0.05805f
C12695 VPWR.t1365 VGND 0.08842f
C12696 VPWR.t1345 VGND 0.02464f
C12697 VPWR.t1723 VGND 0.02189f
C12698 VPWR.n1189 VGND 0.06768f
C12699 VPWR.n1191 VGND 0.08003f
C12700 VPWR.t1722 VGND 0.06817f
C12701 VPWR.t1601 VGND 0.05805f
C12702 VPWR.t1344 VGND 0.08842f
C12703 VPWR.t1599 VGND 0.02464f
C12704 VPWR.t1704 VGND 0.02189f
C12705 VPWR.n1192 VGND 0.06768f
C12706 VPWR.n1194 VGND 0.02304f
C12707 VPWR.n1195 VGND 0.02731f
C12708 VPWR.n1196 VGND 0.02542f
C12709 VPWR.n1197 VGND 0.01268f
C12710 VPWR.n1199 VGND 0.08003f
C12711 VPWR.t1703 VGND 0.06817f
C12712 VPWR.t1579 VGND 0.05805f
C12713 VPWR.t1598 VGND 0.08842f
C12714 VPWR.t1472 VGND 0.02464f
C12715 VPWR.t1545 VGND 0.02189f
C12716 VPWR.n1200 VGND 0.06768f
C12717 VPWR.n1202 VGND 0.08003f
C12718 VPWR.t1544 VGND 0.06817f
C12719 VPWR.t1426 VGND 0.05805f
C12720 VPWR.t1471 VGND 0.08842f
C12721 VPWR.t1446 VGND 0.02464f
C12722 VPWR.t1441 VGND 0.02189f
C12723 VPWR.n1203 VGND 0.06768f
C12724 VPWR.n1205 VGND 0.08003f
C12725 VPWR.t1440 VGND 0.06817f
C12726 VPWR.t1709 VGND 0.05805f
C12727 VPWR.t1445 VGND 0.08842f
C12728 VPWR.t1685 VGND 0.02464f
C12729 VPWR.t1696 VGND 0.02189f
C12730 VPWR.n1206 VGND 0.06768f
C12731 VPWR.n1208 VGND 0.02304f
C12732 VPWR.n1209 VGND 0.02731f
C12733 VPWR.n1210 VGND 0.02542f
C12734 VPWR.n1211 VGND 0.01268f
C12735 VPWR.n1213 VGND 0.08003f
C12736 VPWR.t1695 VGND 0.06817f
C12737 VPWR.t1666 VGND 0.05805f
C12738 VPWR.t1684 VGND 0.08842f
C12739 VPWR.t1577 VGND 0.02464f
C12740 VPWR.t1656 VGND 0.02189f
C12741 VPWR.n1214 VGND 0.06768f
C12742 VPWR.n1216 VGND 0.08003f
C12743 VPWR.t1655 VGND 0.06817f
C12744 VPWR.t1443 VGND 0.05805f
C12745 VPWR.t1576 VGND 0.08842f
C12746 VPWR.t1418 VGND 0.02464f
C12747 VPWR.t1548 VGND 0.02189f
C12748 VPWR.n1217 VGND 0.06768f
C12749 VPWR.n1219 VGND 0.08003f
C12750 VPWR.t1547 VGND 0.06817f
C12751 VPWR.t1428 VGND 0.05805f
C12752 VPWR.t1417 VGND 0.08842f
C12753 VPWR.n1220 VGND 0.08003f
C12754 VPWR.n1222 VGND 0.01268f
C12755 VPWR.n1224 VGND 0.0225f
C12756 VPWR.t1585 VGND 0.01981f
C12757 VPWR.n1226 VGND 0.04233f
C12758 VPWR.t506 VGND 0.02189f
C12759 VPWR.n1227 VGND 0.0347f
C12760 VPWR.t1448 VGND 0.10732f
C12761 VPWR.t1433 VGND 0.05805f
C12762 VPWR.t895 VGND 0.06817f
C12763 VPWR.n1228 VGND 0.0225f
C12764 VPWR.t1449 VGND 0.01981f
C12765 VPWR.n1230 VGND 0.04233f
C12766 VPWR.t896 VGND 0.02189f
C12767 VPWR.n1231 VGND 0.0347f
C12768 VPWR.n1232 VGND -0.0138f
C12769 VPWR.n1233 VGND 0.03466f
C12770 VPWR.t398 VGND 0.72151f
C12771 VPWR.n1234 VGND 0.39351f
C12772 VPWR.t47 VGND 0.72151f
C12773 VPWR.n1235 VGND 0.30604f
C12774 VPWR.n1236 VGND 0.21505f
C12775 VPWR.t743 VGND 0.04227f
C12776 VPWR.t628 VGND 0.0106f
C12777 VPWR.t631 VGND 0.0106f
C12778 VPWR.n1238 VGND 0.02326f
C12779 VPWR.t1311 VGND 0.0106f
C12780 VPWR.t1768 VGND 0.0106f
C12781 VPWR.n1239 VGND 0.02322f
C12782 VPWR.t53 VGND 0.0106f
C12783 VPWR.t52 VGND 0.0106f
C12784 VPWR.n1240 VGND 0.02322f
C12785 VPWR.n1241 VGND 0.07706f
C12786 VPWR.n1242 VGND 0.13446f
C12787 VPWR.n1243 VGND 0.04257f
C12788 VPWR.n1244 VGND 0.03127f
C12789 VPWR.t48 VGND 0.0106f
C12790 VPWR.t54 VGND 0.0106f
C12791 VPWR.n1245 VGND 0.02326f
C12792 VPWR.n1246 VGND 0.09541f
C12793 VPWR.n1248 VGND 0.01206f
C12794 VPWR.n1249 VGND 0.01413f
C12795 VPWR.n1250 VGND 0.02072f
C12796 VPWR.t742 VGND 0.04227f
C12797 VPWR.n1251 VGND 0.11136f
C12798 VPWR.t1854 VGND 0.04226f
C12799 VPWR.t80 VGND 0.04226f
C12800 VPWR.n1253 VGND 0.09943f
C12801 VPWR.n1254 VGND 0.2482f
C12802 VPWR.n1255 VGND 1.21348f
C12803 VPWR.n1256 VGND 0.03466f
C12804 VPWR.t229 VGND 0.72151f
C12805 VPWR.n1257 VGND 0.39351f
C12806 VPWR.t157 VGND 0.72151f
C12807 VPWR.n1258 VGND 0.30604f
C12808 VPWR.n1259 VGND 0.21698f
C12809 VPWR.t415 VGND 0.0106f
C12810 VPWR.t413 VGND 0.0106f
C12811 VPWR.n1261 VGND 0.02326f
C12812 VPWR.t412 VGND 0.0106f
C12813 VPWR.t409 VGND 0.0106f
C12814 VPWR.n1262 VGND 0.02322f
C12815 VPWR.t1845 VGND 0.0106f
C12816 VPWR.t1846 VGND 0.0106f
C12817 VPWR.n1263 VGND 0.02322f
C12818 VPWR.n1264 VGND 0.07706f
C12819 VPWR.n1265 VGND 0.13446f
C12820 VPWR.n1266 VGND 0.04257f
C12821 VPWR.n1267 VGND 0.03127f
C12822 VPWR.t1030 VGND 0.0106f
C12823 VPWR.t158 VGND 0.0106f
C12824 VPWR.n1268 VGND 0.02326f
C12825 VPWR.n1269 VGND 0.09541f
C12826 VPWR.n1271 VGND 0.01206f
C12827 VPWR.n1272 VGND 0.01413f
C12828 VPWR.n1273 VGND 0.02034f
C12829 VPWR.t744 VGND 0.04221f
C12830 VPWR.n1275 VGND 0.04512f
C12831 VPWR.t550 VGND 0.0423f
C12832 VPWR.n1277 VGND 0.06737f
C12833 VPWR.n1278 VGND 0.2482f
C12834 VPWR.n1279 VGND 1.21348f
C12835 VPWR.n1280 VGND 0.03466f
C12836 VPWR.t234 VGND 0.72151f
C12837 VPWR.n1281 VGND 0.39351f
C12838 VPWR.t81 VGND 0.72151f
C12839 VPWR.n1282 VGND 0.30604f
C12840 VPWR.n1283 VGND 0.21698f
C12841 VPWR.t918 VGND 0.0106f
C12842 VPWR.t916 VGND 0.0106f
C12843 VPWR.n1285 VGND 0.02326f
C12844 VPWR.t915 VGND 0.0106f
C12845 VPWR.t914 VGND 0.0106f
C12846 VPWR.n1286 VGND 0.02322f
C12847 VPWR.t757 VGND 0.0106f
C12848 VPWR.t764 VGND 0.0106f
C12849 VPWR.n1287 VGND 0.02322f
C12850 VPWR.n1288 VGND 0.07706f
C12851 VPWR.n1289 VGND 0.13446f
C12852 VPWR.n1290 VGND 0.04257f
C12853 VPWR.n1291 VGND 0.03127f
C12854 VPWR.t761 VGND 0.0106f
C12855 VPWR.t758 VGND 0.0106f
C12856 VPWR.n1292 VGND 0.02326f
C12857 VPWR.n1293 VGND 0.09541f
C12858 VPWR.n1295 VGND 0.01206f
C12859 VPWR.n1296 VGND 0.01413f
C12860 VPWR.n1297 VGND 0.02034f
C12861 VPWR.n1298 VGND 0.01034f
C12862 VPWR.t1855 VGND 0.0423f
C12863 VPWR.t82 VGND 0.0423f
C12864 VPWR.n1300 VGND 0.12493f
C12865 VPWR.n1301 VGND 0.2482f
C12866 VPWR.n1302 VGND 1.21348f
C12867 VPWR.t1199 VGND 0.04223f
C12868 VPWR.t748 VGND 0.0423f
C12869 VPWR.t1201 VGND 0.04194f
C12870 VPWR.n1303 VGND 0.10875f
C12871 VPWR.t397 VGND 0.04146f
C12872 VPWR.n1304 VGND 0.0501f
C12873 VPWR.n1305 VGND 0.03466f
C12874 VPWR.t1120 VGND 0.03991f
C12875 VPWR.n1306 VGND 0.03796f
C12876 VPWR.t1193 VGND 0.0106f
C12877 VPWR.t231 VGND 0.0106f
C12878 VPWR.n1307 VGND 0.02315f
C12879 VPWR.t331 VGND 0.03708f
C12880 VPWR.n1308 VGND 0.05562f
C12881 VPWR.n1309 VGND 0.03466f
C12882 VPWR.t394 VGND 0.04225f
C12883 VPWR.n1310 VGND 0.05319f
C12884 VPWR.n1311 VGND 0.02034f
C12885 VPWR.n1312 VGND 0.03466f
C12886 VPWR.t233 VGND 0.0106f
C12887 VPWR.t444 VGND 0.0106f
C12888 VPWR.n1314 VGND 0.02315f
C12889 VPWR.n1315 VGND 0.03393f
C12890 VPWR.n1317 VGND 0.02599f
C12891 VPWR.n1318 VGND 0.02599f
C12892 VPWR.n1319 VGND 0.03466f
C12893 VPWR.t984 VGND 0.0106f
C12894 VPWR.t1197 VGND 0.0106f
C12895 VPWR.n1321 VGND 0.02315f
C12896 VPWR.n1322 VGND 0.02666f
C12897 VPWR.t934 VGND 0.0106f
C12898 VPWR.t1767 VGND 0.0106f
C12899 VPWR.n1323 VGND 0.02315f
C12900 VPWR.n1324 VGND 0.02946f
C12901 VPWR.n1326 VGND 0.03146f
C12902 VPWR.n1327 VGND 0.01187f
C12903 VPWR.t1232 VGND 0.03554f
C12904 VPWR.t1198 VGND 0.07996f
C12905 VPWR.t747 VGND 0.09329f
C12906 VPWR.t1200 VGND 0.17324f
C12907 VPWR.t393 VGND 0.09321f
C12908 VPWR.t443 VGND 0.10581f
C12909 VPWR.t232 VGND 0.10287f
C12910 VPWR.t230 VGND 0.16452f
C12911 VPWR.t1192 VGND 0.13993f
C12912 VPWR.t330 VGND 0.09329f
C12913 VPWR.t1196 VGND 0.09329f
C12914 VPWR.t1766 VGND 0.09329f
C12915 VPWR.t983 VGND 0.09329f
C12916 VPWR.t933 VGND 0.09329f
C12917 VPWR.t1119 VGND 0.09329f
C12918 VPWR.t396 VGND 0.09217f
C12919 VPWR.n1329 VGND 0.31703f
C12920 VPWR.n1330 VGND 0.12882f
C12921 VPWR.n1331 VGND 0.01413f
C12922 VPWR.n1332 VGND 0.02599f
C12923 VPWR.n1333 VGND 0.03127f
C12924 VPWR.n1335 VGND 0.04701f
C12925 VPWR.n1336 VGND 0.23407f
C12926 VPWR.n1337 VGND 1.21348f
C12927 VPWR.t160 VGND 0.04155f
C12928 VPWR.t745 VGND 0.04143f
C12929 VPWR.t746 VGND 0.04226f
C12930 VPWR.n1338 VGND 0.05889f
C12931 VPWR.t1312 VGND 0.04034f
C12932 VPWR.t55 VGND 0.04034f
C12933 VPWR.n1339 VGND 0.07319f
C12934 VPWR.n1340 VGND 0.03466f
C12935 VPWR.n1342 VGND 0.03466f
C12936 VPWR.t629 VGND 0.0106f
C12937 VPWR.t1327 VGND 0.0106f
C12938 VPWR.n1343 VGND 0.02315f
C12939 VPWR.t56 VGND 0.0106f
C12940 VPWR.t937 VGND 0.0106f
C12941 VPWR.n1344 VGND 0.02315f
C12942 VPWR.n1345 VGND 0.04717f
C12943 VPWR.t939 VGND 0.04225f
C12944 VPWR.t445 VGND 0.04225f
C12945 VPWR.n1346 VGND 0.09738f
C12946 VPWR.n1347 VGND 0.02034f
C12947 VPWR.n1348 VGND 0.03466f
C12948 VPWR.t1329 VGND 0.0106f
C12949 VPWR.t333 VGND 0.0106f
C12950 VPWR.n1350 VGND 0.02315f
C12951 VPWR.t954 VGND 0.0106f
C12952 VPWR.t1764 VGND 0.0106f
C12953 VPWR.n1351 VGND 0.02315f
C12954 VPWR.n1352 VGND 0.05331f
C12955 VPWR.n1354 VGND 0.03466f
C12956 VPWR.n1355 VGND 0.03466f
C12957 VPWR.n1356 VGND 0.03466f
C12958 VPWR.t1769 VGND 0.0106f
C12959 VPWR.t630 VGND 0.0106f
C12960 VPWR.n1358 VGND 0.02315f
C12961 VPWR.t51 VGND 0.0106f
C12962 VPWR.t50 VGND 0.0106f
C12963 VPWR.n1359 VGND 0.02315f
C12964 VPWR.n1360 VGND 0.04717f
C12965 VPWR.n1363 VGND 0.03466f
C12966 VPWR.n1364 VGND 0.02599f
C12967 VPWR.t159 VGND 0.72151f
C12968 VPWR.n1366 VGND 0.39351f
C12969 VPWR.t49 VGND 0.72151f
C12970 VPWR.n1367 VGND 0.30604f
C12971 VPWR.n1368 VGND 0.21505f
C12972 VPWR.n1369 VGND 0.01413f
C12973 VPWR.n1370 VGND 0.02599f
C12974 VPWR.n1371 VGND 0.03146f
C12975 VPWR.n1373 VGND 0.04309f
C12976 VPWR.n1374 VGND 0.05837f
C12977 VPWR.n1375 VGND 0.23388f
C12978 VPWR.n1376 VGND 1.21348f
C12979 VPWR.t501 VGND 0.04221f
C12980 VPWR.t269 VGND 0.04221f
C12981 VPWR.n1377 VGND 0.01034f
C12982 VPWR.t411 VGND 0.04034f
C12983 VPWR.t156 VGND 0.04034f
C12984 VPWR.n1378 VGND 0.07319f
C12985 VPWR.n1379 VGND 0.03466f
C12986 VPWR.n1381 VGND 0.03466f
C12987 VPWR.t416 VGND 0.0106f
C12988 VPWR.t952 VGND 0.0106f
C12989 VPWR.n1382 VGND 0.02315f
C12990 VPWR.t1028 VGND 0.0106f
C12991 VPWR.t446 VGND 0.0106f
C12992 VPWR.n1383 VGND 0.02315f
C12993 VPWR.n1384 VGND 0.04717f
C12994 VPWR.t447 VGND 0.04225f
C12995 VPWR.t936 VGND 0.04225f
C12996 VPWR.n1385 VGND 0.09738f
C12997 VPWR.n1386 VGND 0.02034f
C12998 VPWR.n1387 VGND 0.03466f
C12999 VPWR.t956 VGND 0.0106f
C13000 VPWR.t1765 VGND 0.0106f
C13001 VPWR.n1389 VGND 0.02315f
C13002 VPWR.t1326 VGND 0.0106f
C13003 VPWR.t449 VGND 0.0106f
C13004 VPWR.n1390 VGND 0.02315f
C13005 VPWR.n1391 VGND 0.05331f
C13006 VPWR.n1393 VGND 0.03466f
C13007 VPWR.n1394 VGND 0.03466f
C13008 VPWR.n1395 VGND 0.03466f
C13009 VPWR.t417 VGND 0.0106f
C13010 VPWR.t414 VGND 0.0106f
C13011 VPWR.n1397 VGND 0.02315f
C13012 VPWR.t1847 VGND 0.0106f
C13013 VPWR.t1029 VGND 0.0106f
C13014 VPWR.n1398 VGND 0.02315f
C13015 VPWR.n1399 VGND 0.04717f
C13016 VPWR.n1402 VGND 0.03466f
C13017 VPWR.n1403 VGND 0.02599f
C13018 VPWR.t410 VGND 0.72151f
C13019 VPWR.n1405 VGND 0.39351f
C13020 VPWR.t155 VGND 0.72151f
C13021 VPWR.n1406 VGND 0.30604f
C13022 VPWR.n1407 VGND 0.21698f
C13023 VPWR.n1408 VGND 0.01413f
C13024 VPWR.n1409 VGND 0.02599f
C13025 VPWR.n1410 VGND 0.03146f
C13026 VPWR.n1412 VGND 0.08532f
C13027 VPWR.n1413 VGND 0.23765f
C13028 VPWR.n1414 VGND 1.21348f
C13029 VPWR.t917 VGND 0.04034f
C13030 VPWR.t759 VGND 0.04034f
C13031 VPWR.n1415 VGND 0.07319f
C13032 VPWR.n1416 VGND 0.03466f
C13033 VPWR.n1418 VGND 0.03466f
C13034 VPWR.t912 VGND 0.0106f
C13035 VPWR.t1328 VGND 0.0106f
C13036 VPWR.n1419 VGND 0.02315f
C13037 VPWR.t760 VGND 0.0106f
C13038 VPWR.t392 VGND 0.0106f
C13039 VPWR.n1420 VGND 0.02315f
C13040 VPWR.n1421 VGND 0.04717f
C13041 VPWR.t953 VGND 0.04225f
C13042 VPWR.t950 VGND 0.04225f
C13043 VPWR.n1422 VGND 0.09738f
C13044 VPWR.n1423 VGND 0.02034f
C13045 VPWR.n1424 VGND 0.03466f
C13046 VPWR.t448 VGND 0.0106f
C13047 VPWR.t390 VGND 0.0106f
C13048 VPWR.n1426 VGND 0.02315f
C13049 VPWR.t395 VGND 0.0106f
C13050 VPWR.t935 VGND 0.0106f
C13051 VPWR.n1427 VGND 0.02315f
C13052 VPWR.n1428 VGND 0.05331f
C13053 VPWR.n1430 VGND 0.03466f
C13054 VPWR.n1431 VGND 0.03466f
C13055 VPWR.n1432 VGND 0.03466f
C13056 VPWR.t913 VGND 0.0106f
C13057 VPWR.t911 VGND 0.0106f
C13058 VPWR.n1434 VGND 0.02315f
C13059 VPWR.t763 VGND 0.0106f
C13060 VPWR.t762 VGND 0.0106f
C13061 VPWR.n1435 VGND 0.02315f
C13062 VPWR.n1436 VGND 0.04717f
C13063 VPWR.n1439 VGND 0.03466f
C13064 VPWR.n1440 VGND 0.02599f
C13065 VPWR.t389 VGND 0.55347f
C13066 VPWR.n1442 VGND 0.31666f
C13067 VPWR.t391 VGND 0.55347f
C13068 VPWR.n1443 VGND 0.24813f
C13069 VPWR.n1444 VGND 0.20802f
C13070 VPWR.n1445 VGND 0.31801f
C13071 VPWR.n1446 VGND 4.62393f
C13072 VPWR.n1447 VGND 6.76927f
C13073 VPWR.n1448 VGND 0.06176f
C13074 VPWR.n1449 VGND 0.81338f
C13075 VPWR.n1450 VGND 0.74646f
C13076 VPWR.n1451 VGND 0.04794f
C13077 VPWR.n1452 VGND 0.04023f
C13078 VPWR.n1453 VGND 0.02048f
C13079 VPWR.n1454 VGND 0.01403f
C13080 VPWR.n1455 VGND 0.04617f
C13081 VPWR.n1456 VGND 0.0574f
C13082 VPWR.n1457 VGND 0.06785f
C13083 VPWR.n1458 VGND 0.02048f
C13084 VPWR.n1459 VGND 0.01403f
C13085 VPWR.n1460 VGND 0.04617f
C13086 VPWR.n1461 VGND 0.07207f
C13087 VPWR.n1462 VGND 0.06785f
C13088 VPWR.n1463 VGND 0.04856f
C13089 VPWR.n1464 VGND 0.04023f
C13090 VPWR.n1465 VGND 0.10289f
C13091 VPWR.n1466 VGND 0.01329f
C13092 VPWR.n1468 VGND 0.08003f
C13093 VPWR.t1609 VGND 0.08842f
C13094 VPWR.t1564 VGND 0.05805f
C13095 VPWR.t1892 VGND 0.06817f
C13096 VPWR.n1469 VGND 0.0225f
C13097 VPWR.t1610 VGND 0.01981f
C13098 VPWR.n1471 VGND 0.04233f
C13099 VPWR.t1893 VGND 0.02189f
C13100 VPWR.n1472 VGND 0.0347f
C13101 VPWR.n1473 VGND 0.01329f
C13102 VPWR.n1475 VGND 0.08003f
C13103 VPWR.t1711 VGND 0.08842f
C13104 VPWR.t1693 VGND 0.05805f
C13105 VPWR.t825 VGND 0.06817f
C13106 VPWR.n1476 VGND 0.0225f
C13107 VPWR.t1712 VGND 0.01981f
C13108 VPWR.n1478 VGND 0.04233f
C13109 VPWR.t826 VGND 0.02189f
C13110 VPWR.n1479 VGND 0.0347f
C13111 VPWR.n1481 VGND 0.08003f
C13112 VPWR.t1482 VGND 0.08842f
C13113 VPWR.t1349 VGND 0.05805f
C13114 VPWR.t149 VGND 0.06817f
C13115 VPWR.n1482 VGND 0.0225f
C13116 VPWR.t1483 VGND 0.01981f
C13117 VPWR.n1484 VGND 0.04233f
C13118 VPWR.t150 VGND 0.02189f
C13119 VPWR.n1485 VGND 0.0347f
C13120 VPWR.n1487 VGND 0.06176f
C13121 VPWR.n1488 VGND -0.0138f
C13122 VPWR.n1489 VGND 0.10289f
C13123 VPWR.n1490 VGND 0.01329f
C13124 VPWR.n1492 VGND 0.08003f
C13125 VPWR.t1584 VGND 0.08842f
C13126 VPWR.t1459 VGND 0.05805f
C13127 VPWR.t505 VGND 0.06817f
C13128 VPWR.t1614 VGND 0.05805f
C13129 VPWR.t1606 VGND 0.08842f
C13130 VPWR.n1493 VGND 0.08003f
C13131 VPWR.n1495 VGND 0.01329f
C13132 VPWR.n1496 VGND 0.04023f
C13133 VPWR.n1497 VGND 0.10289f
C13134 VPWR.n1498 VGND -0.0138f
C13135 VPWR.n1499 VGND 0.06176f
C13136 VPWR.n1500 VGND 0.06176f
C13137 VPWR.n1501 VGND -0.0138f
C13138 VPWR.n1502 VGND 0.04023f
C13139 VPWR.n1503 VGND 0.10289f
C13140 VPWR.n1504 VGND 0.01329f
C13141 VPWR.n1506 VGND 0.08003f
C13142 VPWR.t1357 VGND 0.08842f
C13143 VPWR.t1616 VGND 0.05805f
C13144 VPWR.t485 VGND 0.06817f
C13145 VPWR.t1464 VGND 0.05805f
C13146 VPWR.t1479 VGND 0.08842f
C13147 VPWR.n1507 VGND 0.08003f
C13148 VPWR.n1509 VGND 0.01329f
C13149 VPWR.n1510 VGND 0.04023f
C13150 VPWR.n1511 VGND 0.10289f
C13151 VPWR.n1512 VGND -0.0138f
C13152 VPWR.n1513 VGND 0.06176f
C13153 VPWR.n1514 VGND 0.06176f
C13154 VPWR.n1515 VGND -0.0138f
C13155 VPWR.n1516 VGND 0.04023f
C13156 VPWR.n1517 VGND 0.10289f
C13157 VPWR.n1518 VGND 0.01329f
C13158 VPWR.n1520 VGND 0.08003f
C13159 VPWR.t1620 VGND 0.08842f
C13160 VPWR.t1494 VGND 0.05805f
C13161 VPWR.t1107 VGND 0.06817f
C13162 VPWR.t1612 VGND 0.05805f
C13163 VPWR.t1636 VGND 0.08842f
C13164 VPWR.n1521 VGND 0.08003f
C13165 VPWR.n1523 VGND 0.01329f
C13166 VPWR.n1524 VGND 0.04023f
C13167 VPWR.n1525 VGND 0.10289f
C13168 VPWR.n1526 VGND -0.0138f
C13169 VPWR.n1527 VGND 0.06176f
C13170 VPWR.n1528 VGND 0.06176f
C13171 VPWR.n1529 VGND 0.06176f
C13172 VPWR.n1530 VGND 0.06176f
C13173 VPWR.n1531 VGND -0.0138f
C13174 VPWR.n1532 VGND 0.10289f
C13175 VPWR.n1533 VGND 0.01329f
C13176 VPWR.n1535 VGND 0.08003f
C13177 VPWR.t220 VGND 0.06817f
C13178 VPWR.t1363 VGND 0.05805f
C13179 VPWR.t1379 VGND 0.08842f
C13180 VPWR.n1536 VGND 0.08003f
C13181 VPWR.n1538 VGND 0.01329f
C13182 VPWR.n1539 VGND 0.10289f
C13183 VPWR.n1540 VGND 0.04023f
C13184 VPWR.n1541 VGND 0.04856f
C13185 VPWR.n1542 VGND 0.06785f
C13186 VPWR.n1543 VGND 0.02048f
C13187 VPWR.n1544 VGND 0.01403f
C13188 VPWR.n1545 VGND 0.04617f
C13189 VPWR.n1546 VGND 0.07207f
C13190 VPWR.n1547 VGND 0.06785f
C13191 VPWR.n1548 VGND 0.02048f
C13192 VPWR.n1549 VGND 0.01403f
C13193 VPWR.n1550 VGND 0.04617f
C13194 VPWR.n1551 VGND 0.07207f
C13195 VPWR.n1552 VGND 0.06785f
C13196 VPWR.n1553 VGND 0.02048f
C13197 VPWR.n1554 VGND 0.01403f
C13198 VPWR.n1555 VGND 0.04617f
C13199 VPWR.n1556 VGND 0.07207f
C13200 VPWR.n1557 VGND 0.06785f
C13201 VPWR.n1558 VGND 0.02048f
C13202 VPWR.n1559 VGND 0.01403f
C13203 VPWR.n1560 VGND 0.04617f
C13204 VPWR.n1561 VGND 0.07207f
C13205 VPWR.n1562 VGND 0.06785f
C13206 VPWR.n1563 VGND 0.02048f
C13207 VPWR.n1564 VGND 0.01403f
C13208 VPWR.n1565 VGND 0.04617f
C13209 VPWR.n1566 VGND 0.07207f
C13210 VPWR.n1567 VGND 0.06785f
C13211 VPWR.n1568 VGND 0.02048f
C13212 VPWR.n1569 VGND 0.01403f
C13213 VPWR.n1570 VGND 0.04617f
C13214 VPWR.n1571 VGND 0.07207f
C13215 VPWR.n1572 VGND 0.06785f
C13216 VPWR.n1573 VGND 0.02048f
C13217 VPWR.n1574 VGND 0.01403f
C13218 VPWR.n1575 VGND 0.04617f
C13219 VPWR.n1576 VGND 0.07207f
C13220 VPWR.n1577 VGND 0.06785f
C13221 VPWR.n1578 VGND 0.02048f
C13222 VPWR.n1579 VGND 0.01403f
C13223 VPWR.n1580 VGND 0.04617f
C13224 VPWR.n1581 VGND 0.07207f
C13225 VPWR.n1582 VGND 0.06785f
C13226 VPWR.n1583 VGND 0.04856f
C13227 VPWR.n1584 VGND 0.04023f
C13228 VPWR.n1585 VGND 0.10289f
C13229 VPWR.n1586 VGND -0.0138f
C13230 VPWR.n1587 VGND 0.06176f
C13231 VPWR.n1588 VGND 0.06176f
C13232 VPWR.n1589 VGND -0.0138f
C13233 VPWR.n1591 VGND 0.01268f
C13234 VPWR.n1593 VGND 0.08003f
C13235 VPWR.t1506 VGND 0.06817f
C13236 VPWR.t1387 VGND 0.05805f
C13237 VPWR.t1420 VGND 0.08842f
C13238 VPWR.n1594 VGND 0.08003f
C13239 VPWR.n1596 VGND 0.01268f
C13240 VPWR.n1597 VGND 0.02542f
C13241 VPWR.n1598 VGND 0.02304f
C13242 VPWR.n1599 VGND 0.02731f
C13243 VPWR.n1601 VGND 0.02047f
C13244 VPWR.n1602 VGND 0.02084f
C13245 VPWR.n1603 VGND 0.01313f
C13246 VPWR.n1605 VGND 0.01347f
C13247 VPWR.n1606 VGND 0.01763f
C13248 VPWR.n1607 VGND 0.17544f
C13249 VPWR.n1608 VGND 0.13004f
C13250 VPWR.n1609 VGND 0.01763f
C13251 VPWR.n1610 VGND 0.01313f
C13252 VPWR.n1611 VGND 0.02213f
C13253 VPWR.n1612 VGND 0.02429f
C13254 VPWR.n1613 VGND 0.02542f
C13255 VPWR.n1614 VGND 0.02304f
C13256 VPWR.n1615 VGND 0.02731f
C13257 VPWR.n1617 VGND 0.02047f
C13258 VPWR.n1618 VGND 0.02084f
C13259 VPWR.n1619 VGND 0.01347f
C13260 VPWR.n1620 VGND 0.01763f
C13261 VPWR.n1621 VGND 0.01313f
C13262 VPWR.n1622 VGND 0.02213f
C13263 VPWR.n1623 VGND 0.02429f
C13264 VPWR.n1624 VGND 0.02542f
C13265 VPWR.n1625 VGND 0.02304f
C13266 VPWR.n1626 VGND 0.02731f
C13267 VPWR.n1628 VGND 0.02047f
C13268 VPWR.n1629 VGND 0.02084f
C13269 VPWR.n1630 VGND 0.01313f
C13270 VPWR.n1632 VGND 0.01347f
C13271 VPWR.n1633 VGND 0.01763f
C13272 VPWR.n1634 VGND 0.13004f
C13273 VPWR.n1635 VGND 0.13004f
C13274 VPWR.n1636 VGND 0.01763f
C13275 VPWR.n1637 VGND 0.01313f
C13276 VPWR.n1638 VGND 0.02213f
C13277 VPWR.n1639 VGND 0.02429f
C13278 VPWR.n1640 VGND 0.02542f
C13279 VPWR.n1641 VGND 0.02304f
C13280 VPWR.n1642 VGND 0.02731f
C13281 VPWR.n1644 VGND 0.02047f
C13282 VPWR.n1645 VGND 0.02084f
C13283 VPWR.n1646 VGND 0.01347f
C13284 VPWR.n1647 VGND 0.01763f
C13285 VPWR.n1648 VGND 0.01313f
C13286 VPWR.n1649 VGND 0.02213f
C13287 VPWR.n1650 VGND 0.02429f
C13288 VPWR.n1651 VGND 0.02542f
C13289 VPWR.n1652 VGND 0.02304f
C13290 VPWR.n1653 VGND 0.02731f
C13291 VPWR.n1655 VGND 0.02047f
C13292 VPWR.n1656 VGND 0.02084f
C13293 VPWR.n1657 VGND 0.01313f
C13294 VPWR.n1659 VGND 0.01347f
C13295 VPWR.n1660 VGND 0.01763f
C13296 VPWR.n1661 VGND 0.13004f
C13297 VPWR.n1662 VGND 0.13004f
C13298 VPWR.n1663 VGND 0.01763f
C13299 VPWR.n1664 VGND 0.01313f
C13300 VPWR.n1665 VGND 0.02213f
C13301 VPWR.n1666 VGND 0.02429f
C13302 VPWR.n1667 VGND 0.02542f
C13303 VPWR.n1668 VGND 0.02304f
C13304 VPWR.n1669 VGND 0.02731f
C13305 VPWR.n1671 VGND 0.02047f
C13306 VPWR.n1672 VGND 0.02084f
C13307 VPWR.n1673 VGND 0.01347f
C13308 VPWR.n1674 VGND 0.01763f
C13309 VPWR.n1675 VGND 0.01313f
C13310 VPWR.n1676 VGND 0.02213f
C13311 VPWR.n1677 VGND 0.02429f
C13312 VPWR.n1678 VGND 0.02542f
C13313 VPWR.n1679 VGND 0.02304f
C13314 VPWR.n1680 VGND 0.02731f
C13315 VPWR.n1682 VGND 0.02047f
C13316 VPWR.n1683 VGND 0.02084f
C13317 VPWR.n1684 VGND 0.01313f
C13318 VPWR.n1686 VGND 0.01347f
C13319 VPWR.n1687 VGND 0.01763f
C13320 VPWR.n1688 VGND 0.13004f
C13321 VPWR.n1689 VGND 0.13004f
C13322 VPWR.n1690 VGND 0.01763f
C13323 VPWR.n1691 VGND 0.01313f
C13324 VPWR.n1692 VGND 0.02213f
C13325 VPWR.n1693 VGND 0.02429f
C13326 VPWR.n1694 VGND 0.02542f
C13327 VPWR.n1695 VGND 0.02304f
C13328 VPWR.n1696 VGND 0.02731f
C13329 VPWR.n1698 VGND 0.02047f
C13330 VPWR.n1699 VGND 0.02084f
C13331 VPWR.n1700 VGND 0.01347f
C13332 VPWR.n1701 VGND 0.01763f
C13333 VPWR.n1702 VGND 0.01313f
C13334 VPWR.n1703 VGND 0.02213f
C13335 VPWR.n1704 VGND 0.02429f
C13336 VPWR.n1705 VGND 0.02542f
C13337 VPWR.n1706 VGND 0.02304f
C13338 VPWR.n1707 VGND 0.02731f
C13339 VPWR.n1709 VGND 0.02047f
C13340 VPWR.n1710 VGND 0.02084f
C13341 VPWR.n1711 VGND 0.01313f
C13342 VPWR.n1713 VGND 0.01347f
C13343 VPWR.n1714 VGND 0.01763f
C13344 VPWR.n1715 VGND 0.13004f
C13345 VPWR.n1716 VGND 0.02213f
C13346 VPWR.n1717 VGND 0.02429f
C13347 VPWR.n1718 VGND 0.02304f
C13348 VPWR.n1719 VGND 0.02731f
C13349 VPWR.n1721 VGND 0.02047f
C13350 VPWR.n1722 VGND 0.02084f
C13351 VPWR.n1723 VGND 0.01313f
C13352 VPWR.n1725 VGND 0.01347f
C13353 VPWR.n1726 VGND 0.01763f
C13354 VPWR.n1727 VGND 0.1565f
C13355 VPWR.n1728 VGND 0.01879f
C13356 VPWR.n1729 VGND 0.01313f
C13357 VPWR.n1730 VGND 0.02047f
C13358 VPWR.n1731 VGND 0.02084f
C13359 VPWR.n1733 VGND 0.02304f
C13360 VPWR.n1734 VGND 0.02731f
C13361 VPWR.n1735 VGND 0.02542f
C13362 VPWR.n1737 VGND 0.01268f
C13363 VPWR.n1739 VGND 0.08003f
C13364 VPWR.t1623 VGND 0.06817f
C13365 VPWR.t1502 VGND 0.05805f
C13366 VPWR.t1631 VGND 0.08842f
C13367 VPWR.n1740 VGND 0.08003f
C13368 VPWR.n1742 VGND 0.01268f
C13369 VPWR.n1744 VGND 0.04023f
C13370 VPWR.n1745 VGND 0.0225f
C13371 VPWR.t1374 VGND 0.01981f
C13372 VPWR.n1747 VGND 0.04233f
C13373 VPWR.t1027 VGND 0.02189f
C13374 VPWR.n1748 VGND 0.0347f
C13375 VPWR.t1644 VGND 0.05805f
C13376 VPWR.t1026 VGND 0.06817f
C13377 VPWR.t1682 VGND 0.05805f
C13378 VPWR.t1423 VGND 0.08842f
C13379 VPWR.n1749 VGND 0.08003f
C13380 VPWR.n1751 VGND 0.01329f
C13381 VPWR.n1752 VGND 0.10289f
C13382 VPWR.n1753 VGND -0.0138f
C13383 VPWR.n1754 VGND 0.06176f
C13384 VPWR.n1755 VGND 0.06176f
C13385 VPWR.n1756 VGND -0.0138f
C13386 VPWR.n1757 VGND 0.10289f
C13387 VPWR.n1758 VGND 0.01329f
C13388 VPWR.n1760 VGND 0.08003f
C13389 VPWR.t541 VGND 0.06817f
C13390 VPWR.t1626 VGND 0.05805f
C13391 VPWR.t1550 VGND 0.08842f
C13392 VPWR.n1761 VGND 0.08003f
C13393 VPWR.n1763 VGND 0.01329f
C13394 VPWR.n1764 VGND 0.10289f
C13395 VPWR.n1765 VGND 0.04023f
C13396 VPWR.n1766 VGND 0.04856f
C13397 VPWR.n1767 VGND 0.06785f
C13398 VPWR.n1768 VGND 0.02048f
C13399 VPWR.n1769 VGND 0.01403f
C13400 VPWR.n1770 VGND 0.04617f
C13401 VPWR.n1771 VGND 0.07207f
C13402 VPWR.n1772 VGND 0.06785f
C13403 VPWR.n1773 VGND 0.02048f
C13404 VPWR.n1774 VGND 0.01403f
C13405 VPWR.n1775 VGND 0.04617f
C13406 VPWR.n1776 VGND 0.07207f
C13407 VPWR.n1777 VGND 0.02048f
C13408 VPWR.n1778 VGND 0.01403f
C13409 VPWR.n1779 VGND 0.04616f
C13410 VPWR.n1780 VGND 0.038f
C13411 VPWR.n1781 VGND 0.02048f
C13412 VPWR.n1782 VGND 0.01403f
C13413 VPWR.n1783 VGND 0.04617f
C13414 VPWR.n1784 VGND 0.07207f
C13415 VPWR.n1785 VGND 0.06785f
C13416 VPWR.n1786 VGND 0.04856f
C13417 VPWR.n1787 VGND 0.04023f
C13418 VPWR.n1788 VGND 0.10289f
C13419 VPWR.n1789 VGND 0.01329f
C13420 VPWR.n1791 VGND 0.08003f
C13421 VPWR.t1531 VGND 0.08842f
C13422 VPWR.t1514 VGND 0.05805f
C13423 VPWR.t1639 VGND 0.0986f
C13424 VPWR.n1792 VGND 0.05634f
C13425 VPWR.n1793 VGND 0.01329f
C13426 VPWR.n1794 VGND 0.10289f
C13427 VPWR.n1795 VGND 0.12172f
C13428 VPWR.n1796 VGND 0.75117f
C13429 VPWR.n1797 VGND 0.06176f
C13430 VPWR.n1798 VGND 0.06176f
C13431 VPWR.n1799 VGND 0.06176f
C13432 VPWR.n1800 VGND 0.06176f
C13433 VPWR.n1801 VGND 0.06176f
C13434 VPWR.n1802 VGND 0.06176f
C13435 VPWR.n1803 VGND 0.06176f
C13436 VPWR.n1804 VGND 0.06176f
C13437 VPWR.n1805 VGND 0.06176f
C13438 VPWR.n1806 VGND 0.06176f
C13439 VPWR.n1807 VGND 0.06176f
C13440 VPWR.n1808 VGND 0.06176f
C13441 VPWR.n1809 VGND 0.06176f
C13442 VPWR.n1810 VGND 0.06176f
C13443 VPWR.n1811 VGND 0.06176f
C13444 VPWR.n1812 VGND 0.14325f
C13445 VPWR.n1813 VGND 0.75117f
C13446 VPWR.n1814 VGND 0.75117f
C13447 VPWR.n1815 VGND 0.14325f
C13448 VPWR.n1816 VGND 0.10289f
C13449 VPWR.n1817 VGND 0.01329f
C13450 VPWR.n1818 VGND 0.05634f
C13451 VPWR.t1676 VGND 0.0986f
C13452 VPWR.t622 VGND 0.05805f
C13453 VPWR.t1002 VGND 0.08842f
C13454 VPWR.n1819 VGND 0.08003f
C13455 VPWR.n1821 VGND 0.01329f
C13456 VPWR.n1822 VGND 0.10289f
C13457 VPWR.n1823 VGND 0.06176f
C13458 VPWR.n1824 VGND 0.06176f
C13459 VPWR.n1825 VGND 0.10289f
C13460 VPWR.n1826 VGND 0.01329f
C13461 VPWR.n1828 VGND 0.08003f
C13462 VPWR.t1790 VGND 0.06817f
C13463 VPWR.t975 VGND 0.05805f
C13464 VPWR.t1246 VGND 0.08842f
C13465 VPWR.n1829 VGND 0.08003f
C13466 VPWR.n1831 VGND 0.01329f
C13467 VPWR.n1832 VGND 0.10289f
C13468 VPWR.n1833 VGND 0.06176f
C13469 VPWR.n1834 VGND 0.06176f
C13470 VPWR.n1835 VGND 0.10289f
C13471 VPWR.n1836 VGND 0.01329f
C13472 VPWR.n1838 VGND 0.08003f
C13473 VPWR.t1804 VGND 0.06817f
C13474 VPWR.t627 VGND 0.05805f
C13475 VPWR.t525 VGND 0.08842f
C13476 VPWR.n1839 VGND 0.08003f
C13477 VPWR.n1841 VGND 0.01329f
C13478 VPWR.n1842 VGND 0.10289f
C13479 VPWR.n1843 VGND 0.06176f
C13480 VPWR.n1844 VGND 0.06176f
C13481 VPWR.n1845 VGND 0.10289f
C13482 VPWR.n1846 VGND 0.01329f
C13483 VPWR.n1848 VGND 0.08003f
C13484 VPWR.t381 VGND 0.06817f
C13485 VPWR.t979 VGND 0.05805f
C13486 VPWR.t1894 VGND 0.08842f
C13487 VPWR.n1849 VGND 0.08003f
C13488 VPWR.n1851 VGND 0.01329f
C13489 VPWR.n1852 VGND 0.10289f
C13490 VPWR.n1853 VGND 0.06176f
C13491 VPWR.n1854 VGND 0.06176f
C13492 VPWR.n1855 VGND 0.10289f
C13493 VPWR.n1856 VGND 0.01329f
C13494 VPWR.n1858 VGND 0.08003f
C13495 VPWR.t851 VGND 0.06817f
C13496 VPWR.t624 VGND 0.05805f
C13497 VPWR.t1736 VGND 0.08842f
C13498 VPWR.n1859 VGND 0.08003f
C13499 VPWR.n1861 VGND 0.01329f
C13500 VPWR.n1862 VGND 0.10289f
C13501 VPWR.n1863 VGND 0.06176f
C13502 VPWR.n1864 VGND 0.06176f
C13503 VPWR.n1865 VGND 0.10289f
C13504 VPWR.n1866 VGND 0.01329f
C13505 VPWR.n1868 VGND 0.08003f
C13506 VPWR.t1760 VGND 0.06817f
C13507 VPWR.t978 VGND 0.05805f
C13508 VPWR.t658 VGND 0.08842f
C13509 VPWR.n1869 VGND 0.08003f
C13510 VPWR.n1871 VGND 0.01329f
C13511 VPWR.n1872 VGND 0.10289f
C13512 VPWR.n1873 VGND 0.06176f
C13513 VPWR.n1874 VGND 0.06176f
C13514 VPWR.n1875 VGND 0.10289f
C13515 VPWR.n1876 VGND 0.01329f
C13516 VPWR.n1878 VGND 0.08003f
C13517 VPWR.t1039 VGND 0.06817f
C13518 VPWR.t1771 VGND 0.05805f
C13519 VPWR.t797 VGND 0.08842f
C13520 VPWR.n1879 VGND 0.08003f
C13521 VPWR.n1881 VGND 0.01329f
C13522 VPWR.n1882 VGND 0.10289f
C13523 VPWR.n1883 VGND 0.06176f
C13524 VPWR.n1884 VGND 0.06176f
C13525 VPWR.n1885 VGND 0.10289f
C13526 VPWR.n1886 VGND 0.01329f
C13527 VPWR.n1888 VGND 0.08003f
C13528 VPWR.t1216 VGND 0.06817f
C13529 VPWR.t980 VGND 0.05805f
C13530 VPWR.t909 VGND 0.08842f
C13531 VPWR.n1889 VGND 0.08003f
C13532 VPWR.n1891 VGND 0.01329f
C13533 VPWR.n1892 VGND 0.10289f
C13534 VPWR.n1893 VGND 0.06176f
C13535 VPWR.n1894 VGND 0.74646f
C13536 VPWR.n1895 VGND 0.14325f
C13537 VPWR.n1896 VGND 0.06176f
C13538 VPWR.n1897 VGND 0.06176f
C13539 VPWR.n1898 VGND 0.06176f
C13540 VPWR.n1899 VGND 0.06176f
C13541 VPWR.n1900 VGND 0.06176f
C13542 VPWR.n1901 VGND 0.06176f
C13543 VPWR.n1902 VGND 0.06176f
C13544 VPWR.n1903 VGND 0.06176f
C13545 VPWR.n1904 VGND 0.06176f
C13546 VPWR.n1905 VGND 0.06176f
C13547 VPWR.n1906 VGND 0.06176f
C13548 VPWR.n1907 VGND 0.06176f
C13549 VPWR.n1908 VGND 0.06176f
C13550 VPWR.n1909 VGND 0.06176f
C13551 VPWR.n1910 VGND 0.06176f
C13552 VPWR.n1911 VGND 0.74646f
C13553 VPWR.n1912 VGND 0.74646f
C13554 VPWR.n1913 VGND 0.06176f
C13555 VPWR.n1914 VGND 0.10289f
C13556 VPWR.n1915 VGND 0.01329f
C13557 VPWR.n1917 VGND 0.08003f
C13558 VPWR.t481 VGND 0.08842f
C13559 VPWR.t662 VGND 0.05805f
C13560 VPWR.t143 VGND 0.06817f
C13561 VPWR.t293 VGND 0.05805f
C13562 VPWR.t511 VGND 0.08842f
C13563 VPWR.n1918 VGND 0.08003f
C13564 VPWR.n1920 VGND 0.01329f
C13565 VPWR.n1921 VGND 0.10289f
C13566 VPWR.n1922 VGND 0.06176f
C13567 VPWR.n1923 VGND 0.06176f
C13568 VPWR.n1924 VGND 0.10289f
C13569 VPWR.n1925 VGND 0.01329f
C13570 VPWR.n1927 VGND 0.08003f
C13571 VPWR.t815 VGND 0.08842f
C13572 VPWR.t292 VGND 0.05805f
C13573 VPWR.t634 VGND 0.06817f
C13574 VPWR.t666 VGND 0.05805f
C13575 VPWR.t1330 VGND 0.08842f
C13576 VPWR.n1928 VGND 0.08003f
C13577 VPWR.n1930 VGND 0.01329f
C13578 VPWR.n1931 VGND 0.10289f
C13579 VPWR.n1932 VGND 0.06176f
C13580 VPWR.n1933 VGND 0.06176f
C13581 VPWR.n1934 VGND 0.10289f
C13582 VPWR.n1935 VGND 0.01329f
C13583 VPWR.n1937 VGND 0.08003f
C13584 VPWR.t1202 VGND 0.08842f
C13585 VPWR.t282 VGND 0.05805f
C13586 VPWR.t1812 VGND 0.06817f
C13587 VPWR.t281 VGND 0.05805f
C13588 VPWR.t59 VGND 0.08842f
C13589 VPWR.n1938 VGND 0.08003f
C13590 VPWR.n1940 VGND 0.01329f
C13591 VPWR.n1941 VGND 0.10289f
C13592 VPWR.n1942 VGND 0.06176f
C13593 VPWR.n1943 VGND 0.06176f
C13594 VPWR.n1944 VGND 0.10289f
C13595 VPWR.n1945 VGND 0.01329f
C13596 VPWR.n1947 VGND 0.08003f
C13597 VPWR.t1863 VGND 0.08842f
C13598 VPWR.t665 VGND 0.05805f
C13599 VPWR.t573 VGND 0.06817f
C13600 VPWR.t664 VGND 0.05805f
C13601 VPWR.t597 VGND 0.08842f
C13602 VPWR.n1948 VGND 0.08003f
C13603 VPWR.n1950 VGND 0.01329f
C13604 VPWR.n1951 VGND 0.10289f
C13605 VPWR.n1952 VGND 0.06176f
C13606 VPWR.n1953 VGND 0.06176f
C13607 VPWR.n1954 VGND 0.10289f
C13608 VPWR.n1955 VGND 0.01329f
C13609 VPWR.n1957 VGND 0.08003f
C13610 VPWR.t1220 VGND 0.08842f
C13611 VPWR.t283 VGND 0.05805f
C13612 VPWR.t344 VGND 0.06817f
C13613 VPWR.t291 VGND 0.05805f
C13614 VPWR.t338 VGND 0.08842f
C13615 VPWR.n1958 VGND 0.08003f
C13616 VPWR.n1960 VGND 0.01329f
C13617 VPWR.n1961 VGND 0.10289f
C13618 VPWR.n1962 VGND 0.06176f
C13619 VPWR.n1963 VGND 0.06176f
C13620 VPWR.n1964 VGND 0.10289f
C13621 VPWR.n1965 VGND 0.01329f
C13622 VPWR.n1967 VGND 0.08003f
C13623 VPWR.t1839 VGND 0.08842f
C13624 VPWR.t290 VGND 0.05805f
C13625 VPWR.t1808 VGND 0.06817f
C13626 VPWR.t296 VGND 0.05805f
C13627 VPWR.t921 VGND 0.08842f
C13628 VPWR.n1968 VGND 0.08003f
C13629 VPWR.n1970 VGND 0.01329f
C13630 VPWR.n1971 VGND 0.10289f
C13631 VPWR.n1972 VGND 0.06176f
C13632 VPWR.n1973 VGND 0.06176f
C13633 VPWR.n1974 VGND 0.10289f
C13634 VPWR.n1975 VGND 0.01329f
C13635 VPWR.n1977 VGND 0.08003f
C13636 VPWR.t1291 VGND 0.08842f
C13637 VPWR.t295 VGND 0.05805f
C13638 VPWR.t12 VGND 0.06817f
C13639 VPWR.t294 VGND 0.05805f
C13640 VPWR.t24 VGND 0.08842f
C13641 VPWR.n1978 VGND 0.08003f
C13642 VPWR.n1980 VGND 0.01329f
C13643 VPWR.n1981 VGND 0.10289f
C13644 VPWR.n1982 VGND 0.06176f
C13645 VPWR.n1983 VGND 0.06176f
C13646 VPWR.n1984 VGND 0.10289f
C13647 VPWR.n1985 VGND 0.01329f
C13648 VPWR.n1987 VGND 0.08003f
C13649 VPWR.t867 VGND 0.08842f
C13650 VPWR.t663 VGND 0.05805f
C13651 VPWR.t1384 VGND 0.0986f
C13652 VPWR.n1988 VGND 0.05634f
C13653 VPWR.n1989 VGND 0.01329f
C13654 VPWR.n1990 VGND 0.10289f
C13655 VPWR.n1991 VGND 0.14325f
C13656 VPWR.n1992 VGND 0.75117f
C13657 VPWR.n1993 VGND 0.06176f
C13658 VPWR.n1994 VGND 0.06176f
C13659 VPWR.n1995 VGND 0.06176f
C13660 VPWR.n1996 VGND 0.06176f
C13661 VPWR.n1997 VGND 0.06176f
C13662 VPWR.n1998 VGND 0.06176f
C13663 VPWR.n1999 VGND 0.06176f
C13664 VPWR.n2000 VGND 0.06176f
C13665 VPWR.n2001 VGND 0.06176f
C13666 VPWR.n2002 VGND 0.06176f
C13667 VPWR.n2003 VGND 0.06176f
C13668 VPWR.n2004 VGND 0.06176f
C13669 VPWR.n2005 VGND 0.06176f
C13670 VPWR.n2006 VGND 0.06176f
C13671 VPWR.n2007 VGND 0.06176f
C13672 VPWR.n2008 VGND 0.14325f
C13673 VPWR.n2009 VGND 0.75117f
C13674 VPWR.n2010 VGND 0.75117f
C13675 VPWR.n2011 VGND 0.14325f
C13676 VPWR.n2012 VGND 0.10289f
C13677 VPWR.n2013 VGND 0.01329f
C13678 VPWR.n2014 VGND 0.05634f
C13679 VPWR.t1456 VGND 0.0986f
C13680 VPWR.t26 VGND 0.05805f
C13681 VPWR.t183 VGND 0.08842f
C13682 VPWR.n2015 VGND 0.08003f
C13683 VPWR.n2017 VGND 0.01329f
C13684 VPWR.n2018 VGND 0.10289f
C13685 VPWR.n2019 VGND 0.06176f
C13686 VPWR.n2020 VGND 0.06176f
C13687 VPWR.n2021 VGND 0.10289f
C13688 VPWR.n2022 VGND 0.01329f
C13689 VPWR.n2024 VGND 0.08003f
C13690 VPWR.t20 VGND 0.06817f
C13691 VPWR.t1302 VGND 0.05805f
C13692 VPWR.t1279 VGND 0.08842f
C13693 VPWR.n2025 VGND 0.08003f
C13694 VPWR.n2027 VGND 0.01329f
C13695 VPWR.n2028 VGND 0.10289f
C13696 VPWR.n2029 VGND 0.06176f
C13697 VPWR.n2030 VGND 0.06176f
C13698 VPWR.n2031 VGND 0.10289f
C13699 VPWR.n2032 VGND 0.01329f
C13700 VPWR.n2034 VGND 0.08003f
C13701 VPWR.t1078 VGND 0.06817f
C13702 VPWR.t1297 VGND 0.05805f
C13703 VPWR.t1113 VGND 0.08842f
C13704 VPWR.n2035 VGND 0.08003f
C13705 VPWR.n2037 VGND 0.01329f
C13706 VPWR.n2038 VGND 0.10289f
C13707 VPWR.n2039 VGND 0.06176f
C13708 VPWR.n2040 VGND 0.06176f
C13709 VPWR.n2041 VGND 0.10289f
C13710 VPWR.n2042 VGND 0.01329f
C13711 VPWR.n2044 VGND 0.08003f
C13712 VPWR.t334 VGND 0.06817f
C13713 VPWR.t1264 VGND 0.05805f
C13714 VPWR.t855 VGND 0.08842f
C13715 VPWR.n2045 VGND 0.08003f
C13716 VPWR.n2047 VGND 0.01329f
C13717 VPWR.n2048 VGND 0.10289f
C13718 VPWR.n2049 VGND 0.06176f
C13719 VPWR.n2050 VGND 0.06176f
C13720 VPWR.n2051 VGND 0.10289f
C13721 VPWR.n2052 VGND 0.01329f
C13722 VPWR.n2054 VGND 0.08003f
C13723 VPWR.t67 VGND 0.06817f
C13724 VPWR.t28 VGND 0.05805f
C13725 VPWR.t1857 VGND 0.08842f
C13726 VPWR.n2055 VGND 0.08003f
C13727 VPWR.n2057 VGND 0.01329f
C13728 VPWR.n2058 VGND 0.10289f
C13729 VPWR.n2059 VGND 0.06176f
C13730 VPWR.n2060 VGND 0.06176f
C13731 VPWR.n2061 VGND 0.10289f
C13732 VPWR.n2062 VGND 0.01329f
C13733 VPWR.n2064 VGND 0.08003f
C13734 VPWR.t1165 VGND 0.06817f
C13735 VPWR.t1263 VGND 0.05805f
C13736 VPWR.t1127 VGND 0.08842f
C13737 VPWR.n2065 VGND 0.08003f
C13738 VPWR.n2067 VGND 0.01329f
C13739 VPWR.n2068 VGND 0.10289f
C13740 VPWR.n2069 VGND 0.06176f
C13741 VPWR.n2070 VGND 0.06176f
C13742 VPWR.n2071 VGND 0.10289f
C13743 VPWR.n2072 VGND 0.01329f
C13744 VPWR.n2074 VGND 0.08003f
C13745 VPWR.t1338 VGND 0.06817f
C13746 VPWR.t1299 VGND 0.05805f
C13747 VPWR.t823 VGND 0.08842f
C13748 VPWR.n2075 VGND 0.08003f
C13749 VPWR.n2077 VGND 0.01329f
C13750 VPWR.n2078 VGND 0.10289f
C13751 VPWR.n2079 VGND 0.06176f
C13752 VPWR.n2080 VGND 0.06176f
C13753 VPWR.n2081 VGND 0.10289f
C13754 VPWR.n2082 VGND 0.01329f
C13755 VPWR.n2084 VGND 0.08003f
C13756 VPWR.t507 VGND 0.06817f
C13757 VPWR.t1265 VGND 0.05805f
C13758 VPWR.t1724 VGND 0.08842f
C13759 VPWR.n2085 VGND 0.08003f
C13760 VPWR.n2087 VGND 0.01329f
C13761 VPWR.n2088 VGND 0.10289f
C13762 VPWR.n2089 VGND 0.06176f
C13763 VPWR.n2090 VGND 0.74646f
C13764 VPWR.n2091 VGND 0.14325f
C13765 VPWR.n2092 VGND 0.06176f
C13766 VPWR.n2093 VGND 0.06176f
C13767 VPWR.n2094 VGND 0.06176f
C13768 VPWR.n2095 VGND 0.06176f
C13769 VPWR.n2096 VGND 0.06176f
C13770 VPWR.n2097 VGND 0.06176f
C13771 VPWR.n2098 VGND 0.06176f
C13772 VPWR.n2099 VGND 0.06176f
C13773 VPWR.n2100 VGND 0.06176f
C13774 VPWR.n2101 VGND 0.06176f
C13775 VPWR.n2102 VGND 0.06176f
C13776 VPWR.n2103 VGND 0.06176f
C13777 VPWR.n2104 VGND 0.06176f
C13778 VPWR.n2105 VGND 0.06176f
C13779 VPWR.n2106 VGND 0.06176f
C13780 VPWR.n2107 VGND 0.74646f
C13781 VPWR.n2108 VGND 0.74646f
C13782 VPWR.n2109 VGND 0.06176f
C13783 VPWR.n2110 VGND 0.10289f
C13784 VPWR.n2111 VGND 0.01329f
C13785 VPWR.n2113 VGND 0.08003f
C13786 VPWR.t479 VGND 0.08842f
C13787 VPWR.t100 VGND 0.05805f
C13788 VPWR.t141 VGND 0.06817f
C13789 VPWR.t502 VGND 0.05805f
C13790 VPWR.t509 VGND 0.08842f
C13791 VPWR.n2114 VGND 0.08003f
C13792 VPWR.n2116 VGND 0.01329f
C13793 VPWR.n2117 VGND 0.10289f
C13794 VPWR.n2118 VGND 0.06176f
C13795 VPWR.n2119 VGND 0.06176f
C13796 VPWR.n2120 VGND 0.10289f
C13797 VPWR.n2121 VGND 0.01329f
C13798 VPWR.n2123 VGND 0.08003f
C13799 VPWR.t817 VGND 0.08842f
C13800 VPWR.t839 VGND 0.05805f
C13801 VPWR.t687 VGND 0.06817f
C13802 VPWR.t567 VGND 0.05805f
C13803 VPWR.t379 VGND 0.08842f
C13804 VPWR.n2124 VGND 0.08003f
C13805 VPWR.n2126 VGND 0.01329f
C13806 VPWR.n2127 VGND 0.10289f
C13807 VPWR.n2128 VGND 0.06176f
C13808 VPWR.n2129 VGND 0.06176f
C13809 VPWR.n2130 VGND 0.10289f
C13810 VPWR.n2131 VGND 0.01329f
C13811 VPWR.n2133 VGND 0.08003f
C13812 VPWR.t139 VGND 0.08842f
C13813 VPWR.t319 VGND 0.05805f
C13814 VPWR.t63 VGND 0.06817f
C13815 VPWR.t318 VGND 0.05805f
C13816 VPWR.t57 VGND 0.08842f
C13817 VPWR.n2134 VGND 0.08003f
C13818 VPWR.n2136 VGND 0.01329f
C13819 VPWR.n2137 VGND 0.10289f
C13820 VPWR.n2138 VGND 0.06176f
C13821 VPWR.n2139 VGND 0.06176f
C13822 VPWR.n2140 VGND 0.10289f
C13823 VPWR.n2141 VGND 0.01329f
C13824 VPWR.n2143 VGND 0.08003f
C13825 VPWR.t1861 VGND 0.08842f
C13826 VPWR.t566 VGND 0.05805f
C13827 VPWR.t571 VGND 0.06817f
C13828 VPWR.t565 VGND 0.05805f
C13829 VPWR.t595 VGND 0.08842f
C13830 VPWR.n2144 VGND 0.08003f
C13831 VPWR.n2146 VGND 0.01329f
C13832 VPWR.n2147 VGND 0.10289f
C13833 VPWR.n2148 VGND 0.06176f
C13834 VPWR.n2149 VGND 0.06176f
C13835 VPWR.n2150 VGND 0.10289f
C13836 VPWR.n2151 VGND 0.01329f
C13837 VPWR.n2153 VGND 0.08003f
C13838 VPWR.t1218 VGND 0.08842f
C13839 VPWR.t320 VGND 0.05805f
C13840 VPWR.t342 VGND 0.06817f
C13841 VPWR.t838 VGND 0.05805f
C13842 VPWR.t336 VGND 0.08842f
C13843 VPWR.n2154 VGND 0.08003f
C13844 VPWR.n2156 VGND 0.01329f
C13845 VPWR.n2157 VGND 0.10289f
C13846 VPWR.n2158 VGND 0.06176f
C13847 VPWR.n2159 VGND 0.06176f
C13848 VPWR.n2160 VGND 0.10289f
C13849 VPWR.n2161 VGND 0.01329f
C13850 VPWR.n2163 VGND 0.08003f
C13851 VPWR.t1837 VGND 0.08842f
C13852 VPWR.t837 VGND 0.05805f
C13853 VPWR.t1806 VGND 0.06817f
C13854 VPWR.t317 VGND 0.05805f
C13855 VPWR.t919 VGND 0.08842f
C13856 VPWR.n2164 VGND 0.08003f
C13857 VPWR.n2166 VGND 0.01329f
C13858 VPWR.n2167 VGND 0.10289f
C13859 VPWR.n2168 VGND 0.06176f
C13860 VPWR.n2169 VGND 0.06176f
C13861 VPWR.n2170 VGND 0.10289f
C13862 VPWR.n2171 VGND 0.01329f
C13863 VPWR.n2173 VGND 0.08003f
C13864 VPWR.t1289 VGND 0.08842f
C13865 VPWR.t504 VGND 0.05805f
C13866 VPWR.t10 VGND 0.06817f
C13867 VPWR.t503 VGND 0.05805f
C13868 VPWR.t22 VGND 0.08842f
C13869 VPWR.n2174 VGND 0.08003f
C13870 VPWR.n2176 VGND 0.01329f
C13871 VPWR.n2177 VGND 0.10289f
C13872 VPWR.n2178 VGND 0.06176f
C13873 VPWR.n2179 VGND 0.06176f
C13874 VPWR.n2180 VGND 0.10289f
C13875 VPWR.n2181 VGND 0.01329f
C13876 VPWR.n2183 VGND 0.08003f
C13877 VPWR.t165 VGND 0.08842f
C13878 VPWR.t101 VGND 0.05805f
C13879 VPWR.t1389 VGND 0.0986f
C13880 VPWR.n2184 VGND 0.05634f
C13881 VPWR.n2185 VGND 0.01329f
C13882 VPWR.n2186 VGND 0.10289f
C13883 VPWR.n2187 VGND 0.14325f
C13884 VPWR.n2188 VGND 0.75117f
C13885 VPWR.n2189 VGND 0.06176f
C13886 VPWR.n2190 VGND 0.06176f
C13887 VPWR.n2191 VGND 0.06176f
C13888 VPWR.n2192 VGND 0.06176f
C13889 VPWR.n2193 VGND 0.06176f
C13890 VPWR.n2194 VGND 0.06176f
C13891 VPWR.n2195 VGND 0.06176f
C13892 VPWR.n2196 VGND 0.06176f
C13893 VPWR.n2197 VGND 0.06176f
C13894 VPWR.n2198 VGND 0.06176f
C13895 VPWR.n2199 VGND 0.06176f
C13896 VPWR.n2200 VGND 0.06176f
C13897 VPWR.n2201 VGND 0.06176f
C13898 VPWR.n2202 VGND 0.06176f
C13899 VPWR.n2203 VGND 0.06176f
C13900 VPWR.n2204 VGND 0.14325f
C13901 VPWR.n2205 VGND 0.75117f
C13902 VPWR.n2206 VGND 0.75117f
C13903 VPWR.n2207 VGND 0.14325f
C13904 VPWR.n2208 VGND 0.10289f
C13905 VPWR.n2209 VGND 0.01329f
C13906 VPWR.n2210 VGND 0.05634f
C13907 VPWR.t1555 VGND 0.0986f
C13908 VPWR.t865 VGND 0.05805f
C13909 VPWR.t203 VGND 0.08842f
C13910 VPWR.n2211 VGND 0.08003f
C13911 VPWR.n2213 VGND 0.01329f
C13912 VPWR.n2214 VGND 0.10289f
C13913 VPWR.n2215 VGND 0.06176f
C13914 VPWR.n2216 VGND 0.06176f
C13915 VPWR.n2217 VGND 0.10289f
C13916 VPWR.n2218 VGND 0.01329f
C13917 VPWR.n2220 VGND 0.08003f
C13918 VPWR.t41 VGND 0.06817f
C13919 VPWR.t859 VGND 0.05805f
C13920 VPWR.t971 VGND 0.08842f
C13921 VPWR.n2221 VGND 0.08003f
C13922 VPWR.n2223 VGND 0.01329f
C13923 VPWR.n2224 VGND 0.10289f
C13924 VPWR.n2225 VGND 0.06176f
C13925 VPWR.n2226 VGND 0.06176f
C13926 VPWR.n2227 VGND 0.10289f
C13927 VPWR.n2228 VGND 0.01329f
C13928 VPWR.n2230 VGND 0.08003f
C13929 VPWR.t1149 VGND 0.06817f
C13930 VPWR.t1773 VGND 0.05805f
C13931 VPWR.t706 VGND 0.08842f
C13932 VPWR.n2231 VGND 0.08003f
C13933 VPWR.n2233 VGND 0.01329f
C13934 VPWR.n2234 VGND 0.10289f
C13935 VPWR.n2235 VGND 0.06176f
C13936 VPWR.n2236 VGND 0.06176f
C13937 VPWR.n2237 VGND 0.10289f
C13938 VPWR.n2238 VGND 0.01329f
C13939 VPWR.n2240 VGND 0.08003f
C13940 VPWR.t427 VGND 0.06817f
C13941 VPWR.t863 VGND 0.05805f
C13942 VPWR.t519 VGND 0.08842f
C13943 VPWR.n2241 VGND 0.08003f
C13944 VPWR.n2243 VGND 0.01329f
C13945 VPWR.n2244 VGND 0.10289f
C13946 VPWR.n2245 VGND 0.06176f
C13947 VPWR.n2246 VGND 0.06176f
C13948 VPWR.n2247 VGND 0.10289f
C13949 VPWR.n2248 VGND 0.01329f
C13950 VPWR.n2250 VGND 0.08003f
C13951 VPWR.t6 VGND 0.06817f
C13952 VPWR.t999 VGND 0.05805f
C13953 VPWR.t491 VGND 0.08842f
C13954 VPWR.n2251 VGND 0.08003f
C13955 VPWR.n2253 VGND 0.01329f
C13956 VPWR.n2254 VGND 0.10289f
C13957 VPWR.n2255 VGND 0.06176f
C13958 VPWR.n2256 VGND 0.06176f
C13959 VPWR.n2257 VGND 0.10289f
C13960 VPWR.n2258 VGND 0.01329f
C13961 VPWR.n2260 VGND 0.08003f
C13962 VPWR.t1170 VGND 0.06817f
C13963 VPWR.t862 VGND 0.05805f
C13964 VPWR.t1320 VGND 0.08842f
C13965 VPWR.n2261 VGND 0.08003f
C13966 VPWR.n2263 VGND 0.01329f
C13967 VPWR.n2264 VGND 0.10289f
C13968 VPWR.n2265 VGND 0.06176f
C13969 VPWR.n2266 VGND 0.06176f
C13970 VPWR.n2267 VGND 0.10289f
C13971 VPWR.n2268 VGND 0.01329f
C13972 VPWR.n2270 VGND 0.08003f
C13973 VPWR.t375 VGND 0.06817f
C13974 VPWR.t1775 VGND 0.05805f
C13975 VPWR.t781 VGND 0.08842f
C13976 VPWR.n2271 VGND 0.08003f
C13977 VPWR.n2273 VGND 0.01329f
C13978 VPWR.n2274 VGND 0.10289f
C13979 VPWR.n2275 VGND 0.06176f
C13980 VPWR.n2276 VGND 0.06176f
C13981 VPWR.n2277 VGND 0.10289f
C13982 VPWR.n2278 VGND 0.01329f
C13983 VPWR.n2280 VGND 0.08003f
C13984 VPWR.t267 VGND 0.06817f
C13985 VPWR.t864 VGND 0.05805f
C13986 VPWR.t1910 VGND 0.08842f
C13987 VPWR.n2281 VGND 0.08003f
C13988 VPWR.n2283 VGND 0.01329f
C13989 VPWR.n2284 VGND 0.10289f
C13990 VPWR.n2285 VGND 0.06176f
C13991 VPWR.n2286 VGND 0.74646f
C13992 VPWR.n2287 VGND 0.14325f
C13993 VPWR.n2288 VGND 0.06176f
C13994 VPWR.n2289 VGND 0.06176f
C13995 VPWR.n2290 VGND 0.06176f
C13996 VPWR.n2291 VGND 0.06176f
C13997 VPWR.n2292 VGND 0.06176f
C13998 VPWR.n2293 VGND 0.06176f
C13999 VPWR.n2294 VGND 0.06176f
C14000 VPWR.n2295 VGND 0.06176f
C14001 VPWR.n2296 VGND 0.06176f
C14002 VPWR.n2297 VGND 0.06176f
C14003 VPWR.n2298 VGND 0.06176f
C14004 VPWR.n2299 VGND 0.06176f
C14005 VPWR.n2300 VGND 0.06176f
C14006 VPWR.n2301 VGND 0.06176f
C14007 VPWR.n2302 VGND 0.06176f
C14008 VPWR.n2303 VGND 0.74646f
C14009 VPWR.n2304 VGND 0.74646f
C14010 VPWR.n2305 VGND 0.06176f
C14011 VPWR.n2306 VGND 0.10289f
C14012 VPWR.n2307 VGND 0.01329f
C14013 VPWR.n2309 VGND 0.08003f
C14014 VPWR.t957 VGND 0.08842f
C14015 VPWR.t130 VGND 0.05805f
C14016 VPWR.t1133 VGND 0.06817f
C14017 VPWR.t1823 VGND 0.05805f
C14018 VPWR.t1129 VGND 0.08842f
C14019 VPWR.n2310 VGND 0.08003f
C14020 VPWR.n2312 VGND 0.01329f
C14021 VPWR.n2313 VGND 0.10289f
C14022 VPWR.n2314 VGND 0.06176f
C14023 VPWR.n2315 VGND 0.06176f
C14024 VPWR.n2316 VGND 0.10289f
C14025 VPWR.n2317 VGND 0.01329f
C14026 VPWR.n2319 VGND 0.08003f
C14027 VPWR.t827 VGND 0.08842f
C14028 VPWR.t1822 VGND 0.05805f
C14029 VPWR.t1336 VGND 0.06817f
C14030 VPWR.t1267 VGND 0.05805f
C14031 VPWR.t153 VGND 0.08842f
C14032 VPWR.n2320 VGND 0.08003f
C14033 VPWR.n2322 VGND 0.01329f
C14034 VPWR.n2323 VGND 0.10289f
C14035 VPWR.n2324 VGND 0.06176f
C14036 VPWR.n2325 VGND 0.06176f
C14037 VPWR.n2326 VGND 0.10289f
C14038 VPWR.n2327 VGND 0.01329f
C14039 VPWR.n2329 VGND 0.08003f
C14040 VPWR.t1121 VGND 0.08842f
C14041 VPWR.t454 VGND 0.05805f
C14042 VPWR.t1161 VGND 0.06817f
C14043 VPWR.t453 VGND 0.05805f
C14044 VPWR.t1176 VGND 0.08842f
C14045 VPWR.n2330 VGND 0.08003f
C14046 VPWR.n2332 VGND 0.01329f
C14047 VPWR.n2333 VGND 0.10289f
C14048 VPWR.n2334 VGND 0.06176f
C14049 VPWR.n2335 VGND 0.06176f
C14050 VPWR.n2336 VGND 0.10289f
C14051 VPWR.n2337 VGND 0.01329f
C14052 VPWR.n2339 VGND 0.08003f
C14053 VPWR.t1256 VGND 0.08842f
C14054 VPWR.t1266 VGND 0.05805f
C14055 VPWR.t603 VGND 0.06817f
C14056 VPWR.t132 VGND 0.05805f
C14057 VPWR.t736 VGND 0.08842f
C14058 VPWR.n2340 VGND 0.08003f
C14059 VPWR.n2342 VGND 0.01329f
C14060 VPWR.n2343 VGND 0.10289f
C14061 VPWR.n2344 VGND 0.06176f
C14062 VPWR.n2345 VGND 0.06176f
C14063 VPWR.n2346 VGND 0.10289f
C14064 VPWR.n2347 VGND 0.01329f
C14065 VPWR.n2349 VGND 0.08003f
C14066 VPWR.t579 VGND 0.08842f
C14067 VPWR.t455 VGND 0.05805f
C14068 VPWR.t439 VGND 0.06817f
C14069 VPWR.t1821 VGND 0.05805f
C14070 VPWR.t431 VGND 0.08842f
C14071 VPWR.n2350 VGND 0.08003f
C14072 VPWR.n2352 VGND 0.01329f
C14073 VPWR.n2353 VGND 0.10289f
C14074 VPWR.n2354 VGND 0.06176f
C14075 VPWR.n2355 VGND 0.06176f
C14076 VPWR.n2356 VGND 0.10289f
C14077 VPWR.n2357 VGND 0.01329f
C14078 VPWR.n2359 VGND 0.08003f
C14079 VPWR.t1914 VGND 0.08842f
C14080 VPWR.t1820 VGND 0.05805f
C14081 VPWR.t94 VGND 0.06817f
C14082 VPWR.t452 VGND 0.05805f
C14083 VPWR.t1780 VGND 0.08842f
C14084 VPWR.n2360 VGND 0.08003f
C14085 VPWR.n2362 VGND 0.01329f
C14086 VPWR.n2363 VGND 0.10289f
C14087 VPWR.n2364 VGND 0.06176f
C14088 VPWR.n2365 VGND 0.06176f
C14089 VPWR.n2366 VGND 0.10289f
C14090 VPWR.n2367 VGND 0.01329f
C14091 VPWR.n2369 VGND 0.08003f
C14092 VPWR.t545 VGND 0.08842f
C14093 VPWR.t451 VGND 0.05805f
C14094 VPWR.t891 VGND 0.06817f
C14095 VPWR.t450 VGND 0.05805f
C14096 VPWR.t883 VGND 0.08842f
C14097 VPWR.n2370 VGND 0.08003f
C14098 VPWR.n2372 VGND 0.01329f
C14099 VPWR.n2373 VGND 0.10289f
C14100 VPWR.n2374 VGND 0.06176f
C14101 VPWR.n2375 VGND 0.06176f
C14102 VPWR.n2376 VGND 0.10289f
C14103 VPWR.n2377 VGND 0.01329f
C14104 VPWR.n2379 VGND 0.08003f
C14105 VPWR.t181 VGND 0.08842f
C14106 VPWR.t131 VGND 0.05805f
C14107 VPWR.t1488 VGND 0.0986f
C14108 VPWR.n2380 VGND 0.05634f
C14109 VPWR.n2381 VGND 0.01329f
C14110 VPWR.n2382 VGND 0.10289f
C14111 VPWR.n2383 VGND 0.14325f
C14112 VPWR.n2384 VGND 0.75117f
C14113 VPWR.n2385 VGND 0.06176f
C14114 VPWR.n2386 VGND 0.06176f
C14115 VPWR.n2387 VGND 0.06176f
C14116 VPWR.n2388 VGND 0.06176f
C14117 VPWR.n2389 VGND 0.06176f
C14118 VPWR.n2390 VGND 0.06176f
C14119 VPWR.n2391 VGND 0.06176f
C14120 VPWR.n2392 VGND 0.06176f
C14121 VPWR.n2393 VGND 0.06176f
C14122 VPWR.n2394 VGND 0.06176f
C14123 VPWR.n2395 VGND 0.06176f
C14124 VPWR.n2396 VGND 0.06176f
C14125 VPWR.n2397 VGND 0.06176f
C14126 VPWR.n2398 VGND 0.06176f
C14127 VPWR.n2399 VGND 0.06176f
C14128 VPWR.n2400 VGND 0.14325f
C14129 VPWR.n2401 VGND 0.75117f
C14130 VPWR.n2402 VGND 0.75117f
C14131 VPWR.n2403 VGND 0.14325f
C14132 VPWR.n2404 VGND 0.10289f
C14133 VPWR.n2405 VGND 0.01329f
C14134 VPWR.n2406 VGND 0.05634f
C14135 VPWR.t1658 VGND 0.0986f
C14136 VPWR.t1181 VGND 0.05805f
C14137 VPWR.t1008 VGND 0.08842f
C14138 VPWR.n2407 VGND 0.08003f
C14139 VPWR.n2409 VGND 0.01329f
C14140 VPWR.n2410 VGND 0.10289f
C14141 VPWR.n2411 VGND 0.06176f
C14142 VPWR.n2412 VGND 0.06176f
C14143 VPWR.n2413 VGND 0.10289f
C14144 VPWR.n2414 VGND 0.01329f
C14145 VPWR.n2416 VGND 0.08003f
C14146 VPWR.t1024 VGND 0.06817f
C14147 VPWR.t456 VGND 0.05805f
C14148 VPWR.t1250 VGND 0.08842f
C14149 VPWR.n2417 VGND 0.08003f
C14150 VPWR.n2419 VGND 0.01329f
C14151 VPWR.n2420 VGND 0.10289f
C14152 VPWR.n2421 VGND 0.06176f
C14153 VPWR.n2422 VGND 0.06176f
C14154 VPWR.n2423 VGND 0.10289f
C14155 VPWR.n2424 VGND 0.01329f
C14156 VPWR.n2426 VGND 0.08003f
C14157 VPWR.t1157 VGND 0.06817f
C14158 VPWR.t1922 VGND 0.05805f
C14159 VPWR.t531 VGND 0.08842f
C14160 VPWR.n2427 VGND 0.08003f
C14161 VPWR.n2429 VGND 0.01329f
C14162 VPWR.n2430 VGND 0.10289f
C14163 VPWR.n2431 VGND 0.06176f
C14164 VPWR.n2432 VGND 0.06176f
C14165 VPWR.n2433 VGND 0.10289f
C14166 VPWR.n2434 VGND 0.01329f
C14167 VPWR.n2436 VGND 0.08003f
C14168 VPWR.t385 VGND 0.06817f
C14169 VPWR.t460 VGND 0.05805f
C14170 VPWR.t1900 VGND 0.08842f
C14171 VPWR.n2437 VGND 0.08003f
C14172 VPWR.n2439 VGND 0.01329f
C14173 VPWR.n2440 VGND 0.10289f
C14174 VPWR.n2441 VGND 0.06176f
C14175 VPWR.n2442 VGND 0.06176f
C14176 VPWR.n2443 VGND 0.10289f
C14177 VPWR.n2444 VGND 0.01329f
C14178 VPWR.n2446 VGND 0.08003f
C14179 VPWR.t288 VGND 0.06817f
C14180 VPWR.t1183 VGND 0.05805f
C14181 VPWR.t1742 VGND 0.08842f
C14182 VPWR.n2447 VGND 0.08003f
C14183 VPWR.n2449 VGND 0.01329f
C14184 VPWR.n2450 VGND 0.10289f
C14185 VPWR.n2451 VGND 0.06176f
C14186 VPWR.n2452 VGND 0.06176f
C14187 VPWR.n2453 VGND 0.10289f
C14188 VPWR.n2454 VGND 0.01329f
C14189 VPWR.n2456 VGND 0.08003f
C14190 VPWR.t695 VGND 0.06817f
C14191 VPWR.t459 VGND 0.05805f
C14192 VPWR.t401 VGND 0.08842f
C14193 VPWR.n2457 VGND 0.08003f
C14194 VPWR.n2459 VGND 0.01329f
C14195 VPWR.n2460 VGND 0.10289f
C14196 VPWR.n2461 VGND 0.06176f
C14197 VPWR.n2462 VGND 0.06176f
C14198 VPWR.n2463 VGND 0.10289f
C14199 VPWR.n2464 VGND 0.01329f
C14200 VPWR.n2466 VGND 0.08003f
C14201 VPWR.t1045 VGND 0.06817f
C14202 VPWR.t1924 VGND 0.05805f
C14203 VPWR.t793 VGND 0.08842f
C14204 VPWR.n2467 VGND 0.08003f
C14205 VPWR.n2469 VGND 0.01329f
C14206 VPWR.n2470 VGND 0.10289f
C14207 VPWR.n2471 VGND 0.06176f
C14208 VPWR.n2472 VGND 0.06176f
C14209 VPWR.n2473 VGND 0.10289f
C14210 VPWR.n2474 VGND 0.01329f
C14211 VPWR.n2476 VGND 0.08003f
C14212 VPWR.t1139 VGND 0.06817f
C14213 VPWR.t1180 VGND 0.05805f
C14214 VPWR.t899 VGND 0.08842f
C14215 VPWR.n2477 VGND 0.08003f
C14216 VPWR.n2479 VGND 0.01329f
C14217 VPWR.n2480 VGND 0.10289f
C14218 VPWR.n2481 VGND 0.06176f
C14219 VPWR.n2482 VGND 0.74646f
C14220 VPWR.n2483 VGND 0.14325f
C14221 VPWR.n2484 VGND 0.06176f
C14222 VPWR.n2485 VGND 0.06176f
C14223 VPWR.n2486 VGND 0.06176f
C14224 VPWR.n2487 VGND 0.06176f
C14225 VPWR.n2488 VGND 0.06176f
C14226 VPWR.n2489 VGND 0.06176f
C14227 VPWR.n2490 VGND 0.06176f
C14228 VPWR.n2491 VGND 0.06176f
C14229 VPWR.n2492 VGND 0.06176f
C14230 VPWR.n2493 VGND 0.06176f
C14231 VPWR.n2494 VGND 0.06176f
C14232 VPWR.n2495 VGND 0.06176f
C14233 VPWR.n2496 VGND 0.06176f
C14234 VPWR.n2497 VGND 0.06176f
C14235 VPWR.n2498 VGND 0.06176f
C14236 VPWR.n2499 VGND 0.74646f
C14237 VPWR.n2500 VGND 0.42248f
C14238 VPWR.n2501 VGND 0.06176f
C14239 VPWR.n2502 VGND 0.064f
C14240 VPWR.n2504 VGND 0.01268f
C14241 VPWR.n2506 VGND 0.08003f
C14242 VPWR.t1537 VGND 0.08842f
C14243 VPWR.t1504 VGND 0.05805f
C14244 VPWR.t1628 VGND 0.06817f
C14245 VPWR.t1634 VGND 0.05805f
C14246 VPWR.t1649 VGND 0.08842f
C14247 VPWR.n2507 VGND 0.08003f
C14248 VPWR.n2509 VGND 0.01268f
C14249 VPWR.n2511 VGND 0.064f
C14250 VPWR.n2512 VGND 0.06176f
C14251 VPWR.n2513 VGND 0.06176f
C14252 VPWR.n2514 VGND 0.064f
C14253 VPWR.n2516 VGND 0.01268f
C14254 VPWR.n2518 VGND 0.08003f
C14255 VPWR.t1414 VGND 0.08842f
C14256 VPWR.t1674 VGND 0.05805f
C14257 VPWR.t1408 VGND 0.06817f
C14258 VPWR.t1398 VGND 0.05805f
C14259 VPWR.t1525 VGND 0.08842f
C14260 VPWR.n2519 VGND 0.08003f
C14261 VPWR.n2521 VGND 0.01268f
C14262 VPWR.n2523 VGND 0.064f
C14263 VPWR.n2524 VGND 0.06176f
C14264 VPWR.n2525 VGND 0.06176f
C14265 VPWR.n2526 VGND 0.064f
C14266 VPWR.n2528 VGND 0.01268f
C14267 VPWR.n2530 VGND 0.08003f
C14268 VPWR.t1534 VGND 0.08842f
C14269 VPWR.t1542 VGND 0.05805f
C14270 VPWR.t1671 VGND 0.06817f
C14271 VPWR.t1566 VGND 0.05805f
C14272 VPWR.t1690 VGND 0.08842f
C14273 VPWR.n2531 VGND 0.08003f
C14274 VPWR.n2533 VGND 0.01268f
C14275 VPWR.n2535 VGND 0.064f
C14276 VPWR.n2536 VGND 0.06176f
C14277 VPWR.n2537 VGND 0.06176f
C14278 VPWR.n2538 VGND 0.064f
C14279 VPWR.n2540 VGND 0.01268f
C14280 VPWR.n2542 VGND 0.08003f
C14281 VPWR.t1411 VGND 0.08842f
C14282 VPWR.t1403 VGND 0.05805f
C14283 VPWR.t1430 VGND 0.06817f
C14284 VPWR.t1438 VGND 0.05805f
C14285 VPWR.t1571 VGND 0.08842f
C14286 VPWR.n2543 VGND 0.08003f
C14287 VPWR.n2545 VGND 0.01268f
C14288 VPWR.n2547 VGND 0.064f
C14289 VPWR.n2548 VGND 0.06176f
C14290 VPWR.n2549 VGND 0.06176f
C14291 VPWR.n2550 VGND 0.064f
C14292 VPWR.n2552 VGND 0.01268f
C14293 VPWR.n2554 VGND 0.08003f
C14294 VPWR.t1587 VGND 0.08842f
C14295 VPWR.t1540 VGND 0.05805f
C14296 VPWR.t1668 VGND 0.06817f
C14297 VPWR.t1701 VGND 0.05805f
C14298 VPWR.t1717 VGND 0.08842f
C14299 VPWR.n2555 VGND 0.08003f
C14300 VPWR.n2557 VGND 0.01268f
C14301 VPWR.n2559 VGND 0.064f
C14302 VPWR.n2560 VGND 0.06176f
C14303 VPWR.n2561 VGND 0.06176f
C14304 VPWR.n2562 VGND 0.064f
C14305 VPWR.n2564 VGND 0.01268f
C14306 VPWR.n2566 VGND 0.08003f
C14307 VPWR.t1461 VGND 0.08842f
C14308 VPWR.t1720 VGND 0.05805f
C14309 VPWR.t1453 VGND 0.06817f
C14310 VPWR.t1574 VGND 0.05805f
C14311 VPWR.t1491 VGND 0.08842f
C14312 VPWR.n2567 VGND 0.08003f
C14313 VPWR.n2569 VGND 0.01268f
C14314 VPWR.n2571 VGND 0.064f
C14315 VPWR.n2572 VGND 0.06176f
C14316 VPWR.n2573 VGND 0.06176f
C14317 VPWR.n2574 VGND 0.064f
C14318 VPWR.n2576 VGND 0.01268f
C14319 VPWR.n2578 VGND 0.08003f
C14320 VPWR.t1341 VGND 0.08842f
C14321 VPWR.t1593 VGND 0.05805f
C14322 VPWR.t1714 VGND 0.06817f
C14323 VPWR.t1618 VGND 0.05805f
C14324 VPWR.t1360 VGND 0.08842f
C14325 VPWR.n2579 VGND 0.08003f
C14326 VPWR.n2581 VGND 0.01268f
C14327 VPWR.n2583 VGND 0.064f
C14328 VPWR.n2584 VGND 0.06176f
C14329 VPWR.n2585 VGND 0.06176f
C14330 VPWR.n2586 VGND 0.064f
C14331 VPWR.n2588 VGND 0.01268f
C14332 VPWR.n2590 VGND 0.08003f
C14333 VPWR.t1485 VGND 0.08842f
C14334 VPWR.t1469 VGND 0.05805f
C14335 VPWR.t1590 VGND 0.0986f
C14336 VPWR.n2591 VGND 0.05631f
C14337 VPWR.n2592 VGND 0.01256f
C14338 VPWR.n2594 VGND 0.08026f
C14339 VPWR.n2595 VGND 0.14325f
C14340 VPWR.n2596 VGND 1.96905f
C14341 VPWR.n2597 VGND 0.80188f
C14342 VPWR.n2598 VGND 0.33599f
C14343 VPWR.t117 VGND 0.04034f
C14344 VPWR.t989 VGND 0.04034f
C14345 VPWR.n2599 VGND 0.07319f
C14346 VPWR.n2600 VGND 0.03466f
C14347 VPWR.t115 VGND 0.0106f
C14348 VPWR.t123 VGND 0.0106f
C14349 VPWR.n2601 VGND 0.02274f
C14350 VPWR.t994 VGND 0.0106f
C14351 VPWR.t988 VGND 0.0106f
C14352 VPWR.n2602 VGND 0.02274f
C14353 VPWR.n2604 VGND 0.03466f
C14354 VPWR.t1830 VGND 0.0106f
C14355 VPWR.t246 VGND 0.0106f
C14356 VPWR.n2605 VGND 0.02274f
C14357 VPWR.t240 VGND 0.0106f
C14358 VPWR.t325 VGND 0.0106f
C14359 VPWR.n2606 VGND 0.02274f
C14360 VPWR.t252 VGND 0.04225f
C14361 VPWR.t298 VGND 0.04225f
C14362 VPWR.n2607 VGND 0.09744f
C14363 VPWR.n2608 VGND 0.03127f
C14364 VPWR.n2609 VGND 0.01007f
C14365 VPWR.n2610 VGND 0.04572f
C14366 VPWR.t297 VGND 0.0106f
C14367 VPWR.t121 VGND 0.0106f
C14368 VPWR.n2612 VGND 0.02274f
C14369 VPWR.t254 VGND 0.0106f
C14370 VPWR.t992 VGND 0.0106f
C14371 VPWR.n2613 VGND 0.02274f
C14372 VPWR.n2614 VGND 0.04572f
C14373 VPWR.n2615 VGND 0.01054f
C14374 VPWR.n2616 VGND 0.03466f
C14375 VPWR.n2617 VGND 0.03466f
C14376 VPWR.n2618 VGND 0.03466f
C14377 VPWR.n2620 VGND 0.04572f
C14378 VPWR.n2623 VGND 0.03466f
C14379 VPWR.n2624 VGND 0.02599f
C14380 VPWR.t251 VGND 0.1266f
C14381 VPWR.t239 VGND 0.18657f
C14382 VPWR.t245 VGND 0.18657f
C14383 VPWR.t253 VGND 0.18657f
C14384 VPWR.t120 VGND 0.18657f
C14385 VPWR.t114 VGND 0.18657f
C14386 VPWR.t122 VGND 0.18657f
C14387 VPWR.t116 VGND 0.41537f
C14388 VPWR.n2626 VGND 0.45337f
C14389 VPWR.n2627 VGND 0.01319f
C14390 VPWR.n2628 VGND 0.7952f
C14391 VPWR.n2629 VGND 0.03466f
C14392 VPWR.t299 VGND 0.1266f
C14393 VPWR.t235 VGND 0.18657f
C14394 VPWR.t214 VGND 0.18657f
C14395 VPWR.t270 VGND 0.18657f
C14396 VPWR.t461 VGND 0.18657f
C14397 VPWR.t471 VGND 0.18657f
C14398 VPWR.t463 VGND 0.18657f
C14399 VPWR.t473 VGND 0.30651f
C14400 VPWR.t738 VGND 0.32539f
C14401 VPWR.n2630 VGND 0.45918f
C14402 VPWR.n2631 VGND 0.13062f
C14403 VPWR.n2632 VGND 0.03466f
C14404 VPWR.t472 VGND 0.0106f
C14405 VPWR.t464 VGND 0.0106f
C14406 VPWR.n2633 VGND 0.02274f
C14407 VPWR.t750 VGND 0.0106f
C14408 VPWR.t756 VGND 0.0106f
C14409 VPWR.n2634 VGND 0.02274f
C14410 VPWR.n2635 VGND 0.04572f
C14411 VPWR.n2636 VGND 0.03466f
C14412 VPWR.t314 VGND 0.0106f
C14413 VPWR.t462 VGND 0.0106f
C14414 VPWR.n2637 VGND 0.02274f
C14415 VPWR.t271 VGND 0.0106f
C14416 VPWR.t754 VGND 0.0106f
C14417 VPWR.n2638 VGND 0.02274f
C14418 VPWR.t300 VGND 0.04225f
C14419 VPWR.t315 VGND 0.04225f
C14420 VPWR.n2640 VGND 0.09744f
C14421 VPWR.t280 VGND 0.0106f
C14422 VPWR.t242 VGND 0.0106f
C14423 VPWR.n2641 VGND 0.02274f
C14424 VPWR.t236 VGND 0.0106f
C14425 VPWR.t215 VGND 0.0106f
C14426 VPWR.n2642 VGND 0.02274f
C14427 VPWR.n2643 VGND 0.04572f
C14428 VPWR.n2644 VGND 0.01007f
C14429 VPWR.n2645 VGND 0.03127f
C14430 VPWR.n2646 VGND 0.03466f
C14431 VPWR.n2647 VGND 0.03466f
C14432 VPWR.n2648 VGND 0.01054f
C14433 VPWR.n2649 VGND 0.04572f
C14434 VPWR.n2652 VGND 0.03466f
C14435 VPWR.n2653 VGND 0.03466f
C14436 VPWR.t474 VGND 0.04034f
C14437 VPWR.t752 VGND 0.04034f
C14438 VPWR.n2656 VGND 0.07319f
C14439 VPWR.n2658 VGND 0.02599f
C14440 VPWR.n2659 VGND 0.01319f
C14441 VPWR.n2660 VGND 0.02599f
C14442 VPWR.n2661 VGND 0.01034f
C14443 VPWR.t840 VGND 0.04221f
C14444 VPWR.t739 VGND 0.04221f
C14445 VPWR.n2663 VGND 0.08532f
C14446 VPWR.n2664 VGND 0.02411f
C14447 VPWR.n2665 VGND 1.21026f
C14448 VPWR.n2666 VGND 0.03466f
C14449 VPWR.t1853 VGND 0.04143f
C14450 VPWR.t276 VGND 0.1266f
C14451 VPWR.t226 VGND 0.18657f
C14452 VPWR.t309 VGND 0.18657f
C14453 VPWR.t274 VGND 0.18657f
C14454 VPWR.t648 VGND 0.18657f
C14455 VPWR.t642 VGND 0.18657f
C14456 VPWR.t650 VGND 0.18657f
C14457 VPWR.t644 VGND 0.30651f
C14458 VPWR.t1233 VGND 0.11772f
C14459 VPWR.t1852 VGND 0.09329f
C14460 VPWR.t135 VGND 0.20767f
C14461 VPWR.n2667 VGND 0.40698f
C14462 VPWR.n2668 VGND 0.12868f
C14463 VPWR.n2669 VGND 0.03466f
C14464 VPWR.t927 VGND 0.0106f
C14465 VPWR.t931 VGND 0.0106f
C14466 VPWR.n2670 VGND 0.02274f
C14467 VPWR.t643 VGND 0.0106f
C14468 VPWR.t651 VGND 0.0106f
C14469 VPWR.n2671 VGND 0.02274f
C14470 VPWR.n2672 VGND 0.04572f
C14471 VPWR.n2673 VGND 0.03466f
C14472 VPWR.t275 VGND 0.0106f
C14473 VPWR.t930 VGND 0.0106f
C14474 VPWR.n2674 VGND 0.02274f
C14475 VPWR.t324 VGND 0.0106f
C14476 VPWR.t649 VGND 0.0106f
C14477 VPWR.n2675 VGND 0.02274f
C14478 VPWR.t316 VGND 0.04225f
C14479 VPWR.t277 VGND 0.04225f
C14480 VPWR.n2677 VGND 0.09744f
C14481 VPWR.t238 VGND 0.0106f
C14482 VPWR.t310 VGND 0.0106f
C14483 VPWR.n2678 VGND 0.02274f
C14484 VPWR.t227 VGND 0.0106f
C14485 VPWR.t1835 VGND 0.0106f
C14486 VPWR.n2679 VGND 0.02274f
C14487 VPWR.n2680 VGND 0.04572f
C14488 VPWR.n2681 VGND 0.01007f
C14489 VPWR.n2682 VGND 0.03127f
C14490 VPWR.n2683 VGND 0.03466f
C14491 VPWR.n2684 VGND 0.03466f
C14492 VPWR.n2685 VGND 0.01054f
C14493 VPWR.n2686 VGND 0.04572f
C14494 VPWR.n2689 VGND 0.03466f
C14495 VPWR.n2690 VGND 0.03466f
C14496 VPWR.t928 VGND 0.04034f
C14497 VPWR.t645 VGND 0.04034f
C14498 VPWR.n2693 VGND 0.07319f
C14499 VPWR.n2695 VGND 0.02599f
C14500 VPWR.n2696 VGND 0.01319f
C14501 VPWR.n2697 VGND 0.02599f
C14502 VPWR.t136 VGND 0.04226f
C14503 VPWR.n2698 VGND 0.05889f
C14504 VPWR.n2700 VGND 0.04309f
C14505 VPWR.t1234 VGND 0.04154f
C14506 VPWR.n2701 VGND 0.05384f
C14507 VPWR.n2702 VGND 0.02053f
C14508 VPWR.n2703 VGND 1.21026f
C14509 VPWR.n2704 VGND 0.03466f
C14510 VPWR.t272 VGND 0.0718f
C14511 VPWR.t223 VGND 0.10581f
C14512 VPWR.t1833 VGND 0.10287f
C14513 VPWR.t322 VGND 0.16452f
C14514 VPWR.t1088 VGND 0.13993f
C14515 VPWR.t248 VGND 0.09329f
C14516 VPWR.t1082 VGND 0.09329f
C14517 VPWR.t302 VGND 0.09329f
C14518 VPWR.t1090 VGND 0.09329f
C14519 VPWR.t243 VGND 0.09329f
C14520 VPWR.t1084 VGND 0.09329f
C14521 VPWR.t311 VGND 0.12993f
C14522 VPWR.t1235 VGND 0.0733f
C14523 VPWR.t189 VGND 0.07996f
C14524 VPWR.t133 VGND 0.09329f
C14525 VPWR.t191 VGND 0.17324f
C14526 VPWR.n2705 VGND 0.27927f
C14527 VPWR.n2706 VGND 0.12882f
C14528 VPWR.t192 VGND 0.04194f
C14529 VPWR.n2707 VGND 0.03466f
C14530 VPWR.t312 VGND 0.04146f
C14531 VPWR.t1085 VGND 0.03991f
C14532 VPWR.t303 VGND 0.0106f
C14533 VPWR.t244 VGND 0.0106f
C14534 VPWR.n2708 VGND 0.02274f
C14535 VPWR.t1083 VGND 0.0106f
C14536 VPWR.t1091 VGND 0.0106f
C14537 VPWR.n2709 VGND 0.02274f
C14538 VPWR.n2710 VGND 0.02593f
C14539 VPWR.n2711 VGND 0.03466f
C14540 VPWR.t323 VGND 0.0106f
C14541 VPWR.t1089 VGND 0.0106f
C14542 VPWR.n2712 VGND 0.02274f
C14543 VPWR.t273 VGND 0.04225f
C14544 VPWR.n2714 VGND 0.05325f
C14545 VPWR.t224 VGND 0.0106f
C14546 VPWR.t1834 VGND 0.0106f
C14547 VPWR.n2715 VGND 0.02274f
C14548 VPWR.n2716 VGND 0.02593f
C14549 VPWR.n2717 VGND 0.01007f
C14550 VPWR.n2718 VGND 0.03127f
C14551 VPWR.n2719 VGND 0.03466f
C14552 VPWR.n2720 VGND 0.03466f
C14553 VPWR.n2721 VGND 0.01054f
C14554 VPWR.n2722 VGND 0.02533f
C14555 VPWR.t249 VGND 0.03708f
C14556 VPWR.n2723 VGND 0.02956f
C14557 VPWR.n2725 VGND 0.03466f
C14558 VPWR.n2726 VGND 0.03466f
C14559 VPWR.n2727 VGND 0.02873f
C14560 VPWR.n2729 VGND 0.03803f
C14561 VPWR.n2730 VGND 0.0501f
C14562 VPWR.n2732 VGND 0.02053f
C14563 VPWR.n2733 VGND 0.01319f
C14564 VPWR.n2734 VGND 0.02599f
C14565 VPWR.t134 VGND 0.0423f
C14566 VPWR.n2735 VGND 0.10875f
C14567 VPWR.t190 VGND 0.04223f
C14568 VPWR.n2737 VGND 0.04701f
C14569 VPWR.n2738 VGND 0.02034f
C14570 VPWR.n2739 VGND 1.21026f
C14571 VPWR.n2740 VGND 0.03127f
C14572 VPWR.t279 VGND 0.49308f
C14573 VPWR.t228 VGND 0.18657f
C14574 VPWR.t321 VGND 0.18657f
C14575 VPWR.t222 VGND 0.18657f
C14576 VPWR.t124 VGND 0.18657f
C14577 VPWR.t118 VGND 0.18657f
C14578 VPWR.t126 VGND 0.18657f
C14579 VPWR.t128 VGND 0.1688f
C14580 VPWR.t43 VGND 0.40868f
C14581 VPWR.t1098 VGND 0.11327f
C14582 VPWR.n2741 VGND 0.24485f
C14583 VPWR.n2742 VGND 0.13062f
C14584 VPWR.t125 VGND 0.0106f
C14585 VPWR.t119 VGND 0.0106f
C14586 VPWR.n2743 VGND 0.02322f
C14587 VPWR.t991 VGND 0.0106f
C14588 VPWR.t990 VGND 0.0106f
C14589 VPWR.n2744 VGND 0.02322f
C14590 VPWR.n2745 VGND 0.08815f
C14591 VPWR.n2746 VGND 0.07146f
C14592 VPWR.t127 VGND 0.0106f
C14593 VPWR.t129 VGND 0.0106f
C14594 VPWR.n2747 VGND 0.02326f
C14595 VPWR.t993 VGND 0.0106f
C14596 VPWR.t987 VGND 0.0106f
C14597 VPWR.n2748 VGND 0.02326f
C14598 VPWR.n2749 VGND 0.09662f
C14599 VPWR.n2751 VGND 0.27909f
C14600 VPWR.n2752 VGND 0.01319f
C14601 VPWR.n2753 VGND 0.01206f
C14602 VPWR.n2754 VGND 0.01034f
C14603 VPWR.t44 VGND 0.0423f
C14604 VPWR.t836 VGND 0.0423f
C14605 VPWR.n2756 VGND 0.12493f
C14606 VPWR.n2757 VGND 0.02599f
C14607 VPWR.n2758 VGND 1.21026f
C14608 VPWR.n2759 VGND 0.03127f
C14609 VPWR.t237 VGND 0.49308f
C14610 VPWR.t1832 VGND 0.18657f
C14611 VPWR.t301 VGND 0.18657f
C14612 VPWR.t1831 VGND 0.18657f
C14613 VPWR.t465 VGND 0.18657f
C14614 VPWR.t475 VGND 0.18657f
C14615 VPWR.t467 VGND 0.18657f
C14616 VPWR.t469 VGND 0.1688f
C14617 VPWR.t833 VGND 0.36315f
C14618 VPWR.t1100 VGND 0.07996f
C14619 VPWR.t1104 VGND 0.07885f
C14620 VPWR.n2760 VGND 0.24374f
C14621 VPWR.n2761 VGND 0.13062f
C14622 VPWR.t466 VGND 0.0106f
C14623 VPWR.t476 VGND 0.0106f
C14624 VPWR.n2762 VGND 0.02322f
C14625 VPWR.t749 VGND 0.0106f
C14626 VPWR.t755 VGND 0.0106f
C14627 VPWR.n2763 VGND 0.02322f
C14628 VPWR.n2764 VGND 0.08815f
C14629 VPWR.n2765 VGND 0.07146f
C14630 VPWR.t468 VGND 0.0106f
C14631 VPWR.t470 VGND 0.0106f
C14632 VPWR.n2766 VGND 0.02326f
C14633 VPWR.t751 VGND 0.0106f
C14634 VPWR.t753 VGND 0.0106f
C14635 VPWR.n2767 VGND 0.02326f
C14636 VPWR.n2768 VGND 0.09662f
C14637 VPWR.n2770 VGND 0.27909f
C14638 VPWR.n2771 VGND 0.01319f
C14639 VPWR.n2772 VGND 0.01187f
C14640 VPWR.t1101 VGND 0.04221f
C14641 VPWR.n2774 VGND 0.04512f
C14642 VPWR.t834 VGND 0.0423f
C14643 VPWR.n2776 VGND 0.06737f
C14644 VPWR.n2777 VGND 0.02599f
C14645 VPWR.n2778 VGND 1.21026f
C14646 VPWR.n2779 VGND 0.03164f
C14647 VPWR.t225 VGND 0.49308f
C14648 VPWR.t250 VGND 0.18657f
C14649 VPWR.t278 VGND 0.18657f
C14650 VPWR.t241 VGND 0.18657f
C14651 VPWR.t652 VGND 0.18657f
C14652 VPWR.t646 VGND 0.18657f
C14653 VPWR.t638 VGND 0.18657f
C14654 VPWR.t640 VGND 0.1688f
C14655 VPWR.t45 VGND 0.38647f
C14656 VPWR.t1096 VGND 0.13327f
C14657 VPWR.n2780 VGND 0.24262f
C14658 VPWR.n2781 VGND 0.12868f
C14659 VPWR.t1099 VGND 0.04227f
C14660 VPWR.t932 VGND 0.0106f
C14661 VPWR.t929 VGND 0.0106f
C14662 VPWR.n2782 VGND 0.02322f
C14663 VPWR.t653 VGND 0.0106f
C14664 VPWR.t647 VGND 0.0106f
C14665 VPWR.n2783 VGND 0.02322f
C14666 VPWR.n2784 VGND 0.08815f
C14667 VPWR.n2785 VGND 0.07146f
C14668 VPWR.t925 VGND 0.0106f
C14669 VPWR.t926 VGND 0.0106f
C14670 VPWR.n2786 VGND 0.02326f
C14671 VPWR.t639 VGND 0.0106f
C14672 VPWR.t641 VGND 0.0106f
C14673 VPWR.n2787 VGND 0.02326f
C14674 VPWR.n2788 VGND 0.09662f
C14675 VPWR.n2790 VGND 0.27909f
C14676 VPWR.n2791 VGND 0.01319f
C14677 VPWR.n2792 VGND 0.01168f
C14678 VPWR.t1097 VGND 0.04227f
C14679 VPWR.n2793 VGND 0.11136f
C14680 VPWR.t46 VGND 0.04226f
C14681 VPWR.t835 VGND 0.04226f
C14682 VPWR.n2795 VGND 0.09943f
C14683 VPWR.n2796 VGND 0.02599f
C14684 VPWR.n2797 VGND 1.21026f
C14685 VPWR.n2798 VGND 0.03164f
C14686 VPWR.t832 VGND 0.04226f
C14687 VPWR.n2799 VGND 0.01168f
C14688 VPWR.t1103 VGND 0.04227f
C14689 VPWR.n2800 VGND 0.01319f
C14690 VPWR.t247 VGND 0.27964f
C14691 VPWR.t313 VGND 0.10581f
C14692 VPWR.t326 VGND 0.10581f
C14693 VPWR.t213 VGND 0.10581f
C14694 VPWR.t1086 VGND 0.10581f
C14695 VPWR.t1080 VGND 0.10581f
C14696 VPWR.t1092 VGND 0.10581f
C14697 VPWR.t1094 VGND 0.09573f
C14698 VPWR.t831 VGND 0.21918f
C14699 VPWR.t1102 VGND 0.07558f
C14700 VPWR.n2801 VGND 0.13503f
C14701 VPWR.t1093 VGND 0.0106f
C14702 VPWR.t1095 VGND 0.0106f
C14703 VPWR.n2802 VGND 0.02326f
C14704 VPWR.n2803 VGND 0.05725f
C14705 VPWR.t1087 VGND 0.0106f
C14706 VPWR.t1081 VGND 0.0106f
C14707 VPWR.n2804 VGND 0.02421f
C14708 VPWR.n2805 VGND 0.12927f
C14709 VPWR.n2806 VGND 0.27909f
C14710 VPWR.n2808 VGND 0.07145f
C14711 VPWR.n2809 VGND 0.06272f
C14712 VPWR.n2811 VGND 0.05435f
C14713 VPWR.n2812 VGND 0.02599f
C14714 VPWR.n2813 VGND 1.76121f
C14715 VPWR.n2814 VGND 1.42636f
C14716 VPWR.t194 VGND 0.02149f
C14717 VPWR.n2815 VGND 0.09631f
C14718 VPWR.n2816 VGND 0.21199f
C14719 VPWR.n2817 VGND 0.0559f
C14720 VPWR.n2818 VGND 0.02655f
C14721 VPWR.n2819 VGND 0.03242f
C14722 VPWR.n2820 VGND 0.06571f
C14723 VPWR.n2821 VGND 0.08566f
C14724 VPWR.n2822 VGND 0.06571f
C14725 VPWR.t668 VGND 2.0669f
C14726 VPWR.t193 VGND 0.65281f
C14727 VPWR.n2823 VGND 0.08633f
C14728 VPWR.n2824 VGND 0.34157f
C14729 VPWR.t669 VGND 0.02148f
C14730 VPWR.n2825 VGND 0.1315f
C14731 VPWR.n2826 VGND 0.01328f
C14732 VPWR.n2827 VGND 0.07245f
C14733 VPWR.n2828 VGND 0.06504f
C14734 VPWR.n2829 VGND 0.08633f
C14735 VPWR.n2830 VGND 0.05437f
C14736 VPWR.t1071 VGND 0.02148f
C14737 VPWR.n2831 VGND 0.1315f
C14738 VPWR.n2832 VGND 0.01328f
C14739 VPWR.n2833 VGND 0.08633f
C14740 VPWR.n2834 VGND 0.0565f
C14741 VPWR.n2835 VGND 0.06443f
C14742 VPWR.n2836 VGND 1.23519f
C14743 VPWR.n2837 VGND 0.06443f
C14744 VPWR.n2838 VGND 0.0565f
C14745 VPWR.n2839 VGND 0.08633f
C14746 VPWR.n2840 VGND 0.07238f
C14747 VPWR.n2841 VGND 0.05987f
C14748 VPWR.n2842 VGND 0.74248f
C14749 VPWR.n2843 VGND 0.04672f
C14750 VPWR.n2844 VGND 0.06535f
C14751 VPWR.n2845 VGND 0.04543f
C14752 VPWR.n2846 VGND 0.01328f
C14753 VPWR.n2847 VGND 0.04672f
C14754 VPWR.n2848 VGND 0.03587f
C14755 VPWR.n2849 VGND 0.12835f
C14756 VPWR.n2850 VGND 0.05056f
C14757 VPWR.n2851 VGND 0.03242f
C14758 VPWR.t693 VGND 0.25559f
C14759 VPWR.n2852 VGND 0.05987f
C14760 VPWR.n2853 VGND 0.07238f
C14761 VPWR.n2854 VGND 0.02655f
C14762 VPWR.n2855 VGND 1.49593f
C14763 VPWR.n2856 VGND 0.02655f
C14764 VPWR.n2857 VGND 0.02655f
C14765 VPWR.n2858 VGND 0.06598f
C14766 VPWR.n2859 VGND 0.03622f
C14767 VPWR.n2860 VGND 0.28054f
C14768 VPWR.n2861 VGND 0.23083f
C14769 VPWR.t694 VGND 0.02147f
C14770 VPWR.n2862 VGND 0.16245f
C14771 VPWR.n2863 VGND 2.5721f
C14772 XThR.Tn[2].t11 VGND 0.01796f
C14773 XThR.Tn[2].t5 VGND 0.01796f
C14774 XThR.Tn[2].n0 VGND 0.03626f
C14775 XThR.Tn[2].t4 VGND 0.01796f
C14776 XThR.Tn[2].t2 VGND 0.01796f
C14777 XThR.Tn[2].n1 VGND 0.04242f
C14778 XThR.Tn[2].n2 VGND 0.12726f
C14779 XThR.Tn[2].t3 VGND 0.01168f
C14780 XThR.Tn[2].t6 VGND 0.01168f
C14781 XThR.Tn[2].n3 VGND 0.02659f
C14782 XThR.Tn[2].t9 VGND 0.01168f
C14783 XThR.Tn[2].t10 VGND 0.01168f
C14784 XThR.Tn[2].n4 VGND 0.0443f
C14785 XThR.Tn[2].t8 VGND 0.01168f
C14786 XThR.Tn[2].t7 VGND 0.01168f
C14787 XThR.Tn[2].n5 VGND 0.02659f
C14788 XThR.Tn[2].n6 VGND 0.12662f
C14789 XThR.Tn[2].t1 VGND 0.01168f
C14790 XThR.Tn[2].t0 VGND 0.01168f
C14791 XThR.Tn[2].n7 VGND 0.02659f
C14792 XThR.Tn[2].n8 VGND 0.07828f
C14793 XThR.Tn[2].n9 VGND 0.08834f
C14794 XThR.Tn[2].t21 VGND 0.01404f
C14795 XThR.Tn[2].t14 VGND 0.01537f
C14796 XThR.Tn[2].n10 VGND 0.03754f
C14797 XThR.Tn[2].n11 VGND 0.07211f
C14798 XThR.Tn[2].t40 VGND 0.01404f
C14799 XThR.Tn[2].t31 VGND 0.01537f
C14800 XThR.Tn[2].n12 VGND 0.03754f
C14801 XThR.Tn[2].t55 VGND 0.01399f
C14802 XThR.Tn[2].t66 VGND 0.01532f
C14803 XThR.Tn[2].n13 VGND 0.03906f
C14804 XThR.Tn[2].n14 VGND 0.02744f
C14805 XThR.Tn[2].n16 VGND 0.08806f
C14806 XThR.Tn[2].t15 VGND 0.01404f
C14807 XThR.Tn[2].t67 VGND 0.01537f
C14808 XThR.Tn[2].n17 VGND 0.03754f
C14809 XThR.Tn[2].t30 VGND 0.01399f
C14810 XThR.Tn[2].t43 VGND 0.01532f
C14811 XThR.Tn[2].n18 VGND 0.03906f
C14812 XThR.Tn[2].n19 VGND 0.02744f
C14813 XThR.Tn[2].n21 VGND 0.08806f
C14814 XThR.Tn[2].t32 VGND 0.01404f
C14815 XThR.Tn[2].t23 VGND 0.01537f
C14816 XThR.Tn[2].n22 VGND 0.03754f
C14817 XThR.Tn[2].t47 VGND 0.01399f
C14818 XThR.Tn[2].t60 VGND 0.01532f
C14819 XThR.Tn[2].n23 VGND 0.03906f
C14820 XThR.Tn[2].n24 VGND 0.02744f
C14821 XThR.Tn[2].n26 VGND 0.08806f
C14822 XThR.Tn[2].t58 VGND 0.01404f
C14823 XThR.Tn[2].t50 VGND 0.01537f
C14824 XThR.Tn[2].n27 VGND 0.03754f
C14825 XThR.Tn[2].t16 VGND 0.01399f
C14826 XThR.Tn[2].t28 VGND 0.01532f
C14827 XThR.Tn[2].n28 VGND 0.03906f
C14828 XThR.Tn[2].n29 VGND 0.02744f
C14829 XThR.Tn[2].n31 VGND 0.08806f
C14830 XThR.Tn[2].t34 VGND 0.01404f
C14831 XThR.Tn[2].t25 VGND 0.01537f
C14832 XThR.Tn[2].n32 VGND 0.03754f
C14833 XThR.Tn[2].t48 VGND 0.01399f
C14834 XThR.Tn[2].t62 VGND 0.01532f
C14835 XThR.Tn[2].n33 VGND 0.03906f
C14836 XThR.Tn[2].n34 VGND 0.02744f
C14837 XThR.Tn[2].n36 VGND 0.08806f
C14838 XThR.Tn[2].t70 VGND 0.01404f
C14839 XThR.Tn[2].t41 VGND 0.01537f
C14840 XThR.Tn[2].n37 VGND 0.03754f
C14841 XThR.Tn[2].t22 VGND 0.01399f
C14842 XThR.Tn[2].t20 VGND 0.01532f
C14843 XThR.Tn[2].n38 VGND 0.03906f
C14844 XThR.Tn[2].n39 VGND 0.02744f
C14845 XThR.Tn[2].n41 VGND 0.08806f
C14846 XThR.Tn[2].t39 VGND 0.01404f
C14847 XThR.Tn[2].t35 VGND 0.01537f
C14848 XThR.Tn[2].n42 VGND 0.03754f
C14849 XThR.Tn[2].t54 VGND 0.01399f
C14850 XThR.Tn[2].t12 VGND 0.01532f
C14851 XThR.Tn[2].n43 VGND 0.03906f
C14852 XThR.Tn[2].n44 VGND 0.02744f
C14853 XThR.Tn[2].n46 VGND 0.08806f
C14854 XThR.Tn[2].t44 VGND 0.01404f
C14855 XThR.Tn[2].t49 VGND 0.01537f
C14856 XThR.Tn[2].n47 VGND 0.03754f
C14857 XThR.Tn[2].t57 VGND 0.01399f
C14858 XThR.Tn[2].t27 VGND 0.01532f
C14859 XThR.Tn[2].n48 VGND 0.03906f
C14860 XThR.Tn[2].n49 VGND 0.02744f
C14861 XThR.Tn[2].n51 VGND 0.08806f
C14862 XThR.Tn[2].t61 VGND 0.01404f
C14863 XThR.Tn[2].t69 VGND 0.01537f
C14864 XThR.Tn[2].n52 VGND 0.03754f
C14865 XThR.Tn[2].t18 VGND 0.01399f
C14866 XThR.Tn[2].t45 VGND 0.01532f
C14867 XThR.Tn[2].n53 VGND 0.03906f
C14868 XThR.Tn[2].n54 VGND 0.02744f
C14869 XThR.Tn[2].n56 VGND 0.08806f
C14870 XThR.Tn[2].t52 VGND 0.01404f
C14871 XThR.Tn[2].t26 VGND 0.01537f
C14872 XThR.Tn[2].n57 VGND 0.03754f
C14873 XThR.Tn[2].t68 VGND 0.01399f
C14874 XThR.Tn[2].t63 VGND 0.01532f
C14875 XThR.Tn[2].n58 VGND 0.03906f
C14876 XThR.Tn[2].n59 VGND 0.02744f
C14877 XThR.Tn[2].n61 VGND 0.08806f
C14878 XThR.Tn[2].t73 VGND 0.01404f
C14879 XThR.Tn[2].t64 VGND 0.01537f
C14880 XThR.Tn[2].n62 VGND 0.03754f
C14881 XThR.Tn[2].t24 VGND 0.01399f
C14882 XThR.Tn[2].t37 VGND 0.01532f
C14883 XThR.Tn[2].n63 VGND 0.03906f
C14884 XThR.Tn[2].n64 VGND 0.02744f
C14885 XThR.Tn[2].n66 VGND 0.08806f
C14886 XThR.Tn[2].t42 VGND 0.01404f
C14887 XThR.Tn[2].t36 VGND 0.01537f
C14888 XThR.Tn[2].n67 VGND 0.03754f
C14889 XThR.Tn[2].t56 VGND 0.01399f
C14890 XThR.Tn[2].t13 VGND 0.01532f
C14891 XThR.Tn[2].n68 VGND 0.03906f
C14892 XThR.Tn[2].n69 VGND 0.02744f
C14893 XThR.Tn[2].n71 VGND 0.08806f
C14894 XThR.Tn[2].t59 VGND 0.01404f
C14895 XThR.Tn[2].t51 VGND 0.01537f
C14896 XThR.Tn[2].n72 VGND 0.03754f
C14897 XThR.Tn[2].t17 VGND 0.01399f
C14898 XThR.Tn[2].t29 VGND 0.01532f
C14899 XThR.Tn[2].n73 VGND 0.03906f
C14900 XThR.Tn[2].n74 VGND 0.02744f
C14901 XThR.Tn[2].n76 VGND 0.08806f
C14902 XThR.Tn[2].t19 VGND 0.01404f
C14903 XThR.Tn[2].t72 VGND 0.01537f
C14904 XThR.Tn[2].n77 VGND 0.03754f
C14905 XThR.Tn[2].t33 VGND 0.01399f
C14906 XThR.Tn[2].t46 VGND 0.01532f
C14907 XThR.Tn[2].n78 VGND 0.03906f
C14908 XThR.Tn[2].n79 VGND 0.02744f
C14909 XThR.Tn[2].n81 VGND 0.08806f
C14910 XThR.Tn[2].t53 VGND 0.01404f
C14911 XThR.Tn[2].t65 VGND 0.01537f
C14912 XThR.Tn[2].n82 VGND 0.03754f
C14913 XThR.Tn[2].t71 VGND 0.01399f
C14914 XThR.Tn[2].t38 VGND 0.01532f
C14915 XThR.Tn[2].n83 VGND 0.03906f
C14916 XThR.Tn[2].n84 VGND 0.02744f
C14917 XThR.Tn[2].n86 VGND 0.08806f
C14918 XThR.Tn[2].n87 VGND 0.08002f
C14919 XThR.Tn[2].n88 VGND 0.17341f
.ends

