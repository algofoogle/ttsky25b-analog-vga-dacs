magic
tech sky130A
magscale 1 2
timestamp 1762784779
<< metal1 >>
rect 10136 38319 10216 38324
rect 6305 38314 10216 38319
rect 6305 38256 10148 38314
rect 10206 38256 10216 38314
rect 6305 38249 10216 38256
rect 6320 37812 6360 38249
rect 10136 38244 10216 38249
rect 6910 38170 10216 38180
rect 6910 38112 10148 38170
rect 10206 38112 10216 38170
rect 6910 38100 10216 38112
rect 6930 37808 6970 38100
rect 10136 38029 10216 38038
rect 8486 38028 10216 38029
rect 8486 37970 10148 38028
rect 10206 37970 10216 38028
rect 8486 37968 10216 37970
rect 8496 37812 8536 37968
rect 10136 37958 10216 37968
rect 10136 37889 10216 37898
rect 8568 37888 10216 37889
rect 8568 37830 10148 37888
rect 10206 37830 10216 37888
rect 8568 37828 10216 37830
rect 8578 37812 8618 37828
rect 10136 37818 10216 37828
rect 18204 30729 18284 30734
rect 18194 30724 18284 30729
rect 18194 30666 18216 30724
rect 18274 30666 18284 30724
rect 18194 30659 18284 30666
rect 18204 30654 18284 30659
rect 18194 30580 18284 30590
rect 18194 30522 18216 30580
rect 18274 30522 18284 30580
rect 18194 30510 18284 30522
rect 18204 29039 18284 29048
rect 18194 29038 18284 29039
rect 18194 28980 18216 29038
rect 18274 28980 18284 29038
rect 18194 28978 18284 28980
rect 18204 28968 18284 28978
rect 18204 28487 18284 28496
rect 18194 28486 18284 28487
rect 18194 28428 18216 28486
rect 18274 28428 18284 28486
rect 18194 28426 18284 28428
rect 18204 28416 18284 28426
rect 10136 25605 10216 25610
rect 6305 25600 10216 25605
rect 6305 25542 10148 25600
rect 10206 25542 10216 25600
rect 6305 25535 10216 25542
rect 6320 25098 6360 25535
rect 10136 25530 10216 25535
rect 6910 25456 10216 25466
rect 6910 25398 10148 25456
rect 10206 25398 10216 25456
rect 6910 25386 10216 25398
rect 6930 25094 6970 25386
rect 10136 25315 10216 25324
rect 8486 25314 10216 25315
rect 8486 25256 10148 25314
rect 10206 25256 10216 25314
rect 8486 25254 10216 25256
rect 8496 25098 8536 25254
rect 10136 25244 10216 25254
rect 10136 25175 10216 25184
rect 8568 25174 10216 25175
rect 8568 25116 10148 25174
rect 10206 25116 10216 25174
rect 8568 25114 10216 25116
rect 8578 25098 8618 25114
rect 10136 25104 10216 25114
rect 18204 18015 18284 18020
rect 18194 18010 18284 18015
rect 18194 17952 18216 18010
rect 18274 17952 18284 18010
rect 18194 17945 18284 17952
rect 18204 17940 18284 17945
rect 18194 17866 18284 17876
rect 18194 17808 18216 17866
rect 18274 17808 18284 17866
rect 18194 17796 18284 17808
rect 18204 16325 18284 16334
rect 18194 16324 18284 16325
rect 18194 16266 18216 16324
rect 18274 16266 18284 16324
rect 18194 16264 18284 16266
rect 18204 16254 18284 16264
rect 18204 15773 18284 15782
rect 18194 15772 18284 15773
rect 18194 15714 18216 15772
rect 18274 15714 18284 15772
rect 18194 15712 18284 15714
rect 18204 15702 18284 15712
rect 10136 12891 10216 12896
rect 6305 12886 10216 12891
rect 6305 12828 10148 12886
rect 10206 12828 10216 12886
rect 6305 12821 10216 12828
rect 6320 12384 6360 12821
rect 10136 12816 10216 12821
rect 6910 12742 10216 12752
rect 6910 12684 10148 12742
rect 10206 12684 10216 12742
rect 6910 12672 10216 12684
rect 6930 12380 6970 12672
rect 10136 12601 10216 12610
rect 8486 12600 10216 12601
rect 8486 12542 10148 12600
rect 10206 12542 10216 12600
rect 8486 12540 10216 12542
rect 8496 12384 8536 12540
rect 10136 12530 10216 12540
rect 10136 12461 10216 12470
rect 8568 12460 10216 12461
rect 8568 12402 10148 12460
rect 10206 12402 10216 12460
rect 8568 12400 10216 12402
rect 8578 12384 8618 12400
rect 10136 12390 10216 12400
rect 18204 5301 18284 5306
rect 18194 5296 18284 5301
rect 18194 5238 18216 5296
rect 18274 5238 18284 5296
rect 18194 5231 18284 5238
rect 18204 5226 18284 5231
rect 18194 5152 18284 5162
rect 18194 5094 18216 5152
rect 18274 5094 18284 5152
rect 18194 5082 18284 5094
rect 18204 3611 18284 3620
rect 18194 3610 18284 3611
rect 18194 3552 18216 3610
rect 18274 3552 18284 3610
rect 18194 3550 18284 3552
rect 18204 3540 18284 3550
rect 18204 3059 18284 3068
rect 18194 3058 18284 3059
rect 18194 3000 18216 3058
rect 18274 3000 18284 3058
rect 18194 2998 18284 3000
rect 18204 2988 18284 2998
<< via1 >>
rect 10148 38256 10206 38314
rect 10148 38112 10206 38170
rect 10148 37970 10206 38028
rect 10148 37830 10206 37888
rect 18216 30666 18274 30724
rect 18216 30522 18274 30580
rect 18216 28980 18274 29038
rect 18216 28428 18274 28486
rect 10148 25542 10206 25600
rect 10148 25398 10206 25456
rect 10148 25256 10206 25314
rect 10148 25116 10206 25174
rect 18216 17952 18274 18010
rect 18216 17808 18274 17866
rect 18216 16266 18274 16324
rect 18216 15714 18274 15772
rect 10148 12828 10206 12886
rect 10148 12684 10206 12742
rect 10148 12542 10206 12600
rect 10148 12402 10206 12460
rect 18216 5238 18274 5296
rect 18216 5094 18274 5152
rect 18216 3552 18274 3610
rect 18216 3000 18274 3058
<< metal2 >>
rect 21028 44902 21112 44912
rect 21028 44800 21038 44902
rect 21102 44800 21112 44902
rect 21028 44790 21112 44800
rect 21580 44902 21664 44912
rect 21580 44800 21590 44902
rect 21654 44800 21664 44902
rect 21580 44790 21664 44800
rect 22132 44902 22216 44912
rect 22132 44800 22142 44902
rect 22206 44800 22216 44902
rect 22132 44790 22216 44800
rect 22684 44902 22768 44912
rect 22684 44800 22694 44902
rect 22758 44800 22768 44902
rect 22684 44790 22768 44800
rect 23236 44902 23320 44912
rect 23236 44800 23246 44902
rect 23310 44800 23320 44902
rect 23236 44790 23320 44800
rect 23788 44902 23872 44912
rect 23788 44800 23798 44902
rect 23862 44800 23872 44902
rect 23788 44790 23872 44800
rect 24340 44902 24424 44912
rect 24340 44800 24350 44902
rect 24414 44800 24424 44902
rect 24340 44790 24424 44800
rect 24892 44902 24976 44912
rect 24892 44800 24902 44902
rect 24966 44800 24976 44902
rect 24892 44790 24976 44800
rect 25444 44902 25528 44912
rect 25444 44800 25454 44902
rect 25518 44800 25528 44902
rect 25444 44790 25528 44800
rect 25996 44902 26080 44912
rect 25996 44800 26006 44902
rect 26070 44800 26080 44902
rect 25996 44790 26080 44800
rect 26548 44902 26632 44912
rect 26548 44800 26558 44902
rect 26622 44800 26632 44902
rect 26548 44790 26632 44800
rect 27100 44902 27184 44912
rect 27100 44800 27110 44902
rect 27174 44800 27184 44902
rect 27100 44790 27184 44800
rect 27652 44902 27736 44912
rect 27652 44800 27662 44902
rect 27726 44800 27736 44902
rect 27652 44790 27736 44800
rect 28204 44902 28288 44912
rect 28204 44800 28214 44902
rect 28278 44800 28288 44902
rect 28204 44790 28288 44800
rect 28756 44902 28840 44912
rect 28756 44800 28766 44902
rect 28830 44800 28840 44902
rect 28756 44790 28840 44800
rect 29308 44902 29392 44912
rect 29308 44800 29318 44902
rect 29382 44800 29392 44902
rect 29308 44790 29392 44800
rect 21038 44758 21102 44790
rect 21590 44758 21654 44790
rect 22142 44758 22206 44790
rect 22694 44758 22758 44790
rect 23246 44758 23310 44790
rect 23798 44758 23862 44790
rect 24350 44758 24414 44790
rect 24902 44758 24966 44790
rect 25454 44758 25518 44790
rect 26006 44758 26070 44790
rect 26558 44758 26622 44790
rect 27110 44758 27174 44790
rect 27662 44758 27726 44790
rect 28214 44758 28278 44790
rect 28766 44758 28830 44790
rect 29318 44758 29382 44790
rect 10136 38314 10216 38324
rect 10136 38256 10148 38314
rect 10206 38256 10216 38314
rect 10136 38244 10216 38256
rect 10136 38170 10216 38180
rect 10136 38112 10148 38170
rect 10206 38112 10216 38170
rect 10136 38100 10216 38112
rect 10136 38028 10216 38038
rect 10136 37970 10148 38028
rect 10206 37970 10216 38028
rect 10136 37958 10216 37970
rect 10136 37888 10216 37898
rect 10136 37830 10148 37888
rect 10206 37830 10216 37888
rect 10136 37818 10216 37830
rect 18532 36972 18608 36982
rect 18532 36966 18542 36972
rect 18208 36920 18542 36966
rect 18532 36916 18542 36920
rect 18598 36916 18608 36972
rect 18532 36906 18608 36916
rect 18532 36698 18608 36708
rect 18532 36694 18542 36698
rect 18208 36648 18542 36694
rect 18532 36642 18542 36648
rect 18598 36642 18608 36698
rect 18532 36632 18608 36642
rect 18532 36426 18608 36436
rect 18532 36422 18542 36426
rect 18208 36376 18542 36422
rect 18532 36370 18542 36376
rect 18598 36370 18608 36426
rect 18532 36360 18608 36370
rect 18204 30724 18284 30734
rect 18204 30666 18216 30724
rect 18274 30666 18284 30724
rect 18204 30654 18284 30666
rect 18204 30580 18284 30590
rect 18204 30522 18216 30580
rect 18274 30522 18284 30580
rect 18204 30510 18284 30522
rect 18204 29038 18284 29048
rect 18204 28980 18216 29038
rect 18274 28980 18284 29038
rect 18204 28968 18284 28980
rect 18204 28486 18284 28496
rect 18204 28428 18216 28486
rect 18274 28428 18284 28486
rect 18204 28416 18284 28428
rect 10136 25600 10216 25610
rect 10136 25542 10148 25600
rect 10206 25542 10216 25600
rect 10136 25530 10216 25542
rect 10136 25456 10216 25466
rect 10136 25398 10148 25456
rect 10206 25398 10216 25456
rect 10136 25386 10216 25398
rect 10136 25314 10216 25324
rect 10136 25256 10148 25314
rect 10206 25256 10216 25314
rect 10136 25244 10216 25256
rect 10136 25174 10216 25184
rect 10136 25116 10148 25174
rect 10206 25116 10216 25174
rect 10136 25104 10216 25116
rect 18412 24258 18488 24268
rect 18412 24252 18422 24258
rect 18208 24206 18422 24252
rect 18412 24202 18422 24206
rect 18478 24202 18488 24258
rect 18412 24192 18488 24202
rect 18412 23984 18488 23994
rect 18412 23980 18422 23984
rect 18208 23934 18422 23980
rect 18412 23928 18422 23934
rect 18478 23928 18488 23984
rect 18412 23918 18488 23928
rect 18412 23712 18488 23722
rect 18412 23708 18422 23712
rect 18208 23662 18422 23708
rect 18412 23656 18422 23662
rect 18478 23656 18488 23712
rect 18412 23646 18488 23656
rect 18204 18010 18284 18020
rect 18204 17952 18216 18010
rect 18274 17952 18284 18010
rect 18204 17940 18284 17952
rect 18204 17866 18284 17876
rect 18204 17808 18216 17866
rect 18274 17808 18284 17866
rect 18204 17796 18284 17808
rect 18204 16324 18284 16334
rect 18204 16266 18216 16324
rect 18274 16266 18284 16324
rect 18204 16254 18284 16266
rect 18204 15772 18284 15782
rect 18204 15714 18216 15772
rect 18274 15714 18284 15772
rect 18204 15702 18284 15714
rect 10136 12886 10216 12896
rect 10136 12828 10148 12886
rect 10206 12828 10216 12886
rect 10136 12816 10216 12828
rect 10136 12742 10216 12752
rect 10136 12684 10148 12742
rect 10206 12684 10216 12742
rect 10136 12672 10216 12684
rect 10136 12600 10216 12610
rect 10136 12542 10148 12600
rect 10206 12542 10216 12600
rect 10136 12530 10216 12542
rect 10136 12460 10216 12470
rect 10136 12402 10148 12460
rect 10206 12402 10216 12460
rect 10136 12390 10216 12402
rect 18412 11544 18488 11554
rect 18412 11538 18422 11544
rect 18208 11492 18422 11538
rect 18412 11488 18422 11492
rect 18478 11488 18488 11544
rect 18412 11478 18488 11488
rect 18412 11270 18488 11280
rect 18412 11266 18422 11270
rect 18208 11220 18422 11266
rect 18412 11214 18422 11220
rect 18478 11214 18488 11270
rect 18412 11204 18488 11214
rect 18412 10998 18488 11008
rect 18412 10994 18422 10998
rect 18208 10948 18422 10994
rect 18412 10942 18422 10948
rect 18478 10942 18488 10998
rect 18412 10932 18488 10942
rect 18204 5296 18284 5306
rect 18204 5238 18216 5296
rect 18274 5238 18284 5296
rect 18204 5226 18284 5238
rect 18204 5152 18284 5162
rect 18204 5094 18216 5152
rect 18274 5094 18284 5152
rect 18204 5082 18284 5094
rect 18204 3610 18284 3620
rect 18204 3552 18216 3610
rect 18274 3552 18284 3610
rect 18204 3540 18284 3552
rect 18204 3058 18284 3068
rect 18204 3000 18216 3058
rect 18274 3000 18284 3058
rect 18204 2988 18284 3000
<< via2 >>
rect 21038 44800 21102 44902
rect 21590 44800 21654 44902
rect 22142 44800 22206 44902
rect 22694 44800 22758 44902
rect 23246 44800 23310 44902
rect 23798 44800 23862 44902
rect 24350 44800 24414 44902
rect 24902 44800 24966 44902
rect 25454 44800 25518 44902
rect 26006 44800 26070 44902
rect 26558 44800 26622 44902
rect 27110 44800 27174 44902
rect 27662 44800 27726 44902
rect 28214 44800 28278 44902
rect 28766 44800 28830 44902
rect 29318 44800 29382 44902
rect 10148 38256 10206 38314
rect 10148 38112 10206 38170
rect 10148 37970 10206 38028
rect 10148 37830 10206 37888
rect 18542 36916 18598 36972
rect 18542 36642 18598 36698
rect 18542 36370 18598 36426
rect 18216 30666 18274 30724
rect 18216 30522 18274 30580
rect 18216 28980 18274 29038
rect 18216 28428 18274 28486
rect 10148 25542 10206 25600
rect 10148 25398 10206 25456
rect 10148 25256 10206 25314
rect 10148 25116 10206 25174
rect 18422 24202 18478 24258
rect 18422 23928 18478 23984
rect 18422 23656 18478 23712
rect 18216 17952 18274 18010
rect 18216 17808 18274 17866
rect 18216 16266 18274 16324
rect 18216 15714 18274 15772
rect 10148 12828 10206 12886
rect 10148 12684 10206 12742
rect 10148 12542 10206 12600
rect 10148 12402 10206 12460
rect 18422 11488 18478 11544
rect 18422 11214 18478 11270
rect 18422 10942 18478 10998
rect 18216 5238 18274 5296
rect 18216 5094 18274 5152
rect 18216 3552 18274 3610
rect 18216 3000 18274 3058
<< metal3 >>
rect 9722 44846 9728 44910
rect 9792 44846 9798 44910
rect 21028 44906 21112 44912
rect 9730 44642 9790 44846
rect 21028 44796 21034 44906
rect 21106 44796 21112 44906
rect 21028 44790 21112 44796
rect 21580 44906 21664 44912
rect 21580 44796 21586 44906
rect 21658 44796 21664 44906
rect 21580 44790 21664 44796
rect 22132 44906 22216 44912
rect 22132 44796 22138 44906
rect 22210 44796 22216 44906
rect 22132 44790 22216 44796
rect 22684 44906 22768 44912
rect 22684 44796 22690 44906
rect 22762 44796 22768 44906
rect 22684 44790 22768 44796
rect 23236 44906 23320 44912
rect 23236 44796 23242 44906
rect 23314 44796 23320 44906
rect 23236 44790 23320 44796
rect 23788 44906 23872 44912
rect 23788 44796 23794 44906
rect 23866 44796 23872 44906
rect 23788 44790 23872 44796
rect 24340 44906 24424 44912
rect 24340 44796 24346 44906
rect 24418 44796 24424 44906
rect 24340 44790 24424 44796
rect 24892 44906 24976 44912
rect 24892 44796 24898 44906
rect 24970 44796 24976 44906
rect 24892 44790 24976 44796
rect 25444 44906 25528 44912
rect 25444 44796 25450 44906
rect 25522 44796 25528 44906
rect 25444 44790 25528 44796
rect 25996 44906 26080 44912
rect 25996 44796 26002 44906
rect 26074 44796 26080 44906
rect 25996 44790 26080 44796
rect 26548 44906 26632 44912
rect 26548 44796 26554 44906
rect 26626 44796 26632 44906
rect 26548 44790 26632 44796
rect 27100 44906 27184 44912
rect 27100 44796 27106 44906
rect 27178 44796 27184 44906
rect 27100 44790 27184 44796
rect 27652 44906 27736 44912
rect 27652 44796 27658 44906
rect 27730 44796 27736 44906
rect 27652 44790 27736 44796
rect 28204 44906 28288 44912
rect 28204 44796 28210 44906
rect 28282 44796 28288 44906
rect 28204 44790 28288 44796
rect 28756 44906 28840 44912
rect 28756 44796 28762 44906
rect 28834 44796 28840 44906
rect 28756 44790 28840 44796
rect 29308 44906 29392 44912
rect 29308 44796 29314 44906
rect 29386 44796 29392 44906
rect 29308 44790 29392 44796
rect 540 44582 9790 44642
rect 540 44044 616 44582
rect 540 43980 546 44044
rect 610 43980 616 44044
rect 909 43840 915 44210
rect 1283 44190 30425 44210
rect 1283 43930 23690 44190
rect 24000 43930 30090 44190
rect 30400 43930 30425 44190
rect 1283 43840 30425 43930
rect 159 43290 165 43660
rect 533 43290 19530 43660
rect 23010 43290 23360 43370
rect 29410 43290 29770 43380
rect 19130 43280 29770 43290
rect 19130 42980 23030 43280
rect 23340 42980 29430 43280
rect 29740 42980 29770 43280
rect 19130 42970 29770 42980
rect 13798 42640 19490 42644
rect 13798 42528 18794 42640
rect 18926 42528 19490 42640
rect 13798 42524 19490 42528
rect 13798 42368 19490 42372
rect 13798 42256 18242 42368
rect 18374 42256 19490 42368
rect 13798 42252 19490 42256
rect 13798 42096 19490 42100
rect 13798 41984 17690 42096
rect 17822 41984 19490 42096
rect 13798 41980 19490 41984
rect 13798 41824 19490 41828
rect 13798 41712 17138 41824
rect 17270 41712 19490 41824
rect 13798 41708 19490 41712
rect 13798 41552 19490 41556
rect 13798 41440 16586 41552
rect 16718 41440 19490 41552
rect 13798 41436 19490 41440
rect 13798 41280 19490 41284
rect 13798 41168 16034 41280
rect 16166 41168 19490 41280
rect 13798 41164 19490 41168
rect 13798 41008 19490 41012
rect 13798 40896 15482 41008
rect 15614 40896 19490 41008
rect 13798 40892 19490 40896
rect 13798 40736 19490 40740
rect 13798 40624 14930 40736
rect 15062 40624 19490 40736
rect 13798 40620 19490 40624
rect 13798 40464 19490 40468
rect 13798 40352 14378 40464
rect 14510 40352 19490 40464
rect 13798 40348 19490 40352
rect 13798 40192 19490 40196
rect 13798 40080 13826 40192
rect 13958 40080 19490 40192
rect 13798 40076 19490 40080
rect 10136 38316 10216 38324
rect 10136 38314 19131 38316
rect 10136 38256 10148 38314
rect 10206 38256 19131 38314
rect 10136 38254 19131 38256
rect 10136 38244 10216 38254
rect 10136 38172 10216 38180
rect 10136 38170 18959 38172
rect 10136 38112 10148 38170
rect 10206 38112 18959 38170
rect 10136 38110 18959 38112
rect 10136 38100 10216 38110
rect 10136 38030 10216 38038
rect 10136 38028 18789 38030
rect 10136 37970 10148 38028
rect 10206 37970 18789 38028
rect 10136 37968 18789 37970
rect 10136 37958 10216 37968
rect 10136 37890 10216 37898
rect 10136 37888 18536 37890
rect 10136 37830 10148 37888
rect 10206 37830 18536 37888
rect 10136 37828 18536 37830
rect 10136 37818 10216 37828
rect 0 37744 1840 37754
rect 0 36940 10 37744
rect 710 36940 1840 37744
rect 18474 37179 18536 37828
rect 18727 37453 18789 37968
rect 18897 37737 18959 38110
rect 19069 37991 19131 38254
rect 19069 37929 19490 37991
rect 18897 37675 19490 37737
rect 18727 37391 19490 37453
rect 18474 37117 19490 37179
rect 18532 36980 18608 36982
rect 18532 36972 19284 36980
rect 18532 36916 18542 36972
rect 18598 36916 19284 36972
rect 18532 36908 19284 36916
rect 18532 36906 18608 36908
rect 18532 36706 18608 36708
rect 18532 36698 19104 36706
rect 18532 36642 18542 36698
rect 18598 36642 19104 36698
rect 18532 36634 19104 36642
rect 18532 36632 18608 36634
rect 18532 36434 18608 36436
rect 18532 36426 18914 36434
rect 18532 36370 18542 36426
rect 18598 36370 18914 36426
rect 18532 36362 18914 36370
rect 18532 36360 18608 36362
rect 0 34946 10 35960
rect 710 34946 1840 35960
rect 18363 35652 18541 35657
rect 17132 35472 17138 35652
rect 17316 35651 18542 35652
rect 17316 35473 18363 35651
rect 18541 35473 18542 35651
rect 17316 35472 18542 35473
rect 18363 35467 18541 35472
rect 18842 35272 18914 36362
rect 19032 35542 19104 36634
rect 19212 35812 19284 36908
rect 19212 35740 19490 35812
rect 19032 35470 19490 35542
rect 18842 35200 19490 35272
rect 0 34936 1840 34946
rect 18204 30726 18284 30734
rect 18204 30724 19030 30726
rect 18204 30666 18216 30724
rect 18274 30666 19030 30724
rect 18204 30664 19030 30666
rect 18204 30654 18284 30664
rect 18204 30582 18284 30590
rect 18204 30580 18849 30582
rect 18204 30522 18216 30580
rect 18274 30522 18849 30580
rect 18204 30520 18849 30522
rect 18204 30510 18284 30520
rect 18787 29551 18849 30520
rect 18968 29831 19030 30664
rect 18968 29769 19490 29831
rect 18787 29489 19490 29551
rect 18783 29213 19490 29275
rect 18204 29040 18284 29048
rect 18783 29040 18845 29213
rect 18204 29038 18845 29040
rect 18204 28980 18216 29038
rect 18274 28980 18845 29038
rect 18204 28978 18845 28980
rect 18204 28968 18284 28978
rect 18987 28951 19490 29013
rect 18204 28488 18284 28496
rect 18987 28488 19049 28951
rect 18204 28486 19049 28488
rect 18204 28428 18216 28486
rect 18274 28428 19049 28486
rect 18204 28426 19049 28428
rect 18204 28416 18284 28426
rect 19129 26722 19307 26727
rect 17054 26542 17060 26722
rect 17238 26721 19308 26722
rect 17238 26543 19129 26721
rect 19307 26543 19308 26721
rect 17238 26542 19308 26543
rect 19129 26537 19307 26542
rect 10136 25602 10216 25610
rect 10136 25600 19190 25602
rect 10136 25542 10148 25600
rect 10206 25542 19190 25600
rect 10136 25540 19190 25542
rect 10136 25530 10216 25540
rect 10136 25458 10216 25466
rect 10136 25456 19057 25458
rect 10136 25398 10148 25456
rect 10206 25398 19057 25456
rect 10136 25396 19057 25398
rect 10136 25386 10216 25396
rect 10136 25316 10216 25324
rect 10136 25314 18899 25316
rect 10136 25256 10148 25314
rect 10206 25256 18899 25314
rect 10136 25254 18899 25256
rect 10136 25244 10216 25254
rect 10136 25176 10216 25184
rect 10136 25174 18729 25176
rect 10136 25116 10148 25174
rect 10206 25116 18729 25174
rect 10136 25114 18729 25116
rect 10136 25104 10216 25114
rect 0 25030 1840 25040
rect 0 24120 10 25030
rect 710 24120 1840 25030
rect 18667 24461 18729 25114
rect 18837 24655 18899 25254
rect 18995 24927 19057 25396
rect 19128 25211 19190 25540
rect 19128 25149 19490 25211
rect 18995 24865 19490 24927
rect 18837 24593 19490 24655
rect 18667 24399 19207 24461
rect 19145 24387 19207 24399
rect 19145 24325 19490 24387
rect 18412 24266 18488 24268
rect 18412 24258 19016 24266
rect 18412 24202 18422 24258
rect 18478 24202 19016 24258
rect 18412 24194 19016 24202
rect 18412 24192 18488 24194
rect 18944 24120 19016 24194
rect 18944 24048 19490 24120
rect 18412 23992 18488 23994
rect 18412 23984 18870 23992
rect 18412 23928 18422 23984
rect 18478 23928 18870 23984
rect 18412 23920 18870 23928
rect 18412 23918 18488 23920
rect 18798 23850 18870 23920
rect 18798 23778 19490 23850
rect 18412 23720 18488 23722
rect 18412 23712 18740 23720
rect 18412 23656 18422 23712
rect 18478 23656 18740 23712
rect 18412 23648 18740 23656
rect 18412 23646 18488 23648
rect 18668 23582 18740 23648
rect 18668 23510 19490 23582
rect 0 22232 10 23140
rect 710 22232 1840 23140
rect 0 22222 1840 22232
rect 18721 18071 19490 18133
rect 18204 18012 18284 18020
rect 18721 18012 18783 18071
rect 18204 18010 18783 18012
rect 18204 17952 18216 18010
rect 18274 17952 18783 18010
rect 18204 17950 18783 17952
rect 18204 17940 18284 17950
rect 18204 17868 18284 17876
rect 18204 17866 19490 17868
rect 18204 17808 18216 17866
rect 18274 17808 19490 17866
rect 18204 17806 19490 17808
rect 18204 17796 18284 17806
rect 18811 17519 19490 17581
rect 18204 16326 18284 16334
rect 18811 16326 18873 17519
rect 18204 16324 18873 16326
rect 18204 16266 18216 16324
rect 18274 16266 18873 16324
rect 18204 16264 18873 16266
rect 19069 17259 19490 17321
rect 18204 16254 18284 16264
rect 18204 15774 18284 15782
rect 19069 15774 19131 17259
rect 18204 15772 19131 15774
rect 18204 15714 18216 15772
rect 18274 15714 19131 15772
rect 18204 15712 19131 15714
rect 18204 15702 18284 15712
rect 18760 13998 18960 14010
rect 17320 13818 17326 13998
rect 17504 13997 18960 13998
rect 17504 13819 18777 13997
rect 18955 13819 18960 13997
rect 17504 13818 18960 13819
rect 18760 13810 18960 13818
rect 17814 13447 19490 13509
rect 10136 12888 10216 12896
rect 17814 12888 17876 13447
rect 10136 12886 17876 12888
rect 10136 12828 10148 12886
rect 10206 12828 17876 12886
rect 10136 12826 17876 12828
rect 17957 13175 19490 13237
rect 10136 12816 10216 12826
rect 10136 12744 10216 12752
rect 17957 12744 18019 13175
rect 10136 12742 18019 12744
rect 10136 12684 10148 12742
rect 10206 12684 18019 12742
rect 10136 12682 18019 12684
rect 18117 12905 19490 12967
rect 10136 12672 10216 12682
rect 10136 12602 10216 12610
rect 18117 12602 18179 12905
rect 10136 12600 18179 12602
rect 10136 12542 10148 12600
rect 10206 12542 18179 12600
rect 10136 12540 18179 12542
rect 18303 12631 19490 12693
rect 10136 12530 10216 12540
rect 10136 12462 10216 12470
rect 18303 12462 18365 12631
rect 10136 12460 18365 12462
rect 10136 12402 10148 12460
rect 10206 12402 18365 12460
rect 10136 12400 18365 12402
rect 10136 12390 10216 12400
rect 18754 12356 19490 12428
rect 0 12316 1840 12326
rect 0 11380 10 12316
rect 710 11380 1840 12316
rect 18412 11552 18488 11554
rect 18754 11552 18826 12356
rect 18412 11544 18826 11552
rect 18412 11488 18422 11544
rect 18478 11488 18826 11544
rect 18412 11480 18826 11488
rect 19002 12078 19490 12150
rect 18412 11478 18488 11480
rect 18412 11278 18488 11280
rect 19002 11278 19074 12078
rect 18412 11270 19074 11278
rect 18412 11214 18422 11270
rect 18478 11214 19074 11270
rect 18412 11206 19074 11214
rect 19174 11814 19490 11886
rect 18412 11204 18488 11206
rect 18412 11006 18488 11008
rect 19174 11006 19246 11814
rect 18412 10998 19246 11006
rect 18412 10942 18422 10998
rect 18478 10942 19246 10998
rect 18412 10934 19246 10942
rect 18412 10932 18488 10934
rect 0 9518 10 10400
rect 710 9518 1840 10400
rect 0 9508 1840 9518
rect 18705 6373 19490 6435
rect 18204 5298 18284 5306
rect 18705 5298 18767 6373
rect 18204 5296 18767 5298
rect 18204 5238 18216 5296
rect 18274 5238 18767 5296
rect 18204 5236 18767 5238
rect 18871 6101 19490 6163
rect 18204 5226 18284 5236
rect 18204 5154 18284 5162
rect 18871 5154 18933 6101
rect 18204 5152 18933 5154
rect 18204 5094 18216 5152
rect 18274 5094 18933 5152
rect 18204 5092 18933 5094
rect 19053 5833 19490 5895
rect 18204 5082 18284 5092
rect 18204 3612 18284 3620
rect 19053 3612 19115 5833
rect 18204 3610 19115 3612
rect 18204 3552 18216 3610
rect 18274 3552 19115 3610
rect 18204 3550 19115 3552
rect 19219 5561 19490 5623
rect 18204 3540 18284 3550
rect 18204 3060 18284 3068
rect 19219 3060 19281 5561
rect 18204 3058 19281 3060
rect 18204 3000 18216 3058
rect 18274 3000 19281 3058
rect 18204 2998 19281 3000
rect 18204 2988 18284 2998
rect 18791 464 18969 469
rect 18174 284 18180 464
rect 18358 463 18970 464
rect 18358 285 18791 463
rect 18969 285 18970 463
rect 18358 284 18970 285
rect 18791 279 18969 284
<< via3 >>
rect 9728 44846 9792 44910
rect 21034 44902 21106 44906
rect 21034 44800 21038 44902
rect 21038 44800 21102 44902
rect 21102 44800 21106 44902
rect 21034 44796 21106 44800
rect 21586 44902 21658 44906
rect 21586 44800 21590 44902
rect 21590 44800 21654 44902
rect 21654 44800 21658 44902
rect 21586 44796 21658 44800
rect 22138 44902 22210 44906
rect 22138 44800 22142 44902
rect 22142 44800 22206 44902
rect 22206 44800 22210 44902
rect 22138 44796 22210 44800
rect 22690 44902 22762 44906
rect 22690 44800 22694 44902
rect 22694 44800 22758 44902
rect 22758 44800 22762 44902
rect 22690 44796 22762 44800
rect 23242 44902 23314 44906
rect 23242 44800 23246 44902
rect 23246 44800 23310 44902
rect 23310 44800 23314 44902
rect 23242 44796 23314 44800
rect 23794 44902 23866 44906
rect 23794 44800 23798 44902
rect 23798 44800 23862 44902
rect 23862 44800 23866 44902
rect 23794 44796 23866 44800
rect 24346 44902 24418 44906
rect 24346 44800 24350 44902
rect 24350 44800 24414 44902
rect 24414 44800 24418 44902
rect 24346 44796 24418 44800
rect 24898 44902 24970 44906
rect 24898 44800 24902 44902
rect 24902 44800 24966 44902
rect 24966 44800 24970 44902
rect 24898 44796 24970 44800
rect 25450 44902 25522 44906
rect 25450 44800 25454 44902
rect 25454 44800 25518 44902
rect 25518 44800 25522 44902
rect 25450 44796 25522 44800
rect 26002 44902 26074 44906
rect 26002 44800 26006 44902
rect 26006 44800 26070 44902
rect 26070 44800 26074 44902
rect 26002 44796 26074 44800
rect 26554 44902 26626 44906
rect 26554 44800 26558 44902
rect 26558 44800 26622 44902
rect 26622 44800 26626 44902
rect 26554 44796 26626 44800
rect 27106 44902 27178 44906
rect 27106 44800 27110 44902
rect 27110 44800 27174 44902
rect 27174 44800 27178 44902
rect 27106 44796 27178 44800
rect 27658 44902 27730 44906
rect 27658 44800 27662 44902
rect 27662 44800 27726 44902
rect 27726 44800 27730 44902
rect 27658 44796 27730 44800
rect 28210 44902 28282 44906
rect 28210 44800 28214 44902
rect 28214 44800 28278 44902
rect 28278 44800 28282 44902
rect 28210 44796 28282 44800
rect 28762 44902 28834 44906
rect 28762 44800 28766 44902
rect 28766 44800 28830 44902
rect 28830 44800 28834 44902
rect 28762 44796 28834 44800
rect 29314 44902 29386 44906
rect 29314 44800 29318 44902
rect 29318 44800 29382 44902
rect 29382 44800 29386 44902
rect 29314 44796 29386 44800
rect 546 43980 610 44044
rect 915 43840 1283 44210
rect 23690 43930 24000 44190
rect 30090 43930 30400 44190
rect 165 43290 533 43660
rect 23030 42980 23340 43280
rect 29430 42980 29740 43280
rect 18794 42528 18926 42640
rect 18242 42256 18374 42368
rect 17690 41984 17822 42096
rect 17138 41712 17270 41824
rect 16586 41440 16718 41552
rect 16034 41168 16166 41280
rect 15482 40896 15614 41008
rect 14930 40624 15062 40736
rect 14378 40352 14510 40464
rect 13826 40080 13958 40192
rect 10 36940 710 37744
rect 10 34946 710 35960
rect 17138 35472 17316 35652
rect 18363 35473 18541 35651
rect 17060 26542 17238 26722
rect 19129 26543 19307 26721
rect 10 24120 710 25030
rect 10 22232 710 23140
rect 17326 13818 17504 13998
rect 18777 13819 18955 13997
rect 10 11380 710 12316
rect 10 9518 710 10400
rect 18180 284 18358 464
rect 18791 285 18969 463
<< metal4 >>
rect 6134 44804 6194 45152
rect 6686 44804 6746 45152
rect 7238 44804 7298 45152
rect 7790 44804 7850 45152
rect 8342 44804 8402 45152
rect 8894 44804 8954 45152
rect 9446 44908 9506 45152
rect 9727 44910 9793 44911
rect 9727 44908 9728 44910
rect 9446 44848 9728 44908
rect 9727 44846 9728 44848
rect 9792 44908 9793 44910
rect 9998 44908 10058 45152
rect 9792 44848 10058 44908
rect 9792 44846 9793 44848
rect 9727 44845 9793 44846
rect 10550 44804 10610 45152
rect 11102 44804 11162 45152
rect 11654 44804 11714 45152
rect 12206 44804 12266 45152
rect 12758 44804 12818 45152
rect 13310 44804 13370 45152
rect 13862 44858 13922 45152
rect 14414 44858 14474 45152
rect 14966 44858 15026 45152
rect 15518 44858 15578 45152
rect 16070 44858 16130 45152
rect 16622 44858 16682 45152
rect 17174 44858 17234 45152
rect 17726 44858 17786 45152
rect 18278 44858 18338 45152
rect 18830 44858 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44912 21098 45152
rect 21590 44912 21650 45152
rect 22142 44912 22202 45152
rect 22694 44912 22754 45152
rect 23246 44912 23306 45152
rect 23798 44912 23858 45152
rect 24350 44912 24410 45152
rect 24902 44912 24962 45152
rect 25454 44912 25514 45152
rect 26006 44912 26066 45152
rect 26558 44912 26618 45152
rect 27110 44912 27170 45152
rect 27662 44912 27722 45152
rect 28214 44912 28274 45152
rect 28766 44912 28826 45152
rect 29318 44912 29378 45152
rect 21028 44906 21112 44912
rect 800 44704 9360 44804
rect 10144 44704 13440 44804
rect 800 44556 13440 44704
rect 800 44210 1520 44556
rect 0 44044 720 44152
rect 0 43980 546 44044
rect 610 43980 720 44044
rect 0 43660 720 43980
rect 0 43290 165 43660
rect 533 43290 720 43660
rect 0 37744 720 43290
rect 0 36940 10 37744
rect 710 36940 720 37744
rect 0 35960 720 36940
rect 0 34946 10 35960
rect 710 34946 720 35960
rect 0 25030 720 34946
rect 0 24120 10 25030
rect 710 24120 720 25030
rect 0 23140 720 24120
rect 0 22232 10 23140
rect 710 22232 720 23140
rect 0 12316 720 22232
rect 0 11380 10 12316
rect 710 11380 720 12316
rect 0 10400 720 11380
rect 0 9518 10 10400
rect 710 9518 720 10400
rect 0 1000 720 9518
rect 800 43840 915 44210
rect 1283 43840 1520 44210
rect 800 1000 1520 43840
rect 13822 40192 13962 44858
rect 13822 40080 13826 40192
rect 13958 40080 13962 40192
rect 13822 40028 13962 40080
rect 14374 40464 14514 44858
rect 14374 40352 14378 40464
rect 14510 40352 14514 40464
rect 14374 40028 14514 40352
rect 14926 40736 15066 44858
rect 14926 40624 14930 40736
rect 15062 40624 15066 40736
rect 14926 40028 15066 40624
rect 15478 41008 15618 44858
rect 15478 40896 15482 41008
rect 15614 40896 15618 41008
rect 15478 40028 15618 40896
rect 16030 41280 16170 44858
rect 16030 41168 16034 41280
rect 16166 41168 16170 41280
rect 16030 40028 16170 41168
rect 16582 41552 16722 44858
rect 16582 41440 16586 41552
rect 16718 41440 16722 41552
rect 16582 40028 16722 41440
rect 17134 41824 17274 44858
rect 17134 41712 17138 41824
rect 17270 41712 17274 41824
rect 17134 40028 17274 41712
rect 17686 42096 17826 44858
rect 17686 41984 17690 42096
rect 17822 41984 17826 42096
rect 17686 40028 17826 41984
rect 18238 42368 18378 44858
rect 18238 42256 18242 42368
rect 18374 42256 18378 42368
rect 18238 40028 18378 42256
rect 18790 42640 18930 44858
rect 21028 44796 21034 44906
rect 21106 44796 21112 44906
rect 21028 44790 21112 44796
rect 21580 44906 21664 44912
rect 21580 44796 21586 44906
rect 21658 44796 21664 44906
rect 21580 44790 21664 44796
rect 22132 44906 22216 44912
rect 22132 44796 22138 44906
rect 22210 44796 22216 44906
rect 22132 44790 22216 44796
rect 22684 44906 22768 44912
rect 22684 44796 22690 44906
rect 22762 44796 22768 44906
rect 22684 44790 22768 44796
rect 23236 44906 23320 44912
rect 23236 44796 23242 44906
rect 23314 44796 23320 44906
rect 23236 44790 23320 44796
rect 23788 44906 23872 44912
rect 23788 44796 23794 44906
rect 23866 44796 23872 44906
rect 23788 44790 23872 44796
rect 24340 44906 24424 44912
rect 24340 44796 24346 44906
rect 24418 44796 24424 44906
rect 24340 44790 24424 44796
rect 24892 44906 24976 44912
rect 24892 44796 24898 44906
rect 24970 44796 24976 44906
rect 24892 44790 24976 44796
rect 25444 44906 25528 44912
rect 25444 44796 25450 44906
rect 25522 44796 25528 44906
rect 25444 44790 25528 44796
rect 25996 44906 26080 44912
rect 25996 44796 26002 44906
rect 26074 44796 26080 44906
rect 25996 44790 26080 44796
rect 26548 44906 26632 44912
rect 26548 44796 26554 44906
rect 26626 44796 26632 44906
rect 26548 44790 26632 44796
rect 27100 44906 27184 44912
rect 27100 44796 27106 44906
rect 27178 44796 27184 44906
rect 27100 44790 27184 44796
rect 27652 44906 27736 44912
rect 27652 44796 27658 44906
rect 27730 44796 27736 44906
rect 27652 44790 27736 44796
rect 28204 44906 28288 44912
rect 28204 44796 28210 44906
rect 28282 44796 28288 44906
rect 28204 44790 28288 44796
rect 28756 44906 28840 44912
rect 28756 44796 28762 44906
rect 28834 44796 28840 44906
rect 28756 44790 28840 44796
rect 29308 44906 29392 44912
rect 29308 44796 29314 44906
rect 29386 44796 29392 44906
rect 29308 44790 29392 44796
rect 18790 42528 18794 42640
rect 18926 42528 18930 42640
rect 18790 40028 18930 42528
rect 23024 43280 23344 44200
rect 23024 42980 23030 43280
rect 23340 42980 23344 43280
rect 17137 35652 17317 35653
rect 15123 35613 17029 35626
rect 17137 35613 17138 35652
rect 15123 35536 17138 35613
rect 16973 35511 17138 35536
rect 17137 35472 17138 35511
rect 17316 35472 17317 35652
rect 17137 35471 17317 35472
rect 18362 35651 18542 35652
rect 18362 35473 18363 35651
rect 18541 35473 18542 35651
rect 17059 26722 17239 26723
rect 14942 26542 17060 26722
rect 17238 26542 17239 26722
rect 17059 26541 17239 26542
rect 17325 13998 17505 13999
rect 14942 13818 17326 13998
rect 17504 13818 17505 13998
rect 17325 13817 17505 13818
rect 14952 1120 15896 1300
rect 15716 464 15896 1120
rect 18362 756 18542 35473
rect 19120 26721 19320 26722
rect 19120 26543 19129 26721
rect 19307 26543 19320 26721
rect 19120 26542 19320 26543
rect 18760 13997 18960 14010
rect 18760 13819 18777 13997
rect 18955 13819 18960 13997
rect 18760 13810 18960 13819
rect 18776 884 18956 13810
rect 19128 1070 19308 26542
rect 19128 894 19880 1070
rect 23024 1000 23344 42980
rect 23684 44190 24004 44200
rect 23684 43930 23690 44190
rect 24000 43930 24004 44190
rect 23684 1000 24004 43930
rect 29424 43280 29744 44200
rect 29424 42980 29430 43280
rect 29740 42980 29744 43280
rect 29424 1000 29744 42980
rect 30084 44190 30404 44200
rect 30084 43930 30090 44190
rect 30400 43930 30404 44190
rect 30084 1000 30404 43930
rect 19128 890 30542 894
rect 18776 838 19012 884
rect 18776 806 19040 838
rect 18776 778 19076 806
rect 18820 760 19076 778
rect 18362 576 18662 756
rect 18820 744 19550 760
rect 18854 698 19550 744
rect 19700 714 30542 890
rect 18896 576 19550 698
rect 18179 464 18359 465
rect 15716 284 18180 464
rect 18358 284 18359 464
rect 18179 283 18359 284
rect 18482 210 18662 576
rect 19350 550 19550 576
rect 18790 463 19240 464
rect 18790 285 18791 463
rect 18969 285 19240 463
rect 19350 370 23490 550
rect 18790 284 19240 285
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18482 0 18950 210
rect 19060 180 19240 284
rect 22510 180 22820 210
rect 19060 0 22820 180
rect 23310 180 23490 370
rect 26350 180 26678 210
rect 23310 0 26678 180
rect 30362 0 30542 714
use controller_wrapper  controller_wrapper_0
timestamp 1762784779
transform 1 0 19368 0 1 900
box 0 496 12775 43900
use csdac255  dac_blue
timestamp 1762784779
transform -1 0 16108 0 1 1000
box -2130 0 14828 11424
use csdac255  dac_green
timestamp 1762784779
transform -1 0 16108 0 1 13714
box -2130 0 14828 11424
use csdac255  dac_red
timestamp 1762784779
transform -1 0 16108 0 1 26428
box -2130 0 14828 11424
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 0 1000 720 44152 0 FreeSans 3200 90 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1520 44152 0 FreeSans 3200 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 30084 1000 30404 44200 0 FreeSans 1600 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 29424 1000 29744 44200 0 FreeSans 1600 90 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 23684 1000 24004 44200 0 FreeSans 1600 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 23024 1000 23344 44200 0 FreeSans 1600 90 0 0 VDPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
