magic
tech sky130A
timestamp 1762784779
<< nwell >>
rect 0 0 837 287
<< pmos >>
rect 91 101 141 186
rect 187 101 287 186
rect 317 101 517 186
rect 546 101 746 186
<< pdiff >>
rect 62 182 91 186
rect 62 105 68 182
rect 85 105 91 182
rect 62 101 91 105
rect 141 182 187 186
rect 141 105 147 182
rect 181 105 187 182
rect 141 101 187 105
rect 287 182 317 186
rect 287 105 293 182
rect 311 105 317 182
rect 287 101 317 105
rect 517 182 546 186
rect 517 106 523 182
rect 540 106 546 182
rect 517 101 546 106
rect 746 182 775 186
rect 746 105 752 182
rect 769 105 775 182
rect 746 101 775 105
<< pdiffc >>
rect 68 105 85 182
rect 147 105 181 182
rect 293 105 311 182
rect 523 106 540 182
rect 752 105 769 182
<< nsubdiff >>
rect 18 252 52 269
rect 785 252 819 269
rect 18 235 35 252
rect 802 235 819 252
rect 18 35 35 52
rect 802 35 819 52
rect 18 18 52 35
rect 785 18 819 35
<< nsubdiffcont >>
rect 52 252 785 269
rect 18 52 35 235
rect 802 52 819 235
rect 52 18 785 35
<< poly >>
rect 91 227 141 236
rect 91 210 102 227
rect 130 210 141 227
rect 91 186 141 210
rect 187 227 287 236
rect 187 210 198 227
rect 276 210 287 227
rect 187 186 287 210
rect 317 227 517 236
rect 317 210 328 227
rect 506 210 517 227
rect 317 186 517 210
rect 546 227 746 236
rect 546 210 557 227
rect 735 210 746 227
rect 546 186 746 210
rect 91 77 141 101
rect 91 60 102 77
rect 130 60 141 77
rect 91 51 141 60
rect 187 77 287 101
rect 187 60 198 77
rect 276 60 287 77
rect 187 51 287 60
rect 317 77 517 101
rect 317 60 328 77
rect 506 60 517 77
rect 317 51 517 60
rect 546 77 746 101
rect 546 60 557 77
rect 735 60 746 77
rect 546 51 746 60
<< polycont >>
rect 102 210 130 227
rect 198 210 276 227
rect 328 210 506 227
rect 557 210 735 227
rect 102 60 130 77
rect 198 60 276 77
rect 328 60 506 77
rect 557 60 735 77
<< locali >>
rect 18 252 52 269
rect 785 252 819 269
rect 18 235 35 252
rect 102 229 130 235
rect 102 227 105 229
rect 127 227 130 229
rect 35 103 60 190
rect 82 182 85 190
rect 82 103 85 105
rect 35 97 85 103
rect 102 77 130 210
rect 198 229 276 235
rect 198 227 201 229
rect 223 227 276 229
rect 198 202 276 210
rect 147 184 181 190
rect 147 182 153 184
rect 175 182 181 184
rect 147 103 153 105
rect 175 103 181 105
rect 147 97 181 103
rect 102 52 130 60
rect 198 85 226 202
rect 293 184 311 252
rect 802 235 819 252
rect 198 77 276 85
rect 198 52 276 60
rect 18 35 35 52
rect 293 35 311 105
rect 328 229 506 235
rect 328 227 336 229
rect 358 227 506 229
rect 328 202 506 210
rect 557 227 735 235
rect 557 202 735 210
rect 328 85 356 202
rect 519 184 544 190
rect 519 103 520 184
rect 542 103 544 184
rect 519 97 544 103
rect 634 85 658 202
rect 752 187 802 190
rect 752 182 755 187
rect 752 100 755 105
rect 777 100 802 187
rect 752 97 802 100
rect 328 77 506 85
rect 328 52 506 60
rect 557 81 735 85
rect 557 77 693 81
rect 732 77 735 81
rect 557 55 693 60
rect 732 55 735 60
rect 557 52 735 55
rect 802 35 819 52
rect 18 18 52 35
rect 785 18 819 35
<< viali >>
rect 105 227 127 229
rect 105 210 127 227
rect 60 182 82 190
rect 60 105 68 182
rect 68 105 82 182
rect 60 103 82 105
rect 201 227 223 229
rect 201 210 223 227
rect 153 182 175 184
rect 153 105 175 182
rect 153 103 175 105
rect 1119 237 1288 254
rect 293 182 311 184
rect 293 105 311 182
rect 336 227 358 229
rect 336 210 358 227
rect 520 182 542 184
rect 520 106 523 182
rect 523 106 540 182
rect 540 106 542 182
rect 520 103 542 106
rect 755 182 777 187
rect 755 105 769 182
rect 769 105 777 182
rect 755 100 777 105
rect 693 77 732 81
rect 693 60 732 77
rect 693 55 732 60
rect 926 41 943 58
<< metal1 >>
rect 29 269 85 287
rect 29 190 85 241
rect 102 229 130 287
rect 102 210 105 229
rect 127 210 130 229
rect 102 204 130 210
rect 198 229 226 287
rect 198 210 201 229
rect 223 210 226 229
rect 198 204 226 210
rect 288 269 316 287
rect 29 103 60 190
rect 82 103 85 190
rect 29 97 85 103
rect 147 97 150 190
rect 178 97 181 190
rect 288 184 316 241
rect 333 229 361 287
rect 333 210 336 229
rect 358 210 361 229
rect 333 204 361 210
rect 752 269 780 287
rect 288 105 293 184
rect 311 105 316 184
rect 288 97 316 105
rect 514 186 549 190
rect 514 101 518 186
rect 545 101 549 186
rect 514 97 549 101
rect 752 187 780 241
rect 1116 254 1291 287
rect 1116 237 1119 254
rect 1288 237 1291 254
rect 752 100 755 187
rect 777 100 780 187
rect 752 94 780 100
rect 955 187 1017 190
rect 955 100 958 187
rect 1014 139 1017 187
rect 1116 167 1291 237
rect 1305 139 1335 167
rect 1014 100 1335 139
rect 690 83 735 87
rect 690 40 693 83
rect 732 40 735 83
rect 955 80 1335 100
rect 835 35 838 65
rect 864 58 951 65
rect 864 41 926 58
rect 943 41 951 58
rect 864 35 951 41
rect 1031 0 1088 80
<< via1 >>
rect 29 241 85 269
rect 288 241 316 269
rect 150 184 178 190
rect 150 103 153 184
rect 153 103 175 184
rect 175 103 178 184
rect 150 97 178 103
rect 752 241 780 269
rect 518 184 545 186
rect 518 103 520 184
rect 520 103 542 184
rect 542 103 545 184
rect 518 101 545 103
rect 958 100 1014 187
rect 693 81 732 83
rect 693 55 732 81
rect 693 40 732 55
rect 838 35 864 65
<< metal2 >>
rect 26 241 29 269
rect 85 241 288 269
rect 316 241 752 269
rect 780 241 783 269
rect 147 97 150 190
rect 178 187 1017 190
rect 178 186 958 187
rect 178 101 518 186
rect 545 101 958 186
rect 178 100 958 101
rect 1014 100 1017 187
rect 178 97 1017 100
rect 690 40 693 83
rect 732 60 735 83
rect 835 60 838 65
rect 732 40 838 60
rect 835 35 838 40
rect 864 35 867 65
use sky130_fd_pr__nfet_g5v0d10v5_VRH6W2  Mmirror
timestamp 1762784779
transform 0 1 1161 -1 0 139
box -139 -259 139 259
<< labels >>
flabel metal1 29 269 85 287 0 FreeSans 96 0 0 0 VPWR
port 9 nsew
flabel metal1 102 269 130 287 0 FreeSans 52 0 0 0 bias[2]
port 12 nsew
flabel metal1 198 269 226 287 0 FreeSans 52 0 0 0 bias[1]
port 13 nsew
flabel metal1 333 269 361 287 0 FreeSans 52 0 0 0 bias[0]
port 14 nsew
flabel metal1 1117 265 1186 287 0 FreeSans 96 0 0 0 VGND
port 15 nsew
flabel metal1 1031 0 1088 22 0 FreeSans 80 0 0 0 Vbias
port 17 nsew
<< end >>
