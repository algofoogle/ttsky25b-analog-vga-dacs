magic
tech sky130A
magscale 1 2
timestamp 1762665665
<< viali >>
rect 1777 42857 1811 42891
rect 3893 42857 3927 42891
rect 5273 42857 5307 42891
rect 10609 42857 10643 42891
rect 1133 42789 1167 42823
rect 6009 42789 6043 42823
rect 9045 42789 9079 42823
rect 10225 42789 10259 42823
rect 10425 42789 10459 42823
rect 10701 42789 10735 42823
rect 1869 42721 1903 42755
rect 3065 42721 3099 42755
rect 3985 42721 4019 42755
rect 6193 42721 6227 42755
rect 7297 42721 7331 42755
rect 8401 42721 8435 42755
rect 8585 42721 8619 42755
rect 8677 42721 8711 42755
rect 8769 42721 8803 42755
rect 9229 42721 9263 42755
rect 9413 42721 9447 42755
rect 9505 42721 9539 42755
rect 9689 42721 9723 42755
rect 2053 42653 2087 42687
rect 2789 42653 2823 42687
rect 3341 42653 3375 42687
rect 4261 42653 4295 42687
rect 5365 42653 5399 42687
rect 5457 42653 5491 42687
rect 6469 42653 6503 42687
rect 7573 42653 7607 42687
rect 1317 42585 1351 42619
rect 5825 42585 5859 42619
rect 9597 42585 9631 42619
rect 1409 42517 1443 42551
rect 4905 42517 4939 42551
rect 8953 42517 8987 42551
rect 10057 42517 10091 42551
rect 10241 42517 10275 42551
rect 6837 42245 6871 42279
rect 9781 42245 9815 42279
rect 2789 42177 2823 42211
rect 6101 42177 6135 42211
rect 7573 42177 7607 42211
rect 10609 42177 10643 42211
rect 1225 42109 1259 42143
rect 1317 42109 1351 42143
rect 1584 42109 1618 42143
rect 3249 42109 3283 42143
rect 4997 42109 5031 42143
rect 5641 42109 5675 42143
rect 6193 42109 6227 42143
rect 7113 42109 7147 42143
rect 7389 42109 7423 42143
rect 8401 42109 8435 42143
rect 2973 42041 3007 42075
rect 4752 42041 4786 42075
rect 7665 42041 7699 42075
rect 7757 42041 7791 42075
rect 7849 42041 7883 42075
rect 8033 42041 8067 42075
rect 8668 42041 8702 42075
rect 1041 41973 1075 42007
rect 2697 41973 2731 42007
rect 3433 41973 3467 42007
rect 3617 41973 3651 42007
rect 5089 41973 5123 42007
rect 8217 41973 8251 42007
rect 9965 41973 9999 42007
rect 3954 41701 3988 41735
rect 5457 41701 5491 41735
rect 5641 41701 5675 41735
rect 10425 41701 10459 41735
rect 1225 41633 1259 41667
rect 1317 41633 1351 41667
rect 1573 41633 1607 41667
rect 3249 41633 3283 41667
rect 3709 41633 3743 41667
rect 5273 41633 5307 41667
rect 5825 41633 5859 41667
rect 6009 41633 6043 41667
rect 7389 41633 7423 41667
rect 7757 41633 7791 41667
rect 8125 41633 8159 41667
rect 8217 41633 8251 41667
rect 8401 41633 8435 41667
rect 9790 41633 9824 41667
rect 10057 41633 10091 41667
rect 10609 41633 10643 41667
rect 3065 41565 3099 41599
rect 3157 41565 3191 41599
rect 5089 41497 5123 41531
rect 8677 41497 8711 41531
rect 1041 41429 1075 41463
rect 2697 41429 2731 41463
rect 3617 41429 3651 41463
rect 5917 41429 5951 41463
rect 8585 41429 8619 41463
rect 10241 41429 10275 41463
rect 1041 41225 1075 41259
rect 9229 41225 9263 41259
rect 3433 41157 3467 41191
rect 6837 41157 6871 41191
rect 3709 41089 3743 41123
rect 6101 41089 6135 41123
rect 1225 41021 1259 41055
rect 1593 41021 1627 41055
rect 1685 41021 1719 41055
rect 3249 41021 3283 41055
rect 5365 41021 5399 41055
rect 5917 41021 5951 41055
rect 8217 41021 8251 41055
rect 8585 41021 8619 41055
rect 8769 41021 8803 41055
rect 8861 41021 8895 41055
rect 8953 41021 8987 41055
rect 9321 41021 9355 41055
rect 1317 40953 1351 40987
rect 1409 40953 1443 40987
rect 1930 40953 1964 40987
rect 3976 40953 4010 40987
rect 7950 40953 7984 40987
rect 9588 40953 9622 40987
rect 3065 40885 3099 40919
rect 5089 40885 5123 40919
rect 5273 40885 5307 40919
rect 6653 40885 6687 40919
rect 10701 40885 10735 40919
rect 3341 40681 3375 40715
rect 4445 40681 4479 40715
rect 5457 40681 5491 40715
rect 7221 40681 7255 40715
rect 7941 40681 7975 40715
rect 8585 40681 8619 40715
rect 10149 40681 10183 40715
rect 6653 40613 6687 40647
rect 7021 40613 7055 40647
rect 8401 40613 8435 40647
rect 1133 40545 1167 40579
rect 1501 40545 1535 40579
rect 1849 40545 1883 40579
rect 3065 40545 3099 40579
rect 5457 40545 5491 40579
rect 7481 40545 7515 40579
rect 7757 40545 7791 40579
rect 8677 40545 8711 40579
rect 8944 40545 8978 40579
rect 10425 40545 10459 40579
rect 10517 40545 10551 40579
rect 10609 40545 10643 40579
rect 10793 40545 10827 40579
rect 1593 40477 1627 40511
rect 3893 40477 3927 40511
rect 4537 40477 4571 40511
rect 4721 40477 4755 40511
rect 4905 40477 4939 40511
rect 5549 40477 5583 40511
rect 6101 40477 6135 40511
rect 7573 40477 7607 40511
rect 8033 40477 8067 40511
rect 7389 40409 7423 40443
rect 949 40341 983 40375
rect 1317 40341 1351 40375
rect 2973 40341 3007 40375
rect 3157 40341 3191 40375
rect 4077 40341 4111 40375
rect 7205 40341 7239 40375
rect 8401 40341 8435 40375
rect 10057 40341 10091 40375
rect 1501 40137 1535 40171
rect 3985 40137 4019 40171
rect 8677 40137 8711 40171
rect 9045 40137 9079 40171
rect 9229 40137 9263 40171
rect 9781 40137 9815 40171
rect 5733 40069 5767 40103
rect 1317 40001 1351 40035
rect 2881 40001 2915 40035
rect 3433 40001 3467 40035
rect 4629 40001 4663 40035
rect 7113 40001 7147 40035
rect 10057 40001 10091 40035
rect 1225 39933 1259 39967
rect 1685 39933 1719 39967
rect 1869 39933 1903 39967
rect 1961 39933 1995 39967
rect 2053 39933 2087 39967
rect 2329 39933 2363 39967
rect 4077 39933 4111 39967
rect 4813 39933 4847 39967
rect 5181 39933 5215 39967
rect 5457 39933 5491 39967
rect 5641 39933 5675 39967
rect 7757 39933 7791 39967
rect 7941 39933 7975 39967
rect 8401 39933 8435 39967
rect 9137 39933 9171 39967
rect 9413 39933 9447 39967
rect 10241 39933 10275 39967
rect 4997 39865 5031 39899
rect 5089 39865 5123 39899
rect 6846 39865 6880 39899
rect 8677 39865 8711 39899
rect 8769 39865 8803 39899
rect 9781 39865 9815 39899
rect 10425 39865 10459 39899
rect 10701 39865 10735 39899
rect 2237 39797 2271 39831
rect 5365 39797 5399 39831
rect 5549 39797 5583 39831
rect 7205 39797 7239 39831
rect 8125 39797 8159 39831
rect 8493 39797 8527 39831
rect 8861 39797 8895 39831
rect 9965 39797 9999 39831
rect 10609 39797 10643 39831
rect 1685 39593 1719 39627
rect 4169 39593 4203 39627
rect 6653 39593 6687 39627
rect 7113 39593 7147 39627
rect 7757 39593 7791 39627
rect 10793 39593 10827 39627
rect 4077 39525 4111 39559
rect 7021 39525 7055 39559
rect 1317 39457 1351 39491
rect 1409 39457 1443 39491
rect 1593 39457 1627 39491
rect 2412 39457 2446 39491
rect 3893 39457 3927 39491
rect 4537 39457 4571 39491
rect 4997 39457 5031 39491
rect 5825 39457 5859 39491
rect 6009 39457 6043 39491
rect 6285 39457 6319 39491
rect 6469 39457 6503 39491
rect 7481 39457 7515 39491
rect 7665 39457 7699 39491
rect 7849 39457 7883 39491
rect 8125 39457 8159 39491
rect 8953 39457 8987 39491
rect 9321 39457 9355 39491
rect 9680 39457 9714 39491
rect 2145 39389 2179 39423
rect 3709 39389 3743 39423
rect 4629 39389 4663 39423
rect 4813 39389 4847 39423
rect 5641 39389 5675 39423
rect 7297 39389 7331 39423
rect 8401 39389 8435 39423
rect 9413 39389 9447 39423
rect 1133 39253 1167 39287
rect 1869 39253 1903 39287
rect 3525 39253 3559 39287
rect 8033 39253 8067 39287
rect 8493 39253 8527 39287
rect 8677 39253 8711 39287
rect 8769 39253 8803 39287
rect 9229 39253 9263 39287
rect 949 39049 983 39083
rect 3249 39049 3283 39083
rect 5733 39049 5767 39083
rect 6837 39049 6871 39083
rect 8125 39049 8159 39083
rect 9137 39049 9171 39083
rect 9781 39049 9815 39083
rect 1409 38981 1443 39015
rect 3065 38981 3099 39015
rect 5181 38981 5215 39015
rect 9689 38981 9723 39015
rect 1685 38913 1719 38947
rect 5365 38913 5399 38947
rect 7021 38913 7055 38947
rect 7113 38913 7147 38947
rect 7849 38913 7883 38947
rect 857 38845 891 38879
rect 1041 38845 1075 38879
rect 3433 38845 3467 38879
rect 3525 38845 3559 38879
rect 3801 38845 3835 38879
rect 5549 38845 5583 38879
rect 5825 38845 5859 38879
rect 6561 38845 6595 38879
rect 7389 38845 7423 38879
rect 7481 38845 7515 38879
rect 7665 38845 7699 38879
rect 7757 38845 7791 38879
rect 7941 38845 7975 38879
rect 8585 38845 8619 38879
rect 8677 38845 8711 38879
rect 8861 38845 8895 38879
rect 8953 38845 8987 38879
rect 9413 38845 9447 38879
rect 9505 38845 9539 38879
rect 9965 38845 9999 38879
rect 10149 38845 10183 38879
rect 10425 38845 10459 38879
rect 1133 38777 1167 38811
rect 1930 38777 1964 38811
rect 4068 38777 4102 38811
rect 9045 38777 9079 38811
rect 10609 38777 10643 38811
rect 1593 38709 1627 38743
rect 5917 38709 5951 38743
rect 7205 38709 7239 38743
rect 8401 38709 8435 38743
rect 10241 38709 10275 38743
rect 1317 38505 1351 38539
rect 1777 38505 1811 38539
rect 3985 38505 4019 38539
rect 6193 38505 6227 38539
rect 7297 38505 7331 38539
rect 8217 38505 8251 38539
rect 9137 38505 9171 38539
rect 10425 38505 10459 38539
rect 949 38437 983 38471
rect 2136 38437 2170 38471
rect 3709 38437 3743 38471
rect 6285 38437 6319 38471
rect 7665 38437 7699 38471
rect 1179 38403 1213 38437
rect 1593 38369 1627 38403
rect 3433 38369 3467 38403
rect 3617 38369 3651 38403
rect 3801 38369 3835 38403
rect 5201 38369 5235 38403
rect 5457 38369 5491 38403
rect 6837 38369 6871 38403
rect 7113 38369 7147 38403
rect 7573 38369 7607 38403
rect 7757 38369 7791 38403
rect 8033 38369 8067 38403
rect 8401 38369 8435 38403
rect 8861 38369 8895 38403
rect 9505 38369 9539 38403
rect 9965 38369 9999 38403
rect 10241 38369 10275 38403
rect 10517 38369 10551 38403
rect 1409 38301 1443 38335
rect 1869 38301 1903 38335
rect 6377 38301 6411 38335
rect 6929 38301 6963 38335
rect 8677 38301 8711 38335
rect 8769 38301 8803 38335
rect 9229 38301 9263 38335
rect 10149 38301 10183 38335
rect 5825 38233 5859 38267
rect 7389 38233 7423 38267
rect 8585 38233 8619 38267
rect 1133 38165 1167 38199
rect 3249 38165 3283 38199
rect 4077 38165 4111 38199
rect 7021 38165 7055 38199
rect 7941 38165 7975 38199
rect 9321 38165 9355 38199
rect 9689 38165 9723 38199
rect 9965 38165 9999 38199
rect 10701 38165 10735 38199
rect 949 37961 983 37995
rect 2145 37961 2179 37995
rect 2513 37961 2547 37995
rect 2973 37961 3007 37995
rect 7205 37961 7239 37995
rect 7389 37961 7423 37995
rect 7849 37961 7883 37995
rect 8401 37961 8435 37995
rect 8861 37961 8895 37995
rect 9597 37961 9631 37995
rect 3249 37893 3283 37927
rect 1869 37825 1903 37859
rect 3801 37825 3835 37859
rect 4813 37825 4847 37859
rect 6929 37825 6963 37859
rect 7941 37825 7975 37859
rect 8953 37825 8987 37859
rect 9597 37825 9631 37859
rect 1133 37757 1167 37791
rect 1593 37757 1627 37791
rect 1777 37757 1811 37791
rect 1961 37757 1995 37791
rect 2329 37757 2363 37791
rect 2789 37757 2823 37791
rect 3617 37757 3651 37791
rect 5549 37757 5583 37791
rect 6009 37757 6043 37791
rect 6745 37757 6779 37791
rect 7757 37757 7791 37791
rect 8217 37757 8251 37791
rect 8677 37757 8711 37791
rect 8769 37757 8803 37791
rect 9137 37757 9171 37791
rect 9395 37757 9429 37791
rect 10701 37757 10735 37791
rect 4629 37689 4663 37723
rect 6561 37689 6595 37723
rect 7021 37689 7055 37723
rect 7237 37689 7271 37723
rect 9873 37689 9907 37723
rect 1409 37621 1443 37655
rect 3709 37621 3743 37655
rect 4261 37621 4295 37655
rect 4721 37621 4755 37655
rect 6377 37621 6411 37655
rect 7573 37621 7607 37655
rect 9229 37621 9263 37655
rect 10149 37621 10183 37655
rect 2881 37417 2915 37451
rect 4261 37417 4295 37451
rect 4721 37417 4755 37451
rect 5089 37417 5123 37451
rect 6561 37417 6595 37451
rect 8217 37417 8251 37451
rect 8861 37417 8895 37451
rect 1317 37349 1351 37383
rect 3801 37349 3835 37383
rect 6469 37349 6503 37383
rect 9045 37349 9079 37383
rect 9496 37349 9530 37383
rect 1133 37281 1167 37315
rect 1409 37281 1443 37315
rect 1676 37281 1710 37315
rect 3249 37281 3283 37315
rect 3709 37281 3743 37315
rect 3893 37281 3927 37315
rect 3985 37281 4019 37315
rect 4169 37281 4203 37315
rect 4629 37281 4663 37315
rect 5273 37281 5307 37315
rect 5365 37281 5399 37315
rect 5457 37281 5491 37315
rect 5641 37281 5675 37315
rect 5825 37281 5859 37315
rect 6009 37281 6043 37315
rect 6285 37281 6319 37315
rect 7297 37281 7331 37315
rect 7481 37281 7515 37315
rect 7665 37281 7699 37315
rect 8309 37281 8343 37315
rect 8953 37281 8987 37315
rect 9137 37281 9171 37315
rect 949 37213 983 37247
rect 3341 37213 3375 37247
rect 3433 37213 3467 37247
rect 4813 37213 4847 37247
rect 7205 37213 7239 37247
rect 7941 37213 7975 37247
rect 8585 37213 8619 37247
rect 9229 37213 9263 37247
rect 2789 37145 2823 37179
rect 4169 37145 4203 37179
rect 7297 37077 7331 37111
rect 7757 37077 7791 37111
rect 8401 37077 8435 37111
rect 10609 37077 10643 37111
rect 1041 36873 1075 36907
rect 5457 36873 5491 36907
rect 9505 36873 9539 36907
rect 10333 36873 10367 36907
rect 7297 36805 7331 36839
rect 9045 36805 9079 36839
rect 10149 36805 10183 36839
rect 1225 36737 1259 36771
rect 3341 36737 3375 36771
rect 8493 36737 8527 36771
rect 9413 36737 9447 36771
rect 949 36669 983 36703
rect 1133 36669 1167 36703
rect 1501 36669 1535 36703
rect 3985 36669 4019 36703
rect 4252 36669 4286 36703
rect 5641 36669 5675 36703
rect 5825 36669 5859 36703
rect 6009 36669 6043 36703
rect 6193 36669 6227 36703
rect 6561 36669 6595 36703
rect 7481 36669 7515 36703
rect 7757 36669 7791 36703
rect 7941 36669 7975 36703
rect 8033 36669 8067 36703
rect 8401 36669 8435 36703
rect 8585 36669 8619 36703
rect 9137 36669 9171 36703
rect 9505 36669 9539 36703
rect 10609 36669 10643 36703
rect 10793 36669 10827 36703
rect 2881 36601 2915 36635
rect 5733 36601 5767 36635
rect 7665 36601 7699 36635
rect 8677 36601 8711 36635
rect 8861 36601 8895 36635
rect 9873 36601 9907 36635
rect 10057 36601 10091 36635
rect 10301 36601 10335 36635
rect 10517 36601 10551 36635
rect 3893 36533 3927 36567
rect 5365 36533 5399 36567
rect 7205 36533 7239 36567
rect 7849 36533 7883 36567
rect 8217 36533 8251 36567
rect 9229 36533 9263 36567
rect 9689 36533 9723 36567
rect 10701 36533 10735 36567
rect 2421 36329 2455 36363
rect 3341 36329 3375 36363
rect 3801 36329 3835 36363
rect 5365 36329 5399 36363
rect 5549 36329 5583 36363
rect 7573 36329 7607 36363
rect 8217 36329 8251 36363
rect 9153 36329 9187 36363
rect 10793 36329 10827 36363
rect 4230 36261 4264 36295
rect 8953 36261 8987 36295
rect 9658 36261 9692 36295
rect 1041 36193 1075 36227
rect 1297 36193 1331 36227
rect 2881 36193 2915 36227
rect 2973 36193 3007 36227
rect 3617 36193 3651 36227
rect 3801 36193 3835 36227
rect 3985 36193 4019 36227
rect 5457 36193 5491 36227
rect 5641 36193 5675 36227
rect 6009 36193 6043 36227
rect 7849 36193 7883 36227
rect 8125 36193 8159 36227
rect 8309 36193 8343 36227
rect 8401 36193 8435 36227
rect 8585 36193 8619 36227
rect 8677 36193 8711 36227
rect 9413 36193 9447 36227
rect 2789 36125 2823 36159
rect 5825 36125 5859 36159
rect 6285 36125 6319 36159
rect 7113 36125 7147 36159
rect 7481 36125 7515 36159
rect 8033 36125 8067 36159
rect 6193 36057 6227 36091
rect 9321 36057 9355 36091
rect 8585 35989 8619 36023
rect 8769 35989 8803 36023
rect 9137 35989 9171 36023
rect 1409 35785 1443 35819
rect 8493 35785 8527 35819
rect 8769 35785 8803 35819
rect 9597 35785 9631 35819
rect 10057 35785 10091 35819
rect 3433 35717 3467 35751
rect 5733 35717 5767 35751
rect 1133 35649 1167 35683
rect 1501 35649 1535 35683
rect 3709 35649 3743 35683
rect 8125 35649 8159 35683
rect 9137 35649 9171 35683
rect 9229 35649 9263 35683
rect 1041 35581 1075 35615
rect 1757 35581 1791 35615
rect 3525 35581 3559 35615
rect 4353 35581 4387 35615
rect 6377 35581 6411 35615
rect 7573 35581 7607 35615
rect 7941 35581 7975 35615
rect 8585 35581 8619 35615
rect 8953 35581 8987 35615
rect 10517 35581 10551 35615
rect 4261 35513 4295 35547
rect 4598 35513 4632 35547
rect 6561 35513 6595 35547
rect 9965 35513 9999 35547
rect 2881 35445 2915 35479
rect 5825 35445 5859 35479
rect 7757 35445 7791 35479
rect 9597 35445 9631 35479
rect 9781 35445 9815 35479
rect 10609 35445 10643 35479
rect 2881 35241 2915 35275
rect 4077 35241 4111 35275
rect 4537 35241 4571 35275
rect 4905 35241 4939 35275
rect 6469 35241 6503 35275
rect 8677 35241 8711 35275
rect 9413 35241 9447 35275
rect 3801 35173 3835 35207
rect 6745 35173 6779 35207
rect 8585 35173 8619 35207
rect 10526 35173 10560 35207
rect 1317 35105 1351 35139
rect 1593 35105 1627 35139
rect 2421 35105 2455 35139
rect 2881 35105 2915 35139
rect 3065 35105 3099 35139
rect 3157 35105 3191 35139
rect 3893 35105 3927 35139
rect 4149 35105 4183 35139
rect 4261 35105 4295 35139
rect 5365 35105 5399 35139
rect 5549 35105 5583 35139
rect 6009 35105 6043 35139
rect 6101 35105 6135 35139
rect 6837 35105 6871 35139
rect 7389 35105 7423 35139
rect 8125 35105 8159 35139
rect 8309 35105 8343 35139
rect 8953 35105 8987 35139
rect 1685 35037 1719 35071
rect 2237 35037 2271 35071
rect 2329 35037 2363 35071
rect 4997 35037 5031 35071
rect 5089 35037 5123 35071
rect 6193 35037 6227 35071
rect 6285 35037 6319 35071
rect 7113 35037 7147 35071
rect 7941 35037 7975 35071
rect 9045 35037 9079 35071
rect 10793 35037 10827 35071
rect 1961 34969 1995 35003
rect 4445 34969 4479 35003
rect 8493 34969 8527 35003
rect 8861 34969 8895 35003
rect 1133 34901 1167 34935
rect 2789 34901 2823 34935
rect 5457 34901 5491 34935
rect 1317 34697 1351 34731
rect 2973 34697 3007 34731
rect 4445 34697 4479 34731
rect 5089 34697 5123 34731
rect 5181 34697 5215 34731
rect 5549 34697 5583 34731
rect 7113 34697 7147 34731
rect 10057 34697 10091 34731
rect 10517 34629 10551 34663
rect 10793 34629 10827 34663
rect 3985 34561 4019 34595
rect 5273 34561 5307 34595
rect 6837 34561 6871 34595
rect 8493 34561 8527 34595
rect 1133 34493 1167 34527
rect 2441 34493 2475 34527
rect 2697 34493 2731 34527
rect 2789 34493 2823 34527
rect 3341 34493 3375 34527
rect 3801 34493 3835 34527
rect 4077 34493 4111 34527
rect 4537 34493 4571 34527
rect 4721 34493 4755 34527
rect 4813 34493 4847 34527
rect 4905 34493 4939 34527
rect 5181 34493 5215 34527
rect 6285 34493 6319 34527
rect 6469 34493 6503 34527
rect 6653 34493 6687 34527
rect 6929 34493 6963 34527
rect 7113 34493 7147 34527
rect 7481 34493 7515 34527
rect 7573 34493 7607 34527
rect 7757 34493 7791 34527
rect 8033 34493 8067 34527
rect 8217 34493 8251 34527
rect 8401 34493 8435 34527
rect 8585 34493 8619 34527
rect 8677 34493 8711 34527
rect 10241 34493 10275 34527
rect 10333 34493 10367 34527
rect 10609 34493 10643 34527
rect 10793 34493 10827 34527
rect 3525 34425 3559 34459
rect 8922 34425 8956 34459
rect 10517 34425 10551 34459
rect 949 34357 983 34391
rect 5733 34357 5767 34391
rect 8217 34357 8251 34391
rect 5825 34153 5859 34187
rect 7573 34153 7607 34187
rect 8861 34153 8895 34187
rect 9597 34153 9631 34187
rect 10425 34153 10459 34187
rect 9229 34085 9263 34119
rect 10149 34085 10183 34119
rect 1584 34017 1618 34051
rect 3424 34017 3458 34051
rect 4905 34017 4939 34051
rect 5089 34017 5123 34051
rect 5181 34017 5215 34051
rect 5365 34017 5399 34051
rect 5641 34017 5675 34051
rect 6938 34017 6972 34051
rect 7205 34017 7239 34051
rect 7757 34017 7791 34051
rect 7849 34017 7883 34051
rect 8033 34017 8067 34051
rect 8585 34017 8619 34051
rect 8953 34017 8987 34051
rect 9413 34017 9447 34051
rect 9873 34017 9907 34051
rect 10701 34017 10735 34051
rect 1317 33949 1351 33983
rect 3157 33949 3191 33983
rect 4997 33949 5031 33983
rect 8217 33949 8251 33983
rect 9689 33949 9723 33983
rect 10425 33949 10459 33983
rect 4537 33881 4571 33915
rect 5549 33881 5583 33915
rect 8125 33881 8159 33915
rect 8401 33881 8435 33915
rect 10609 33881 10643 33915
rect 2697 33813 2731 33847
rect 5273 33813 5307 33847
rect 8217 33813 8251 33847
rect 10241 33813 10275 33847
rect 1961 33609 1995 33643
rect 3525 33609 3559 33643
rect 5273 33609 5307 33643
rect 8125 33609 8159 33643
rect 2789 33541 2823 33575
rect 5457 33541 5491 33575
rect 6009 33541 6043 33575
rect 9597 33541 9631 33575
rect 10333 33541 10367 33575
rect 1685 33473 1719 33507
rect 2513 33473 2547 33507
rect 4077 33473 4111 33507
rect 5844 33473 5878 33507
rect 9321 33473 9355 33507
rect 1133 33405 1167 33439
rect 1317 33405 1351 33439
rect 1409 33405 1443 33439
rect 1501 33405 1535 33439
rect 3065 33405 3099 33439
rect 3893 33405 3927 33439
rect 5089 33405 5123 33439
rect 5549 33405 5583 33439
rect 5641 33405 5675 33439
rect 5733 33405 5767 33439
rect 5927 33405 5961 33439
rect 6285 33405 6319 33439
rect 6377 33405 6411 33439
rect 6531 33405 6565 33439
rect 7481 33405 7515 33439
rect 7849 33405 7883 33439
rect 8033 33405 8067 33439
rect 8217 33405 8251 33439
rect 8401 33405 8435 33439
rect 8493 33405 8527 33439
rect 8769 33405 8803 33439
rect 8861 33405 8895 33439
rect 10057 33405 10091 33439
rect 10149 33405 10183 33439
rect 10425 33405 10459 33439
rect 1685 33337 1719 33371
rect 2789 33337 2823 33371
rect 6009 33337 6043 33371
rect 6837 33337 6871 33371
rect 8677 33337 8711 33371
rect 10333 33337 10367 33371
rect 949 33269 983 33303
rect 2329 33269 2363 33303
rect 2421 33269 2455 33303
rect 2973 33269 3007 33303
rect 3985 33269 4019 33303
rect 6193 33269 6227 33303
rect 6745 33269 6779 33303
rect 9045 33269 9079 33303
rect 9781 33269 9815 33303
rect 10609 33269 10643 33303
rect 2881 33065 2915 33099
rect 7757 33065 7791 33099
rect 8861 33065 8895 33099
rect 9137 33065 9171 33099
rect 10701 33065 10735 33099
rect 949 32997 983 33031
rect 3341 32997 3375 33031
rect 6377 32997 6411 33031
rect 9045 32997 9079 33031
rect 10250 32997 10284 33031
rect 1133 32929 1167 32963
rect 1593 32929 1627 32963
rect 1777 32929 1811 32963
rect 2145 32929 2179 32963
rect 2697 32929 2731 32963
rect 2973 32929 3007 32963
rect 3157 32929 3191 32963
rect 3617 32929 3651 32963
rect 3709 32929 3743 32963
rect 3893 32929 3927 32963
rect 4261 32929 4295 32963
rect 4353 32929 4387 32963
rect 4537 32929 4571 32963
rect 5273 32929 5307 32963
rect 5549 32929 5583 32963
rect 5917 32929 5951 32963
rect 6101 32929 6135 32963
rect 6193 32929 6227 32963
rect 6837 32929 6871 32963
rect 7021 32929 7055 32963
rect 7481 32929 7515 32963
rect 8217 32929 8251 32963
rect 8401 32929 8435 32963
rect 8493 32929 8527 32963
rect 8677 32929 8711 32963
rect 8769 32929 8803 32963
rect 10609 32929 10643 32963
rect 10793 32929 10827 32963
rect 6745 32861 6779 32895
rect 7297 32861 7331 32895
rect 7941 32861 7975 32895
rect 8033 32861 8067 32895
rect 8125 32861 8159 32895
rect 10517 32861 10551 32895
rect 1317 32793 1351 32827
rect 4445 32793 4479 32827
rect 6009 32793 6043 32827
rect 8401 32793 8435 32827
rect 9045 32793 9079 32827
rect 2513 32725 2547 32759
rect 4077 32725 4111 32759
rect 4721 32725 4755 32759
rect 5089 32725 5123 32759
rect 5457 32725 5491 32759
rect 6469 32725 6503 32759
rect 6837 32725 6871 32759
rect 7113 32725 7147 32759
rect 7665 32725 7699 32759
rect 2513 32521 2547 32555
rect 6101 32521 6135 32555
rect 6285 32521 6319 32555
rect 7113 32521 7147 32555
rect 9413 32521 9447 32555
rect 6653 32453 6687 32487
rect 8769 32453 8803 32487
rect 2237 32385 2271 32419
rect 5917 32385 5951 32419
rect 6929 32385 6963 32419
rect 7389 32385 7423 32419
rect 8217 32385 8251 32419
rect 10793 32385 10827 32419
rect 1981 32317 2015 32351
rect 2881 32317 2915 32351
rect 3801 32317 3835 32351
rect 5273 32317 5307 32351
rect 6101 32317 6135 32351
rect 6469 32317 6503 32351
rect 6561 32317 6595 32351
rect 6745 32317 6779 32351
rect 7481 32317 7515 32351
rect 8493 32317 8527 32351
rect 8585 32317 8619 32351
rect 8953 32317 8987 32351
rect 9045 32317 9079 32351
rect 9229 32317 9263 32351
rect 2513 32249 2547 32283
rect 3617 32249 3651 32283
rect 4068 32249 4102 32283
rect 5641 32249 5675 32283
rect 7021 32249 7055 32283
rect 8033 32249 8067 32283
rect 10526 32249 10560 32283
rect 857 32181 891 32215
rect 2329 32181 2363 32215
rect 3525 32181 3559 32215
rect 5181 32181 5215 32215
rect 5457 32181 5491 32215
rect 7665 32181 7699 32215
rect 3801 31977 3835 32011
rect 5641 31977 5675 32011
rect 6193 31977 6227 32011
rect 7021 31977 7055 32011
rect 7113 31977 7147 32011
rect 8217 31977 8251 32011
rect 10701 31977 10735 32011
rect 3893 31909 3927 31943
rect 5825 31909 5859 31943
rect 8953 31909 8987 31943
rect 9505 31909 9539 31943
rect 949 31841 983 31875
rect 1205 31841 1239 31875
rect 2421 31841 2455 31875
rect 2688 31841 2722 31875
rect 4905 31841 4939 31875
rect 5273 31841 5307 31875
rect 6009 31841 6043 31875
rect 6469 31841 6503 31875
rect 6837 31841 6871 31875
rect 7297 31841 7331 31875
rect 7389 31841 7423 31875
rect 7481 31841 7515 31875
rect 7757 31841 7791 31875
rect 7941 31841 7975 31875
rect 8033 31841 8067 31875
rect 8493 31841 8527 31875
rect 9137 31841 9171 31875
rect 10241 31841 10275 31875
rect 10425 31841 10459 31875
rect 10517 31841 10551 31875
rect 5181 31773 5215 31807
rect 5365 31773 5399 31807
rect 5457 31773 5491 31807
rect 6377 31773 6411 31807
rect 9965 31773 9999 31807
rect 10057 31773 10091 31807
rect 10149 31773 10183 31807
rect 10701 31773 10735 31807
rect 2329 31705 2363 31739
rect 7665 31705 7699 31739
rect 8769 31705 8803 31739
rect 9781 31705 9815 31739
rect 6745 31637 6779 31671
rect 8033 31637 8067 31671
rect 8401 31637 8435 31671
rect 9505 31637 9539 31671
rect 9689 31637 9723 31671
rect 1133 31433 1167 31467
rect 1317 31433 1351 31467
rect 4813 31433 4847 31467
rect 5641 31433 5675 31467
rect 6009 31433 6043 31467
rect 6561 31433 6595 31467
rect 6929 31433 6963 31467
rect 7113 31433 7147 31467
rect 8769 31433 8803 31467
rect 4629 31365 4663 31399
rect 5273 31297 5307 31331
rect 5365 31297 5399 31331
rect 6837 31297 6871 31331
rect 1593 31229 1627 31263
rect 1869 31229 1903 31263
rect 2145 31229 2179 31263
rect 2421 31229 2455 31263
rect 2605 31229 2639 31263
rect 2697 31229 2731 31263
rect 2789 31229 2823 31263
rect 3249 31229 3283 31263
rect 4997 31229 5031 31263
rect 5089 31229 5123 31263
rect 6193 31229 6227 31263
rect 6377 31229 6411 31263
rect 6653 31229 6687 31263
rect 6929 31229 6963 31263
rect 7849 31229 7883 31263
rect 9882 31229 9916 31263
rect 10149 31229 10183 31263
rect 949 31161 983 31195
rect 1165 31161 1199 31195
rect 2329 31161 2363 31195
rect 3065 31161 3099 31195
rect 3494 31161 3528 31195
rect 5457 31161 5491 31195
rect 5733 31161 5767 31195
rect 5917 31161 5951 31195
rect 7297 31161 7331 31195
rect 8033 31161 8067 31195
rect 8585 31161 8619 31195
rect 10333 31161 10367 31195
rect 1409 31093 1443 31127
rect 1777 31093 1811 31127
rect 1961 31093 1995 31127
rect 7389 31093 7423 31127
rect 8217 31093 8251 31127
rect 8493 31093 8527 31127
rect 10425 31093 10459 31127
rect 1041 30889 1075 30923
rect 3157 30889 3191 30923
rect 3325 30889 3359 30923
rect 4077 30889 4111 30923
rect 5549 30889 5583 30923
rect 6377 30889 6411 30923
rect 6561 30889 6595 30923
rect 9413 30889 9447 30923
rect 1209 30821 1243 30855
rect 1409 30821 1443 30855
rect 1869 30821 1903 30855
rect 2513 30821 2547 30855
rect 3525 30821 3559 30855
rect 10526 30821 10560 30855
rect 1685 30753 1719 30787
rect 1961 30753 1995 30787
rect 2053 30753 2087 30787
rect 2145 30753 2179 30787
rect 2329 30753 2363 30787
rect 2789 30753 2823 30787
rect 5365 30753 5399 30787
rect 5457 30753 5491 30787
rect 5825 30753 5859 30787
rect 6469 30753 6503 30787
rect 6653 30753 6687 30787
rect 7389 30753 7423 30787
rect 7573 30753 7607 30787
rect 8033 30753 8067 30787
rect 8217 30753 8251 30787
rect 8309 30753 8343 30787
rect 8953 30753 8987 30787
rect 3065 30685 3099 30719
rect 6101 30685 6135 30719
rect 7113 30685 7147 30719
rect 7297 30685 7331 30719
rect 10793 30685 10827 30719
rect 8125 30617 8159 30651
rect 1225 30549 1259 30583
rect 1501 30549 1535 30583
rect 2605 30549 2639 30583
rect 2973 30549 3007 30583
rect 3341 30549 3375 30583
rect 6193 30549 6227 30583
rect 6929 30549 6963 30583
rect 7665 30549 7699 30583
rect 9229 30549 9263 30583
rect 1501 30345 1535 30379
rect 2973 30345 3007 30379
rect 3985 30345 4019 30379
rect 4997 30345 5031 30379
rect 5181 30345 5215 30379
rect 5917 30345 5951 30379
rect 6193 30345 6227 30379
rect 9689 30345 9723 30379
rect 10425 30345 10459 30379
rect 3341 30277 3375 30311
rect 4169 30277 4203 30311
rect 1961 30141 1995 30175
rect 2237 30141 2271 30175
rect 2789 30141 2823 30175
rect 2881 30141 2915 30175
rect 3065 30141 3099 30175
rect 3249 30141 3283 30175
rect 3433 30141 3467 30175
rect 3617 30141 3651 30175
rect 4353 30141 4387 30175
rect 4537 30141 4571 30175
rect 4629 30141 4663 30175
rect 4905 30141 4939 30175
rect 5825 30141 5859 30175
rect 6009 30141 6043 30175
rect 6101 30141 6135 30175
rect 6469 30141 6503 30175
rect 6745 30141 6779 30175
rect 6929 30141 6963 30175
rect 7021 30141 7055 30175
rect 7113 30141 7147 30175
rect 7849 30141 7883 30175
rect 7941 30141 7975 30175
rect 8033 30141 8067 30175
rect 8217 30141 8251 30175
rect 1225 30073 1259 30107
rect 1685 30073 1719 30107
rect 3985 30073 4019 30107
rect 5365 30073 5399 30107
rect 8401 30073 8435 30107
rect 10609 30073 10643 30107
rect 4445 30005 4479 30039
rect 5457 30005 5491 30039
rect 6653 30005 6687 30039
rect 7389 30005 7423 30039
rect 7573 30005 7607 30039
rect 10241 30005 10275 30039
rect 10409 30005 10443 30039
rect 3157 29801 3191 29835
rect 4261 29801 4295 29835
rect 4905 29801 4939 29835
rect 5825 29801 5859 29835
rect 7297 29801 7331 29835
rect 8033 29801 8067 29835
rect 8953 29801 8987 29835
rect 949 29733 983 29767
rect 2789 29733 2823 29767
rect 3433 29733 3467 29767
rect 3525 29733 3559 29767
rect 6009 29733 6043 29767
rect 10088 29733 10122 29767
rect 1685 29665 1719 29699
rect 1777 29665 1811 29699
rect 1869 29665 1903 29699
rect 2053 29665 2087 29699
rect 2421 29665 2455 29699
rect 2697 29665 2731 29699
rect 2881 29665 2915 29699
rect 3893 29665 3927 29699
rect 4997 29665 5031 29699
rect 5641 29665 5675 29699
rect 6193 29665 6227 29699
rect 6285 29665 6319 29699
rect 6469 29665 6503 29699
rect 6653 29665 6687 29699
rect 7021 29665 7055 29699
rect 7481 29665 7515 29699
rect 7573 29665 7607 29699
rect 7849 29665 7883 29699
rect 8585 29665 8619 29699
rect 8769 29665 8803 29699
rect 8861 29665 8895 29699
rect 10425 29665 10459 29699
rect 10518 29665 10552 29699
rect 1225 29597 1259 29631
rect 2145 29597 2179 29631
rect 4721 29597 4755 29631
rect 7757 29597 7791 29631
rect 8309 29597 8343 29631
rect 10333 29597 10367 29631
rect 1133 29529 1167 29563
rect 2053 29529 2087 29563
rect 2237 29461 2271 29495
rect 2605 29461 2639 29495
rect 4445 29461 4479 29495
rect 5365 29461 5399 29495
rect 5549 29461 5583 29495
rect 6285 29461 6319 29495
rect 7021 29461 7055 29495
rect 7205 29461 7239 29495
rect 8493 29461 8527 29495
rect 10609 29461 10643 29495
rect 2329 29257 2363 29291
rect 6009 29257 6043 29291
rect 6745 29257 6779 29291
rect 6929 29257 6963 29291
rect 8217 29257 8251 29291
rect 9137 29257 9171 29291
rect 857 29189 891 29223
rect 4721 29189 4755 29223
rect 5089 29189 5123 29223
rect 8125 29189 8159 29223
rect 8677 29189 8711 29223
rect 8769 29189 8803 29223
rect 1777 29121 1811 29155
rect 2237 29121 2271 29155
rect 9413 29121 9447 29155
rect 1041 29053 1075 29087
rect 1133 29053 1167 29087
rect 2053 29053 2087 29087
rect 2513 29053 2547 29087
rect 2773 29053 2807 29087
rect 2873 29047 2907 29081
rect 3065 29053 3099 29087
rect 3801 29053 3835 29087
rect 5365 29053 5399 29087
rect 5825 29053 5859 29087
rect 6101 29053 6135 29087
rect 6377 29053 6411 29087
rect 6561 29053 6595 29087
rect 6837 29053 6871 29087
rect 7113 29053 7147 29087
rect 7297 29053 7331 29087
rect 7389 29053 7423 29087
rect 7849 29053 7883 29087
rect 8217 29053 8251 29087
rect 8493 29053 8527 29087
rect 857 28985 891 29019
rect 1225 28985 1259 29019
rect 3433 28985 3467 29019
rect 3709 28985 3743 29019
rect 4169 28985 4203 29019
rect 4537 28985 4571 29019
rect 5641 28985 5675 29019
rect 7757 28985 7791 29019
rect 7941 28985 7975 29019
rect 9658 28985 9692 29019
rect 2697 28917 2731 28951
rect 2881 28917 2915 28951
rect 4905 28917 4939 28951
rect 6285 28917 6319 28951
rect 6561 28917 6595 28951
rect 9137 28917 9171 28951
rect 9321 28917 9355 28951
rect 10793 28917 10827 28951
rect 1041 28713 1075 28747
rect 3433 28713 3467 28747
rect 4077 28713 4111 28747
rect 5181 28713 5215 28747
rect 6101 28713 6135 28747
rect 7665 28713 7699 28747
rect 8585 28713 8619 28747
rect 10083 28713 10117 28747
rect 1225 28645 1259 28679
rect 5365 28645 5399 28679
rect 7205 28645 7239 28679
rect 9413 28645 9447 28679
rect 9873 28645 9907 28679
rect 857 28577 891 28611
rect 1133 28577 1167 28611
rect 2053 28577 2087 28611
rect 2237 28577 2271 28611
rect 2329 28577 2363 28611
rect 2513 28577 2547 28611
rect 2605 28577 2639 28611
rect 2789 28577 2823 28611
rect 2881 28577 2915 28611
rect 2973 28577 3007 28611
rect 3617 28577 3651 28611
rect 3893 28577 3927 28611
rect 4169 28577 4203 28611
rect 4629 28577 4663 28611
rect 5089 28577 5123 28611
rect 5457 28577 5491 28611
rect 5641 28577 5675 28611
rect 6377 28577 6411 28611
rect 6469 28577 6503 28611
rect 6837 28577 6871 28611
rect 7573 28577 7607 28611
rect 7757 28577 7791 28611
rect 8125 28577 8159 28611
rect 8217 28577 8251 28611
rect 8401 28577 8435 28611
rect 8861 28577 8895 28611
rect 8953 28577 8987 28611
rect 9045 28577 9079 28611
rect 9229 28577 9263 28611
rect 10517 28577 10551 28611
rect 10701 28577 10735 28611
rect 1777 28509 1811 28543
rect 4721 28509 4755 28543
rect 4905 28509 4939 28543
rect 10333 28509 10367 28543
rect 3709 28441 3743 28475
rect 4261 28441 4295 28475
rect 8677 28441 8711 28475
rect 10241 28441 10275 28475
rect 857 28373 891 28407
rect 2421 28373 2455 28407
rect 3249 28373 3283 28407
rect 5365 28373 5399 28407
rect 5549 28373 5583 28407
rect 7389 28373 7423 28407
rect 7941 28373 7975 28407
rect 9505 28373 9539 28407
rect 10079 28373 10113 28407
rect 3249 28169 3283 28203
rect 3617 28169 3651 28203
rect 4169 28169 4203 28203
rect 857 28101 891 28135
rect 5917 28101 5951 28135
rect 8033 28101 8067 28135
rect 1225 28033 1259 28067
rect 2697 28033 2731 28067
rect 2789 28033 2823 28067
rect 3709 28033 3743 28067
rect 3801 28033 3835 28067
rect 8585 28033 8619 28067
rect 9229 28033 9263 28067
rect 9413 28033 9447 28067
rect 9505 28033 9539 28067
rect 9689 28033 9723 28067
rect 10149 28033 10183 28067
rect 10609 28033 10643 28067
rect 857 27965 891 27999
rect 1133 27965 1167 27999
rect 1409 27965 1443 27999
rect 1685 27965 1719 27999
rect 2329 27965 2363 27999
rect 2513 27965 2547 27999
rect 2881 27965 2915 27999
rect 3065 27965 3099 27999
rect 3433 27965 3467 27999
rect 3985 27965 4019 27999
rect 4261 27965 4295 27999
rect 4905 27965 4939 27999
rect 4997 27965 5031 27999
rect 6561 27965 6595 27999
rect 8217 27965 8251 27999
rect 9597 27965 9631 27999
rect 10241 27965 10275 27999
rect 2237 27897 2271 27931
rect 2973 27897 3007 27931
rect 5365 27897 5399 27931
rect 5733 27897 5767 27931
rect 6285 27897 6319 27931
rect 6653 27897 6687 27931
rect 7021 27897 7055 27931
rect 8677 27897 8711 27931
rect 1041 27829 1075 27863
rect 4629 27829 4663 27863
rect 7389 27829 7423 27863
rect 7573 27829 7607 27863
rect 8769 27829 8803 27863
rect 9137 27829 9171 27863
rect 2421 27625 2455 27659
rect 3249 27625 3283 27659
rect 5273 27625 5307 27659
rect 8033 27625 8067 27659
rect 1041 27557 1075 27591
rect 4160 27557 4194 27591
rect 6377 27557 6411 27591
rect 6745 27557 6779 27591
rect 7113 27557 7147 27591
rect 7481 27557 7515 27591
rect 8217 27557 8251 27591
rect 8309 27557 8343 27591
rect 1225 27489 1259 27523
rect 1869 27489 1903 27523
rect 2145 27489 2179 27523
rect 2605 27489 2639 27523
rect 2697 27489 2731 27523
rect 3617 27489 3651 27523
rect 3893 27489 3927 27523
rect 5549 27489 5583 27523
rect 5825 27489 5859 27523
rect 6653 27489 6687 27523
rect 7941 27489 7975 27523
rect 8493 27489 8527 27523
rect 8769 27489 8803 27523
rect 8953 27489 8987 27523
rect 9229 27489 9263 27523
rect 9485 27489 9519 27523
rect 1317 27421 1351 27455
rect 2329 27421 2363 27455
rect 2789 27421 2823 27455
rect 2881 27421 2915 27455
rect 3433 27421 3467 27455
rect 3525 27421 3559 27455
rect 3709 27421 3743 27455
rect 8677 27353 8711 27387
rect 857 27285 891 27319
rect 5457 27285 5491 27319
rect 5917 27285 5951 27319
rect 7665 27285 7699 27319
rect 8217 27285 8251 27319
rect 9137 27285 9171 27319
rect 10609 27285 10643 27319
rect 3893 27081 3927 27115
rect 7849 27081 7883 27115
rect 8493 27081 8527 27115
rect 6193 27013 6227 27047
rect 1685 26945 1719 26979
rect 2237 26945 2271 26979
rect 2605 26945 2639 26979
rect 2697 26945 2731 26979
rect 4261 26945 4295 26979
rect 8677 26945 8711 26979
rect 1133 26877 1167 26911
rect 1225 26877 1259 26911
rect 1409 26877 1443 26911
rect 2329 26877 2363 26911
rect 2513 26877 2547 26911
rect 2881 26877 2915 26911
rect 3617 26877 3651 26911
rect 4077 26877 4111 26911
rect 4353 26877 4387 26911
rect 4445 26877 4479 26911
rect 4629 26877 4663 26911
rect 5641 26877 5675 26911
rect 6561 26877 6595 26911
rect 6837 26877 6871 26911
rect 6929 26877 6963 26911
rect 7021 26877 7055 26911
rect 7205 26877 7239 26911
rect 8401 26877 8435 26911
rect 8769 26877 8803 26911
rect 8861 26877 8895 26911
rect 9045 26877 9079 26911
rect 9137 26877 9171 26911
rect 10793 26877 10827 26911
rect 4905 26809 4939 26843
rect 5181 26809 5215 26843
rect 5273 26809 5307 26843
rect 6009 26809 6043 26843
rect 7481 26809 7515 26843
rect 7665 26809 7699 26843
rect 7941 26809 7975 26843
rect 9321 26809 9355 26843
rect 10526 26809 10560 26843
rect 949 26741 983 26775
rect 3065 26741 3099 26775
rect 6469 26741 6503 26775
rect 6653 26741 6687 26775
rect 7297 26741 7331 26775
rect 8677 26741 8711 26775
rect 9413 26741 9447 26775
rect 1041 26537 1075 26571
rect 2053 26537 2087 26571
rect 8217 26537 8251 26571
rect 3065 26469 3099 26503
rect 7021 26469 7055 26503
rect 857 26401 891 26435
rect 1041 26401 1075 26435
rect 1409 26401 1443 26435
rect 1685 26401 1719 26435
rect 1961 26401 1995 26435
rect 2237 26401 2271 26435
rect 2513 26401 2547 26435
rect 2697 26401 2731 26435
rect 3249 26401 3283 26435
rect 5089 26401 5123 26435
rect 5365 26401 5399 26435
rect 5825 26401 5859 26435
rect 6469 26401 6503 26435
rect 6561 26401 6595 26435
rect 6653 26401 6687 26435
rect 7205 26401 7239 26435
rect 7481 26401 7515 26435
rect 7665 26401 7699 26435
rect 7757 26401 7791 26435
rect 8033 26401 8067 26435
rect 8585 26401 8619 26435
rect 9321 26401 9355 26435
rect 9505 26401 9539 26435
rect 9873 26401 9907 26435
rect 10517 26401 10551 26435
rect 5641 26333 5675 26367
rect 6377 26333 6411 26367
rect 7849 26333 7883 26367
rect 9413 26333 9447 26367
rect 9781 26333 9815 26367
rect 10333 26333 10367 26367
rect 1869 26265 1903 26299
rect 5181 26265 5215 26299
rect 6009 26265 6043 26299
rect 10241 26265 10275 26299
rect 1225 26197 1259 26231
rect 1501 26197 1535 26231
rect 3617 26197 3651 26231
rect 5549 26197 5583 26231
rect 6193 26197 6227 26231
rect 6837 26197 6871 26231
rect 10701 26197 10735 26231
rect 949 25993 983 26027
rect 2973 25993 3007 26027
rect 4721 25993 4755 26027
rect 5549 25993 5583 26027
rect 9781 25993 9815 26027
rect 3249 25925 3283 25959
rect 5641 25925 5675 25959
rect 1225 25857 1259 25891
rect 1777 25857 1811 25891
rect 4077 25857 4111 25891
rect 5089 25857 5123 25891
rect 5181 25857 5215 25891
rect 7665 25857 7699 25891
rect 1133 25789 1167 25823
rect 2053 25789 2087 25823
rect 2237 25789 2271 25823
rect 2421 25789 2455 25823
rect 2513 25789 2547 25823
rect 2624 25789 2658 25823
rect 2789 25789 2823 25823
rect 3425 25767 3459 25801
rect 3525 25789 3559 25823
rect 3709 25789 3743 25823
rect 3801 25789 3835 25823
rect 4813 25789 4847 25823
rect 4997 25789 5031 25823
rect 5365 25789 5399 25823
rect 5825 25789 5859 25823
rect 6101 25789 6135 25823
rect 6193 25789 6227 25823
rect 6837 25789 6871 25823
rect 6929 25789 6963 25823
rect 7021 25789 7055 25823
rect 7205 25789 7239 25823
rect 7297 25779 7331 25813
rect 7481 25789 7515 25823
rect 7573 25789 7607 25823
rect 7849 25789 7883 25823
rect 8493 25789 8527 25823
rect 10517 25789 10551 25823
rect 10701 25789 10735 25823
rect 4261 25721 4295 25755
rect 6009 25721 6043 25755
rect 4353 25653 4387 25687
rect 6377 25653 6411 25687
rect 6561 25653 6595 25687
rect 8033 25653 8067 25687
rect 10333 25653 10367 25687
rect 1133 25449 1167 25483
rect 3341 25449 3375 25483
rect 4629 25449 4663 25483
rect 4813 25449 4847 25483
rect 6469 25449 6503 25483
rect 8585 25449 8619 25483
rect 8953 25449 8987 25483
rect 3157 25381 3191 25415
rect 3617 25381 3651 25415
rect 4445 25381 4479 25415
rect 9597 25381 9631 25415
rect 857 25313 891 25347
rect 1777 25313 1811 25347
rect 2053 25313 2087 25347
rect 2237 25313 2271 25347
rect 2513 25313 2547 25347
rect 3065 25313 3099 25347
rect 3433 25313 3467 25347
rect 3801 25313 3835 25347
rect 3985 25313 4019 25347
rect 4165 25315 4199 25349
rect 4333 25313 4367 25347
rect 4705 25319 4739 25353
rect 5089 25313 5123 25347
rect 5365 25313 5399 25347
rect 6009 25313 6043 25347
rect 6285 25313 6319 25347
rect 6653 25313 6687 25347
rect 6837 25313 6871 25347
rect 6929 25313 6963 25347
rect 7021 25313 7055 25347
rect 7205 25313 7239 25347
rect 7481 25313 7515 25347
rect 7757 25313 7791 25347
rect 7849 25313 7883 25347
rect 8033 25313 8067 25347
rect 8493 25313 8527 25347
rect 9137 25313 9171 25347
rect 9229 25313 9263 25347
rect 1133 25245 1167 25279
rect 1225 25245 1259 25279
rect 2697 25245 2731 25279
rect 2789 25245 2823 25279
rect 3249 25245 3283 25279
rect 4077 25245 4111 25279
rect 4813 25245 4847 25279
rect 5641 25245 5675 25279
rect 7665 25245 7699 25279
rect 8677 25245 8711 25279
rect 9505 25245 9539 25279
rect 10149 25245 10183 25279
rect 949 25177 983 25211
rect 5181 25177 5215 25211
rect 5549 25177 5583 25211
rect 6193 25177 6227 25211
rect 7297 25177 7331 25211
rect 2329 25109 2363 25143
rect 4445 25109 4479 25143
rect 4997 25109 5031 25143
rect 5825 25109 5859 25143
rect 8125 25109 8159 25143
rect 10793 25109 10827 25143
rect 3249 24905 3283 24939
rect 4077 24905 4111 24939
rect 8217 24905 8251 24939
rect 1961 24837 1995 24871
rect 7849 24837 7883 24871
rect 1501 24769 1535 24803
rect 1685 24769 1719 24803
rect 3525 24769 3559 24803
rect 8769 24769 8803 24803
rect 10333 24769 10367 24803
rect 1777 24701 1811 24735
rect 2145 24701 2179 24735
rect 2421 24701 2455 24735
rect 2605 24701 2639 24735
rect 2697 24701 2731 24735
rect 3249 24701 3283 24735
rect 3433 24701 3467 24735
rect 3709 24701 3743 24735
rect 4261 24701 4295 24735
rect 4721 24701 4755 24735
rect 4813 24701 4847 24735
rect 4997 24701 5031 24735
rect 5181 24701 5215 24735
rect 5917 24701 5951 24735
rect 6009 24701 6043 24735
rect 6837 24701 6871 24735
rect 7113 24701 7147 24735
rect 7205 24701 7239 24735
rect 7389 24701 7423 24735
rect 7481 24701 7515 24735
rect 7573 24701 7607 24735
rect 7941 24701 7975 24735
rect 8033 24701 8067 24735
rect 8217 24701 8251 24735
rect 10057 24701 10091 24735
rect 10609 24701 10643 24735
rect 10793 24701 10827 24735
rect 2881 24633 2915 24667
rect 3893 24633 3927 24667
rect 4537 24633 4571 24667
rect 5273 24633 5307 24667
rect 5457 24633 5491 24667
rect 8401 24633 8435 24667
rect 8585 24633 8619 24667
rect 9045 24633 9079 24667
rect 9229 24633 9263 24667
rect 1317 24565 1351 24599
rect 2329 24565 2363 24599
rect 5089 24565 5123 24599
rect 5641 24565 5675 24599
rect 6193 24565 6227 24599
rect 8861 24565 8895 24599
rect 9413 24565 9447 24599
rect 10701 24565 10735 24599
rect 6285 24361 6319 24395
rect 6929 24361 6963 24395
rect 7849 24361 7883 24395
rect 9321 24361 9355 24395
rect 10149 24361 10183 24395
rect 10701 24361 10735 24395
rect 1225 24293 1259 24327
rect 3985 24293 4019 24327
rect 4169 24293 4203 24327
rect 4629 24293 4663 24327
rect 5273 24293 5307 24327
rect 5365 24293 5399 24327
rect 5483 24293 5517 24327
rect 8953 24293 8987 24327
rect 9045 24293 9079 24327
rect 1777 24225 1811 24259
rect 2053 24225 2087 24259
rect 2329 24225 2363 24259
rect 2513 24225 2547 24259
rect 2881 24225 2915 24259
rect 3065 24225 3099 24259
rect 4813 24225 4847 24259
rect 5181 24225 5215 24259
rect 6193 24225 6227 24259
rect 6837 24225 6871 24259
rect 7205 24225 7239 24259
rect 7389 24225 7423 24259
rect 7481 24225 7515 24259
rect 7665 24225 7699 24259
rect 7757 24225 7791 24259
rect 8033 24225 8067 24259
rect 8309 24225 8343 24259
rect 8677 24225 8711 24259
rect 8769 24225 8803 24259
rect 9169 24225 9203 24259
rect 10241 24225 10275 24259
rect 10609 24225 10643 24259
rect 10793 24225 10827 24259
rect 2237 24157 2271 24191
rect 2789 24157 2823 24191
rect 3157 24157 3191 24191
rect 3433 24157 3467 24191
rect 3617 24157 3651 24191
rect 3709 24157 3743 24191
rect 5641 24157 5675 24191
rect 6377 24157 6411 24191
rect 8217 24157 8251 24191
rect 9689 24157 9723 24191
rect 9781 24157 9815 24191
rect 3065 24089 3099 24123
rect 4353 24089 4387 24123
rect 5825 24089 5859 24123
rect 8493 24089 8527 24123
rect 2697 24021 2731 24055
rect 4445 24021 4479 24055
rect 4997 24021 5031 24055
rect 9505 24021 9539 24055
rect 10425 24021 10459 24055
rect 4169 23817 4203 23851
rect 5089 23817 5123 23851
rect 7573 23817 7607 23851
rect 8401 23817 8435 23851
rect 10333 23817 10367 23851
rect 10609 23817 10643 23851
rect 2697 23749 2731 23783
rect 4721 23749 4755 23783
rect 1777 23681 1811 23715
rect 2329 23681 2363 23715
rect 3249 23681 3283 23715
rect 6469 23681 6503 23715
rect 6837 23681 6871 23715
rect 6929 23681 6963 23715
rect 7757 23681 7791 23715
rect 9413 23681 9447 23715
rect 2053 23613 2087 23647
rect 2237 23613 2271 23647
rect 2513 23613 2547 23647
rect 2789 23613 2823 23647
rect 3433 23613 3467 23647
rect 3617 23613 3651 23647
rect 3709 23613 3743 23647
rect 4077 23613 4111 23647
rect 4353 23613 4387 23647
rect 4629 23613 4663 23647
rect 4905 23613 4939 23647
rect 5181 23613 5215 23647
rect 5273 23613 5307 23647
rect 5457 23613 5491 23647
rect 6173 23613 6207 23647
rect 6377 23613 6411 23647
rect 6653 23613 6687 23647
rect 6745 23613 6779 23647
rect 7297 23613 7331 23647
rect 7389 23613 7423 23647
rect 7647 23613 7681 23647
rect 8585 23613 8619 23647
rect 8677 23613 8711 23647
rect 8953 23613 8987 23647
rect 9045 23613 9079 23647
rect 9137 23613 9171 23647
rect 9229 23613 9263 23647
rect 9505 23613 9539 23647
rect 9873 23613 9907 23647
rect 10057 23613 10091 23647
rect 10241 23613 10275 23647
rect 10425 23613 10459 23647
rect 10517 23613 10551 23647
rect 10701 23613 10735 23647
rect 1225 23545 1259 23579
rect 4537 23545 4571 23579
rect 5365 23545 5399 23579
rect 6091 23545 6125 23579
rect 6285 23545 6319 23579
rect 7113 23545 7147 23579
rect 7941 23545 7975 23579
rect 8769 23545 8803 23579
rect 9413 23545 9447 23579
rect 3985 23477 4019 23511
rect 9689 23477 9723 23511
rect 9873 23477 9907 23511
rect 1317 23273 1351 23307
rect 5089 23273 5123 23307
rect 9137 23273 9171 23307
rect 9229 23273 9263 23307
rect 10333 23273 10367 23307
rect 2789 23205 2823 23239
rect 7573 23205 7607 23239
rect 8217 23205 8251 23239
rect 1133 23137 1167 23171
rect 1501 23137 1535 23171
rect 1961 23137 1995 23171
rect 2145 23137 2179 23171
rect 2237 23137 2271 23171
rect 2329 23137 2363 23171
rect 2421 23137 2455 23171
rect 2605 23137 2639 23171
rect 3433 23137 3467 23171
rect 3801 23137 3835 23171
rect 3893 23137 3927 23171
rect 4261 23137 4295 23171
rect 4721 23137 4755 23171
rect 5273 23137 5307 23171
rect 5825 23137 5859 23171
rect 5917 23137 5951 23171
rect 6101 23137 6135 23171
rect 6193 23137 6227 23171
rect 6285 23137 6319 23171
rect 6561 23137 6595 23171
rect 6745 23137 6779 23171
rect 6837 23137 6871 23171
rect 7021 23137 7055 23171
rect 7113 23137 7147 23171
rect 7389 23137 7423 23171
rect 7941 23137 7975 23171
rect 8493 23137 8527 23171
rect 8677 23137 8711 23171
rect 8769 23137 8803 23171
rect 8861 23137 8895 23171
rect 9597 23137 9631 23171
rect 10149 23137 10183 23171
rect 1685 23069 1719 23103
rect 4813 23069 4847 23103
rect 5549 23069 5583 23103
rect 7205 23069 7239 23103
rect 9505 23069 9539 23103
rect 9873 23069 9907 23103
rect 8033 23001 8067 23035
rect 9965 23001 9999 23035
rect 949 22933 983 22967
rect 1777 22933 1811 22967
rect 4077 22933 4111 22967
rect 5457 22933 5491 22967
rect 6469 22933 6503 22967
rect 6653 22933 6687 22967
rect 7757 22933 7791 22967
rect 949 22729 983 22763
rect 2053 22729 2087 22763
rect 2237 22729 2271 22763
rect 3617 22729 3651 22763
rect 4353 22729 4387 22763
rect 4813 22729 4847 22763
rect 5917 22729 5951 22763
rect 6377 22729 6411 22763
rect 6837 22729 6871 22763
rect 7665 22729 7699 22763
rect 9597 22729 9631 22763
rect 5181 22661 5215 22695
rect 8677 22661 8711 22695
rect 10241 22661 10275 22695
rect 1225 22593 1259 22627
rect 7481 22593 7515 22627
rect 8033 22593 8067 22627
rect 10057 22593 10091 22627
rect 10517 22593 10551 22627
rect 1133 22525 1167 22559
rect 1685 22525 1719 22559
rect 1777 22525 1811 22559
rect 1869 22525 1903 22559
rect 2421 22525 2455 22559
rect 2697 22525 2731 22559
rect 3065 22525 3099 22559
rect 3249 22525 3283 22559
rect 4169 22525 4203 22559
rect 4997 22525 5031 22559
rect 5181 22525 5215 22559
rect 5365 22525 5399 22559
rect 6101 22525 6135 22559
rect 6561 22525 6595 22559
rect 7849 22525 7883 22559
rect 8125 22525 8159 22559
rect 8401 22525 8435 22559
rect 8585 22525 8619 22559
rect 8953 22525 8987 22559
rect 9045 22525 9079 22559
rect 9137 22525 9171 22559
rect 9321 22525 9355 22559
rect 9965 22525 9999 22559
rect 10609 22525 10643 22559
rect 3985 22457 4019 22491
rect 4445 22457 4479 22491
rect 4629 22457 4663 22491
rect 6285 22457 6319 22491
rect 6745 22457 6779 22491
rect 7297 22457 7331 22491
rect 2605 22389 2639 22423
rect 2881 22389 2915 22423
rect 3617 22389 3651 22423
rect 3801 22389 3835 22423
rect 5549 22389 5583 22423
rect 7205 22389 7239 22423
rect 8493 22389 8527 22423
rect 2329 22185 2363 22219
rect 2881 22185 2915 22219
rect 4445 22185 4479 22219
rect 5181 22185 5215 22219
rect 5641 22185 5675 22219
rect 8125 22185 8159 22219
rect 10425 22185 10459 22219
rect 4813 22117 4847 22151
rect 7573 22117 7607 22151
rect 8401 22117 8435 22151
rect 8493 22117 8527 22151
rect 1777 22049 1811 22083
rect 2053 22049 2087 22083
rect 2513 22049 2547 22083
rect 2697 22049 2731 22083
rect 2789 22049 2823 22083
rect 3065 22049 3099 22083
rect 3157 22049 3191 22083
rect 3433 22049 3467 22083
rect 3709 22049 3743 22083
rect 3801 22049 3835 22083
rect 3893 22049 3927 22083
rect 4261 22049 4295 22083
rect 4537 22049 4571 22083
rect 4997 22049 5031 22083
rect 5089 22049 5123 22083
rect 5273 22049 5307 22083
rect 5365 22049 5399 22083
rect 7665 22049 7699 22083
rect 8309 22049 8343 22083
rect 8677 22049 8711 22083
rect 8769 22071 8803 22105
rect 8953 22049 8987 22083
rect 9137 22049 9171 22083
rect 9689 22049 9723 22083
rect 9965 22049 9999 22083
rect 10149 22049 10183 22083
rect 10425 22049 10459 22083
rect 10609 22049 10643 22083
rect 1225 21981 1259 22015
rect 2237 21981 2271 22015
rect 3525 21981 3559 22015
rect 3985 21981 4019 22015
rect 5457 21981 5491 22015
rect 5641 21981 5675 22015
rect 8861 21981 8895 22015
rect 9413 21981 9447 22015
rect 10333 21981 10367 22015
rect 6285 21913 6319 21947
rect 3341 21845 3375 21879
rect 4629 21845 4663 21879
rect 7849 21845 7883 21879
rect 9321 21845 9355 21879
rect 9505 21845 9539 21879
rect 9873 21845 9907 21879
rect 1041 21641 1075 21675
rect 1501 21641 1535 21675
rect 3341 21641 3375 21675
rect 4537 21641 4571 21675
rect 6377 21641 6411 21675
rect 8861 21641 8895 21675
rect 9873 21641 9907 21675
rect 3617 21573 3651 21607
rect 5733 21573 5767 21607
rect 6193 21573 6227 21607
rect 7021 21573 7055 21607
rect 9597 21573 9631 21607
rect 5273 21505 5307 21539
rect 5457 21505 5491 21539
rect 6561 21505 6595 21539
rect 6745 21505 6779 21539
rect 6837 21505 6871 21539
rect 7665 21505 7699 21539
rect 1225 21437 1259 21471
rect 1409 21437 1443 21471
rect 1685 21437 1719 21471
rect 1869 21437 1903 21471
rect 1961 21437 1995 21471
rect 2605 21437 2639 21471
rect 2789 21437 2823 21471
rect 3065 21437 3099 21471
rect 3249 21437 3283 21471
rect 3433 21437 3467 21471
rect 3617 21437 3651 21471
rect 4261 21437 4295 21471
rect 5918 21437 5952 21471
rect 6009 21437 6043 21471
rect 6285 21437 6319 21471
rect 6653 21437 6687 21471
rect 7389 21437 7423 21471
rect 8217 21437 8251 21471
rect 8401 21437 8435 21471
rect 9234 21437 9268 21471
rect 9413 21437 9447 21471
rect 9781 21437 9815 21471
rect 9965 21437 9999 21471
rect 2421 21369 2455 21403
rect 2973 21369 3007 21403
rect 4721 21369 4755 21403
rect 8033 21369 8067 21403
rect 8861 21369 8895 21403
rect 9045 21369 9079 21403
rect 9137 21369 9171 21403
rect 2145 21301 2179 21335
rect 4353 21301 4387 21335
rect 4521 21301 4555 21335
rect 4813 21301 4847 21335
rect 5181 21301 5215 21335
rect 7481 21301 7515 21335
rect 7849 21301 7883 21335
rect 8585 21301 8619 21335
rect 1317 21097 1351 21131
rect 1869 21097 1903 21131
rect 7113 21097 7147 21131
rect 10149 21097 10183 21131
rect 3341 21029 3375 21063
rect 4813 21029 4847 21063
rect 4997 21029 5031 21063
rect 5825 21029 5859 21063
rect 1501 20961 1535 20995
rect 1685 20961 1719 20995
rect 1777 20961 1811 20995
rect 2053 20961 2087 20995
rect 2329 20961 2363 20995
rect 2605 20961 2639 20995
rect 2789 20961 2823 20995
rect 3157 20961 3191 20995
rect 3617 20961 3651 20995
rect 3709 20961 3743 20995
rect 3893 20961 3927 20995
rect 4077 20961 4111 20995
rect 4169 20961 4203 20995
rect 4353 20961 4387 20995
rect 5089 20961 5123 20995
rect 5273 20961 5307 20995
rect 5641 20961 5675 20995
rect 6009 20961 6043 20995
rect 6193 20961 6227 20995
rect 6285 20961 6319 20995
rect 6469 20961 6503 20995
rect 6561 20961 6595 20995
rect 6837 20961 6871 20995
rect 7297 20961 7331 20995
rect 7481 20961 7515 20995
rect 7665 20961 7699 20995
rect 7849 20961 7883 20995
rect 9229 20961 9263 20995
rect 9505 20961 9539 20995
rect 9965 20961 9999 20995
rect 10241 20961 10275 20995
rect 2881 20893 2915 20927
rect 2973 20893 3007 20927
rect 5365 20893 5399 20927
rect 6653 20893 6687 20927
rect 7573 20893 7607 20927
rect 8861 20893 8895 20927
rect 8953 20893 8987 20927
rect 9597 20893 9631 20927
rect 9689 20893 9723 20927
rect 9781 20893 9815 20927
rect 2237 20825 2271 20859
rect 3801 20825 3835 20859
rect 5273 20825 5307 20859
rect 5457 20825 5491 20859
rect 8769 20825 8803 20859
rect 2421 20757 2455 20791
rect 3433 20757 3467 20791
rect 4537 20757 4571 20791
rect 4629 20757 4663 20791
rect 5549 20757 5583 20791
rect 7021 20757 7055 20791
rect 9137 20757 9171 20791
rect 9321 20757 9355 20791
rect 9965 20757 9999 20791
rect 2697 20553 2731 20587
rect 5457 20553 5491 20587
rect 5549 20553 5583 20587
rect 7481 20553 7515 20587
rect 7665 20553 7699 20587
rect 9413 20553 9447 20587
rect 3249 20485 3283 20519
rect 4169 20485 4203 20519
rect 1225 20417 1259 20451
rect 1777 20417 1811 20451
rect 4629 20417 4663 20451
rect 5365 20417 5399 20451
rect 6469 20417 6503 20451
rect 6837 20417 6871 20451
rect 7849 20417 7883 20451
rect 9045 20417 9079 20451
rect 9689 20417 9723 20451
rect 10333 20417 10367 20451
rect 2053 20349 2087 20383
rect 2237 20349 2271 20383
rect 2513 20349 2547 20383
rect 2789 20349 2823 20383
rect 3433 20349 3467 20383
rect 3709 20349 3743 20383
rect 4077 20349 4111 20383
rect 4353 20349 4387 20383
rect 4445 20349 4479 20383
rect 4905 20349 4939 20383
rect 4997 20349 5031 20383
rect 5089 20349 5123 20383
rect 5181 20349 5215 20383
rect 5641 20349 5675 20383
rect 6193 20349 6227 20383
rect 7665 20349 7699 20383
rect 8493 20349 8527 20383
rect 8953 20349 8987 20383
rect 9137 20349 9171 20383
rect 9781 20349 9815 20383
rect 10425 20349 10459 20383
rect 3617 20281 3651 20315
rect 6285 20281 6319 20315
rect 6929 20281 6963 20315
rect 7941 20281 7975 20315
rect 2329 20213 2363 20247
rect 4721 20213 4755 20247
rect 5825 20213 5859 20247
rect 7021 20213 7055 20247
rect 7389 20213 7423 20247
rect 8585 20213 8619 20247
rect 10057 20213 10091 20247
rect 2605 20009 2639 20043
rect 3157 20009 3191 20043
rect 3525 20009 3559 20043
rect 4813 20009 4847 20043
rect 5273 20009 5307 20043
rect 4629 19941 4663 19975
rect 6561 19941 6595 19975
rect 7757 19941 7791 19975
rect 9689 19941 9723 19975
rect 1777 19873 1811 19907
rect 2053 19873 2087 19907
rect 2789 19873 2823 19907
rect 3341 19873 3375 19907
rect 3617 19873 3651 19907
rect 3893 19873 3927 19907
rect 4169 19873 4203 19907
rect 4261 19873 4295 19907
rect 4445 19873 4479 19907
rect 4537 19873 4571 19907
rect 4721 19873 4755 19907
rect 5181 19873 5215 19907
rect 6285 19873 6319 19907
rect 6377 19873 6411 19907
rect 6745 19873 6779 19907
rect 7113 19873 7147 19907
rect 7297 19873 7331 19907
rect 8217 19873 8251 19907
rect 8401 19873 8435 19907
rect 8953 19873 8987 19907
rect 9137 19873 9171 19907
rect 1225 19805 1259 19839
rect 2237 19805 2271 19839
rect 3065 19805 3099 19839
rect 4077 19805 4111 19839
rect 5457 19805 5491 19839
rect 6101 19805 6135 19839
rect 6193 19805 6227 19839
rect 6929 19805 6963 19839
rect 7021 19805 7055 19839
rect 7849 19805 7883 19839
rect 8033 19805 8067 19839
rect 8585 19805 8619 19839
rect 8677 19805 8711 19839
rect 2973 19737 3007 19771
rect 3709 19737 3743 19771
rect 7389 19737 7423 19771
rect 9965 19737 9999 19771
rect 5917 19669 5951 19703
rect 8953 19669 8987 19703
rect 10149 19669 10183 19703
rect 2329 19465 2363 19499
rect 3985 19465 4019 19499
rect 6745 19465 6779 19499
rect 7665 19465 7699 19499
rect 8677 19465 8711 19499
rect 10241 19465 10275 19499
rect 3617 19397 3651 19431
rect 6285 19397 6319 19431
rect 1225 19329 1259 19363
rect 2789 19329 2823 19363
rect 3249 19329 3283 19363
rect 5089 19329 5123 19363
rect 5181 19329 5215 19363
rect 5457 19329 5491 19363
rect 5825 19329 5859 19363
rect 7205 19329 7239 19363
rect 10333 19329 10367 19363
rect 1041 19261 1075 19295
rect 1133 19261 1167 19295
rect 1777 19261 1811 19295
rect 2053 19261 2087 19295
rect 2237 19261 2271 19295
rect 2513 19261 2547 19295
rect 2697 19261 2731 19295
rect 3433 19261 3467 19295
rect 3525 19261 3559 19295
rect 3801 19261 3835 19295
rect 4077 19261 4111 19295
rect 4813 19261 4847 19295
rect 4997 19261 5031 19295
rect 5273 19261 5307 19295
rect 5641 19261 5675 19295
rect 5733 19261 5767 19295
rect 6009 19261 6043 19295
rect 6101 19261 6135 19295
rect 6469 19261 6503 19295
rect 6561 19261 6595 19295
rect 6837 19261 6871 19295
rect 6929 19261 6963 19295
rect 7113 19261 7147 19295
rect 7297 19261 7331 19295
rect 7481 19261 7515 19295
rect 8033 19261 8067 19295
rect 8861 19261 8895 19295
rect 8953 19261 8987 19295
rect 9137 19261 9171 19295
rect 9229 19261 9263 19295
rect 9505 19261 9539 19295
rect 9781 19261 9815 19295
rect 9977 19261 10011 19295
rect 10609 19261 10643 19295
rect 857 19193 891 19227
rect 4353 19193 4387 19227
rect 4537 19193 4571 19227
rect 5825 19193 5859 19227
rect 955 19125 989 19159
rect 3249 19125 3283 19159
rect 4169 19125 4203 19159
rect 5457 19125 5491 19159
rect 7849 19125 7883 19159
rect 9321 19125 9355 19159
rect 10057 19125 10091 19159
rect 3249 18921 3283 18955
rect 4077 18921 4111 18955
rect 6929 18921 6963 18955
rect 8401 18921 8435 18955
rect 10333 18921 10367 18955
rect 10609 18921 10643 18955
rect 857 18853 891 18887
rect 4997 18853 5031 18887
rect 6837 18853 6871 18887
rect 7297 18853 7331 18887
rect 9413 18853 9447 18887
rect 10701 18853 10735 18887
rect 1041 18785 1075 18819
rect 1133 18785 1167 18819
rect 1225 18785 1259 18819
rect 1777 18785 1811 18819
rect 2053 18785 2087 18819
rect 2329 18785 2363 18819
rect 2513 18785 2547 18819
rect 2697 18785 2731 18819
rect 3065 18785 3099 18819
rect 3341 18785 3375 18819
rect 3709 18785 3743 18819
rect 3893 18785 3927 18819
rect 4169 18785 4203 18819
rect 4353 18785 4387 18819
rect 4905 18785 4939 18819
rect 5273 18785 5307 18819
rect 6101 18785 6135 18819
rect 6193 18785 6227 18819
rect 6469 18785 6503 18819
rect 6653 18785 6687 18819
rect 7113 18785 7147 18819
rect 8033 18785 8067 18819
rect 8953 18785 8987 18819
rect 9965 18785 9999 18819
rect 10149 18785 10183 18819
rect 10425 18785 10459 18819
rect 2237 18717 2271 18751
rect 2789 18717 2823 18751
rect 4997 18717 5031 18751
rect 5917 18717 5951 18751
rect 7941 18717 7975 18751
rect 9045 18717 9079 18751
rect 9321 18717 9355 18751
rect 9873 18717 9907 18751
rect 4537 18649 4571 18683
rect 4721 18649 4755 18683
rect 5181 18649 5215 18683
rect 9689 18649 9723 18683
rect 857 18581 891 18615
rect 2881 18581 2915 18615
rect 6009 18581 6043 18615
rect 2053 18377 2087 18411
rect 5549 18377 5583 18411
rect 5825 18377 5859 18411
rect 1409 18309 1443 18343
rect 3893 18309 3927 18343
rect 5457 18309 5491 18343
rect 9045 18309 9079 18343
rect 2145 18241 2179 18275
rect 2329 18241 2363 18275
rect 2421 18241 2455 18275
rect 3801 18241 3835 18275
rect 4353 18241 4387 18275
rect 5549 18241 5583 18275
rect 5733 18241 5767 18275
rect 7757 18241 7791 18275
rect 8677 18241 8711 18275
rect 10333 18241 10367 18275
rect 1225 18173 1259 18207
rect 1501 18173 1535 18207
rect 1593 18173 1627 18207
rect 1685 18173 1719 18207
rect 1869 18173 1903 18207
rect 3249 18173 3283 18207
rect 3341 18173 3375 18207
rect 3525 18173 3559 18207
rect 3617 18173 3651 18207
rect 4077 18173 4111 18207
rect 4261 18173 4295 18207
rect 4445 18173 4479 18207
rect 4629 18151 4663 18185
rect 4905 18173 4939 18207
rect 5365 18173 5399 18207
rect 6081 18173 6115 18207
rect 6193 18173 6227 18207
rect 6285 18173 6319 18207
rect 6469 18173 6503 18207
rect 7297 18173 7331 18207
rect 7481 18173 7515 18207
rect 7573 18173 7607 18207
rect 7665 18173 7699 18207
rect 7849 18173 7883 18207
rect 9321 18173 9355 18207
rect 9505 18173 9539 18207
rect 2789 18105 2823 18139
rect 4721 18105 4755 18139
rect 6653 18105 6687 18139
rect 1041 18037 1075 18071
rect 5089 18037 5123 18071
rect 6929 18037 6963 18071
rect 7113 18037 7147 18071
rect 9137 18037 9171 18071
rect 3709 17833 3743 17867
rect 5825 17833 5859 17867
rect 8033 17833 8067 17867
rect 8401 17765 8435 17799
rect 9045 17765 9079 17799
rect 1317 17697 1351 17731
rect 1593 17697 1627 17731
rect 1869 17697 1903 17731
rect 2145 17697 2179 17731
rect 2329 17697 2363 17731
rect 2605 17697 2639 17731
rect 2881 17697 2915 17731
rect 3065 17697 3099 17731
rect 3341 17697 3375 17731
rect 3525 17697 3559 17731
rect 3617 17697 3651 17731
rect 3893 17697 3927 17731
rect 4445 17697 4479 17731
rect 4629 17697 4663 17731
rect 4813 17697 4847 17731
rect 4997 17697 5031 17731
rect 5089 17697 5123 17731
rect 5273 17697 5307 17731
rect 5365 17697 5399 17731
rect 5641 17697 5675 17731
rect 6009 17697 6043 17731
rect 6101 17697 6135 17731
rect 6377 17697 6411 17731
rect 6469 17695 6503 17729
rect 6653 17697 6687 17731
rect 7021 17697 7055 17731
rect 7205 17697 7239 17731
rect 7297 17697 7331 17731
rect 7481 17697 7515 17731
rect 7576 17697 7610 17731
rect 7665 17697 7699 17731
rect 7849 17697 7883 17731
rect 8309 17697 8343 17731
rect 8493 17697 8527 17731
rect 8677 17697 8711 17731
rect 8769 17697 8803 17731
rect 9413 17697 9447 17731
rect 10057 17697 10091 17731
rect 4077 17629 4111 17663
rect 4169 17629 4203 17663
rect 4721 17629 4755 17663
rect 6745 17629 6779 17663
rect 6837 17629 6871 17663
rect 9597 17629 9631 17663
rect 1501 17561 1535 17595
rect 1685 17561 1719 17595
rect 4261 17561 4295 17595
rect 5549 17561 5583 17595
rect 6285 17561 6319 17595
rect 9873 17561 9907 17595
rect 1133 17493 1167 17527
rect 2421 17493 2455 17527
rect 3157 17493 3191 17527
rect 8125 17493 8159 17527
rect 9137 17493 9171 17527
rect 2329 17289 2363 17323
rect 3617 17289 3651 17323
rect 5641 17289 5675 17323
rect 3341 17221 3375 17255
rect 1777 17153 1811 17187
rect 3525 17153 3559 17187
rect 6837 17153 6871 17187
rect 7021 17153 7055 17187
rect 9413 17153 9447 17187
rect 2053 17085 2087 17119
rect 2237 17085 2271 17119
rect 2605 17085 2639 17119
rect 2697 17085 2731 17119
rect 2789 17085 2823 17119
rect 2973 17085 3007 17119
rect 3249 17085 3283 17119
rect 3801 17085 3835 17119
rect 3893 17085 3927 17119
rect 4077 17085 4111 17119
rect 4169 17085 4203 17119
rect 4445 17085 4479 17119
rect 4629 17085 4663 17119
rect 4721 17085 4755 17119
rect 4813 17085 4847 17119
rect 4997 17085 5031 17119
rect 5457 17085 5491 17119
rect 5825 17085 5859 17119
rect 5917 17085 5951 17119
rect 6101 17085 6135 17119
rect 6193 17085 6227 17119
rect 7389 17085 7423 17119
rect 7573 17085 7607 17119
rect 7665 17085 7699 17119
rect 7757 17085 7791 17119
rect 7941 17085 7975 17119
rect 8953 17085 8987 17119
rect 1225 17017 1259 17051
rect 5089 17017 5123 17051
rect 5273 17017 5307 17051
rect 6745 17017 6779 17051
rect 8861 17017 8895 17051
rect 9137 17017 9171 17051
rect 9680 17017 9714 17051
rect 3525 16949 3559 16983
rect 4261 16949 4295 16983
rect 6377 16949 6411 16983
rect 7205 16949 7239 16983
rect 8585 16949 8619 16983
rect 8769 16949 8803 16983
rect 10793 16949 10827 16983
rect 4997 16745 5031 16779
rect 5825 16745 5859 16779
rect 6469 16745 6503 16779
rect 7297 16745 7331 16779
rect 8217 16745 8251 16779
rect 8775 16745 8809 16779
rect 8861 16745 8895 16779
rect 9597 16745 9631 16779
rect 10425 16745 10459 16779
rect 7113 16677 7147 16711
rect 7573 16677 7607 16711
rect 7757 16677 7791 16711
rect 8401 16677 8435 16711
rect 9413 16677 9447 16711
rect 1777 16609 1811 16643
rect 2053 16609 2087 16643
rect 2605 16609 2639 16643
rect 3341 16609 3375 16643
rect 3433 16609 3467 16643
rect 4169 16609 4203 16643
rect 5089 16609 5123 16643
rect 6009 16609 6043 16643
rect 6101 16609 6135 16643
rect 6193 16609 6227 16643
rect 6285 16609 6319 16643
rect 6653 16609 6687 16643
rect 6837 16609 6871 16643
rect 6929 16609 6963 16643
rect 8125 16609 8159 16643
rect 8677 16609 8711 16643
rect 8953 16609 8987 16643
rect 9045 16609 9079 16643
rect 9873 16609 9907 16643
rect 9965 16609 9999 16643
rect 10333 16609 10367 16643
rect 10517 16609 10551 16643
rect 1225 16541 1259 16575
rect 2237 16541 2271 16575
rect 2421 16541 2455 16575
rect 2881 16541 2915 16575
rect 3525 16541 3559 16575
rect 3893 16541 3927 16575
rect 4077 16541 4111 16575
rect 5181 16541 5215 16575
rect 7389 16541 7423 16575
rect 10057 16541 10091 16575
rect 10149 16541 10183 16575
rect 8401 16473 8435 16507
rect 9689 16473 9723 16507
rect 2789 16405 2823 16439
rect 2973 16405 3007 16439
rect 4537 16405 4571 16439
rect 4629 16405 4663 16439
rect 9413 16405 9447 16439
rect 1133 16201 1167 16235
rect 2421 16201 2455 16235
rect 4077 16201 4111 16235
rect 8401 16201 8435 16235
rect 9229 16201 9263 16235
rect 10057 16201 10091 16235
rect 3249 16133 3283 16167
rect 9045 16133 9079 16167
rect 1593 16065 1627 16099
rect 3709 16065 3743 16099
rect 3801 16065 3835 16099
rect 4261 16065 4295 16099
rect 4353 16065 4387 16099
rect 4445 16065 4479 16099
rect 4537 16065 4571 16099
rect 4813 16065 4847 16099
rect 8677 16065 8711 16099
rect 1317 15997 1351 16031
rect 1501 15997 1535 16031
rect 1777 15997 1811 16031
rect 2053 15997 2087 16031
rect 2697 15997 2731 16031
rect 2789 15997 2823 16031
rect 2881 15997 2915 16031
rect 3065 15997 3099 16031
rect 3617 15997 3651 16031
rect 4721 15997 4755 16031
rect 4905 15997 4939 16031
rect 8585 15997 8619 16031
rect 8769 15997 8803 16031
rect 8861 15997 8895 16031
rect 9229 15997 9263 16031
rect 9597 15997 9631 16031
rect 9689 15997 9723 16031
rect 9873 15929 9907 15963
rect 1961 15861 1995 15895
rect 2421 15657 2455 15691
rect 2881 15657 2915 15691
rect 3341 15657 3375 15691
rect 4353 15657 4387 15691
rect 6193 15657 6227 15691
rect 7757 15657 7791 15691
rect 8585 15657 8619 15691
rect 9137 15657 9171 15691
rect 9321 15657 9355 15691
rect 10241 15657 10275 15691
rect 3617 15589 3651 15623
rect 6469 15589 6503 15623
rect 9689 15589 9723 15623
rect 10393 15589 10427 15623
rect 10609 15589 10643 15623
rect 2145 15521 2179 15555
rect 2697 15521 2731 15555
rect 2973 15521 3007 15555
rect 3065 15521 3099 15555
rect 3249 15521 3283 15555
rect 3525 15521 3559 15555
rect 3709 15521 3743 15555
rect 3893 15521 3927 15555
rect 3985 15521 4019 15555
rect 4537 15521 4571 15555
rect 4813 15521 4847 15555
rect 6377 15521 6411 15555
rect 6561 15521 6595 15555
rect 6745 15521 6779 15555
rect 6837 15521 6871 15555
rect 7389 15521 7423 15555
rect 7849 15521 7883 15555
rect 8033 15521 8067 15555
rect 8125 15521 8159 15555
rect 8401 15521 8435 15555
rect 8677 15521 8711 15555
rect 8861 15521 8895 15555
rect 8953 15521 8987 15555
rect 9229 15521 9263 15555
rect 9505 15521 9539 15555
rect 9965 15521 9999 15555
rect 2421 15453 2455 15487
rect 2513 15453 2547 15487
rect 7481 15453 7515 15487
rect 10149 15453 10183 15487
rect 3065 15385 3099 15419
rect 4629 15385 4663 15419
rect 4721 15385 4755 15419
rect 8953 15385 8987 15419
rect 2237 15317 2271 15351
rect 7849 15317 7883 15351
rect 9781 15317 9815 15351
rect 10425 15317 10459 15351
rect 2237 15113 2271 15147
rect 5181 15113 5215 15147
rect 5365 15113 5399 15147
rect 6469 15113 6503 15147
rect 8677 15113 8711 15147
rect 8861 15113 8895 15147
rect 10149 15113 10183 15147
rect 3801 15045 3835 15079
rect 4905 15045 4939 15079
rect 9137 15045 9171 15079
rect 9229 15045 9263 15079
rect 1225 14977 1259 15011
rect 1869 14977 1903 15011
rect 2789 14977 2823 15011
rect 6653 14977 6687 15011
rect 7481 14977 7515 15011
rect 7573 14977 7607 15011
rect 7849 14977 7883 15011
rect 8769 14977 8803 15011
rect 9965 14977 9999 15011
rect 1409 14909 1443 14943
rect 1685 14909 1719 14943
rect 1777 14909 1811 14943
rect 2053 14909 2087 14943
rect 2329 14909 2363 14943
rect 2513 14909 2547 14943
rect 2697 14909 2731 14943
rect 2881 14909 2915 14943
rect 3065 14909 3099 14943
rect 4077 14909 4111 14943
rect 4629 14909 4663 14943
rect 4905 14909 4939 14943
rect 5089 14909 5123 14943
rect 5825 14909 5859 14943
rect 5917 14909 5951 14943
rect 6285 14909 6319 14943
rect 6745 14909 6779 14943
rect 7389 14909 7423 14943
rect 7665 14909 7699 14943
rect 8217 14909 8251 14943
rect 8493 14909 8527 14943
rect 8585 14909 8619 14943
rect 9045 14909 9079 14943
rect 9321 14909 9355 14943
rect 9873 14909 9907 14943
rect 10333 14909 10367 14943
rect 10425 14909 10459 14943
rect 10517 14909 10551 14943
rect 3341 14841 3375 14875
rect 3525 14841 3559 14875
rect 3801 14841 3835 14875
rect 5549 14841 5583 14875
rect 6101 14841 6135 14875
rect 6193 14841 6227 14875
rect 8033 14841 8067 14875
rect 1593 14773 1627 14807
rect 3709 14773 3743 14807
rect 3985 14773 4019 14807
rect 5349 14773 5383 14807
rect 7113 14773 7147 14807
rect 7205 14773 7239 14807
rect 9505 14773 9539 14807
rect 10701 14773 10735 14807
rect 1869 14569 1903 14603
rect 2973 14569 3007 14603
rect 3065 14569 3099 14603
rect 5273 14569 5307 14603
rect 6377 14569 6411 14603
rect 7757 14569 7791 14603
rect 8033 14569 8067 14603
rect 8670 14569 8704 14603
rect 9229 14569 9263 14603
rect 10241 14569 10275 14603
rect 10425 14569 10459 14603
rect 5549 14501 5583 14535
rect 6469 14501 6503 14535
rect 7573 14501 7607 14535
rect 8861 14501 8895 14535
rect 9045 14501 9079 14535
rect 1501 14433 1535 14467
rect 2329 14433 2363 14467
rect 2513 14433 2547 14467
rect 2605 14433 2639 14467
rect 2697 14433 2731 14467
rect 3341 14433 3375 14467
rect 3433 14433 3467 14467
rect 3525 14433 3559 14467
rect 3703 14433 3737 14467
rect 4169 14433 4203 14467
rect 4721 14433 4755 14467
rect 4997 14433 5031 14467
rect 5457 14433 5491 14467
rect 5641 14433 5675 14467
rect 6034 14433 6068 14467
rect 6561 14433 6595 14467
rect 6837 14433 6871 14467
rect 6929 14433 6963 14467
rect 7849 14433 7883 14467
rect 7941 14433 7975 14467
rect 8125 14433 8159 14467
rect 8309 14433 8343 14467
rect 8401 14433 8435 14467
rect 8493 14433 8527 14467
rect 8585 14433 8619 14467
rect 8769 14433 8803 14467
rect 9137 14433 9171 14467
rect 9597 14433 9631 14467
rect 9873 14433 9907 14467
rect 10057 14433 10091 14467
rect 10333 14433 10367 14467
rect 10517 14433 10551 14467
rect 1409 14365 1443 14399
rect 3985 14365 4019 14399
rect 4077 14365 4111 14399
rect 4261 14365 4295 14399
rect 5917 14365 5951 14399
rect 6653 14365 6687 14399
rect 7021 14365 7055 14399
rect 7481 14365 7515 14399
rect 9505 14365 9539 14399
rect 7113 14297 7147 14331
rect 7573 14297 7607 14331
rect 3801 14229 3835 14263
rect 5089 14229 5123 14263
rect 8861 14229 8895 14263
rect 1501 14025 1535 14059
rect 2421 14025 2455 14059
rect 3801 14025 3835 14059
rect 6469 14025 6503 14059
rect 9781 14025 9815 14059
rect 2789 13957 2823 13991
rect 4261 13957 4295 13991
rect 5181 13957 5215 13991
rect 8953 13957 8987 13991
rect 9597 13957 9631 13991
rect 1225 13889 1259 13923
rect 2053 13889 2087 13923
rect 3617 13889 3651 13923
rect 4721 13889 4755 13923
rect 9413 13889 9447 13923
rect 1133 13821 1167 13855
rect 2145 13821 2179 13855
rect 3525 13821 3559 13855
rect 4813 13821 4847 13855
rect 6193 13821 6227 13855
rect 6469 13821 6503 13855
rect 9321 13821 9355 13855
rect 3065 13753 3099 13787
rect 4537 13753 4571 13787
rect 9749 13753 9783 13787
rect 9965 13753 9999 13787
rect 2605 13685 2639 13719
rect 4077 13685 4111 13719
rect 6285 13685 6319 13719
rect 1593 13481 1627 13515
rect 1961 13481 1995 13515
rect 6101 13481 6135 13515
rect 4261 13413 4295 13447
rect 8677 13413 8711 13447
rect 1777 13345 1811 13379
rect 2053 13345 2087 13379
rect 2605 13345 2639 13379
rect 3157 13345 3191 13379
rect 3249 13345 3283 13379
rect 3433 13345 3467 13379
rect 3525 13345 3559 13379
rect 3617 13345 3651 13379
rect 3801 13345 3835 13379
rect 3985 13345 4019 13379
rect 4077 13345 4111 13379
rect 4445 13345 4479 13379
rect 4629 13345 4663 13379
rect 4905 13345 4939 13379
rect 5089 13345 5123 13379
rect 6745 13345 6779 13379
rect 7573 13345 7607 13379
rect 7941 13345 7975 13379
rect 8125 13345 8159 13379
rect 8401 13345 8435 13379
rect 8493 13345 8527 13379
rect 9413 13345 9447 13379
rect 2329 13277 2363 13311
rect 4353 13277 4387 13311
rect 6837 13277 6871 13311
rect 2421 13209 2455 13243
rect 4261 13209 4295 13243
rect 2789 13141 2823 13175
rect 2973 13141 3007 13175
rect 3709 13141 3743 13175
rect 4813 13141 4847 13175
rect 4997 13141 5031 13175
rect 7665 13141 7699 13175
rect 8677 13141 8711 13175
rect 9229 13141 9263 13175
rect 3065 12937 3099 12971
rect 3709 12937 3743 12971
rect 9137 12937 9171 12971
rect 10333 12937 10367 12971
rect 5273 12869 5307 12903
rect 8953 12869 8987 12903
rect 2053 12801 2087 12835
rect 2513 12801 2547 12835
rect 3893 12801 3927 12835
rect 4721 12801 4755 12835
rect 8493 12801 8527 12835
rect 9505 12801 9539 12835
rect 9597 12801 9631 12835
rect 9873 12801 9907 12835
rect 10057 12801 10091 12835
rect 10517 12801 10551 12835
rect 1225 12733 1259 12767
rect 1685 12733 1719 12767
rect 3249 12733 3283 12767
rect 3525 12733 3559 12767
rect 4537 12733 4571 12767
rect 6009 12733 6043 12767
rect 6101 12733 6135 12767
rect 6653 12733 6687 12767
rect 6929 12733 6963 12767
rect 7113 12733 7147 12767
rect 7573 12733 7607 12767
rect 7757 12733 7791 12767
rect 7849 12733 7883 12767
rect 7941 12733 7975 12767
rect 8125 12733 8159 12767
rect 8585 12733 8619 12767
rect 9321 12733 9355 12767
rect 9413 12733 9447 12767
rect 9965 12733 9999 12767
rect 10149 12733 10183 12767
rect 10425 12733 10459 12767
rect 10609 12733 10643 12767
rect 2697 12665 2731 12699
rect 5089 12665 5123 12699
rect 7205 12665 7239 12699
rect 7297 12665 7331 12699
rect 8033 12665 8067 12699
rect 2605 12597 2639 12631
rect 3341 12597 3375 12631
rect 7389 12597 7423 12631
rect 2697 12393 2731 12427
rect 2881 12393 2915 12427
rect 4077 12393 4111 12427
rect 4261 12393 4295 12427
rect 5365 12393 5399 12427
rect 6561 12393 6595 12427
rect 9505 12393 9539 12427
rect 10241 12393 10275 12427
rect 2237 12325 2271 12359
rect 3433 12325 3467 12359
rect 4813 12325 4847 12359
rect 6101 12325 6135 12359
rect 8309 12325 8343 12359
rect 8861 12325 8895 12359
rect 10609 12325 10643 12359
rect 1593 12257 1627 12291
rect 1961 12257 1995 12291
rect 2421 12257 2455 12291
rect 2878 12257 2912 12291
rect 3617 12257 3651 12291
rect 3801 12257 3835 12291
rect 3893 12257 3927 12291
rect 4258 12257 4292 12291
rect 4997 12257 5031 12291
rect 5089 12257 5123 12291
rect 5181 12257 5215 12291
rect 5457 12257 5491 12291
rect 6285 12257 6319 12291
rect 6377 12257 6411 12291
rect 6745 12257 6779 12291
rect 7297 12257 7331 12291
rect 7481 12257 7515 12291
rect 7757 12257 7791 12291
rect 8033 12257 8067 12291
rect 8217 12257 8251 12291
rect 8493 12257 8527 12291
rect 8769 12257 8803 12291
rect 8953 12257 8987 12291
rect 9137 12257 9171 12291
rect 9321 12257 9355 12291
rect 9781 12257 9815 12291
rect 10425 12257 10459 12291
rect 2237 12189 2271 12223
rect 3341 12189 3375 12223
rect 4721 12189 4755 12223
rect 7021 12189 7055 12223
rect 8677 12189 8711 12223
rect 9873 12189 9907 12223
rect 4813 12121 4847 12155
rect 5181 12121 5215 12155
rect 7573 12121 7607 12155
rect 10149 12121 10183 12155
rect 1409 12053 1443 12087
rect 2053 12053 2087 12087
rect 2513 12053 2547 12087
rect 3249 12053 3283 12087
rect 4629 12053 4663 12087
rect 6101 12053 6135 12087
rect 6929 12053 6963 12087
rect 7389 12053 7423 12087
rect 2605 11849 2639 11883
rect 3249 11849 3283 11883
rect 3801 11849 3835 11883
rect 6193 11849 6227 11883
rect 6745 11849 6779 11883
rect 7297 11849 7331 11883
rect 8125 11849 8159 11883
rect 8861 11849 8895 11883
rect 10241 11849 10275 11883
rect 7941 11713 7975 11747
rect 8677 11713 8711 11747
rect 9045 11713 9079 11747
rect 9597 11713 9631 11747
rect 10333 11713 10367 11747
rect 1593 11645 1627 11679
rect 1961 11645 1995 11679
rect 2605 11645 2639 11679
rect 2789 11645 2823 11679
rect 3433 11645 3467 11679
rect 3709 11645 3743 11679
rect 3801 11645 3835 11679
rect 3985 11645 4019 11679
rect 5917 11645 5951 11679
rect 6193 11645 6227 11679
rect 6929 11645 6963 11679
rect 7205 11645 7239 11679
rect 7297 11645 7331 11679
rect 7481 11645 7515 11679
rect 7665 11645 7699 11679
rect 7849 11645 7883 11679
rect 8198 11645 8232 11679
rect 8585 11645 8619 11679
rect 9505 11645 9539 11679
rect 9689 11645 9723 11679
rect 10057 11645 10091 11679
rect 10609 11645 10643 11679
rect 7113 11577 7147 11611
rect 7757 11577 7791 11611
rect 9229 11577 9263 11611
rect 9413 11577 9447 11611
rect 10425 11577 10459 11611
rect 1409 11509 1443 11543
rect 1777 11509 1811 11543
rect 3617 11509 3651 11543
rect 6009 11509 6043 11543
rect 7941 11509 7975 11543
rect 9873 11509 9907 11543
rect 10793 11509 10827 11543
rect 1777 11305 1811 11339
rect 3065 11305 3099 11339
rect 4721 11305 4755 11339
rect 4905 11305 4939 11339
rect 6193 11305 6227 11339
rect 9413 11305 9447 11339
rect 10057 11305 10091 11339
rect 10149 11305 10183 11339
rect 2697 11237 2731 11271
rect 5457 11237 5491 11271
rect 8861 11237 8895 11271
rect 1685 11169 1719 11203
rect 1869 11169 1903 11203
rect 2145 11169 2179 11203
rect 2605 11169 2639 11203
rect 2881 11169 2915 11203
rect 4261 11169 4295 11203
rect 4353 11169 4387 11203
rect 4537 11169 4571 11203
rect 4819 11169 4853 11203
rect 4997 11169 5031 11203
rect 5365 11169 5399 11203
rect 5641 11169 5675 11203
rect 5825 11169 5859 11203
rect 6009 11169 6043 11203
rect 6561 11169 6595 11203
rect 8677 11169 8711 11203
rect 8953 11169 8987 11203
rect 9229 11169 9263 11203
rect 9413 11169 9447 11203
rect 9873 11169 9907 11203
rect 10057 11169 10091 11203
rect 10149 11169 10183 11203
rect 10333 11169 10367 11203
rect 2237 11101 2271 11135
rect 6653 11101 6687 11135
rect 6929 11101 6963 11135
rect 2513 11033 2547 11067
rect 5641 11033 5675 11067
rect 8493 11033 8527 11067
rect 1869 10761 1903 10795
rect 2237 10761 2271 10795
rect 2513 10761 2547 10795
rect 6377 10761 6411 10795
rect 7573 10761 7607 10795
rect 4261 10693 4295 10727
rect 4997 10693 5031 10727
rect 5825 10693 5859 10727
rect 1225 10625 1259 10659
rect 1777 10625 1811 10659
rect 3985 10625 4019 10659
rect 5549 10625 5583 10659
rect 6561 10625 6595 10659
rect 7849 10625 7883 10659
rect 1133 10557 1167 10591
rect 1317 10557 1351 10591
rect 1409 10557 1443 10591
rect 2053 10557 2087 10591
rect 2329 10557 2363 10591
rect 2421 10557 2455 10591
rect 2605 10557 2639 10591
rect 3893 10557 3927 10591
rect 5273 10557 5307 10591
rect 5457 10557 5491 10591
rect 5641 10557 5675 10591
rect 5733 10557 5767 10591
rect 5917 10557 5951 10591
rect 6193 10557 6227 10591
rect 6469 10557 6503 10591
rect 6929 10557 6963 10591
rect 7205 10557 7239 10591
rect 7389 10557 7423 10591
rect 7481 10557 7515 10591
rect 7665 10557 7699 10591
rect 7757 10557 7791 10591
rect 7941 10557 7975 10591
rect 8953 10557 8987 10591
rect 9137 10557 9171 10591
rect 9597 10557 9631 10591
rect 9781 10557 9815 10591
rect 1593 10489 1627 10523
rect 4997 10489 5031 10523
rect 5181 10489 5215 10523
rect 6745 10489 6779 10523
rect 7021 10489 7055 10523
rect 6009 10421 6043 10455
rect 8953 10421 8987 10455
rect 9781 10421 9815 10455
rect 3341 10217 3375 10251
rect 5273 10217 5307 10251
rect 5549 10217 5583 10251
rect 7021 10217 7055 10251
rect 9229 10217 9263 10251
rect 10425 10217 10459 10251
rect 3157 10149 3191 10183
rect 5365 10149 5399 10183
rect 7481 10149 7515 10183
rect 1409 10081 1443 10115
rect 1869 10081 1903 10115
rect 2053 10081 2087 10115
rect 3065 10081 3099 10115
rect 3249 10081 3283 10115
rect 3525 10081 3559 10115
rect 3801 10081 3835 10115
rect 3893 10081 3927 10115
rect 4077 10081 4111 10115
rect 4353 10081 4387 10115
rect 4537 10081 4571 10115
rect 4905 10081 4939 10115
rect 5641 10081 5675 10115
rect 6193 10081 6227 10115
rect 6377 10081 6411 10115
rect 6653 10081 6687 10115
rect 6837 10081 6871 10115
rect 7113 10081 7147 10115
rect 7297 10081 7331 10115
rect 8861 10081 8895 10115
rect 9597 10081 9631 10115
rect 10241 10081 10275 10115
rect 10517 10081 10551 10115
rect 10701 10081 10735 10115
rect 1501 10013 1535 10047
rect 2329 10013 2363 10047
rect 4261 10013 4295 10047
rect 4997 10013 5031 10047
rect 8953 10013 8987 10047
rect 9505 10013 9539 10047
rect 10057 10013 10091 10047
rect 10609 10013 10643 10047
rect 3709 9945 3743 9979
rect 4445 9945 4479 9979
rect 5365 9945 5399 9979
rect 6009 9945 6043 9979
rect 9965 9945 9999 9979
rect 1685 9877 1719 9911
rect 2237 9877 2271 9911
rect 5181 9673 5215 9707
rect 6193 9673 6227 9707
rect 6377 9673 6411 9707
rect 6745 9673 6779 9707
rect 8953 9673 8987 9707
rect 9965 9673 9999 9707
rect 1961 9605 1995 9639
rect 2605 9605 2639 9639
rect 4353 9605 4387 9639
rect 6009 9605 6043 9639
rect 1685 9537 1719 9571
rect 2329 9537 2363 9571
rect 4077 9537 4111 9571
rect 5733 9537 5767 9571
rect 8677 9537 8711 9571
rect 9229 9537 9263 9571
rect 9321 9537 9355 9571
rect 9413 9537 9447 9571
rect 1593 9469 1627 9503
rect 2237 9469 2271 9503
rect 2697 9469 2731 9503
rect 2881 9469 2915 9503
rect 3985 9469 4019 9503
rect 4445 9469 4479 9503
rect 4629 9469 4663 9503
rect 4905 9469 4939 9503
rect 5089 9469 5123 9503
rect 5181 9469 5215 9503
rect 5365 9469 5399 9503
rect 5641 9469 5675 9503
rect 6653 9469 6687 9503
rect 6837 9469 6871 9503
rect 8585 9469 8619 9503
rect 9505 9469 9539 9503
rect 10149 9469 10183 9503
rect 10333 9469 10367 9503
rect 2789 9401 2823 9435
rect 6345 9401 6379 9435
rect 6561 9401 6595 9435
rect 9045 9333 9079 9367
rect 1317 9129 1351 9163
rect 2329 9129 2363 9163
rect 4077 9129 4111 9163
rect 4721 9129 4755 9163
rect 4905 9129 4939 9163
rect 7297 9129 7331 9163
rect 9137 9129 9171 9163
rect 2145 9061 2179 9095
rect 2513 9061 2547 9095
rect 3341 9061 3375 9095
rect 9229 9061 9263 9095
rect 1685 8993 1719 9027
rect 1961 8993 1995 9027
rect 2421 8993 2455 9027
rect 2605 8993 2639 9027
rect 3249 8993 3283 9027
rect 3433 8993 3467 9027
rect 3709 8993 3743 9027
rect 3893 8993 3927 9027
rect 3985 8993 4019 9027
rect 4077 8993 4111 9027
rect 4261 8993 4295 9027
rect 4353 8993 4387 9027
rect 4537 8993 4571 9027
rect 4813 8993 4847 9027
rect 4997 8993 5031 9027
rect 7481 8993 7515 9027
rect 8953 8993 8987 9027
rect 9413 8993 9447 9027
rect 1593 8925 1627 8959
rect 7757 8925 7791 8959
rect 8033 8925 8067 8959
rect 8125 8925 8159 8959
rect 8217 8925 8251 8959
rect 8309 8925 8343 8959
rect 8769 8925 8803 8959
rect 9689 8925 9723 8959
rect 3525 8857 3559 8891
rect 7665 8789 7699 8823
rect 7849 8789 7883 8823
rect 9597 8789 9631 8823
rect 4169 8585 4203 8619
rect 8401 8585 8435 8619
rect 8861 8585 8895 8619
rect 9597 8585 9631 8619
rect 10609 8585 10643 8619
rect 2053 8517 2087 8551
rect 8217 8517 8251 8551
rect 1593 8449 1627 8483
rect 7389 8449 7423 8483
rect 7665 8449 7699 8483
rect 10517 8449 10551 8483
rect 1685 8381 1719 8415
rect 7297 8381 7331 8415
rect 8677 8381 8711 8415
rect 8769 8381 8803 8415
rect 8953 8381 8987 8415
rect 9321 8381 9355 8415
rect 9505 8381 9539 8415
rect 9781 8381 9815 8415
rect 9965 8381 9999 8415
rect 10057 8381 10091 8415
rect 10609 8381 10643 8415
rect 10793 8381 10827 8415
rect 3801 8313 3835 8347
rect 3985 8313 4019 8347
rect 7849 8313 7883 8347
rect 8033 8313 8067 8347
rect 8401 8313 8435 8347
rect 8585 8313 8619 8347
rect 10149 8313 10183 8347
rect 10333 8313 10367 8347
rect 9321 8245 9355 8279
rect 2605 8041 2639 8075
rect 9413 8041 9447 8075
rect 6285 7973 6319 8007
rect 7113 7973 7147 8007
rect 8493 7973 8527 8007
rect 8769 7973 8803 8007
rect 9045 7973 9079 8007
rect 9245 7973 9279 8007
rect 1593 7905 1627 7939
rect 1961 7905 1995 7939
rect 6469 7905 6503 7939
rect 6653 7905 6687 7939
rect 7205 7905 7239 7939
rect 7481 7905 7515 7939
rect 7665 7905 7699 7939
rect 7757 7905 7791 7939
rect 8401 7903 8435 7937
rect 8585 7905 8619 7939
rect 8677 7905 8711 7939
rect 8953 7905 8987 7939
rect 9689 7905 9723 7939
rect 10333 7905 10367 7939
rect 10425 7905 10459 7939
rect 10609 7905 10643 7939
rect 10793 7905 10827 7939
rect 6745 7837 6779 7871
rect 7849 7837 7883 7871
rect 8309 7837 8343 7871
rect 9781 7837 9815 7871
rect 10149 7837 10183 7871
rect 8125 7769 8159 7803
rect 8953 7769 8987 7803
rect 10057 7769 10091 7803
rect 6929 7701 6963 7735
rect 7297 7701 7331 7735
rect 9229 7701 9263 7735
rect 10609 7701 10643 7735
rect 1041 7497 1075 7531
rect 2881 7497 2915 7531
rect 5365 7497 5399 7531
rect 6745 7497 6779 7531
rect 7573 7497 7607 7531
rect 7665 7497 7699 7531
rect 9045 7497 9079 7531
rect 10517 7497 10551 7531
rect 949 7429 983 7463
rect 1777 7429 1811 7463
rect 2421 7429 2455 7463
rect 1133 7361 1167 7395
rect 1501 7361 1535 7395
rect 1961 7361 1995 7395
rect 2973 7361 3007 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 7021 7361 7055 7395
rect 9229 7361 9263 7395
rect 857 7293 891 7327
rect 1409 7293 1443 7327
rect 2053 7293 2087 7327
rect 2697 7293 2731 7327
rect 3433 7293 3467 7327
rect 3617 7293 3651 7327
rect 4629 7293 4663 7327
rect 4813 7293 4847 7327
rect 5549 7293 5583 7327
rect 5733 7293 5767 7327
rect 5917 7293 5951 7327
rect 6101 7293 6135 7327
rect 6193 7293 6227 7327
rect 6377 7293 6411 7327
rect 6653 7293 6687 7327
rect 6828 7295 6862 7329
rect 6929 7293 6963 7327
rect 7113 7293 7147 7327
rect 7297 7293 7331 7327
rect 7389 7293 7423 7327
rect 8033 7293 8067 7327
rect 9321 7293 9355 7327
rect 9597 7293 9631 7327
rect 9781 7293 9815 7327
rect 10057 7293 10091 7327
rect 10333 7293 10367 7327
rect 10517 7293 10551 7327
rect 7849 7225 7883 7259
rect 2513 7157 2547 7191
rect 3801 7157 3835 7191
rect 4721 7157 4755 7191
rect 6285 7157 6319 7191
rect 10241 7157 10275 7191
rect 2237 6953 2271 6987
rect 5641 6953 5675 6987
rect 6929 6953 6963 6987
rect 7941 6953 7975 6987
rect 9413 6953 9447 6987
rect 1225 6817 1259 6851
rect 1685 6817 1719 6851
rect 1869 6817 1903 6851
rect 2053 6817 2087 6851
rect 2145 6817 2179 6851
rect 2237 6817 2271 6851
rect 2421 6817 2455 6851
rect 2513 6817 2547 6851
rect 2697 6817 2731 6851
rect 2789 6817 2823 6851
rect 2973 6817 3007 6851
rect 3249 6817 3283 6851
rect 3893 6817 3927 6851
rect 4353 6817 4387 6851
rect 4537 6817 4571 6851
rect 4813 6817 4847 6851
rect 4997 6817 5031 6851
rect 5273 6817 5307 6851
rect 6009 6817 6043 6851
rect 6285 6817 6319 6851
rect 6561 6817 6595 6851
rect 7205 6817 7239 6851
rect 7757 6817 7791 6851
rect 8033 6817 8067 6851
rect 8125 6817 8159 6851
rect 8309 6817 8343 6851
rect 9321 6817 9355 6851
rect 9597 6817 9631 6851
rect 1317 6749 1351 6783
rect 1593 6749 1627 6783
rect 3157 6749 3191 6783
rect 3801 6749 3835 6783
rect 5365 6749 5399 6783
rect 5825 6749 5859 6783
rect 6653 6749 6687 6783
rect 7021 6749 7055 6783
rect 7481 6749 7515 6783
rect 2513 6681 2547 6715
rect 3617 6681 3651 6715
rect 4261 6681 4295 6715
rect 6193 6681 6227 6715
rect 2973 6613 3007 6647
rect 7389 6613 7423 6647
rect 7573 6613 7607 6647
rect 8125 6613 8159 6647
rect 9781 6613 9815 6647
rect 2421 6409 2455 6443
rect 3709 6409 3743 6443
rect 4721 6409 4755 6443
rect 4997 6409 5031 6443
rect 5365 6409 5399 6443
rect 6377 6409 6411 6443
rect 7113 6409 7147 6443
rect 3433 6341 3467 6375
rect 3801 6341 3835 6375
rect 4353 6273 4387 6307
rect 7021 6273 7055 6307
rect 2145 6205 2179 6239
rect 2237 6205 2271 6239
rect 3249 6205 3283 6239
rect 3433 6205 3467 6239
rect 3801 6205 3835 6239
rect 3985 6205 4019 6239
rect 4537 6205 4571 6239
rect 4813 6205 4847 6239
rect 4997 6205 5031 6239
rect 5549 6205 5583 6239
rect 5825 6205 5859 6239
rect 6469 6205 6503 6239
rect 6653 6205 6687 6239
rect 6837 6205 6871 6239
rect 6929 6205 6963 6239
rect 7205 6205 7239 6239
rect 7297 6205 7331 6239
rect 8953 6205 8987 6239
rect 9137 6205 9171 6239
rect 9229 6205 9263 6239
rect 5733 6137 5767 6171
rect 6009 6137 6043 6171
rect 6193 6137 6227 6171
rect 1777 6069 1811 6103
rect 8769 6069 8803 6103
rect 1317 5865 1351 5899
rect 2697 5865 2731 5899
rect 7481 5865 7515 5899
rect 8125 5865 8159 5899
rect 9321 5865 9355 5899
rect 10425 5865 10459 5899
rect 2881 5797 2915 5831
rect 9689 5797 9723 5831
rect 10241 5797 10275 5831
rect 1225 5729 1259 5763
rect 1409 5729 1443 5763
rect 1685 5729 1719 5763
rect 2329 5729 2363 5763
rect 2789 5729 2823 5763
rect 2973 5729 3007 5763
rect 6193 5729 6227 5763
rect 7021 5729 7055 5763
rect 7665 5729 7699 5763
rect 7849 5729 7883 5763
rect 7941 5729 7975 5763
rect 8033 5729 8067 5763
rect 8217 5729 8251 5763
rect 9505 5729 9539 5763
rect 9781 5729 9815 5763
rect 10057 5729 10091 5763
rect 10333 5729 10367 5763
rect 10517 5729 10551 5763
rect 10609 5729 10643 5763
rect 10793 5729 10827 5763
rect 1777 5661 1811 5695
rect 2237 5661 2271 5695
rect 6285 5661 6319 5695
rect 6929 5661 6963 5695
rect 9873 5661 9907 5695
rect 2053 5593 2087 5627
rect 7389 5593 7423 5627
rect 5825 5525 5859 5559
rect 10701 5525 10735 5559
rect 2145 5321 2179 5355
rect 6929 5321 6963 5355
rect 7021 5321 7055 5355
rect 9413 5321 9447 5355
rect 3801 5253 3835 5287
rect 5825 5253 5859 5287
rect 9597 5253 9631 5287
rect 10609 5253 10643 5287
rect 3525 5185 3559 5219
rect 6653 5185 6687 5219
rect 8769 5185 8803 5219
rect 9873 5185 9907 5219
rect 10701 5185 10735 5219
rect 2421 5117 2455 5151
rect 2513 5117 2547 5151
rect 3433 5117 3467 5151
rect 4905 5117 4939 5151
rect 5089 5117 5123 5151
rect 5365 5117 5399 5151
rect 5457 5117 5491 5151
rect 5580 5117 5614 5151
rect 6285 5117 6319 5151
rect 6561 5117 6595 5151
rect 7205 5117 7239 5151
rect 7297 5117 7331 5151
rect 7849 5117 7883 5151
rect 8033 5117 8067 5151
rect 8401 5117 8435 5151
rect 8861 5117 8895 5151
rect 9045 5117 9079 5151
rect 9229 5117 9263 5151
rect 9321 5117 9355 5151
rect 9505 5117 9539 5151
rect 9965 5117 9999 5151
rect 10425 5117 10459 5151
rect 1777 5049 1811 5083
rect 1961 5049 1995 5083
rect 5273 5049 5307 5083
rect 5917 5049 5951 5083
rect 6101 5049 6135 5083
rect 8585 5049 8619 5083
rect 2237 4981 2271 5015
rect 7941 4981 7975 5015
rect 10241 4981 10275 5015
rect 2053 4777 2087 4811
rect 2789 4777 2823 4811
rect 3157 4777 3191 4811
rect 3709 4777 3743 4811
rect 5365 4777 5399 4811
rect 7849 4777 7883 4811
rect 8309 4777 8343 4811
rect 8953 4777 8987 4811
rect 9965 4777 9999 4811
rect 10609 4777 10643 4811
rect 2237 4709 2271 4743
rect 4169 4709 4203 4743
rect 8217 4709 8251 4743
rect 8461 4709 8495 4743
rect 8677 4709 8711 4743
rect 9597 4709 9631 4743
rect 9781 4709 9815 4743
rect 10241 4709 10275 4743
rect 1132 4641 1166 4675
rect 1225 4641 1259 4675
rect 1501 4641 1535 4675
rect 1961 4641 1995 4675
rect 2329 4641 2363 4675
rect 2513 4641 2547 4675
rect 2697 4641 2731 4675
rect 2973 4641 3007 4675
rect 3249 4641 3283 4675
rect 3341 4641 3375 4675
rect 3495 4641 3529 4675
rect 3801 4641 3835 4675
rect 3985 4641 4019 4675
rect 4997 4641 5031 4675
rect 5181 4641 5215 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 9321 4641 9355 4675
rect 10057 4641 10091 4675
rect 10517 4641 10551 4675
rect 10701 4641 10735 4675
rect 857 4573 891 4607
rect 1409 4573 1443 4607
rect 7205 4573 7239 4607
rect 9413 4573 9447 4607
rect 10425 4573 10459 4607
rect 1869 4505 1903 4539
rect 7665 4505 7699 4539
rect 2237 4437 2271 4471
rect 8493 4437 8527 4471
rect 1409 4233 1443 4267
rect 3985 4233 4019 4267
rect 8677 4233 8711 4267
rect 3065 4165 3099 4199
rect 3801 4165 3835 4199
rect 5181 4165 5215 4199
rect 6929 4165 6963 4199
rect 7849 4165 7883 4199
rect 2145 4097 2179 4131
rect 2421 4097 2455 4131
rect 2605 4097 2639 4131
rect 3525 4097 3559 4131
rect 4169 4097 4203 4131
rect 4813 4097 4847 4131
rect 5549 4097 5583 4131
rect 9505 4097 9539 4131
rect 9873 4097 9907 4131
rect 2053 4029 2087 4063
rect 2697 4029 2731 4063
rect 3433 4029 3467 4063
rect 4261 4029 4295 4063
rect 4537 4029 4571 4063
rect 4721 4029 4755 4063
rect 4997 4029 5031 4063
rect 5089 4029 5123 4063
rect 5365 4029 5399 4063
rect 5641 4029 5675 4063
rect 5733 4029 5767 4063
rect 6653 4029 6687 4063
rect 6929 4029 6963 4063
rect 7849 4029 7883 4063
rect 8033 4029 8067 4063
rect 8125 4029 8159 4063
rect 8493 4029 8527 4063
rect 8677 4029 8711 4063
rect 8953 4029 8987 4063
rect 9229 4029 9263 4063
rect 9413 4029 9447 4063
rect 9689 4029 9723 4063
rect 9965 4029 9999 4063
rect 10149 4029 10183 4063
rect 1593 3961 1627 3995
rect 1777 3961 1811 3995
rect 4813 3961 4847 3995
rect 5917 3961 5951 3995
rect 10057 3961 10091 3995
rect 4721 3893 4755 3927
rect 6101 3893 6135 3927
rect 6745 3893 6779 3927
rect 8769 3893 8803 3927
rect 3709 3689 3743 3723
rect 2405 3621 2439 3655
rect 2605 3621 2639 3655
rect 6561 3621 6595 3655
rect 9045 3621 9079 3655
rect 3341 3553 3375 3587
rect 4353 3553 4387 3587
rect 4537 3553 4571 3587
rect 4629 3553 4663 3587
rect 4813 3553 4847 3587
rect 5273 3553 5307 3587
rect 6193 3553 6227 3587
rect 6469 3553 6503 3587
rect 6653 3553 6687 3587
rect 8033 3553 8067 3587
rect 8309 3553 8343 3587
rect 8861 3553 8895 3587
rect 9137 3553 9171 3587
rect 9505 3553 9539 3587
rect 3249 3485 3283 3519
rect 5365 3485 5399 3519
rect 5641 3485 5675 3519
rect 6101 3485 6135 3519
rect 8217 3485 8251 3519
rect 8493 3417 8527 3451
rect 2237 3349 2271 3383
rect 2421 3349 2455 3383
rect 4445 3349 4479 3383
rect 4997 3349 5031 3383
rect 5917 3349 5951 3383
rect 7849 3349 7883 3383
rect 8677 3349 8711 3383
rect 9321 3349 9355 3383
rect 9689 3349 9723 3383
rect 2881 3145 2915 3179
rect 5641 3145 5675 3179
rect 7205 3145 7239 3179
rect 8125 3145 8159 3179
rect 8769 3145 8803 3179
rect 10425 3145 10459 3179
rect 10701 3145 10735 3179
rect 2513 3077 2547 3111
rect 3433 3077 3467 3111
rect 5825 3077 5859 3111
rect 1041 3009 1075 3043
rect 5181 3009 5215 3043
rect 9045 3009 9079 3043
rect 3249 2941 3283 2975
rect 5273 2941 5307 2975
rect 5733 2941 5767 2975
rect 5917 2941 5951 2975
rect 8401 2941 8435 2975
rect 10517 2941 10551 2975
rect 1308 2873 1342 2907
rect 7189 2873 7223 2907
rect 7389 2873 7423 2907
rect 7849 2873 7883 2907
rect 8769 2873 8803 2907
rect 9290 2873 9324 2907
rect 2421 2805 2455 2839
rect 2881 2805 2915 2839
rect 3065 2805 3099 2839
rect 7021 2805 7055 2839
rect 8953 2805 8987 2839
rect 1593 2601 1627 2635
rect 3249 2601 3283 2635
rect 7941 2601 7975 2635
rect 8033 2601 8067 2635
rect 1133 2533 1167 2567
rect 1501 2533 1535 2567
rect 1777 2533 1811 2567
rect 2237 2533 2271 2567
rect 3801 2533 3835 2567
rect 9657 2533 9691 2567
rect 9873 2533 9907 2567
rect 1317 2465 1351 2499
rect 2421 2465 2455 2499
rect 2789 2465 2823 2499
rect 2973 2465 3007 2499
rect 3433 2465 3467 2499
rect 4353 2465 4387 2499
rect 6561 2465 6595 2499
rect 6828 2465 6862 2499
rect 9157 2465 9191 2499
rect 9413 2465 9447 2499
rect 2881 2397 2915 2431
rect 3065 2397 3099 2431
rect 2145 2329 2179 2363
rect 9505 2329 9539 2363
rect 1777 2261 1811 2295
rect 2605 2261 2639 2295
rect 3801 2261 3835 2295
rect 3985 2261 4019 2295
rect 4169 2261 4203 2295
rect 9689 2261 9723 2295
rect 1593 2057 1627 2091
rect 3709 2057 3743 2091
rect 5181 2057 5215 2091
rect 6929 2057 6963 2091
rect 7113 2057 7147 2091
rect 8769 2057 8803 2091
rect 8953 2057 8987 2091
rect 6561 1989 6595 2023
rect 8033 1989 8067 2023
rect 1225 1921 1259 1955
rect 7481 1921 7515 1955
rect 7573 1921 7607 1955
rect 7757 1921 7791 1955
rect 1409 1853 1443 1887
rect 3065 1853 3099 1887
rect 3801 1853 3835 1887
rect 7665 1853 7699 1887
rect 7941 1853 7975 1887
rect 8125 1853 8159 1887
rect 8585 1853 8619 1887
rect 9045 1853 9079 1887
rect 2820 1785 2854 1819
rect 3341 1785 3375 1819
rect 3525 1785 3559 1819
rect 4068 1785 4102 1819
rect 6929 1785 6963 1819
rect 8401 1785 8435 1819
rect 1685 1717 1719 1751
rect 7297 1717 7331 1751
rect 2789 1513 2823 1547
rect 2881 1513 2915 1547
rect 2237 1445 2271 1479
rect 4537 1445 4571 1479
rect 2145 1377 2179 1411
rect 2329 1377 2363 1411
rect 2605 1377 2639 1411
rect 3994 1377 4028 1411
rect 2421 1309 2455 1343
rect 4261 1309 4295 1343
rect 4353 1309 4387 1343
rect 3249 969 3283 1003
rect 3433 969 3467 1003
rect 3401 697 3435 731
rect 3617 697 3651 731
<< metal1 >>
rect 5810 43596 5816 43648
rect 5868 43636 5874 43648
rect 10502 43636 10508 43648
rect 5868 43608 10508 43636
rect 5868 43596 5874 43608
rect 10502 43596 10508 43608
rect 10560 43596 10566 43648
rect 552 43002 11132 43024
rect 552 42950 4322 43002
rect 4374 42950 4386 43002
rect 4438 42950 4450 43002
rect 4502 42950 4514 43002
rect 4566 42950 4578 43002
rect 4630 42950 10722 43002
rect 10774 42950 10786 43002
rect 10838 42950 10850 43002
rect 10902 42950 10914 43002
rect 10966 42950 10978 43002
rect 11030 42950 11132 43002
rect 552 42928 11132 42950
rect 1762 42848 1768 42900
rect 1820 42888 1826 42900
rect 2130 42888 2136 42900
rect 1820 42860 2136 42888
rect 1820 42848 1826 42860
rect 2130 42848 2136 42860
rect 2188 42848 2194 42900
rect 3881 42891 3939 42897
rect 3881 42857 3893 42891
rect 3927 42888 3939 42891
rect 5261 42891 5319 42897
rect 5261 42888 5273 42891
rect 3927 42860 5273 42888
rect 3927 42857 3939 42860
rect 3881 42851 3939 42857
rect 5261 42857 5273 42860
rect 5307 42857 5319 42891
rect 10597 42891 10655 42897
rect 10597 42888 10609 42891
rect 5261 42851 5319 42857
rect 9140 42860 10609 42888
rect 1121 42823 1179 42829
rect 1121 42789 1133 42823
rect 1167 42820 1179 42823
rect 5626 42820 5632 42832
rect 1167 42792 5632 42820
rect 1167 42789 1179 42792
rect 1121 42783 1179 42789
rect 5626 42780 5632 42792
rect 5684 42780 5690 42832
rect 5997 42823 6055 42829
rect 5997 42789 6009 42823
rect 6043 42820 6055 42823
rect 6638 42820 6644 42832
rect 6043 42792 6644 42820
rect 6043 42789 6055 42792
rect 5997 42783 6055 42789
rect 6638 42780 6644 42792
rect 6696 42780 6702 42832
rect 9033 42823 9091 42829
rect 9033 42820 9045 42823
rect 6886 42792 9045 42820
rect 1857 42755 1915 42761
rect 1857 42721 1869 42755
rect 1903 42752 1915 42755
rect 2314 42752 2320 42764
rect 1903 42724 2320 42752
rect 1903 42721 1915 42724
rect 1857 42715 1915 42721
rect 2314 42712 2320 42724
rect 2372 42712 2378 42764
rect 3050 42712 3056 42764
rect 3108 42712 3114 42764
rect 3878 42712 3884 42764
rect 3936 42752 3942 42764
rect 3973 42755 4031 42761
rect 3973 42752 3985 42755
rect 3936 42724 3985 42752
rect 3936 42712 3942 42724
rect 3973 42721 3985 42724
rect 4019 42721 4031 42755
rect 3973 42715 4031 42721
rect 4356 42724 6132 42752
rect 2038 42644 2044 42696
rect 2096 42644 2102 42696
rect 2777 42687 2835 42693
rect 2777 42653 2789 42687
rect 2823 42653 2835 42687
rect 2777 42647 2835 42653
rect 3329 42687 3387 42693
rect 3329 42653 3341 42687
rect 3375 42653 3387 42687
rect 3329 42647 3387 42653
rect 1305 42619 1363 42625
rect 1305 42585 1317 42619
rect 1351 42616 1363 42619
rect 1351 42588 2084 42616
rect 1351 42585 1363 42588
rect 1305 42579 1363 42585
rect 1397 42551 1455 42557
rect 1397 42517 1409 42551
rect 1443 42548 1455 42551
rect 1578 42548 1584 42560
rect 1443 42520 1584 42548
rect 1443 42517 1455 42520
rect 1397 42511 1455 42517
rect 1578 42508 1584 42520
rect 1636 42508 1642 42560
rect 2056 42548 2084 42588
rect 2130 42576 2136 42628
rect 2188 42616 2194 42628
rect 2792 42616 2820 42647
rect 2188 42588 2820 42616
rect 3344 42616 3372 42647
rect 4246 42644 4252 42696
rect 4304 42644 4310 42696
rect 4356 42628 4384 42724
rect 4706 42644 4712 42696
rect 4764 42684 4770 42696
rect 5353 42687 5411 42693
rect 5353 42684 5365 42687
rect 4764 42656 5365 42684
rect 4764 42644 4770 42656
rect 5353 42653 5365 42656
rect 5399 42653 5411 42687
rect 5353 42647 5411 42653
rect 5445 42687 5503 42693
rect 5445 42653 5457 42687
rect 5491 42653 5503 42687
rect 6104 42684 6132 42724
rect 6178 42712 6184 42764
rect 6236 42712 6242 42764
rect 6886 42752 6914 42792
rect 9033 42789 9045 42792
rect 9079 42789 9091 42823
rect 9033 42783 9091 42789
rect 6380 42724 6914 42752
rect 6380 42684 6408 42724
rect 7190 42712 7196 42764
rect 7248 42752 7254 42764
rect 7285 42755 7343 42761
rect 7285 42752 7297 42755
rect 7248 42724 7297 42752
rect 7248 42712 7254 42724
rect 7285 42721 7297 42724
rect 7331 42721 7343 42755
rect 7285 42715 7343 42721
rect 8386 42712 8392 42764
rect 8444 42712 8450 42764
rect 8478 42712 8484 42764
rect 8536 42752 8542 42764
rect 8573 42755 8631 42761
rect 8573 42752 8585 42755
rect 8536 42724 8585 42752
rect 8536 42712 8542 42724
rect 8573 42721 8585 42724
rect 8619 42721 8631 42755
rect 8573 42715 8631 42721
rect 8662 42712 8668 42764
rect 8720 42712 8726 42764
rect 8757 42755 8815 42761
rect 8757 42721 8769 42755
rect 8803 42752 8815 42755
rect 8846 42752 8852 42764
rect 8803 42724 8852 42752
rect 8803 42721 8815 42724
rect 8757 42715 8815 42721
rect 8846 42712 8852 42724
rect 8904 42752 8910 42764
rect 9140 42752 9168 42860
rect 10597 42857 10609 42860
rect 10643 42857 10655 42891
rect 10597 42851 10655 42857
rect 10213 42823 10271 42829
rect 10213 42789 10225 42823
rect 10259 42820 10271 42823
rect 10318 42820 10324 42832
rect 10259 42792 10324 42820
rect 10259 42789 10271 42792
rect 10213 42783 10271 42789
rect 10318 42780 10324 42792
rect 10376 42780 10382 42832
rect 10413 42823 10471 42829
rect 10413 42789 10425 42823
rect 10459 42789 10471 42823
rect 10413 42783 10471 42789
rect 8904 42724 9168 42752
rect 8904 42712 8910 42724
rect 9214 42712 9220 42764
rect 9272 42712 9278 42764
rect 9401 42755 9459 42761
rect 9401 42721 9413 42755
rect 9447 42752 9459 42755
rect 9493 42755 9551 42761
rect 9493 42752 9505 42755
rect 9447 42724 9505 42752
rect 9447 42721 9459 42724
rect 9401 42715 9459 42721
rect 9493 42721 9505 42724
rect 9539 42721 9551 42755
rect 9493 42715 9551 42721
rect 9677 42755 9735 42761
rect 9677 42721 9689 42755
rect 9723 42721 9735 42755
rect 10428 42752 10456 42783
rect 10502 42780 10508 42832
rect 10560 42820 10566 42832
rect 10689 42823 10747 42829
rect 10689 42820 10701 42823
rect 10560 42792 10701 42820
rect 10560 42780 10566 42792
rect 10689 42789 10701 42792
rect 10735 42789 10747 42823
rect 10689 42783 10747 42789
rect 10594 42752 10600 42764
rect 10428 42724 10600 42752
rect 9677 42715 9735 42721
rect 6104 42656 6408 42684
rect 6457 42687 6515 42693
rect 5445 42647 5503 42653
rect 6457 42653 6469 42687
rect 6503 42653 6515 42687
rect 6457 42647 6515 42653
rect 4338 42616 4344 42628
rect 3344 42588 4344 42616
rect 2188 42576 2194 42588
rect 4338 42576 4344 42588
rect 4396 42576 4402 42628
rect 4798 42576 4804 42628
rect 4856 42616 4862 42628
rect 5460 42616 5488 42647
rect 4856 42588 5488 42616
rect 4856 42576 4862 42588
rect 5810 42576 5816 42628
rect 5868 42576 5874 42628
rect 6178 42576 6184 42628
rect 6236 42616 6242 42628
rect 6472 42616 6500 42647
rect 7006 42644 7012 42696
rect 7064 42684 7070 42696
rect 7561 42687 7619 42693
rect 7561 42684 7573 42687
rect 7064 42656 7573 42684
rect 7064 42644 7070 42656
rect 7561 42653 7573 42656
rect 7607 42653 7619 42687
rect 7561 42647 7619 42653
rect 7742 42644 7748 42696
rect 7800 42684 7806 42696
rect 9692 42684 9720 42715
rect 10594 42712 10600 42724
rect 10652 42712 10658 42764
rect 7800 42656 9720 42684
rect 7800 42644 7806 42656
rect 6236 42588 6500 42616
rect 6236 42576 6242 42588
rect 7650 42576 7656 42628
rect 7708 42616 7714 42628
rect 9585 42619 9643 42625
rect 9585 42616 9597 42619
rect 7708 42588 9597 42616
rect 7708 42576 7714 42588
rect 9585 42585 9597 42588
rect 9631 42585 9643 42619
rect 9585 42579 9643 42585
rect 9766 42576 9772 42628
rect 9824 42616 9830 42628
rect 9824 42588 10272 42616
rect 9824 42576 9830 42588
rect 2498 42548 2504 42560
rect 2056 42520 2504 42548
rect 2498 42508 2504 42520
rect 2556 42508 2562 42560
rect 4890 42508 4896 42560
rect 4948 42508 4954 42560
rect 5350 42508 5356 42560
rect 5408 42548 5414 42560
rect 8941 42551 8999 42557
rect 8941 42548 8953 42551
rect 5408 42520 8953 42548
rect 5408 42508 5414 42520
rect 8941 42517 8953 42520
rect 8987 42517 8999 42551
rect 8941 42511 8999 42517
rect 9030 42508 9036 42560
rect 9088 42548 9094 42560
rect 10244 42557 10272 42588
rect 10045 42551 10103 42557
rect 10045 42548 10057 42551
rect 9088 42520 10057 42548
rect 9088 42508 9094 42520
rect 10045 42517 10057 42520
rect 10091 42517 10103 42551
rect 10045 42511 10103 42517
rect 10229 42551 10287 42557
rect 10229 42517 10241 42551
rect 10275 42517 10287 42551
rect 10229 42511 10287 42517
rect 552 42458 11132 42480
rect 552 42406 3662 42458
rect 3714 42406 3726 42458
rect 3778 42406 3790 42458
rect 3842 42406 3854 42458
rect 3906 42406 3918 42458
rect 3970 42406 10062 42458
rect 10114 42406 10126 42458
rect 10178 42406 10190 42458
rect 10242 42406 10254 42458
rect 10306 42406 10318 42458
rect 10370 42406 11132 42458
rect 552 42384 11132 42406
rect 6546 42304 6552 42356
rect 6604 42344 6610 42356
rect 8386 42344 8392 42356
rect 6604 42316 8392 42344
rect 6604 42304 6610 42316
rect 8386 42304 8392 42316
rect 8444 42304 8450 42356
rect 8662 42304 8668 42356
rect 8720 42344 8726 42356
rect 9122 42344 9128 42356
rect 8720 42316 9128 42344
rect 8720 42304 8726 42316
rect 9122 42304 9128 42316
rect 9180 42304 9186 42356
rect 6825 42279 6883 42285
rect 6825 42245 6837 42279
rect 6871 42276 6883 42279
rect 9769 42279 9827 42285
rect 6871 42248 7420 42276
rect 6871 42245 6883 42248
rect 6825 42239 6883 42245
rect 2777 42211 2835 42217
rect 2777 42177 2789 42211
rect 2823 42208 2835 42211
rect 2958 42208 2964 42220
rect 2823 42180 2964 42208
rect 2823 42177 2835 42180
rect 2777 42171 2835 42177
rect 2958 42168 2964 42180
rect 3016 42168 3022 42220
rect 6086 42168 6092 42220
rect 6144 42168 6150 42220
rect 7392 42152 7420 42248
rect 9769 42245 9781 42279
rect 9815 42276 9827 42279
rect 10502 42276 10508 42288
rect 9815 42248 10508 42276
rect 9815 42245 9827 42248
rect 9769 42239 9827 42245
rect 10502 42236 10508 42248
rect 10560 42236 10566 42288
rect 7561 42211 7619 42217
rect 7561 42177 7573 42211
rect 7607 42208 7619 42211
rect 7650 42208 7656 42220
rect 7607 42180 7656 42208
rect 7607 42177 7619 42180
rect 7561 42171 7619 42177
rect 7650 42168 7656 42180
rect 7708 42168 7714 42220
rect 8110 42168 8116 42220
rect 8168 42208 8174 42220
rect 8168 42180 8524 42208
rect 8168 42168 8174 42180
rect 1210 42100 1216 42152
rect 1268 42100 1274 42152
rect 1305 42143 1363 42149
rect 1305 42109 1317 42143
rect 1351 42140 1363 42143
rect 1394 42140 1400 42152
rect 1351 42112 1400 42140
rect 1351 42109 1363 42112
rect 1305 42103 1363 42109
rect 1394 42100 1400 42112
rect 1452 42100 1458 42152
rect 1578 42149 1584 42152
rect 1572 42140 1584 42149
rect 1539 42112 1584 42140
rect 1572 42103 1584 42112
rect 1578 42100 1584 42103
rect 1636 42100 1642 42152
rect 2866 42100 2872 42152
rect 2924 42140 2930 42152
rect 3237 42143 3295 42149
rect 3237 42140 3249 42143
rect 2924 42112 3249 42140
rect 2924 42100 2930 42112
rect 3237 42109 3249 42112
rect 3283 42109 3295 42143
rect 3237 42103 3295 42109
rect 3694 42100 3700 42152
rect 3752 42140 3758 42152
rect 4985 42143 5043 42149
rect 4985 42140 4997 42143
rect 3752 42112 4997 42140
rect 3752 42100 3758 42112
rect 4985 42109 4997 42112
rect 5031 42109 5043 42143
rect 4985 42103 5043 42109
rect 5629 42143 5687 42149
rect 5629 42109 5641 42143
rect 5675 42109 5687 42143
rect 5629 42103 5687 42109
rect 2961 42075 3019 42081
rect 2961 42041 2973 42075
rect 3007 42072 3019 42075
rect 4154 42072 4160 42084
rect 3007 42044 4160 42072
rect 3007 42041 3019 42044
rect 2961 42035 3019 42041
rect 4154 42032 4160 42044
rect 4212 42032 4218 42084
rect 4740 42075 4798 42081
rect 4740 42041 4752 42075
rect 4786 42072 4798 42075
rect 4890 42072 4896 42084
rect 4786 42044 4896 42072
rect 4786 42041 4798 42044
rect 4740 42035 4798 42041
rect 4890 42032 4896 42044
rect 4948 42032 4954 42084
rect 566 41964 572 42016
rect 624 42004 630 42016
rect 1029 42007 1087 42013
rect 1029 42004 1041 42007
rect 624 41976 1041 42004
rect 624 41964 630 41976
rect 1029 41973 1041 41976
rect 1075 41973 1087 42007
rect 1029 41967 1087 41973
rect 2685 42007 2743 42013
rect 2685 41973 2697 42007
rect 2731 42004 2743 42007
rect 2774 42004 2780 42016
rect 2731 41976 2780 42004
rect 2731 41973 2743 41976
rect 2685 41967 2743 41973
rect 2774 41964 2780 41976
rect 2832 41964 2838 42016
rect 3050 41964 3056 42016
rect 3108 42004 3114 42016
rect 3421 42007 3479 42013
rect 3421 42004 3433 42007
rect 3108 41976 3433 42004
rect 3108 41964 3114 41976
rect 3421 41973 3433 41976
rect 3467 41973 3479 42007
rect 3421 41967 3479 41973
rect 3605 42007 3663 42013
rect 3605 41973 3617 42007
rect 3651 42004 3663 42007
rect 4338 42004 4344 42016
rect 3651 41976 4344 42004
rect 3651 41973 3663 41976
rect 3605 41967 3663 41973
rect 4338 41964 4344 41976
rect 4396 41964 4402 42016
rect 5074 41964 5080 42016
rect 5132 41964 5138 42016
rect 5644 42004 5672 42103
rect 5994 42100 6000 42152
rect 6052 42140 6058 42152
rect 6181 42143 6239 42149
rect 6181 42140 6193 42143
rect 6052 42112 6193 42140
rect 6052 42100 6058 42112
rect 6181 42109 6193 42112
rect 6227 42109 6239 42143
rect 7101 42143 7159 42149
rect 7101 42140 7113 42143
rect 6181 42103 6239 42109
rect 6886 42112 7113 42140
rect 5718 42032 5724 42084
rect 5776 42072 5782 42084
rect 6886 42072 6914 42112
rect 7101 42109 7113 42112
rect 7147 42109 7159 42143
rect 7101 42103 7159 42109
rect 7374 42100 7380 42152
rect 7432 42100 7438 42152
rect 8386 42100 8392 42152
rect 8444 42100 8450 42152
rect 8496 42140 8524 42180
rect 9674 42168 9680 42220
rect 9732 42208 9738 42220
rect 10594 42208 10600 42220
rect 9732 42180 10600 42208
rect 9732 42168 9738 42180
rect 10594 42168 10600 42180
rect 10652 42168 10658 42220
rect 9692 42140 9720 42168
rect 8496 42112 9720 42140
rect 5776 42044 6914 42072
rect 5776 42032 5782 42044
rect 7558 42032 7564 42084
rect 7616 42072 7622 42084
rect 7653 42075 7711 42081
rect 7653 42072 7665 42075
rect 7616 42044 7665 42072
rect 7616 42032 7622 42044
rect 7653 42041 7665 42044
rect 7699 42041 7711 42075
rect 7653 42035 7711 42041
rect 7742 42032 7748 42084
rect 7800 42032 7806 42084
rect 8662 42081 8668 42084
rect 7837 42075 7895 42081
rect 7837 42041 7849 42075
rect 7883 42041 7895 42075
rect 7837 42035 7895 42041
rect 8021 42075 8079 42081
rect 8021 42041 8033 42075
rect 8067 42072 8079 42075
rect 8067 42044 8622 42072
rect 8067 42041 8079 42044
rect 8021 42035 8079 42041
rect 6454 42004 6460 42016
rect 5644 41976 6460 42004
rect 6454 41964 6460 41976
rect 6512 42004 6518 42016
rect 7852 42004 7880 42035
rect 6512 41976 7880 42004
rect 6512 41964 6518 41976
rect 8202 41964 8208 42016
rect 8260 41964 8266 42016
rect 8594 42004 8622 42044
rect 8656 42035 8668 42081
rect 8662 42032 8668 42035
rect 8720 42032 8726 42084
rect 9766 42004 9772 42016
rect 8594 41976 9772 42004
rect 9766 41964 9772 41976
rect 9824 41964 9830 42016
rect 9950 41964 9956 42016
rect 10008 41964 10014 42016
rect 552 41914 11132 41936
rect 552 41862 4322 41914
rect 4374 41862 4386 41914
rect 4438 41862 4450 41914
rect 4502 41862 4514 41914
rect 4566 41862 4578 41914
rect 4630 41862 10722 41914
rect 10774 41862 10786 41914
rect 10838 41862 10850 41914
rect 10902 41862 10914 41914
rect 10966 41862 10978 41914
rect 11030 41862 11132 41914
rect 552 41840 11132 41862
rect 3694 41800 3700 41812
rect 2746 41772 3700 41800
rect 1394 41732 1400 41744
rect 1320 41704 1400 41732
rect 1118 41624 1124 41676
rect 1176 41664 1182 41676
rect 1320 41673 1348 41704
rect 1394 41692 1400 41704
rect 1452 41732 1458 41744
rect 2222 41732 2228 41744
rect 1452 41704 2228 41732
rect 1452 41692 1458 41704
rect 2222 41692 2228 41704
rect 2280 41732 2286 41744
rect 2746 41732 2774 41772
rect 3694 41760 3700 41772
rect 3752 41760 3758 41812
rect 8110 41800 8116 41812
rect 5460 41772 8116 41800
rect 2280 41704 2774 41732
rect 2280 41692 2286 41704
rect 3326 41692 3332 41744
rect 3384 41732 3390 41744
rect 3942 41735 4000 41741
rect 3942 41732 3954 41735
rect 3384 41704 3954 41732
rect 3384 41692 3390 41704
rect 3942 41701 3954 41704
rect 3988 41701 4000 41735
rect 5350 41732 5356 41744
rect 3942 41695 4000 41701
rect 5092 41704 5356 41732
rect 1213 41667 1271 41673
rect 1213 41664 1225 41667
rect 1176 41636 1225 41664
rect 1176 41624 1182 41636
rect 1213 41633 1225 41636
rect 1259 41633 1271 41667
rect 1213 41627 1271 41633
rect 1305 41667 1363 41673
rect 1305 41633 1317 41667
rect 1351 41633 1363 41667
rect 1561 41667 1619 41673
rect 1561 41664 1573 41667
rect 1305 41627 1363 41633
rect 1412 41636 1573 41664
rect 750 41556 756 41608
rect 808 41596 814 41608
rect 1412 41596 1440 41636
rect 1561 41633 1573 41636
rect 1607 41633 1619 41667
rect 1561 41627 1619 41633
rect 3234 41624 3240 41676
rect 3292 41624 3298 41676
rect 3694 41624 3700 41676
rect 3752 41624 3758 41676
rect 5092 41664 5120 41704
rect 5350 41692 5356 41704
rect 5408 41692 5414 41744
rect 5460 41741 5488 41772
rect 8110 41760 8116 41772
rect 8168 41760 8174 41812
rect 8386 41760 8392 41812
rect 8444 41800 8450 41812
rect 8444 41772 9536 41800
rect 8444 41760 8450 41772
rect 9508 41744 9536 41772
rect 9766 41760 9772 41812
rect 9824 41800 9830 41812
rect 10686 41800 10692 41812
rect 9824 41772 10692 41800
rect 9824 41760 9830 41772
rect 10686 41760 10692 41772
rect 10744 41760 10750 41812
rect 5445 41735 5503 41741
rect 5445 41701 5457 41735
rect 5491 41701 5503 41735
rect 5445 41695 5503 41701
rect 5629 41735 5687 41741
rect 5629 41701 5641 41735
rect 5675 41732 5687 41735
rect 5675 41704 6040 41732
rect 5675 41701 5687 41704
rect 5629 41695 5687 41701
rect 6012 41676 6040 41704
rect 6638 41692 6644 41744
rect 6696 41692 6702 41744
rect 7650 41692 7656 41744
rect 7708 41732 7714 41744
rect 9030 41732 9036 41744
rect 7708 41704 7788 41732
rect 7708 41692 7714 41704
rect 3804 41636 5120 41664
rect 808 41568 1440 41596
rect 3053 41599 3111 41605
rect 808 41556 814 41568
rect 3053 41565 3065 41599
rect 3099 41565 3111 41599
rect 3053 41559 3111 41565
rect 3145 41599 3203 41605
rect 3145 41565 3157 41599
rect 3191 41596 3203 41599
rect 3804 41596 3832 41636
rect 5166 41624 5172 41676
rect 5224 41664 5230 41676
rect 5261 41667 5319 41673
rect 5261 41664 5273 41667
rect 5224 41636 5273 41664
rect 5224 41624 5230 41636
rect 5261 41633 5273 41636
rect 5307 41633 5319 41667
rect 5261 41627 5319 41633
rect 5718 41624 5724 41676
rect 5776 41664 5782 41676
rect 5813 41667 5871 41673
rect 5813 41664 5825 41667
rect 5776 41636 5825 41664
rect 5776 41624 5782 41636
rect 5813 41633 5825 41636
rect 5859 41633 5871 41667
rect 5813 41627 5871 41633
rect 5994 41624 6000 41676
rect 6052 41624 6058 41676
rect 7374 41624 7380 41676
rect 7432 41624 7438 41676
rect 7760 41673 7788 41704
rect 8128 41704 9036 41732
rect 7745 41667 7803 41673
rect 7745 41633 7757 41667
rect 7791 41633 7803 41667
rect 7745 41627 7803 41633
rect 7834 41624 7840 41676
rect 7892 41664 7898 41676
rect 8128 41673 8156 41704
rect 9030 41692 9036 41704
rect 9088 41692 9094 41744
rect 9490 41692 9496 41744
rect 9548 41732 9554 41744
rect 10413 41735 10471 41741
rect 9548 41704 10088 41732
rect 9548 41692 9554 41704
rect 8113 41667 8171 41673
rect 8113 41664 8125 41667
rect 7892 41636 8125 41664
rect 7892 41624 7898 41636
rect 8113 41633 8125 41636
rect 8159 41633 8171 41667
rect 8113 41627 8171 41633
rect 8205 41667 8263 41673
rect 8205 41633 8217 41667
rect 8251 41664 8263 41667
rect 8251 41636 8340 41664
rect 8251 41633 8263 41636
rect 8205 41627 8263 41633
rect 3191 41568 3832 41596
rect 8312 41596 8340 41636
rect 8386 41624 8392 41676
rect 8444 41624 8450 41676
rect 9214 41664 9220 41676
rect 8496 41636 9220 41664
rect 8496 41596 8524 41636
rect 9214 41624 9220 41636
rect 9272 41624 9278 41676
rect 9766 41624 9772 41676
rect 9824 41673 9830 41676
rect 10060 41673 10088 41704
rect 10413 41701 10425 41735
rect 10459 41732 10471 41735
rect 11054 41732 11060 41744
rect 10459 41704 11060 41732
rect 10459 41701 10471 41704
rect 10413 41695 10471 41701
rect 11054 41692 11060 41704
rect 11112 41692 11118 41744
rect 9824 41627 9836 41673
rect 10045 41667 10103 41673
rect 10045 41633 10057 41667
rect 10091 41633 10103 41667
rect 10045 41627 10103 41633
rect 9824 41624 9830 41627
rect 10594 41624 10600 41676
rect 10652 41624 10658 41676
rect 8312 41568 8524 41596
rect 3191 41565 3203 41568
rect 3145 41559 3203 41565
rect 3068 41528 3096 41559
rect 5077 41531 5135 41537
rect 3068 41500 3740 41528
rect 1026 41420 1032 41472
rect 1084 41420 1090 41472
rect 1578 41420 1584 41472
rect 1636 41460 1642 41472
rect 2685 41463 2743 41469
rect 2685 41460 2697 41463
rect 1636 41432 2697 41460
rect 1636 41420 1642 41432
rect 2685 41429 2697 41432
rect 2731 41429 2743 41463
rect 2685 41423 2743 41429
rect 3418 41420 3424 41472
rect 3476 41460 3482 41472
rect 3605 41463 3663 41469
rect 3605 41460 3617 41463
rect 3476 41432 3617 41460
rect 3476 41420 3482 41432
rect 3605 41429 3617 41432
rect 3651 41429 3663 41463
rect 3712 41460 3740 41500
rect 5077 41497 5089 41531
rect 5123 41528 5135 41531
rect 6454 41528 6460 41540
rect 5123 41500 6460 41528
rect 5123 41497 5135 41500
rect 5077 41491 5135 41497
rect 6454 41488 6460 41500
rect 6512 41488 6518 41540
rect 4798 41460 4804 41472
rect 3712 41432 4804 41460
rect 3605 41423 3663 41429
rect 4798 41420 4804 41432
rect 4856 41420 4862 41472
rect 5902 41420 5908 41472
rect 5960 41420 5966 41472
rect 7650 41420 7656 41472
rect 7708 41460 7714 41472
rect 8496 41460 8524 41568
rect 8665 41531 8723 41537
rect 8665 41497 8677 41531
rect 8711 41528 8723 41531
rect 8754 41528 8760 41540
rect 8711 41500 8760 41528
rect 8711 41497 8723 41500
rect 8665 41491 8723 41497
rect 8754 41488 8760 41500
rect 8812 41488 8818 41540
rect 7708 41432 8524 41460
rect 7708 41420 7714 41432
rect 8570 41420 8576 41472
rect 8628 41420 8634 41472
rect 9858 41420 9864 41472
rect 9916 41460 9922 41472
rect 10229 41463 10287 41469
rect 10229 41460 10241 41463
rect 9916 41432 10241 41460
rect 9916 41420 9922 41432
rect 10229 41429 10241 41432
rect 10275 41429 10287 41463
rect 10229 41423 10287 41429
rect 552 41370 11132 41392
rect 552 41318 3662 41370
rect 3714 41318 3726 41370
rect 3778 41318 3790 41370
rect 3842 41318 3854 41370
rect 3906 41318 3918 41370
rect 3970 41318 10062 41370
rect 10114 41318 10126 41370
rect 10178 41318 10190 41370
rect 10242 41318 10254 41370
rect 10306 41318 10318 41370
rect 10370 41318 11132 41370
rect 552 41296 11132 41318
rect 1029 41259 1087 41265
rect 1029 41225 1041 41259
rect 1075 41256 1087 41259
rect 4706 41256 4712 41268
rect 1075 41228 4712 41256
rect 1075 41225 1087 41228
rect 1029 41219 1087 41225
rect 4706 41216 4712 41228
rect 4764 41216 4770 41268
rect 8478 41256 8484 41268
rect 6288 41228 8484 41256
rect 198 41148 204 41200
rect 256 41188 262 41200
rect 1486 41188 1492 41200
rect 256 41160 1492 41188
rect 256 41148 262 41160
rect 1486 41148 1492 41160
rect 1544 41148 1550 41200
rect 1670 41148 1676 41200
rect 1728 41148 1734 41200
rect 2682 41148 2688 41200
rect 2740 41188 2746 41200
rect 3421 41191 3479 41197
rect 3421 41188 3433 41191
rect 2740 41160 3433 41188
rect 2740 41148 2746 41160
rect 3421 41157 3433 41160
rect 3467 41157 3479 41191
rect 3421 41151 3479 41157
rect 4890 41148 4896 41200
rect 4948 41188 4954 41200
rect 6288 41188 6316 41228
rect 8478 41216 8484 41228
rect 8536 41216 8542 41268
rect 8846 41216 8852 41268
rect 8904 41256 8910 41268
rect 9030 41256 9036 41268
rect 8904 41228 9036 41256
rect 8904 41216 8910 41228
rect 9030 41216 9036 41228
rect 9088 41216 9094 41268
rect 9217 41259 9275 41265
rect 9217 41225 9229 41259
rect 9263 41256 9275 41259
rect 9674 41256 9680 41268
rect 9263 41228 9680 41256
rect 9263 41225 9275 41228
rect 9217 41219 9275 41225
rect 9674 41216 9680 41228
rect 9732 41216 9738 41268
rect 4948 41160 6316 41188
rect 4948 41148 4954 41160
rect 6730 41148 6736 41200
rect 6788 41188 6794 41200
rect 6825 41191 6883 41197
rect 6825 41188 6837 41191
rect 6788 41160 6837 41188
rect 6788 41148 6794 41160
rect 6825 41157 6837 41160
rect 6871 41157 6883 41191
rect 8570 41188 8576 41200
rect 6825 41151 6883 41157
rect 8404 41160 8576 41188
rect 1688 41120 1716 41148
rect 1228 41092 1716 41120
rect 1228 41061 1256 41092
rect 3510 41080 3516 41132
rect 3568 41120 3574 41132
rect 3697 41123 3755 41129
rect 3697 41120 3709 41123
rect 3568 41092 3709 41120
rect 3568 41080 3574 41092
rect 3697 41089 3709 41092
rect 3743 41089 3755 41123
rect 3697 41083 3755 41089
rect 6086 41080 6092 41132
rect 6144 41080 6150 41132
rect 8404 41064 8432 41160
rect 8570 41148 8576 41160
rect 8628 41148 8634 41200
rect 1213 41055 1271 41061
rect 1213 41021 1225 41055
rect 1259 41021 1271 41055
rect 1213 41015 1271 41021
rect 1578 41012 1584 41064
rect 1636 41012 1642 41064
rect 1673 41055 1731 41061
rect 1673 41021 1685 41055
rect 1719 41052 1731 41055
rect 2222 41052 2228 41064
rect 1719 41024 2228 41052
rect 1719 41021 1731 41024
rect 1673 41015 1731 41021
rect 2222 41012 2228 41024
rect 2280 41012 2286 41064
rect 2774 41012 2780 41064
rect 2832 41052 2838 41064
rect 3237 41055 3295 41061
rect 3237 41052 3249 41055
rect 2832 41024 3249 41052
rect 2832 41012 2838 41024
rect 3237 41021 3249 41024
rect 3283 41021 3295 41055
rect 3237 41015 3295 41021
rect 4982 41012 4988 41064
rect 5040 41052 5046 41064
rect 5353 41055 5411 41061
rect 5353 41052 5365 41055
rect 5040 41024 5365 41052
rect 5040 41012 5046 41024
rect 5353 41021 5365 41024
rect 5399 41021 5411 41055
rect 5353 41015 5411 41021
rect 5902 41012 5908 41064
rect 5960 41012 5966 41064
rect 8205 41055 8263 41061
rect 8205 41021 8217 41055
rect 8251 41052 8263 41055
rect 8294 41052 8300 41064
rect 8251 41024 8300 41052
rect 8251 41021 8263 41024
rect 8205 41015 8263 41021
rect 8294 41012 8300 41024
rect 8352 41012 8358 41064
rect 8386 41012 8392 41064
rect 8444 41012 8450 41064
rect 8570 41012 8576 41064
rect 8628 41012 8634 41064
rect 8754 41012 8760 41064
rect 8812 41012 8818 41064
rect 8846 41012 8852 41064
rect 8904 41012 8910 41064
rect 8941 41055 8999 41061
rect 8941 41021 8953 41055
rect 8987 41052 8999 41055
rect 9214 41052 9220 41064
rect 8987 41024 9220 41052
rect 8987 41021 8999 41024
rect 8941 41015 8999 41021
rect 9214 41012 9220 41024
rect 9272 41012 9278 41064
rect 9309 41055 9367 41061
rect 9309 41021 9321 41055
rect 9355 41052 9367 41055
rect 9398 41052 9404 41064
rect 9355 41024 9404 41052
rect 9355 41021 9367 41024
rect 9309 41015 9367 41021
rect 9398 41012 9404 41024
rect 9456 41012 9462 41064
rect 1305 40987 1363 40993
rect 1305 40953 1317 40987
rect 1351 40953 1363 40987
rect 1305 40947 1363 40953
rect 1397 40987 1455 40993
rect 1397 40953 1409 40987
rect 1443 40984 1455 40987
rect 1486 40984 1492 40996
rect 1443 40956 1492 40984
rect 1443 40953 1455 40956
rect 1397 40947 1455 40953
rect 382 40876 388 40928
rect 440 40916 446 40928
rect 658 40916 664 40928
rect 440 40888 664 40916
rect 440 40876 446 40888
rect 658 40876 664 40888
rect 716 40876 722 40928
rect 1320 40916 1348 40947
rect 1486 40944 1492 40956
rect 1544 40944 1550 40996
rect 1762 40944 1768 40996
rect 1820 40984 1826 40996
rect 1918 40987 1976 40993
rect 1918 40984 1930 40987
rect 1820 40956 1930 40984
rect 1820 40944 1826 40956
rect 1918 40953 1930 40956
rect 1964 40953 1976 40987
rect 3964 40987 4022 40993
rect 1918 40947 1976 40953
rect 3068 40956 3924 40984
rect 2038 40916 2044 40928
rect 1320 40888 2044 40916
rect 2038 40876 2044 40888
rect 2096 40876 2102 40928
rect 3068 40925 3096 40956
rect 3053 40919 3111 40925
rect 3053 40885 3065 40919
rect 3099 40885 3111 40919
rect 3896 40916 3924 40956
rect 3964 40953 3976 40987
rect 4010 40984 4022 40987
rect 4062 40984 4068 40996
rect 4010 40956 4068 40984
rect 4010 40953 4022 40956
rect 3964 40947 4022 40953
rect 4062 40944 4068 40956
rect 4120 40944 4126 40996
rect 7926 40944 7932 40996
rect 7984 40993 7990 40996
rect 7984 40947 7996 40993
rect 9576 40987 9634 40993
rect 9576 40953 9588 40987
rect 9622 40984 9634 40987
rect 10134 40984 10140 40996
rect 9622 40956 10140 40984
rect 9622 40953 9634 40956
rect 9576 40947 9634 40953
rect 7984 40944 7990 40947
rect 10134 40944 10140 40956
rect 10192 40944 10198 40996
rect 4890 40916 4896 40928
rect 3896 40888 4896 40916
rect 3053 40879 3111 40885
rect 4890 40876 4896 40888
rect 4948 40876 4954 40928
rect 4982 40876 4988 40928
rect 5040 40916 5046 40928
rect 5077 40919 5135 40925
rect 5077 40916 5089 40919
rect 5040 40888 5089 40916
rect 5040 40876 5046 40888
rect 5077 40885 5089 40888
rect 5123 40916 5135 40919
rect 5166 40916 5172 40928
rect 5123 40888 5172 40916
rect 5123 40885 5135 40888
rect 5077 40879 5135 40885
rect 5166 40876 5172 40888
rect 5224 40876 5230 40928
rect 5258 40876 5264 40928
rect 5316 40876 5322 40928
rect 5350 40876 5356 40928
rect 5408 40916 5414 40928
rect 6546 40916 6552 40928
rect 5408 40888 6552 40916
rect 5408 40876 5414 40888
rect 6546 40876 6552 40888
rect 6604 40876 6610 40928
rect 6638 40876 6644 40928
rect 6696 40876 6702 40928
rect 10318 40876 10324 40928
rect 10376 40916 10382 40928
rect 10686 40916 10692 40928
rect 10376 40888 10692 40916
rect 10376 40876 10382 40888
rect 10686 40876 10692 40888
rect 10744 40876 10750 40928
rect 552 40826 11132 40848
rect 552 40774 4322 40826
rect 4374 40774 4386 40826
rect 4438 40774 4450 40826
rect 4502 40774 4514 40826
rect 4566 40774 4578 40826
rect 4630 40774 10722 40826
rect 10774 40774 10786 40826
rect 10838 40774 10850 40826
rect 10902 40774 10914 40826
rect 10966 40774 10978 40826
rect 11030 40774 11132 40826
rect 552 40752 11132 40774
rect 658 40672 664 40724
rect 716 40712 722 40724
rect 716 40684 2084 40712
rect 716 40672 722 40684
rect 2056 40644 2084 40684
rect 3234 40672 3240 40724
rect 3292 40712 3298 40724
rect 3329 40715 3387 40721
rect 3329 40712 3341 40715
rect 3292 40684 3341 40712
rect 3292 40672 3298 40684
rect 3329 40681 3341 40684
rect 3375 40681 3387 40715
rect 3329 40675 3387 40681
rect 4433 40715 4491 40721
rect 4433 40681 4445 40715
rect 4479 40712 4491 40715
rect 5074 40712 5080 40724
rect 4479 40684 5080 40712
rect 4479 40681 4491 40684
rect 4433 40675 4491 40681
rect 5074 40672 5080 40684
rect 5132 40672 5138 40724
rect 5445 40715 5503 40721
rect 5445 40681 5457 40715
rect 5491 40712 5503 40715
rect 6086 40712 6092 40724
rect 5491 40684 6092 40712
rect 5491 40681 5503 40684
rect 5445 40675 5503 40681
rect 6086 40672 6092 40684
rect 6144 40672 6150 40724
rect 6546 40672 6552 40724
rect 6604 40712 6610 40724
rect 7209 40715 7267 40721
rect 7209 40712 7221 40715
rect 6604 40684 7221 40712
rect 6604 40672 6610 40684
rect 7209 40681 7221 40684
rect 7255 40712 7267 40715
rect 7834 40712 7840 40724
rect 7255 40684 7840 40712
rect 7255 40681 7267 40684
rect 7209 40675 7267 40681
rect 7834 40672 7840 40684
rect 7892 40672 7898 40724
rect 7926 40672 7932 40724
rect 7984 40672 7990 40724
rect 8478 40712 8484 40724
rect 8312 40684 8484 40712
rect 2056 40616 6040 40644
rect 1121 40579 1179 40585
rect 1121 40545 1133 40579
rect 1167 40576 1179 40579
rect 1302 40576 1308 40588
rect 1167 40548 1308 40576
rect 1167 40545 1179 40548
rect 1121 40539 1179 40545
rect 1302 40536 1308 40548
rect 1360 40536 1366 40588
rect 1486 40536 1492 40588
rect 1544 40536 1550 40588
rect 1670 40536 1676 40588
rect 1728 40576 1734 40588
rect 1837 40579 1895 40585
rect 1837 40576 1849 40579
rect 1728 40548 1849 40576
rect 1728 40536 1734 40548
rect 1837 40545 1849 40548
rect 1883 40545 1895 40579
rect 1837 40539 1895 40545
rect 3053 40579 3111 40585
rect 3053 40545 3065 40579
rect 3099 40576 3111 40579
rect 3234 40576 3240 40588
rect 3099 40548 3240 40576
rect 3099 40545 3111 40548
rect 3053 40539 3111 40545
rect 3234 40536 3240 40548
rect 3292 40536 3298 40588
rect 4982 40576 4988 40588
rect 3896 40548 4988 40576
rect 1394 40468 1400 40520
rect 1452 40508 1458 40520
rect 1581 40511 1639 40517
rect 1581 40508 1593 40511
rect 1452 40480 1593 40508
rect 1452 40468 1458 40480
rect 1581 40477 1593 40480
rect 1627 40477 1639 40511
rect 1581 40471 1639 40477
rect 3510 40468 3516 40520
rect 3568 40508 3574 40520
rect 3896 40517 3924 40548
rect 4982 40536 4988 40548
rect 5040 40536 5046 40588
rect 5074 40536 5080 40588
rect 5132 40576 5138 40588
rect 5445 40579 5503 40585
rect 5445 40576 5457 40579
rect 5132 40548 5457 40576
rect 5132 40536 5138 40548
rect 5445 40545 5457 40548
rect 5491 40545 5503 40579
rect 6012 40562 6040 40616
rect 6178 40604 6184 40656
rect 6236 40644 6242 40656
rect 6641 40647 6699 40653
rect 6641 40644 6653 40647
rect 6236 40616 6653 40644
rect 6236 40604 6242 40616
rect 6641 40613 6653 40616
rect 6687 40613 6699 40647
rect 6641 40607 6699 40613
rect 7009 40647 7067 40653
rect 7009 40613 7021 40647
rect 7055 40644 7067 40647
rect 8312 40644 8340 40684
rect 8478 40672 8484 40684
rect 8536 40672 8542 40724
rect 8573 40715 8631 40721
rect 8573 40681 8585 40715
rect 8619 40712 8631 40715
rect 8662 40712 8668 40724
rect 8619 40684 8668 40712
rect 8619 40681 8631 40684
rect 8573 40675 8631 40681
rect 8662 40672 8668 40684
rect 8720 40672 8726 40724
rect 8938 40672 8944 40724
rect 8996 40712 9002 40724
rect 9398 40712 9404 40724
rect 8996 40684 9404 40712
rect 8996 40672 9002 40684
rect 9398 40672 9404 40684
rect 9456 40672 9462 40724
rect 10134 40672 10140 40724
rect 10192 40672 10198 40724
rect 7055 40616 8340 40644
rect 7055 40613 7067 40616
rect 7009 40607 7067 40613
rect 8386 40604 8392 40656
rect 8444 40604 8450 40656
rect 8588 40616 9076 40644
rect 5445 40539 5503 40545
rect 6730 40536 6736 40588
rect 6788 40576 6794 40588
rect 7469 40579 7527 40585
rect 7469 40576 7481 40579
rect 6788 40548 7481 40576
rect 6788 40536 6794 40548
rect 7469 40545 7481 40548
rect 7515 40545 7527 40579
rect 7469 40539 7527 40545
rect 7745 40579 7803 40585
rect 7745 40545 7757 40579
rect 7791 40576 7803 40579
rect 8294 40576 8300 40588
rect 7791 40548 8300 40576
rect 7791 40545 7803 40548
rect 7745 40539 7803 40545
rect 8294 40536 8300 40548
rect 8352 40536 8358 40588
rect 8478 40536 8484 40588
rect 8536 40576 8542 40588
rect 8588 40576 8616 40616
rect 8536 40548 8616 40576
rect 8536 40536 8542 40548
rect 8662 40536 8668 40588
rect 8720 40536 8726 40588
rect 8938 40585 8944 40588
rect 8932 40539 8944 40585
rect 8938 40536 8944 40539
rect 8996 40536 9002 40588
rect 9048 40576 9076 40616
rect 9122 40604 9128 40656
rect 9180 40644 9186 40656
rect 9180 40616 10824 40644
rect 9180 40604 9186 40616
rect 10134 40576 10140 40588
rect 9048 40548 10140 40576
rect 10134 40536 10140 40548
rect 10192 40536 10198 40588
rect 10318 40576 10324 40588
rect 10244 40548 10324 40576
rect 3881 40511 3939 40517
rect 3881 40508 3893 40511
rect 3568 40480 3893 40508
rect 3568 40468 3574 40480
rect 3881 40477 3893 40480
rect 3927 40477 3939 40511
rect 3881 40471 3939 40477
rect 4522 40468 4528 40520
rect 4580 40468 4586 40520
rect 4709 40511 4767 40517
rect 4709 40477 4721 40511
rect 4755 40508 4767 40511
rect 4798 40508 4804 40520
rect 4755 40480 4804 40508
rect 4755 40477 4767 40480
rect 4709 40471 4767 40477
rect 4798 40468 4804 40480
rect 4856 40468 4862 40520
rect 4890 40468 4896 40520
rect 4948 40468 4954 40520
rect 5537 40511 5595 40517
rect 5537 40477 5549 40511
rect 5583 40508 5595 40511
rect 5810 40508 5816 40520
rect 5583 40480 5816 40508
rect 5583 40477 5595 40480
rect 5537 40471 5595 40477
rect 5810 40468 5816 40480
rect 5868 40508 5874 40520
rect 6089 40511 6147 40517
rect 6089 40508 6101 40511
rect 5868 40480 6101 40508
rect 5868 40468 5874 40480
rect 6089 40477 6101 40480
rect 6135 40477 6147 40511
rect 6089 40471 6147 40477
rect 7561 40511 7619 40517
rect 7561 40477 7573 40511
rect 7607 40508 7619 40511
rect 8021 40511 8079 40517
rect 8021 40508 8033 40511
rect 7607 40480 8033 40508
rect 7607 40477 7619 40480
rect 7561 40471 7619 40477
rect 8021 40477 8033 40480
rect 8067 40508 8079 40511
rect 8386 40508 8392 40520
rect 8067 40480 8392 40508
rect 8067 40477 8079 40480
rect 8021 40471 8079 40477
rect 2590 40400 2596 40452
rect 2648 40440 2654 40452
rect 2866 40440 2872 40452
rect 2648 40412 2872 40440
rect 2648 40400 2654 40412
rect 2866 40400 2872 40412
rect 2924 40400 2930 40452
rect 5626 40400 5632 40452
rect 5684 40440 5690 40452
rect 7377 40443 7435 40449
rect 5684 40412 7236 40440
rect 5684 40400 5690 40412
rect 934 40332 940 40384
rect 992 40332 998 40384
rect 1302 40332 1308 40384
rect 1360 40332 1366 40384
rect 1854 40332 1860 40384
rect 1912 40372 1918 40384
rect 2961 40375 3019 40381
rect 2961 40372 2973 40375
rect 1912 40344 2973 40372
rect 1912 40332 1918 40344
rect 2961 40341 2973 40344
rect 3007 40341 3019 40375
rect 2961 40335 3019 40341
rect 3050 40332 3056 40384
rect 3108 40372 3114 40384
rect 3145 40375 3203 40381
rect 3145 40372 3157 40375
rect 3108 40344 3157 40372
rect 3108 40332 3114 40344
rect 3145 40341 3157 40344
rect 3191 40341 3203 40375
rect 3145 40335 3203 40341
rect 4065 40375 4123 40381
rect 4065 40341 4077 40375
rect 4111 40372 4123 40375
rect 4614 40372 4620 40384
rect 4111 40344 4620 40372
rect 4111 40341 4123 40344
rect 4065 40335 4123 40341
rect 4614 40332 4620 40344
rect 4672 40332 4678 40384
rect 7208 40381 7236 40412
rect 7377 40409 7389 40443
rect 7423 40440 7435 40443
rect 7576 40440 7604 40471
rect 8386 40468 8392 40480
rect 8444 40468 8450 40520
rect 9674 40468 9680 40520
rect 9732 40508 9738 40520
rect 10244 40508 10272 40548
rect 10318 40536 10324 40548
rect 10376 40576 10382 40588
rect 10413 40579 10471 40585
rect 10413 40576 10425 40579
rect 10376 40548 10425 40576
rect 10376 40536 10382 40548
rect 10413 40545 10425 40548
rect 10459 40545 10471 40579
rect 10413 40539 10471 40545
rect 10505 40579 10563 40585
rect 10505 40545 10517 40579
rect 10551 40545 10563 40579
rect 10505 40539 10563 40545
rect 10597 40579 10655 40585
rect 10597 40545 10609 40579
rect 10643 40576 10655 40579
rect 10686 40576 10692 40588
rect 10643 40548 10692 40576
rect 10643 40545 10655 40548
rect 10597 40539 10655 40545
rect 10520 40508 10548 40539
rect 10686 40536 10692 40548
rect 10744 40536 10750 40588
rect 10796 40585 10824 40616
rect 10781 40579 10839 40585
rect 10781 40545 10793 40579
rect 10827 40545 10839 40579
rect 10781 40539 10839 40545
rect 9732 40480 10272 40508
rect 10428 40480 10548 40508
rect 9732 40468 9738 40480
rect 10428 40452 10456 40480
rect 7423 40412 7604 40440
rect 7423 40409 7435 40412
rect 7377 40403 7435 40409
rect 10410 40400 10416 40452
rect 10468 40400 10474 40452
rect 7193 40375 7251 40381
rect 7193 40341 7205 40375
rect 7239 40372 7251 40375
rect 8018 40372 8024 40384
rect 7239 40344 8024 40372
rect 7239 40341 7251 40344
rect 7193 40335 7251 40341
rect 8018 40332 8024 40344
rect 8076 40332 8082 40384
rect 8389 40375 8447 40381
rect 8389 40341 8401 40375
rect 8435 40372 8447 40375
rect 8570 40372 8576 40384
rect 8435 40344 8576 40372
rect 8435 40341 8447 40344
rect 8389 40335 8447 40341
rect 8570 40332 8576 40344
rect 8628 40372 8634 40384
rect 9030 40372 9036 40384
rect 8628 40344 9036 40372
rect 8628 40332 8634 40344
rect 9030 40332 9036 40344
rect 9088 40332 9094 40384
rect 9582 40332 9588 40384
rect 9640 40372 9646 40384
rect 10045 40375 10103 40381
rect 10045 40372 10057 40375
rect 9640 40344 10057 40372
rect 9640 40332 9646 40344
rect 10045 40341 10057 40344
rect 10091 40341 10103 40375
rect 10045 40335 10103 40341
rect 10134 40332 10140 40384
rect 10192 40372 10198 40384
rect 10502 40372 10508 40384
rect 10192 40344 10508 40372
rect 10192 40332 10198 40344
rect 10502 40332 10508 40344
rect 10560 40332 10566 40384
rect 552 40282 11132 40304
rect 552 40230 3662 40282
rect 3714 40230 3726 40282
rect 3778 40230 3790 40282
rect 3842 40230 3854 40282
rect 3906 40230 3918 40282
rect 3970 40230 10062 40282
rect 10114 40230 10126 40282
rect 10178 40230 10190 40282
rect 10242 40230 10254 40282
rect 10306 40230 10318 40282
rect 10370 40230 11132 40282
rect 552 40208 11132 40230
rect 1489 40171 1547 40177
rect 1489 40137 1501 40171
rect 1535 40168 1547 40171
rect 2590 40168 2596 40180
rect 1535 40140 2596 40168
rect 1535 40137 1547 40140
rect 1489 40131 1547 40137
rect 2590 40128 2596 40140
rect 2648 40128 2654 40180
rect 3050 40128 3056 40180
rect 3108 40168 3114 40180
rect 3694 40168 3700 40180
rect 3108 40140 3700 40168
rect 3108 40128 3114 40140
rect 3694 40128 3700 40140
rect 3752 40128 3758 40180
rect 3973 40171 4031 40177
rect 3973 40137 3985 40171
rect 4019 40168 4031 40171
rect 4062 40168 4068 40180
rect 4019 40140 4068 40168
rect 4019 40137 4031 40140
rect 3973 40131 4031 40137
rect 4062 40128 4068 40140
rect 4120 40128 4126 40180
rect 4890 40128 4896 40180
rect 4948 40168 4954 40180
rect 8202 40168 8208 40180
rect 4948 40140 8208 40168
rect 4948 40128 4954 40140
rect 8202 40128 8208 40140
rect 8260 40128 8266 40180
rect 8294 40128 8300 40180
rect 8352 40168 8358 40180
rect 8665 40171 8723 40177
rect 8665 40168 8677 40171
rect 8352 40140 8677 40168
rect 8352 40128 8358 40140
rect 8665 40137 8677 40140
rect 8711 40137 8723 40171
rect 8665 40131 8723 40137
rect 8846 40128 8852 40180
rect 8904 40168 8910 40180
rect 9033 40171 9091 40177
rect 9033 40168 9045 40171
rect 8904 40140 9045 40168
rect 8904 40128 8910 40140
rect 9033 40137 9045 40140
rect 9079 40137 9091 40171
rect 9033 40131 9091 40137
rect 9217 40171 9275 40177
rect 9217 40137 9229 40171
rect 9263 40168 9275 40171
rect 9398 40168 9404 40180
rect 9263 40140 9404 40168
rect 9263 40137 9275 40140
rect 9217 40131 9275 40137
rect 9398 40128 9404 40140
rect 9456 40128 9462 40180
rect 9769 40171 9827 40177
rect 9769 40137 9781 40171
rect 9815 40137 9827 40171
rect 9769 40131 9827 40137
rect 2038 40060 2044 40112
rect 2096 40100 2102 40112
rect 3234 40100 3240 40112
rect 2096 40072 3240 40100
rect 2096 40060 2102 40072
rect 3234 40060 3240 40072
rect 3292 40060 3298 40112
rect 5721 40103 5779 40109
rect 3344 40072 3556 40100
rect 1305 40035 1363 40041
rect 1305 40001 1317 40035
rect 1351 40032 1363 40035
rect 1351 40004 2774 40032
rect 1351 40001 1363 40004
rect 1305 39995 1363 40001
rect 1213 39967 1271 39973
rect 1213 39933 1225 39967
rect 1259 39933 1271 39967
rect 1213 39927 1271 39933
rect 1228 39896 1256 39927
rect 1578 39924 1584 39976
rect 1636 39964 1642 39976
rect 1673 39967 1731 39973
rect 1673 39964 1685 39967
rect 1636 39936 1685 39964
rect 1636 39924 1642 39936
rect 1673 39933 1685 39936
rect 1719 39933 1731 39967
rect 1673 39927 1731 39933
rect 1854 39924 1860 39976
rect 1912 39924 1918 39976
rect 1946 39924 1952 39976
rect 2004 39924 2010 39976
rect 2038 39924 2044 39976
rect 2096 39924 2102 39976
rect 2314 39924 2320 39976
rect 2372 39924 2378 39976
rect 2746 39964 2774 40004
rect 2866 39992 2872 40044
rect 2924 39992 2930 40044
rect 3344 40032 3372 40072
rect 3252 40004 3372 40032
rect 3252 39964 3280 40004
rect 3418 39992 3424 40044
rect 3476 39992 3482 40044
rect 3528 40032 3556 40072
rect 5721 40069 5733 40103
rect 5767 40069 5779 40103
rect 5721 40063 5779 40069
rect 3528 40004 4568 40032
rect 2746 39936 3280 39964
rect 3326 39924 3332 39976
rect 3384 39964 3390 39976
rect 4065 39967 4123 39973
rect 4065 39964 4077 39967
rect 3384 39936 4077 39964
rect 3384 39924 3390 39936
rect 4065 39933 4077 39936
rect 4111 39933 4123 39967
rect 4540 39964 4568 40004
rect 4614 39992 4620 40044
rect 4672 39992 4678 40044
rect 5736 40032 5764 40063
rect 8018 40060 8024 40112
rect 8076 40100 8082 40112
rect 9784 40100 9812 40131
rect 11238 40100 11244 40112
rect 8076 40072 9812 40100
rect 9876 40072 11244 40100
rect 8076 40060 8082 40072
rect 7101 40035 7159 40041
rect 4724 40004 5856 40032
rect 4724 39964 4752 40004
rect 4540 39936 4752 39964
rect 4801 39967 4859 39973
rect 4065 39927 4123 39933
rect 4801 39933 4813 39967
rect 4847 39933 4859 39967
rect 4801 39927 4859 39933
rect 2682 39896 2688 39908
rect 1228 39868 2688 39896
rect 2682 39856 2688 39868
rect 2740 39896 2746 39908
rect 2958 39896 2964 39908
rect 2740 39868 2964 39896
rect 2740 39856 2746 39868
rect 2958 39856 2964 39868
rect 3016 39856 3022 39908
rect 3050 39856 3056 39908
rect 3108 39896 3114 39908
rect 4816 39896 4844 39927
rect 5166 39924 5172 39976
rect 5224 39924 5230 39976
rect 5442 39924 5448 39976
rect 5500 39924 5506 39976
rect 5629 39967 5687 39973
rect 5629 39933 5641 39967
rect 5675 39964 5687 39967
rect 5828 39964 5856 40004
rect 7101 40001 7113 40035
rect 7147 40032 7159 40035
rect 8570 40032 8576 40044
rect 7147 40004 8576 40032
rect 7147 40001 7159 40004
rect 7101 39995 7159 40001
rect 8570 39992 8576 40004
rect 8628 39992 8634 40044
rect 9876 40032 9904 40072
rect 11238 40060 11244 40072
rect 11296 40060 11302 40112
rect 9324 40004 9904 40032
rect 7745 39967 7803 39973
rect 7745 39964 7757 39967
rect 5675 39936 5764 39964
rect 5828 39936 7757 39964
rect 5675 39933 5687 39936
rect 5629 39927 5687 39933
rect 3108 39868 4844 39896
rect 4985 39899 5043 39905
rect 3108 39856 3114 39868
rect 4985 39865 4997 39899
rect 5031 39865 5043 39899
rect 4985 39859 5043 39865
rect 2225 39831 2283 39837
rect 2225 39797 2237 39831
rect 2271 39828 2283 39831
rect 4522 39828 4528 39840
rect 2271 39800 4528 39828
rect 2271 39797 2283 39800
rect 2225 39791 2283 39797
rect 4522 39788 4528 39800
rect 4580 39788 4586 39840
rect 4706 39788 4712 39840
rect 4764 39828 4770 39840
rect 5000 39828 5028 39859
rect 5074 39856 5080 39908
rect 5132 39856 5138 39908
rect 5184 39896 5212 39924
rect 5736 39896 5764 39936
rect 7745 39933 7757 39936
rect 7791 39933 7803 39967
rect 7745 39927 7803 39933
rect 7834 39924 7840 39976
rect 7892 39964 7898 39976
rect 7929 39967 7987 39973
rect 7929 39964 7941 39967
rect 7892 39936 7941 39964
rect 7892 39924 7898 39936
rect 7929 39933 7941 39936
rect 7975 39933 7987 39967
rect 7929 39927 7987 39933
rect 8386 39924 8392 39976
rect 8444 39924 8450 39976
rect 9125 39967 9183 39973
rect 9125 39933 9137 39967
rect 9171 39964 9183 39967
rect 9324 39964 9352 40004
rect 10042 39992 10048 40044
rect 10100 40032 10106 40044
rect 11054 40032 11060 40044
rect 10100 40004 11060 40032
rect 10100 39992 10106 40004
rect 11054 39992 11060 40004
rect 11112 39992 11118 40044
rect 9171 39936 9352 39964
rect 9401 39967 9459 39973
rect 9171 39933 9183 39936
rect 9125 39927 9183 39933
rect 9401 39933 9413 39967
rect 9447 39966 9459 39967
rect 10229 39967 10287 39973
rect 9447 39964 9536 39966
rect 9447 39938 10180 39964
rect 9447 39933 9459 39938
rect 9508 39936 10180 39938
rect 9401 39927 9459 39933
rect 6454 39896 6460 39908
rect 5184 39868 5672 39896
rect 5736 39868 6460 39896
rect 4764 39800 5028 39828
rect 4764 39788 4770 39800
rect 5350 39788 5356 39840
rect 5408 39788 5414 39840
rect 5534 39788 5540 39840
rect 5592 39788 5598 39840
rect 5644 39828 5672 39868
rect 6454 39856 6460 39868
rect 6512 39856 6518 39908
rect 6638 39856 6644 39908
rect 6696 39896 6702 39908
rect 6834 39899 6892 39905
rect 6834 39896 6846 39899
rect 6696 39868 6846 39896
rect 6696 39856 6702 39868
rect 6834 39865 6846 39868
rect 6880 39865 6892 39899
rect 6834 39859 6892 39865
rect 8662 39856 8668 39908
rect 8720 39856 8726 39908
rect 8754 39856 8760 39908
rect 8812 39856 8818 39908
rect 7006 39828 7012 39840
rect 5644 39800 7012 39828
rect 7006 39788 7012 39800
rect 7064 39788 7070 39840
rect 7098 39788 7104 39840
rect 7156 39828 7162 39840
rect 7193 39831 7251 39837
rect 7193 39828 7205 39831
rect 7156 39800 7205 39828
rect 7156 39788 7162 39800
rect 7193 39797 7205 39800
rect 7239 39797 7251 39831
rect 7193 39791 7251 39797
rect 8110 39788 8116 39840
rect 8168 39788 8174 39840
rect 8478 39788 8484 39840
rect 8536 39788 8542 39840
rect 8570 39788 8576 39840
rect 8628 39828 8634 39840
rect 8849 39831 8907 39837
rect 8849 39828 8861 39831
rect 8628 39800 8861 39828
rect 8628 39788 8634 39800
rect 8849 39797 8861 39800
rect 8895 39797 8907 39831
rect 8849 39791 8907 39797
rect 8938 39788 8944 39840
rect 8996 39828 9002 39840
rect 9692 39828 9720 39936
rect 9769 39899 9827 39905
rect 9769 39865 9781 39899
rect 9815 39896 9827 39899
rect 9858 39896 9864 39908
rect 9815 39868 9864 39896
rect 9815 39865 9827 39868
rect 9769 39859 9827 39865
rect 9858 39856 9864 39868
rect 9916 39856 9922 39908
rect 10152 39896 10180 39936
rect 10229 39933 10241 39967
rect 10275 39964 10287 39967
rect 10594 39964 10600 39976
rect 10275 39936 10600 39964
rect 10275 39933 10287 39936
rect 10229 39927 10287 39933
rect 10594 39924 10600 39936
rect 10652 39924 10658 39976
rect 10410 39896 10416 39908
rect 10152 39868 10416 39896
rect 10410 39856 10416 39868
rect 10468 39856 10474 39908
rect 10686 39856 10692 39908
rect 10744 39896 10750 39908
rect 11146 39896 11152 39908
rect 10744 39868 11152 39896
rect 10744 39856 10750 39868
rect 11146 39856 11152 39868
rect 11204 39856 11210 39908
rect 8996 39800 9720 39828
rect 8996 39788 9002 39800
rect 9950 39788 9956 39840
rect 10008 39788 10014 39840
rect 10226 39788 10232 39840
rect 10284 39828 10290 39840
rect 10597 39831 10655 39837
rect 10597 39828 10609 39831
rect 10284 39800 10609 39828
rect 10284 39788 10290 39800
rect 10597 39797 10609 39800
rect 10643 39797 10655 39831
rect 10597 39791 10655 39797
rect 552 39738 11132 39760
rect 552 39686 4322 39738
rect 4374 39686 4386 39738
rect 4438 39686 4450 39738
rect 4502 39686 4514 39738
rect 4566 39686 4578 39738
rect 4630 39686 10722 39738
rect 10774 39686 10786 39738
rect 10838 39686 10850 39738
rect 10902 39686 10914 39738
rect 10966 39686 10978 39738
rect 11030 39686 11132 39738
rect 552 39664 11132 39686
rect 1578 39584 1584 39636
rect 1636 39584 1642 39636
rect 1670 39584 1676 39636
rect 1728 39584 1734 39636
rect 4154 39584 4160 39636
rect 4212 39584 4218 39636
rect 4706 39584 4712 39636
rect 4764 39624 4770 39636
rect 6546 39624 6552 39636
rect 4764 39596 6552 39624
rect 4764 39584 4770 39596
rect 6546 39584 6552 39596
rect 6604 39584 6610 39636
rect 6638 39584 6644 39636
rect 6696 39584 6702 39636
rect 7098 39584 7104 39636
rect 7156 39584 7162 39636
rect 7374 39584 7380 39636
rect 7432 39624 7438 39636
rect 7745 39627 7803 39633
rect 7745 39624 7757 39627
rect 7432 39596 7757 39624
rect 7432 39584 7438 39596
rect 7745 39593 7757 39596
rect 7791 39624 7803 39627
rect 8938 39624 8944 39636
rect 7791 39596 8944 39624
rect 7791 39593 7803 39596
rect 7745 39587 7803 39593
rect 8938 39584 8944 39596
rect 8996 39624 9002 39636
rect 9582 39624 9588 39636
rect 8996 39596 9588 39624
rect 8996 39584 9002 39596
rect 9582 39584 9588 39596
rect 9640 39584 9646 39636
rect 9766 39624 9772 39636
rect 9692 39596 9772 39624
rect 1596 39556 1624 39584
rect 1946 39556 1952 39568
rect 1596 39528 1952 39556
rect 1946 39516 1952 39528
rect 2004 39516 2010 39568
rect 2038 39516 2044 39568
rect 2096 39556 2102 39568
rect 3142 39556 3148 39568
rect 2096 39528 3148 39556
rect 2096 39516 2102 39528
rect 3142 39516 3148 39528
rect 3200 39556 3206 39568
rect 3602 39556 3608 39568
rect 3200 39528 3608 39556
rect 3200 39516 3206 39528
rect 3602 39516 3608 39528
rect 3660 39516 3666 39568
rect 4065 39559 4123 39565
rect 4065 39525 4077 39559
rect 4111 39556 4123 39559
rect 5442 39556 5448 39568
rect 4111 39528 5448 39556
rect 4111 39525 4123 39528
rect 4065 39519 4123 39525
rect 5442 39516 5448 39528
rect 5500 39556 5506 39568
rect 7009 39559 7067 39565
rect 5500 39528 6040 39556
rect 5500 39516 5506 39528
rect 566 39448 572 39500
rect 624 39488 630 39500
rect 1305 39491 1363 39497
rect 1305 39488 1317 39491
rect 624 39460 1317 39488
rect 624 39448 630 39460
rect 1305 39457 1317 39460
rect 1351 39457 1363 39491
rect 1305 39451 1363 39457
rect 1397 39491 1455 39497
rect 1397 39457 1409 39491
rect 1443 39457 1455 39491
rect 1397 39451 1455 39457
rect 1412 39352 1440 39451
rect 1578 39448 1584 39500
rect 1636 39448 1642 39500
rect 2406 39497 2412 39500
rect 2400 39488 2412 39497
rect 2367 39460 2412 39488
rect 2400 39451 2412 39460
rect 2406 39448 2412 39451
rect 2464 39448 2470 39500
rect 3881 39491 3939 39497
rect 3881 39457 3893 39491
rect 3927 39457 3939 39491
rect 3881 39451 3939 39457
rect 4525 39491 4583 39497
rect 4525 39457 4537 39491
rect 4571 39488 4583 39491
rect 4985 39491 5043 39497
rect 4985 39488 4997 39491
rect 4571 39460 4997 39488
rect 4571 39457 4583 39460
rect 4525 39451 4583 39457
rect 4985 39457 4997 39460
rect 5031 39457 5043 39491
rect 4985 39451 5043 39457
rect 1486 39380 1492 39432
rect 1544 39420 1550 39432
rect 2133 39423 2191 39429
rect 2133 39420 2145 39423
rect 1544 39392 2145 39420
rect 1544 39380 1550 39392
rect 2133 39389 2145 39392
rect 2179 39389 2191 39423
rect 2133 39383 2191 39389
rect 3697 39423 3755 39429
rect 3697 39389 3709 39423
rect 3743 39389 3755 39423
rect 3697 39383 3755 39389
rect 1670 39352 1676 39364
rect 1412 39324 1676 39352
rect 1670 39312 1676 39324
rect 1728 39312 1734 39364
rect 1118 39244 1124 39296
rect 1176 39244 1182 39296
rect 1854 39244 1860 39296
rect 1912 39244 1918 39296
rect 3326 39244 3332 39296
rect 3384 39284 3390 39296
rect 3513 39287 3571 39293
rect 3513 39284 3525 39287
rect 3384 39256 3525 39284
rect 3384 39244 3390 39256
rect 3513 39253 3525 39256
rect 3559 39253 3571 39287
rect 3712 39284 3740 39383
rect 3896 39352 3924 39451
rect 5074 39448 5080 39500
rect 5132 39488 5138 39500
rect 5132 39460 5764 39488
rect 5132 39448 5138 39460
rect 4062 39380 4068 39432
rect 4120 39420 4126 39432
rect 4617 39423 4675 39429
rect 4617 39420 4629 39423
rect 4120 39392 4629 39420
rect 4120 39380 4126 39392
rect 4617 39389 4629 39392
rect 4663 39389 4675 39423
rect 4617 39383 4675 39389
rect 4798 39380 4804 39432
rect 4856 39380 4862 39432
rect 4890 39380 4896 39432
rect 4948 39420 4954 39432
rect 5258 39420 5264 39432
rect 4948 39392 5264 39420
rect 4948 39380 4954 39392
rect 5258 39380 5264 39392
rect 5316 39380 5322 39432
rect 5626 39420 5632 39432
rect 5368 39392 5632 39420
rect 5368 39352 5396 39392
rect 5626 39380 5632 39392
rect 5684 39380 5690 39432
rect 5736 39420 5764 39460
rect 5810 39448 5816 39500
rect 5868 39448 5874 39500
rect 6012 39497 6040 39528
rect 7009 39525 7021 39559
rect 7055 39556 7067 39559
rect 9692 39556 9720 39596
rect 9766 39584 9772 39596
rect 9824 39584 9830 39636
rect 10781 39627 10839 39633
rect 10781 39593 10793 39627
rect 10827 39624 10839 39627
rect 11054 39624 11060 39636
rect 10827 39596 11060 39624
rect 10827 39593 10839 39596
rect 10781 39587 10839 39593
rect 11054 39584 11060 39596
rect 11112 39584 11118 39636
rect 7055 39528 9720 39556
rect 7055 39525 7067 39528
rect 7009 39519 7067 39525
rect 5997 39491 6055 39497
rect 5997 39457 6009 39491
rect 6043 39457 6055 39491
rect 5997 39451 6055 39457
rect 6086 39448 6092 39500
rect 6144 39488 6150 39500
rect 6273 39491 6331 39497
rect 6273 39488 6285 39491
rect 6144 39460 6285 39488
rect 6144 39448 6150 39460
rect 6273 39457 6285 39460
rect 6319 39457 6331 39491
rect 6273 39451 6331 39457
rect 6454 39448 6460 39500
rect 6512 39448 6518 39500
rect 7098 39448 7104 39500
rect 7156 39488 7162 39500
rect 7466 39488 7472 39500
rect 7156 39460 7472 39488
rect 7156 39448 7162 39460
rect 7466 39448 7472 39460
rect 7524 39448 7530 39500
rect 7558 39448 7564 39500
rect 7616 39488 7622 39500
rect 7653 39491 7711 39497
rect 7653 39488 7665 39491
rect 7616 39460 7665 39488
rect 7616 39448 7622 39460
rect 7653 39457 7665 39460
rect 7699 39457 7711 39491
rect 7653 39451 7711 39457
rect 7742 39448 7748 39500
rect 7800 39488 7806 39500
rect 7837 39491 7895 39497
rect 7837 39488 7849 39491
rect 7800 39460 7849 39488
rect 7800 39448 7806 39460
rect 7837 39457 7849 39460
rect 7883 39457 7895 39491
rect 8113 39491 8171 39497
rect 8113 39488 8125 39491
rect 7837 39451 7895 39457
rect 8036 39460 8125 39488
rect 7190 39420 7196 39432
rect 5736 39392 7196 39420
rect 7190 39380 7196 39392
rect 7248 39380 7254 39432
rect 7282 39380 7288 39432
rect 7340 39380 7346 39432
rect 6914 39352 6920 39364
rect 3896 39324 5396 39352
rect 5460 39324 6920 39352
rect 5460 39284 5488 39324
rect 6914 39312 6920 39324
rect 6972 39312 6978 39364
rect 3712 39256 5488 39284
rect 3513 39247 3571 39253
rect 5718 39244 5724 39296
rect 5776 39284 5782 39296
rect 8036 39293 8064 39460
rect 8113 39457 8125 39460
rect 8159 39457 8171 39491
rect 8113 39451 8171 39457
rect 8202 39448 8208 39500
rect 8260 39488 8266 39500
rect 8260 39460 8340 39488
rect 8260 39448 8266 39460
rect 8312 39352 8340 39460
rect 8938 39448 8944 39500
rect 8996 39448 9002 39500
rect 9030 39448 9036 39500
rect 9088 39488 9094 39500
rect 9309 39491 9367 39497
rect 9309 39488 9321 39491
rect 9088 39460 9321 39488
rect 9088 39448 9094 39460
rect 9309 39457 9321 39460
rect 9355 39457 9367 39491
rect 9309 39451 9367 39457
rect 9668 39491 9726 39497
rect 9668 39457 9680 39491
rect 9714 39488 9726 39491
rect 9950 39488 9956 39500
rect 9714 39460 9956 39488
rect 9714 39457 9726 39460
rect 9668 39451 9726 39457
rect 9950 39448 9956 39460
rect 10008 39448 10014 39500
rect 8389 39423 8447 39429
rect 8389 39389 8401 39423
rect 8435 39420 8447 39423
rect 8478 39420 8484 39432
rect 8435 39392 8484 39420
rect 8435 39389 8447 39392
rect 8389 39383 8447 39389
rect 8478 39380 8484 39392
rect 8536 39420 8542 39432
rect 9048 39420 9076 39448
rect 8536 39392 9076 39420
rect 8536 39380 8542 39392
rect 9398 39380 9404 39432
rect 9456 39380 9462 39432
rect 8312 39324 9260 39352
rect 8496 39293 8524 39324
rect 8021 39287 8079 39293
rect 8021 39284 8033 39287
rect 5776 39256 8033 39284
rect 5776 39244 5782 39256
rect 8021 39253 8033 39256
rect 8067 39253 8079 39287
rect 8021 39247 8079 39253
rect 8481 39287 8539 39293
rect 8481 39253 8493 39287
rect 8527 39253 8539 39287
rect 8481 39247 8539 39253
rect 8662 39244 8668 39296
rect 8720 39244 8726 39296
rect 8757 39287 8815 39293
rect 8757 39253 8769 39287
rect 8803 39284 8815 39287
rect 8846 39284 8852 39296
rect 8803 39256 8852 39284
rect 8803 39253 8815 39256
rect 8757 39247 8815 39253
rect 8846 39244 8852 39256
rect 8904 39244 8910 39296
rect 9232 39293 9260 39324
rect 9217 39287 9275 39293
rect 9217 39253 9229 39287
rect 9263 39284 9275 39287
rect 9674 39284 9680 39296
rect 9263 39256 9680 39284
rect 9263 39253 9275 39256
rect 9217 39247 9275 39253
rect 9674 39244 9680 39256
rect 9732 39284 9738 39296
rect 10042 39284 10048 39296
rect 9732 39256 10048 39284
rect 9732 39244 9738 39256
rect 10042 39244 10048 39256
rect 10100 39244 10106 39296
rect 552 39194 11132 39216
rect 552 39142 3662 39194
rect 3714 39142 3726 39194
rect 3778 39142 3790 39194
rect 3842 39142 3854 39194
rect 3906 39142 3918 39194
rect 3970 39142 10062 39194
rect 10114 39142 10126 39194
rect 10178 39142 10190 39194
rect 10242 39142 10254 39194
rect 10306 39142 10318 39194
rect 10370 39142 11132 39194
rect 552 39120 11132 39142
rect 658 39040 664 39092
rect 716 39080 722 39092
rect 937 39083 995 39089
rect 937 39080 949 39083
rect 716 39052 949 39080
rect 716 39040 722 39052
rect 937 39049 949 39052
rect 983 39049 995 39083
rect 937 39043 995 39049
rect 1854 39040 1860 39092
rect 1912 39080 1918 39092
rect 3237 39083 3295 39089
rect 3237 39080 3249 39083
rect 1912 39052 3249 39080
rect 1912 39040 1918 39052
rect 3237 39049 3249 39052
rect 3283 39049 3295 39083
rect 3237 39043 3295 39049
rect 3694 39040 3700 39092
rect 3752 39080 3758 39092
rect 5074 39080 5080 39092
rect 3752 39052 5080 39080
rect 3752 39040 3758 39052
rect 5074 39040 5080 39052
rect 5132 39040 5138 39092
rect 5718 39040 5724 39092
rect 5776 39040 5782 39092
rect 5902 39040 5908 39092
rect 5960 39080 5966 39092
rect 5960 39052 6776 39080
rect 5960 39040 5966 39052
rect 6748 39024 6776 39052
rect 6822 39040 6828 39092
rect 6880 39040 6886 39092
rect 7282 39040 7288 39092
rect 7340 39080 7346 39092
rect 8113 39083 8171 39089
rect 8113 39080 8125 39083
rect 7340 39052 8125 39080
rect 7340 39040 7346 39052
rect 8113 39049 8125 39052
rect 8159 39049 8171 39083
rect 8113 39043 8171 39049
rect 8294 39040 8300 39092
rect 8352 39040 8358 39092
rect 8386 39040 8392 39092
rect 8444 39080 8450 39092
rect 9125 39083 9183 39089
rect 9125 39080 9137 39083
rect 8444 39052 9137 39080
rect 8444 39040 8450 39052
rect 1394 38972 1400 39024
rect 1452 38972 1458 39024
rect 3050 38972 3056 39024
rect 3108 38972 3114 39024
rect 5169 39015 5227 39021
rect 5169 38981 5181 39015
rect 5215 39012 5227 39015
rect 5626 39012 5632 39024
rect 5215 38984 5632 39012
rect 5215 38981 5227 38984
rect 5169 38975 5227 38981
rect 5626 38972 5632 38984
rect 5684 39012 5690 39024
rect 6638 39012 6644 39024
rect 5684 38984 6644 39012
rect 5684 38972 5690 38984
rect 6638 38972 6644 38984
rect 6696 38972 6702 39024
rect 6730 38972 6736 39024
rect 6788 39012 6794 39024
rect 8202 39012 8208 39024
rect 6788 38984 8208 39012
rect 6788 38972 6794 38984
rect 1302 38944 1308 38956
rect 860 38916 1308 38944
rect 860 38885 888 38916
rect 1302 38904 1308 38916
rect 1360 38904 1366 38956
rect 1486 38904 1492 38956
rect 1544 38944 1550 38956
rect 7116 38953 7144 38984
rect 8202 38972 8208 38984
rect 8260 38972 8266 39024
rect 1673 38947 1731 38953
rect 1673 38944 1685 38947
rect 1544 38916 1685 38944
rect 1544 38904 1550 38916
rect 1673 38913 1685 38916
rect 1719 38913 1731 38947
rect 5353 38947 5411 38953
rect 1673 38907 1731 38913
rect 2746 38916 3832 38944
rect 845 38879 903 38885
rect 845 38845 857 38879
rect 891 38845 903 38879
rect 845 38839 903 38845
rect 1026 38836 1032 38888
rect 1084 38836 1090 38888
rect 1688 38876 1716 38907
rect 2746 38876 2774 38916
rect 3804 38885 3832 38916
rect 5353 38913 5365 38947
rect 5399 38944 5411 38947
rect 7009 38947 7067 38953
rect 7009 38944 7021 38947
rect 5399 38916 7021 38944
rect 5399 38913 5411 38916
rect 5353 38907 5411 38913
rect 7009 38913 7021 38916
rect 7055 38913 7067 38947
rect 7009 38907 7067 38913
rect 7101 38947 7159 38953
rect 7101 38913 7113 38947
rect 7147 38913 7159 38947
rect 7101 38907 7159 38913
rect 7190 38904 7196 38956
rect 7248 38944 7254 38956
rect 7837 38947 7895 38953
rect 7248 38916 7788 38944
rect 7248 38904 7254 38916
rect 7760 38888 7788 38916
rect 7837 38913 7849 38947
rect 7883 38944 7895 38947
rect 8312 38944 8340 39040
rect 7883 38916 8340 38944
rect 7883 38913 7895 38916
rect 7837 38907 7895 38913
rect 8386 38904 8392 38956
rect 8444 38944 8450 38956
rect 8444 38916 8616 38944
rect 8444 38904 8450 38916
rect 1688 38848 2774 38876
rect 3421 38879 3479 38885
rect 3421 38845 3433 38879
rect 3467 38845 3479 38879
rect 3421 38839 3479 38845
rect 3513 38879 3571 38885
rect 3513 38845 3525 38879
rect 3559 38845 3571 38879
rect 3513 38839 3571 38845
rect 3789 38879 3847 38885
rect 3789 38845 3801 38879
rect 3835 38876 3847 38879
rect 3878 38876 3884 38888
rect 3835 38848 3884 38876
rect 3835 38845 3847 38848
rect 3789 38839 3847 38845
rect 1118 38768 1124 38820
rect 1176 38768 1182 38820
rect 1918 38811 1976 38817
rect 1918 38808 1930 38811
rect 1596 38780 1930 38808
rect 1596 38749 1624 38780
rect 1918 38777 1930 38780
rect 1964 38808 1976 38811
rect 3436 38808 3464 38839
rect 1964 38780 3464 38808
rect 1964 38777 1976 38780
rect 1918 38771 1976 38777
rect 1581 38743 1639 38749
rect 1581 38709 1593 38743
rect 1627 38709 1639 38743
rect 1581 38703 1639 38709
rect 1670 38700 1676 38752
rect 1728 38740 1734 38752
rect 3528 38740 3556 38839
rect 3878 38836 3884 38848
rect 3936 38836 3942 38888
rect 5537 38879 5595 38885
rect 5537 38845 5549 38879
rect 5583 38845 5595 38879
rect 5537 38839 5595 38845
rect 5813 38879 5871 38885
rect 5813 38845 5825 38879
rect 5859 38876 5871 38879
rect 5902 38876 5908 38888
rect 5859 38848 5908 38876
rect 5859 38845 5871 38848
rect 5813 38839 5871 38845
rect 4056 38811 4114 38817
rect 4056 38777 4068 38811
rect 4102 38808 4114 38811
rect 4154 38808 4160 38820
rect 4102 38780 4160 38808
rect 4102 38777 4114 38780
rect 4056 38771 4114 38777
rect 4154 38768 4160 38780
rect 4212 38768 4218 38820
rect 5552 38808 5580 38839
rect 5902 38836 5908 38848
rect 5960 38836 5966 38888
rect 6549 38879 6607 38885
rect 6549 38845 6561 38879
rect 6595 38876 6607 38879
rect 6730 38876 6736 38888
rect 6595 38848 6736 38876
rect 6595 38845 6607 38848
rect 6549 38839 6607 38845
rect 6730 38836 6736 38848
rect 6788 38836 6794 38888
rect 7282 38836 7288 38888
rect 7340 38876 7346 38888
rect 7377 38879 7435 38885
rect 7377 38876 7389 38879
rect 7340 38848 7389 38876
rect 7340 38836 7346 38848
rect 7377 38845 7389 38848
rect 7423 38845 7435 38879
rect 7377 38839 7435 38845
rect 6822 38808 6828 38820
rect 5552 38780 6828 38808
rect 6822 38768 6828 38780
rect 6880 38768 6886 38820
rect 7392 38808 7420 38839
rect 7466 38836 7472 38888
rect 7524 38836 7530 38888
rect 7558 38836 7564 38888
rect 7616 38876 7622 38888
rect 7653 38879 7711 38885
rect 7653 38876 7665 38879
rect 7616 38848 7665 38876
rect 7616 38836 7622 38848
rect 7653 38845 7665 38848
rect 7699 38845 7711 38879
rect 7653 38839 7711 38845
rect 7742 38836 7748 38888
rect 7800 38836 7806 38888
rect 7926 38836 7932 38888
rect 7984 38836 7990 38888
rect 8202 38836 8208 38888
rect 8260 38878 8266 38888
rect 8294 38878 8300 38888
rect 8260 38848 8300 38878
rect 8260 38836 8266 38848
rect 8294 38836 8300 38848
rect 8352 38836 8358 38888
rect 8588 38885 8616 38916
rect 8671 38885 8699 39052
rect 9125 39049 9137 39052
rect 9171 39080 9183 39083
rect 9582 39080 9588 39092
rect 9171 39052 9588 39080
rect 9171 39049 9183 39052
rect 9125 39043 9183 39049
rect 9582 39040 9588 39052
rect 9640 39040 9646 39092
rect 9766 39040 9772 39092
rect 9824 39040 9830 39092
rect 8938 38972 8944 39024
rect 8996 38972 9002 39024
rect 9677 39015 9735 39021
rect 9677 38981 9689 39015
rect 9723 39012 9735 39015
rect 9950 39012 9956 39024
rect 9723 38984 9956 39012
rect 9723 38981 9735 38984
rect 9677 38975 9735 38981
rect 9950 38972 9956 38984
rect 10008 38972 10014 39024
rect 8956 38944 8984 38972
rect 8956 38916 9536 38944
rect 8573 38879 8631 38885
rect 8573 38845 8585 38879
rect 8619 38845 8631 38879
rect 8573 38839 8631 38845
rect 8665 38879 8723 38885
rect 8665 38845 8677 38879
rect 8711 38845 8723 38879
rect 8665 38839 8723 38845
rect 8846 38836 8852 38888
rect 8904 38836 8910 38888
rect 8938 38836 8944 38888
rect 8996 38836 9002 38888
rect 9508 38885 9536 38916
rect 9582 38904 9588 38956
rect 9640 38944 9646 38956
rect 9640 38916 10456 38944
rect 9640 38904 9646 38916
rect 9401 38879 9459 38885
rect 9401 38845 9413 38879
rect 9447 38845 9459 38879
rect 9401 38839 9459 38845
rect 9493 38879 9551 38885
rect 9493 38845 9505 38879
rect 9539 38845 9551 38879
rect 9493 38839 9551 38845
rect 9033 38811 9091 38817
rect 9033 38808 9045 38811
rect 7392 38780 9045 38808
rect 9033 38777 9045 38780
rect 9079 38777 9091 38811
rect 9416 38808 9444 38839
rect 9858 38836 9864 38888
rect 9916 38876 9922 38888
rect 9953 38879 10011 38885
rect 9953 38876 9965 38879
rect 9916 38848 9965 38876
rect 9916 38836 9922 38848
rect 9953 38845 9965 38848
rect 9999 38845 10011 38879
rect 9953 38839 10011 38845
rect 10134 38836 10140 38888
rect 10192 38836 10198 38888
rect 10428 38885 10456 38916
rect 10413 38879 10471 38885
rect 10413 38845 10425 38879
rect 10459 38845 10471 38879
rect 10413 38839 10471 38845
rect 9674 38808 9680 38820
rect 9416 38780 9680 38808
rect 9033 38771 9091 38777
rect 9674 38768 9680 38780
rect 9732 38768 9738 38820
rect 10597 38811 10655 38817
rect 10597 38808 10609 38811
rect 10428 38780 10609 38808
rect 10428 38752 10456 38780
rect 10597 38777 10609 38780
rect 10643 38777 10655 38811
rect 10597 38771 10655 38777
rect 1728 38712 3556 38740
rect 1728 38700 1734 38712
rect 5902 38700 5908 38752
rect 5960 38700 5966 38752
rect 7098 38700 7104 38752
rect 7156 38740 7162 38752
rect 7193 38743 7251 38749
rect 7193 38740 7205 38743
rect 7156 38712 7205 38740
rect 7156 38700 7162 38712
rect 7193 38709 7205 38712
rect 7239 38740 7251 38743
rect 8294 38740 8300 38752
rect 7239 38712 8300 38740
rect 7239 38709 7251 38712
rect 7193 38703 7251 38709
rect 8294 38700 8300 38712
rect 8352 38700 8358 38752
rect 8389 38743 8447 38749
rect 8389 38709 8401 38743
rect 8435 38740 8447 38743
rect 8478 38740 8484 38752
rect 8435 38712 8484 38740
rect 8435 38709 8447 38712
rect 8389 38703 8447 38709
rect 8478 38700 8484 38712
rect 8536 38700 8542 38752
rect 8662 38700 8668 38752
rect 8720 38740 8726 38752
rect 9306 38740 9312 38752
rect 8720 38712 9312 38740
rect 8720 38700 8726 38712
rect 9306 38700 9312 38712
rect 9364 38700 9370 38752
rect 10226 38700 10232 38752
rect 10284 38700 10290 38752
rect 10410 38700 10416 38752
rect 10468 38700 10474 38752
rect 552 38650 11132 38672
rect 552 38598 4322 38650
rect 4374 38598 4386 38650
rect 4438 38598 4450 38650
rect 4502 38598 4514 38650
rect 4566 38598 4578 38650
rect 4630 38598 10722 38650
rect 10774 38598 10786 38650
rect 10838 38598 10850 38650
rect 10902 38598 10914 38650
rect 10966 38598 10978 38650
rect 11030 38598 11132 38650
rect 552 38576 11132 38598
rect 750 38496 756 38548
rect 808 38536 814 38548
rect 1305 38539 1363 38545
rect 1305 38536 1317 38539
rect 808 38508 1317 38536
rect 808 38496 814 38508
rect 1305 38505 1317 38508
rect 1351 38505 1363 38539
rect 1305 38499 1363 38505
rect 1762 38496 1768 38548
rect 1820 38496 1826 38548
rect 2406 38536 2412 38548
rect 1872 38508 2412 38536
rect 937 38471 995 38477
rect 937 38437 949 38471
rect 983 38437 995 38471
rect 937 38431 995 38437
rect 1167 38437 1225 38443
rect 952 38332 980 38431
rect 1167 38403 1179 38437
rect 1213 38434 1225 38437
rect 1213 38403 1236 38434
rect 1167 38400 1236 38403
rect 1302 38400 1308 38412
rect 1167 38397 1308 38400
rect 1208 38372 1308 38397
rect 1302 38360 1308 38372
rect 1360 38400 1366 38412
rect 1581 38403 1639 38409
rect 1581 38400 1593 38403
rect 1360 38372 1593 38400
rect 1360 38360 1366 38372
rect 1581 38369 1593 38372
rect 1627 38400 1639 38403
rect 1872 38400 1900 38508
rect 2406 38496 2412 38508
rect 2464 38496 2470 38548
rect 3786 38496 3792 38548
rect 3844 38536 3850 38548
rect 3973 38539 4031 38545
rect 3973 38536 3985 38539
rect 3844 38508 3985 38536
rect 3844 38496 3850 38508
rect 3973 38505 3985 38508
rect 4019 38505 4031 38539
rect 3973 38499 4031 38505
rect 5350 38496 5356 38548
rect 5408 38536 5414 38548
rect 5408 38508 5856 38536
rect 5408 38496 5414 38508
rect 2124 38471 2182 38477
rect 2124 38437 2136 38471
rect 2170 38468 2182 38471
rect 2314 38468 2320 38480
rect 2170 38440 2320 38468
rect 2170 38437 2182 38440
rect 2124 38431 2182 38437
rect 2314 38428 2320 38440
rect 2372 38428 2378 38480
rect 3234 38428 3240 38480
rect 3292 38468 3298 38480
rect 3694 38468 3700 38480
rect 3292 38440 3700 38468
rect 3292 38428 3298 38440
rect 3694 38428 3700 38440
rect 3752 38428 3758 38480
rect 4062 38428 4068 38480
rect 4120 38468 4126 38480
rect 5828 38468 5856 38508
rect 5902 38496 5908 38548
rect 5960 38536 5966 38548
rect 6181 38539 6239 38545
rect 6181 38536 6193 38539
rect 5960 38508 6193 38536
rect 5960 38496 5966 38508
rect 6181 38505 6193 38508
rect 6227 38505 6239 38539
rect 6181 38499 6239 38505
rect 7285 38539 7343 38545
rect 7285 38505 7297 38539
rect 7331 38536 7343 38539
rect 7466 38536 7472 38548
rect 7331 38508 7472 38536
rect 7331 38505 7343 38508
rect 7285 38499 7343 38505
rect 7466 38496 7472 38508
rect 7524 38496 7530 38548
rect 7742 38496 7748 38548
rect 7800 38536 7806 38548
rect 8205 38539 8263 38545
rect 8205 38536 8217 38539
rect 7800 38508 8217 38536
rect 7800 38496 7806 38508
rect 8205 38505 8217 38508
rect 8251 38536 8263 38539
rect 8251 38508 8800 38536
rect 8251 38505 8263 38508
rect 8205 38499 8263 38505
rect 6273 38471 6331 38477
rect 6273 38468 6285 38471
rect 4120 38440 5488 38468
rect 5828 38440 6285 38468
rect 4120 38428 4126 38440
rect 1627 38372 1900 38400
rect 1627 38369 1639 38372
rect 1581 38363 1639 38369
rect 1946 38360 1952 38412
rect 2004 38400 2010 38412
rect 3421 38403 3479 38409
rect 3421 38400 3433 38403
rect 2004 38372 3433 38400
rect 2004 38360 2010 38372
rect 3421 38369 3433 38372
rect 3467 38369 3479 38403
rect 3421 38363 3479 38369
rect 1397 38335 1455 38341
rect 1397 38332 1409 38335
rect 952 38304 1409 38332
rect 1397 38301 1409 38304
rect 1443 38301 1455 38335
rect 1397 38295 1455 38301
rect 382 38224 388 38276
rect 440 38264 446 38276
rect 1412 38264 1440 38295
rect 1486 38292 1492 38344
rect 1544 38332 1550 38344
rect 1857 38335 1915 38341
rect 1857 38332 1869 38335
rect 1544 38304 1869 38332
rect 1544 38292 1550 38304
rect 1857 38301 1869 38304
rect 1903 38301 1915 38335
rect 3436 38332 3464 38363
rect 3510 38360 3516 38412
rect 3568 38400 3574 38412
rect 3605 38403 3663 38409
rect 3605 38400 3617 38403
rect 3568 38372 3617 38400
rect 3568 38360 3574 38372
rect 3605 38369 3617 38372
rect 3651 38369 3663 38403
rect 3605 38363 3663 38369
rect 3786 38360 3792 38412
rect 3844 38360 3850 38412
rect 4706 38400 4712 38412
rect 4448 38372 4712 38400
rect 4448 38332 4476 38372
rect 4706 38360 4712 38372
rect 4764 38360 4770 38412
rect 5460 38409 5488 38440
rect 6273 38437 6285 38440
rect 6319 38437 6331 38471
rect 7374 38468 7380 38480
rect 6273 38431 6331 38437
rect 6748 38440 7380 38468
rect 5189 38403 5247 38409
rect 5189 38369 5201 38403
rect 5235 38400 5247 38403
rect 5445 38403 5503 38409
rect 5235 38372 5396 38400
rect 5235 38369 5247 38372
rect 5189 38363 5247 38369
rect 3436 38304 4476 38332
rect 5368 38332 5396 38372
rect 5445 38369 5457 38403
rect 5491 38369 5503 38403
rect 5445 38363 5503 38369
rect 5626 38360 5632 38412
rect 5684 38400 5690 38412
rect 6748 38400 6776 38440
rect 5684 38372 6776 38400
rect 6825 38403 6883 38409
rect 5684 38360 5690 38372
rect 6825 38369 6837 38403
rect 6871 38400 6883 38403
rect 7006 38400 7012 38412
rect 6871 38372 7012 38400
rect 6871 38369 6883 38372
rect 6825 38363 6883 38369
rect 7006 38360 7012 38372
rect 7064 38360 7070 38412
rect 7116 38409 7144 38440
rect 7374 38428 7380 38440
rect 7432 38428 7438 38480
rect 7653 38471 7711 38477
rect 7653 38437 7665 38471
rect 7699 38468 7711 38471
rect 8294 38468 8300 38480
rect 7699 38440 8300 38468
rect 7699 38437 7711 38440
rect 7653 38431 7711 38437
rect 8294 38428 8300 38440
rect 8352 38428 8358 38480
rect 8772 38468 8800 38508
rect 8938 38496 8944 38548
rect 8996 38536 9002 38548
rect 9125 38539 9183 38545
rect 9125 38536 9137 38539
rect 8996 38508 9137 38536
rect 8996 38496 9002 38508
rect 9125 38505 9137 38508
rect 9171 38505 9183 38539
rect 9125 38499 9183 38505
rect 9214 38496 9220 38548
rect 9272 38496 9278 38548
rect 9858 38496 9864 38548
rect 9916 38536 9922 38548
rect 10413 38539 10471 38545
rect 10413 38536 10425 38539
rect 9916 38508 10425 38536
rect 9916 38496 9922 38508
rect 10413 38505 10425 38508
rect 10459 38505 10471 38539
rect 10413 38499 10471 38505
rect 9232 38468 9260 38496
rect 8772 38440 9260 38468
rect 7101 38403 7159 38409
rect 7101 38369 7113 38403
rect 7147 38369 7159 38403
rect 7101 38363 7159 38369
rect 7282 38360 7288 38412
rect 7340 38400 7346 38412
rect 7561 38403 7619 38409
rect 7561 38400 7573 38403
rect 7340 38372 7573 38400
rect 7340 38360 7346 38372
rect 7561 38369 7573 38372
rect 7607 38400 7619 38403
rect 7607 38372 7696 38400
rect 7607 38369 7619 38372
rect 7561 38363 7619 38369
rect 5368 38304 5856 38332
rect 1857 38295 1915 38301
rect 1670 38264 1676 38276
rect 440 38236 1348 38264
rect 1412 38236 1676 38264
rect 440 38224 446 38236
rect 1118 38156 1124 38208
rect 1176 38156 1182 38208
rect 1320 38196 1348 38236
rect 1670 38224 1676 38236
rect 1728 38224 1734 38276
rect 2958 38224 2964 38276
rect 3016 38264 3022 38276
rect 4430 38264 4436 38276
rect 3016 38236 4436 38264
rect 3016 38224 3022 38236
rect 4430 38224 4436 38236
rect 4488 38224 4494 38276
rect 5828 38273 5856 38304
rect 6270 38292 6276 38344
rect 6328 38332 6334 38344
rect 6365 38335 6423 38341
rect 6365 38332 6377 38335
rect 6328 38304 6377 38332
rect 6328 38292 6334 38304
rect 6365 38301 6377 38304
rect 6411 38301 6423 38335
rect 6365 38295 6423 38301
rect 6914 38292 6920 38344
rect 6972 38292 6978 38344
rect 5813 38267 5871 38273
rect 5813 38233 5825 38267
rect 5859 38233 5871 38267
rect 5813 38227 5871 38233
rect 7098 38224 7104 38276
rect 7156 38264 7162 38276
rect 7377 38267 7435 38273
rect 7377 38264 7389 38267
rect 7156 38236 7389 38264
rect 7156 38224 7162 38236
rect 7377 38233 7389 38236
rect 7423 38233 7435 38267
rect 7668 38264 7696 38372
rect 7742 38360 7748 38412
rect 7800 38360 7806 38412
rect 8018 38360 8024 38412
rect 8076 38360 8082 38412
rect 8386 38360 8392 38412
rect 8444 38360 8450 38412
rect 8849 38403 8907 38409
rect 8849 38369 8861 38403
rect 8895 38400 8907 38403
rect 8938 38400 8944 38412
rect 8895 38372 8944 38400
rect 8895 38369 8907 38372
rect 8849 38363 8907 38369
rect 8938 38360 8944 38372
rect 8996 38360 9002 38412
rect 9232 38400 9260 38440
rect 9674 38428 9680 38480
rect 9732 38468 9738 38480
rect 9732 38440 10272 38468
rect 9732 38428 9738 38440
rect 10244 38409 10272 38440
rect 9493 38403 9551 38409
rect 9493 38400 9505 38403
rect 9232 38372 9505 38400
rect 9493 38369 9505 38372
rect 9539 38369 9551 38403
rect 9493 38363 9551 38369
rect 9953 38403 10011 38409
rect 9953 38369 9965 38403
rect 9999 38369 10011 38403
rect 9953 38363 10011 38369
rect 10229 38403 10287 38409
rect 10229 38369 10241 38403
rect 10275 38369 10287 38403
rect 10229 38363 10287 38369
rect 7760 38332 7788 38360
rect 8665 38335 8723 38341
rect 8665 38332 8677 38335
rect 7760 38304 8677 38332
rect 8665 38301 8677 38304
rect 8711 38301 8723 38335
rect 8665 38295 8723 38301
rect 8757 38335 8815 38341
rect 8757 38301 8769 38335
rect 8803 38332 8815 38335
rect 9217 38335 9275 38341
rect 9217 38332 9229 38335
rect 8803 38304 9229 38332
rect 8803 38301 8815 38304
rect 8757 38295 8815 38301
rect 9217 38301 9229 38304
rect 9263 38332 9275 38335
rect 9306 38332 9312 38344
rect 9263 38304 9312 38332
rect 9263 38301 9275 38304
rect 9217 38295 9275 38301
rect 9306 38292 9312 38304
rect 9364 38292 9370 38344
rect 8573 38267 8631 38273
rect 8573 38264 8585 38267
rect 7668 38236 8585 38264
rect 7377 38227 7435 38233
rect 8573 38233 8585 38236
rect 8619 38233 8631 38267
rect 8573 38227 8631 38233
rect 9122 38224 9128 38276
rect 9180 38264 9186 38276
rect 9968 38264 9996 38363
rect 10502 38360 10508 38412
rect 10560 38360 10566 38412
rect 10042 38292 10048 38344
rect 10100 38332 10106 38344
rect 10137 38335 10195 38341
rect 10137 38332 10149 38335
rect 10100 38304 10149 38332
rect 10100 38292 10106 38304
rect 10137 38301 10149 38304
rect 10183 38301 10195 38335
rect 10137 38295 10195 38301
rect 9180 38236 9996 38264
rect 10152 38264 10180 38295
rect 10502 38264 10508 38276
rect 10152 38236 10508 38264
rect 9180 38224 9186 38236
rect 10502 38224 10508 38236
rect 10560 38224 10566 38276
rect 2498 38196 2504 38208
rect 1320 38168 2504 38196
rect 2498 38156 2504 38168
rect 2556 38156 2562 38208
rect 3237 38199 3295 38205
rect 3237 38165 3249 38199
rect 3283 38196 3295 38199
rect 3510 38196 3516 38208
rect 3283 38168 3516 38196
rect 3283 38165 3295 38168
rect 3237 38159 3295 38165
rect 3510 38156 3516 38168
rect 3568 38156 3574 38208
rect 4065 38199 4123 38205
rect 4065 38165 4077 38199
rect 4111 38196 4123 38199
rect 4154 38196 4160 38208
rect 4111 38168 4160 38196
rect 4111 38165 4123 38168
rect 4065 38159 4123 38165
rect 4154 38156 4160 38168
rect 4212 38196 4218 38208
rect 6730 38196 6736 38208
rect 4212 38168 6736 38196
rect 4212 38156 4218 38168
rect 6730 38156 6736 38168
rect 6788 38156 6794 38208
rect 7009 38199 7067 38205
rect 7009 38165 7021 38199
rect 7055 38196 7067 38199
rect 7282 38196 7288 38208
rect 7055 38168 7288 38196
rect 7055 38165 7067 38168
rect 7009 38159 7067 38165
rect 7282 38156 7288 38168
rect 7340 38196 7346 38208
rect 7466 38196 7472 38208
rect 7340 38168 7472 38196
rect 7340 38156 7346 38168
rect 7466 38156 7472 38168
rect 7524 38156 7530 38208
rect 7650 38156 7656 38208
rect 7708 38196 7714 38208
rect 7929 38199 7987 38205
rect 7929 38196 7941 38199
rect 7708 38168 7941 38196
rect 7708 38156 7714 38168
rect 7929 38165 7941 38168
rect 7975 38165 7987 38199
rect 7929 38159 7987 38165
rect 8110 38156 8116 38208
rect 8168 38196 8174 38208
rect 9214 38196 9220 38208
rect 8168 38168 9220 38196
rect 8168 38156 8174 38168
rect 9214 38156 9220 38168
rect 9272 38196 9278 38208
rect 9309 38199 9367 38205
rect 9309 38196 9321 38199
rect 9272 38168 9321 38196
rect 9272 38156 9278 38168
rect 9309 38165 9321 38168
rect 9355 38165 9367 38199
rect 9309 38159 9367 38165
rect 9677 38199 9735 38205
rect 9677 38165 9689 38199
rect 9723 38196 9735 38199
rect 9766 38196 9772 38208
rect 9723 38168 9772 38196
rect 9723 38165 9735 38168
rect 9677 38159 9735 38165
rect 9766 38156 9772 38168
rect 9824 38156 9830 38208
rect 9950 38156 9956 38208
rect 10008 38196 10014 38208
rect 10226 38196 10232 38208
rect 10008 38168 10232 38196
rect 10008 38156 10014 38168
rect 10226 38156 10232 38168
rect 10284 38156 10290 38208
rect 10318 38156 10324 38208
rect 10376 38196 10382 38208
rect 10689 38199 10747 38205
rect 10689 38196 10701 38199
rect 10376 38168 10701 38196
rect 10376 38156 10382 38168
rect 10689 38165 10701 38168
rect 10735 38196 10747 38199
rect 11054 38196 11060 38208
rect 10735 38168 11060 38196
rect 10735 38165 10747 38168
rect 10689 38159 10747 38165
rect 11054 38156 11060 38168
rect 11112 38156 11118 38208
rect 552 38106 11132 38128
rect 552 38054 3662 38106
rect 3714 38054 3726 38106
rect 3778 38054 3790 38106
rect 3842 38054 3854 38106
rect 3906 38054 3918 38106
rect 3970 38054 10062 38106
rect 10114 38054 10126 38106
rect 10178 38054 10190 38106
rect 10242 38054 10254 38106
rect 10306 38054 10318 38106
rect 10370 38054 11132 38106
rect 552 38032 11132 38054
rect 842 37952 848 38004
rect 900 37992 906 38004
rect 937 37995 995 38001
rect 937 37992 949 37995
rect 900 37964 949 37992
rect 900 37952 906 37964
rect 937 37961 949 37964
rect 983 37961 995 37995
rect 937 37955 995 37961
rect 2130 37952 2136 38004
rect 2188 37952 2194 38004
rect 2498 37952 2504 38004
rect 2556 37952 2562 38004
rect 2958 37952 2964 38004
rect 3016 37952 3022 38004
rect 3050 37952 3056 38004
rect 3108 37992 3114 38004
rect 3326 37992 3332 38004
rect 3108 37964 3332 37992
rect 3108 37952 3114 37964
rect 3326 37952 3332 37964
rect 3384 37952 3390 38004
rect 3878 37952 3884 38004
rect 3936 37992 3942 38004
rect 5626 37992 5632 38004
rect 3936 37964 5632 37992
rect 3936 37952 3942 37964
rect 5626 37952 5632 37964
rect 5684 37952 5690 38004
rect 7193 37995 7251 38001
rect 7193 37961 7205 37995
rect 7239 37961 7251 37995
rect 7193 37955 7251 37961
rect 7377 37995 7435 38001
rect 7377 37961 7389 37995
rect 7423 37992 7435 37995
rect 7558 37992 7564 38004
rect 7423 37964 7564 37992
rect 7423 37961 7435 37964
rect 7377 37955 7435 37961
rect 1118 37884 1124 37936
rect 1176 37884 1182 37936
rect 2406 37884 2412 37936
rect 2464 37924 2470 37936
rect 3237 37927 3295 37933
rect 3237 37924 3249 37927
rect 2464 37896 3249 37924
rect 2464 37884 2470 37896
rect 3237 37893 3249 37896
rect 3283 37893 3295 37927
rect 3237 37887 3295 37893
rect 3970 37884 3976 37936
rect 4028 37924 4034 37936
rect 7208 37924 7236 37955
rect 7558 37952 7564 37964
rect 7616 37952 7622 38004
rect 7837 37995 7895 38001
rect 7837 37961 7849 37995
rect 7883 37961 7895 37995
rect 7837 37955 7895 37961
rect 7742 37924 7748 37936
rect 4028 37896 6960 37924
rect 7208 37896 7748 37924
rect 4028 37884 4034 37896
rect 1136 37856 1164 37884
rect 1857 37859 1915 37865
rect 1857 37856 1869 37859
rect 1136 37828 1869 37856
rect 1857 37825 1869 37828
rect 1903 37825 1915 37859
rect 1857 37819 1915 37825
rect 3326 37816 3332 37868
rect 3384 37856 3390 37868
rect 3789 37859 3847 37865
rect 3789 37856 3801 37859
rect 3384 37828 3801 37856
rect 3384 37816 3390 37828
rect 3789 37825 3801 37828
rect 3835 37825 3847 37859
rect 3789 37819 3847 37825
rect 4798 37816 4804 37868
rect 4856 37856 4862 37868
rect 6270 37856 6276 37868
rect 4856 37828 6276 37856
rect 4856 37816 4862 37828
rect 6270 37816 6276 37828
rect 6328 37816 6334 37868
rect 6932 37865 6960 37896
rect 7742 37884 7748 37896
rect 7800 37884 7806 37936
rect 7852 37924 7880 37955
rect 7926 37952 7932 38004
rect 7984 37992 7990 38004
rect 8389 37995 8447 38001
rect 8389 37992 8401 37995
rect 7984 37964 8401 37992
rect 7984 37952 7990 37964
rect 8389 37961 8401 37964
rect 8435 37961 8447 37995
rect 8389 37955 8447 37961
rect 8849 37995 8907 38001
rect 8849 37961 8861 37995
rect 8895 37992 8907 37995
rect 9122 37992 9128 38004
rect 8895 37964 9128 37992
rect 8895 37961 8907 37964
rect 8849 37955 8907 37961
rect 9122 37952 9128 37964
rect 9180 37952 9186 38004
rect 9582 37952 9588 38004
rect 9640 37952 9646 38004
rect 8110 37924 8116 37936
rect 7852 37896 8116 37924
rect 8110 37884 8116 37896
rect 8168 37884 8174 37936
rect 10502 37924 10508 37936
rect 8496 37896 8800 37924
rect 6917 37859 6975 37865
rect 6917 37825 6929 37859
rect 6963 37856 6975 37859
rect 7098 37856 7104 37868
rect 6963 37828 7104 37856
rect 6963 37825 6975 37828
rect 6917 37819 6975 37825
rect 7098 37816 7104 37828
rect 7156 37816 7162 37868
rect 7929 37859 7987 37865
rect 7929 37825 7941 37859
rect 7975 37856 7987 37859
rect 8496 37856 8524 37896
rect 7975 37828 8524 37856
rect 7975 37825 7987 37828
rect 7929 37819 7987 37825
rect 8570 37816 8576 37868
rect 8628 37856 8634 37868
rect 8772 37856 8800 37896
rect 9508 37896 10508 37924
rect 8941 37859 8999 37865
rect 8628 37828 8708 37856
rect 8772 37828 8892 37856
rect 8628 37816 8634 37828
rect 106 37748 112 37800
rect 164 37788 170 37800
rect 1121 37791 1179 37797
rect 1121 37788 1133 37791
rect 164 37760 1133 37788
rect 164 37748 170 37760
rect 1121 37757 1133 37760
rect 1167 37757 1179 37791
rect 1121 37751 1179 37757
rect 1578 37748 1584 37800
rect 1636 37748 1642 37800
rect 1765 37791 1823 37797
rect 1765 37757 1777 37791
rect 1811 37757 1823 37791
rect 1765 37751 1823 37757
rect 1596 37720 1624 37748
rect 1136 37692 1624 37720
rect 1780 37720 1808 37751
rect 1946 37748 1952 37800
rect 2004 37748 2010 37800
rect 2314 37748 2320 37800
rect 2372 37748 2378 37800
rect 2777 37791 2835 37797
rect 2777 37788 2789 37791
rect 2424 37760 2789 37788
rect 1854 37720 1860 37732
rect 1780 37692 1860 37720
rect 1136 37664 1164 37692
rect 1854 37680 1860 37692
rect 1912 37680 1918 37732
rect 2130 37680 2136 37732
rect 2188 37720 2194 37732
rect 2424 37720 2452 37760
rect 2777 37757 2789 37760
rect 2823 37757 2835 37791
rect 2777 37751 2835 37757
rect 3602 37748 3608 37800
rect 3660 37748 3666 37800
rect 4246 37748 4252 37800
rect 4304 37748 4310 37800
rect 4706 37748 4712 37800
rect 4764 37788 4770 37800
rect 5442 37788 5448 37800
rect 4764 37760 5448 37788
rect 4764 37748 4770 37760
rect 5442 37748 5448 37760
rect 5500 37748 5506 37800
rect 5534 37748 5540 37800
rect 5592 37748 5598 37800
rect 5997 37791 6055 37797
rect 5997 37757 6009 37791
rect 6043 37788 6055 37791
rect 6086 37788 6092 37800
rect 6043 37760 6092 37788
rect 6043 37757 6055 37760
rect 5997 37751 6055 37757
rect 6086 37748 6092 37760
rect 6144 37748 6150 37800
rect 6730 37748 6736 37800
rect 6788 37748 6794 37800
rect 6822 37748 6828 37800
rect 6880 37788 6886 37800
rect 7745 37791 7803 37797
rect 6880 37760 7052 37788
rect 6880 37748 6886 37760
rect 2188 37692 2452 37720
rect 2188 37680 2194 37692
rect 2498 37680 2504 37732
rect 2556 37720 2562 37732
rect 4264 37720 4292 37748
rect 2556 37692 4292 37720
rect 4617 37723 4675 37729
rect 2556 37680 2562 37692
rect 4617 37689 4629 37723
rect 4663 37720 4675 37723
rect 6178 37720 6184 37732
rect 4663 37692 6184 37720
rect 4663 37689 4675 37692
rect 4617 37683 4675 37689
rect 6178 37680 6184 37692
rect 6236 37680 6242 37732
rect 6270 37680 6276 37732
rect 6328 37720 6334 37732
rect 7024 37729 7052 37760
rect 7745 37757 7757 37791
rect 7791 37757 7803 37791
rect 7745 37751 7803 37757
rect 8205 37791 8263 37797
rect 8205 37757 8217 37791
rect 8251 37788 8263 37791
rect 8386 37788 8392 37800
rect 8251 37760 8392 37788
rect 8251 37757 8263 37760
rect 8205 37751 8263 37757
rect 6549 37723 6607 37729
rect 6549 37720 6561 37723
rect 6328 37692 6561 37720
rect 6328 37680 6334 37692
rect 6549 37689 6561 37692
rect 6595 37689 6607 37723
rect 6549 37683 6607 37689
rect 7009 37723 7067 37729
rect 7009 37689 7021 37723
rect 7055 37689 7067 37723
rect 7009 37683 7067 37689
rect 7225 37723 7283 37729
rect 7225 37689 7237 37723
rect 7271 37720 7283 37723
rect 7760 37720 7788 37751
rect 8386 37748 8392 37760
rect 8444 37748 8450 37800
rect 8680 37797 8708 37828
rect 8665 37791 8723 37797
rect 8665 37757 8677 37791
rect 8711 37757 8723 37791
rect 8665 37751 8723 37757
rect 8757 37791 8815 37797
rect 8757 37757 8769 37791
rect 8803 37757 8815 37791
rect 8757 37751 8815 37757
rect 7271 37692 7604 37720
rect 7760 37692 8294 37720
rect 7271 37689 7283 37692
rect 7225 37683 7283 37689
rect 1118 37612 1124 37664
rect 1176 37612 1182 37664
rect 1397 37655 1455 37661
rect 1397 37621 1409 37655
rect 1443 37652 1455 37655
rect 1670 37652 1676 37664
rect 1443 37624 1676 37652
rect 1443 37621 1455 37624
rect 1397 37615 1455 37621
rect 1670 37612 1676 37624
rect 1728 37612 1734 37664
rect 3050 37612 3056 37664
rect 3108 37652 3114 37664
rect 3697 37655 3755 37661
rect 3697 37652 3709 37655
rect 3108 37624 3709 37652
rect 3108 37612 3114 37624
rect 3697 37621 3709 37624
rect 3743 37621 3755 37655
rect 3697 37615 3755 37621
rect 4246 37612 4252 37664
rect 4304 37612 4310 37664
rect 4706 37612 4712 37664
rect 4764 37612 4770 37664
rect 6365 37655 6423 37661
rect 6365 37621 6377 37655
rect 6411 37652 6423 37655
rect 6730 37652 6736 37664
rect 6411 37624 6736 37652
rect 6411 37621 6423 37624
rect 6365 37615 6423 37621
rect 6730 37612 6736 37624
rect 6788 37612 6794 37664
rect 7576 37661 7604 37692
rect 7561 37655 7619 37661
rect 7561 37621 7573 37655
rect 7607 37621 7619 37655
rect 8266 37652 8294 37692
rect 8772 37664 8800 37751
rect 8864 37720 8892 37828
rect 8941 37825 8953 37859
rect 8987 37856 8999 37859
rect 9508 37856 9536 37896
rect 10502 37884 10508 37896
rect 10560 37884 10566 37936
rect 8987 37828 9536 37856
rect 9585 37859 9643 37865
rect 8987 37825 8999 37828
rect 8941 37819 8999 37825
rect 9585 37825 9597 37859
rect 9631 37856 9643 37859
rect 9858 37856 9864 37868
rect 9631 37828 9864 37856
rect 9631 37825 9643 37828
rect 9585 37819 9643 37825
rect 9858 37816 9864 37828
rect 9916 37816 9922 37868
rect 9122 37748 9128 37800
rect 9180 37748 9186 37800
rect 9398 37797 9404 37800
rect 9383 37791 9404 37797
rect 9383 37757 9395 37791
rect 9383 37751 9404 37757
rect 9398 37748 9404 37751
rect 9456 37748 9462 37800
rect 9950 37788 9956 37800
rect 9784 37760 9956 37788
rect 9784 37720 9812 37760
rect 9950 37748 9956 37760
rect 10008 37748 10014 37800
rect 10502 37748 10508 37800
rect 10560 37788 10566 37800
rect 10689 37791 10747 37797
rect 10689 37788 10701 37791
rect 10560 37760 10701 37788
rect 10560 37748 10566 37760
rect 10689 37757 10701 37760
rect 10735 37757 10747 37791
rect 10689 37751 10747 37757
rect 8864 37692 9812 37720
rect 9858 37680 9864 37732
rect 9916 37720 9922 37732
rect 10410 37720 10416 37732
rect 9916 37692 10416 37720
rect 9916 37680 9922 37692
rect 10410 37680 10416 37692
rect 10468 37680 10474 37732
rect 8662 37652 8668 37664
rect 8266 37624 8668 37652
rect 7561 37615 7619 37621
rect 8662 37612 8668 37624
rect 8720 37612 8726 37664
rect 8754 37612 8760 37664
rect 8812 37612 8818 37664
rect 9217 37655 9275 37661
rect 9217 37621 9229 37655
rect 9263 37652 9275 37655
rect 9306 37652 9312 37664
rect 9263 37624 9312 37652
rect 9263 37621 9275 37624
rect 9217 37615 9275 37621
rect 9306 37612 9312 37624
rect 9364 37612 9370 37664
rect 9398 37612 9404 37664
rect 9456 37652 9462 37664
rect 10137 37655 10195 37661
rect 10137 37652 10149 37655
rect 9456 37624 10149 37652
rect 9456 37612 9462 37624
rect 10137 37621 10149 37624
rect 10183 37621 10195 37655
rect 10137 37615 10195 37621
rect 552 37562 11132 37584
rect 552 37510 4322 37562
rect 4374 37510 4386 37562
rect 4438 37510 4450 37562
rect 4502 37510 4514 37562
rect 4566 37510 4578 37562
rect 4630 37510 10722 37562
rect 10774 37510 10786 37562
rect 10838 37510 10850 37562
rect 10902 37510 10914 37562
rect 10966 37510 10978 37562
rect 11030 37510 11132 37562
rect 552 37488 11132 37510
rect 1026 37408 1032 37460
rect 1084 37448 1090 37460
rect 2869 37451 2927 37457
rect 2869 37448 2881 37451
rect 1084 37420 2881 37448
rect 1084 37408 1090 37420
rect 2869 37417 2881 37420
rect 2915 37417 2927 37451
rect 2869 37411 2927 37417
rect 3326 37408 3332 37460
rect 3384 37448 3390 37460
rect 4249 37451 4307 37457
rect 4249 37448 4261 37451
rect 3384 37420 4261 37448
rect 3384 37408 3390 37420
rect 4249 37417 4261 37420
rect 4295 37417 4307 37451
rect 4249 37411 4307 37417
rect 4709 37451 4767 37457
rect 4709 37417 4721 37451
rect 4755 37448 4767 37451
rect 5077 37451 5135 37457
rect 5077 37448 5089 37451
rect 4755 37420 5089 37448
rect 4755 37417 4767 37420
rect 4709 37411 4767 37417
rect 5077 37417 5089 37420
rect 5123 37417 5135 37451
rect 5077 37411 5135 37417
rect 5810 37408 5816 37460
rect 5868 37408 5874 37460
rect 6178 37408 6184 37460
rect 6236 37448 6242 37460
rect 6549 37451 6607 37457
rect 6549 37448 6561 37451
rect 6236 37420 6561 37448
rect 6236 37408 6242 37420
rect 6549 37417 6561 37420
rect 6595 37417 6607 37451
rect 6549 37411 6607 37417
rect 6914 37408 6920 37460
rect 6972 37448 6978 37460
rect 7834 37448 7840 37460
rect 6972 37420 7840 37448
rect 6972 37408 6978 37420
rect 7834 37408 7840 37420
rect 7892 37408 7898 37460
rect 8202 37408 8208 37460
rect 8260 37408 8266 37460
rect 8754 37408 8760 37460
rect 8812 37448 8818 37460
rect 8849 37451 8907 37457
rect 8849 37448 8861 37451
rect 8812 37420 8861 37448
rect 8812 37408 8818 37420
rect 8849 37417 8861 37420
rect 8895 37417 8907 37451
rect 8849 37411 8907 37417
rect 9122 37408 9128 37460
rect 9180 37448 9186 37460
rect 9180 37420 9536 37448
rect 9180 37408 9186 37420
rect 1305 37383 1363 37389
rect 1305 37349 1317 37383
rect 1351 37380 1363 37383
rect 1578 37380 1584 37392
rect 1351 37352 1584 37380
rect 1351 37349 1363 37352
rect 1305 37343 1363 37349
rect 1578 37340 1584 37352
rect 1636 37340 1642 37392
rect 3418 37340 3424 37392
rect 3476 37380 3482 37392
rect 3789 37383 3847 37389
rect 3476 37352 3740 37380
rect 3476 37340 3482 37352
rect 1118 37272 1124 37324
rect 1176 37272 1182 37324
rect 1397 37315 1455 37321
rect 1397 37281 1409 37315
rect 1443 37312 1455 37315
rect 1486 37312 1492 37324
rect 1443 37284 1492 37312
rect 1443 37281 1455 37284
rect 1397 37275 1455 37281
rect 1486 37272 1492 37284
rect 1544 37272 1550 37324
rect 1670 37321 1676 37324
rect 1664 37312 1676 37321
rect 1631 37284 1676 37312
rect 1664 37275 1676 37284
rect 1670 37272 1676 37275
rect 1728 37272 1734 37324
rect 2866 37272 2872 37324
rect 2924 37312 2930 37324
rect 3712 37321 3740 37352
rect 3789 37349 3801 37383
rect 3835 37380 3847 37383
rect 5828 37380 5856 37408
rect 3835 37352 5856 37380
rect 3835 37349 3847 37352
rect 3789 37343 3847 37349
rect 6086 37340 6092 37392
rect 6144 37380 6150 37392
rect 6457 37383 6515 37389
rect 6457 37380 6469 37383
rect 6144 37352 6469 37380
rect 6144 37340 6150 37352
rect 6457 37349 6469 37352
rect 6503 37349 6515 37383
rect 6457 37343 6515 37349
rect 7190 37340 7196 37392
rect 7248 37380 7254 37392
rect 9033 37383 9091 37389
rect 7248 37352 7788 37380
rect 7248 37340 7254 37352
rect 3237 37315 3295 37321
rect 3237 37312 3249 37315
rect 2924 37284 3249 37312
rect 2924 37272 2930 37284
rect 3237 37281 3249 37284
rect 3283 37281 3295 37315
rect 3237 37275 3295 37281
rect 3697 37315 3755 37321
rect 3697 37281 3709 37315
rect 3743 37281 3755 37315
rect 3697 37275 3755 37281
rect 3878 37272 3884 37324
rect 3936 37272 3942 37324
rect 3970 37272 3976 37324
rect 4028 37272 4034 37324
rect 4154 37272 4160 37324
rect 4212 37272 4218 37324
rect 4617 37315 4675 37321
rect 4617 37281 4629 37315
rect 4663 37312 4675 37315
rect 5166 37312 5172 37324
rect 4663 37284 5172 37312
rect 4663 37281 4675 37284
rect 4617 37275 4675 37281
rect 5166 37272 5172 37284
rect 5224 37272 5230 37324
rect 5258 37272 5264 37324
rect 5316 37272 5322 37324
rect 5350 37272 5356 37324
rect 5408 37272 5414 37324
rect 5442 37272 5448 37324
rect 5500 37272 5506 37324
rect 5626 37272 5632 37324
rect 5684 37272 5690 37324
rect 5813 37315 5871 37321
rect 5813 37281 5825 37315
rect 5859 37281 5871 37315
rect 5813 37275 5871 37281
rect 5997 37315 6055 37321
rect 5997 37281 6009 37315
rect 6043 37281 6055 37315
rect 5997 37275 6055 37281
rect 937 37247 995 37253
rect 937 37213 949 37247
rect 983 37244 995 37247
rect 983 37216 1440 37244
rect 983 37213 995 37216
rect 937 37207 995 37213
rect 1412 37108 1440 37216
rect 2682 37204 2688 37256
rect 2740 37244 2746 37256
rect 3329 37247 3387 37253
rect 3329 37244 3341 37247
rect 2740 37216 3341 37244
rect 2740 37204 2746 37216
rect 3329 37213 3341 37216
rect 3375 37213 3387 37247
rect 3329 37207 3387 37213
rect 3418 37204 3424 37256
rect 3476 37204 3482 37256
rect 4798 37204 4804 37256
rect 4856 37244 4862 37256
rect 5074 37244 5080 37256
rect 4856 37216 5080 37244
rect 4856 37204 4862 37216
rect 5074 37204 5080 37216
rect 5132 37204 5138 37256
rect 2777 37179 2835 37185
rect 2777 37145 2789 37179
rect 2823 37176 2835 37179
rect 4157 37179 4215 37185
rect 2823 37148 4108 37176
rect 2823 37145 2835 37148
rect 2777 37139 2835 37145
rect 1762 37108 1768 37120
rect 1412 37080 1768 37108
rect 1762 37068 1768 37080
rect 1820 37068 1826 37120
rect 4080 37108 4108 37148
rect 4157 37145 4169 37179
rect 4203 37176 4215 37179
rect 5534 37176 5540 37188
rect 4203 37148 5540 37176
rect 4203 37145 4215 37148
rect 4157 37139 4215 37145
rect 5534 37136 5540 37148
rect 5592 37176 5598 37188
rect 5828 37176 5856 37275
rect 6012 37244 6040 37275
rect 6270 37272 6276 37324
rect 6328 37272 6334 37324
rect 6638 37272 6644 37324
rect 6696 37312 6702 37324
rect 7285 37315 7343 37321
rect 7285 37312 7297 37315
rect 6696 37284 7297 37312
rect 6696 37272 6702 37284
rect 7285 37281 7297 37284
rect 7331 37281 7343 37315
rect 7285 37275 7343 37281
rect 7374 37272 7380 37324
rect 7432 37312 7438 37324
rect 7469 37315 7527 37321
rect 7469 37312 7481 37315
rect 7432 37284 7481 37312
rect 7432 37272 7438 37284
rect 7469 37281 7481 37284
rect 7515 37281 7527 37315
rect 7469 37275 7527 37281
rect 7650 37272 7656 37324
rect 7708 37272 7714 37324
rect 7760 37312 7788 37352
rect 9033 37349 9045 37383
rect 9079 37380 9091 37383
rect 9214 37380 9220 37392
rect 9079 37352 9220 37380
rect 9079 37349 9091 37352
rect 9033 37343 9091 37349
rect 9214 37340 9220 37352
rect 9272 37340 9278 37392
rect 9508 37389 9536 37420
rect 9484 37383 9542 37389
rect 9484 37349 9496 37383
rect 9530 37349 9542 37383
rect 9484 37343 9542 37349
rect 8297 37315 8355 37321
rect 7760 37284 8156 37312
rect 6546 37244 6552 37256
rect 6012 37216 6552 37244
rect 6546 37204 6552 37216
rect 6604 37204 6610 37256
rect 6914 37204 6920 37256
rect 6972 37244 6978 37256
rect 7193 37247 7251 37253
rect 7193 37244 7205 37247
rect 6972 37216 7205 37244
rect 6972 37204 6978 37216
rect 7193 37213 7205 37216
rect 7239 37244 7251 37247
rect 7929 37247 7987 37253
rect 7239 37216 7880 37244
rect 7239 37213 7251 37216
rect 7193 37207 7251 37213
rect 5592 37148 5856 37176
rect 5592 37136 5598 37148
rect 7006 37136 7012 37188
rect 7064 37176 7070 37188
rect 7374 37176 7380 37188
rect 7064 37148 7380 37176
rect 7064 37136 7070 37148
rect 7374 37136 7380 37148
rect 7432 37176 7438 37188
rect 7852 37176 7880 37216
rect 7929 37213 7941 37247
rect 7975 37244 7987 37247
rect 8018 37244 8024 37256
rect 7975 37216 8024 37244
rect 7975 37213 7987 37216
rect 7929 37207 7987 37213
rect 8018 37204 8024 37216
rect 8076 37204 8082 37256
rect 8128 37244 8156 37284
rect 8297 37281 8309 37315
rect 8343 37312 8355 37315
rect 8386 37312 8392 37324
rect 8343 37284 8392 37312
rect 8343 37281 8355 37284
rect 8297 37275 8355 37281
rect 8386 37272 8392 37284
rect 8444 37272 8450 37324
rect 8846 37272 8852 37324
rect 8904 37312 8910 37324
rect 8941 37315 8999 37321
rect 8941 37312 8953 37315
rect 8904 37284 8953 37312
rect 8904 37272 8910 37284
rect 8941 37281 8953 37284
rect 8987 37281 8999 37315
rect 8941 37275 8999 37281
rect 9125 37315 9183 37321
rect 9125 37281 9137 37315
rect 9171 37312 9183 37315
rect 11054 37312 11060 37324
rect 9171 37284 11060 37312
rect 9171 37281 9183 37284
rect 9125 37275 9183 37281
rect 11054 37272 11060 37284
rect 11112 37272 11118 37324
rect 8573 37247 8631 37253
rect 8573 37244 8585 37247
rect 8128 37216 8585 37244
rect 8573 37213 8585 37216
rect 8619 37213 8631 37247
rect 8573 37207 8631 37213
rect 9217 37247 9275 37253
rect 9217 37213 9229 37247
rect 9263 37213 9275 37247
rect 9217 37207 9275 37213
rect 8110 37176 8116 37188
rect 7432 37148 7788 37176
rect 7852 37148 8116 37176
rect 7432 37136 7438 37148
rect 4614 37108 4620 37120
rect 4080 37080 4620 37108
rect 4614 37068 4620 37080
rect 4672 37068 4678 37120
rect 6454 37068 6460 37120
rect 6512 37108 6518 37120
rect 7760 37117 7788 37148
rect 8110 37136 8116 37148
rect 8168 37136 8174 37188
rect 7285 37111 7343 37117
rect 7285 37108 7297 37111
rect 6512 37080 7297 37108
rect 6512 37068 6518 37080
rect 7285 37077 7297 37080
rect 7331 37077 7343 37111
rect 7285 37071 7343 37077
rect 7745 37111 7803 37117
rect 7745 37077 7757 37111
rect 7791 37077 7803 37111
rect 7745 37071 7803 37077
rect 8294 37068 8300 37120
rect 8352 37108 8358 37120
rect 8389 37111 8447 37117
rect 8389 37108 8401 37111
rect 8352 37080 8401 37108
rect 8352 37068 8358 37080
rect 8389 37077 8401 37080
rect 8435 37077 8447 37111
rect 8588 37108 8616 37207
rect 8938 37136 8944 37188
rect 8996 37176 9002 37188
rect 9232 37176 9260 37207
rect 8996 37148 9260 37176
rect 8996 37136 9002 37148
rect 10502 37108 10508 37120
rect 8588 37080 10508 37108
rect 8389 37071 8447 37077
rect 10502 37068 10508 37080
rect 10560 37108 10566 37120
rect 10597 37111 10655 37117
rect 10597 37108 10609 37111
rect 10560 37080 10609 37108
rect 10560 37068 10566 37080
rect 10597 37077 10609 37080
rect 10643 37077 10655 37111
rect 10597 37071 10655 37077
rect 552 37018 11132 37040
rect 552 36966 3662 37018
rect 3714 36966 3726 37018
rect 3778 36966 3790 37018
rect 3842 36966 3854 37018
rect 3906 36966 3918 37018
rect 3970 36966 10062 37018
rect 10114 36966 10126 37018
rect 10178 36966 10190 37018
rect 10242 36966 10254 37018
rect 10306 36966 10318 37018
rect 10370 36966 11132 37018
rect 552 36944 11132 36966
rect 1029 36907 1087 36913
rect 1029 36873 1041 36907
rect 1075 36904 1087 36907
rect 1118 36904 1124 36916
rect 1075 36876 1124 36904
rect 1075 36873 1087 36876
rect 1029 36867 1087 36873
rect 1118 36864 1124 36876
rect 1176 36864 1182 36916
rect 4706 36864 4712 36916
rect 4764 36904 4770 36916
rect 5445 36907 5503 36913
rect 5445 36904 5457 36907
rect 4764 36876 5457 36904
rect 4764 36864 4770 36876
rect 5445 36873 5457 36876
rect 5491 36873 5503 36907
rect 5445 36867 5503 36873
rect 5552 36876 6040 36904
rect 5552 36836 5580 36876
rect 5000 36808 5580 36836
rect 1213 36771 1271 36777
rect 1213 36737 1225 36771
rect 1259 36768 1271 36771
rect 1394 36768 1400 36780
rect 1259 36740 1400 36768
rect 1259 36737 1271 36740
rect 1213 36731 1271 36737
rect 1394 36728 1400 36740
rect 1452 36728 1458 36780
rect 3326 36728 3332 36780
rect 3384 36728 3390 36780
rect 937 36703 995 36709
rect 937 36669 949 36703
rect 983 36669 995 36703
rect 937 36663 995 36669
rect 952 36632 980 36663
rect 1026 36660 1032 36712
rect 1084 36700 1090 36712
rect 1121 36703 1179 36709
rect 1121 36700 1133 36703
rect 1084 36672 1133 36700
rect 1084 36660 1090 36672
rect 1121 36669 1133 36672
rect 1167 36669 1179 36703
rect 1121 36663 1179 36669
rect 1489 36703 1547 36709
rect 1489 36669 1501 36703
rect 1535 36700 1547 36703
rect 1762 36700 1768 36712
rect 1535 36672 1768 36700
rect 1535 36669 1547 36672
rect 1489 36663 1547 36669
rect 1762 36660 1768 36672
rect 1820 36660 1826 36712
rect 3973 36703 4031 36709
rect 3973 36669 3985 36703
rect 4019 36700 4031 36703
rect 4062 36700 4068 36712
rect 4019 36672 4068 36700
rect 4019 36669 4031 36672
rect 3973 36663 4031 36669
rect 4062 36660 4068 36672
rect 4120 36660 4126 36712
rect 4246 36709 4252 36712
rect 4240 36700 4252 36709
rect 4207 36672 4252 36700
rect 4240 36663 4252 36672
rect 4246 36660 4252 36663
rect 4304 36660 4310 36712
rect 1302 36632 1308 36644
rect 952 36604 1308 36632
rect 1302 36592 1308 36604
rect 1360 36592 1366 36644
rect 2866 36592 2872 36644
rect 2924 36592 2930 36644
rect 3510 36592 3516 36644
rect 3568 36632 3574 36644
rect 5000 36632 5028 36808
rect 5902 36768 5908 36780
rect 5736 36740 5908 36768
rect 5350 36660 5356 36712
rect 5408 36660 5414 36712
rect 5629 36703 5687 36709
rect 5629 36669 5641 36703
rect 5675 36700 5687 36703
rect 5736 36700 5764 36740
rect 5902 36728 5908 36740
rect 5960 36728 5966 36780
rect 5675 36672 5764 36700
rect 5675 36669 5687 36672
rect 5629 36663 5687 36669
rect 5810 36660 5816 36712
rect 5868 36660 5874 36712
rect 6012 36709 6040 36876
rect 9122 36864 9128 36916
rect 9180 36904 9186 36916
rect 9493 36907 9551 36913
rect 9493 36904 9505 36907
rect 9180 36876 9505 36904
rect 9180 36864 9186 36876
rect 9493 36873 9505 36876
rect 9539 36873 9551 36907
rect 9493 36867 9551 36873
rect 9858 36864 9864 36916
rect 9916 36904 9922 36916
rect 10318 36904 10324 36916
rect 9916 36876 10324 36904
rect 9916 36864 9922 36876
rect 10318 36864 10324 36876
rect 10376 36864 10382 36916
rect 7285 36839 7343 36845
rect 7285 36805 7297 36839
rect 7331 36836 7343 36839
rect 7374 36836 7380 36848
rect 7331 36808 7380 36836
rect 7331 36805 7343 36808
rect 7285 36799 7343 36805
rect 7374 36796 7380 36808
rect 7432 36796 7438 36848
rect 7926 36796 7932 36848
rect 7984 36796 7990 36848
rect 9033 36839 9091 36845
rect 9033 36805 9045 36839
rect 9079 36836 9091 36839
rect 9674 36836 9680 36848
rect 9079 36808 9680 36836
rect 9079 36805 9091 36808
rect 9033 36799 9091 36805
rect 9674 36796 9680 36808
rect 9732 36796 9738 36848
rect 10137 36839 10195 36845
rect 10137 36805 10149 36839
rect 10183 36836 10195 36839
rect 10594 36836 10600 36848
rect 10183 36808 10600 36836
rect 10183 36805 10195 36808
rect 10137 36799 10195 36805
rect 6086 36728 6092 36780
rect 6144 36768 6150 36780
rect 7944 36768 7972 36796
rect 8481 36771 8539 36777
rect 6144 36740 7880 36768
rect 7944 36740 8064 36768
rect 6144 36728 6150 36740
rect 5997 36703 6055 36709
rect 5997 36669 6009 36703
rect 6043 36669 6055 36703
rect 5997 36663 6055 36669
rect 6178 36660 6184 36712
rect 6236 36660 6242 36712
rect 6546 36660 6552 36712
rect 6604 36660 6610 36712
rect 7190 36660 7196 36712
rect 7248 36700 7254 36712
rect 7469 36703 7527 36709
rect 7469 36700 7481 36703
rect 7248 36672 7481 36700
rect 7248 36660 7254 36672
rect 7469 36669 7481 36672
rect 7515 36669 7527 36703
rect 7745 36703 7803 36709
rect 7745 36700 7757 36703
rect 7469 36663 7527 36669
rect 7576 36672 7757 36700
rect 3568 36604 5028 36632
rect 5368 36632 5396 36660
rect 5721 36635 5779 36641
rect 5721 36632 5733 36635
rect 5368 36604 5733 36632
rect 3568 36592 3574 36604
rect 5721 36601 5733 36604
rect 5767 36632 5779 36635
rect 6638 36632 6644 36644
rect 5767 36604 6644 36632
rect 5767 36601 5779 36604
rect 5721 36595 5779 36601
rect 6638 36592 6644 36604
rect 6696 36592 6702 36644
rect 7098 36592 7104 36644
rect 7156 36632 7162 36644
rect 7576 36632 7604 36672
rect 7745 36669 7757 36672
rect 7791 36669 7803 36703
rect 7745 36663 7803 36669
rect 7156 36604 7604 36632
rect 7653 36635 7711 36641
rect 7156 36592 7162 36604
rect 7653 36601 7665 36635
rect 7699 36632 7711 36635
rect 7852 36632 7880 36740
rect 7926 36660 7932 36712
rect 7984 36660 7990 36712
rect 8036 36709 8064 36740
rect 8481 36737 8493 36771
rect 8527 36768 8539 36771
rect 9401 36771 9459 36777
rect 8527 36740 9168 36768
rect 8527 36737 8539 36740
rect 8481 36731 8539 36737
rect 9140 36712 9168 36740
rect 9401 36737 9413 36771
rect 9447 36768 9459 36771
rect 10152 36768 10180 36799
rect 10594 36796 10600 36808
rect 10652 36796 10658 36848
rect 11238 36768 11244 36780
rect 9447 36740 10180 36768
rect 10612 36740 11244 36768
rect 9447 36737 9459 36740
rect 9401 36731 9459 36737
rect 8021 36703 8079 36709
rect 8021 36669 8033 36703
rect 8067 36669 8079 36703
rect 8021 36663 8079 36669
rect 8386 36660 8392 36712
rect 8444 36660 8450 36712
rect 8573 36703 8631 36709
rect 8573 36669 8585 36703
rect 8619 36700 8631 36703
rect 8754 36700 8760 36712
rect 8619 36672 8760 36700
rect 8619 36669 8631 36672
rect 8573 36663 8631 36669
rect 8754 36660 8760 36672
rect 8812 36700 8818 36712
rect 8812 36672 9076 36700
rect 8812 36660 8818 36672
rect 8404 36632 8432 36660
rect 7699 36604 8432 36632
rect 7699 36601 7711 36604
rect 7653 36595 7711 36601
rect 8662 36592 8668 36644
rect 8720 36592 8726 36644
rect 8849 36635 8907 36641
rect 8849 36601 8861 36635
rect 8895 36601 8907 36635
rect 9048 36632 9076 36672
rect 9122 36660 9128 36712
rect 9180 36660 9186 36712
rect 9306 36660 9312 36712
rect 9364 36700 9370 36712
rect 9493 36703 9551 36709
rect 9493 36700 9505 36703
rect 9364 36672 9505 36700
rect 9364 36660 9370 36672
rect 9493 36669 9505 36672
rect 9539 36669 9551 36703
rect 9493 36663 9551 36669
rect 9600 36672 10088 36700
rect 9600 36632 9628 36672
rect 9048 36604 9628 36632
rect 8849 36595 8907 36601
rect 3878 36524 3884 36576
rect 3936 36524 3942 36576
rect 5353 36567 5411 36573
rect 5353 36533 5365 36567
rect 5399 36564 5411 36567
rect 6914 36564 6920 36576
rect 5399 36536 6920 36564
rect 5399 36533 5411 36536
rect 5353 36527 5411 36533
rect 6914 36524 6920 36536
rect 6972 36524 6978 36576
rect 7193 36567 7251 36573
rect 7193 36533 7205 36567
rect 7239 36564 7251 36567
rect 7558 36564 7564 36576
rect 7239 36536 7564 36564
rect 7239 36533 7251 36536
rect 7193 36527 7251 36533
rect 7558 36524 7564 36536
rect 7616 36524 7622 36576
rect 7742 36524 7748 36576
rect 7800 36564 7806 36576
rect 7837 36567 7895 36573
rect 7837 36564 7849 36567
rect 7800 36536 7849 36564
rect 7800 36524 7806 36536
rect 7837 36533 7849 36536
rect 7883 36533 7895 36567
rect 7837 36527 7895 36533
rect 8202 36524 8208 36576
rect 8260 36524 8266 36576
rect 8294 36524 8300 36576
rect 8352 36564 8358 36576
rect 8864 36564 8892 36595
rect 9858 36592 9864 36644
rect 9916 36592 9922 36644
rect 10060 36641 10088 36672
rect 10134 36660 10140 36712
rect 10192 36700 10198 36712
rect 10612 36709 10640 36740
rect 11238 36728 11244 36740
rect 11296 36728 11302 36780
rect 10597 36703 10655 36709
rect 10597 36700 10609 36703
rect 10192 36672 10609 36700
rect 10192 36660 10198 36672
rect 10597 36669 10609 36672
rect 10643 36669 10655 36703
rect 10597 36663 10655 36669
rect 10686 36660 10692 36712
rect 10744 36700 10750 36712
rect 10781 36703 10839 36709
rect 10781 36700 10793 36703
rect 10744 36672 10793 36700
rect 10744 36660 10750 36672
rect 10781 36669 10793 36672
rect 10827 36669 10839 36703
rect 10781 36663 10839 36669
rect 10045 36635 10103 36641
rect 10045 36601 10057 36635
rect 10091 36632 10103 36635
rect 10289 36635 10347 36641
rect 10289 36632 10301 36635
rect 10091 36604 10301 36632
rect 10091 36601 10103 36604
rect 10045 36595 10103 36601
rect 10289 36601 10301 36604
rect 10335 36601 10347 36635
rect 10289 36595 10347 36601
rect 10502 36592 10508 36644
rect 10560 36592 10566 36644
rect 8352 36536 8892 36564
rect 8352 36524 8358 36536
rect 9214 36524 9220 36576
rect 9272 36564 9278 36576
rect 9490 36564 9496 36576
rect 9272 36536 9496 36564
rect 9272 36524 9278 36536
rect 9490 36524 9496 36536
rect 9548 36524 9554 36576
rect 9674 36524 9680 36576
rect 9732 36524 9738 36576
rect 9950 36524 9956 36576
rect 10008 36564 10014 36576
rect 10689 36567 10747 36573
rect 10689 36564 10701 36567
rect 10008 36536 10701 36564
rect 10008 36524 10014 36536
rect 10689 36533 10701 36536
rect 10735 36533 10747 36567
rect 10689 36527 10747 36533
rect 552 36474 11132 36496
rect 552 36422 4322 36474
rect 4374 36422 4386 36474
rect 4438 36422 4450 36474
rect 4502 36422 4514 36474
rect 4566 36422 4578 36474
rect 4630 36422 10722 36474
rect 10774 36422 10786 36474
rect 10838 36422 10850 36474
rect 10902 36422 10914 36474
rect 10966 36422 10978 36474
rect 11030 36422 11132 36474
rect 552 36400 11132 36422
rect 2409 36363 2467 36369
rect 2409 36329 2421 36363
rect 2455 36360 2467 36363
rect 2682 36360 2688 36372
rect 2455 36332 2688 36360
rect 2455 36329 2467 36332
rect 2409 36323 2467 36329
rect 2682 36320 2688 36332
rect 2740 36320 2746 36372
rect 3329 36363 3387 36369
rect 3329 36329 3341 36363
rect 3375 36329 3387 36363
rect 3329 36323 3387 36329
rect 1394 36292 1400 36304
rect 1044 36264 1400 36292
rect 1044 36233 1072 36264
rect 1394 36252 1400 36264
rect 1452 36252 1458 36304
rect 1762 36252 1768 36304
rect 1820 36292 1826 36304
rect 3344 36292 3372 36323
rect 3786 36320 3792 36372
rect 3844 36320 3850 36372
rect 5166 36320 5172 36372
rect 5224 36360 5230 36372
rect 5353 36363 5411 36369
rect 5353 36360 5365 36363
rect 5224 36332 5365 36360
rect 5224 36320 5230 36332
rect 5353 36329 5365 36332
rect 5399 36329 5411 36363
rect 5353 36323 5411 36329
rect 5537 36363 5595 36369
rect 5537 36329 5549 36363
rect 5583 36360 5595 36363
rect 6178 36360 6184 36372
rect 5583 36332 6184 36360
rect 5583 36329 5595 36332
rect 5537 36323 5595 36329
rect 6178 36320 6184 36332
rect 6236 36320 6242 36372
rect 6546 36320 6552 36372
rect 6604 36360 6610 36372
rect 7561 36363 7619 36369
rect 7561 36360 7573 36363
rect 6604 36332 7573 36360
rect 6604 36320 6610 36332
rect 7561 36329 7573 36332
rect 7607 36329 7619 36363
rect 7561 36323 7619 36329
rect 7926 36320 7932 36372
rect 7984 36360 7990 36372
rect 8205 36363 8263 36369
rect 8205 36360 8217 36363
rect 7984 36332 8217 36360
rect 7984 36320 7990 36332
rect 8205 36329 8217 36332
rect 8251 36329 8263 36363
rect 8205 36323 8263 36329
rect 8386 36320 8392 36372
rect 8444 36320 8450 36372
rect 9122 36320 9128 36372
rect 9180 36369 9186 36372
rect 9180 36363 9199 36369
rect 9187 36329 9199 36363
rect 9180 36323 9199 36329
rect 9180 36320 9186 36323
rect 10318 36320 10324 36372
rect 10376 36360 10382 36372
rect 10781 36363 10839 36369
rect 10781 36360 10793 36363
rect 10376 36332 10793 36360
rect 10376 36320 10382 36332
rect 10781 36329 10793 36332
rect 10827 36329 10839 36363
rect 10781 36323 10839 36329
rect 1820 36264 3372 36292
rect 1820 36252 1826 36264
rect 3418 36252 3424 36304
rect 3476 36292 3482 36304
rect 3476 36264 3832 36292
rect 3476 36252 3482 36264
rect 1029 36227 1087 36233
rect 1029 36193 1041 36227
rect 1075 36193 1087 36227
rect 1029 36187 1087 36193
rect 1118 36184 1124 36236
rect 1176 36224 1182 36236
rect 1285 36227 1343 36233
rect 1285 36224 1297 36227
rect 1176 36196 1297 36224
rect 1176 36184 1182 36196
rect 1285 36193 1297 36196
rect 1331 36193 1343 36227
rect 1285 36187 1343 36193
rect 2866 36184 2872 36236
rect 2924 36184 2930 36236
rect 2961 36227 3019 36233
rect 2961 36193 2973 36227
rect 3007 36224 3019 36227
rect 3142 36224 3148 36236
rect 3007 36196 3148 36224
rect 3007 36193 3019 36196
rect 2961 36187 3019 36193
rect 3142 36184 3148 36196
rect 3200 36184 3206 36236
rect 2222 36116 2228 36168
rect 2280 36156 2286 36168
rect 2777 36159 2835 36165
rect 2777 36156 2789 36159
rect 2280 36128 2789 36156
rect 2280 36116 2286 36128
rect 2777 36125 2789 36128
rect 2823 36156 2835 36159
rect 3436 36156 3464 36252
rect 3510 36184 3516 36236
rect 3568 36224 3574 36236
rect 3804 36233 3832 36264
rect 3878 36252 3884 36304
rect 3936 36292 3942 36304
rect 4218 36295 4276 36301
rect 4218 36292 4230 36295
rect 3936 36264 4230 36292
rect 3936 36252 3942 36264
rect 4218 36261 4230 36264
rect 4264 36261 4276 36295
rect 6270 36292 6276 36304
rect 4218 36255 4276 36261
rect 5644 36264 6276 36292
rect 3605 36227 3663 36233
rect 3605 36224 3617 36227
rect 3568 36196 3617 36224
rect 3568 36184 3574 36196
rect 3605 36193 3617 36196
rect 3651 36193 3663 36227
rect 3605 36187 3663 36193
rect 3789 36227 3847 36233
rect 3789 36193 3801 36227
rect 3835 36224 3847 36227
rect 3973 36227 4031 36233
rect 3835 36196 3924 36224
rect 3835 36193 3847 36196
rect 3789 36187 3847 36193
rect 2823 36128 3464 36156
rect 2823 36125 2835 36128
rect 2777 36119 2835 36125
rect 1026 35980 1032 36032
rect 1084 36020 1090 36032
rect 3142 36020 3148 36032
rect 1084 35992 3148 36020
rect 1084 35980 1090 35992
rect 3142 35980 3148 35992
rect 3200 35980 3206 36032
rect 3896 36020 3924 36196
rect 3973 36193 3985 36227
rect 4019 36224 4031 36227
rect 4062 36224 4068 36236
rect 4019 36196 4068 36224
rect 4019 36193 4031 36196
rect 3973 36187 4031 36193
rect 4062 36184 4068 36196
rect 4120 36184 4126 36236
rect 5445 36227 5503 36233
rect 5445 36193 5457 36227
rect 5491 36224 5503 36227
rect 5534 36224 5540 36236
rect 5491 36196 5540 36224
rect 5491 36193 5503 36196
rect 5445 36187 5503 36193
rect 5534 36184 5540 36196
rect 5592 36184 5598 36236
rect 5644 36233 5672 36264
rect 6270 36252 6276 36264
rect 6328 36252 6334 36304
rect 8404 36292 8432 36320
rect 6564 36264 7880 36292
rect 5629 36227 5687 36233
rect 5629 36193 5641 36227
rect 5675 36193 5687 36227
rect 5997 36227 6055 36233
rect 5997 36224 6009 36227
rect 5629 36187 5687 36193
rect 5736 36196 6009 36224
rect 4890 36020 4896 36032
rect 3896 35992 4896 36020
rect 4890 35980 4896 35992
rect 4948 36020 4954 36032
rect 5350 36020 5356 36032
rect 4948 35992 5356 36020
rect 4948 35980 4954 35992
rect 5350 35980 5356 35992
rect 5408 35980 5414 36032
rect 5736 36020 5764 36196
rect 5997 36193 6009 36196
rect 6043 36193 6055 36227
rect 5997 36187 6055 36193
rect 6086 36184 6092 36236
rect 6144 36184 6150 36236
rect 5813 36159 5871 36165
rect 5813 36125 5825 36159
rect 5859 36156 5871 36159
rect 6104 36156 6132 36184
rect 5859 36128 6132 36156
rect 5859 36125 5871 36128
rect 5813 36119 5871 36125
rect 6270 36116 6276 36168
rect 6328 36116 6334 36168
rect 6454 36116 6460 36168
rect 6512 36156 6518 36168
rect 6564 36156 6592 36264
rect 7742 36224 7748 36236
rect 7222 36196 7748 36224
rect 7742 36184 7748 36196
rect 7800 36184 7806 36236
rect 7852 36233 7880 36264
rect 8312 36264 8432 36292
rect 7837 36227 7895 36233
rect 7837 36193 7849 36227
rect 7883 36193 7895 36227
rect 7837 36187 7895 36193
rect 8110 36184 8116 36236
rect 8168 36184 8174 36236
rect 8312 36233 8340 36264
rect 8938 36252 8944 36304
rect 8996 36252 9002 36304
rect 9646 36295 9704 36301
rect 9646 36292 9658 36295
rect 9324 36264 9658 36292
rect 8297 36227 8355 36233
rect 8297 36193 8309 36227
rect 8343 36193 8355 36227
rect 8297 36187 8355 36193
rect 8389 36227 8447 36233
rect 8389 36193 8401 36227
rect 8435 36224 8447 36227
rect 8478 36224 8484 36236
rect 8435 36196 8484 36224
rect 8435 36193 8447 36196
rect 8389 36187 8447 36193
rect 8478 36184 8484 36196
rect 8536 36184 8542 36236
rect 8573 36227 8631 36233
rect 8573 36193 8585 36227
rect 8619 36193 8631 36227
rect 8573 36187 8631 36193
rect 7101 36159 7159 36165
rect 7101 36156 7113 36159
rect 6512 36128 7113 36156
rect 6512 36116 6518 36128
rect 7101 36125 7113 36128
rect 7147 36125 7159 36159
rect 7101 36119 7159 36125
rect 7469 36159 7527 36165
rect 7469 36125 7481 36159
rect 7515 36125 7527 36159
rect 7760 36156 7788 36184
rect 8021 36159 8079 36165
rect 8021 36156 8033 36159
rect 7760 36128 8033 36156
rect 7469 36119 7527 36125
rect 8021 36125 8033 36128
rect 8067 36125 8079 36159
rect 8021 36119 8079 36125
rect 6181 36091 6239 36097
rect 6181 36057 6193 36091
rect 6227 36088 6239 36091
rect 7484 36088 7512 36119
rect 8588 36088 8616 36187
rect 8662 36184 8668 36236
rect 8720 36224 8726 36236
rect 9122 36224 9128 36236
rect 8720 36196 9128 36224
rect 8720 36184 8726 36196
rect 9122 36184 9128 36196
rect 9180 36184 9186 36236
rect 9324 36214 9352 36264
rect 9646 36261 9658 36264
rect 9692 36261 9704 36295
rect 9646 36255 9704 36261
rect 9232 36186 9352 36214
rect 6227 36060 7512 36088
rect 7576 36060 8616 36088
rect 9232 36088 9260 36186
rect 9398 36184 9404 36236
rect 9456 36184 9462 36236
rect 9490 36184 9496 36236
rect 9548 36224 9554 36236
rect 9950 36224 9956 36236
rect 9548 36196 9956 36224
rect 9548 36184 9554 36196
rect 9950 36184 9956 36196
rect 10008 36184 10014 36236
rect 9309 36091 9367 36097
rect 9309 36088 9321 36091
rect 9232 36060 9321 36088
rect 6227 36057 6239 36060
rect 6181 36051 6239 36057
rect 7116 36032 7144 36060
rect 6914 36020 6920 36032
rect 5736 35992 6920 36020
rect 6914 35980 6920 35992
rect 6972 35980 6978 36032
rect 7098 35980 7104 36032
rect 7156 35980 7162 36032
rect 7466 35980 7472 36032
rect 7524 36020 7530 36032
rect 7576 36020 7604 36060
rect 9309 36057 9321 36060
rect 9355 36057 9367 36091
rect 9309 36051 9367 36057
rect 7524 35992 7604 36020
rect 7524 35980 7530 35992
rect 8386 35980 8392 36032
rect 8444 36020 8450 36032
rect 8573 36023 8631 36029
rect 8573 36020 8585 36023
rect 8444 35992 8585 36020
rect 8444 35980 8450 35992
rect 8573 35989 8585 35992
rect 8619 35989 8631 36023
rect 8573 35983 8631 35989
rect 8662 35980 8668 36032
rect 8720 36020 8726 36032
rect 8757 36023 8815 36029
rect 8757 36020 8769 36023
rect 8720 35992 8769 36020
rect 8720 35980 8726 35992
rect 8757 35989 8769 35992
rect 8803 36020 8815 36023
rect 9030 36020 9036 36032
rect 8803 35992 9036 36020
rect 8803 35989 8815 35992
rect 8757 35983 8815 35989
rect 9030 35980 9036 35992
rect 9088 35980 9094 36032
rect 9125 36023 9183 36029
rect 9125 35989 9137 36023
rect 9171 36020 9183 36023
rect 9674 36020 9680 36032
rect 9171 35992 9680 36020
rect 9171 35989 9183 35992
rect 9125 35983 9183 35989
rect 9674 35980 9680 35992
rect 9732 35980 9738 36032
rect 552 35930 11132 35952
rect 552 35878 3662 35930
rect 3714 35878 3726 35930
rect 3778 35878 3790 35930
rect 3842 35878 3854 35930
rect 3906 35878 3918 35930
rect 3970 35878 10062 35930
rect 10114 35878 10126 35930
rect 10178 35878 10190 35930
rect 10242 35878 10254 35930
rect 10306 35878 10318 35930
rect 10370 35878 11132 35930
rect 552 35856 11132 35878
rect 1397 35819 1455 35825
rect 1397 35785 1409 35819
rect 1443 35816 1455 35819
rect 3878 35816 3884 35828
rect 1443 35788 3884 35816
rect 1443 35785 1455 35788
rect 1397 35779 1455 35785
rect 3878 35776 3884 35788
rect 3936 35776 3942 35828
rect 3970 35776 3976 35828
rect 4028 35816 4034 35828
rect 5442 35816 5448 35828
rect 4028 35788 5448 35816
rect 4028 35776 4034 35788
rect 5442 35776 5448 35788
rect 5500 35816 5506 35828
rect 7282 35816 7288 35828
rect 5500 35788 7288 35816
rect 5500 35776 5506 35788
rect 7282 35776 7288 35788
rect 7340 35776 7346 35828
rect 7834 35776 7840 35828
rect 7892 35816 7898 35828
rect 8481 35819 8539 35825
rect 8481 35816 8493 35819
rect 7892 35788 8493 35816
rect 7892 35776 7898 35788
rect 8481 35785 8493 35788
rect 8527 35785 8539 35819
rect 8481 35779 8539 35785
rect 8754 35776 8760 35828
rect 8812 35816 8818 35828
rect 9214 35816 9220 35828
rect 8812 35788 9220 35816
rect 8812 35776 8818 35788
rect 9214 35776 9220 35788
rect 9272 35776 9278 35828
rect 9585 35819 9643 35825
rect 9585 35785 9597 35819
rect 9631 35816 9643 35819
rect 10045 35819 10103 35825
rect 10045 35816 10057 35819
rect 9631 35788 10057 35816
rect 9631 35785 9643 35788
rect 9585 35779 9643 35785
rect 10045 35785 10057 35788
rect 10091 35785 10103 35819
rect 10045 35779 10103 35785
rect 3421 35751 3479 35757
rect 3421 35717 3433 35751
rect 3467 35748 3479 35751
rect 4062 35748 4068 35760
rect 3467 35720 4068 35748
rect 3467 35717 3479 35720
rect 3421 35711 3479 35717
rect 4062 35708 4068 35720
rect 4120 35708 4126 35760
rect 5721 35751 5779 35757
rect 5721 35717 5733 35751
rect 5767 35748 5779 35751
rect 5767 35720 6224 35748
rect 5767 35717 5779 35720
rect 5721 35711 5779 35717
rect 1121 35683 1179 35689
rect 1121 35649 1133 35683
rect 1167 35680 1179 35683
rect 1167 35652 1440 35680
rect 1167 35649 1179 35652
rect 1121 35643 1179 35649
rect 1029 35615 1087 35621
rect 1029 35581 1041 35615
rect 1075 35612 1087 35615
rect 1302 35612 1308 35624
rect 1075 35584 1308 35612
rect 1075 35581 1087 35584
rect 1029 35575 1087 35581
rect 1302 35572 1308 35584
rect 1360 35572 1366 35624
rect 1412 35544 1440 35652
rect 1486 35640 1492 35692
rect 1544 35640 1550 35692
rect 3697 35683 3755 35689
rect 3697 35649 3709 35683
rect 3743 35680 3755 35683
rect 4246 35680 4252 35692
rect 3743 35652 4252 35680
rect 3743 35649 3755 35652
rect 3697 35643 3755 35649
rect 4246 35640 4252 35652
rect 4304 35640 4310 35692
rect 6196 35624 6224 35720
rect 6638 35708 6644 35760
rect 6696 35748 6702 35760
rect 9600 35748 9628 35779
rect 6696 35720 9628 35748
rect 6696 35708 6702 35720
rect 8113 35683 8171 35689
rect 6932 35652 7972 35680
rect 1578 35572 1584 35624
rect 1636 35612 1642 35624
rect 1745 35615 1803 35621
rect 1745 35612 1757 35615
rect 1636 35584 1757 35612
rect 1636 35572 1642 35584
rect 1745 35581 1757 35584
rect 1791 35581 1803 35615
rect 1745 35575 1803 35581
rect 3513 35615 3571 35621
rect 3513 35581 3525 35615
rect 3559 35612 3571 35615
rect 3970 35612 3976 35624
rect 3559 35584 3976 35612
rect 3559 35581 3571 35584
rect 3513 35575 3571 35581
rect 3970 35572 3976 35584
rect 4028 35572 4034 35624
rect 4154 35572 4160 35624
rect 4212 35612 4218 35624
rect 4341 35615 4399 35621
rect 4341 35612 4353 35615
rect 4212 35584 4353 35612
rect 4212 35572 4218 35584
rect 4341 35581 4353 35584
rect 4387 35581 4399 35615
rect 4341 35575 4399 35581
rect 5166 35572 5172 35624
rect 5224 35572 5230 35624
rect 6178 35572 6184 35624
rect 6236 35612 6242 35624
rect 6365 35615 6423 35621
rect 6365 35612 6377 35615
rect 6236 35584 6377 35612
rect 6236 35572 6242 35584
rect 6365 35581 6377 35584
rect 6411 35581 6423 35615
rect 6932 35612 6960 35652
rect 7944 35621 7972 35652
rect 8113 35649 8125 35683
rect 8159 35680 8171 35683
rect 8294 35680 8300 35692
rect 8159 35652 8300 35680
rect 8159 35649 8171 35652
rect 8113 35643 8171 35649
rect 6365 35575 6423 35581
rect 6472 35598 6960 35612
rect 7561 35615 7619 35621
rect 6472 35584 6946 35598
rect 1412 35516 1808 35544
rect 1780 35488 1808 35516
rect 3050 35504 3056 35556
rect 3108 35544 3114 35556
rect 4249 35547 4307 35553
rect 3108 35516 4200 35544
rect 3108 35504 3114 35516
rect 1762 35436 1768 35488
rect 1820 35436 1826 35488
rect 2869 35479 2927 35485
rect 2869 35445 2881 35479
rect 2915 35476 2927 35479
rect 3142 35476 3148 35488
rect 2915 35448 3148 35476
rect 2915 35445 2927 35448
rect 2869 35439 2927 35445
rect 3142 35436 3148 35448
rect 3200 35436 3206 35488
rect 4172 35476 4200 35516
rect 4249 35513 4261 35547
rect 4295 35544 4307 35547
rect 4586 35547 4644 35553
rect 4586 35544 4598 35547
rect 4295 35516 4598 35544
rect 4295 35513 4307 35516
rect 4249 35507 4307 35513
rect 4586 35513 4598 35516
rect 4632 35513 4644 35547
rect 5184 35544 5212 35572
rect 6472 35544 6500 35584
rect 7561 35581 7573 35615
rect 7607 35581 7619 35615
rect 7561 35575 7619 35581
rect 7929 35615 7987 35621
rect 7929 35581 7941 35615
rect 7975 35581 7987 35615
rect 7929 35575 7987 35581
rect 5184 35516 6500 35544
rect 4586 35507 4644 35513
rect 6546 35504 6552 35556
rect 6604 35504 6610 35556
rect 7576 35544 7604 35575
rect 8128 35544 8156 35643
rect 8294 35640 8300 35652
rect 8352 35680 8358 35692
rect 9030 35680 9036 35692
rect 8352 35652 9036 35680
rect 8352 35640 8358 35652
rect 9030 35640 9036 35652
rect 9088 35680 9094 35692
rect 9125 35683 9183 35689
rect 9125 35680 9137 35683
rect 9088 35652 9137 35680
rect 9088 35640 9094 35652
rect 9125 35649 9137 35652
rect 9171 35649 9183 35683
rect 9125 35643 9183 35649
rect 9214 35640 9220 35692
rect 9272 35640 9278 35692
rect 8570 35572 8576 35624
rect 8628 35572 8634 35624
rect 8938 35572 8944 35624
rect 8996 35572 9002 35624
rect 9674 35572 9680 35624
rect 9732 35612 9738 35624
rect 10505 35615 10563 35621
rect 10505 35612 10517 35615
rect 9732 35584 10517 35612
rect 9732 35572 9738 35584
rect 10505 35581 10517 35584
rect 10551 35581 10563 35615
rect 10505 35575 10563 35581
rect 9953 35547 10011 35553
rect 9953 35544 9965 35547
rect 7576 35516 8156 35544
rect 9508 35516 9965 35544
rect 9508 35488 9536 35516
rect 9953 35513 9965 35516
rect 9999 35513 10011 35547
rect 9953 35507 10011 35513
rect 4798 35476 4804 35488
rect 4172 35448 4804 35476
rect 4798 35436 4804 35448
rect 4856 35436 4862 35488
rect 4982 35436 4988 35488
rect 5040 35476 5046 35488
rect 5166 35476 5172 35488
rect 5040 35448 5172 35476
rect 5040 35436 5046 35448
rect 5166 35436 5172 35448
rect 5224 35436 5230 35488
rect 5810 35436 5816 35488
rect 5868 35436 5874 35488
rect 5994 35436 6000 35488
rect 6052 35476 6058 35488
rect 7745 35479 7803 35485
rect 7745 35476 7757 35479
rect 6052 35448 7757 35476
rect 6052 35436 6058 35448
rect 7745 35445 7757 35448
rect 7791 35445 7803 35479
rect 7745 35439 7803 35445
rect 8202 35436 8208 35488
rect 8260 35476 8266 35488
rect 9490 35476 9496 35488
rect 8260 35448 9496 35476
rect 8260 35436 8266 35448
rect 9490 35436 9496 35448
rect 9548 35436 9554 35488
rect 9582 35436 9588 35488
rect 9640 35436 9646 35488
rect 9766 35436 9772 35488
rect 9824 35436 9830 35488
rect 10410 35436 10416 35488
rect 10468 35476 10474 35488
rect 10597 35479 10655 35485
rect 10597 35476 10609 35479
rect 10468 35448 10609 35476
rect 10468 35436 10474 35448
rect 10597 35445 10609 35448
rect 10643 35445 10655 35479
rect 10597 35439 10655 35445
rect 552 35386 11132 35408
rect 552 35334 4322 35386
rect 4374 35334 4386 35386
rect 4438 35334 4450 35386
rect 4502 35334 4514 35386
rect 4566 35334 4578 35386
rect 4630 35334 10722 35386
rect 10774 35334 10786 35386
rect 10838 35334 10850 35386
rect 10902 35334 10914 35386
rect 10966 35334 10978 35386
rect 11030 35334 11132 35386
rect 552 35312 11132 35334
rect 2774 35232 2780 35284
rect 2832 35272 2838 35284
rect 2869 35275 2927 35281
rect 2869 35272 2881 35275
rect 2832 35244 2881 35272
rect 2832 35232 2838 35244
rect 2869 35241 2881 35244
rect 2915 35241 2927 35275
rect 4065 35275 4123 35281
rect 4065 35272 4077 35275
rect 2869 35235 2927 35241
rect 3068 35244 4077 35272
rect 566 35164 572 35216
rect 624 35204 630 35216
rect 3068 35204 3096 35244
rect 3344 35216 3372 35244
rect 4065 35241 4077 35244
rect 4111 35241 4123 35275
rect 4065 35235 4123 35241
rect 4246 35232 4252 35284
rect 4304 35272 4310 35284
rect 4525 35275 4583 35281
rect 4525 35272 4537 35275
rect 4304 35244 4537 35272
rect 4304 35232 4310 35244
rect 4525 35241 4537 35244
rect 4571 35241 4583 35275
rect 4525 35235 4583 35241
rect 4893 35275 4951 35281
rect 4893 35241 4905 35275
rect 4939 35272 4951 35275
rect 5810 35272 5816 35284
rect 4939 35244 5816 35272
rect 4939 35241 4951 35244
rect 4893 35235 4951 35241
rect 5810 35232 5816 35244
rect 5868 35232 5874 35284
rect 6454 35232 6460 35284
rect 6512 35232 6518 35284
rect 6914 35232 6920 35284
rect 6972 35272 6978 35284
rect 8018 35272 8024 35284
rect 6972 35244 8024 35272
rect 6972 35232 6978 35244
rect 8018 35232 8024 35244
rect 8076 35272 8082 35284
rect 8662 35272 8668 35284
rect 8076 35244 8668 35272
rect 8076 35232 8082 35244
rect 8662 35232 8668 35244
rect 8720 35232 8726 35284
rect 9030 35232 9036 35284
rect 9088 35272 9094 35284
rect 9401 35275 9459 35281
rect 9401 35272 9413 35275
rect 9088 35244 9413 35272
rect 9088 35232 9094 35244
rect 9401 35241 9413 35244
rect 9447 35241 9459 35275
rect 9401 35235 9459 35241
rect 624 35176 3096 35204
rect 624 35164 630 35176
rect 3326 35164 3332 35216
rect 3384 35164 3390 35216
rect 3418 35164 3424 35216
rect 3476 35164 3482 35216
rect 3789 35207 3847 35213
rect 3789 35173 3801 35207
rect 3835 35204 3847 35207
rect 5626 35204 5632 35216
rect 3835 35176 5632 35204
rect 3835 35173 3847 35176
rect 3789 35167 3847 35173
rect 5626 35164 5632 35176
rect 5684 35164 5690 35216
rect 6362 35204 6368 35216
rect 5920 35176 6368 35204
rect 1118 35096 1124 35148
rect 1176 35136 1182 35148
rect 1305 35139 1363 35145
rect 1305 35136 1317 35139
rect 1176 35108 1317 35136
rect 1176 35096 1182 35108
rect 1305 35105 1317 35108
rect 1351 35105 1363 35139
rect 1305 35099 1363 35105
rect 1578 35096 1584 35148
rect 1636 35096 1642 35148
rect 1762 35096 1768 35148
rect 1820 35136 1826 35148
rect 2409 35139 2467 35145
rect 2409 35136 2421 35139
rect 1820 35108 2421 35136
rect 1820 35096 1826 35108
rect 2409 35105 2421 35108
rect 2455 35136 2467 35139
rect 2498 35136 2504 35148
rect 2455 35108 2504 35136
rect 2455 35105 2467 35108
rect 2409 35099 2467 35105
rect 2498 35096 2504 35108
rect 2556 35096 2562 35148
rect 2866 35096 2872 35148
rect 2924 35096 2930 35148
rect 3050 35096 3056 35148
rect 3108 35096 3114 35148
rect 3142 35096 3148 35148
rect 3200 35096 3206 35148
rect 3436 35136 3464 35164
rect 3881 35139 3939 35145
rect 3881 35136 3893 35139
rect 3436 35108 3893 35136
rect 3881 35105 3893 35108
rect 3927 35136 3939 35139
rect 3970 35136 3976 35148
rect 3927 35108 3976 35136
rect 3927 35105 3939 35108
rect 3881 35099 3939 35105
rect 3970 35096 3976 35108
rect 4028 35096 4034 35148
rect 4137 35139 4195 35145
rect 4137 35105 4149 35139
rect 4183 35105 4195 35139
rect 4137 35099 4195 35105
rect 4249 35139 4307 35145
rect 4249 35105 4261 35139
rect 4295 35136 4307 35139
rect 5258 35136 5264 35148
rect 4295 35108 5264 35136
rect 4295 35105 4307 35108
rect 4249 35099 4307 35105
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35068 1731 35071
rect 1854 35068 1860 35080
rect 1719 35040 1860 35068
rect 1719 35037 1731 35040
rect 1673 35031 1731 35037
rect 1854 35028 1860 35040
rect 1912 35028 1918 35080
rect 2222 35028 2228 35080
rect 2280 35028 2286 35080
rect 2314 35028 2320 35080
rect 2372 35068 2378 35080
rect 3418 35068 3424 35080
rect 2372 35040 3424 35068
rect 2372 35028 2378 35040
rect 3418 35028 3424 35040
rect 3476 35028 3482 35080
rect 4152 35068 4180 35099
rect 5258 35096 5264 35108
rect 5316 35096 5322 35148
rect 5353 35139 5411 35145
rect 5353 35105 5365 35139
rect 5399 35136 5411 35139
rect 5442 35136 5448 35148
rect 5399 35108 5448 35136
rect 5399 35105 5411 35108
rect 5353 35099 5411 35105
rect 5442 35096 5448 35108
rect 5500 35096 5506 35148
rect 5537 35139 5595 35145
rect 5537 35105 5549 35139
rect 5583 35136 5595 35139
rect 5920 35136 5948 35176
rect 6362 35164 6368 35176
rect 6420 35164 6426 35216
rect 6733 35207 6791 35213
rect 6733 35173 6745 35207
rect 6779 35204 6791 35207
rect 7190 35204 7196 35216
rect 6779 35176 7196 35204
rect 6779 35173 6791 35176
rect 6733 35167 6791 35173
rect 7190 35164 7196 35176
rect 7248 35164 7254 35216
rect 8573 35207 8631 35213
rect 8573 35173 8585 35207
rect 8619 35204 8631 35207
rect 9122 35204 9128 35216
rect 8619 35176 9128 35204
rect 8619 35173 8631 35176
rect 8573 35167 8631 35173
rect 9122 35164 9128 35176
rect 9180 35164 9186 35216
rect 9766 35164 9772 35216
rect 9824 35204 9830 35216
rect 10514 35207 10572 35213
rect 10514 35204 10526 35207
rect 9824 35176 10526 35204
rect 9824 35164 9830 35176
rect 10514 35173 10526 35176
rect 10560 35173 10572 35207
rect 10514 35167 10572 35173
rect 5583 35108 5948 35136
rect 5583 35105 5595 35108
rect 5537 35099 5595 35105
rect 5994 35096 6000 35148
rect 6052 35096 6058 35148
rect 6089 35139 6147 35145
rect 6089 35105 6101 35139
rect 6135 35136 6147 35139
rect 6638 35136 6644 35148
rect 6135 35108 6644 35136
rect 6135 35105 6147 35108
rect 6089 35099 6147 35105
rect 6638 35096 6644 35108
rect 6696 35096 6702 35148
rect 6822 35096 6828 35148
rect 6880 35096 6886 35148
rect 7374 35096 7380 35148
rect 7432 35096 7438 35148
rect 7466 35096 7472 35148
rect 7524 35136 7530 35148
rect 8113 35139 8171 35145
rect 8113 35136 8125 35139
rect 7524 35108 8125 35136
rect 7524 35096 7530 35108
rect 8113 35105 8125 35108
rect 8159 35136 8171 35139
rect 8202 35136 8208 35148
rect 8159 35108 8208 35136
rect 8159 35105 8171 35108
rect 8113 35099 8171 35105
rect 8202 35096 8208 35108
rect 8260 35096 8266 35148
rect 8294 35096 8300 35148
rect 8352 35096 8358 35148
rect 8846 35136 8852 35148
rect 8404 35108 8852 35136
rect 4338 35068 4344 35080
rect 4152 35040 4344 35068
rect 4338 35028 4344 35040
rect 4396 35028 4402 35080
rect 4982 35028 4988 35080
rect 5040 35028 5046 35080
rect 5074 35028 5080 35080
rect 5132 35028 5138 35080
rect 6178 35028 6184 35080
rect 6236 35028 6242 35080
rect 6273 35071 6331 35077
rect 6273 35037 6285 35071
rect 6319 35068 6331 35071
rect 6546 35068 6552 35080
rect 6319 35040 6552 35068
rect 6319 35037 6331 35040
rect 6273 35031 6331 35037
rect 6546 35028 6552 35040
rect 6604 35068 6610 35080
rect 7101 35071 7159 35077
rect 7101 35068 7113 35071
rect 6604 35040 7113 35068
rect 6604 35028 6610 35040
rect 7101 35037 7113 35040
rect 7147 35037 7159 35071
rect 7101 35031 7159 35037
rect 7742 35028 7748 35080
rect 7800 35068 7806 35080
rect 7929 35071 7987 35077
rect 7929 35068 7941 35071
rect 7800 35040 7941 35068
rect 7800 35028 7806 35040
rect 7929 35037 7941 35040
rect 7975 35037 7987 35071
rect 7929 35031 7987 35037
rect 1949 35003 2007 35009
rect 1949 34969 1961 35003
rect 1995 35000 2007 35003
rect 4433 35003 4491 35009
rect 1995 34972 4384 35000
rect 1995 34969 2007 34972
rect 1949 34963 2007 34969
rect 1118 34892 1124 34944
rect 1176 34892 1182 34944
rect 2590 34892 2596 34944
rect 2648 34932 2654 34944
rect 2777 34935 2835 34941
rect 2777 34932 2789 34935
rect 2648 34904 2789 34932
rect 2648 34892 2654 34904
rect 2777 34901 2789 34904
rect 2823 34901 2835 34935
rect 4356 34932 4384 34972
rect 4433 34969 4445 35003
rect 4479 35000 4491 35003
rect 5092 35000 5120 35028
rect 4479 34972 5120 35000
rect 4479 34969 4491 34972
rect 4433 34963 4491 34969
rect 5166 34960 5172 35012
rect 5224 35000 5230 35012
rect 5224 34972 5488 35000
rect 5224 34960 5230 34972
rect 5350 34932 5356 34944
rect 4356 34904 5356 34932
rect 2777 34895 2835 34901
rect 5350 34892 5356 34904
rect 5408 34892 5414 34944
rect 5460 34941 5488 34972
rect 5994 34960 6000 35012
rect 6052 35000 6058 35012
rect 6052 34972 8064 35000
rect 6052 34960 6058 34972
rect 8036 34944 8064 34972
rect 8202 34960 8208 35012
rect 8260 35000 8266 35012
rect 8404 35000 8432 35108
rect 8846 35096 8852 35108
rect 8904 35096 8910 35148
rect 8938 35096 8944 35148
rect 8996 35096 9002 35148
rect 8754 35028 8760 35080
rect 8812 35068 8818 35080
rect 9033 35071 9091 35077
rect 9033 35068 9045 35071
rect 8812 35040 9045 35068
rect 8812 35028 8818 35040
rect 9033 35037 9045 35040
rect 9079 35037 9091 35071
rect 9033 35031 9091 35037
rect 10781 35071 10839 35077
rect 10781 35037 10793 35071
rect 10827 35037 10839 35071
rect 10781 35031 10839 35037
rect 8260 34972 8432 35000
rect 8481 35003 8539 35009
rect 8260 34960 8266 34972
rect 8481 34969 8493 35003
rect 8527 35000 8539 35003
rect 8849 35003 8907 35009
rect 8849 35000 8861 35003
rect 8527 34972 8861 35000
rect 8527 34969 8539 34972
rect 8481 34963 8539 34969
rect 8849 34969 8861 34972
rect 8895 35000 8907 35003
rect 9306 35000 9312 35012
rect 8895 34972 9312 35000
rect 8895 34969 8907 34972
rect 8849 34963 8907 34969
rect 9306 34960 9312 34972
rect 9364 34960 9370 35012
rect 5445 34935 5503 34941
rect 5445 34901 5457 34935
rect 5491 34901 5503 34935
rect 5445 34895 5503 34901
rect 8018 34892 8024 34944
rect 8076 34932 8082 34944
rect 10410 34932 10416 34944
rect 8076 34904 10416 34932
rect 8076 34892 8082 34904
rect 10410 34892 10416 34904
rect 10468 34892 10474 34944
rect 10502 34892 10508 34944
rect 10560 34932 10566 34944
rect 10796 34932 10824 35031
rect 10560 34904 10824 34932
rect 10560 34892 10566 34904
rect 552 34842 11132 34864
rect 552 34790 3662 34842
rect 3714 34790 3726 34842
rect 3778 34790 3790 34842
rect 3842 34790 3854 34842
rect 3906 34790 3918 34842
rect 3970 34790 10062 34842
rect 10114 34790 10126 34842
rect 10178 34790 10190 34842
rect 10242 34790 10254 34842
rect 10306 34790 10318 34842
rect 10370 34790 11132 34842
rect 552 34768 11132 34790
rect 1302 34688 1308 34740
rect 1360 34728 1366 34740
rect 2314 34728 2320 34740
rect 1360 34700 2320 34728
rect 1360 34688 1366 34700
rect 2314 34688 2320 34700
rect 2372 34688 2378 34740
rect 2682 34688 2688 34740
rect 2740 34728 2746 34740
rect 2961 34731 3019 34737
rect 2961 34728 2973 34731
rect 2740 34700 2973 34728
rect 2740 34688 2746 34700
rect 2961 34697 2973 34700
rect 3007 34697 3019 34731
rect 2961 34691 3019 34697
rect 3602 34688 3608 34740
rect 3660 34728 3666 34740
rect 4338 34728 4344 34740
rect 3660 34700 4344 34728
rect 3660 34688 3666 34700
rect 4338 34688 4344 34700
rect 4396 34688 4402 34740
rect 4433 34731 4491 34737
rect 4433 34697 4445 34731
rect 4479 34728 4491 34731
rect 4479 34700 4936 34728
rect 4479 34697 4491 34700
rect 4433 34691 4491 34697
rect 2866 34620 2872 34672
rect 2924 34660 2930 34672
rect 2924 34632 4476 34660
rect 2924 34620 2930 34632
rect 2958 34592 2964 34604
rect 2792 34564 2964 34592
rect 198 34484 204 34536
rect 256 34524 262 34536
rect 474 34524 480 34536
rect 256 34496 480 34524
rect 256 34484 262 34496
rect 474 34484 480 34496
rect 532 34524 538 34536
rect 1121 34527 1179 34533
rect 1121 34524 1133 34527
rect 532 34496 1133 34524
rect 532 34484 538 34496
rect 1121 34493 1133 34496
rect 1167 34493 1179 34527
rect 1121 34487 1179 34493
rect 2429 34527 2487 34533
rect 2429 34493 2441 34527
rect 2475 34524 2487 34527
rect 2590 34524 2596 34536
rect 2475 34496 2596 34524
rect 2475 34493 2487 34496
rect 2429 34487 2487 34493
rect 2590 34484 2596 34496
rect 2648 34484 2654 34536
rect 2792 34533 2820 34564
rect 2958 34552 2964 34564
rect 3016 34552 3022 34604
rect 3970 34552 3976 34604
rect 4028 34592 4034 34604
rect 4246 34592 4252 34604
rect 4028 34564 4252 34592
rect 4028 34552 4034 34564
rect 4246 34552 4252 34564
rect 4304 34552 4310 34604
rect 2685 34527 2743 34533
rect 2685 34493 2697 34527
rect 2731 34493 2743 34527
rect 2685 34487 2743 34493
rect 2777 34527 2835 34533
rect 2777 34493 2789 34527
rect 2823 34493 2835 34527
rect 2777 34487 2835 34493
rect 2700 34456 2728 34487
rect 3050 34484 3056 34536
rect 3108 34524 3114 34536
rect 3329 34527 3387 34533
rect 3329 34524 3341 34527
rect 3108 34496 3341 34524
rect 3108 34484 3114 34496
rect 3329 34493 3341 34496
rect 3375 34493 3387 34527
rect 3329 34487 3387 34493
rect 3418 34484 3424 34536
rect 3476 34524 3482 34536
rect 3786 34524 3792 34536
rect 3476 34496 3792 34524
rect 3476 34484 3482 34496
rect 3786 34484 3792 34496
rect 3844 34484 3850 34536
rect 4062 34484 4068 34536
rect 4120 34484 4126 34536
rect 3142 34456 3148 34468
rect 2700 34428 3148 34456
rect 3142 34416 3148 34428
rect 3200 34416 3206 34468
rect 3510 34416 3516 34468
rect 3568 34416 3574 34468
rect 4448 34456 4476 34632
rect 4614 34620 4620 34672
rect 4672 34660 4678 34672
rect 4672 34632 4752 34660
rect 4672 34620 4678 34632
rect 4525 34527 4583 34533
rect 4525 34493 4537 34527
rect 4571 34524 4583 34527
rect 4614 34524 4620 34536
rect 4571 34496 4620 34524
rect 4571 34493 4583 34496
rect 4525 34487 4583 34493
rect 4614 34484 4620 34496
rect 4672 34484 4678 34536
rect 4724 34533 4752 34632
rect 4908 34592 4936 34700
rect 4982 34688 4988 34740
rect 5040 34728 5046 34740
rect 5077 34731 5135 34737
rect 5077 34728 5089 34731
rect 5040 34700 5089 34728
rect 5040 34688 5046 34700
rect 5077 34697 5089 34700
rect 5123 34697 5135 34731
rect 5077 34691 5135 34697
rect 5166 34688 5172 34740
rect 5224 34688 5230 34740
rect 5258 34688 5264 34740
rect 5316 34728 5322 34740
rect 5537 34731 5595 34737
rect 5537 34728 5549 34731
rect 5316 34700 5549 34728
rect 5316 34688 5322 34700
rect 5537 34697 5549 34700
rect 5583 34697 5595 34731
rect 5537 34691 5595 34697
rect 7101 34731 7159 34737
rect 7101 34697 7113 34731
rect 7147 34728 7159 34731
rect 8938 34728 8944 34740
rect 7147 34700 8944 34728
rect 7147 34697 7159 34700
rect 7101 34691 7159 34697
rect 8938 34688 8944 34700
rect 8996 34688 9002 34740
rect 9306 34688 9312 34740
rect 9364 34728 9370 34740
rect 10045 34731 10103 34737
rect 10045 34728 10057 34731
rect 9364 34700 10057 34728
rect 9364 34688 9370 34700
rect 10045 34697 10057 34700
rect 10091 34697 10103 34731
rect 10045 34691 10103 34697
rect 6178 34620 6184 34672
rect 6236 34660 6242 34672
rect 8386 34660 8392 34672
rect 6236 34632 8392 34660
rect 6236 34620 6242 34632
rect 5261 34595 5319 34601
rect 5261 34592 5273 34595
rect 4908 34564 5273 34592
rect 4709 34527 4767 34533
rect 4709 34493 4721 34527
rect 4755 34493 4767 34527
rect 4709 34487 4767 34493
rect 4798 34484 4804 34536
rect 4856 34484 4862 34536
rect 4908 34533 4936 34564
rect 5261 34561 5273 34564
rect 5307 34561 5319 34595
rect 5261 34555 5319 34561
rect 4893 34527 4951 34533
rect 4893 34493 4905 34527
rect 4939 34493 4951 34527
rect 4893 34487 4951 34493
rect 5169 34527 5227 34533
rect 5169 34493 5181 34527
rect 5215 34524 5227 34527
rect 5350 34524 5356 34536
rect 5215 34496 5356 34524
rect 5215 34493 5227 34496
rect 5169 34487 5227 34493
rect 5350 34484 5356 34496
rect 5408 34484 5414 34536
rect 6270 34484 6276 34536
rect 6328 34484 6334 34536
rect 6457 34527 6515 34533
rect 6457 34493 6469 34527
rect 6503 34524 6515 34527
rect 6564 34524 6592 34632
rect 8386 34620 8392 34632
rect 8444 34620 8450 34672
rect 9950 34620 9956 34672
rect 10008 34660 10014 34672
rect 10505 34663 10563 34669
rect 10505 34660 10517 34663
rect 10008 34632 10517 34660
rect 10008 34620 10014 34632
rect 10505 34629 10517 34632
rect 10551 34629 10563 34663
rect 10505 34623 10563 34629
rect 10781 34663 10839 34669
rect 10781 34629 10793 34663
rect 10827 34660 10839 34663
rect 11054 34660 11060 34672
rect 10827 34632 11060 34660
rect 10827 34629 10839 34632
rect 10781 34623 10839 34629
rect 11054 34620 11060 34632
rect 11112 34620 11118 34672
rect 6825 34595 6883 34601
rect 6825 34561 6837 34595
rect 6871 34592 6883 34595
rect 8481 34595 8539 34601
rect 8481 34592 8493 34595
rect 6871 34564 7604 34592
rect 6871 34561 6883 34564
rect 6825 34555 6883 34561
rect 6503 34496 6592 34524
rect 6503 34493 6515 34496
rect 6457 34487 6515 34493
rect 6638 34484 6644 34536
rect 6696 34484 6702 34536
rect 6914 34484 6920 34536
rect 6972 34484 6978 34536
rect 7101 34527 7159 34533
rect 7101 34493 7113 34527
rect 7147 34524 7159 34527
rect 7282 34524 7288 34536
rect 7147 34496 7288 34524
rect 7147 34493 7159 34496
rect 7101 34487 7159 34493
rect 7282 34484 7288 34496
rect 7340 34484 7346 34536
rect 7374 34484 7380 34536
rect 7432 34524 7438 34536
rect 7576 34533 7604 34564
rect 7668 34564 8493 34592
rect 7469 34527 7527 34533
rect 7469 34524 7481 34527
rect 7432 34496 7481 34524
rect 7432 34484 7438 34496
rect 7469 34493 7481 34496
rect 7515 34493 7527 34527
rect 7469 34487 7527 34493
rect 7561 34527 7619 34533
rect 7561 34493 7573 34527
rect 7607 34493 7619 34527
rect 7561 34487 7619 34493
rect 5258 34456 5264 34468
rect 4448 34428 5264 34456
rect 5258 34416 5264 34428
rect 5316 34416 5322 34468
rect 7484 34456 7512 34487
rect 7668 34456 7696 34564
rect 8481 34561 8493 34564
rect 8527 34561 8539 34595
rect 10410 34592 10416 34604
rect 8481 34555 8539 34561
rect 10336 34564 10416 34592
rect 10336 34536 10364 34564
rect 10410 34552 10416 34564
rect 10468 34552 10474 34604
rect 7745 34527 7803 34533
rect 7745 34493 7757 34527
rect 7791 34524 7803 34527
rect 7834 34524 7840 34536
rect 7791 34496 7840 34524
rect 7791 34493 7803 34496
rect 7745 34487 7803 34493
rect 7834 34484 7840 34496
rect 7892 34484 7898 34536
rect 8018 34484 8024 34536
rect 8076 34484 8082 34536
rect 8110 34484 8116 34536
rect 8168 34524 8174 34536
rect 8205 34527 8263 34533
rect 8205 34524 8217 34527
rect 8168 34496 8217 34524
rect 8168 34484 8174 34496
rect 8205 34493 8217 34496
rect 8251 34493 8263 34527
rect 8205 34487 8263 34493
rect 8386 34484 8392 34536
rect 8444 34484 8450 34536
rect 8570 34484 8576 34536
rect 8628 34484 8634 34536
rect 8662 34484 8668 34536
rect 8720 34524 8726 34536
rect 8720 34496 9076 34524
rect 8720 34484 8726 34496
rect 7484 34428 7696 34456
rect 7760 34428 8524 34456
rect 934 34348 940 34400
rect 992 34348 998 34400
rect 2774 34348 2780 34400
rect 2832 34388 2838 34400
rect 3528 34388 3556 34416
rect 2832 34360 3556 34388
rect 2832 34348 2838 34360
rect 4890 34348 4896 34400
rect 4948 34388 4954 34400
rect 5442 34388 5448 34400
rect 4948 34360 5448 34388
rect 4948 34348 4954 34360
rect 5442 34348 5448 34360
rect 5500 34348 5506 34400
rect 5626 34348 5632 34400
rect 5684 34388 5690 34400
rect 5721 34391 5779 34397
rect 5721 34388 5733 34391
rect 5684 34360 5733 34388
rect 5684 34348 5690 34360
rect 5721 34357 5733 34360
rect 5767 34357 5779 34391
rect 5721 34351 5779 34357
rect 6546 34348 6552 34400
rect 6604 34388 6610 34400
rect 7760 34388 7788 34428
rect 6604 34360 7788 34388
rect 8205 34391 8263 34397
rect 6604 34348 6610 34360
rect 8205 34357 8217 34391
rect 8251 34388 8263 34391
rect 8386 34388 8392 34400
rect 8251 34360 8392 34388
rect 8251 34357 8263 34360
rect 8205 34351 8263 34357
rect 8386 34348 8392 34360
rect 8444 34348 8450 34400
rect 8496 34388 8524 34428
rect 8754 34416 8760 34468
rect 8812 34456 8818 34468
rect 8910 34459 8968 34465
rect 8910 34456 8922 34459
rect 8812 34428 8922 34456
rect 8812 34416 8818 34428
rect 8910 34425 8922 34428
rect 8956 34425 8968 34459
rect 9048 34456 9076 34496
rect 10134 34484 10140 34536
rect 10192 34524 10198 34536
rect 10229 34527 10287 34533
rect 10229 34524 10241 34527
rect 10192 34496 10241 34524
rect 10192 34484 10198 34496
rect 10229 34493 10241 34496
rect 10275 34493 10287 34527
rect 10229 34487 10287 34493
rect 10318 34484 10324 34536
rect 10376 34484 10382 34536
rect 10594 34484 10600 34536
rect 10652 34484 10658 34536
rect 10781 34527 10839 34533
rect 10781 34493 10793 34527
rect 10827 34524 10839 34527
rect 10962 34524 10968 34536
rect 10827 34496 10968 34524
rect 10827 34493 10839 34496
rect 10781 34487 10839 34493
rect 10962 34484 10968 34496
rect 11020 34484 11026 34536
rect 9398 34456 9404 34468
rect 9048 34428 9404 34456
rect 8910 34419 8968 34425
rect 9398 34416 9404 34428
rect 9456 34456 9462 34468
rect 10410 34456 10416 34468
rect 9456 34428 10416 34456
rect 9456 34416 9462 34428
rect 10410 34416 10416 34428
rect 10468 34416 10474 34468
rect 10505 34459 10563 34465
rect 10505 34425 10517 34459
rect 10551 34425 10563 34459
rect 10505 34419 10563 34425
rect 10226 34388 10232 34400
rect 8496 34360 10232 34388
rect 10226 34348 10232 34360
rect 10284 34348 10290 34400
rect 10520 34388 10548 34419
rect 10594 34388 10600 34400
rect 10520 34360 10600 34388
rect 10594 34348 10600 34360
rect 10652 34348 10658 34400
rect 552 34298 11132 34320
rect 552 34246 4322 34298
rect 4374 34246 4386 34298
rect 4438 34246 4450 34298
rect 4502 34246 4514 34298
rect 4566 34246 4578 34298
rect 4630 34246 10722 34298
rect 10774 34246 10786 34298
rect 10838 34246 10850 34298
rect 10902 34246 10914 34298
rect 10966 34246 10978 34298
rect 11030 34246 11132 34298
rect 552 34224 11132 34246
rect 5350 34184 5356 34196
rect 5092 34156 5356 34184
rect 1026 34076 1032 34128
rect 1084 34116 1090 34128
rect 1084 34088 2452 34116
rect 1084 34076 1090 34088
rect 1572 34051 1630 34057
rect 1572 34017 1584 34051
rect 1618 34048 1630 34051
rect 1946 34048 1952 34060
rect 1618 34020 1952 34048
rect 1618 34017 1630 34020
rect 1572 34011 1630 34017
rect 1946 34008 1952 34020
rect 2004 34008 2010 34060
rect 1302 33940 1308 33992
rect 1360 33940 1366 33992
rect 2424 33980 2452 34088
rect 2498 34076 2504 34128
rect 2556 34116 2562 34128
rect 2556 34088 4844 34116
rect 2556 34076 2562 34088
rect 3418 34057 3424 34060
rect 3412 34011 3424 34057
rect 3418 34008 3424 34011
rect 3476 34008 3482 34060
rect 2424 33952 3104 33980
rect 1578 33804 1584 33856
rect 1636 33844 1642 33856
rect 2498 33844 2504 33856
rect 1636 33816 2504 33844
rect 1636 33804 1642 33816
rect 2498 33804 2504 33816
rect 2556 33844 2562 33856
rect 2685 33847 2743 33853
rect 2685 33844 2697 33847
rect 2556 33816 2697 33844
rect 2556 33804 2562 33816
rect 2685 33813 2697 33816
rect 2731 33844 2743 33847
rect 2958 33844 2964 33856
rect 2731 33816 2964 33844
rect 2731 33813 2743 33816
rect 2685 33807 2743 33813
rect 2958 33804 2964 33816
rect 3016 33804 3022 33856
rect 3076 33844 3104 33952
rect 3142 33940 3148 33992
rect 3200 33940 3206 33992
rect 4522 33872 4528 33924
rect 4580 33872 4586 33924
rect 4816 33912 4844 34088
rect 4890 34008 4896 34060
rect 4948 34008 4954 34060
rect 5092 34057 5120 34156
rect 5350 34144 5356 34156
rect 5408 34144 5414 34196
rect 5813 34187 5871 34193
rect 5813 34153 5825 34187
rect 5859 34184 5871 34187
rect 6270 34184 6276 34196
rect 5859 34156 6276 34184
rect 5859 34153 5871 34156
rect 5813 34147 5871 34153
rect 6270 34144 6276 34156
rect 6328 34144 6334 34196
rect 7561 34187 7619 34193
rect 7561 34153 7573 34187
rect 7607 34184 7619 34187
rect 7607 34156 8800 34184
rect 7607 34153 7619 34156
rect 7561 34147 7619 34153
rect 8662 34116 8668 34128
rect 7208 34088 8668 34116
rect 5077 34051 5135 34057
rect 5077 34017 5089 34051
rect 5123 34017 5135 34051
rect 5077 34011 5135 34017
rect 5166 34008 5172 34060
rect 5224 34008 5230 34060
rect 5258 34008 5264 34060
rect 5316 34048 5322 34060
rect 5353 34051 5411 34057
rect 5353 34048 5365 34051
rect 5316 34020 5365 34048
rect 5316 34008 5322 34020
rect 5353 34017 5365 34020
rect 5399 34017 5411 34051
rect 5353 34011 5411 34017
rect 5626 34008 5632 34060
rect 5684 34008 5690 34060
rect 5810 34008 5816 34060
rect 5868 34048 5874 34060
rect 6926 34051 6984 34057
rect 6926 34048 6938 34051
rect 5868 34020 6938 34048
rect 5868 34008 5874 34020
rect 6926 34017 6938 34020
rect 6972 34017 6984 34051
rect 6926 34011 6984 34017
rect 7098 34008 7104 34060
rect 7156 34008 7162 34060
rect 7208 34057 7236 34088
rect 8662 34076 8668 34088
rect 8720 34076 8726 34128
rect 8772 34060 8800 34156
rect 8846 34144 8852 34196
rect 8904 34144 8910 34196
rect 8938 34144 8944 34196
rect 8996 34184 9002 34196
rect 8996 34156 9260 34184
rect 8996 34144 9002 34156
rect 9232 34125 9260 34156
rect 9398 34144 9404 34196
rect 9456 34144 9462 34196
rect 9582 34144 9588 34196
rect 9640 34144 9646 34196
rect 10413 34187 10471 34193
rect 10413 34153 10425 34187
rect 10459 34184 10471 34187
rect 10594 34184 10600 34196
rect 10459 34156 10600 34184
rect 10459 34153 10471 34156
rect 10413 34147 10471 34153
rect 10594 34144 10600 34156
rect 10652 34144 10658 34196
rect 9217 34119 9275 34125
rect 9217 34085 9229 34119
rect 9263 34085 9275 34119
rect 9416 34116 9444 34144
rect 10137 34119 10195 34125
rect 10137 34116 10149 34119
rect 9416 34088 10149 34116
rect 9217 34079 9275 34085
rect 10137 34085 10149 34088
rect 10183 34085 10195 34119
rect 10137 34079 10195 34085
rect 7193 34051 7251 34057
rect 7193 34017 7205 34051
rect 7239 34017 7251 34051
rect 7193 34011 7251 34017
rect 7374 34008 7380 34060
rect 7432 34048 7438 34060
rect 7745 34051 7803 34057
rect 7745 34048 7757 34051
rect 7432 34020 7757 34048
rect 7432 34008 7438 34020
rect 7745 34017 7757 34020
rect 7791 34017 7803 34051
rect 7745 34011 7803 34017
rect 7834 34008 7840 34060
rect 7892 34008 7898 34060
rect 8021 34051 8079 34057
rect 8021 34017 8033 34051
rect 8067 34048 8079 34051
rect 8478 34048 8484 34060
rect 8067 34020 8484 34048
rect 8067 34017 8079 34020
rect 8021 34011 8079 34017
rect 4985 33983 5043 33989
rect 4985 33949 4997 33983
rect 5031 33980 5043 33983
rect 6086 33980 6092 33992
rect 5031 33952 6092 33980
rect 5031 33949 5043 33952
rect 4985 33943 5043 33949
rect 6086 33940 6092 33952
rect 6144 33940 6150 33992
rect 7116 33980 7144 34008
rect 8036 33980 8064 34011
rect 8478 34008 8484 34020
rect 8536 34008 8542 34060
rect 8573 34051 8631 34057
rect 8573 34017 8585 34051
rect 8619 34048 8631 34051
rect 8754 34048 8760 34060
rect 8619 34020 8760 34048
rect 8619 34017 8631 34020
rect 8573 34011 8631 34017
rect 8754 34008 8760 34020
rect 8812 34008 8818 34060
rect 8938 34008 8944 34060
rect 8996 34008 9002 34060
rect 9030 34008 9036 34060
rect 9088 34048 9094 34060
rect 9401 34051 9459 34057
rect 9401 34048 9413 34051
rect 9088 34020 9413 34048
rect 9088 34008 9094 34020
rect 9401 34017 9413 34020
rect 9447 34017 9459 34051
rect 9401 34011 9459 34017
rect 9766 34008 9772 34060
rect 9824 34048 9830 34060
rect 9861 34051 9919 34057
rect 9861 34048 9873 34051
rect 9824 34020 9873 34048
rect 9824 34008 9830 34020
rect 9861 34017 9873 34020
rect 9907 34017 9919 34051
rect 9861 34011 9919 34017
rect 10318 34008 10324 34060
rect 10376 34048 10382 34060
rect 10689 34051 10747 34057
rect 10689 34048 10701 34051
rect 10376 34020 10701 34048
rect 10376 34008 10382 34020
rect 10689 34017 10701 34020
rect 10735 34017 10747 34051
rect 10689 34011 10747 34017
rect 7116 33952 8064 33980
rect 8202 33940 8208 33992
rect 8260 33940 8266 33992
rect 8846 33980 8852 33992
rect 8312 33952 8852 33980
rect 5537 33915 5595 33921
rect 5537 33912 5549 33915
rect 4816 33884 5549 33912
rect 5537 33881 5549 33884
rect 5583 33912 5595 33915
rect 5718 33912 5724 33924
rect 5583 33884 5724 33912
rect 5583 33881 5595 33884
rect 5537 33875 5595 33881
rect 5718 33872 5724 33884
rect 5776 33872 5782 33924
rect 8113 33915 8171 33921
rect 8113 33881 8125 33915
rect 8159 33912 8171 33915
rect 8312 33912 8340 33952
rect 8846 33940 8852 33952
rect 8904 33980 8910 33992
rect 9677 33983 9735 33989
rect 9677 33980 9689 33983
rect 8904 33952 9689 33980
rect 8904 33940 8910 33952
rect 9677 33949 9689 33952
rect 9723 33949 9735 33983
rect 9677 33943 9735 33949
rect 10413 33983 10471 33989
rect 10413 33949 10425 33983
rect 10459 33980 10471 33983
rect 10459 33952 10732 33980
rect 10459 33949 10471 33952
rect 10413 33943 10471 33949
rect 10704 33924 10732 33952
rect 8159 33884 8340 33912
rect 8389 33915 8447 33921
rect 8159 33881 8171 33884
rect 8113 33875 8171 33881
rect 8389 33881 8401 33915
rect 8435 33912 8447 33915
rect 8435 33884 8616 33912
rect 8435 33881 8447 33884
rect 8389 33875 8447 33881
rect 5261 33847 5319 33853
rect 5261 33844 5273 33847
rect 3076 33816 5273 33844
rect 5261 33813 5273 33816
rect 5307 33813 5319 33847
rect 5261 33807 5319 33813
rect 5994 33804 6000 33856
rect 6052 33844 6058 33856
rect 6822 33844 6828 33856
rect 6052 33816 6828 33844
rect 6052 33804 6058 33816
rect 6822 33804 6828 33816
rect 6880 33804 6886 33856
rect 6914 33804 6920 33856
rect 6972 33844 6978 33856
rect 7650 33844 7656 33856
rect 6972 33816 7656 33844
rect 6972 33804 6978 33816
rect 7650 33804 7656 33816
rect 7708 33804 7714 33856
rect 8202 33804 8208 33856
rect 8260 33804 8266 33856
rect 8588 33844 8616 33884
rect 9306 33872 9312 33924
rect 9364 33912 9370 33924
rect 10134 33912 10140 33924
rect 9364 33884 10140 33912
rect 9364 33872 9370 33884
rect 10134 33872 10140 33884
rect 10192 33912 10198 33924
rect 10597 33915 10655 33921
rect 10597 33912 10609 33915
rect 10192 33884 10609 33912
rect 10192 33872 10198 33884
rect 10597 33881 10609 33884
rect 10643 33881 10655 33915
rect 10597 33875 10655 33881
rect 10686 33872 10692 33924
rect 10744 33872 10750 33924
rect 8754 33844 8760 33856
rect 8588 33816 8760 33844
rect 8754 33804 8760 33816
rect 8812 33804 8818 33856
rect 10226 33804 10232 33856
rect 10284 33844 10290 33856
rect 10410 33844 10416 33856
rect 10284 33816 10416 33844
rect 10284 33804 10290 33816
rect 10410 33804 10416 33816
rect 10468 33804 10474 33856
rect 552 33754 11132 33776
rect 552 33702 3662 33754
rect 3714 33702 3726 33754
rect 3778 33702 3790 33754
rect 3842 33702 3854 33754
rect 3906 33702 3918 33754
rect 3970 33702 10062 33754
rect 10114 33702 10126 33754
rect 10178 33702 10190 33754
rect 10242 33702 10254 33754
rect 10306 33702 10318 33754
rect 10370 33702 11132 33754
rect 552 33680 11132 33702
rect 1946 33600 1952 33652
rect 2004 33600 2010 33652
rect 3418 33600 3424 33652
rect 3476 33640 3482 33652
rect 3513 33643 3571 33649
rect 3513 33640 3525 33643
rect 3476 33612 3525 33640
rect 3476 33600 3482 33612
rect 3513 33609 3525 33612
rect 3559 33609 3571 33643
rect 3513 33603 3571 33609
rect 5261 33643 5319 33649
rect 5261 33609 5273 33643
rect 5307 33640 5319 33643
rect 5534 33640 5540 33652
rect 5307 33612 5540 33640
rect 5307 33609 5319 33612
rect 5261 33603 5319 33609
rect 5534 33600 5540 33612
rect 5592 33600 5598 33652
rect 6914 33640 6920 33652
rect 5920 33612 6920 33640
rect 2314 33532 2320 33584
rect 2372 33572 2378 33584
rect 2777 33575 2835 33581
rect 2777 33572 2789 33575
rect 2372 33544 2789 33572
rect 2372 33532 2378 33544
rect 2777 33541 2789 33544
rect 2823 33541 2835 33575
rect 2777 33535 2835 33541
rect 5445 33575 5503 33581
rect 5445 33541 5457 33575
rect 5491 33572 5503 33575
rect 5920 33572 5948 33612
rect 6914 33600 6920 33612
rect 6972 33600 6978 33652
rect 7650 33600 7656 33652
rect 7708 33640 7714 33652
rect 8113 33643 8171 33649
rect 8113 33640 8125 33643
rect 7708 33612 8125 33640
rect 7708 33600 7714 33612
rect 8113 33609 8125 33612
rect 8159 33609 8171 33643
rect 8294 33640 8300 33652
rect 8113 33603 8171 33609
rect 8266 33600 8300 33640
rect 8352 33600 8358 33652
rect 8662 33600 8668 33652
rect 8720 33640 8726 33652
rect 9306 33640 9312 33652
rect 8720 33612 9312 33640
rect 8720 33600 8726 33612
rect 9306 33600 9312 33612
rect 9364 33600 9370 33652
rect 10686 33640 10692 33652
rect 9793 33612 10692 33640
rect 5491 33544 5948 33572
rect 5997 33575 6055 33581
rect 5491 33541 5503 33544
rect 5445 33535 5503 33541
rect 5997 33541 6009 33575
rect 6043 33541 6055 33575
rect 8266 33572 8294 33600
rect 9214 33572 9220 33584
rect 8266 33544 8432 33572
rect 5997 33535 6055 33541
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33504 1731 33507
rect 1946 33504 1952 33516
rect 1719 33476 1952 33504
rect 1719 33473 1731 33476
rect 1673 33467 1731 33473
rect 1946 33464 1952 33476
rect 2004 33464 2010 33516
rect 2222 33464 2228 33516
rect 2280 33504 2286 33516
rect 2501 33507 2559 33513
rect 2501 33504 2513 33507
rect 2280 33476 2513 33504
rect 2280 33464 2286 33476
rect 2501 33473 2513 33476
rect 2547 33504 2559 33507
rect 4065 33507 4123 33513
rect 4065 33504 4077 33507
rect 2547 33476 4077 33504
rect 2547 33473 2559 33476
rect 2501 33467 2559 33473
rect 4065 33473 4077 33476
rect 4111 33473 4123 33507
rect 4065 33467 4123 33473
rect 5810 33464 5816 33516
rect 5868 33513 5874 33516
rect 5868 33507 5890 33513
rect 5878 33473 5890 33507
rect 5868 33467 5890 33473
rect 5868 33464 5874 33467
rect 1118 33396 1124 33448
rect 1176 33396 1182 33448
rect 1305 33439 1363 33445
rect 1305 33405 1317 33439
rect 1351 33436 1363 33439
rect 1394 33436 1400 33448
rect 1351 33408 1400 33436
rect 1351 33405 1363 33408
rect 1305 33399 1363 33405
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1489 33439 1547 33445
rect 1489 33405 1501 33439
rect 1535 33436 1547 33439
rect 3050 33436 3056 33448
rect 1535 33408 3056 33436
rect 1535 33405 1547 33408
rect 1489 33399 1547 33405
rect 3050 33396 3056 33408
rect 3108 33396 3114 33448
rect 3881 33439 3939 33445
rect 3881 33405 3893 33439
rect 3927 33436 3939 33439
rect 4246 33436 4252 33448
rect 3927 33408 4252 33436
rect 3927 33405 3939 33408
rect 3881 33399 3939 33405
rect 4246 33396 4252 33408
rect 4304 33396 4310 33448
rect 5074 33396 5080 33448
rect 5132 33396 5138 33448
rect 5534 33396 5540 33448
rect 5592 33396 5598 33448
rect 5629 33439 5687 33445
rect 5629 33405 5641 33439
rect 5675 33405 5687 33439
rect 5629 33399 5687 33405
rect 1673 33371 1731 33377
rect 1673 33337 1685 33371
rect 1719 33368 1731 33371
rect 2777 33371 2835 33377
rect 2777 33368 2789 33371
rect 1719 33340 2789 33368
rect 1719 33337 1731 33340
rect 1673 33331 1731 33337
rect 2777 33337 2789 33340
rect 2823 33337 2835 33371
rect 5644 33368 5672 33399
rect 5718 33396 5724 33448
rect 5776 33396 5782 33448
rect 5915 33439 5973 33445
rect 5915 33405 5927 33439
rect 5961 33436 5973 33439
rect 6012 33436 6040 33535
rect 8404 33504 8432 33544
rect 8772 33544 9220 33572
rect 7852 33476 8156 33504
rect 8404 33476 8524 33504
rect 7852 33448 7880 33476
rect 5961 33408 6040 33436
rect 5961 33405 5973 33408
rect 5915 33399 5973 33405
rect 6270 33396 6276 33448
rect 6328 33396 6334 33448
rect 6362 33396 6368 33448
rect 6420 33396 6426 33448
rect 6546 33445 6552 33448
rect 6519 33439 6552 33445
rect 6519 33405 6531 33439
rect 6519 33399 6552 33405
rect 6546 33396 6552 33399
rect 6604 33396 6610 33448
rect 7098 33396 7104 33448
rect 7156 33436 7162 33448
rect 7469 33439 7527 33445
rect 7469 33436 7481 33439
rect 7156 33408 7481 33436
rect 7156 33396 7162 33408
rect 7469 33405 7481 33408
rect 7515 33405 7527 33439
rect 7469 33399 7527 33405
rect 7834 33396 7840 33448
rect 7892 33396 7898 33448
rect 7926 33396 7932 33448
rect 7984 33438 7990 33448
rect 8021 33439 8079 33445
rect 8021 33438 8033 33439
rect 7984 33410 8033 33438
rect 7984 33396 7990 33410
rect 8021 33405 8033 33410
rect 8067 33405 8079 33439
rect 8021 33399 8079 33405
rect 5994 33368 6000 33380
rect 5644 33340 6000 33368
rect 2777 33331 2835 33337
rect 5994 33328 6000 33340
rect 6052 33328 6058 33380
rect 6825 33371 6883 33377
rect 6825 33368 6837 33371
rect 6104 33340 6837 33368
rect 842 33260 848 33312
rect 900 33300 906 33312
rect 937 33303 995 33309
rect 937 33300 949 33303
rect 900 33272 949 33300
rect 900 33260 906 33272
rect 937 33269 949 33272
rect 983 33269 995 33303
rect 937 33263 995 33269
rect 2038 33260 2044 33312
rect 2096 33300 2102 33312
rect 2317 33303 2375 33309
rect 2317 33300 2329 33303
rect 2096 33272 2329 33300
rect 2096 33260 2102 33272
rect 2317 33269 2329 33272
rect 2363 33269 2375 33303
rect 2317 33263 2375 33269
rect 2409 33303 2467 33309
rect 2409 33269 2421 33303
rect 2455 33300 2467 33303
rect 2498 33300 2504 33312
rect 2455 33272 2504 33300
rect 2455 33269 2467 33272
rect 2409 33263 2467 33269
rect 2498 33260 2504 33272
rect 2556 33260 2562 33312
rect 2958 33260 2964 33312
rect 3016 33260 3022 33312
rect 3970 33260 3976 33312
rect 4028 33300 4034 33312
rect 4522 33300 4528 33312
rect 4028 33272 4528 33300
rect 4028 33260 4034 33272
rect 4522 33260 4528 33272
rect 4580 33260 4586 33312
rect 5166 33260 5172 33312
rect 5224 33300 5230 33312
rect 6104 33300 6132 33340
rect 6825 33337 6837 33340
rect 6871 33368 6883 33371
rect 7374 33368 7380 33380
rect 6871 33340 7380 33368
rect 6871 33337 6883 33340
rect 6825 33331 6883 33337
rect 7374 33328 7380 33340
rect 7432 33328 7438 33380
rect 8128 33368 8156 33476
rect 8205 33439 8263 33445
rect 8205 33405 8217 33439
rect 8251 33438 8263 33439
rect 8294 33438 8300 33450
rect 8251 33410 8300 33438
rect 8251 33405 8263 33410
rect 8205 33399 8263 33405
rect 8294 33398 8300 33410
rect 8352 33398 8358 33450
rect 8386 33396 8392 33448
rect 8444 33396 8450 33448
rect 8496 33445 8524 33476
rect 8772 33445 8800 33544
rect 9214 33532 9220 33544
rect 9272 33532 9278 33584
rect 9585 33575 9643 33581
rect 9585 33572 9597 33575
rect 9416 33544 9597 33572
rect 9309 33507 9367 33513
rect 9309 33504 9321 33507
rect 9232 33476 9321 33504
rect 8481 33439 8539 33445
rect 8481 33405 8493 33439
rect 8527 33405 8539 33439
rect 8481 33399 8539 33405
rect 8757 33439 8815 33445
rect 8757 33405 8769 33439
rect 8803 33405 8815 33439
rect 8757 33399 8815 33405
rect 8849 33439 8907 33445
rect 8849 33405 8861 33439
rect 8895 33405 8907 33439
rect 8849 33399 8907 33405
rect 8128 33340 8524 33368
rect 5224 33272 6132 33300
rect 6181 33303 6239 33309
rect 5224 33260 5230 33272
rect 6181 33269 6193 33303
rect 6227 33300 6239 33303
rect 6362 33300 6368 33312
rect 6227 33272 6368 33300
rect 6227 33269 6239 33272
rect 6181 33263 6239 33269
rect 6362 33260 6368 33272
rect 6420 33260 6426 33312
rect 6733 33303 6791 33309
rect 6733 33269 6745 33303
rect 6779 33300 6791 33303
rect 7098 33300 7104 33312
rect 6779 33272 7104 33300
rect 6779 33269 6791 33272
rect 6733 33263 6791 33269
rect 7098 33260 7104 33272
rect 7156 33260 7162 33312
rect 7650 33260 7656 33312
rect 7708 33300 7714 33312
rect 7834 33300 7840 33312
rect 7708 33272 7840 33300
rect 7708 33260 7714 33272
rect 7834 33260 7840 33272
rect 7892 33260 7898 33312
rect 8496 33300 8524 33340
rect 8570 33328 8576 33380
rect 8628 33368 8634 33380
rect 8665 33371 8723 33377
rect 8665 33368 8677 33371
rect 8628 33340 8677 33368
rect 8628 33328 8634 33340
rect 8665 33337 8677 33340
rect 8711 33337 8723 33371
rect 8665 33331 8723 33337
rect 8864 33300 8892 33399
rect 9232 33312 9260 33476
rect 9309 33473 9321 33476
rect 9355 33473 9367 33507
rect 9309 33467 9367 33473
rect 9416 33436 9444 33544
rect 9585 33541 9597 33544
rect 9631 33572 9643 33575
rect 9793 33572 9821 33612
rect 10686 33600 10692 33612
rect 10744 33600 10750 33652
rect 9631 33544 9821 33572
rect 9631 33541 9643 33544
rect 9585 33535 9643 33541
rect 9858 33532 9864 33584
rect 9916 33572 9922 33584
rect 10321 33575 10379 33581
rect 10321 33572 10333 33575
rect 9916 33544 10333 33572
rect 9916 33532 9922 33544
rect 10321 33541 10333 33544
rect 10367 33541 10379 33575
rect 10321 33535 10379 33541
rect 10410 33532 10416 33584
rect 10468 33532 10474 33584
rect 9766 33504 9772 33516
rect 9324 33408 9444 33436
rect 9499 33476 9772 33504
rect 9324 33380 9352 33408
rect 9306 33328 9312 33380
rect 9364 33328 9370 33380
rect 8496 33272 8892 33300
rect 9030 33260 9036 33312
rect 9088 33260 9094 33312
rect 9214 33260 9220 33312
rect 9272 33300 9278 33312
rect 9499 33300 9527 33476
rect 9766 33464 9772 33476
rect 9824 33464 9830 33516
rect 10428 33504 10456 33532
rect 10152 33476 10456 33504
rect 10152 33448 10180 33476
rect 9582 33396 9588 33448
rect 9640 33436 9646 33448
rect 10045 33439 10103 33445
rect 10045 33436 10057 33439
rect 9640 33408 10057 33436
rect 9640 33396 9646 33408
rect 10045 33405 10057 33408
rect 10091 33405 10103 33439
rect 10045 33399 10103 33405
rect 10134 33396 10140 33448
rect 10192 33396 10198 33448
rect 10410 33396 10416 33448
rect 10468 33396 10474 33448
rect 10321 33371 10379 33377
rect 10321 33337 10333 33371
rect 10367 33337 10379 33371
rect 10321 33331 10379 33337
rect 9272 33272 9527 33300
rect 9272 33260 9278 33272
rect 9766 33260 9772 33312
rect 9824 33260 9830 33312
rect 10336 33300 10364 33331
rect 10410 33300 10416 33312
rect 10336 33272 10416 33300
rect 10410 33260 10416 33272
rect 10468 33260 10474 33312
rect 10597 33303 10655 33309
rect 10597 33269 10609 33303
rect 10643 33300 10655 33303
rect 11238 33300 11244 33312
rect 10643 33272 11244 33300
rect 10643 33269 10655 33272
rect 10597 33263 10655 33269
rect 11238 33260 11244 33272
rect 11296 33260 11302 33312
rect 552 33210 11132 33232
rect 552 33158 4322 33210
rect 4374 33158 4386 33210
rect 4438 33158 4450 33210
rect 4502 33158 4514 33210
rect 4566 33158 4578 33210
rect 4630 33158 10722 33210
rect 10774 33158 10786 33210
rect 10838 33158 10850 33210
rect 10902 33158 10914 33210
rect 10966 33158 10978 33210
rect 11030 33158 11132 33210
rect 552 33136 11132 33158
rect 842 33056 848 33108
rect 900 33096 906 33108
rect 2869 33099 2927 33105
rect 2869 33096 2881 33099
rect 900 33068 2881 33096
rect 900 33056 906 33068
rect 2869 33065 2881 33068
rect 2915 33065 2927 33099
rect 2869 33059 2927 33065
rect 4338 33056 4344 33108
rect 4396 33096 4402 33108
rect 6730 33096 6736 33108
rect 4396 33068 6736 33096
rect 4396 33056 4402 33068
rect 937 33031 995 33037
rect 937 32997 949 33031
rect 983 33028 995 33031
rect 3329 33031 3387 33037
rect 3329 33028 3341 33031
rect 983 33000 1808 33028
rect 983 32997 995 33000
rect 937 32991 995 32997
rect 1118 32920 1124 32972
rect 1176 32960 1182 32972
rect 1486 32960 1492 32972
rect 1176 32932 1492 32960
rect 1176 32920 1182 32932
rect 1486 32920 1492 32932
rect 1544 32920 1550 32972
rect 1578 32920 1584 32972
rect 1636 32920 1642 32972
rect 1780 32969 1808 33000
rect 2884 33000 3341 33028
rect 1765 32963 1823 32969
rect 1765 32929 1777 32963
rect 1811 32960 1823 32963
rect 2038 32960 2044 32972
rect 1811 32932 2044 32960
rect 1811 32929 1823 32932
rect 1765 32923 1823 32929
rect 2038 32920 2044 32932
rect 2096 32920 2102 32972
rect 2130 32920 2136 32972
rect 2188 32920 2194 32972
rect 2682 32920 2688 32972
rect 2740 32920 2746 32972
rect 1394 32852 1400 32904
rect 1452 32892 1458 32904
rect 2884 32892 2912 33000
rect 3329 32997 3341 33000
rect 3375 33028 3387 33031
rect 5810 33028 5816 33040
rect 3375 33000 5816 33028
rect 3375 32997 3387 33000
rect 3329 32991 3387 32997
rect 5810 32988 5816 33000
rect 5868 32988 5874 33040
rect 2961 32963 3019 32969
rect 2961 32929 2973 32963
rect 3007 32960 3019 32963
rect 3050 32960 3056 32972
rect 3007 32932 3056 32960
rect 3007 32929 3019 32932
rect 2961 32923 3019 32929
rect 3050 32920 3056 32932
rect 3108 32920 3114 32972
rect 3145 32963 3203 32969
rect 3145 32929 3157 32963
rect 3191 32929 3203 32963
rect 3145 32923 3203 32929
rect 1452 32864 2912 32892
rect 1452 32852 1458 32864
rect 1305 32827 1363 32833
rect 1305 32793 1317 32827
rect 1351 32824 1363 32827
rect 1762 32824 1768 32836
rect 1351 32796 1768 32824
rect 1351 32793 1363 32796
rect 1305 32787 1363 32793
rect 1762 32784 1768 32796
rect 1820 32824 1826 32836
rect 2958 32824 2964 32836
rect 1820 32796 2964 32824
rect 1820 32784 1826 32796
rect 2958 32784 2964 32796
rect 3016 32824 3022 32836
rect 3160 32824 3188 32923
rect 3510 32920 3516 32972
rect 3568 32960 3574 32972
rect 3605 32963 3663 32969
rect 3605 32960 3617 32963
rect 3568 32932 3617 32960
rect 3568 32920 3574 32932
rect 3605 32929 3617 32932
rect 3651 32929 3663 32963
rect 3605 32923 3663 32929
rect 3694 32920 3700 32972
rect 3752 32920 3758 32972
rect 3881 32963 3939 32969
rect 3881 32929 3893 32963
rect 3927 32929 3939 32963
rect 3881 32923 3939 32929
rect 3896 32892 3924 32923
rect 4246 32920 4252 32972
rect 4304 32920 4310 32972
rect 4338 32920 4344 32972
rect 4396 32920 4402 32972
rect 4525 32963 4583 32969
rect 4525 32929 4537 32963
rect 4571 32960 4583 32963
rect 4890 32960 4896 32972
rect 4571 32932 4896 32960
rect 4571 32929 4583 32932
rect 4525 32923 4583 32929
rect 4890 32920 4896 32932
rect 4948 32920 4954 32972
rect 5261 32963 5319 32969
rect 5261 32929 5273 32963
rect 5307 32929 5319 32963
rect 5261 32923 5319 32929
rect 5276 32892 5304 32923
rect 5534 32920 5540 32972
rect 5592 32920 5598 32972
rect 5902 32920 5908 32972
rect 5960 32920 5966 32972
rect 6104 32969 6132 33068
rect 6730 33056 6736 33068
rect 6788 33056 6794 33108
rect 6822 33056 6828 33108
rect 6880 33096 6886 33108
rect 7745 33099 7803 33105
rect 7745 33096 7757 33099
rect 6880 33068 7757 33096
rect 6880 33056 6886 33068
rect 7745 33065 7757 33068
rect 7791 33065 7803 33099
rect 7745 33059 7803 33065
rect 7852 33068 8248 33096
rect 6365 33031 6423 33037
rect 6365 32997 6377 33031
rect 6411 33028 6423 33031
rect 6411 33000 7512 33028
rect 6411 32997 6423 33000
rect 6365 32991 6423 32997
rect 7484 32972 7512 33000
rect 7558 32988 7564 33040
rect 7616 33028 7622 33040
rect 7852 33028 7880 33068
rect 7616 33000 7880 33028
rect 7616 32988 7622 33000
rect 8018 32988 8024 33040
rect 8076 33028 8082 33040
rect 8076 33000 8156 33028
rect 8076 32988 8082 33000
rect 6089 32963 6147 32969
rect 6089 32929 6101 32963
rect 6135 32929 6147 32963
rect 6089 32923 6147 32929
rect 6181 32963 6239 32969
rect 6181 32929 6193 32963
rect 6227 32929 6239 32963
rect 6181 32923 6239 32929
rect 5626 32892 5632 32904
rect 3896 32864 5632 32892
rect 5626 32852 5632 32864
rect 5684 32852 5690 32904
rect 5718 32852 5724 32904
rect 5776 32892 5782 32904
rect 6196 32892 6224 32923
rect 6822 32920 6828 32972
rect 6880 32920 6886 32972
rect 7006 32920 7012 32972
rect 7064 32920 7070 32972
rect 7466 32920 7472 32972
rect 7524 32920 7530 32972
rect 5776 32864 6224 32892
rect 5776 32852 5782 32864
rect 6362 32852 6368 32904
rect 6420 32892 6426 32904
rect 6420 32864 6684 32892
rect 6420 32852 6426 32864
rect 4433 32827 4491 32833
rect 4433 32824 4445 32827
rect 3016 32796 3188 32824
rect 3988 32796 4445 32824
rect 3016 32784 3022 32796
rect 2038 32716 2044 32768
rect 2096 32756 2102 32768
rect 2406 32756 2412 32768
rect 2096 32728 2412 32756
rect 2096 32716 2102 32728
rect 2406 32716 2412 32728
rect 2464 32716 2470 32768
rect 2498 32716 2504 32768
rect 2556 32716 2562 32768
rect 2682 32716 2688 32768
rect 2740 32756 2746 32768
rect 3988 32756 4016 32796
rect 4433 32793 4445 32796
rect 4479 32824 4491 32827
rect 4614 32824 4620 32836
rect 4479 32796 4620 32824
rect 4479 32793 4491 32796
rect 4433 32787 4491 32793
rect 4614 32784 4620 32796
rect 4672 32784 4678 32836
rect 5994 32784 6000 32836
rect 6052 32784 6058 32836
rect 6546 32824 6552 32836
rect 6380 32796 6552 32824
rect 2740 32728 4016 32756
rect 2740 32716 2746 32728
rect 4062 32716 4068 32768
rect 4120 32716 4126 32768
rect 4709 32759 4767 32765
rect 4709 32725 4721 32759
rect 4755 32756 4767 32759
rect 4982 32756 4988 32768
rect 4755 32728 4988 32756
rect 4755 32725 4767 32728
rect 4709 32719 4767 32725
rect 4982 32716 4988 32728
rect 5040 32716 5046 32768
rect 5074 32716 5080 32768
rect 5132 32716 5138 32768
rect 5445 32759 5503 32765
rect 5445 32725 5457 32759
rect 5491 32756 5503 32759
rect 5902 32756 5908 32768
rect 5491 32728 5908 32756
rect 5491 32725 5503 32728
rect 5445 32719 5503 32725
rect 5902 32716 5908 32728
rect 5960 32756 5966 32768
rect 6380 32756 6408 32796
rect 6546 32784 6552 32796
rect 6604 32784 6610 32836
rect 5960 32728 6408 32756
rect 6457 32759 6515 32765
rect 5960 32716 5966 32728
rect 6457 32725 6469 32759
rect 6503 32756 6515 32759
rect 6656 32756 6684 32864
rect 6730 32852 6736 32904
rect 6788 32852 6794 32904
rect 7285 32895 7343 32901
rect 7285 32861 7297 32895
rect 7331 32861 7343 32895
rect 7285 32855 7343 32861
rect 7300 32824 7328 32855
rect 7926 32852 7932 32904
rect 7984 32852 7990 32904
rect 8018 32852 8024 32904
rect 8076 32852 8082 32904
rect 8128 32901 8156 33000
rect 8220 32969 8248 33068
rect 8846 33056 8852 33108
rect 8904 33056 8910 33108
rect 9125 33099 9183 33105
rect 9125 33096 9137 33099
rect 8956 33068 9137 33096
rect 8294 32988 8300 33040
rect 8352 33028 8358 33040
rect 8956 33028 8984 33068
rect 9125 33065 9137 33068
rect 9171 33096 9183 33099
rect 9674 33096 9680 33108
rect 9171 33068 9680 33096
rect 9171 33065 9183 33068
rect 9125 33059 9183 33065
rect 9674 33056 9680 33068
rect 9732 33096 9738 33108
rect 10594 33096 10600 33108
rect 9732 33068 10600 33096
rect 9732 33056 9738 33068
rect 10594 33056 10600 33068
rect 10652 33056 10658 33108
rect 10689 33099 10747 33105
rect 10689 33065 10701 33099
rect 10735 33096 10747 33099
rect 10870 33096 10876 33108
rect 10735 33068 10876 33096
rect 10735 33065 10747 33068
rect 10689 33059 10747 33065
rect 10870 33056 10876 33068
rect 10928 33056 10934 33108
rect 8352 33000 8984 33028
rect 8352 32988 8358 33000
rect 9030 32988 9036 33040
rect 9088 32988 9094 33040
rect 9950 32988 9956 33040
rect 10008 33028 10014 33040
rect 10238 33031 10296 33037
rect 10238 33028 10250 33031
rect 10008 33000 10250 33028
rect 10008 32988 10014 33000
rect 10238 32997 10250 33000
rect 10284 32997 10296 33031
rect 11330 33028 11336 33040
rect 10238 32991 10296 32997
rect 10612 33000 11336 33028
rect 8205 32963 8263 32969
rect 8205 32929 8217 32963
rect 8251 32929 8263 32963
rect 8205 32923 8263 32929
rect 8386 32920 8392 32972
rect 8444 32920 8450 32972
rect 8481 32963 8539 32969
rect 8481 32929 8493 32963
rect 8527 32929 8539 32963
rect 8481 32923 8539 32929
rect 8113 32895 8171 32901
rect 8113 32861 8125 32895
rect 8159 32861 8171 32895
rect 8113 32855 8171 32861
rect 8294 32852 8300 32904
rect 8352 32892 8358 32904
rect 8496 32892 8524 32923
rect 8662 32920 8668 32972
rect 8720 32920 8726 32972
rect 8754 32920 8760 32972
rect 8812 32920 8818 32972
rect 9674 32960 9680 32972
rect 9048 32932 9680 32960
rect 8352 32864 8524 32892
rect 8352 32852 8358 32864
rect 7374 32824 7380 32836
rect 7300 32796 7380 32824
rect 7374 32784 7380 32796
rect 7432 32824 7438 32836
rect 9048 32833 9076 32932
rect 9674 32920 9680 32932
rect 9732 32920 9738 32972
rect 10612 32969 10640 33000
rect 11330 32988 11336 33000
rect 11388 32988 11394 33040
rect 10597 32963 10655 32969
rect 10597 32929 10609 32963
rect 10643 32929 10655 32963
rect 10597 32923 10655 32929
rect 10781 32963 10839 32969
rect 10781 32929 10793 32963
rect 10827 32960 10839 32963
rect 10827 32932 10916 32960
rect 10827 32929 10839 32932
rect 10781 32923 10839 32929
rect 10502 32852 10508 32904
rect 10560 32892 10566 32904
rect 10560 32864 10824 32892
rect 10560 32852 10566 32864
rect 10796 32836 10824 32864
rect 8389 32827 8447 32833
rect 8389 32824 8401 32827
rect 7432 32796 8401 32824
rect 7432 32784 7438 32796
rect 8389 32793 8401 32796
rect 8435 32793 8447 32827
rect 8389 32787 8447 32793
rect 9033 32827 9091 32833
rect 9033 32793 9045 32827
rect 9079 32793 9091 32827
rect 9033 32787 9091 32793
rect 10778 32784 10784 32836
rect 10836 32784 10842 32836
rect 6730 32756 6736 32768
rect 6503 32728 6736 32756
rect 6503 32725 6515 32728
rect 6457 32719 6515 32725
rect 6730 32716 6736 32728
rect 6788 32716 6794 32768
rect 6825 32759 6883 32765
rect 6825 32725 6837 32759
rect 6871 32756 6883 32759
rect 6914 32756 6920 32768
rect 6871 32728 6920 32756
rect 6871 32725 6883 32728
rect 6825 32719 6883 32725
rect 6914 32716 6920 32728
rect 6972 32716 6978 32768
rect 7098 32716 7104 32768
rect 7156 32716 7162 32768
rect 7282 32716 7288 32768
rect 7340 32756 7346 32768
rect 7653 32759 7711 32765
rect 7653 32756 7665 32759
rect 7340 32728 7665 32756
rect 7340 32716 7346 32728
rect 7653 32725 7665 32728
rect 7699 32725 7711 32759
rect 7653 32719 7711 32725
rect 7834 32716 7840 32768
rect 7892 32756 7898 32768
rect 8570 32756 8576 32768
rect 7892 32728 8576 32756
rect 7892 32716 7898 32728
rect 8570 32716 8576 32728
rect 8628 32756 8634 32768
rect 10888 32756 10916 32932
rect 8628 32728 10916 32756
rect 8628 32716 8634 32728
rect 552 32666 11132 32688
rect 552 32614 3662 32666
rect 3714 32614 3726 32666
rect 3778 32614 3790 32666
rect 3842 32614 3854 32666
rect 3906 32614 3918 32666
rect 3970 32614 10062 32666
rect 10114 32614 10126 32666
rect 10178 32614 10190 32666
rect 10242 32614 10254 32666
rect 10306 32614 10318 32666
rect 10370 32614 11132 32666
rect 552 32592 11132 32614
rect 1946 32512 1952 32564
rect 2004 32552 2010 32564
rect 2501 32555 2559 32561
rect 2501 32552 2513 32555
rect 2004 32524 2513 32552
rect 2004 32512 2010 32524
rect 2424 32496 2452 32524
rect 2501 32521 2513 32524
rect 2547 32521 2559 32555
rect 2501 32515 2559 32521
rect 3510 32512 3516 32564
rect 3568 32552 3574 32564
rect 5902 32552 5908 32564
rect 3568 32524 5908 32552
rect 3568 32512 3574 32524
rect 5902 32512 5908 32524
rect 5960 32512 5966 32564
rect 6086 32512 6092 32564
rect 6144 32512 6150 32564
rect 6273 32555 6331 32561
rect 6273 32521 6285 32555
rect 6319 32552 6331 32555
rect 6914 32552 6920 32564
rect 6319 32524 6920 32552
rect 6319 32521 6331 32524
rect 6273 32515 6331 32521
rect 6914 32512 6920 32524
rect 6972 32512 6978 32564
rect 7098 32512 7104 32564
rect 7156 32552 7162 32564
rect 7834 32552 7840 32564
rect 7156 32524 7840 32552
rect 7156 32512 7162 32524
rect 7834 32512 7840 32524
rect 7892 32512 7898 32564
rect 8202 32512 8208 32564
rect 8260 32552 8266 32564
rect 9401 32555 9459 32561
rect 9401 32552 9413 32555
rect 8260 32524 9413 32552
rect 8260 32512 8266 32524
rect 9401 32521 9413 32524
rect 9447 32521 9459 32555
rect 10502 32552 10508 32564
rect 9401 32515 9459 32521
rect 9600 32524 10508 32552
rect 9600 32496 9628 32524
rect 10502 32512 10508 32524
rect 10560 32552 10566 32564
rect 10870 32552 10876 32564
rect 10560 32524 10876 32552
rect 10560 32512 10566 32524
rect 10870 32512 10876 32524
rect 10928 32512 10934 32564
rect 2406 32444 2412 32496
rect 2464 32444 2470 32496
rect 3234 32444 3240 32496
rect 3292 32484 3298 32496
rect 3694 32484 3700 32496
rect 3292 32456 3700 32484
rect 3292 32444 3298 32456
rect 3694 32444 3700 32456
rect 3752 32444 3758 32496
rect 5534 32444 5540 32496
rect 5592 32484 5598 32496
rect 5592 32456 6132 32484
rect 5592 32444 5598 32456
rect 2225 32419 2283 32425
rect 2225 32385 2237 32419
rect 2271 32416 2283 32419
rect 2271 32388 3280 32416
rect 2271 32385 2283 32388
rect 2225 32379 2283 32385
rect 3252 32360 3280 32388
rect 5810 32376 5816 32428
rect 5868 32416 5874 32428
rect 5905 32419 5963 32425
rect 5905 32416 5917 32419
rect 5868 32388 5917 32416
rect 5868 32376 5874 32388
rect 5905 32385 5917 32388
rect 5951 32385 5963 32419
rect 5905 32379 5963 32385
rect 1969 32351 2027 32357
rect 1969 32317 1981 32351
rect 2015 32348 2027 32351
rect 2314 32348 2320 32360
rect 2015 32320 2320 32348
rect 2015 32317 2027 32320
rect 1969 32311 2027 32317
rect 2314 32308 2320 32320
rect 2372 32308 2378 32360
rect 2682 32348 2688 32360
rect 2424 32320 2688 32348
rect 1302 32240 1308 32292
rect 1360 32280 1366 32292
rect 2424 32280 2452 32320
rect 2682 32308 2688 32320
rect 2740 32308 2746 32360
rect 2866 32308 2872 32360
rect 2924 32308 2930 32360
rect 3234 32308 3240 32360
rect 3292 32348 3298 32360
rect 3789 32351 3847 32357
rect 3789 32348 3801 32351
rect 3292 32320 3801 32348
rect 3292 32308 3298 32320
rect 3789 32317 3801 32320
rect 3835 32317 3847 32351
rect 3789 32311 3847 32317
rect 3878 32308 3884 32360
rect 3936 32348 3942 32360
rect 5258 32348 5264 32360
rect 3936 32320 5264 32348
rect 3936 32308 3942 32320
rect 5258 32308 5264 32320
rect 5316 32308 5322 32360
rect 5442 32308 5448 32360
rect 5500 32308 5506 32360
rect 1360 32252 2452 32280
rect 1360 32240 1366 32252
rect 2498 32240 2504 32292
rect 2556 32240 2562 32292
rect 3605 32283 3663 32289
rect 3605 32249 3617 32283
rect 3651 32249 3663 32283
rect 3605 32243 3663 32249
rect 4056 32283 4114 32289
rect 4056 32249 4068 32283
rect 4102 32280 4114 32283
rect 4798 32280 4804 32292
rect 4102 32252 4804 32280
rect 4102 32249 4114 32252
rect 4056 32243 4114 32249
rect 14 32172 20 32224
rect 72 32212 78 32224
rect 845 32215 903 32221
rect 845 32212 857 32215
rect 72 32184 857 32212
rect 72 32172 78 32184
rect 845 32181 857 32184
rect 891 32212 903 32215
rect 1578 32212 1584 32224
rect 891 32184 1584 32212
rect 891 32181 903 32184
rect 845 32175 903 32181
rect 1578 32172 1584 32184
rect 1636 32172 1642 32224
rect 2317 32215 2375 32221
rect 2317 32181 2329 32215
rect 2363 32212 2375 32215
rect 2682 32212 2688 32224
rect 2363 32184 2688 32212
rect 2363 32181 2375 32184
rect 2317 32175 2375 32181
rect 2682 32172 2688 32184
rect 2740 32172 2746 32224
rect 3510 32172 3516 32224
rect 3568 32172 3574 32224
rect 3620 32212 3648 32243
rect 4798 32240 4804 32252
rect 4856 32240 4862 32292
rect 5460 32280 5488 32308
rect 5629 32283 5687 32289
rect 5629 32280 5641 32283
rect 5460 32252 5641 32280
rect 5629 32249 5641 32252
rect 5675 32280 5687 32283
rect 5810 32280 5816 32292
rect 5675 32252 5816 32280
rect 5675 32249 5687 32252
rect 5629 32243 5687 32249
rect 5810 32240 5816 32252
rect 5868 32240 5874 32292
rect 5920 32280 5948 32379
rect 6104 32357 6132 32456
rect 6454 32444 6460 32496
rect 6512 32484 6518 32496
rect 6641 32487 6699 32493
rect 6641 32484 6653 32487
rect 6512 32456 6653 32484
rect 6512 32444 6518 32456
rect 6641 32453 6653 32456
rect 6687 32453 6699 32487
rect 8018 32484 8024 32496
rect 6641 32447 6699 32453
rect 6932 32456 8024 32484
rect 6178 32376 6184 32428
rect 6236 32416 6242 32428
rect 6932 32425 6960 32456
rect 8018 32444 8024 32456
rect 8076 32444 8082 32496
rect 8220 32456 8616 32484
rect 6917 32419 6975 32425
rect 6236 32388 6500 32416
rect 6236 32376 6242 32388
rect 6089 32351 6147 32357
rect 6089 32317 6101 32351
rect 6135 32348 6147 32351
rect 6270 32348 6276 32360
rect 6135 32320 6276 32348
rect 6135 32317 6147 32320
rect 6089 32311 6147 32317
rect 6270 32308 6276 32320
rect 6328 32308 6334 32360
rect 6472 32357 6500 32388
rect 6917 32385 6929 32419
rect 6963 32385 6975 32419
rect 6917 32379 6975 32385
rect 7374 32376 7380 32428
rect 7432 32376 7438 32428
rect 8220 32425 8248 32456
rect 8205 32419 8263 32425
rect 8205 32385 8217 32419
rect 8251 32385 8263 32419
rect 8205 32379 8263 32385
rect 6457 32351 6515 32357
rect 6457 32317 6469 32351
rect 6503 32317 6515 32351
rect 6457 32311 6515 32317
rect 6546 32308 6552 32360
rect 6604 32308 6610 32360
rect 6733 32351 6791 32357
rect 6733 32317 6745 32351
rect 6779 32348 6791 32351
rect 7190 32348 7196 32360
rect 6779 32320 7196 32348
rect 6779 32317 6791 32320
rect 6733 32311 6791 32317
rect 7190 32308 7196 32320
rect 7248 32308 7254 32360
rect 7466 32308 7472 32360
rect 7524 32308 7530 32360
rect 8294 32348 8300 32360
rect 7576 32320 8300 32348
rect 6178 32280 6184 32292
rect 5920 32252 6184 32280
rect 6178 32240 6184 32252
rect 6236 32240 6242 32292
rect 7006 32240 7012 32292
rect 7064 32240 7070 32292
rect 4430 32212 4436 32224
rect 3620 32184 4436 32212
rect 4430 32172 4436 32184
rect 4488 32172 4494 32224
rect 5169 32215 5227 32221
rect 5169 32181 5181 32215
rect 5215 32212 5227 32215
rect 5350 32212 5356 32224
rect 5215 32184 5356 32212
rect 5215 32181 5227 32184
rect 5169 32175 5227 32181
rect 5350 32172 5356 32184
rect 5408 32172 5414 32224
rect 5445 32215 5503 32221
rect 5445 32181 5457 32215
rect 5491 32212 5503 32215
rect 5534 32212 5540 32224
rect 5491 32184 5540 32212
rect 5491 32181 5503 32184
rect 5445 32175 5503 32181
rect 5534 32172 5540 32184
rect 5592 32212 5598 32224
rect 7576 32212 7604 32320
rect 8294 32308 8300 32320
rect 8352 32308 8358 32360
rect 8588 32357 8616 32456
rect 8662 32444 8668 32496
rect 8720 32484 8726 32496
rect 8757 32487 8815 32493
rect 8757 32484 8769 32487
rect 8720 32456 8769 32484
rect 8720 32444 8726 32456
rect 8757 32453 8769 32456
rect 8803 32453 8815 32487
rect 8757 32447 8815 32453
rect 9030 32444 9036 32496
rect 9088 32484 9094 32496
rect 9582 32484 9588 32496
rect 9088 32456 9588 32484
rect 9088 32444 9094 32456
rect 9582 32444 9588 32456
rect 9640 32444 9646 32496
rect 9490 32416 9496 32428
rect 8956 32388 9496 32416
rect 8956 32360 8984 32388
rect 9490 32376 9496 32388
rect 9548 32376 9554 32428
rect 10778 32376 10784 32428
rect 10836 32376 10842 32428
rect 8481 32351 8539 32357
rect 8481 32317 8493 32351
rect 8527 32317 8539 32351
rect 8481 32311 8539 32317
rect 8573 32351 8631 32357
rect 8573 32317 8585 32351
rect 8619 32348 8631 32351
rect 8662 32348 8668 32360
rect 8619 32320 8668 32348
rect 8619 32317 8631 32320
rect 8573 32311 8631 32317
rect 8021 32283 8079 32289
rect 8021 32249 8033 32283
rect 8067 32280 8079 32283
rect 8202 32280 8208 32292
rect 8067 32252 8208 32280
rect 8067 32249 8079 32252
rect 8021 32243 8079 32249
rect 8202 32240 8208 32252
rect 8260 32240 8266 32292
rect 8386 32240 8392 32292
rect 8444 32280 8450 32292
rect 8496 32280 8524 32311
rect 8662 32308 8668 32320
rect 8720 32308 8726 32360
rect 8938 32308 8944 32360
rect 8996 32308 9002 32360
rect 9033 32351 9091 32357
rect 9033 32317 9045 32351
rect 9079 32317 9091 32351
rect 9033 32311 9091 32317
rect 9217 32351 9275 32357
rect 9217 32317 9229 32351
rect 9263 32348 9275 32351
rect 9306 32348 9312 32360
rect 9263 32320 9312 32348
rect 9263 32317 9275 32320
rect 9217 32311 9275 32317
rect 8846 32280 8852 32292
rect 8444 32252 8852 32280
rect 8444 32240 8450 32252
rect 8846 32240 8852 32252
rect 8904 32240 8910 32292
rect 9048 32280 9076 32311
rect 9306 32308 9312 32320
rect 9364 32308 9370 32360
rect 9582 32308 9588 32360
rect 9640 32348 9646 32360
rect 10796 32348 10824 32376
rect 9640 32320 10824 32348
rect 9640 32308 9646 32320
rect 9122 32280 9128 32292
rect 9048 32252 9128 32280
rect 5592 32184 7604 32212
rect 7653 32215 7711 32221
rect 5592 32172 5598 32184
rect 7653 32181 7665 32215
rect 7699 32212 7711 32215
rect 7926 32212 7932 32224
rect 7699 32184 7932 32212
rect 7699 32181 7711 32184
rect 7653 32175 7711 32181
rect 7926 32172 7932 32184
rect 7984 32212 7990 32224
rect 9048 32212 9076 32252
rect 9122 32240 9128 32252
rect 9180 32240 9186 32292
rect 9766 32240 9772 32292
rect 9824 32280 9830 32292
rect 10514 32283 10572 32289
rect 10514 32280 10526 32283
rect 9824 32252 10526 32280
rect 9824 32240 9830 32252
rect 10514 32249 10526 32252
rect 10560 32249 10572 32283
rect 10514 32243 10572 32249
rect 7984 32184 9076 32212
rect 7984 32172 7990 32184
rect 552 32122 11132 32144
rect 552 32070 4322 32122
rect 4374 32070 4386 32122
rect 4438 32070 4450 32122
rect 4502 32070 4514 32122
rect 4566 32070 4578 32122
rect 4630 32070 10722 32122
rect 10774 32070 10786 32122
rect 10838 32070 10850 32122
rect 10902 32070 10914 32122
rect 10966 32070 10978 32122
rect 11030 32070 11132 32122
rect 552 32048 11132 32070
rect 382 31968 388 32020
rect 440 32008 446 32020
rect 440 31980 3372 32008
rect 440 31968 446 31980
rect 1394 31940 1400 31952
rect 952 31912 1400 31940
rect 952 31881 980 31912
rect 1394 31900 1400 31912
rect 1452 31940 1458 31952
rect 3234 31940 3240 31952
rect 1452 31912 3240 31940
rect 1452 31900 1458 31912
rect 937 31875 995 31881
rect 937 31841 949 31875
rect 983 31841 995 31875
rect 937 31835 995 31841
rect 1026 31832 1032 31884
rect 1084 31872 1090 31884
rect 1193 31875 1251 31881
rect 1193 31872 1205 31875
rect 1084 31844 1205 31872
rect 1084 31832 1090 31844
rect 1193 31841 1205 31844
rect 1239 31841 1251 31875
rect 1193 31835 1251 31841
rect 1946 31832 1952 31884
rect 2004 31872 2010 31884
rect 2222 31872 2228 31884
rect 2004 31844 2228 31872
rect 2004 31832 2010 31844
rect 2222 31832 2228 31844
rect 2280 31832 2286 31884
rect 2424 31881 2452 31912
rect 3234 31900 3240 31912
rect 3292 31900 3298 31952
rect 3344 31940 3372 31980
rect 3786 31968 3792 32020
rect 3844 31968 3850 32020
rect 4706 31968 4712 32020
rect 4764 32008 4770 32020
rect 5534 32008 5540 32020
rect 4764 31980 5540 32008
rect 4764 31968 4770 31980
rect 3881 31943 3939 31949
rect 3881 31940 3893 31943
rect 3344 31912 3893 31940
rect 3881 31909 3893 31912
rect 3927 31909 3939 31943
rect 3881 31903 3939 31909
rect 2682 31881 2688 31884
rect 2409 31875 2467 31881
rect 2409 31841 2421 31875
rect 2455 31841 2467 31875
rect 2676 31872 2688 31881
rect 2643 31844 2688 31872
rect 2409 31835 2467 31841
rect 2676 31835 2688 31844
rect 2682 31832 2688 31835
rect 2740 31832 2746 31884
rect 4430 31832 4436 31884
rect 4488 31832 4494 31884
rect 4932 31881 4960 31980
rect 5534 31968 5540 31980
rect 5592 31968 5598 32020
rect 5629 32011 5687 32017
rect 5629 31977 5641 32011
rect 5675 32008 5687 32011
rect 6181 32011 6239 32017
rect 5675 31980 6132 32008
rect 5675 31977 5687 31980
rect 5629 31971 5687 31977
rect 6104 31952 6132 31980
rect 6181 31977 6193 32011
rect 6227 31977 6239 32011
rect 6181 31971 6239 31977
rect 5718 31940 5724 31952
rect 5368 31912 5724 31940
rect 4893 31875 4960 31881
rect 4893 31841 4905 31875
rect 4939 31844 4960 31875
rect 5261 31875 5319 31881
rect 4939 31841 4951 31844
rect 4893 31835 4951 31841
rect 5261 31841 5273 31875
rect 5307 31872 5319 31875
rect 5368 31872 5396 31912
rect 5718 31900 5724 31912
rect 5776 31900 5782 31952
rect 5810 31900 5816 31952
rect 5868 31900 5874 31952
rect 6086 31900 6092 31952
rect 6144 31900 6150 31952
rect 5307 31844 5396 31872
rect 5997 31875 6055 31881
rect 5307 31841 5319 31844
rect 5261 31835 5319 31841
rect 5997 31841 6009 31875
rect 6043 31841 6055 31875
rect 5997 31835 6055 31841
rect 2130 31764 2136 31816
rect 2188 31804 2194 31816
rect 5169 31807 5227 31813
rect 2188 31776 2360 31804
rect 2188 31764 2194 31776
rect 2332 31745 2360 31776
rect 5169 31773 5181 31807
rect 5215 31804 5227 31807
rect 5353 31807 5411 31813
rect 5215 31776 5304 31804
rect 5215 31773 5227 31776
rect 5169 31767 5227 31773
rect 5276 31748 5304 31776
rect 5353 31773 5365 31807
rect 5399 31773 5411 31807
rect 5353 31767 5411 31773
rect 5445 31807 5503 31813
rect 5445 31773 5457 31807
rect 5491 31804 5503 31807
rect 5810 31804 5816 31816
rect 5491 31776 5816 31804
rect 5491 31773 5503 31776
rect 5445 31767 5503 31773
rect 2317 31739 2375 31745
rect 2317 31705 2329 31739
rect 2363 31736 2375 31739
rect 2363 31708 2397 31736
rect 4724 31708 5212 31736
rect 2363 31705 2375 31708
rect 2317 31699 2375 31705
rect 934 31628 940 31680
rect 992 31668 998 31680
rect 2406 31668 2412 31680
rect 992 31640 2412 31668
rect 992 31628 998 31640
rect 2406 31628 2412 31640
rect 2464 31628 2470 31680
rect 3694 31628 3700 31680
rect 3752 31668 3758 31680
rect 4724 31668 4752 31708
rect 5184 31680 5212 31708
rect 5258 31696 5264 31748
rect 5316 31696 5322 31748
rect 5368 31736 5396 31767
rect 5810 31764 5816 31776
rect 5868 31764 5874 31816
rect 5534 31736 5540 31748
rect 5368 31708 5540 31736
rect 5534 31696 5540 31708
rect 5592 31736 5598 31748
rect 6012 31736 6040 31835
rect 6086 31764 6092 31816
rect 6144 31804 6150 31816
rect 6196 31804 6224 31971
rect 6822 31968 6828 32020
rect 6880 32008 6886 32020
rect 7009 32011 7067 32017
rect 7009 32008 7021 32011
rect 6880 31980 7021 32008
rect 6880 31968 6886 31980
rect 7009 31977 7021 31980
rect 7055 31977 7067 32011
rect 7009 31971 7067 31977
rect 7101 32011 7159 32017
rect 7101 31977 7113 32011
rect 7147 32008 7159 32011
rect 7558 32008 7564 32020
rect 7147 31980 7564 32008
rect 7147 31977 7159 31980
rect 7101 31971 7159 31977
rect 7558 31968 7564 31980
rect 7616 31968 7622 32020
rect 7834 31968 7840 32020
rect 7892 32008 7898 32020
rect 8205 32011 8263 32017
rect 7892 31980 8064 32008
rect 7892 31968 7898 31980
rect 6730 31900 6736 31952
rect 6788 31940 6794 31952
rect 8036 31940 8064 31980
rect 8205 31977 8217 32011
rect 8251 32008 8263 32011
rect 8294 32008 8300 32020
rect 8251 31980 8300 32008
rect 8251 31977 8263 31980
rect 8205 31971 8263 31977
rect 8294 31968 8300 31980
rect 8352 31968 8358 32020
rect 9306 31968 9312 32020
rect 9364 32008 9370 32020
rect 10134 32008 10140 32020
rect 9364 31980 10140 32008
rect 9364 31968 9370 31980
rect 10134 31968 10140 31980
rect 10192 31968 10198 32020
rect 10410 31968 10416 32020
rect 10468 32008 10474 32020
rect 10689 32011 10747 32017
rect 10689 32008 10701 32011
rect 10468 31980 10701 32008
rect 10468 31968 10474 31980
rect 10689 31977 10701 31980
rect 10735 31977 10747 32011
rect 10689 31971 10747 31977
rect 6788 31912 6960 31940
rect 6788 31900 6794 31912
rect 6457 31875 6515 31881
rect 6457 31841 6469 31875
rect 6503 31872 6515 31875
rect 6503 31844 6776 31872
rect 6503 31841 6515 31844
rect 6457 31835 6515 31841
rect 6748 31816 6776 31844
rect 6822 31832 6828 31884
rect 6880 31832 6886 31884
rect 6932 31872 6960 31912
rect 7944 31912 8064 31940
rect 7285 31875 7343 31881
rect 7285 31872 7297 31875
rect 6932 31844 7297 31872
rect 7285 31841 7297 31844
rect 7331 31841 7343 31875
rect 7285 31835 7343 31841
rect 7374 31832 7380 31884
rect 7432 31832 7438 31884
rect 7469 31875 7527 31881
rect 7469 31841 7481 31875
rect 7515 31841 7527 31875
rect 7469 31835 7527 31841
rect 6144 31776 6224 31804
rect 6144 31764 6150 31776
rect 6362 31764 6368 31816
rect 6420 31764 6426 31816
rect 6730 31764 6736 31816
rect 6788 31764 6794 31816
rect 7098 31764 7104 31816
rect 7156 31804 7162 31816
rect 7484 31804 7512 31835
rect 7558 31832 7564 31884
rect 7616 31872 7622 31884
rect 7944 31881 7972 31912
rect 8938 31900 8944 31952
rect 8996 31900 9002 31952
rect 9490 31900 9496 31952
rect 9548 31900 9554 31952
rect 9950 31900 9956 31952
rect 10008 31940 10014 31952
rect 10008 31912 10456 31940
rect 10008 31900 10014 31912
rect 7745 31875 7803 31881
rect 7616 31870 7696 31872
rect 7745 31870 7757 31875
rect 7616 31844 7757 31870
rect 7616 31832 7622 31844
rect 7668 31842 7757 31844
rect 7745 31841 7757 31842
rect 7791 31841 7803 31875
rect 7745 31835 7803 31841
rect 7929 31875 7987 31881
rect 7929 31841 7941 31875
rect 7975 31841 7987 31875
rect 7929 31835 7987 31841
rect 8021 31878 8079 31881
rect 8021 31875 8248 31878
rect 8021 31841 8033 31875
rect 8067 31850 8248 31875
rect 8067 31841 8079 31850
rect 8021 31835 8079 31841
rect 8220 31804 8248 31850
rect 8481 31875 8539 31881
rect 8481 31841 8493 31875
rect 8527 31872 8539 31875
rect 9030 31872 9036 31884
rect 8527 31844 9036 31872
rect 8527 31841 8539 31844
rect 8481 31835 8539 31841
rect 9030 31832 9036 31844
rect 9088 31832 9094 31884
rect 9122 31832 9128 31884
rect 9180 31832 9186 31884
rect 10428 31881 10456 31912
rect 10229 31875 10287 31881
rect 10229 31872 10241 31875
rect 9416 31870 9812 31872
rect 9876 31870 10241 31872
rect 9416 31844 10241 31870
rect 8846 31804 8852 31816
rect 7156 31776 7512 31804
rect 7576 31776 8248 31804
rect 8680 31776 8852 31804
rect 7156 31764 7162 31776
rect 6178 31736 6184 31748
rect 5592 31708 5875 31736
rect 6012 31708 6184 31736
rect 5592 31696 5598 31708
rect 3752 31640 4752 31668
rect 3752 31628 3758 31640
rect 5166 31628 5172 31680
rect 5224 31628 5230 31680
rect 5847 31668 5875 31708
rect 6178 31696 6184 31708
rect 6236 31696 6242 31748
rect 7116 31736 7144 31764
rect 6288 31708 7144 31736
rect 6288 31668 6316 31708
rect 7190 31696 7196 31748
rect 7248 31736 7254 31748
rect 7576 31736 7604 31776
rect 7248 31708 7604 31736
rect 7653 31739 7711 31745
rect 7248 31696 7254 31708
rect 7653 31705 7665 31739
rect 7699 31736 7711 31739
rect 8680 31736 8708 31776
rect 8846 31764 8852 31776
rect 8904 31764 8910 31816
rect 7699 31708 8708 31736
rect 8757 31739 8815 31745
rect 7699 31705 7711 31708
rect 7653 31699 7711 31705
rect 8757 31705 8769 31739
rect 8803 31736 8815 31739
rect 9122 31736 9128 31748
rect 8803 31708 9128 31736
rect 8803 31705 8815 31708
rect 8757 31699 8815 31705
rect 9122 31696 9128 31708
rect 9180 31736 9186 31748
rect 9416 31736 9444 31844
rect 9784 31842 9904 31844
rect 10229 31841 10241 31844
rect 10275 31841 10287 31875
rect 10229 31835 10287 31841
rect 10413 31875 10471 31881
rect 10413 31841 10425 31875
rect 10459 31841 10471 31875
rect 10413 31835 10471 31841
rect 10502 31832 10508 31884
rect 10560 31832 10566 31884
rect 9490 31764 9496 31816
rect 9548 31804 9554 31816
rect 9548 31776 9904 31804
rect 9548 31764 9554 31776
rect 9769 31739 9827 31745
rect 9769 31736 9781 31739
rect 9180 31708 9444 31736
rect 9508 31708 9781 31736
rect 9180 31696 9186 31708
rect 5847 31640 6316 31668
rect 6730 31628 6736 31680
rect 6788 31628 6794 31680
rect 6914 31628 6920 31680
rect 6972 31668 6978 31680
rect 7558 31668 7564 31680
rect 6972 31640 7564 31668
rect 6972 31628 6978 31640
rect 7558 31628 7564 31640
rect 7616 31628 7622 31680
rect 8021 31671 8079 31677
rect 8021 31637 8033 31671
rect 8067 31668 8079 31671
rect 8202 31668 8208 31680
rect 8067 31640 8208 31668
rect 8067 31637 8079 31640
rect 8021 31631 8079 31637
rect 8202 31628 8208 31640
rect 8260 31628 8266 31680
rect 8389 31671 8447 31677
rect 8389 31637 8401 31671
rect 8435 31668 8447 31671
rect 8662 31668 8668 31680
rect 8435 31640 8668 31668
rect 8435 31637 8447 31640
rect 8389 31631 8447 31637
rect 8662 31628 8668 31640
rect 8720 31628 8726 31680
rect 9508 31677 9536 31708
rect 9769 31705 9781 31708
rect 9815 31705 9827 31739
rect 9876 31736 9904 31776
rect 9950 31764 9956 31816
rect 10008 31764 10014 31816
rect 10042 31764 10048 31816
rect 10100 31764 10106 31816
rect 10134 31764 10140 31816
rect 10192 31764 10198 31816
rect 10689 31807 10747 31813
rect 10689 31804 10701 31807
rect 10667 31776 10701 31804
rect 10689 31773 10701 31776
rect 10735 31773 10747 31807
rect 10689 31767 10747 31773
rect 10704 31736 10732 31767
rect 9876 31708 10732 31736
rect 9769 31699 9827 31705
rect 9493 31671 9551 31677
rect 9493 31637 9505 31671
rect 9539 31637 9551 31671
rect 9493 31631 9551 31637
rect 9674 31628 9680 31680
rect 9732 31628 9738 31680
rect 552 31578 11132 31600
rect 552 31526 3662 31578
rect 3714 31526 3726 31578
rect 3778 31526 3790 31578
rect 3842 31526 3854 31578
rect 3906 31526 3918 31578
rect 3970 31526 10062 31578
rect 10114 31526 10126 31578
rect 10178 31526 10190 31578
rect 10242 31526 10254 31578
rect 10306 31526 10318 31578
rect 10370 31526 11132 31578
rect 552 31504 11132 31526
rect 842 31424 848 31476
rect 900 31464 906 31476
rect 1121 31467 1179 31473
rect 1121 31464 1133 31467
rect 900 31436 1133 31464
rect 900 31424 906 31436
rect 1121 31433 1133 31436
rect 1167 31433 1179 31467
rect 1121 31427 1179 31433
rect 1305 31467 1363 31473
rect 1305 31433 1317 31467
rect 1351 31464 1363 31467
rect 2866 31464 2872 31476
rect 1351 31436 2872 31464
rect 1351 31433 1363 31436
rect 1305 31427 1363 31433
rect 2866 31424 2872 31436
rect 2924 31424 2930 31476
rect 3142 31424 3148 31476
rect 3200 31464 3206 31476
rect 4801 31467 4859 31473
rect 4801 31464 4813 31467
rect 3200 31436 4813 31464
rect 3200 31424 3206 31436
rect 4801 31433 4813 31436
rect 4847 31433 4859 31467
rect 4801 31427 4859 31433
rect 5626 31424 5632 31476
rect 5684 31424 5690 31476
rect 5902 31424 5908 31476
rect 5960 31464 5966 31476
rect 5997 31467 6055 31473
rect 5997 31464 6009 31467
rect 5960 31436 6009 31464
rect 5960 31424 5966 31436
rect 5997 31433 6009 31436
rect 6043 31433 6055 31467
rect 5997 31427 6055 31433
rect 6546 31424 6552 31476
rect 6604 31424 6610 31476
rect 6917 31467 6975 31473
rect 6917 31433 6929 31467
rect 6963 31433 6975 31467
rect 6917 31427 6975 31433
rect 7101 31467 7159 31473
rect 7101 31433 7113 31467
rect 7147 31464 7159 31467
rect 7374 31464 7380 31476
rect 7147 31436 7380 31464
rect 7147 31433 7159 31436
rect 7101 31427 7159 31433
rect 2774 31396 2780 31408
rect 1780 31368 2780 31396
rect 1780 31328 1808 31368
rect 2774 31356 2780 31368
rect 2832 31356 2838 31408
rect 1504 31300 1808 31328
rect 1302 31260 1308 31272
rect 952 31232 1308 31260
rect 952 31201 980 31232
rect 1302 31220 1308 31232
rect 1360 31220 1366 31272
rect 937 31195 995 31201
rect 937 31161 949 31195
rect 983 31161 995 31195
rect 937 31155 995 31161
rect 1153 31195 1211 31201
rect 1153 31161 1165 31195
rect 1199 31192 1211 31195
rect 1504 31192 1532 31300
rect 1578 31220 1584 31272
rect 1636 31220 1642 31272
rect 1780 31257 1808 31300
rect 1946 31288 1952 31340
rect 2004 31328 2010 31340
rect 2884 31328 2912 31424
rect 4246 31356 4252 31408
rect 4304 31396 4310 31408
rect 4617 31399 4675 31405
rect 4617 31396 4629 31399
rect 4304 31368 4629 31396
rect 4304 31356 4310 31368
rect 4617 31365 4629 31368
rect 4663 31365 4675 31399
rect 4617 31359 4675 31365
rect 4890 31356 4896 31408
rect 4948 31396 4954 31408
rect 5644 31396 5672 31424
rect 6362 31396 6368 31408
rect 4948 31368 6368 31396
rect 4948 31356 4954 31368
rect 6362 31356 6368 31368
rect 6420 31396 6426 31408
rect 6730 31396 6736 31408
rect 6420 31368 6736 31396
rect 6420 31356 6426 31368
rect 6730 31356 6736 31368
rect 6788 31356 6794 31408
rect 6932 31396 6960 31427
rect 7374 31424 7380 31436
rect 7432 31424 7438 31476
rect 7558 31424 7564 31476
rect 7616 31464 7622 31476
rect 8386 31464 8392 31476
rect 7616 31436 8392 31464
rect 7616 31424 7622 31436
rect 8386 31424 8392 31436
rect 8444 31424 8450 31476
rect 8757 31467 8815 31473
rect 8757 31433 8769 31467
rect 8803 31464 8815 31467
rect 9398 31464 9404 31476
rect 8803 31436 9404 31464
rect 8803 31433 8815 31436
rect 8757 31427 8815 31433
rect 9398 31424 9404 31436
rect 9456 31424 9462 31476
rect 7834 31396 7840 31408
rect 6932 31368 7840 31396
rect 7834 31356 7840 31368
rect 7892 31396 7898 31408
rect 8570 31396 8576 31408
rect 7892 31368 8576 31396
rect 7892 31356 7898 31368
rect 8570 31356 8576 31368
rect 8628 31356 8634 31408
rect 3050 31328 3056 31340
rect 2004 31300 2452 31328
rect 2004 31288 2010 31300
rect 1857 31263 1915 31269
rect 1857 31257 1869 31263
rect 1780 31229 1869 31257
rect 1903 31229 1915 31263
rect 1857 31223 1915 31229
rect 2133 31263 2191 31269
rect 2133 31229 2145 31263
rect 2179 31260 2191 31263
rect 2222 31260 2228 31272
rect 2179 31232 2228 31260
rect 2179 31229 2191 31232
rect 2133 31223 2191 31229
rect 2222 31220 2228 31232
rect 2280 31220 2286 31272
rect 2424 31269 2452 31300
rect 2700 31300 3056 31328
rect 2700 31269 2728 31300
rect 3050 31288 3056 31300
rect 3108 31288 3114 31340
rect 5258 31288 5264 31340
rect 5316 31288 5322 31340
rect 5353 31331 5411 31337
rect 5353 31297 5365 31331
rect 5399 31328 5411 31331
rect 5534 31328 5540 31340
rect 5399 31300 5540 31328
rect 5399 31297 5411 31300
rect 5353 31291 5411 31297
rect 5534 31288 5540 31300
rect 5592 31288 5598 31340
rect 6454 31288 6460 31340
rect 6512 31328 6518 31340
rect 6825 31331 6883 31337
rect 6825 31328 6837 31331
rect 6512 31300 6837 31328
rect 6512 31288 6518 31300
rect 6825 31297 6837 31300
rect 6871 31328 6883 31331
rect 6871 31300 7052 31328
rect 6871 31297 6883 31300
rect 6825 31291 6883 31297
rect 2409 31263 2467 31269
rect 2409 31229 2421 31263
rect 2455 31229 2467 31263
rect 2409 31223 2467 31229
rect 2593 31263 2651 31269
rect 2593 31229 2605 31263
rect 2639 31229 2651 31263
rect 2593 31223 2651 31229
rect 2685 31263 2743 31269
rect 2685 31229 2697 31263
rect 2731 31229 2743 31263
rect 2685 31223 2743 31229
rect 2777 31263 2835 31269
rect 2777 31229 2789 31263
rect 2823 31260 2835 31263
rect 2823 31232 3004 31260
rect 2823 31229 2835 31232
rect 2777 31223 2835 31229
rect 1199 31164 1532 31192
rect 1199 31161 1211 31164
rect 1153 31155 1211 31161
rect 2314 31152 2320 31204
rect 2372 31152 2378 31204
rect 1394 31084 1400 31136
rect 1452 31084 1458 31136
rect 1762 31084 1768 31136
rect 1820 31084 1826 31136
rect 1949 31127 2007 31133
rect 1949 31093 1961 31127
rect 1995 31124 2007 31127
rect 2038 31124 2044 31136
rect 1995 31096 2044 31124
rect 1995 31093 2007 31096
rect 1949 31087 2007 31093
rect 2038 31084 2044 31096
rect 2096 31084 2102 31136
rect 2424 31124 2452 31223
rect 2608 31192 2636 31223
rect 2866 31192 2872 31204
rect 2608 31164 2872 31192
rect 2866 31152 2872 31164
rect 2924 31152 2930 31204
rect 2590 31124 2596 31136
rect 2424 31096 2596 31124
rect 2590 31084 2596 31096
rect 2648 31084 2654 31136
rect 2976 31124 3004 31232
rect 3234 31220 3240 31272
rect 3292 31260 3298 31272
rect 4062 31260 4068 31272
rect 3292 31232 4068 31260
rect 3292 31220 3298 31232
rect 4062 31220 4068 31232
rect 4120 31220 4126 31272
rect 4982 31220 4988 31272
rect 5040 31220 5046 31272
rect 5077 31263 5135 31269
rect 5077 31229 5089 31263
rect 5123 31260 5135 31263
rect 6086 31260 6092 31272
rect 5123 31259 5764 31260
rect 5828 31259 6092 31260
rect 5123 31232 6092 31259
rect 5123 31229 5135 31232
rect 5736 31231 5856 31232
rect 5077 31223 5135 31229
rect 6086 31220 6092 31232
rect 6144 31220 6150 31272
rect 6178 31220 6184 31272
rect 6236 31220 6242 31272
rect 6270 31220 6276 31272
rect 6328 31260 6334 31272
rect 6365 31263 6423 31269
rect 6365 31260 6377 31263
rect 6328 31232 6377 31260
rect 6328 31220 6334 31232
rect 6365 31229 6377 31232
rect 6411 31229 6423 31263
rect 6365 31223 6423 31229
rect 6638 31220 6644 31272
rect 6696 31220 6702 31272
rect 6917 31263 6975 31269
rect 6917 31229 6929 31263
rect 6963 31229 6975 31263
rect 7024 31260 7052 31300
rect 7650 31288 7656 31340
rect 7708 31328 7714 31340
rect 7708 31300 8708 31328
rect 7708 31288 7714 31300
rect 7837 31263 7895 31269
rect 7024 31232 7788 31260
rect 6917 31223 6975 31229
rect 3053 31195 3111 31201
rect 3053 31161 3065 31195
rect 3099 31192 3111 31195
rect 3482 31195 3540 31201
rect 3482 31192 3494 31195
rect 3099 31164 3494 31192
rect 3099 31161 3111 31164
rect 3053 31155 3111 31161
rect 3482 31161 3494 31164
rect 3528 31161 3540 31195
rect 3482 31155 3540 31161
rect 5350 31152 5356 31204
rect 5408 31192 5414 31204
rect 5445 31195 5503 31201
rect 5445 31192 5457 31195
rect 5408 31164 5457 31192
rect 5408 31152 5414 31164
rect 5445 31161 5457 31164
rect 5491 31161 5503 31195
rect 5445 31155 5503 31161
rect 5534 31152 5540 31204
rect 5592 31192 5598 31204
rect 5721 31195 5779 31201
rect 5721 31192 5733 31195
rect 5592 31164 5733 31192
rect 5592 31152 5598 31164
rect 5721 31161 5733 31164
rect 5767 31161 5779 31195
rect 5721 31155 5779 31161
rect 3234 31124 3240 31136
rect 2976 31096 3240 31124
rect 3234 31084 3240 31096
rect 3292 31124 3298 31136
rect 4246 31124 4252 31136
rect 3292 31096 4252 31124
rect 3292 31084 3298 31096
rect 4246 31084 4252 31096
rect 4304 31084 4310 31136
rect 4614 31084 4620 31136
rect 4672 31124 4678 31136
rect 5626 31124 5632 31136
rect 4672 31096 5632 31124
rect 4672 31084 4678 31096
rect 5626 31084 5632 31096
rect 5684 31084 5690 31136
rect 5736 31124 5764 31155
rect 5902 31152 5908 31204
rect 5960 31152 5966 31204
rect 6454 31152 6460 31204
rect 6512 31192 6518 31204
rect 6932 31192 6960 31223
rect 6512 31164 6960 31192
rect 7285 31195 7343 31201
rect 6512 31152 6518 31164
rect 7285 31161 7297 31195
rect 7331 31161 7343 31195
rect 7285 31155 7343 31161
rect 7300 31124 7328 31155
rect 5736 31096 7328 31124
rect 7374 31084 7380 31136
rect 7432 31084 7438 31136
rect 7760 31124 7788 31232
rect 7837 31229 7849 31263
rect 7883 31260 7895 31263
rect 8110 31260 8116 31272
rect 7883 31232 8116 31260
rect 7883 31229 7895 31232
rect 7837 31223 7895 31229
rect 8110 31220 8116 31232
rect 8168 31220 8174 31272
rect 8021 31195 8079 31201
rect 8021 31161 8033 31195
rect 8067 31192 8079 31195
rect 8386 31192 8392 31204
rect 8067 31164 8392 31192
rect 8067 31161 8079 31164
rect 8021 31155 8079 31161
rect 8386 31152 8392 31164
rect 8444 31152 8450 31204
rect 8570 31152 8576 31204
rect 8628 31152 8634 31204
rect 8680 31192 8708 31300
rect 9858 31220 9864 31272
rect 9916 31269 9922 31272
rect 9916 31223 9928 31269
rect 10137 31263 10195 31269
rect 10137 31229 10149 31263
rect 10183 31260 10195 31263
rect 10502 31260 10508 31272
rect 10183 31232 10508 31260
rect 10183 31229 10195 31232
rect 10137 31223 10195 31229
rect 9916 31220 9922 31223
rect 10502 31220 10508 31232
rect 10560 31220 10566 31272
rect 10321 31195 10379 31201
rect 10321 31192 10333 31195
rect 8680 31164 10333 31192
rect 10321 31161 10333 31164
rect 10367 31192 10379 31195
rect 10594 31192 10600 31204
rect 10367 31164 10600 31192
rect 10367 31161 10379 31164
rect 10321 31155 10379 31161
rect 10594 31152 10600 31164
rect 10652 31152 10658 31204
rect 8202 31124 8208 31136
rect 7760 31096 8208 31124
rect 8202 31084 8208 31096
rect 8260 31084 8266 31136
rect 8294 31084 8300 31136
rect 8352 31124 8358 31136
rect 8481 31127 8539 31133
rect 8481 31124 8493 31127
rect 8352 31096 8493 31124
rect 8352 31084 8358 31096
rect 8481 31093 8493 31096
rect 8527 31124 8539 31127
rect 8846 31124 8852 31136
rect 8527 31096 8852 31124
rect 8527 31093 8539 31096
rect 8481 31087 8539 31093
rect 8846 31084 8852 31096
rect 8904 31084 8910 31136
rect 9950 31084 9956 31136
rect 10008 31124 10014 31136
rect 10413 31127 10471 31133
rect 10413 31124 10425 31127
rect 10008 31096 10425 31124
rect 10008 31084 10014 31096
rect 10413 31093 10425 31096
rect 10459 31093 10471 31127
rect 10413 31087 10471 31093
rect 552 31034 11132 31056
rect 552 30982 4322 31034
rect 4374 30982 4386 31034
rect 4438 30982 4450 31034
rect 4502 30982 4514 31034
rect 4566 30982 4578 31034
rect 4630 30982 10722 31034
rect 10774 30982 10786 31034
rect 10838 30982 10850 31034
rect 10902 30982 10914 31034
rect 10966 30982 10978 31034
rect 11030 30982 11132 31034
rect 552 30960 11132 30982
rect 1026 30880 1032 30932
rect 1084 30880 1090 30932
rect 1946 30920 1952 30932
rect 1412 30892 1952 30920
rect 1197 30855 1255 30861
rect 1197 30821 1209 30855
rect 1243 30852 1255 30855
rect 1302 30852 1308 30864
rect 1243 30824 1308 30852
rect 1243 30821 1255 30824
rect 1197 30815 1255 30821
rect 1302 30812 1308 30824
rect 1360 30812 1366 30864
rect 1412 30861 1440 30892
rect 1946 30880 1952 30892
rect 2004 30880 2010 30932
rect 2958 30880 2964 30932
rect 3016 30920 3022 30932
rect 3326 30929 3332 30932
rect 3145 30923 3203 30929
rect 3145 30920 3157 30923
rect 3016 30892 3157 30920
rect 3016 30880 3022 30892
rect 3145 30889 3157 30892
rect 3191 30889 3203 30923
rect 3145 30883 3203 30889
rect 3313 30923 3332 30929
rect 3313 30889 3325 30923
rect 3313 30883 3332 30889
rect 1397 30855 1455 30861
rect 1397 30821 1409 30855
rect 1443 30821 1455 30855
rect 1397 30815 1455 30821
rect 1857 30855 1915 30861
rect 1857 30821 1869 30855
rect 1903 30852 1915 30855
rect 2501 30855 2559 30861
rect 2501 30852 2513 30855
rect 1903 30824 2513 30852
rect 1903 30821 1915 30824
rect 1857 30815 1915 30821
rect 2501 30821 2513 30824
rect 2547 30852 2559 30855
rect 3160 30852 3188 30883
rect 3326 30880 3332 30883
rect 3384 30880 3390 30932
rect 4065 30923 4123 30929
rect 4065 30889 4077 30923
rect 4111 30920 4123 30923
rect 4154 30920 4160 30932
rect 4111 30892 4160 30920
rect 4111 30889 4123 30892
rect 4065 30883 4123 30889
rect 4154 30880 4160 30892
rect 4212 30880 4218 30932
rect 4430 30880 4436 30932
rect 4488 30920 4494 30932
rect 5537 30923 5595 30929
rect 5537 30920 5549 30923
rect 4488 30892 5549 30920
rect 4488 30880 4494 30892
rect 5537 30889 5549 30892
rect 5583 30920 5595 30923
rect 5718 30920 5724 30932
rect 5583 30892 5724 30920
rect 5583 30889 5595 30892
rect 5537 30883 5595 30889
rect 5718 30880 5724 30892
rect 5776 30880 5782 30932
rect 6365 30923 6423 30929
rect 6365 30889 6377 30923
rect 6411 30920 6423 30923
rect 6454 30920 6460 30932
rect 6411 30892 6460 30920
rect 6411 30889 6423 30892
rect 6365 30883 6423 30889
rect 6454 30880 6460 30892
rect 6512 30880 6518 30932
rect 6549 30923 6607 30929
rect 6549 30889 6561 30923
rect 6595 30920 6607 30923
rect 6638 30920 6644 30932
rect 6595 30892 6644 30920
rect 6595 30889 6607 30892
rect 6549 30883 6607 30889
rect 6638 30880 6644 30892
rect 6696 30880 6702 30932
rect 6730 30880 6736 30932
rect 6788 30920 6794 30932
rect 7374 30920 7380 30932
rect 6788 30892 7380 30920
rect 6788 30880 6794 30892
rect 7374 30880 7380 30892
rect 7432 30880 7438 30932
rect 8938 30880 8944 30932
rect 8996 30920 9002 30932
rect 9401 30923 9459 30929
rect 9401 30920 9413 30923
rect 8996 30892 9413 30920
rect 8996 30880 9002 30892
rect 9401 30889 9413 30892
rect 9447 30889 9459 30923
rect 9401 30883 9459 30889
rect 3418 30852 3424 30864
rect 2547 30824 3096 30852
rect 3160 30824 3424 30852
rect 2547 30821 2559 30824
rect 2501 30815 2559 30821
rect 1486 30744 1492 30796
rect 1544 30784 1550 30796
rect 1673 30787 1731 30793
rect 1673 30784 1685 30787
rect 1544 30756 1685 30784
rect 1544 30744 1550 30756
rect 1673 30753 1685 30756
rect 1719 30753 1731 30787
rect 1673 30747 1731 30753
rect 1946 30744 1952 30796
rect 2004 30744 2010 30796
rect 2038 30744 2044 30796
rect 2096 30744 2102 30796
rect 2133 30787 2191 30793
rect 2133 30753 2145 30787
rect 2179 30753 2191 30787
rect 2133 30747 2191 30753
rect 2317 30787 2375 30793
rect 2317 30753 2329 30787
rect 2363 30784 2375 30787
rect 2590 30784 2596 30796
rect 2363 30756 2596 30784
rect 2363 30753 2375 30756
rect 2317 30747 2375 30753
rect 1026 30676 1032 30728
rect 1084 30716 1090 30728
rect 2148 30716 2176 30747
rect 2590 30744 2596 30756
rect 2648 30744 2654 30796
rect 2682 30744 2688 30796
rect 2740 30784 2746 30796
rect 2777 30787 2835 30793
rect 2777 30784 2789 30787
rect 2740 30756 2789 30784
rect 2740 30744 2746 30756
rect 2777 30753 2789 30756
rect 2823 30753 2835 30787
rect 3068 30784 3096 30824
rect 3418 30812 3424 30824
rect 3476 30812 3482 30864
rect 3510 30812 3516 30864
rect 3568 30812 3574 30864
rect 4246 30812 4252 30864
rect 4304 30852 4310 30864
rect 5736 30852 5764 30880
rect 4304 30824 5488 30852
rect 5736 30824 6500 30852
rect 4304 30812 4310 30824
rect 3068 30756 3556 30784
rect 2777 30747 2835 30753
rect 3528 30728 3556 30756
rect 5350 30744 5356 30796
rect 5408 30744 5414 30796
rect 5460 30793 5488 30824
rect 5445 30787 5503 30793
rect 5445 30753 5457 30787
rect 5491 30753 5503 30787
rect 5445 30747 5503 30753
rect 5534 30744 5540 30796
rect 5592 30784 5598 30796
rect 5810 30784 5816 30796
rect 5592 30756 5816 30784
rect 5592 30744 5598 30756
rect 5810 30744 5816 30756
rect 5868 30744 5874 30796
rect 6472 30793 6500 30824
rect 6564 30824 6914 30852
rect 6457 30787 6515 30793
rect 6457 30753 6469 30787
rect 6503 30753 6515 30787
rect 6457 30747 6515 30753
rect 1084 30688 2176 30716
rect 1084 30676 1090 30688
rect 2222 30676 2228 30728
rect 2280 30716 2286 30728
rect 3053 30719 3111 30725
rect 3053 30716 3065 30719
rect 2280 30688 3065 30716
rect 2280 30676 2286 30688
rect 3053 30685 3065 30688
rect 3099 30685 3111 30719
rect 3053 30679 3111 30685
rect 3510 30676 3516 30728
rect 3568 30676 3574 30728
rect 4890 30716 4896 30728
rect 3896 30688 4896 30716
rect 1578 30608 1584 30660
rect 1636 30648 1642 30660
rect 2774 30648 2780 30660
rect 1636 30620 2780 30648
rect 1636 30608 1642 30620
rect 2774 30608 2780 30620
rect 2832 30608 2838 30660
rect 1213 30583 1271 30589
rect 1213 30549 1225 30583
rect 1259 30580 1271 30583
rect 1394 30580 1400 30592
rect 1259 30552 1400 30580
rect 1259 30549 1271 30552
rect 1213 30543 1271 30549
rect 1394 30540 1400 30552
rect 1452 30540 1458 30592
rect 1489 30583 1547 30589
rect 1489 30549 1501 30583
rect 1535 30580 1547 30583
rect 1670 30580 1676 30592
rect 1535 30552 1676 30580
rect 1535 30549 1547 30552
rect 1489 30543 1547 30549
rect 1670 30540 1676 30552
rect 1728 30540 1734 30592
rect 1762 30540 1768 30592
rect 1820 30580 1826 30592
rect 2593 30583 2651 30589
rect 2593 30580 2605 30583
rect 1820 30552 2605 30580
rect 1820 30540 1826 30552
rect 2593 30549 2605 30552
rect 2639 30549 2651 30583
rect 2593 30543 2651 30549
rect 2958 30540 2964 30592
rect 3016 30540 3022 30592
rect 3329 30583 3387 30589
rect 3329 30549 3341 30583
rect 3375 30580 3387 30583
rect 3896 30580 3924 30688
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 4982 30676 4988 30728
rect 5040 30716 5046 30728
rect 6089 30719 6147 30725
rect 6089 30716 6101 30719
rect 5040 30688 6101 30716
rect 5040 30676 5046 30688
rect 6089 30685 6101 30688
rect 6135 30685 6147 30719
rect 6089 30679 6147 30685
rect 6270 30676 6276 30728
rect 6328 30716 6334 30728
rect 6564 30716 6592 30824
rect 6641 30787 6699 30793
rect 6641 30753 6653 30787
rect 6687 30753 6699 30787
rect 6886 30784 6914 30824
rect 7282 30812 7288 30864
rect 7340 30852 7346 30864
rect 7340 30824 7696 30852
rect 7340 30812 7346 30824
rect 7377 30787 7435 30793
rect 7377 30784 7389 30787
rect 6886 30756 7389 30784
rect 6641 30747 6699 30753
rect 7377 30753 7389 30756
rect 7423 30753 7435 30787
rect 7377 30747 7435 30753
rect 6328 30688 6592 30716
rect 6328 30676 6334 30688
rect 3970 30608 3976 30660
rect 4028 30648 4034 30660
rect 4338 30648 4344 30660
rect 4028 30620 4344 30648
rect 4028 30608 4034 30620
rect 4338 30608 4344 30620
rect 4396 30608 4402 30660
rect 5626 30608 5632 30660
rect 5684 30648 5690 30660
rect 6656 30648 6684 30747
rect 7558 30744 7564 30796
rect 7616 30744 7622 30796
rect 7668 30784 7696 30824
rect 7742 30812 7748 30864
rect 7800 30852 7806 30864
rect 7800 30824 8984 30852
rect 7800 30812 7806 30824
rect 8021 30787 8079 30793
rect 8021 30784 8033 30787
rect 7668 30756 8033 30784
rect 8021 30753 8033 30756
rect 8067 30753 8079 30787
rect 8021 30747 8079 30753
rect 8110 30744 8116 30796
rect 8168 30784 8174 30796
rect 8205 30787 8263 30793
rect 8205 30784 8217 30787
rect 8168 30756 8217 30784
rect 8168 30744 8174 30756
rect 8205 30753 8217 30756
rect 8251 30753 8263 30787
rect 8205 30747 8263 30753
rect 8294 30744 8300 30796
rect 8352 30744 8358 30796
rect 8956 30793 8984 30824
rect 9674 30812 9680 30864
rect 9732 30852 9738 30864
rect 10514 30855 10572 30861
rect 10514 30852 10526 30855
rect 9732 30824 10526 30852
rect 9732 30812 9738 30824
rect 10514 30821 10526 30824
rect 10560 30821 10572 30855
rect 10514 30815 10572 30821
rect 8941 30787 8999 30793
rect 8941 30753 8953 30787
rect 8987 30753 8999 30787
rect 8941 30747 8999 30753
rect 7098 30676 7104 30728
rect 7156 30676 7162 30728
rect 7285 30719 7343 30725
rect 7285 30685 7297 30719
rect 7331 30716 7343 30719
rect 9766 30716 9772 30728
rect 7331 30688 9772 30716
rect 7331 30685 7343 30688
rect 7285 30679 7343 30685
rect 9766 30676 9772 30688
rect 9824 30676 9830 30728
rect 10781 30719 10839 30725
rect 10781 30685 10793 30719
rect 10827 30685 10839 30719
rect 10781 30679 10839 30685
rect 5684 30620 6684 30648
rect 5684 30608 5690 30620
rect 7558 30608 7564 30660
rect 7616 30648 7622 30660
rect 8113 30651 8171 30657
rect 8113 30648 8125 30651
rect 7616 30620 8125 30648
rect 7616 30608 7622 30620
rect 8113 30617 8125 30620
rect 8159 30617 8171 30651
rect 8113 30611 8171 30617
rect 3375 30552 3924 30580
rect 3375 30549 3387 30552
rect 3329 30543 3387 30549
rect 4246 30540 4252 30592
rect 4304 30580 4310 30592
rect 4798 30580 4804 30592
rect 4304 30552 4804 30580
rect 4304 30540 4310 30552
rect 4798 30540 4804 30552
rect 4856 30540 4862 30592
rect 6178 30540 6184 30592
rect 6236 30540 6242 30592
rect 6546 30540 6552 30592
rect 6604 30580 6610 30592
rect 6917 30583 6975 30589
rect 6917 30580 6929 30583
rect 6604 30552 6929 30580
rect 6604 30540 6610 30552
rect 6917 30549 6929 30552
rect 6963 30549 6975 30583
rect 6917 30543 6975 30549
rect 7466 30540 7472 30592
rect 7524 30580 7530 30592
rect 7653 30583 7711 30589
rect 7653 30580 7665 30583
rect 7524 30552 7665 30580
rect 7524 30540 7530 30552
rect 7653 30549 7665 30552
rect 7699 30549 7711 30583
rect 7653 30543 7711 30549
rect 8386 30540 8392 30592
rect 8444 30580 8450 30592
rect 8938 30580 8944 30592
rect 8444 30552 8944 30580
rect 8444 30540 8450 30552
rect 8938 30540 8944 30552
rect 8996 30540 9002 30592
rect 9217 30583 9275 30589
rect 9217 30549 9229 30583
rect 9263 30580 9275 30583
rect 9398 30580 9404 30592
rect 9263 30552 9404 30580
rect 9263 30549 9275 30552
rect 9217 30543 9275 30549
rect 9398 30540 9404 30552
rect 9456 30540 9462 30592
rect 10502 30540 10508 30592
rect 10560 30580 10566 30592
rect 10796 30580 10824 30679
rect 10560 30552 10824 30580
rect 10560 30540 10566 30552
rect 552 30490 11132 30512
rect 552 30438 3662 30490
rect 3714 30438 3726 30490
rect 3778 30438 3790 30490
rect 3842 30438 3854 30490
rect 3906 30438 3918 30490
rect 3970 30438 10062 30490
rect 10114 30438 10126 30490
rect 10178 30438 10190 30490
rect 10242 30438 10254 30490
rect 10306 30438 10318 30490
rect 10370 30438 11132 30490
rect 552 30416 11132 30438
rect 14 30336 20 30388
rect 72 30376 78 30388
rect 382 30376 388 30388
rect 72 30348 388 30376
rect 72 30336 78 30348
rect 382 30336 388 30348
rect 440 30336 446 30388
rect 1486 30336 1492 30388
rect 1544 30336 1550 30388
rect 2866 30336 2872 30388
rect 2924 30376 2930 30388
rect 2961 30379 3019 30385
rect 2961 30376 2973 30379
rect 2924 30348 2973 30376
rect 2924 30336 2930 30348
rect 2961 30345 2973 30348
rect 3007 30345 3019 30379
rect 2961 30339 3019 30345
rect 3234 30336 3240 30388
rect 3292 30376 3298 30388
rect 3973 30379 4031 30385
rect 3292 30348 3455 30376
rect 3292 30336 3298 30348
rect 1302 30268 1308 30320
rect 1360 30308 1366 30320
rect 3329 30311 3387 30317
rect 3329 30308 3341 30311
rect 1360 30280 3341 30308
rect 1360 30268 1366 30280
rect 3329 30277 3341 30280
rect 3375 30277 3387 30311
rect 3329 30271 3387 30277
rect 842 30200 848 30252
rect 900 30240 906 30252
rect 3427 30240 3455 30348
rect 3973 30345 3985 30379
rect 4019 30376 4031 30379
rect 4338 30376 4344 30388
rect 4019 30348 4344 30376
rect 4019 30345 4031 30348
rect 3973 30339 4031 30345
rect 4338 30336 4344 30348
rect 4396 30336 4402 30388
rect 4985 30379 5043 30385
rect 4985 30345 4997 30379
rect 5031 30376 5043 30379
rect 5074 30376 5080 30388
rect 5031 30348 5080 30376
rect 5031 30345 5043 30348
rect 4985 30339 5043 30345
rect 5074 30336 5080 30348
rect 5132 30336 5138 30388
rect 5169 30379 5227 30385
rect 5169 30345 5181 30379
rect 5215 30376 5227 30379
rect 5258 30376 5264 30388
rect 5215 30348 5264 30376
rect 5215 30345 5227 30348
rect 5169 30339 5227 30345
rect 5258 30336 5264 30348
rect 5316 30336 5322 30388
rect 5810 30336 5816 30388
rect 5868 30336 5874 30388
rect 5905 30379 5963 30385
rect 5905 30345 5917 30379
rect 5951 30376 5963 30379
rect 6086 30376 6092 30388
rect 5951 30348 6092 30376
rect 5951 30345 5963 30348
rect 5905 30339 5963 30345
rect 6086 30336 6092 30348
rect 6144 30336 6150 30388
rect 6181 30379 6239 30385
rect 6181 30345 6193 30379
rect 6227 30345 6239 30379
rect 6181 30339 6239 30345
rect 4157 30311 4215 30317
rect 4157 30277 4169 30311
rect 4203 30308 4215 30311
rect 4246 30308 4252 30320
rect 4203 30280 4252 30308
rect 4203 30277 4215 30280
rect 4157 30271 4215 30277
rect 4246 30268 4252 30280
rect 4304 30268 4310 30320
rect 5534 30308 5540 30320
rect 4632 30280 5540 30308
rect 900 30212 2728 30240
rect 900 30200 906 30212
rect 1949 30175 2007 30181
rect 1949 30141 1961 30175
rect 1995 30172 2007 30175
rect 2038 30172 2044 30184
rect 1995 30144 2044 30172
rect 1995 30141 2007 30144
rect 1949 30135 2007 30141
rect 2038 30132 2044 30144
rect 2096 30132 2102 30184
rect 2222 30132 2228 30184
rect 2280 30132 2286 30184
rect 1213 30107 1271 30113
rect 1213 30073 1225 30107
rect 1259 30104 1271 30107
rect 1578 30104 1584 30116
rect 1259 30076 1584 30104
rect 1259 30073 1271 30076
rect 1213 30067 1271 30073
rect 1578 30064 1584 30076
rect 1636 30064 1642 30116
rect 1673 30107 1731 30113
rect 1673 30073 1685 30107
rect 1719 30104 1731 30107
rect 1719 30076 2268 30104
rect 1719 30073 1731 30076
rect 1673 30067 1731 30073
rect 2240 30048 2268 30076
rect 2222 29996 2228 30048
rect 2280 29996 2286 30048
rect 2700 30036 2728 30212
rect 3068 30212 3455 30240
rect 2777 30175 2835 30181
rect 2777 30141 2789 30175
rect 2823 30141 2835 30175
rect 2777 30135 2835 30141
rect 2869 30175 2927 30181
rect 2869 30141 2881 30175
rect 2915 30172 2927 30175
rect 2958 30172 2964 30184
rect 2915 30144 2964 30172
rect 2915 30141 2927 30144
rect 2869 30135 2927 30141
rect 2792 30104 2820 30135
rect 2958 30132 2964 30144
rect 3016 30132 3022 30184
rect 3068 30181 3096 30212
rect 3053 30175 3111 30181
rect 3053 30141 3065 30175
rect 3099 30141 3111 30175
rect 3053 30135 3111 30141
rect 3237 30175 3295 30181
rect 3237 30141 3249 30175
rect 3283 30172 3295 30175
rect 3326 30172 3332 30184
rect 3283 30144 3332 30172
rect 3283 30141 3295 30144
rect 3237 30135 3295 30141
rect 3142 30104 3148 30116
rect 2792 30076 3148 30104
rect 3142 30064 3148 30076
rect 3200 30064 3206 30116
rect 3252 30036 3280 30135
rect 3326 30132 3332 30144
rect 3384 30132 3390 30184
rect 3418 30132 3424 30184
rect 3476 30172 3482 30184
rect 3605 30175 3663 30181
rect 3605 30172 3617 30175
rect 3476 30144 3617 30172
rect 3476 30132 3482 30144
rect 3605 30141 3617 30144
rect 3651 30141 3663 30175
rect 3605 30135 3663 30141
rect 3878 30132 3884 30184
rect 3936 30172 3942 30184
rect 4341 30175 4399 30181
rect 4341 30172 4353 30175
rect 3936 30144 4353 30172
rect 3936 30132 3942 30144
rect 4341 30141 4353 30144
rect 4387 30141 4399 30175
rect 4341 30135 4399 30141
rect 4430 30132 4436 30184
rect 4488 30172 4494 30184
rect 4632 30181 4660 30280
rect 5534 30268 5540 30280
rect 5592 30268 5598 30320
rect 5828 30308 5856 30336
rect 6196 30308 6224 30339
rect 6454 30336 6460 30388
rect 6512 30376 6518 30388
rect 7190 30376 7196 30388
rect 6512 30348 7196 30376
rect 6512 30336 6518 30348
rect 7190 30336 7196 30348
rect 7248 30336 7254 30388
rect 8294 30336 8300 30388
rect 8352 30376 8358 30388
rect 9582 30376 9588 30388
rect 8352 30348 9588 30376
rect 8352 30336 8358 30348
rect 9582 30336 9588 30348
rect 9640 30376 9646 30388
rect 9677 30379 9735 30385
rect 9677 30376 9689 30379
rect 9640 30348 9689 30376
rect 9640 30336 9646 30348
rect 9677 30345 9689 30348
rect 9723 30345 9735 30379
rect 10413 30379 10471 30385
rect 10413 30376 10425 30379
rect 9677 30339 9735 30345
rect 9784 30348 10425 30376
rect 5828 30280 6224 30308
rect 6546 30268 6552 30320
rect 6604 30308 6610 30320
rect 6914 30308 6920 30320
rect 6604 30280 6920 30308
rect 6604 30268 6610 30280
rect 6914 30268 6920 30280
rect 6972 30268 6978 30320
rect 8202 30308 8208 30320
rect 7852 30280 8208 30308
rect 4798 30200 4804 30252
rect 4856 30240 4862 30252
rect 5074 30240 5080 30252
rect 4856 30212 5080 30240
rect 4856 30200 4862 30212
rect 5074 30200 5080 30212
rect 5132 30200 5138 30252
rect 5350 30200 5356 30252
rect 5408 30240 5414 30252
rect 7190 30240 7196 30252
rect 5408 30212 6850 30240
rect 5408 30200 5414 30212
rect 4525 30175 4583 30181
rect 4525 30172 4537 30175
rect 4488 30144 4537 30172
rect 4488 30132 4494 30144
rect 4525 30141 4537 30144
rect 4571 30141 4583 30175
rect 4525 30135 4583 30141
rect 4617 30175 4675 30181
rect 4617 30141 4629 30175
rect 4663 30172 4675 30175
rect 4663 30144 4844 30172
rect 4663 30141 4675 30144
rect 4617 30135 4675 30141
rect 4816 30116 4844 30144
rect 4890 30132 4896 30184
rect 4948 30132 4954 30184
rect 5718 30132 5724 30184
rect 5776 30172 5782 30184
rect 5813 30175 5871 30181
rect 5813 30172 5825 30175
rect 5776 30144 5825 30172
rect 5776 30132 5782 30144
rect 5813 30141 5825 30144
rect 5859 30141 5871 30175
rect 5813 30135 5871 30141
rect 5902 30132 5908 30184
rect 5960 30172 5966 30184
rect 5997 30175 6055 30181
rect 5997 30172 6009 30175
rect 5960 30144 6009 30172
rect 5960 30132 5966 30144
rect 5997 30141 6009 30144
rect 6043 30141 6055 30175
rect 5997 30135 6055 30141
rect 6086 30132 6092 30184
rect 6144 30132 6150 30184
rect 6178 30132 6184 30184
rect 6236 30172 6242 30184
rect 6457 30175 6515 30181
rect 6457 30172 6469 30175
rect 6236 30144 6469 30172
rect 6236 30132 6242 30144
rect 6457 30141 6469 30144
rect 6503 30172 6515 30175
rect 6546 30172 6552 30184
rect 6503 30144 6552 30172
rect 6503 30141 6515 30144
rect 6457 30135 6515 30141
rect 6546 30132 6552 30144
rect 6604 30132 6610 30184
rect 6733 30175 6791 30181
rect 6733 30172 6745 30175
rect 6656 30144 6745 30172
rect 3973 30107 4031 30113
rect 3973 30073 3985 30107
rect 4019 30104 4031 30107
rect 4706 30104 4712 30116
rect 4019 30076 4712 30104
rect 4019 30073 4031 30076
rect 3973 30067 4031 30073
rect 4706 30064 4712 30076
rect 4764 30064 4770 30116
rect 4798 30064 4804 30116
rect 4856 30064 4862 30116
rect 5166 30064 5172 30116
rect 5224 30104 5230 30116
rect 5353 30107 5411 30113
rect 5353 30104 5365 30107
rect 5224 30076 5365 30104
rect 5224 30064 5230 30076
rect 5353 30073 5365 30076
rect 5399 30073 5411 30107
rect 5353 30067 5411 30073
rect 2700 30008 3280 30036
rect 4246 29996 4252 30048
rect 4304 30036 4310 30048
rect 4433 30039 4491 30045
rect 4433 30036 4445 30039
rect 4304 30008 4445 30036
rect 4304 29996 4310 30008
rect 4433 30005 4445 30008
rect 4479 30005 4491 30039
rect 4433 29999 4491 30005
rect 5445 30039 5503 30045
rect 5445 30005 5457 30039
rect 5491 30036 5503 30039
rect 5534 30036 5540 30048
rect 5491 30008 5540 30036
rect 5491 30005 5503 30008
rect 5445 29999 5503 30005
rect 5534 29996 5540 30008
rect 5592 29996 5598 30048
rect 6656 30045 6684 30144
rect 6733 30141 6745 30144
rect 6779 30141 6791 30175
rect 6733 30135 6791 30141
rect 6822 30104 6850 30212
rect 7024 30212 7196 30240
rect 6914 30132 6920 30184
rect 6972 30132 6978 30184
rect 7024 30181 7052 30212
rect 7190 30200 7196 30212
rect 7248 30200 7254 30252
rect 7852 30181 7880 30280
rect 8202 30268 8208 30280
rect 8260 30308 8266 30320
rect 9784 30308 9812 30348
rect 10413 30345 10425 30348
rect 10459 30345 10471 30379
rect 10413 30339 10471 30345
rect 8260 30280 9812 30308
rect 8260 30268 8266 30280
rect 8662 30200 8668 30252
rect 8720 30240 8726 30252
rect 8846 30240 8852 30252
rect 8720 30212 8852 30240
rect 8720 30200 8726 30212
rect 8846 30200 8852 30212
rect 8904 30200 8910 30252
rect 7009 30175 7067 30181
rect 7009 30141 7021 30175
rect 7055 30141 7067 30175
rect 7009 30135 7067 30141
rect 7101 30175 7159 30181
rect 7101 30141 7113 30175
rect 7147 30172 7159 30175
rect 7837 30175 7895 30181
rect 7837 30172 7849 30175
rect 7147 30144 7849 30172
rect 7147 30141 7159 30144
rect 7101 30135 7159 30141
rect 7837 30141 7849 30144
rect 7883 30141 7895 30175
rect 7837 30135 7895 30141
rect 7926 30132 7932 30184
rect 7984 30132 7990 30184
rect 8021 30175 8079 30181
rect 8021 30141 8033 30175
rect 8067 30141 8079 30175
rect 8021 30135 8079 30141
rect 8036 30104 8064 30135
rect 8202 30132 8208 30184
rect 8260 30132 8266 30184
rect 9122 30132 9128 30184
rect 9180 30172 9186 30184
rect 9180 30144 10640 30172
rect 9180 30132 9186 30144
rect 8294 30104 8300 30116
rect 6822 30076 7880 30104
rect 8036 30076 8300 30104
rect 6641 30039 6699 30045
rect 6641 30005 6653 30039
rect 6687 30005 6699 30039
rect 6641 29999 6699 30005
rect 7377 30039 7435 30045
rect 7377 30005 7389 30039
rect 7423 30036 7435 30039
rect 7466 30036 7472 30048
rect 7423 30008 7472 30036
rect 7423 30005 7435 30008
rect 7377 29999 7435 30005
rect 7466 29996 7472 30008
rect 7524 29996 7530 30048
rect 7561 30039 7619 30045
rect 7561 30005 7573 30039
rect 7607 30036 7619 30039
rect 7742 30036 7748 30048
rect 7607 30008 7748 30036
rect 7607 30005 7619 30008
rect 7561 29999 7619 30005
rect 7742 29996 7748 30008
rect 7800 29996 7806 30048
rect 7852 30036 7880 30076
rect 8294 30064 8300 30076
rect 8352 30064 8358 30116
rect 8389 30107 8447 30113
rect 8389 30073 8401 30107
rect 8435 30104 8447 30107
rect 8478 30104 8484 30116
rect 8435 30076 8484 30104
rect 8435 30073 8447 30076
rect 8389 30067 8447 30073
rect 8404 30036 8432 30067
rect 8478 30064 8484 30076
rect 8536 30064 8542 30116
rect 9214 30064 9220 30116
rect 9272 30104 9278 30116
rect 10612 30113 10640 30144
rect 10597 30107 10655 30113
rect 9272 30076 10364 30104
rect 9272 30064 9278 30076
rect 7852 30008 8432 30036
rect 10226 29996 10232 30048
rect 10284 29996 10290 30048
rect 10336 30036 10364 30076
rect 10597 30073 10609 30107
rect 10643 30073 10655 30107
rect 10597 30067 10655 30073
rect 10397 30039 10455 30045
rect 10397 30036 10409 30039
rect 10336 30008 10409 30036
rect 10397 30005 10409 30008
rect 10443 30036 10455 30039
rect 11330 30036 11336 30048
rect 10443 30008 11336 30036
rect 10443 30005 10455 30008
rect 10397 29999 10455 30005
rect 11330 29996 11336 30008
rect 11388 29996 11394 30048
rect 552 29946 11132 29968
rect 552 29894 4322 29946
rect 4374 29894 4386 29946
rect 4438 29894 4450 29946
rect 4502 29894 4514 29946
rect 4566 29894 4578 29946
rect 4630 29894 10722 29946
rect 10774 29894 10786 29946
rect 10838 29894 10850 29946
rect 10902 29894 10914 29946
rect 10966 29894 10978 29946
rect 11030 29894 11132 29946
rect 552 29872 11132 29894
rect 2222 29792 2228 29844
rect 2280 29832 2286 29844
rect 2590 29832 2596 29844
rect 2280 29804 2596 29832
rect 2280 29792 2286 29804
rect 2590 29792 2596 29804
rect 2648 29792 2654 29844
rect 2866 29792 2872 29844
rect 2924 29792 2930 29844
rect 3145 29835 3203 29841
rect 3145 29801 3157 29835
rect 3191 29832 3203 29835
rect 4249 29835 4307 29841
rect 3191 29804 4200 29832
rect 3191 29801 3203 29804
rect 3145 29795 3203 29801
rect 937 29767 995 29773
rect 937 29733 949 29767
rect 983 29764 995 29767
rect 2777 29767 2835 29773
rect 2777 29764 2789 29767
rect 983 29736 2789 29764
rect 983 29733 995 29736
rect 937 29727 995 29733
rect 2777 29733 2789 29736
rect 2823 29733 2835 29767
rect 2884 29764 2912 29792
rect 2884 29736 3372 29764
rect 2777 29727 2835 29733
rect 3344 29708 3372 29736
rect 3418 29724 3424 29776
rect 3476 29724 3482 29776
rect 3513 29767 3571 29773
rect 3513 29733 3525 29767
rect 3559 29764 3571 29767
rect 4062 29764 4068 29776
rect 3559 29736 4068 29764
rect 3559 29733 3571 29736
rect 3513 29727 3571 29733
rect 4062 29724 4068 29736
rect 4120 29724 4126 29776
rect 4172 29764 4200 29804
rect 4249 29801 4261 29835
rect 4295 29832 4307 29835
rect 4798 29832 4804 29844
rect 4295 29804 4804 29832
rect 4295 29801 4307 29804
rect 4249 29795 4307 29801
rect 4798 29792 4804 29804
rect 4856 29792 4862 29844
rect 4893 29835 4951 29841
rect 4893 29801 4905 29835
rect 4939 29832 4951 29835
rect 5442 29832 5448 29844
rect 4939 29804 5448 29832
rect 4939 29801 4951 29804
rect 4893 29795 4951 29801
rect 4338 29764 4344 29776
rect 4172 29736 4344 29764
rect 4338 29724 4344 29736
rect 4396 29764 4402 29776
rect 4908 29764 4936 29795
rect 5442 29792 5448 29804
rect 5500 29792 5506 29844
rect 5626 29792 5632 29844
rect 5684 29832 5690 29844
rect 5813 29835 5871 29841
rect 5813 29832 5825 29835
rect 5684 29804 5825 29832
rect 5684 29792 5690 29804
rect 5813 29801 5825 29804
rect 5859 29801 5871 29835
rect 5813 29795 5871 29801
rect 4396 29736 4936 29764
rect 4396 29724 4402 29736
rect 1670 29656 1676 29708
rect 1728 29656 1734 29708
rect 1762 29656 1768 29708
rect 1820 29656 1826 29708
rect 1854 29656 1860 29708
rect 1912 29656 1918 29708
rect 2041 29699 2099 29705
rect 2041 29665 2053 29699
rect 2087 29665 2099 29699
rect 2041 29659 2099 29665
rect 1210 29588 1216 29640
rect 1268 29588 1274 29640
rect 2056 29628 2084 29659
rect 2222 29656 2228 29708
rect 2280 29696 2286 29708
rect 2409 29699 2467 29705
rect 2409 29696 2421 29699
rect 2280 29668 2421 29696
rect 2280 29656 2286 29668
rect 2409 29665 2421 29668
rect 2455 29665 2467 29699
rect 2409 29659 2467 29665
rect 2685 29699 2743 29705
rect 2685 29665 2697 29699
rect 2731 29665 2743 29699
rect 2685 29659 2743 29665
rect 1780 29600 2084 29628
rect 1121 29563 1179 29569
rect 1121 29529 1133 29563
rect 1167 29560 1179 29563
rect 1670 29560 1676 29572
rect 1167 29532 1676 29560
rect 1167 29529 1179 29532
rect 1121 29523 1179 29529
rect 1670 29520 1676 29532
rect 1728 29520 1734 29572
rect 14 29452 20 29504
rect 72 29492 78 29504
rect 1780 29492 1808 29600
rect 2130 29588 2136 29640
rect 2188 29588 2194 29640
rect 2314 29588 2320 29640
rect 2372 29628 2378 29640
rect 2700 29628 2728 29659
rect 2866 29656 2872 29708
rect 2924 29656 2930 29708
rect 3326 29656 3332 29708
rect 3384 29696 3390 29708
rect 3881 29699 3939 29705
rect 3881 29696 3893 29699
rect 3384 29668 3893 29696
rect 3384 29656 3390 29668
rect 3881 29665 3893 29668
rect 3927 29696 3939 29699
rect 4890 29696 4896 29708
rect 3927 29668 4896 29696
rect 3927 29665 3939 29668
rect 3881 29659 3939 29665
rect 4890 29656 4896 29668
rect 4948 29696 4954 29708
rect 4985 29699 5043 29705
rect 4985 29696 4997 29699
rect 4948 29668 4997 29696
rect 4948 29656 4954 29668
rect 4985 29665 4997 29668
rect 5031 29696 5043 29699
rect 5350 29696 5356 29708
rect 5031 29668 5356 29696
rect 5031 29665 5043 29668
rect 4985 29659 5043 29665
rect 5350 29656 5356 29668
rect 5408 29656 5414 29708
rect 5626 29656 5632 29708
rect 5684 29656 5690 29708
rect 2372 29600 2728 29628
rect 3148 29640 3200 29646
rect 2372 29588 2378 29600
rect 4706 29588 4712 29640
rect 4764 29588 4770 29640
rect 3148 29582 3200 29588
rect 2041 29563 2099 29569
rect 2041 29529 2053 29563
rect 2087 29560 2099 29563
rect 5828 29560 5856 29795
rect 6086 29792 6092 29844
rect 6144 29832 6150 29844
rect 6144 29804 6776 29832
rect 6144 29792 6150 29804
rect 5997 29767 6055 29773
rect 5997 29733 6009 29767
rect 6043 29764 6055 29767
rect 6043 29736 6500 29764
rect 6043 29733 6055 29736
rect 5997 29727 6055 29733
rect 6472 29708 6500 29736
rect 6748 29708 6776 29804
rect 7098 29792 7104 29844
rect 7156 29832 7162 29844
rect 7285 29835 7343 29841
rect 7285 29832 7297 29835
rect 7156 29804 7297 29832
rect 7156 29792 7162 29804
rect 7285 29801 7297 29804
rect 7331 29801 7343 29835
rect 7285 29795 7343 29801
rect 8021 29835 8079 29841
rect 8021 29801 8033 29835
rect 8067 29832 8079 29835
rect 8202 29832 8208 29844
rect 8067 29804 8208 29832
rect 8067 29801 8079 29804
rect 8021 29795 8079 29801
rect 8202 29792 8208 29804
rect 8260 29792 8266 29844
rect 8570 29792 8576 29844
rect 8628 29832 8634 29844
rect 8941 29835 8999 29841
rect 8941 29832 8953 29835
rect 8628 29804 8953 29832
rect 8628 29792 8634 29804
rect 8941 29801 8953 29804
rect 8987 29801 8999 29835
rect 9306 29832 9312 29844
rect 8941 29795 8999 29801
rect 9048 29804 9312 29832
rect 9048 29764 9076 29804
rect 9306 29792 9312 29804
rect 9364 29832 9370 29844
rect 11238 29832 11244 29844
rect 9364 29804 11244 29832
rect 9364 29792 9370 29804
rect 11238 29792 11244 29804
rect 11296 29792 11302 29844
rect 6886 29736 8616 29764
rect 6181 29699 6239 29705
rect 6181 29665 6193 29699
rect 6227 29696 6239 29699
rect 6273 29699 6331 29705
rect 6273 29696 6285 29699
rect 6227 29668 6285 29696
rect 6227 29665 6239 29668
rect 6181 29659 6239 29665
rect 6273 29665 6285 29668
rect 6319 29696 6331 29699
rect 6362 29696 6368 29708
rect 6319 29668 6368 29696
rect 6319 29665 6331 29668
rect 6273 29659 6331 29665
rect 6362 29656 6368 29668
rect 6420 29656 6426 29708
rect 6454 29656 6460 29708
rect 6512 29656 6518 29708
rect 6546 29656 6552 29708
rect 6604 29696 6610 29708
rect 6641 29699 6699 29705
rect 6641 29696 6653 29699
rect 6604 29668 6653 29696
rect 6604 29656 6610 29668
rect 6641 29665 6653 29668
rect 6687 29665 6699 29699
rect 6641 29659 6699 29665
rect 6656 29628 6684 29659
rect 6730 29656 6736 29708
rect 6788 29696 6794 29708
rect 6886 29696 6914 29736
rect 7024 29705 7052 29736
rect 6788 29668 6914 29696
rect 7009 29699 7067 29705
rect 6788 29656 6794 29668
rect 7009 29665 7021 29699
rect 7055 29696 7067 29699
rect 7055 29668 7089 29696
rect 7055 29665 7067 29668
rect 7009 29659 7067 29665
rect 7466 29656 7472 29708
rect 7524 29656 7530 29708
rect 7561 29699 7619 29705
rect 7561 29665 7573 29699
rect 7607 29696 7619 29699
rect 7650 29696 7656 29708
rect 7607 29668 7656 29696
rect 7607 29665 7619 29668
rect 7561 29659 7619 29665
rect 7650 29656 7656 29668
rect 7708 29656 7714 29708
rect 7834 29656 7840 29708
rect 7892 29656 7898 29708
rect 8588 29705 8616 29736
rect 8864 29736 9076 29764
rect 8573 29699 8631 29705
rect 8573 29665 8585 29699
rect 8619 29665 8631 29699
rect 8573 29659 8631 29665
rect 6656 29600 7696 29628
rect 6638 29560 6644 29572
rect 2087 29532 3004 29560
rect 5828 29532 6644 29560
rect 2087 29529 2099 29532
rect 2041 29523 2099 29529
rect 2976 29504 3004 29532
rect 6638 29520 6644 29532
rect 6696 29520 6702 29572
rect 7466 29520 7472 29572
rect 7524 29560 7530 29572
rect 7668 29560 7696 29600
rect 7742 29588 7748 29640
rect 7800 29588 7806 29640
rect 8297 29631 8355 29637
rect 8297 29597 8309 29631
rect 8343 29597 8355 29631
rect 8588 29628 8616 29659
rect 8662 29656 8668 29708
rect 8720 29696 8726 29708
rect 8864 29705 8892 29736
rect 9398 29724 9404 29776
rect 9456 29764 9462 29776
rect 9950 29764 9956 29776
rect 9456 29736 9956 29764
rect 9456 29724 9462 29736
rect 9950 29724 9956 29736
rect 10008 29724 10014 29776
rect 10076 29767 10134 29773
rect 10076 29733 10088 29767
rect 10122 29764 10134 29767
rect 10226 29764 10232 29776
rect 10122 29736 10232 29764
rect 10122 29733 10134 29736
rect 10076 29727 10134 29733
rect 10226 29724 10232 29736
rect 10284 29724 10290 29776
rect 10336 29736 10548 29764
rect 8757 29699 8815 29705
rect 8757 29696 8769 29699
rect 8720 29668 8769 29696
rect 8720 29656 8726 29668
rect 8757 29665 8769 29668
rect 8803 29665 8815 29699
rect 8757 29659 8815 29665
rect 8849 29699 8907 29705
rect 8849 29665 8861 29699
rect 8895 29665 8907 29699
rect 10336 29696 10364 29736
rect 10520 29705 10548 29736
rect 8849 29659 8907 29665
rect 9048 29668 10364 29696
rect 10413 29699 10471 29705
rect 8938 29628 8944 29640
rect 8588 29600 8944 29628
rect 8297 29591 8355 29597
rect 8312 29560 8340 29591
rect 8938 29588 8944 29600
rect 8996 29588 9002 29640
rect 8570 29560 8576 29572
rect 7524 29532 8576 29560
rect 7524 29520 7530 29532
rect 8570 29520 8576 29532
rect 8628 29560 8634 29572
rect 9048 29560 9076 29668
rect 10413 29665 10425 29699
rect 10459 29665 10471 29699
rect 10413 29659 10471 29665
rect 10506 29699 10564 29705
rect 10506 29665 10518 29699
rect 10552 29665 10564 29699
rect 10506 29659 10564 29665
rect 10321 29631 10379 29637
rect 10321 29597 10333 29631
rect 10367 29597 10379 29631
rect 10428 29628 10456 29659
rect 10686 29628 10692 29640
rect 10428 29600 10692 29628
rect 10321 29591 10379 29597
rect 8628 29532 9076 29560
rect 10336 29560 10364 29591
rect 10686 29588 10692 29600
rect 10744 29588 10750 29640
rect 10502 29560 10508 29572
rect 10336 29532 10508 29560
rect 8628 29520 8634 29532
rect 72 29464 1808 29492
rect 2225 29495 2283 29501
rect 72 29452 78 29464
rect 2225 29461 2237 29495
rect 2271 29492 2283 29495
rect 2314 29492 2320 29504
rect 2271 29464 2320 29492
rect 2271 29461 2283 29464
rect 2225 29455 2283 29461
rect 2314 29452 2320 29464
rect 2372 29452 2378 29504
rect 2593 29495 2651 29501
rect 2593 29461 2605 29495
rect 2639 29492 2651 29495
rect 2682 29492 2688 29504
rect 2639 29464 2688 29492
rect 2639 29461 2651 29464
rect 2593 29455 2651 29461
rect 2682 29452 2688 29464
rect 2740 29452 2746 29504
rect 2958 29452 2964 29504
rect 3016 29452 3022 29504
rect 4433 29495 4491 29501
rect 4433 29461 4445 29495
rect 4479 29492 4491 29495
rect 4982 29492 4988 29504
rect 4479 29464 4988 29492
rect 4479 29461 4491 29464
rect 4433 29455 4491 29461
rect 4982 29452 4988 29464
rect 5040 29452 5046 29504
rect 5074 29452 5080 29504
rect 5132 29492 5138 29504
rect 5353 29495 5411 29501
rect 5353 29492 5365 29495
rect 5132 29464 5365 29492
rect 5132 29452 5138 29464
rect 5353 29461 5365 29464
rect 5399 29461 5411 29495
rect 5353 29455 5411 29461
rect 5537 29495 5595 29501
rect 5537 29461 5549 29495
rect 5583 29492 5595 29495
rect 5718 29492 5724 29504
rect 5583 29464 5724 29492
rect 5583 29461 5595 29464
rect 5537 29455 5595 29461
rect 5718 29452 5724 29464
rect 5776 29452 5782 29504
rect 6086 29452 6092 29504
rect 6144 29492 6150 29504
rect 6273 29495 6331 29501
rect 6273 29492 6285 29495
rect 6144 29464 6285 29492
rect 6144 29452 6150 29464
rect 6273 29461 6285 29464
rect 6319 29461 6331 29495
rect 6273 29455 6331 29461
rect 6362 29452 6368 29504
rect 6420 29492 6426 29504
rect 6822 29492 6828 29504
rect 6420 29464 6828 29492
rect 6420 29452 6426 29464
rect 6822 29452 6828 29464
rect 6880 29452 6886 29504
rect 7009 29495 7067 29501
rect 7009 29461 7021 29495
rect 7055 29492 7067 29495
rect 7098 29492 7104 29504
rect 7055 29464 7104 29492
rect 7055 29461 7067 29464
rect 7009 29455 7067 29461
rect 7098 29452 7104 29464
rect 7156 29452 7162 29504
rect 7190 29452 7196 29504
rect 7248 29452 7254 29504
rect 8481 29495 8539 29501
rect 8481 29461 8493 29495
rect 8527 29492 8539 29495
rect 9398 29492 9404 29504
rect 8527 29464 9404 29492
rect 8527 29461 8539 29464
rect 8481 29455 8539 29461
rect 9398 29452 9404 29464
rect 9456 29452 9462 29504
rect 9582 29452 9588 29504
rect 9640 29492 9646 29504
rect 9674 29492 9680 29504
rect 9640 29464 9680 29492
rect 9640 29452 9646 29464
rect 9674 29452 9680 29464
rect 9732 29492 9738 29504
rect 10336 29492 10364 29532
rect 10502 29520 10508 29532
rect 10560 29520 10566 29572
rect 9732 29464 10364 29492
rect 9732 29452 9738 29464
rect 10410 29452 10416 29504
rect 10468 29492 10474 29504
rect 10597 29495 10655 29501
rect 10597 29492 10609 29495
rect 10468 29464 10609 29492
rect 10468 29452 10474 29464
rect 10597 29461 10609 29464
rect 10643 29461 10655 29495
rect 10597 29455 10655 29461
rect 552 29402 11132 29424
rect 552 29350 3662 29402
rect 3714 29350 3726 29402
rect 3778 29350 3790 29402
rect 3842 29350 3854 29402
rect 3906 29350 3918 29402
rect 3970 29350 10062 29402
rect 10114 29350 10126 29402
rect 10178 29350 10190 29402
rect 10242 29350 10254 29402
rect 10306 29350 10318 29402
rect 10370 29350 11132 29402
rect 552 29328 11132 29350
rect 1118 29288 1124 29300
rect 768 29260 1124 29288
rect 382 29112 388 29164
rect 440 29112 446 29164
rect 400 28824 428 29112
rect 768 29084 796 29260
rect 1118 29248 1124 29260
rect 1176 29248 1182 29300
rect 1946 29248 1952 29300
rect 2004 29288 2010 29300
rect 2317 29291 2375 29297
rect 2317 29288 2329 29291
rect 2004 29260 2329 29288
rect 2004 29248 2010 29260
rect 2317 29257 2329 29260
rect 2363 29257 2375 29291
rect 2317 29251 2375 29257
rect 5997 29291 6055 29297
rect 5997 29257 6009 29291
rect 6043 29288 6055 29291
rect 6454 29288 6460 29300
rect 6043 29260 6460 29288
rect 6043 29257 6055 29260
rect 5997 29251 6055 29257
rect 6454 29248 6460 29260
rect 6512 29248 6518 29300
rect 6733 29291 6791 29297
rect 6733 29257 6745 29291
rect 6779 29288 6791 29291
rect 6822 29288 6828 29300
rect 6779 29260 6828 29288
rect 6779 29257 6791 29260
rect 6733 29251 6791 29257
rect 6822 29248 6828 29260
rect 6880 29248 6886 29300
rect 6914 29248 6920 29300
rect 6972 29248 6978 29300
rect 7098 29248 7104 29300
rect 7156 29248 7162 29300
rect 7208 29260 7972 29288
rect 845 29223 903 29229
rect 845 29189 857 29223
rect 891 29220 903 29223
rect 1394 29220 1400 29232
rect 891 29192 1400 29220
rect 891 29189 903 29192
rect 845 29183 903 29189
rect 1394 29180 1400 29192
rect 1452 29180 1458 29232
rect 1486 29180 1492 29232
rect 1544 29220 1550 29232
rect 2130 29220 2136 29232
rect 1544 29192 2136 29220
rect 1544 29180 1550 29192
rect 2130 29180 2136 29192
rect 2188 29220 2194 29232
rect 3050 29220 3056 29232
rect 2188 29192 2268 29220
rect 2188 29180 2194 29192
rect 1762 29112 1768 29164
rect 1820 29112 1826 29164
rect 2240 29161 2268 29192
rect 2424 29192 3056 29220
rect 2225 29155 2283 29161
rect 2225 29121 2237 29155
rect 2271 29121 2283 29155
rect 2225 29115 2283 29121
rect 768 29056 980 29084
rect 842 28976 848 29028
rect 900 28976 906 29028
rect 952 29016 980 29056
rect 1026 29044 1032 29096
rect 1084 29044 1090 29096
rect 1118 29044 1124 29096
rect 1176 29044 1182 29096
rect 2041 29087 2099 29093
rect 2041 29053 2053 29087
rect 2087 29084 2099 29087
rect 2424 29084 2452 29192
rect 3050 29180 3056 29192
rect 3108 29180 3114 29232
rect 4614 29180 4620 29232
rect 4672 29220 4678 29232
rect 4709 29223 4767 29229
rect 4709 29220 4721 29223
rect 4672 29192 4721 29220
rect 4672 29180 4678 29192
rect 4709 29189 4721 29192
rect 4755 29189 4767 29223
rect 4709 29183 4767 29189
rect 5074 29180 5080 29232
rect 5132 29180 5138 29232
rect 7116 29220 7144 29248
rect 6104 29192 7144 29220
rect 2516 29124 3004 29152
rect 2516 29093 2544 29124
rect 2087 29056 2452 29084
rect 2501 29087 2559 29093
rect 2087 29053 2099 29056
rect 2041 29047 2099 29053
rect 2501 29053 2513 29087
rect 2547 29053 2559 29087
rect 2761 29087 2819 29093
rect 2761 29084 2773 29087
rect 2501 29047 2559 29053
rect 2608 29056 2773 29084
rect 952 28988 1072 29016
rect 1044 28960 1072 28988
rect 1210 28976 1216 29028
rect 1268 28976 1274 29028
rect 2608 29016 2636 29056
rect 2761 29053 2773 29056
rect 2807 29053 2819 29087
rect 2761 29047 2819 29053
rect 2861 29081 2919 29087
rect 2861 29074 2873 29081
rect 2907 29074 2919 29081
rect 2861 29041 2872 29074
rect 2866 29022 2872 29041
rect 2924 29022 2930 29074
rect 2148 28988 2636 29016
rect 1026 28908 1032 28960
rect 1084 28908 1090 28960
rect 1302 28908 1308 28960
rect 1360 28948 1366 28960
rect 2148 28948 2176 28988
rect 1360 28920 2176 28948
rect 1360 28908 1366 28920
rect 2222 28908 2228 28960
rect 2280 28948 2286 28960
rect 2685 28951 2743 28957
rect 2685 28948 2697 28951
rect 2280 28920 2697 28948
rect 2280 28908 2286 28920
rect 2685 28917 2697 28920
rect 2731 28917 2743 28951
rect 2685 28911 2743 28917
rect 2866 28908 2872 28960
rect 2924 28908 2930 28960
rect 2976 28948 3004 29124
rect 3142 29112 3148 29164
rect 3200 29152 3206 29164
rect 3200 29124 3266 29152
rect 3200 29112 3206 29124
rect 5626 29112 5632 29164
rect 5684 29152 5690 29164
rect 5684 29124 6040 29152
rect 5684 29112 5690 29124
rect 3053 29087 3111 29093
rect 3053 29053 3065 29087
rect 3099 29084 3111 29087
rect 3789 29087 3847 29093
rect 3099 29056 3280 29084
rect 3099 29053 3111 29056
rect 3053 29047 3111 29053
rect 3252 29028 3280 29056
rect 3789 29053 3801 29087
rect 3835 29084 3847 29087
rect 4062 29084 4068 29096
rect 3835 29056 4068 29084
rect 3835 29053 3847 29056
rect 3789 29047 3847 29053
rect 4062 29044 4068 29056
rect 4120 29084 4126 29096
rect 5353 29087 5411 29093
rect 5353 29084 5365 29087
rect 4120 29056 5365 29084
rect 4120 29044 4126 29056
rect 5353 29053 5365 29056
rect 5399 29084 5411 29087
rect 5534 29084 5540 29096
rect 5399 29056 5540 29084
rect 5399 29053 5411 29056
rect 5353 29047 5411 29053
rect 5534 29044 5540 29056
rect 5592 29044 5598 29096
rect 5810 29044 5816 29096
rect 5868 29044 5874 29096
rect 3234 28976 3240 29028
rect 3292 28976 3298 29028
rect 3326 28976 3332 29028
rect 3384 29016 3390 29028
rect 3421 29019 3479 29025
rect 3421 29016 3433 29019
rect 3384 28988 3433 29016
rect 3384 28976 3390 28988
rect 3421 28985 3433 28988
rect 3467 28985 3479 29019
rect 3421 28979 3479 28985
rect 3697 29019 3755 29025
rect 3697 28985 3709 29019
rect 3743 29016 3755 29019
rect 4157 29019 4215 29025
rect 3743 28988 4108 29016
rect 3743 28985 3755 28988
rect 3697 28979 3755 28985
rect 3878 28948 3884 28960
rect 2976 28920 3884 28948
rect 3878 28908 3884 28920
rect 3936 28908 3942 28960
rect 4080 28948 4108 28988
rect 4157 28985 4169 29019
rect 4203 29016 4215 29019
rect 4525 29019 4583 29025
rect 4203 28988 4476 29016
rect 4203 28985 4215 28988
rect 4157 28979 4215 28985
rect 4338 28948 4344 28960
rect 4080 28920 4344 28948
rect 4338 28908 4344 28920
rect 4396 28908 4402 28960
rect 4448 28948 4476 28988
rect 4525 28985 4537 29019
rect 4571 29016 4583 29019
rect 4571 28988 5028 29016
rect 4571 28985 4583 28988
rect 4525 28979 4583 28985
rect 4798 28948 4804 28960
rect 4448 28920 4804 28948
rect 4798 28908 4804 28920
rect 4856 28908 4862 28960
rect 4890 28908 4896 28960
rect 4948 28908 4954 28960
rect 5000 28948 5028 28988
rect 5442 28976 5448 29028
rect 5500 29016 5506 29028
rect 5629 29019 5687 29025
rect 5629 29016 5641 29019
rect 5500 28988 5641 29016
rect 5500 28976 5506 28988
rect 5629 28985 5641 28988
rect 5675 28985 5687 29019
rect 5629 28979 5687 28985
rect 5074 28948 5080 28960
rect 5000 28920 5080 28948
rect 5074 28908 5080 28920
rect 5132 28948 5138 28960
rect 5810 28948 5816 28960
rect 5132 28920 5816 28948
rect 5132 28908 5138 28920
rect 5810 28908 5816 28920
rect 5868 28908 5874 28960
rect 6012 28948 6040 29124
rect 6104 29093 6132 29192
rect 7208 29152 7236 29260
rect 7282 29180 7288 29232
rect 7340 29220 7346 29232
rect 7340 29192 7880 29220
rect 7340 29180 7346 29192
rect 6840 29124 7236 29152
rect 6089 29087 6147 29093
rect 6089 29053 6101 29087
rect 6135 29053 6147 29087
rect 6089 29047 6147 29053
rect 6178 29044 6184 29096
rect 6236 29084 6242 29096
rect 6365 29087 6423 29093
rect 6365 29084 6377 29087
rect 6236 29056 6377 29084
rect 6236 29044 6242 29056
rect 6365 29053 6377 29056
rect 6411 29053 6423 29087
rect 6365 29047 6423 29053
rect 6549 29087 6607 29093
rect 6549 29053 6561 29087
rect 6595 29084 6607 29087
rect 6730 29084 6736 29096
rect 6595 29056 6736 29084
rect 6595 29053 6607 29056
rect 6549 29047 6607 29053
rect 6730 29044 6736 29056
rect 6788 29044 6794 29096
rect 6840 29093 6868 29124
rect 6825 29087 6883 29093
rect 6825 29053 6837 29087
rect 6871 29053 6883 29087
rect 6825 29047 6883 29053
rect 7098 29044 7104 29096
rect 7156 29044 7162 29096
rect 7190 29044 7196 29096
rect 7248 29084 7254 29096
rect 7852 29093 7880 29192
rect 7285 29087 7343 29093
rect 7285 29084 7297 29087
rect 7248 29056 7297 29084
rect 7248 29044 7254 29056
rect 7285 29053 7297 29056
rect 7331 29053 7343 29087
rect 7285 29047 7343 29053
rect 7377 29087 7435 29093
rect 7377 29053 7389 29087
rect 7423 29084 7435 29087
rect 7837 29087 7895 29093
rect 7423 29056 7457 29084
rect 7423 29053 7435 29056
rect 7377 29047 7435 29053
rect 7837 29053 7849 29087
rect 7883 29053 7895 29087
rect 7944 29084 7972 29260
rect 8202 29248 8208 29300
rect 8260 29288 8266 29300
rect 8260 29260 8800 29288
rect 8260 29248 8266 29260
rect 8113 29223 8171 29229
rect 8113 29189 8125 29223
rect 8159 29220 8171 29223
rect 8386 29220 8392 29232
rect 8159 29192 8392 29220
rect 8159 29189 8171 29192
rect 8113 29183 8171 29189
rect 8386 29180 8392 29192
rect 8444 29180 8450 29232
rect 8570 29180 8576 29232
rect 8628 29220 8634 29232
rect 8772 29229 8800 29260
rect 9122 29248 9128 29300
rect 9180 29248 9186 29300
rect 9582 29288 9588 29300
rect 9416 29260 9588 29288
rect 8665 29223 8723 29229
rect 8665 29220 8677 29223
rect 8628 29192 8677 29220
rect 8628 29180 8634 29192
rect 8665 29189 8677 29192
rect 8711 29189 8723 29223
rect 8665 29183 8723 29189
rect 8757 29223 8815 29229
rect 8757 29189 8769 29223
rect 8803 29189 8815 29223
rect 8757 29183 8815 29189
rect 8018 29112 8024 29164
rect 8076 29152 8082 29164
rect 9416 29161 9444 29260
rect 9582 29248 9588 29260
rect 9640 29248 9646 29300
rect 9401 29155 9459 29161
rect 8076 29124 8248 29152
rect 8076 29112 8082 29124
rect 8220 29093 8248 29124
rect 8404 29124 8892 29152
rect 8205 29087 8263 29093
rect 7944 29056 8156 29084
rect 7837 29047 7895 29053
rect 6454 29016 6460 29028
rect 6288 28988 6460 29016
rect 6178 28948 6184 28960
rect 6012 28920 6184 28948
rect 6178 28908 6184 28920
rect 6236 28908 6242 28960
rect 6288 28957 6316 28988
rect 6454 28976 6460 28988
rect 6512 28976 6518 29028
rect 7392 29016 7420 29047
rect 6564 28988 7696 29016
rect 6564 28957 6592 28988
rect 6273 28951 6331 28957
rect 6273 28917 6285 28951
rect 6319 28948 6331 28951
rect 6549 28951 6607 28957
rect 6319 28920 6353 28948
rect 6319 28917 6331 28920
rect 6273 28911 6331 28917
rect 6549 28917 6561 28951
rect 6595 28917 6607 28951
rect 7668 28948 7696 28988
rect 7742 28976 7748 29028
rect 7800 28976 7806 29028
rect 7929 29019 7987 29025
rect 7929 28985 7941 29019
rect 7975 29016 7987 29019
rect 8018 29016 8024 29028
rect 7975 28988 8024 29016
rect 7975 28985 7987 28988
rect 7929 28979 7987 28985
rect 8018 28976 8024 28988
rect 8076 28976 8082 29028
rect 8128 29016 8156 29056
rect 8205 29053 8217 29087
rect 8251 29053 8263 29087
rect 8205 29047 8263 29053
rect 8404 29028 8432 29124
rect 8481 29087 8539 29093
rect 8481 29053 8493 29087
rect 8527 29084 8539 29087
rect 8570 29084 8576 29096
rect 8527 29056 8576 29084
rect 8527 29053 8539 29056
rect 8481 29047 8539 29053
rect 8570 29044 8576 29056
rect 8628 29084 8634 29096
rect 8754 29084 8760 29096
rect 8628 29056 8760 29084
rect 8628 29044 8634 29056
rect 8754 29044 8760 29056
rect 8812 29044 8818 29096
rect 8864 29084 8892 29124
rect 9401 29121 9413 29155
rect 9447 29121 9459 29155
rect 9401 29115 9459 29121
rect 8864 29056 10824 29084
rect 8386 29016 8392 29028
rect 8128 28988 8392 29016
rect 8386 28976 8392 28988
rect 8444 28976 8450 29028
rect 9214 29016 9220 29028
rect 8496 28988 9220 29016
rect 8496 28948 8524 28988
rect 9214 28976 9220 28988
rect 9272 28976 9278 29028
rect 9646 29019 9704 29025
rect 9646 29016 9658 29019
rect 9324 28988 9658 29016
rect 7668 28920 8524 28948
rect 6549 28911 6607 28917
rect 9122 28908 9128 28960
rect 9180 28908 9186 28960
rect 9324 28957 9352 28988
rect 9646 28985 9658 28988
rect 9692 28985 9704 29019
rect 9646 28979 9704 28985
rect 9309 28951 9367 28957
rect 9309 28917 9321 28951
rect 9355 28917 9367 28951
rect 9309 28911 9367 28917
rect 10134 28908 10140 28960
rect 10192 28948 10198 28960
rect 10686 28948 10692 28960
rect 10192 28920 10692 28948
rect 10192 28908 10198 28920
rect 10686 28908 10692 28920
rect 10744 28908 10750 28960
rect 10796 28957 10824 29056
rect 10781 28951 10839 28957
rect 10781 28917 10793 28951
rect 10827 28948 10839 28951
rect 10827 28920 11192 28948
rect 10827 28917 10839 28920
rect 10781 28911 10839 28917
rect 552 28858 11132 28880
rect 382 28772 388 28824
rect 440 28772 446 28824
rect 552 28806 4322 28858
rect 4374 28806 4386 28858
rect 4438 28806 4450 28858
rect 4502 28806 4514 28858
rect 4566 28806 4578 28858
rect 4630 28806 10722 28858
rect 10774 28806 10786 28858
rect 10838 28806 10850 28858
rect 10902 28806 10914 28858
rect 10966 28806 10978 28858
rect 11030 28806 11132 28858
rect 552 28784 11132 28806
rect 1029 28747 1087 28753
rect 1029 28744 1041 28747
rect 32 28716 1041 28744
rect 32 28540 60 28716
rect 1029 28713 1041 28716
rect 1075 28744 1087 28747
rect 1946 28744 1952 28756
rect 1075 28716 1952 28744
rect 1075 28713 1087 28716
rect 1029 28707 1087 28713
rect 1946 28704 1952 28716
rect 2004 28704 2010 28756
rect 2222 28704 2228 28756
rect 2280 28704 2286 28756
rect 2958 28704 2964 28756
rect 3016 28744 3022 28756
rect 3016 28716 3280 28744
rect 3016 28704 3022 28716
rect 106 28636 112 28688
rect 164 28676 170 28688
rect 1213 28679 1271 28685
rect 1213 28676 1225 28679
rect 164 28648 1225 28676
rect 164 28636 170 28648
rect 1213 28645 1225 28648
rect 1259 28676 1271 28679
rect 1302 28676 1308 28688
rect 1259 28648 1308 28676
rect 1259 28645 1271 28648
rect 1213 28639 1271 28645
rect 1302 28636 1308 28648
rect 1360 28636 1366 28688
rect 2240 28676 2268 28704
rect 3252 28676 3280 28716
rect 3326 28704 3332 28756
rect 3384 28744 3390 28756
rect 3421 28747 3479 28753
rect 3421 28744 3433 28747
rect 3384 28716 3433 28744
rect 3384 28704 3390 28716
rect 3421 28713 3433 28716
rect 3467 28713 3479 28747
rect 3421 28707 3479 28713
rect 4062 28704 4068 28756
rect 4120 28744 4126 28756
rect 5169 28747 5227 28753
rect 5169 28744 5181 28747
rect 4120 28716 5181 28744
rect 4120 28704 4126 28716
rect 5169 28713 5181 28716
rect 5215 28713 5227 28747
rect 5169 28707 5227 28713
rect 6089 28747 6147 28753
rect 6089 28713 6101 28747
rect 6135 28744 6147 28747
rect 6270 28744 6276 28756
rect 6135 28716 6276 28744
rect 6135 28713 6147 28716
rect 6089 28707 6147 28713
rect 6270 28704 6276 28716
rect 6328 28704 6334 28756
rect 6914 28704 6920 28756
rect 6972 28744 6978 28756
rect 7653 28747 7711 28753
rect 7653 28744 7665 28747
rect 6972 28716 7665 28744
rect 6972 28704 6978 28716
rect 7653 28713 7665 28716
rect 7699 28713 7711 28747
rect 7653 28707 7711 28713
rect 8573 28747 8631 28753
rect 8573 28713 8585 28747
rect 8619 28744 8631 28747
rect 9122 28744 9128 28756
rect 8619 28716 9128 28744
rect 8619 28713 8631 28716
rect 8573 28707 8631 28713
rect 9122 28704 9128 28716
rect 9180 28704 9186 28756
rect 10071 28747 10129 28753
rect 9232 28716 9996 28744
rect 4890 28676 4896 28688
rect 1504 28648 1992 28676
rect 2240 28648 2452 28676
rect 842 28568 848 28620
rect 900 28568 906 28620
rect 1121 28611 1179 28617
rect 1121 28577 1133 28611
rect 1167 28608 1179 28611
rect 1504 28608 1532 28648
rect 1964 28620 1992 28648
rect 1167 28580 1532 28608
rect 1167 28577 1179 28580
rect 1121 28571 1179 28577
rect 1946 28568 1952 28620
rect 2004 28568 2010 28620
rect 2041 28611 2099 28617
rect 2041 28577 2053 28611
rect 2087 28577 2099 28611
rect 2041 28571 2099 28577
rect 106 28540 112 28552
rect 32 28512 112 28540
rect 106 28500 112 28512
rect 164 28500 170 28552
rect 1762 28500 1768 28552
rect 1820 28500 1826 28552
rect 934 28432 940 28484
rect 992 28472 998 28484
rect 1578 28472 1584 28484
rect 992 28444 1584 28472
rect 992 28432 998 28444
rect 1578 28432 1584 28444
rect 1636 28432 1642 28484
rect 845 28407 903 28413
rect 845 28373 857 28407
rect 891 28404 903 28407
rect 1302 28404 1308 28416
rect 891 28376 1308 28404
rect 891 28373 903 28376
rect 845 28367 903 28373
rect 1302 28364 1308 28376
rect 1360 28364 1366 28416
rect 2056 28404 2084 28571
rect 2130 28568 2136 28620
rect 2188 28608 2194 28620
rect 2225 28611 2283 28617
rect 2225 28608 2237 28611
rect 2188 28580 2237 28608
rect 2188 28568 2194 28580
rect 2225 28577 2237 28580
rect 2271 28577 2283 28611
rect 2225 28571 2283 28577
rect 2317 28611 2375 28617
rect 2317 28577 2329 28611
rect 2363 28577 2375 28611
rect 2317 28571 2375 28577
rect 2130 28432 2136 28484
rect 2188 28472 2194 28484
rect 2332 28472 2360 28571
rect 2424 28540 2452 28648
rect 2516 28648 3004 28676
rect 3252 28648 3455 28676
rect 2516 28617 2544 28648
rect 2501 28611 2559 28617
rect 2501 28577 2513 28611
rect 2547 28577 2559 28611
rect 2501 28571 2559 28577
rect 2593 28611 2651 28617
rect 2593 28577 2605 28611
rect 2639 28577 2651 28611
rect 2593 28571 2651 28577
rect 2777 28611 2835 28617
rect 2777 28577 2789 28611
rect 2823 28577 2835 28611
rect 2777 28571 2835 28577
rect 2608 28540 2636 28571
rect 2792 28540 2820 28571
rect 2866 28568 2872 28620
rect 2924 28568 2930 28620
rect 2976 28617 3004 28648
rect 2961 28611 3019 28617
rect 2961 28577 2973 28611
rect 3007 28608 3019 28611
rect 3326 28608 3332 28620
rect 3007 28580 3332 28608
rect 3007 28577 3019 28580
rect 2961 28571 3019 28577
rect 3326 28568 3332 28580
rect 3384 28568 3390 28620
rect 2424 28512 2636 28540
rect 2700 28512 2820 28540
rect 2188 28444 2360 28472
rect 2188 28432 2194 28444
rect 2222 28404 2228 28416
rect 2056 28376 2228 28404
rect 2222 28364 2228 28376
rect 2280 28364 2286 28416
rect 2406 28364 2412 28416
rect 2464 28364 2470 28416
rect 2700 28404 2728 28512
rect 3234 28500 3240 28552
rect 3292 28540 3298 28552
rect 3427 28540 3455 28648
rect 3896 28648 4896 28676
rect 3602 28568 3608 28620
rect 3660 28568 3666 28620
rect 3896 28617 3924 28648
rect 4890 28636 4896 28648
rect 4948 28676 4954 28688
rect 5353 28679 5411 28685
rect 5353 28676 5365 28679
rect 4948 28648 5365 28676
rect 4948 28636 4954 28648
rect 5353 28645 5365 28648
rect 5399 28645 5411 28679
rect 5810 28676 5816 28688
rect 5353 28639 5411 28645
rect 5644 28648 5816 28676
rect 3881 28611 3939 28617
rect 3881 28577 3893 28611
rect 3927 28577 3939 28611
rect 3881 28571 3939 28577
rect 4157 28611 4215 28617
rect 4157 28577 4169 28611
rect 4203 28608 4215 28611
rect 4246 28608 4252 28620
rect 4203 28580 4252 28608
rect 4203 28577 4215 28580
rect 4157 28571 4215 28577
rect 4246 28568 4252 28580
rect 4304 28568 4310 28620
rect 4614 28568 4620 28620
rect 4672 28568 4678 28620
rect 5077 28611 5135 28617
rect 5077 28577 5089 28611
rect 5123 28577 5135 28611
rect 5077 28571 5135 28577
rect 3292 28512 3455 28540
rect 4264 28540 4292 28568
rect 4264 28512 4384 28540
rect 3292 28500 3298 28512
rect 2774 28432 2780 28484
rect 2832 28472 2838 28484
rect 3697 28475 3755 28481
rect 3697 28472 3709 28475
rect 2832 28444 3709 28472
rect 2832 28432 2838 28444
rect 3697 28441 3709 28444
rect 3743 28441 3755 28475
rect 3697 28435 3755 28441
rect 4246 28432 4252 28484
rect 4304 28432 4310 28484
rect 4356 28472 4384 28512
rect 4430 28500 4436 28552
rect 4488 28540 4494 28552
rect 4709 28543 4767 28549
rect 4709 28540 4721 28543
rect 4488 28512 4721 28540
rect 4488 28500 4494 28512
rect 4709 28509 4721 28512
rect 4755 28509 4767 28543
rect 4709 28503 4767 28509
rect 4893 28543 4951 28549
rect 4893 28509 4905 28543
rect 4939 28540 4951 28543
rect 4982 28540 4988 28552
rect 4939 28512 4988 28540
rect 4939 28509 4951 28512
rect 4893 28503 4951 28509
rect 4982 28500 4988 28512
rect 5040 28500 5046 28552
rect 5092 28472 5120 28571
rect 5442 28568 5448 28620
rect 5500 28568 5506 28620
rect 5644 28617 5672 28648
rect 5810 28636 5816 28648
rect 5868 28636 5874 28688
rect 6288 28648 7144 28676
rect 5629 28611 5687 28617
rect 5629 28577 5641 28611
rect 5675 28577 5687 28611
rect 6288 28608 6316 28648
rect 5629 28571 5687 28577
rect 5736 28580 6316 28608
rect 5736 28540 5764 28580
rect 6362 28568 6368 28620
rect 6420 28568 6426 28620
rect 6454 28568 6460 28620
rect 6512 28568 6518 28620
rect 6546 28568 6552 28620
rect 6604 28608 6610 28620
rect 6825 28611 6883 28617
rect 6825 28608 6837 28611
rect 6604 28580 6837 28608
rect 6604 28568 6610 28580
rect 6825 28577 6837 28580
rect 6871 28577 6883 28611
rect 7006 28606 7012 28620
rect 6825 28571 6883 28577
rect 6932 28578 7012 28606
rect 4356 28444 5120 28472
rect 5368 28512 5764 28540
rect 6932 28526 6960 28578
rect 7006 28568 7012 28578
rect 7064 28568 7070 28620
rect 7116 28608 7144 28648
rect 7190 28636 7196 28688
rect 7248 28636 7254 28688
rect 9232 28676 9260 28716
rect 8220 28648 9260 28676
rect 8220 28620 8248 28648
rect 9398 28636 9404 28688
rect 9456 28636 9462 28688
rect 9490 28636 9496 28688
rect 9548 28676 9554 28688
rect 9861 28679 9919 28685
rect 9861 28676 9873 28679
rect 9548 28648 9873 28676
rect 9548 28636 9554 28648
rect 9861 28645 9873 28648
rect 9907 28645 9919 28679
rect 9968 28676 9996 28716
rect 10071 28713 10083 28747
rect 10117 28744 10129 28747
rect 10117 28716 10640 28744
rect 10117 28713 10129 28716
rect 10071 28707 10129 28713
rect 9968 28648 10548 28676
rect 9861 28639 9919 28645
rect 7561 28611 7619 28617
rect 7561 28608 7573 28611
rect 7116 28580 7573 28608
rect 7561 28577 7573 28580
rect 7607 28577 7619 28611
rect 7561 28571 7619 28577
rect 7650 28568 7656 28620
rect 7708 28608 7714 28620
rect 7745 28611 7803 28617
rect 7745 28608 7757 28611
rect 7708 28580 7757 28608
rect 7708 28568 7714 28580
rect 7745 28577 7757 28580
rect 7791 28577 7803 28611
rect 7745 28571 7803 28577
rect 8113 28611 8171 28617
rect 8113 28577 8125 28611
rect 8159 28577 8171 28611
rect 8113 28571 8171 28577
rect 2958 28404 2964 28416
rect 2700 28376 2964 28404
rect 2958 28364 2964 28376
rect 3016 28364 3022 28416
rect 3237 28407 3295 28413
rect 3237 28373 3249 28407
rect 3283 28404 3295 28407
rect 3602 28404 3608 28416
rect 3283 28376 3608 28404
rect 3283 28373 3295 28376
rect 3237 28367 3295 28373
rect 3602 28364 3608 28376
rect 3660 28364 3666 28416
rect 3878 28364 3884 28416
rect 3936 28404 3942 28416
rect 4338 28404 4344 28416
rect 3936 28376 4344 28404
rect 3936 28364 3942 28376
rect 4338 28364 4344 28376
rect 4396 28364 4402 28416
rect 4522 28364 4528 28416
rect 4580 28404 4586 28416
rect 5368 28413 5396 28512
rect 5353 28407 5411 28413
rect 5353 28404 5365 28407
rect 4580 28376 5365 28404
rect 4580 28364 4586 28376
rect 5353 28373 5365 28376
rect 5399 28373 5411 28407
rect 5353 28367 5411 28373
rect 5442 28364 5448 28416
rect 5500 28404 5506 28416
rect 5537 28407 5595 28413
rect 5537 28404 5549 28407
rect 5500 28376 5549 28404
rect 5500 28364 5506 28376
rect 5537 28373 5549 28376
rect 5583 28373 5595 28407
rect 5537 28367 5595 28373
rect 7374 28364 7380 28416
rect 7432 28364 7438 28416
rect 7650 28364 7656 28416
rect 7708 28404 7714 28416
rect 7929 28407 7987 28413
rect 7929 28404 7941 28407
rect 7708 28376 7941 28404
rect 7708 28364 7714 28376
rect 7929 28373 7941 28376
rect 7975 28373 7987 28407
rect 8128 28404 8156 28571
rect 8202 28568 8208 28620
rect 8260 28568 8266 28620
rect 8386 28568 8392 28620
rect 8444 28568 8450 28620
rect 8570 28568 8576 28620
rect 8628 28608 8634 28620
rect 8849 28611 8907 28617
rect 8849 28608 8861 28611
rect 8628 28580 8861 28608
rect 8628 28568 8634 28580
rect 8849 28577 8861 28580
rect 8895 28577 8907 28611
rect 8849 28571 8907 28577
rect 8864 28540 8892 28571
rect 8938 28568 8944 28620
rect 8996 28568 9002 28620
rect 9033 28611 9091 28617
rect 9033 28577 9045 28611
rect 9079 28608 9091 28611
rect 9122 28608 9128 28620
rect 9079 28580 9128 28608
rect 9079 28577 9091 28580
rect 9033 28571 9091 28577
rect 9122 28568 9128 28580
rect 9180 28568 9186 28620
rect 9217 28611 9275 28617
rect 9217 28577 9229 28611
rect 9263 28608 9275 28611
rect 9950 28608 9956 28620
rect 9263 28580 9956 28608
rect 9263 28577 9275 28580
rect 9217 28571 9275 28577
rect 9950 28568 9956 28580
rect 10008 28608 10014 28620
rect 10410 28608 10416 28620
rect 10008 28580 10416 28608
rect 10008 28568 10014 28580
rect 10410 28568 10416 28580
rect 10468 28568 10474 28620
rect 10520 28617 10548 28648
rect 10505 28611 10563 28617
rect 10505 28577 10517 28611
rect 10551 28577 10563 28611
rect 10505 28571 10563 28577
rect 9306 28540 9312 28552
rect 8864 28512 9312 28540
rect 9306 28500 9312 28512
rect 9364 28500 9370 28552
rect 9398 28500 9404 28552
rect 9456 28540 9462 28552
rect 10321 28543 10379 28549
rect 10321 28540 10333 28543
rect 9456 28512 10333 28540
rect 9456 28500 9462 28512
rect 10321 28509 10333 28512
rect 10367 28509 10379 28543
rect 10612 28540 10640 28716
rect 10689 28611 10747 28617
rect 10689 28577 10701 28611
rect 10735 28608 10747 28611
rect 11164 28608 11192 28920
rect 10735 28580 11192 28608
rect 10735 28577 10747 28580
rect 10689 28571 10747 28577
rect 11330 28540 11336 28552
rect 10612 28512 11336 28540
rect 10321 28503 10379 28509
rect 11330 28500 11336 28512
rect 11388 28500 11394 28552
rect 8294 28432 8300 28484
rect 8352 28472 8358 28484
rect 8665 28475 8723 28481
rect 8665 28472 8677 28475
rect 8352 28444 8677 28472
rect 8352 28432 8358 28444
rect 8665 28441 8677 28444
rect 8711 28441 8723 28475
rect 8665 28435 8723 28441
rect 8754 28432 8760 28484
rect 8812 28472 8818 28484
rect 10229 28475 10287 28481
rect 8812 28444 10114 28472
rect 8812 28432 8818 28444
rect 9306 28404 9312 28416
rect 8128 28376 9312 28404
rect 7929 28367 7987 28373
rect 9306 28364 9312 28376
rect 9364 28364 9370 28416
rect 9490 28364 9496 28416
rect 9548 28364 9554 28416
rect 10086 28413 10114 28444
rect 10229 28441 10241 28475
rect 10275 28472 10287 28475
rect 10502 28472 10508 28484
rect 10275 28444 10508 28472
rect 10275 28441 10287 28444
rect 10229 28435 10287 28441
rect 10502 28432 10508 28444
rect 10560 28432 10566 28484
rect 10067 28407 10125 28413
rect 10067 28373 10079 28407
rect 10113 28373 10125 28407
rect 10067 28367 10125 28373
rect 552 28314 11132 28336
rect 552 28262 3662 28314
rect 3714 28262 3726 28314
rect 3778 28262 3790 28314
rect 3842 28262 3854 28314
rect 3906 28262 3918 28314
rect 3970 28262 10062 28314
rect 10114 28262 10126 28314
rect 10178 28262 10190 28314
rect 10242 28262 10254 28314
rect 10306 28262 10318 28314
rect 10370 28262 11132 28314
rect 552 28240 11132 28262
rect 1854 28160 1860 28212
rect 1912 28200 1918 28212
rect 1912 28172 2728 28200
rect 1912 28160 1918 28172
rect 842 28092 848 28144
rect 900 28132 906 28144
rect 2700 28132 2728 28172
rect 3050 28160 3056 28212
rect 3108 28160 3114 28212
rect 3142 28160 3148 28212
rect 3200 28200 3206 28212
rect 3237 28203 3295 28209
rect 3237 28200 3249 28203
rect 3200 28172 3249 28200
rect 3200 28160 3206 28172
rect 3237 28169 3249 28172
rect 3283 28169 3295 28203
rect 3237 28163 3295 28169
rect 3602 28160 3608 28212
rect 3660 28160 3666 28212
rect 3878 28160 3884 28212
rect 3936 28200 3942 28212
rect 4157 28203 4215 28209
rect 4157 28200 4169 28203
rect 3936 28172 4169 28200
rect 3936 28160 3942 28172
rect 4157 28169 4169 28172
rect 4203 28169 4215 28203
rect 4157 28163 4215 28169
rect 4430 28160 4436 28212
rect 4488 28160 4494 28212
rect 9490 28160 9496 28212
rect 9548 28200 9554 28212
rect 10134 28200 10140 28212
rect 9548 28172 10140 28200
rect 9548 28160 9554 28172
rect 10134 28160 10140 28172
rect 10192 28160 10198 28212
rect 900 28104 1072 28132
rect 2700 28104 2820 28132
rect 900 28092 906 28104
rect 106 27956 112 28008
rect 164 27996 170 28008
rect 845 27999 903 28005
rect 845 27996 857 27999
rect 164 27968 857 27996
rect 164 27956 170 27968
rect 845 27965 857 27968
rect 891 27965 903 27999
rect 845 27959 903 27965
rect 1044 27928 1072 28104
rect 1213 28067 1271 28073
rect 1213 28033 1225 28067
rect 1259 28064 1271 28067
rect 1486 28064 1492 28076
rect 1259 28036 1492 28064
rect 1259 28033 1271 28036
rect 1213 28027 1271 28033
rect 1486 28024 1492 28036
rect 1544 28024 1550 28076
rect 2222 28024 2228 28076
rect 2280 28064 2286 28076
rect 2280 28036 2452 28064
rect 2280 28024 2286 28036
rect 1118 27956 1124 28008
rect 1176 27956 1182 28008
rect 1394 27956 1400 28008
rect 1452 27956 1458 28008
rect 1673 27999 1731 28005
rect 1673 27965 1685 27999
rect 1719 27996 1731 27999
rect 1854 27996 1860 28008
rect 1719 27968 1860 27996
rect 1719 27965 1731 27968
rect 1673 27959 1731 27965
rect 1854 27956 1860 27968
rect 1912 27996 1918 28008
rect 2317 27999 2375 28005
rect 2317 27996 2329 27999
rect 1912 27968 2329 27996
rect 1912 27956 1918 27968
rect 2317 27965 2329 27968
rect 2363 27965 2375 27999
rect 2317 27959 2375 27965
rect 1044 27900 1256 27928
rect 842 27820 848 27872
rect 900 27860 906 27872
rect 1029 27863 1087 27869
rect 1029 27860 1041 27863
rect 900 27832 1041 27860
rect 900 27820 906 27832
rect 1029 27829 1041 27832
rect 1075 27829 1087 27863
rect 1228 27860 1256 27900
rect 1578 27888 1584 27940
rect 1636 27928 1642 27940
rect 2225 27931 2283 27937
rect 2225 27928 2237 27931
rect 1636 27900 2237 27928
rect 1636 27888 1642 27900
rect 2225 27897 2237 27900
rect 2271 27897 2283 27931
rect 2225 27891 2283 27897
rect 2130 27860 2136 27872
rect 1228 27832 2136 27860
rect 1029 27823 1087 27829
rect 2130 27820 2136 27832
rect 2188 27820 2194 27872
rect 2424 27860 2452 28036
rect 2590 28024 2596 28076
rect 2648 28024 2654 28076
rect 2792 28073 2820 28104
rect 2685 28067 2743 28073
rect 2685 28033 2697 28067
rect 2731 28033 2743 28067
rect 2685 28027 2743 28033
rect 2777 28067 2835 28073
rect 2777 28033 2789 28067
rect 2823 28033 2835 28067
rect 3068 28064 3096 28160
rect 4062 28132 4068 28144
rect 3344 28104 4068 28132
rect 3142 28064 3148 28076
rect 3068 28036 3148 28064
rect 2777 28027 2835 28033
rect 2501 27999 2559 28005
rect 2501 27965 2513 27999
rect 2547 27996 2559 27999
rect 2608 27996 2636 28024
rect 2547 27968 2636 27996
rect 2547 27965 2559 27968
rect 2501 27959 2559 27965
rect 2700 27940 2728 28027
rect 3142 28024 3148 28036
rect 3200 28024 3206 28076
rect 2869 27999 2927 28005
rect 2869 27965 2881 27999
rect 2915 27965 2927 27999
rect 2869 27959 2927 27965
rect 3053 27999 3111 28005
rect 3053 27965 3065 27999
rect 3099 27996 3111 27999
rect 3344 27996 3372 28104
rect 4062 28092 4068 28104
rect 4120 28132 4126 28144
rect 4448 28132 4476 28160
rect 4120 28104 4476 28132
rect 5905 28135 5963 28141
rect 4120 28092 4126 28104
rect 5905 28101 5917 28135
rect 5951 28132 5963 28135
rect 6178 28132 6184 28144
rect 5951 28104 6184 28132
rect 5951 28101 5963 28104
rect 5905 28095 5963 28101
rect 6178 28092 6184 28104
rect 6236 28092 6242 28144
rect 8021 28135 8079 28141
rect 8021 28101 8033 28135
rect 8067 28132 8079 28135
rect 8202 28132 8208 28144
rect 8067 28104 8208 28132
rect 8067 28101 8079 28104
rect 8021 28095 8079 28101
rect 8202 28092 8208 28104
rect 8260 28132 8266 28144
rect 11054 28132 11060 28144
rect 8260 28104 8340 28132
rect 8260 28092 8266 28104
rect 3694 28024 3700 28076
rect 3752 28024 3758 28076
rect 3786 28024 3792 28076
rect 3844 28024 3850 28076
rect 4798 28024 4804 28076
rect 4856 28024 4862 28076
rect 7006 28024 7012 28076
rect 7064 28024 7070 28076
rect 3099 27968 3372 27996
rect 3421 27999 3479 28005
rect 3099 27965 3111 27968
rect 3053 27959 3111 27965
rect 3421 27965 3433 27999
rect 3467 27996 3479 27999
rect 3510 27996 3516 28008
rect 3467 27968 3516 27996
rect 3467 27965 3479 27968
rect 3421 27959 3479 27965
rect 2682 27888 2688 27940
rect 2740 27888 2746 27940
rect 2774 27860 2780 27872
rect 2424 27832 2780 27860
rect 2774 27820 2780 27832
rect 2832 27820 2838 27872
rect 2884 27860 2912 27959
rect 3510 27956 3516 27968
rect 3568 27996 3574 28008
rect 3973 27999 4031 28005
rect 3973 27996 3985 27999
rect 3568 27968 3985 27996
rect 3568 27956 3574 27968
rect 3973 27965 3985 27968
rect 4019 27965 4031 27999
rect 3973 27959 4031 27965
rect 4249 27999 4307 28005
rect 4249 27965 4261 27999
rect 4295 27996 4307 27999
rect 4338 27996 4344 28008
rect 4295 27968 4344 27996
rect 4295 27965 4307 27968
rect 4249 27959 4307 27965
rect 4338 27956 4344 27968
rect 4396 27996 4402 28008
rect 4706 27996 4712 28008
rect 4396 27968 4712 27996
rect 4396 27956 4402 27968
rect 4706 27956 4712 27968
rect 4764 27956 4770 28008
rect 4890 27956 4896 28008
rect 4948 27956 4954 28008
rect 4985 27999 5043 28005
rect 4985 27965 4997 27999
rect 5031 27996 5043 27999
rect 6178 27996 6184 28008
rect 5031 27968 5672 27996
rect 5031 27965 5043 27968
rect 4985 27959 5043 27965
rect 5644 27940 5672 27968
rect 5828 27968 6184 27996
rect 2961 27931 3019 27937
rect 2961 27897 2973 27931
rect 3007 27928 3019 27931
rect 4798 27928 4804 27940
rect 3007 27900 4804 27928
rect 3007 27897 3019 27900
rect 2961 27891 3019 27897
rect 4798 27888 4804 27900
rect 4856 27888 4862 27940
rect 5353 27931 5411 27937
rect 5353 27897 5365 27931
rect 5399 27897 5411 27931
rect 5353 27891 5411 27897
rect 4522 27860 4528 27872
rect 2884 27832 4528 27860
rect 4522 27820 4528 27832
rect 4580 27820 4586 27872
rect 4617 27863 4675 27869
rect 4617 27829 4629 27863
rect 4663 27860 4675 27863
rect 5074 27860 5080 27872
rect 4663 27832 5080 27860
rect 4663 27829 4675 27832
rect 4617 27823 4675 27829
rect 5074 27820 5080 27832
rect 5132 27820 5138 27872
rect 5368 27860 5396 27891
rect 5626 27888 5632 27940
rect 5684 27888 5690 27940
rect 5721 27931 5779 27937
rect 5721 27897 5733 27931
rect 5767 27928 5779 27931
rect 5828 27928 5856 27968
rect 6178 27956 6184 27968
rect 6236 27996 6242 28008
rect 6236 27968 6390 27996
rect 6236 27956 6242 27968
rect 5767 27900 5856 27928
rect 5767 27897 5779 27900
rect 5721 27891 5779 27897
rect 5994 27888 6000 27940
rect 6052 27928 6058 27940
rect 6273 27931 6331 27937
rect 6273 27928 6285 27931
rect 6052 27900 6285 27928
rect 6052 27888 6058 27900
rect 6273 27897 6285 27900
rect 6319 27897 6331 27931
rect 6273 27891 6331 27897
rect 5902 27860 5908 27872
rect 5368 27832 5908 27860
rect 5902 27820 5908 27832
rect 5960 27820 5966 27872
rect 6362 27860 6390 27968
rect 6546 27956 6552 28008
rect 6604 27956 6610 28008
rect 6730 27956 6736 28008
rect 6788 27996 6794 28008
rect 7024 27996 7052 28024
rect 6788 27968 7052 27996
rect 6788 27956 6794 27968
rect 8202 27956 8208 28008
rect 8260 27956 8266 28008
rect 8312 27996 8340 28104
rect 8588 28104 11060 28132
rect 8588 28073 8616 28104
rect 11054 28092 11060 28104
rect 11112 28092 11118 28144
rect 8573 28067 8631 28073
rect 8573 28033 8585 28067
rect 8619 28033 8631 28067
rect 8573 28027 8631 28033
rect 8938 28024 8944 28076
rect 8996 28064 9002 28076
rect 9217 28067 9275 28073
rect 9217 28064 9229 28067
rect 8996 28036 9229 28064
rect 8996 28024 9002 28036
rect 9217 28033 9229 28036
rect 9263 28033 9275 28067
rect 9217 28027 9275 28033
rect 9398 28024 9404 28076
rect 9456 28024 9462 28076
rect 9490 28024 9496 28076
rect 9548 28024 9554 28076
rect 9677 28067 9735 28073
rect 9677 28033 9689 28067
rect 9723 28064 9735 28067
rect 9766 28064 9772 28076
rect 9723 28036 9772 28064
rect 9723 28033 9735 28036
rect 9677 28027 9735 28033
rect 9766 28024 9772 28036
rect 9824 28024 9830 28076
rect 9950 28024 9956 28076
rect 10008 28064 10014 28076
rect 10137 28067 10195 28073
rect 10137 28064 10149 28067
rect 10008 28036 10149 28064
rect 10008 28024 10014 28036
rect 10137 28033 10149 28036
rect 10183 28033 10195 28067
rect 10137 28027 10195 28033
rect 10594 28024 10600 28076
rect 10652 28024 10658 28076
rect 9122 27996 9128 28008
rect 8312 27968 9128 27996
rect 9122 27956 9128 27968
rect 9180 27996 9186 28008
rect 9585 27999 9643 28005
rect 9585 27996 9597 27999
rect 9180 27968 9597 27996
rect 9180 27956 9186 27968
rect 9585 27965 9597 27968
rect 9631 27965 9643 27999
rect 9585 27959 9643 27965
rect 10229 27999 10287 28005
rect 10229 27965 10241 27999
rect 10275 27996 10287 27999
rect 10410 27996 10416 28008
rect 10275 27968 10416 27996
rect 10275 27965 10287 27968
rect 10229 27959 10287 27965
rect 10410 27956 10416 27968
rect 10468 27956 10474 28008
rect 6641 27931 6699 27937
rect 6641 27897 6653 27931
rect 6687 27928 6699 27931
rect 6914 27928 6920 27940
rect 6687 27900 6920 27928
rect 6687 27897 6699 27900
rect 6641 27891 6699 27897
rect 6914 27888 6920 27900
rect 6972 27888 6978 27940
rect 7009 27931 7067 27937
rect 7009 27897 7021 27931
rect 7055 27897 7067 27931
rect 7009 27891 7067 27897
rect 7024 27860 7052 27891
rect 7098 27888 7104 27940
rect 7156 27928 7162 27940
rect 7156 27900 7604 27928
rect 7156 27888 7162 27900
rect 6362 27832 7052 27860
rect 7377 27863 7435 27869
rect 7377 27829 7389 27863
rect 7423 27860 7435 27863
rect 7466 27860 7472 27872
rect 7423 27832 7472 27860
rect 7423 27829 7435 27832
rect 7377 27823 7435 27829
rect 7466 27820 7472 27832
rect 7524 27820 7530 27872
rect 7576 27869 7604 27900
rect 8110 27888 8116 27940
rect 8168 27928 8174 27940
rect 8665 27931 8723 27937
rect 8665 27928 8677 27931
rect 8168 27900 8677 27928
rect 8168 27888 8174 27900
rect 8665 27897 8677 27900
rect 8711 27897 8723 27931
rect 8665 27891 8723 27897
rect 9306 27888 9312 27940
rect 9364 27928 9370 27940
rect 9490 27928 9496 27940
rect 9364 27900 9496 27928
rect 9364 27888 9370 27900
rect 9490 27888 9496 27900
rect 9548 27888 9554 27940
rect 9766 27888 9772 27940
rect 9824 27928 9830 27940
rect 10042 27928 10048 27940
rect 9824 27900 10048 27928
rect 9824 27888 9830 27900
rect 10042 27888 10048 27900
rect 10100 27888 10106 27940
rect 7561 27863 7619 27869
rect 7561 27829 7573 27863
rect 7607 27829 7619 27863
rect 7561 27823 7619 27829
rect 8294 27820 8300 27872
rect 8352 27860 8358 27872
rect 8757 27863 8815 27869
rect 8757 27860 8769 27863
rect 8352 27832 8769 27860
rect 8352 27820 8358 27832
rect 8757 27829 8769 27832
rect 8803 27829 8815 27863
rect 8757 27823 8815 27829
rect 9125 27863 9183 27869
rect 9125 27829 9137 27863
rect 9171 27860 9183 27863
rect 9214 27860 9220 27872
rect 9171 27832 9220 27860
rect 9171 27829 9183 27832
rect 9125 27823 9183 27829
rect 9214 27820 9220 27832
rect 9272 27820 9278 27872
rect 552 27770 11132 27792
rect 552 27718 4322 27770
rect 4374 27718 4386 27770
rect 4438 27718 4450 27770
rect 4502 27718 4514 27770
rect 4566 27718 4578 27770
rect 4630 27718 10722 27770
rect 10774 27718 10786 27770
rect 10838 27718 10850 27770
rect 10902 27718 10914 27770
rect 10966 27718 10978 27770
rect 11030 27718 11132 27770
rect 552 27696 11132 27718
rect 1394 27616 1400 27668
rect 1452 27656 1458 27668
rect 1452 27628 1900 27656
rect 1452 27616 1458 27628
rect 1029 27591 1087 27597
rect 1029 27557 1041 27591
rect 1075 27588 1087 27591
rect 1762 27588 1768 27600
rect 1075 27560 1768 27588
rect 1075 27557 1087 27560
rect 1029 27551 1087 27557
rect 1762 27548 1768 27560
rect 1820 27548 1826 27600
rect 1872 27588 1900 27628
rect 1946 27616 1952 27668
rect 2004 27656 2010 27668
rect 2409 27659 2467 27665
rect 2409 27656 2421 27659
rect 2004 27628 2421 27656
rect 2004 27616 2010 27628
rect 2409 27625 2421 27628
rect 2455 27625 2467 27659
rect 3237 27659 3295 27665
rect 3237 27656 3249 27659
rect 2409 27619 2467 27625
rect 2516 27628 3249 27656
rect 2516 27588 2544 27628
rect 3237 27625 3249 27628
rect 3283 27625 3295 27659
rect 3237 27619 3295 27625
rect 4062 27616 4068 27668
rect 4120 27656 4126 27668
rect 5261 27659 5319 27665
rect 5261 27656 5273 27659
rect 4120 27628 5273 27656
rect 4120 27616 4126 27628
rect 5261 27625 5273 27628
rect 5307 27656 5319 27659
rect 5307 27628 5672 27656
rect 5307 27625 5319 27628
rect 5261 27619 5319 27625
rect 1872 27560 2544 27588
rect 2774 27548 2780 27600
rect 2832 27588 2838 27600
rect 3786 27588 3792 27600
rect 2832 27560 3792 27588
rect 2832 27548 2838 27560
rect 3786 27548 3792 27560
rect 3844 27548 3850 27600
rect 4148 27591 4206 27597
rect 4148 27557 4160 27591
rect 4194 27588 4206 27591
rect 4246 27588 4252 27600
rect 4194 27560 4252 27588
rect 4194 27557 4206 27560
rect 4148 27551 4206 27557
rect 4246 27548 4252 27560
rect 4304 27548 4310 27600
rect 4614 27548 4620 27600
rect 4672 27588 4678 27600
rect 4982 27588 4988 27600
rect 4672 27560 4988 27588
rect 4672 27548 4678 27560
rect 4982 27548 4988 27560
rect 5040 27548 5046 27600
rect 5442 27548 5448 27600
rect 5500 27588 5506 27600
rect 5644 27588 5672 27628
rect 5718 27616 5724 27668
rect 5776 27656 5782 27668
rect 8021 27659 8079 27665
rect 8021 27656 8033 27659
rect 5776 27628 8033 27656
rect 5776 27616 5782 27628
rect 8021 27625 8033 27628
rect 8067 27625 8079 27659
rect 8938 27656 8944 27668
rect 8021 27619 8079 27625
rect 8220 27628 8944 27656
rect 5500 27560 5580 27588
rect 5644 27560 5856 27588
rect 5500 27548 5506 27560
rect 14 27480 20 27532
rect 72 27520 78 27532
rect 1213 27523 1271 27529
rect 1213 27520 1225 27523
rect 72 27492 1225 27520
rect 72 27480 78 27492
rect 1213 27489 1225 27492
rect 1259 27520 1271 27523
rect 1259 27492 1716 27520
rect 1259 27489 1271 27492
rect 1213 27483 1271 27489
rect 1305 27455 1363 27461
rect 1305 27421 1317 27455
rect 1351 27452 1363 27455
rect 1578 27452 1584 27464
rect 1351 27424 1584 27452
rect 1351 27421 1363 27424
rect 1305 27415 1363 27421
rect 1578 27412 1584 27424
rect 1636 27412 1642 27464
rect 934 27344 940 27396
rect 992 27384 998 27396
rect 1688 27384 1716 27492
rect 1854 27480 1860 27532
rect 1912 27480 1918 27532
rect 2038 27480 2044 27532
rect 2096 27520 2102 27532
rect 2133 27523 2191 27529
rect 2133 27520 2145 27523
rect 2096 27492 2145 27520
rect 2096 27480 2102 27492
rect 2133 27489 2145 27492
rect 2179 27489 2191 27523
rect 2133 27483 2191 27489
rect 2406 27480 2412 27532
rect 2464 27520 2470 27532
rect 2593 27523 2651 27529
rect 2593 27520 2605 27523
rect 2464 27492 2605 27520
rect 2464 27480 2470 27492
rect 2593 27489 2605 27492
rect 2639 27489 2651 27523
rect 2593 27483 2651 27489
rect 2682 27480 2688 27532
rect 2740 27480 2746 27532
rect 3605 27523 3663 27529
rect 3605 27520 3617 27523
rect 2792 27492 3617 27520
rect 1762 27412 1768 27464
rect 1820 27452 1826 27464
rect 2792 27461 2820 27492
rect 3605 27489 3617 27492
rect 3651 27489 3663 27523
rect 3605 27483 3663 27489
rect 3881 27523 3939 27529
rect 3881 27489 3893 27523
rect 3927 27520 3939 27523
rect 3970 27520 3976 27532
rect 3927 27492 3976 27520
rect 3927 27489 3939 27492
rect 3881 27483 3939 27489
rect 3970 27480 3976 27492
rect 4028 27480 4034 27532
rect 4706 27480 4712 27532
rect 4764 27520 4770 27532
rect 4764 27492 4936 27520
rect 4764 27480 4770 27492
rect 2317 27455 2375 27461
rect 2317 27452 2329 27455
rect 1820 27424 2329 27452
rect 1820 27412 1826 27424
rect 2317 27421 2329 27424
rect 2363 27421 2375 27455
rect 2317 27415 2375 27421
rect 2777 27455 2835 27461
rect 2777 27421 2789 27455
rect 2823 27421 2835 27455
rect 2777 27415 2835 27421
rect 2869 27455 2927 27461
rect 2869 27421 2881 27455
rect 2915 27452 2927 27455
rect 3234 27452 3240 27464
rect 2915 27424 3240 27452
rect 2915 27421 2927 27424
rect 2869 27415 2927 27421
rect 2792 27384 2820 27415
rect 3234 27412 3240 27424
rect 3292 27412 3298 27464
rect 3421 27455 3479 27461
rect 3421 27421 3433 27455
rect 3467 27421 3479 27455
rect 3421 27415 3479 27421
rect 992 27356 1240 27384
rect 992 27344 998 27356
rect 1212 27328 1240 27356
rect 1688 27356 2820 27384
rect 1688 27328 1716 27356
rect 3050 27344 3056 27396
rect 3108 27384 3114 27396
rect 3436 27384 3464 27415
rect 3510 27412 3516 27464
rect 3568 27412 3574 27464
rect 3697 27455 3755 27461
rect 3697 27421 3709 27455
rect 3743 27421 3755 27455
rect 4908 27452 4936 27492
rect 5074 27480 5080 27532
rect 5132 27520 5138 27532
rect 5350 27520 5356 27532
rect 5132 27492 5356 27520
rect 5132 27480 5138 27492
rect 5350 27480 5356 27492
rect 5408 27480 5414 27532
rect 5552 27529 5580 27560
rect 5537 27523 5595 27529
rect 5537 27489 5549 27523
rect 5583 27520 5595 27523
rect 5718 27520 5724 27532
rect 5583 27492 5724 27520
rect 5583 27489 5595 27492
rect 5537 27483 5595 27489
rect 5718 27480 5724 27492
rect 5776 27480 5782 27532
rect 5828 27529 5856 27560
rect 5994 27548 6000 27600
rect 6052 27588 6058 27600
rect 6365 27591 6423 27597
rect 6365 27588 6377 27591
rect 6052 27560 6377 27588
rect 6052 27548 6058 27560
rect 6365 27557 6377 27560
rect 6411 27557 6423 27591
rect 6365 27551 6423 27557
rect 6730 27548 6736 27600
rect 6788 27548 6794 27600
rect 7101 27591 7159 27597
rect 7101 27557 7113 27591
rect 7147 27588 7159 27591
rect 7374 27588 7380 27600
rect 7147 27560 7380 27588
rect 7147 27557 7159 27560
rect 7101 27551 7159 27557
rect 7374 27548 7380 27560
rect 7432 27548 7438 27600
rect 8220 27597 8248 27628
rect 8938 27616 8944 27628
rect 8996 27616 9002 27668
rect 9048 27628 9812 27656
rect 7469 27591 7527 27597
rect 7469 27557 7481 27591
rect 7515 27588 7527 27591
rect 8205 27591 8263 27597
rect 7515 27560 8156 27588
rect 7515 27557 7527 27560
rect 7469 27551 7527 27557
rect 5813 27523 5871 27529
rect 5813 27489 5825 27523
rect 5859 27489 5871 27523
rect 5813 27483 5871 27489
rect 4908 27424 5396 27452
rect 3697 27415 3755 27421
rect 3108 27356 3464 27384
rect 3108 27344 3114 27356
rect 842 27276 848 27328
rect 900 27316 906 27328
rect 1118 27316 1124 27328
rect 900 27288 1124 27316
rect 900 27276 906 27288
rect 1118 27276 1124 27288
rect 1176 27276 1182 27328
rect 1210 27276 1216 27328
rect 1268 27276 1274 27328
rect 1670 27276 1676 27328
rect 1728 27276 1734 27328
rect 2590 27276 2596 27328
rect 2648 27316 2654 27328
rect 2774 27316 2780 27328
rect 2648 27288 2780 27316
rect 2648 27276 2654 27288
rect 2774 27276 2780 27288
rect 2832 27276 2838 27328
rect 3234 27276 3240 27328
rect 3292 27316 3298 27328
rect 3712 27316 3740 27415
rect 5368 27396 5396 27424
rect 5442 27412 5448 27464
rect 5500 27452 5506 27464
rect 5828 27452 5856 27483
rect 6270 27480 6276 27532
rect 6328 27520 6334 27532
rect 6641 27523 6699 27529
rect 6641 27520 6653 27523
rect 6328 27492 6653 27520
rect 6328 27480 6334 27492
rect 6641 27489 6653 27492
rect 6687 27489 6699 27523
rect 6641 27483 6699 27489
rect 7190 27480 7196 27532
rect 7248 27520 7254 27532
rect 7650 27520 7656 27532
rect 7248 27492 7656 27520
rect 7248 27480 7254 27492
rect 7650 27480 7656 27492
rect 7708 27480 7714 27532
rect 7929 27523 7987 27529
rect 7929 27489 7941 27523
rect 7975 27489 7987 27523
rect 7929 27483 7987 27489
rect 5500 27424 5856 27452
rect 5500 27412 5506 27424
rect 5258 27384 5264 27396
rect 4804 27356 5264 27384
rect 3292 27288 3740 27316
rect 3292 27276 3298 27288
rect 4154 27276 4160 27328
rect 4212 27316 4218 27328
rect 4804 27316 4832 27356
rect 5258 27344 5264 27356
rect 5316 27344 5322 27396
rect 5350 27344 5356 27396
rect 5408 27344 5414 27396
rect 5828 27384 5856 27424
rect 6914 27412 6920 27464
rect 6972 27412 6978 27464
rect 7944 27452 7972 27483
rect 8018 27452 8024 27464
rect 7944 27424 8024 27452
rect 8018 27412 8024 27424
rect 8076 27412 8082 27464
rect 8128 27384 8156 27560
rect 8205 27557 8217 27591
rect 8251 27557 8263 27591
rect 8205 27551 8263 27557
rect 8297 27591 8355 27597
rect 8297 27557 8309 27591
rect 8343 27588 8355 27591
rect 9048 27588 9076 27628
rect 9674 27588 9680 27600
rect 8343 27560 9076 27588
rect 9232 27560 9680 27588
rect 8343 27557 8355 27560
rect 8297 27551 8355 27557
rect 8481 27523 8539 27529
rect 8481 27489 8493 27523
rect 8527 27520 8539 27523
rect 8757 27523 8815 27529
rect 8527 27492 8616 27520
rect 8527 27489 8539 27492
rect 8481 27483 8539 27489
rect 8588 27464 8616 27492
rect 8757 27489 8769 27523
rect 8803 27489 8815 27523
rect 8757 27483 8815 27489
rect 8941 27523 8999 27529
rect 8941 27489 8953 27523
rect 8987 27520 8999 27523
rect 9122 27520 9128 27532
rect 8987 27492 9128 27520
rect 8987 27489 8999 27492
rect 8941 27483 8999 27489
rect 8570 27412 8576 27464
rect 8628 27412 8634 27464
rect 8772 27452 8800 27483
rect 9122 27480 9128 27492
rect 9180 27480 9186 27532
rect 9232 27529 9260 27560
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 9784 27588 9812 27628
rect 11238 27588 11244 27600
rect 9784 27560 11244 27588
rect 11238 27548 11244 27560
rect 11296 27548 11302 27600
rect 9217 27523 9275 27529
rect 9217 27489 9229 27523
rect 9263 27489 9275 27523
rect 9473 27523 9531 27529
rect 9473 27520 9485 27523
rect 9217 27483 9275 27489
rect 9324 27492 9485 27520
rect 9324 27452 9352 27492
rect 9473 27489 9485 27492
rect 9519 27489 9531 27523
rect 9473 27483 9531 27489
rect 8772 27424 8984 27452
rect 8956 27396 8984 27424
rect 9048 27424 9352 27452
rect 8294 27384 8300 27396
rect 5828 27356 6100 27384
rect 8128 27356 8300 27384
rect 4212 27288 4832 27316
rect 4212 27276 4218 27288
rect 4982 27276 4988 27328
rect 5040 27316 5046 27328
rect 5445 27319 5503 27325
rect 5445 27316 5457 27319
rect 5040 27288 5457 27316
rect 5040 27276 5046 27288
rect 5445 27285 5457 27288
rect 5491 27285 5503 27319
rect 5445 27279 5503 27285
rect 5810 27276 5816 27328
rect 5868 27316 5874 27328
rect 5905 27319 5963 27325
rect 5905 27316 5917 27319
rect 5868 27288 5917 27316
rect 5868 27276 5874 27288
rect 5905 27285 5917 27288
rect 5951 27285 5963 27319
rect 6072 27316 6100 27356
rect 8294 27344 8300 27356
rect 8352 27344 8358 27396
rect 8665 27387 8723 27393
rect 8665 27353 8677 27387
rect 8711 27384 8723 27387
rect 8754 27384 8760 27396
rect 8711 27356 8760 27384
rect 8711 27353 8723 27356
rect 8665 27347 8723 27353
rect 8754 27344 8760 27356
rect 8812 27344 8818 27396
rect 8938 27344 8944 27396
rect 8996 27344 9002 27396
rect 6178 27316 6184 27328
rect 6072 27288 6184 27316
rect 5905 27279 5963 27285
rect 6178 27276 6184 27288
rect 6236 27276 6242 27328
rect 7650 27276 7656 27328
rect 7708 27316 7714 27328
rect 8110 27316 8116 27328
rect 7708 27288 8116 27316
rect 7708 27276 7714 27288
rect 8110 27276 8116 27288
rect 8168 27276 8174 27328
rect 8205 27319 8263 27325
rect 8205 27285 8217 27319
rect 8251 27316 8263 27319
rect 9048 27316 9076 27424
rect 8251 27288 9076 27316
rect 9125 27319 9183 27325
rect 8251 27285 8263 27288
rect 8205 27279 8263 27285
rect 9125 27285 9137 27319
rect 9171 27316 9183 27319
rect 9490 27316 9496 27328
rect 9171 27288 9496 27316
rect 9171 27285 9183 27288
rect 9125 27279 9183 27285
rect 9490 27276 9496 27288
rect 9548 27276 9554 27328
rect 10597 27319 10655 27325
rect 10597 27285 10609 27319
rect 10643 27316 10655 27319
rect 10686 27316 10692 27328
rect 10643 27288 10692 27316
rect 10643 27285 10655 27288
rect 10597 27279 10655 27285
rect 10686 27276 10692 27288
rect 10744 27276 10750 27328
rect 552 27226 11132 27248
rect 552 27174 3662 27226
rect 3714 27174 3726 27226
rect 3778 27174 3790 27226
rect 3842 27174 3854 27226
rect 3906 27174 3918 27226
rect 3970 27174 10062 27226
rect 10114 27174 10126 27226
rect 10178 27174 10190 27226
rect 10242 27174 10254 27226
rect 10306 27174 10318 27226
rect 10370 27174 11132 27226
rect 552 27152 11132 27174
rect 1210 27072 1216 27124
rect 1268 27112 1274 27124
rect 2682 27112 2688 27124
rect 1268 27084 2688 27112
rect 1268 27072 1274 27084
rect 2682 27072 2688 27084
rect 2740 27072 2746 27124
rect 2774 27072 2780 27124
rect 2832 27112 2838 27124
rect 3418 27112 3424 27124
rect 2832 27084 3424 27112
rect 2832 27072 2838 27084
rect 3418 27072 3424 27084
rect 3476 27112 3482 27124
rect 3881 27115 3939 27121
rect 3881 27112 3893 27115
rect 3476 27084 3893 27112
rect 3476 27072 3482 27084
rect 3881 27081 3893 27084
rect 3927 27081 3939 27115
rect 4246 27112 4252 27124
rect 3881 27075 3939 27081
rect 3988 27084 4252 27112
rect 3988 27044 4016 27084
rect 4246 27072 4252 27084
rect 4304 27072 4310 27124
rect 4706 27072 4712 27124
rect 4764 27072 4770 27124
rect 6914 27072 6920 27124
rect 6972 27112 6978 27124
rect 7190 27112 7196 27124
rect 6972 27084 7196 27112
rect 6972 27072 6978 27084
rect 7190 27072 7196 27084
rect 7248 27072 7254 27124
rect 7282 27072 7288 27124
rect 7340 27112 7346 27124
rect 7466 27112 7472 27124
rect 7340 27084 7472 27112
rect 7340 27072 7346 27084
rect 7466 27072 7472 27084
rect 7524 27112 7530 27124
rect 7837 27115 7895 27121
rect 7837 27112 7849 27115
rect 7524 27084 7849 27112
rect 7524 27072 7530 27084
rect 7837 27081 7849 27084
rect 7883 27081 7895 27115
rect 7837 27075 7895 27081
rect 8481 27115 8539 27121
rect 8481 27081 8493 27115
rect 8527 27112 8539 27115
rect 10134 27112 10140 27124
rect 8527 27084 10140 27112
rect 8527 27081 8539 27084
rect 8481 27075 8539 27081
rect 10134 27072 10140 27084
rect 10192 27072 10198 27124
rect 2516 27016 4016 27044
rect 842 26936 848 26988
rect 900 26976 906 26988
rect 1673 26979 1731 26985
rect 900 26948 1532 26976
rect 900 26936 906 26948
rect 1121 26911 1179 26917
rect 1121 26877 1133 26911
rect 1167 26877 1179 26911
rect 1121 26871 1179 26877
rect 1213 26911 1271 26917
rect 1213 26877 1225 26911
rect 1259 26877 1271 26911
rect 1213 26871 1271 26877
rect 937 26775 995 26781
rect 937 26741 949 26775
rect 983 26772 995 26775
rect 1026 26772 1032 26784
rect 983 26744 1032 26772
rect 983 26741 995 26744
rect 937 26735 995 26741
rect 1026 26732 1032 26744
rect 1084 26732 1090 26784
rect 1136 26772 1164 26871
rect 1228 26840 1256 26871
rect 1302 26868 1308 26920
rect 1360 26908 1366 26920
rect 1397 26911 1455 26917
rect 1397 26908 1409 26911
rect 1360 26880 1409 26908
rect 1360 26868 1366 26880
rect 1397 26877 1409 26880
rect 1443 26877 1455 26911
rect 1504 26908 1532 26948
rect 1673 26945 1685 26979
rect 1719 26976 1731 26979
rect 1854 26976 1860 26988
rect 1719 26948 1860 26976
rect 1719 26945 1731 26948
rect 1673 26939 1731 26945
rect 1854 26936 1860 26948
rect 1912 26936 1918 26988
rect 2225 26979 2283 26985
rect 2225 26945 2237 26979
rect 2271 26976 2283 26979
rect 2406 26976 2412 26988
rect 2271 26948 2412 26976
rect 2271 26945 2283 26948
rect 2225 26939 2283 26945
rect 2406 26936 2412 26948
rect 2464 26936 2470 26988
rect 2516 26917 2544 27016
rect 4062 27004 4068 27056
rect 4120 27004 4126 27056
rect 2590 26936 2596 26988
rect 2648 26936 2654 26988
rect 2685 26979 2743 26985
rect 2685 26945 2697 26979
rect 2731 26976 2743 26979
rect 3510 26976 3516 26988
rect 2731 26948 3516 26976
rect 2731 26945 2743 26948
rect 2685 26939 2743 26945
rect 3510 26936 3516 26948
rect 3568 26936 3574 26988
rect 4080 26976 4108 27004
rect 3620 26948 4108 26976
rect 4249 26979 4307 26985
rect 3620 26920 3648 26948
rect 4249 26945 4261 26979
rect 4295 26976 4307 26979
rect 4522 26976 4528 26988
rect 4295 26948 4528 26976
rect 4295 26945 4307 26948
rect 4249 26939 4307 26945
rect 4522 26936 4528 26948
rect 4580 26936 4586 26988
rect 4724 26962 4752 27072
rect 6181 27047 6239 27053
rect 6181 27013 6193 27047
rect 6227 27044 6239 27047
rect 7374 27044 7380 27056
rect 6227 27016 7380 27044
rect 6227 27013 6239 27016
rect 6181 27007 6239 27013
rect 7374 27004 7380 27016
rect 7432 27004 7438 27056
rect 8018 27004 8024 27056
rect 8076 27044 8082 27056
rect 8076 27016 9516 27044
rect 8076 27004 8082 27016
rect 6362 26976 6368 26988
rect 6072 26948 6368 26976
rect 2317 26911 2375 26917
rect 2317 26908 2329 26911
rect 1504 26880 2329 26908
rect 1397 26871 1455 26877
rect 2317 26877 2329 26880
rect 2363 26877 2375 26911
rect 2317 26871 2375 26877
rect 2501 26911 2559 26917
rect 2501 26877 2513 26911
rect 2547 26877 2559 26911
rect 2501 26871 2559 26877
rect 2869 26911 2927 26917
rect 2869 26877 2881 26911
rect 2915 26877 2927 26911
rect 2869 26871 2927 26877
rect 1762 26840 1768 26852
rect 1228 26812 1768 26840
rect 1762 26800 1768 26812
rect 1820 26800 1826 26852
rect 2406 26800 2412 26852
rect 2464 26840 2470 26852
rect 2884 26840 2912 26871
rect 3602 26868 3608 26920
rect 3660 26868 3666 26920
rect 4062 26868 4068 26920
rect 4120 26868 4126 26920
rect 4338 26868 4344 26920
rect 4396 26868 4402 26920
rect 4433 26911 4491 26917
rect 4433 26877 4445 26911
rect 4479 26877 4491 26911
rect 4433 26871 4491 26877
rect 4617 26911 4675 26917
rect 4617 26877 4629 26911
rect 4663 26908 4675 26911
rect 5534 26908 5540 26920
rect 4663 26880 5540 26908
rect 4663 26877 4675 26880
rect 4617 26871 4675 26877
rect 2464 26812 3464 26840
rect 2464 26800 2470 26812
rect 1210 26772 1216 26784
rect 1136 26744 1216 26772
rect 1210 26732 1216 26744
rect 1268 26732 1274 26784
rect 2498 26732 2504 26784
rect 2556 26772 2562 26784
rect 3053 26775 3111 26781
rect 3053 26772 3065 26775
rect 2556 26744 3065 26772
rect 2556 26732 2562 26744
rect 3053 26741 3065 26744
rect 3099 26741 3111 26775
rect 3436 26772 3464 26812
rect 3694 26800 3700 26852
rect 3752 26840 3758 26852
rect 4356 26840 4384 26868
rect 3752 26812 4384 26840
rect 4448 26840 4476 26871
rect 5534 26868 5540 26880
rect 5592 26868 5598 26920
rect 5629 26911 5687 26917
rect 5629 26877 5641 26911
rect 5675 26908 5687 26911
rect 6072 26908 6100 26948
rect 6362 26936 6368 26948
rect 6420 26936 6426 26988
rect 7742 26976 7748 26988
rect 6840 26948 7748 26976
rect 5675 26880 6100 26908
rect 5675 26877 5687 26880
rect 5629 26871 5687 26877
rect 6454 26868 6460 26920
rect 6512 26908 6518 26920
rect 6549 26911 6607 26917
rect 6549 26908 6561 26911
rect 6512 26880 6561 26908
rect 6512 26868 6518 26880
rect 6549 26877 6561 26880
rect 6595 26908 6607 26911
rect 6730 26908 6736 26920
rect 6595 26880 6736 26908
rect 6595 26877 6607 26880
rect 6549 26871 6607 26877
rect 6730 26868 6736 26880
rect 6788 26868 6794 26920
rect 6840 26917 6868 26948
rect 7742 26936 7748 26948
rect 7800 26936 7806 26988
rect 8665 26979 8723 26985
rect 8665 26945 8677 26979
rect 8711 26976 8723 26979
rect 8938 26976 8944 26988
rect 8711 26948 8944 26976
rect 8711 26945 8723 26948
rect 8665 26939 8723 26945
rect 8938 26936 8944 26948
rect 8996 26936 9002 26988
rect 9306 26936 9312 26988
rect 9364 26936 9370 26988
rect 6825 26911 6883 26917
rect 6825 26877 6837 26911
rect 6871 26877 6883 26911
rect 6825 26871 6883 26877
rect 6914 26868 6920 26920
rect 6972 26868 6978 26920
rect 7009 26911 7067 26917
rect 7009 26877 7021 26911
rect 7055 26908 7067 26911
rect 7098 26908 7104 26920
rect 7055 26880 7104 26908
rect 7055 26877 7067 26880
rect 7009 26871 7067 26877
rect 7098 26868 7104 26880
rect 7156 26868 7162 26920
rect 7190 26868 7196 26920
rect 7248 26868 7254 26920
rect 8018 26868 8024 26920
rect 8076 26908 8082 26920
rect 8294 26908 8300 26920
rect 8076 26880 8300 26908
rect 8076 26868 8082 26880
rect 8294 26868 8300 26880
rect 8352 26908 8358 26920
rect 8389 26911 8447 26917
rect 8389 26908 8401 26911
rect 8352 26880 8401 26908
rect 8352 26868 8358 26880
rect 8389 26877 8401 26880
rect 8435 26877 8447 26911
rect 8389 26871 8447 26877
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 8757 26911 8815 26917
rect 8757 26908 8769 26911
rect 8628 26880 8769 26908
rect 8628 26868 8634 26880
rect 8757 26877 8769 26880
rect 8803 26877 8815 26911
rect 8757 26871 8815 26877
rect 8846 26868 8852 26920
rect 8904 26868 8910 26920
rect 9030 26868 9036 26920
rect 9088 26868 9094 26920
rect 9122 26868 9128 26920
rect 9180 26868 9186 26920
rect 9324 26908 9352 26936
rect 9324 26880 9444 26908
rect 4706 26840 4712 26852
rect 4448 26812 4712 26840
rect 3752 26800 3758 26812
rect 4706 26800 4712 26812
rect 4764 26800 4770 26852
rect 4890 26800 4896 26852
rect 4948 26800 4954 26852
rect 5074 26800 5080 26852
rect 5132 26840 5138 26852
rect 5169 26843 5227 26849
rect 5169 26840 5181 26843
rect 5132 26812 5181 26840
rect 5132 26800 5138 26812
rect 5169 26809 5181 26812
rect 5215 26809 5227 26843
rect 5169 26803 5227 26809
rect 5261 26843 5319 26849
rect 5261 26809 5273 26843
rect 5307 26809 5319 26843
rect 5261 26803 5319 26809
rect 4614 26772 4620 26784
rect 3436 26744 4620 26772
rect 3053 26735 3111 26741
rect 4614 26732 4620 26744
rect 4672 26732 4678 26784
rect 5276 26772 5304 26803
rect 5994 26800 6000 26852
rect 6052 26800 6058 26852
rect 6270 26800 6276 26852
rect 6328 26840 6334 26852
rect 7469 26843 7527 26849
rect 7469 26840 7481 26843
rect 6328 26812 7481 26840
rect 6328 26800 6334 26812
rect 7469 26809 7481 26812
rect 7515 26809 7527 26843
rect 7469 26803 7527 26809
rect 7650 26800 7656 26852
rect 7708 26800 7714 26852
rect 7742 26800 7748 26852
rect 7800 26840 7806 26852
rect 7929 26843 7987 26849
rect 7929 26840 7941 26843
rect 7800 26812 7941 26840
rect 7800 26800 7806 26812
rect 7929 26809 7941 26812
rect 7975 26809 7987 26843
rect 7929 26803 7987 26809
rect 8202 26800 8208 26852
rect 8260 26840 8266 26852
rect 9309 26843 9367 26849
rect 9309 26840 9321 26843
rect 8260 26812 9321 26840
rect 8260 26800 8266 26812
rect 9309 26809 9321 26812
rect 9355 26809 9367 26843
rect 9309 26803 9367 26809
rect 5626 26772 5632 26784
rect 5276 26744 5632 26772
rect 5626 26732 5632 26744
rect 5684 26732 5690 26784
rect 6362 26732 6368 26784
rect 6420 26772 6426 26784
rect 6457 26775 6515 26781
rect 6457 26772 6469 26775
rect 6420 26744 6469 26772
rect 6420 26732 6426 26744
rect 6457 26741 6469 26744
rect 6503 26741 6515 26775
rect 6457 26735 6515 26741
rect 6638 26732 6644 26784
rect 6696 26732 6702 26784
rect 6730 26732 6736 26784
rect 6788 26772 6794 26784
rect 7190 26772 7196 26784
rect 6788 26744 7196 26772
rect 6788 26732 6794 26744
rect 7190 26732 7196 26744
rect 7248 26732 7254 26784
rect 7282 26732 7288 26784
rect 7340 26732 7346 26784
rect 8665 26775 8723 26781
rect 8665 26741 8677 26775
rect 8711 26772 8723 26775
rect 9122 26772 9128 26784
rect 8711 26744 9128 26772
rect 8711 26741 8723 26744
rect 8665 26735 8723 26741
rect 9122 26732 9128 26744
rect 9180 26732 9186 26784
rect 9416 26781 9444 26880
rect 9401 26775 9459 26781
rect 9401 26741 9413 26775
rect 9447 26741 9459 26775
rect 9488 26772 9516 27016
rect 9674 26868 9680 26920
rect 9732 26908 9738 26920
rect 10781 26911 10839 26917
rect 10781 26908 10793 26911
rect 9732 26880 10793 26908
rect 9732 26868 9738 26880
rect 10781 26877 10793 26880
rect 10827 26877 10839 26911
rect 10781 26871 10839 26877
rect 10502 26800 10508 26852
rect 10560 26849 10566 26852
rect 10560 26840 10572 26849
rect 10560 26812 10605 26840
rect 10560 26803 10572 26812
rect 10560 26800 10566 26803
rect 11330 26772 11336 26784
rect 9488 26744 11336 26772
rect 9401 26735 9459 26741
rect 11330 26732 11336 26744
rect 11388 26732 11394 26784
rect 552 26682 11132 26704
rect 552 26630 4322 26682
rect 4374 26630 4386 26682
rect 4438 26630 4450 26682
rect 4502 26630 4514 26682
rect 4566 26630 4578 26682
rect 4630 26630 10722 26682
rect 10774 26630 10786 26682
rect 10838 26630 10850 26682
rect 10902 26630 10914 26682
rect 10966 26630 10978 26682
rect 11030 26630 11132 26682
rect 552 26608 11132 26630
rect 1029 26571 1087 26577
rect 1029 26537 1041 26571
rect 1075 26568 1087 26571
rect 1118 26568 1124 26580
rect 1075 26540 1124 26568
rect 1075 26537 1087 26540
rect 1029 26531 1087 26537
rect 1118 26528 1124 26540
rect 1176 26528 1182 26580
rect 1670 26528 1676 26580
rect 1728 26528 1734 26580
rect 2038 26528 2044 26580
rect 2096 26528 2102 26580
rect 2774 26528 2780 26580
rect 2832 26568 2838 26580
rect 3694 26568 3700 26580
rect 2832 26540 3700 26568
rect 2832 26528 2838 26540
rect 3694 26528 3700 26540
rect 3752 26528 3758 26580
rect 4062 26528 4068 26580
rect 4120 26568 4126 26580
rect 4614 26568 4620 26580
rect 4120 26540 4620 26568
rect 4120 26528 4126 26540
rect 4614 26528 4620 26540
rect 4672 26528 4678 26580
rect 4706 26528 4712 26580
rect 4764 26568 4770 26580
rect 5258 26568 5264 26580
rect 4764 26540 5264 26568
rect 4764 26528 4770 26540
rect 5258 26528 5264 26540
rect 5316 26528 5322 26580
rect 5350 26528 5356 26580
rect 5408 26568 5414 26580
rect 5534 26568 5540 26580
rect 5408 26540 5540 26568
rect 5408 26528 5414 26540
rect 5534 26528 5540 26540
rect 5592 26528 5598 26580
rect 5994 26528 6000 26580
rect 6052 26568 6058 26580
rect 7742 26568 7748 26580
rect 6052 26540 7748 26568
rect 6052 26528 6058 26540
rect 7742 26528 7748 26540
rect 7800 26528 7806 26580
rect 8205 26571 8263 26577
rect 8205 26537 8217 26571
rect 8251 26568 8263 26571
rect 9030 26568 9036 26580
rect 8251 26540 9036 26568
rect 8251 26537 8263 26540
rect 8205 26531 8263 26537
rect 9030 26528 9036 26540
rect 9088 26528 9094 26580
rect 9306 26528 9312 26580
rect 9364 26528 9370 26580
rect 1688 26500 1716 26528
rect 3053 26503 3111 26509
rect 1688 26472 2084 26500
rect 2056 26444 2084 26472
rect 3053 26469 3065 26503
rect 3099 26500 3111 26503
rect 4522 26500 4528 26512
rect 3099 26472 4528 26500
rect 3099 26469 3111 26472
rect 3053 26463 3111 26469
rect 4522 26460 4528 26472
rect 4580 26460 4586 26512
rect 5626 26460 5632 26512
rect 5684 26500 5690 26512
rect 6362 26500 6368 26512
rect 5684 26472 6368 26500
rect 5684 26460 5690 26472
rect 6362 26460 6368 26472
rect 6420 26500 6426 26512
rect 6420 26472 6592 26500
rect 6420 26460 6426 26472
rect 842 26392 848 26444
rect 900 26392 906 26444
rect 1026 26392 1032 26444
rect 1084 26392 1090 26444
rect 1394 26392 1400 26444
rect 1452 26392 1458 26444
rect 1670 26392 1676 26444
rect 1728 26392 1734 26444
rect 1946 26392 1952 26444
rect 2004 26392 2010 26444
rect 2038 26392 2044 26444
rect 2096 26392 2102 26444
rect 2222 26392 2228 26444
rect 2280 26392 2286 26444
rect 2498 26392 2504 26444
rect 2556 26392 2562 26444
rect 2685 26435 2743 26441
rect 2685 26401 2697 26435
rect 2731 26401 2743 26435
rect 2685 26395 2743 26401
rect 3237 26435 3295 26441
rect 3237 26401 3249 26435
rect 3283 26432 3295 26435
rect 4706 26432 4712 26444
rect 3283 26404 4712 26432
rect 3283 26401 3295 26404
rect 3237 26395 3295 26401
rect 2406 26364 2412 26376
rect 1412 26336 2412 26364
rect 1412 26308 1440 26336
rect 2406 26324 2412 26336
rect 2464 26324 2470 26376
rect 1394 26256 1400 26308
rect 1452 26256 1458 26308
rect 1857 26299 1915 26305
rect 1857 26265 1869 26299
rect 1903 26296 1915 26299
rect 2130 26296 2136 26308
rect 1903 26268 2136 26296
rect 1903 26265 1915 26268
rect 1857 26259 1915 26265
rect 2130 26256 2136 26268
rect 2188 26256 2194 26308
rect 2222 26256 2228 26308
rect 2280 26296 2286 26308
rect 2700 26296 2728 26395
rect 4706 26392 4712 26404
rect 4764 26392 4770 26444
rect 5074 26392 5080 26444
rect 5132 26392 5138 26444
rect 5350 26392 5356 26444
rect 5408 26392 5414 26444
rect 5813 26435 5871 26441
rect 5813 26432 5825 26435
rect 5460 26404 5825 26432
rect 3050 26324 3056 26376
rect 3108 26364 3114 26376
rect 5460 26364 5488 26404
rect 5813 26401 5825 26404
rect 5859 26432 5871 26435
rect 6086 26432 6092 26444
rect 5859 26404 6092 26432
rect 5859 26401 5871 26404
rect 5813 26395 5871 26401
rect 6086 26392 6092 26404
rect 6144 26392 6150 26444
rect 6270 26392 6276 26444
rect 6328 26432 6334 26444
rect 6564 26441 6592 26472
rect 7006 26460 7012 26512
rect 7064 26460 7070 26512
rect 8662 26500 8668 26512
rect 7760 26472 8668 26500
rect 6457 26435 6515 26441
rect 6457 26432 6469 26435
rect 6328 26404 6469 26432
rect 6328 26392 6334 26404
rect 6457 26401 6469 26404
rect 6503 26401 6515 26435
rect 6457 26395 6515 26401
rect 6549 26435 6607 26441
rect 6549 26401 6561 26435
rect 6595 26401 6607 26435
rect 6549 26395 6607 26401
rect 6638 26392 6644 26444
rect 6696 26392 6702 26444
rect 7190 26392 7196 26444
rect 7248 26392 7254 26444
rect 7469 26435 7527 26441
rect 7469 26401 7481 26435
rect 7515 26432 7527 26435
rect 7558 26432 7564 26444
rect 7515 26404 7564 26432
rect 7515 26401 7527 26404
rect 7469 26395 7527 26401
rect 7558 26392 7564 26404
rect 7616 26392 7622 26444
rect 7760 26441 7788 26472
rect 8662 26460 8668 26472
rect 8720 26460 8726 26512
rect 9324 26500 9352 26528
rect 9048 26472 9352 26500
rect 9048 26444 9076 26472
rect 9582 26460 9588 26512
rect 9640 26500 9646 26512
rect 9640 26472 9996 26500
rect 9640 26460 9646 26472
rect 7653 26435 7711 26441
rect 7653 26401 7665 26435
rect 7699 26401 7711 26435
rect 7653 26395 7711 26401
rect 7745 26435 7803 26441
rect 7745 26401 7757 26435
rect 7791 26401 7803 26435
rect 7745 26395 7803 26401
rect 8021 26435 8079 26441
rect 8021 26401 8033 26435
rect 8067 26432 8079 26435
rect 8110 26432 8116 26444
rect 8067 26404 8116 26432
rect 8067 26401 8079 26404
rect 8021 26395 8079 26401
rect 3108 26336 5488 26364
rect 3108 26324 3114 26336
rect 5534 26324 5540 26376
rect 5592 26364 5598 26376
rect 5629 26367 5687 26373
rect 5629 26364 5641 26367
rect 5592 26336 5641 26364
rect 5592 26324 5598 26336
rect 5629 26333 5641 26336
rect 5675 26333 5687 26367
rect 5629 26327 5687 26333
rect 6365 26367 6423 26373
rect 6365 26333 6377 26367
rect 6411 26364 6423 26367
rect 6730 26364 6736 26376
rect 6411 26336 6736 26364
rect 6411 26333 6423 26336
rect 6365 26327 6423 26333
rect 2280 26268 3740 26296
rect 2280 26256 2286 26268
rect 1118 26188 1124 26240
rect 1176 26228 1182 26240
rect 1213 26231 1271 26237
rect 1213 26228 1225 26231
rect 1176 26200 1225 26228
rect 1176 26188 1182 26200
rect 1213 26197 1225 26200
rect 1259 26197 1271 26231
rect 1213 26191 1271 26197
rect 1486 26188 1492 26240
rect 1544 26188 1550 26240
rect 1946 26188 1952 26240
rect 2004 26228 2010 26240
rect 2314 26228 2320 26240
rect 2004 26200 2320 26228
rect 2004 26188 2010 26200
rect 2314 26188 2320 26200
rect 2372 26188 2378 26240
rect 2682 26188 2688 26240
rect 2740 26228 2746 26240
rect 3602 26228 3608 26240
rect 2740 26200 3608 26228
rect 2740 26188 2746 26200
rect 3602 26188 3608 26200
rect 3660 26188 3666 26240
rect 3712 26228 3740 26268
rect 3786 26256 3792 26308
rect 3844 26296 3850 26308
rect 5169 26299 5227 26305
rect 5169 26296 5181 26299
rect 3844 26268 5181 26296
rect 3844 26256 3850 26268
rect 5169 26265 5181 26268
rect 5215 26265 5227 26299
rect 5644 26296 5672 26327
rect 6730 26324 6736 26336
rect 6788 26324 6794 26376
rect 5997 26299 6055 26305
rect 5997 26296 6009 26299
rect 5169 26259 5227 26265
rect 5460 26268 6009 26296
rect 5460 26228 5488 26268
rect 5997 26265 6009 26268
rect 6043 26296 6055 26299
rect 6270 26296 6276 26308
rect 6043 26268 6276 26296
rect 6043 26265 6055 26268
rect 5997 26259 6055 26265
rect 6270 26256 6276 26268
rect 6328 26256 6334 26308
rect 6454 26256 6460 26308
rect 6512 26296 6518 26308
rect 7668 26296 7696 26395
rect 8110 26392 8116 26404
rect 8168 26392 8174 26444
rect 8294 26392 8300 26444
rect 8352 26432 8358 26444
rect 8573 26435 8631 26441
rect 8573 26432 8585 26435
rect 8352 26404 8585 26432
rect 8352 26392 8358 26404
rect 8573 26401 8585 26404
rect 8619 26401 8631 26435
rect 8573 26395 8631 26401
rect 9030 26392 9036 26444
rect 9088 26392 9094 26444
rect 9306 26392 9312 26444
rect 9364 26392 9370 26444
rect 9493 26435 9551 26441
rect 9493 26401 9505 26435
rect 9539 26401 9551 26435
rect 9493 26395 9551 26401
rect 9861 26435 9919 26441
rect 9861 26401 9873 26435
rect 9907 26401 9919 26435
rect 9861 26395 9919 26401
rect 7837 26367 7895 26373
rect 7837 26333 7849 26367
rect 7883 26333 7895 26367
rect 9401 26367 9459 26373
rect 9401 26364 9413 26367
rect 7837 26327 7895 26333
rect 8588 26336 9413 26364
rect 6512 26268 7696 26296
rect 6512 26256 6518 26268
rect 3712 26200 5488 26228
rect 5534 26188 5540 26240
rect 5592 26188 5598 26240
rect 6181 26231 6239 26237
rect 6181 26197 6193 26231
rect 6227 26228 6239 26231
rect 6362 26228 6368 26240
rect 6227 26200 6368 26228
rect 6227 26197 6239 26200
rect 6181 26191 6239 26197
rect 6362 26188 6368 26200
rect 6420 26188 6426 26240
rect 6825 26231 6883 26237
rect 6825 26197 6837 26231
rect 6871 26228 6883 26231
rect 7190 26228 7196 26240
rect 6871 26200 7196 26228
rect 6871 26197 6883 26200
rect 6825 26191 6883 26197
rect 7190 26188 7196 26200
rect 7248 26188 7254 26240
rect 7466 26188 7472 26240
rect 7524 26228 7530 26240
rect 7852 26228 7880 26327
rect 8588 26308 8616 26336
rect 9401 26333 9413 26336
rect 9447 26333 9459 26367
rect 9401 26327 9459 26333
rect 8570 26256 8576 26308
rect 8628 26256 8634 26308
rect 9214 26256 9220 26308
rect 9272 26296 9278 26308
rect 9508 26296 9536 26395
rect 9769 26367 9827 26373
rect 9769 26333 9781 26367
rect 9815 26333 9827 26367
rect 9769 26327 9827 26333
rect 9272 26268 9536 26296
rect 9272 26256 9278 26268
rect 7524 26200 7880 26228
rect 7524 26188 7530 26200
rect 9306 26188 9312 26240
rect 9364 26228 9370 26240
rect 9784 26228 9812 26327
rect 9364 26200 9812 26228
rect 9876 26228 9904 26395
rect 9968 26364 9996 26472
rect 10134 26392 10140 26444
rect 10192 26432 10198 26444
rect 10505 26435 10563 26441
rect 10505 26432 10517 26435
rect 10192 26404 10517 26432
rect 10192 26392 10198 26404
rect 10505 26401 10517 26404
rect 10551 26432 10563 26435
rect 11238 26432 11244 26444
rect 10551 26404 11244 26432
rect 10551 26401 10563 26404
rect 10505 26395 10563 26401
rect 11238 26392 11244 26404
rect 11296 26392 11302 26444
rect 10321 26367 10379 26373
rect 10321 26364 10333 26367
rect 9968 26336 10333 26364
rect 10321 26333 10333 26336
rect 10367 26333 10379 26367
rect 10321 26327 10379 26333
rect 9950 26256 9956 26308
rect 10008 26296 10014 26308
rect 10229 26299 10287 26305
rect 10229 26296 10241 26299
rect 10008 26268 10241 26296
rect 10008 26256 10014 26268
rect 10229 26265 10241 26268
rect 10275 26265 10287 26299
rect 10229 26259 10287 26265
rect 10042 26228 10048 26240
rect 9876 26200 10048 26228
rect 9364 26188 9370 26200
rect 10042 26188 10048 26200
rect 10100 26188 10106 26240
rect 10502 26188 10508 26240
rect 10560 26228 10566 26240
rect 10689 26231 10747 26237
rect 10689 26228 10701 26231
rect 10560 26200 10701 26228
rect 10560 26188 10566 26200
rect 10689 26197 10701 26200
rect 10735 26197 10747 26231
rect 10689 26191 10747 26197
rect 552 26138 11132 26160
rect 552 26086 3662 26138
rect 3714 26086 3726 26138
rect 3778 26086 3790 26138
rect 3842 26086 3854 26138
rect 3906 26086 3918 26138
rect 3970 26086 10062 26138
rect 10114 26086 10126 26138
rect 10178 26086 10190 26138
rect 10242 26086 10254 26138
rect 10306 26086 10318 26138
rect 10370 26086 11132 26138
rect 552 26064 11132 26086
rect 937 26027 995 26033
rect 937 25993 949 26027
rect 983 26024 995 26027
rect 1394 26024 1400 26036
rect 983 25996 1400 26024
rect 983 25993 995 25996
rect 937 25987 995 25993
rect 1394 25984 1400 25996
rect 1452 25984 1458 26036
rect 2314 25984 2320 26036
rect 2372 26024 2378 26036
rect 2961 26027 3019 26033
rect 2961 26024 2973 26027
rect 2372 25996 2973 26024
rect 2372 25984 2378 25996
rect 2961 25993 2973 25996
rect 3007 25993 3019 26027
rect 2961 25987 3019 25993
rect 3510 25984 3516 26036
rect 3568 26024 3574 26036
rect 3568 25996 4191 26024
rect 3568 25984 3574 25996
rect 1578 25916 1584 25968
rect 1636 25956 1642 25968
rect 1636 25928 2268 25956
rect 1636 25916 1642 25928
rect 1213 25891 1271 25897
rect 1213 25857 1225 25891
rect 1259 25888 1271 25891
rect 1394 25888 1400 25900
rect 1259 25860 1400 25888
rect 1259 25857 1271 25860
rect 1213 25851 1271 25857
rect 1394 25848 1400 25860
rect 1452 25848 1458 25900
rect 1486 25848 1492 25900
rect 1544 25888 1550 25900
rect 1765 25891 1823 25897
rect 1765 25888 1777 25891
rect 1544 25860 1777 25888
rect 1544 25848 1550 25860
rect 1765 25857 1777 25860
rect 1811 25857 1823 25891
rect 1765 25851 1823 25857
rect 2240 25832 2268 25928
rect 2498 25916 2504 25968
rect 2556 25916 2562 25968
rect 2590 25916 2596 25968
rect 2648 25956 2654 25968
rect 3050 25956 3056 25968
rect 2648 25928 3056 25956
rect 2648 25916 2654 25928
rect 3050 25916 3056 25928
rect 3108 25916 3114 25968
rect 3234 25916 3240 25968
rect 3292 25916 3298 25968
rect 3878 25956 3884 25968
rect 3712 25928 3884 25956
rect 2516 25888 2544 25916
rect 2516 25860 2728 25888
rect 1121 25823 1179 25829
rect 1121 25789 1133 25823
rect 1167 25820 1179 25823
rect 1302 25820 1308 25832
rect 1167 25792 1308 25820
rect 1167 25789 1179 25792
rect 1121 25783 1179 25789
rect 1302 25780 1308 25792
rect 1360 25780 1366 25832
rect 2041 25823 2099 25829
rect 2041 25789 2053 25823
rect 2087 25789 2099 25823
rect 2041 25783 2099 25789
rect 842 25712 848 25764
rect 900 25752 906 25764
rect 2056 25752 2084 25783
rect 2222 25780 2228 25832
rect 2280 25780 2286 25832
rect 2314 25780 2320 25832
rect 2372 25818 2378 25832
rect 2409 25823 2467 25829
rect 2409 25818 2421 25823
rect 2372 25790 2421 25818
rect 2372 25780 2378 25790
rect 2409 25789 2421 25790
rect 2455 25789 2467 25823
rect 2409 25783 2467 25789
rect 2498 25780 2504 25832
rect 2556 25780 2562 25832
rect 2590 25780 2596 25832
rect 2648 25829 2654 25832
rect 2648 25823 2670 25829
rect 2658 25789 2670 25823
rect 2648 25783 2670 25789
rect 2648 25780 2654 25783
rect 2700 25752 2728 25860
rect 3418 25848 3424 25900
rect 3476 25848 3482 25900
rect 3602 25848 3608 25900
rect 3660 25848 3666 25900
rect 2777 25823 2835 25829
rect 2777 25789 2789 25823
rect 2823 25820 2835 25823
rect 2958 25820 2964 25832
rect 2823 25792 2964 25820
rect 2823 25789 2835 25792
rect 2777 25783 2835 25789
rect 900 25724 1900 25752
rect 2056 25724 2728 25752
rect 900 25712 906 25724
rect 1578 25644 1584 25696
rect 1636 25684 1642 25696
rect 1762 25684 1768 25696
rect 1636 25656 1768 25684
rect 1636 25644 1642 25656
rect 1762 25644 1768 25656
rect 1820 25644 1826 25696
rect 1872 25684 1900 25724
rect 2792 25684 2820 25783
rect 2958 25780 2964 25792
rect 3016 25780 3022 25832
rect 3427 25807 3455 25848
rect 3513 25823 3571 25829
rect 3413 25801 3471 25807
rect 3413 25767 3425 25801
rect 3459 25767 3471 25801
rect 3513 25789 3525 25823
rect 3559 25820 3571 25823
rect 3620 25820 3648 25848
rect 3712 25829 3740 25928
rect 3878 25916 3884 25928
rect 3936 25916 3942 25968
rect 3988 25888 4016 25996
rect 4163 25956 4191 25996
rect 4246 25984 4252 26036
rect 4304 26024 4310 26036
rect 4709 26027 4767 26033
rect 4709 26024 4721 26027
rect 4304 25996 4721 26024
rect 4304 25984 4310 25996
rect 4709 25993 4721 25996
rect 4755 25993 4767 26027
rect 5537 26027 5595 26033
rect 5537 26024 5549 26027
rect 4709 25987 4767 25993
rect 4908 25996 5549 26024
rect 4908 25956 4936 25996
rect 5537 25993 5549 25996
rect 5583 25993 5595 26027
rect 6638 26024 6644 26036
rect 5537 25987 5595 25993
rect 5828 25996 6644 26024
rect 4163 25928 4936 25956
rect 4982 25916 4988 25968
rect 5040 25916 5046 25968
rect 5629 25959 5687 25965
rect 5629 25925 5641 25959
rect 5675 25956 5687 25959
rect 5718 25956 5724 25968
rect 5675 25928 5724 25956
rect 5675 25925 5687 25928
rect 5629 25919 5687 25925
rect 5718 25916 5724 25928
rect 5776 25916 5782 25968
rect 4065 25891 4123 25897
rect 4065 25888 4077 25891
rect 3988 25860 4077 25888
rect 4065 25857 4077 25860
rect 4111 25857 4123 25891
rect 5000 25888 5028 25916
rect 5077 25891 5135 25897
rect 5077 25888 5089 25891
rect 5000 25860 5089 25888
rect 4065 25851 4123 25857
rect 5077 25857 5089 25860
rect 5123 25857 5135 25891
rect 5077 25851 5135 25857
rect 5169 25891 5227 25897
rect 5169 25857 5181 25891
rect 5215 25888 5227 25891
rect 5828 25888 5856 25996
rect 6638 25984 6644 25996
rect 6696 25984 6702 26036
rect 6730 25984 6736 26036
rect 6788 26024 6794 26036
rect 7006 26024 7012 26036
rect 6788 25996 7012 26024
rect 6788 25984 6794 25996
rect 7006 25984 7012 25996
rect 7064 25984 7070 26036
rect 8202 26024 8208 26036
rect 7116 25996 8208 26024
rect 6178 25916 6184 25968
rect 6236 25956 6242 25968
rect 6236 25928 6960 25956
rect 6236 25916 6242 25928
rect 5215 25860 5856 25888
rect 5215 25857 5227 25860
rect 5169 25851 5227 25857
rect 5902 25848 5908 25900
rect 5960 25888 5966 25900
rect 6730 25888 6736 25900
rect 5960 25860 6736 25888
rect 5960 25848 5966 25860
rect 6730 25848 6736 25860
rect 6788 25848 6794 25900
rect 3559 25792 3648 25820
rect 3697 25823 3755 25829
rect 3559 25789 3571 25792
rect 3513 25783 3571 25789
rect 3697 25789 3709 25823
rect 3743 25789 3755 25823
rect 3697 25783 3755 25789
rect 3413 25761 3471 25767
rect 1872 25656 2820 25684
rect 3050 25644 3056 25696
rect 3108 25684 3114 25696
rect 3234 25684 3240 25696
rect 3108 25656 3240 25684
rect 3108 25644 3114 25656
rect 3234 25644 3240 25656
rect 3292 25644 3298 25696
rect 3427 25684 3455 25761
rect 3520 25752 3548 25783
rect 3786 25780 3792 25832
rect 3844 25780 3850 25832
rect 3878 25780 3884 25832
rect 3936 25818 3942 25832
rect 4261 25820 4552 25822
rect 3988 25818 4099 25820
rect 4172 25818 4552 25820
rect 3936 25794 4552 25818
rect 3936 25792 4289 25794
rect 3936 25790 4016 25792
rect 4071 25790 4200 25792
rect 3936 25780 3942 25790
rect 4249 25755 4307 25761
rect 4249 25752 4261 25755
rect 3520 25724 4261 25752
rect 4249 25721 4261 25724
rect 4295 25721 4307 25755
rect 4249 25715 4307 25721
rect 4430 25712 4436 25764
rect 4488 25712 4494 25764
rect 3878 25684 3884 25696
rect 3427 25656 3884 25684
rect 3878 25644 3884 25656
rect 3936 25644 3942 25696
rect 4341 25687 4399 25693
rect 4341 25653 4353 25687
rect 4387 25684 4399 25687
rect 4448 25684 4476 25712
rect 4387 25656 4476 25684
rect 4524 25684 4552 25794
rect 4706 25780 4712 25832
rect 4764 25818 4770 25832
rect 4801 25823 4859 25829
rect 4801 25818 4813 25823
rect 4764 25790 4813 25818
rect 4764 25780 4770 25790
rect 4801 25789 4813 25790
rect 4847 25789 4859 25823
rect 4801 25783 4859 25789
rect 4982 25780 4988 25832
rect 5040 25780 5046 25832
rect 5353 25823 5411 25829
rect 5353 25820 5365 25823
rect 5351 25789 5365 25820
rect 5399 25789 5411 25823
rect 5351 25783 5411 25789
rect 4890 25712 4896 25764
rect 4948 25712 4954 25764
rect 4798 25684 4804 25696
rect 4524 25656 4804 25684
rect 4387 25653 4399 25656
rect 4341 25647 4399 25653
rect 4798 25644 4804 25656
rect 4856 25644 4862 25696
rect 4908 25684 4936 25712
rect 5351 25684 5379 25783
rect 5718 25780 5724 25832
rect 5776 25820 5782 25832
rect 5813 25823 5871 25829
rect 5813 25820 5825 25823
rect 5776 25792 5825 25820
rect 5776 25780 5782 25792
rect 5813 25789 5825 25792
rect 5859 25789 5871 25823
rect 5813 25783 5871 25789
rect 6086 25780 6092 25832
rect 6144 25780 6150 25832
rect 6181 25823 6239 25829
rect 6181 25789 6193 25823
rect 6227 25820 6239 25823
rect 6546 25820 6552 25832
rect 6227 25792 6552 25820
rect 6227 25789 6239 25792
rect 6181 25783 6239 25789
rect 6546 25780 6552 25792
rect 6604 25780 6610 25832
rect 6638 25780 6644 25832
rect 6696 25820 6702 25832
rect 6932 25829 6960 25928
rect 6825 25823 6883 25829
rect 6825 25820 6837 25823
rect 6696 25792 6837 25820
rect 6696 25780 6702 25792
rect 6825 25789 6837 25792
rect 6871 25789 6883 25823
rect 6825 25783 6883 25789
rect 6917 25823 6975 25829
rect 6917 25789 6929 25823
rect 6963 25789 6975 25823
rect 6917 25783 6975 25789
rect 7009 25823 7067 25829
rect 7009 25789 7021 25823
rect 7055 25820 7067 25823
rect 7116 25820 7144 25996
rect 8202 25984 8208 25996
rect 8260 25984 8266 26036
rect 8294 25984 8300 26036
rect 8352 26024 8358 26036
rect 9582 26024 9588 26036
rect 8352 25996 9588 26024
rect 8352 25984 8358 25996
rect 9582 25984 9588 25996
rect 9640 26024 9646 26036
rect 9769 26027 9827 26033
rect 9769 26024 9781 26027
rect 9640 25996 9781 26024
rect 9640 25984 9646 25996
rect 9769 25993 9781 25996
rect 9815 25993 9827 26027
rect 9769 25987 9827 25993
rect 7558 25916 7564 25968
rect 7616 25956 7622 25968
rect 7616 25928 7696 25956
rect 7616 25916 7622 25928
rect 7282 25848 7288 25900
rect 7340 25848 7346 25900
rect 7668 25897 7696 25928
rect 9030 25916 9036 25968
rect 9088 25956 9094 25968
rect 10042 25956 10048 25968
rect 9088 25928 10048 25956
rect 9088 25916 9094 25928
rect 10042 25916 10048 25928
rect 10100 25916 10106 25968
rect 7653 25891 7711 25897
rect 7653 25888 7665 25891
rect 7392 25860 7665 25888
rect 7055 25792 7144 25820
rect 7055 25789 7067 25792
rect 7009 25783 7067 25789
rect 7190 25780 7196 25832
rect 7248 25780 7254 25832
rect 7300 25819 7328 25848
rect 7285 25813 7343 25819
rect 5997 25755 6055 25761
rect 5997 25721 6009 25755
rect 6043 25752 6055 25755
rect 7208 25752 7236 25780
rect 7285 25779 7297 25813
rect 7331 25779 7343 25813
rect 7285 25773 7343 25779
rect 7392 25764 7420 25860
rect 7653 25857 7665 25860
rect 7699 25857 7711 25891
rect 8386 25888 8392 25900
rect 7653 25851 7711 25857
rect 7760 25860 8392 25888
rect 7469 25823 7527 25829
rect 7469 25789 7481 25823
rect 7515 25789 7527 25823
rect 7469 25783 7527 25789
rect 6043 25724 7236 25752
rect 6043 25721 6055 25724
rect 5997 25715 6055 25721
rect 7374 25712 7380 25764
rect 7432 25712 7438 25764
rect 4908 25656 5379 25684
rect 5718 25644 5724 25696
rect 5776 25684 5782 25696
rect 6365 25687 6423 25693
rect 6365 25684 6377 25687
rect 5776 25656 6377 25684
rect 5776 25644 5782 25656
rect 6365 25653 6377 25656
rect 6411 25653 6423 25687
rect 6365 25647 6423 25653
rect 6546 25644 6552 25696
rect 6604 25644 6610 25696
rect 6730 25644 6736 25696
rect 6788 25684 6794 25696
rect 7282 25684 7288 25696
rect 6788 25656 7288 25684
rect 6788 25644 6794 25656
rect 7282 25644 7288 25656
rect 7340 25684 7346 25696
rect 7484 25684 7512 25783
rect 7558 25780 7564 25832
rect 7616 25820 7622 25832
rect 7760 25820 7788 25860
rect 8386 25848 8392 25860
rect 8444 25848 8450 25900
rect 7616 25792 7788 25820
rect 7616 25780 7622 25792
rect 7834 25780 7840 25832
rect 7892 25780 7898 25832
rect 8478 25780 8484 25832
rect 8536 25780 8542 25832
rect 10502 25780 10508 25832
rect 10560 25780 10566 25832
rect 10594 25780 10600 25832
rect 10652 25820 10658 25832
rect 10689 25823 10747 25829
rect 10689 25820 10701 25823
rect 10652 25792 10701 25820
rect 10652 25780 10658 25792
rect 10689 25789 10701 25792
rect 10735 25789 10747 25823
rect 10689 25783 10747 25789
rect 7340 25656 7512 25684
rect 7340 25644 7346 25656
rect 8018 25644 8024 25696
rect 8076 25644 8082 25696
rect 9030 25644 9036 25696
rect 9088 25684 9094 25696
rect 10321 25687 10379 25693
rect 10321 25684 10333 25687
rect 9088 25656 10333 25684
rect 9088 25644 9094 25656
rect 10321 25653 10333 25656
rect 10367 25653 10379 25687
rect 10321 25647 10379 25653
rect 552 25594 11132 25616
rect 552 25542 4322 25594
rect 4374 25542 4386 25594
rect 4438 25542 4450 25594
rect 4502 25542 4514 25594
rect 4566 25542 4578 25594
rect 4630 25542 10722 25594
rect 10774 25542 10786 25594
rect 10838 25542 10850 25594
rect 10902 25542 10914 25594
rect 10966 25542 10978 25594
rect 11030 25542 11132 25594
rect 552 25520 11132 25542
rect 1121 25483 1179 25489
rect 1121 25449 1133 25483
rect 1167 25480 1179 25483
rect 2498 25480 2504 25492
rect 1167 25452 2504 25480
rect 1167 25449 1179 25452
rect 1121 25443 1179 25449
rect 2498 25440 2504 25452
rect 2556 25440 2562 25492
rect 2958 25440 2964 25492
rect 3016 25480 3022 25492
rect 3329 25483 3387 25489
rect 3016 25452 3280 25480
rect 3016 25440 3022 25452
rect 1578 25372 1584 25424
rect 1636 25412 1642 25424
rect 1636 25384 2360 25412
rect 1636 25372 1642 25384
rect 845 25347 903 25353
rect 845 25313 857 25347
rect 891 25344 903 25347
rect 934 25344 940 25356
rect 891 25316 940 25344
rect 891 25313 903 25316
rect 845 25307 903 25313
rect 934 25304 940 25316
rect 992 25304 998 25356
rect 1486 25304 1492 25356
rect 1544 25344 1550 25356
rect 1765 25347 1823 25353
rect 1765 25344 1777 25347
rect 1544 25316 1777 25344
rect 1544 25304 1550 25316
rect 1765 25313 1777 25316
rect 1811 25313 1823 25347
rect 1765 25307 1823 25313
rect 2041 25347 2099 25353
rect 2041 25313 2053 25347
rect 2087 25313 2099 25347
rect 2041 25307 2099 25313
rect 1118 25236 1124 25288
rect 1176 25236 1182 25288
rect 1210 25236 1216 25288
rect 1268 25236 1274 25288
rect 842 25168 848 25220
rect 900 25208 906 25220
rect 937 25211 995 25217
rect 937 25208 949 25211
rect 900 25180 949 25208
rect 900 25168 906 25180
rect 937 25177 949 25180
rect 983 25177 995 25211
rect 1136 25208 1164 25236
rect 1578 25208 1584 25220
rect 1136 25180 1584 25208
rect 937 25171 995 25177
rect 1578 25168 1584 25180
rect 1636 25168 1642 25220
rect 2056 25208 2084 25307
rect 2222 25304 2228 25356
rect 2280 25304 2286 25356
rect 2332 25344 2360 25384
rect 2406 25372 2412 25424
rect 2464 25412 2470 25424
rect 2464 25384 2636 25412
rect 2464 25372 2470 25384
rect 2501 25347 2559 25353
rect 2501 25344 2513 25347
rect 2332 25316 2513 25344
rect 2501 25313 2513 25316
rect 2547 25313 2559 25347
rect 2608 25344 2636 25384
rect 2774 25372 2780 25424
rect 2832 25412 2838 25424
rect 3145 25415 3203 25421
rect 3145 25412 3157 25415
rect 2832 25384 3157 25412
rect 2832 25372 2838 25384
rect 3145 25381 3157 25384
rect 3191 25381 3203 25415
rect 3252 25412 3280 25452
rect 3329 25449 3341 25483
rect 3375 25480 3387 25483
rect 3375 25452 4568 25480
rect 3375 25449 3387 25452
rect 3329 25443 3387 25449
rect 3605 25415 3663 25421
rect 3605 25412 3617 25415
rect 3252 25384 3617 25412
rect 3145 25375 3203 25381
rect 3605 25381 3617 25384
rect 3651 25381 3663 25415
rect 3605 25375 3663 25381
rect 2958 25344 2964 25356
rect 2608 25316 2964 25344
rect 2501 25307 2559 25313
rect 2958 25304 2964 25316
rect 3016 25304 3022 25356
rect 3050 25304 3056 25356
rect 3108 25304 3114 25356
rect 2130 25236 2136 25288
rect 2188 25276 2194 25288
rect 2685 25279 2743 25285
rect 2685 25276 2697 25279
rect 2188 25248 2697 25276
rect 2188 25236 2194 25248
rect 2685 25245 2697 25248
rect 2731 25245 2743 25279
rect 2685 25239 2743 25245
rect 2774 25236 2780 25288
rect 2832 25236 2838 25288
rect 3160 25208 3188 25375
rect 3694 25372 3700 25424
rect 3752 25412 3758 25424
rect 4433 25415 4491 25421
rect 4433 25412 4445 25415
rect 3752 25384 4445 25412
rect 3752 25372 3758 25384
rect 4433 25381 4445 25384
rect 4479 25381 4491 25415
rect 4540 25412 4568 25452
rect 4614 25440 4620 25492
rect 4672 25440 4678 25492
rect 4798 25440 4804 25492
rect 4856 25440 4862 25492
rect 5534 25440 5540 25492
rect 5592 25480 5598 25492
rect 6457 25483 6515 25489
rect 6457 25480 6469 25483
rect 5592 25452 6469 25480
rect 5592 25440 5598 25452
rect 6457 25449 6469 25452
rect 6503 25449 6515 25483
rect 6457 25443 6515 25449
rect 6914 25440 6920 25492
rect 6972 25440 6978 25492
rect 7282 25440 7288 25492
rect 7340 25440 7346 25492
rect 7650 25440 7656 25492
rect 7708 25480 7714 25492
rect 8478 25480 8484 25492
rect 7708 25452 8484 25480
rect 7708 25440 7714 25452
rect 8478 25440 8484 25452
rect 8536 25440 8542 25492
rect 8570 25440 8576 25492
rect 8628 25440 8634 25492
rect 8846 25440 8852 25492
rect 8904 25480 8910 25492
rect 8941 25483 8999 25489
rect 8941 25480 8953 25483
rect 8904 25452 8953 25480
rect 8904 25440 8910 25452
rect 8941 25449 8953 25452
rect 8987 25449 8999 25483
rect 8941 25443 8999 25449
rect 9490 25440 9496 25492
rect 9548 25480 9554 25492
rect 9766 25480 9772 25492
rect 9548 25452 9772 25480
rect 9548 25440 9554 25452
rect 9766 25440 9772 25452
rect 9824 25440 9830 25492
rect 6178 25412 6184 25424
rect 4540 25384 4629 25412
rect 4433 25375 4491 25381
rect 3418 25304 3424 25356
rect 3476 25304 3482 25356
rect 3789 25347 3847 25353
rect 3789 25344 3801 25347
rect 3712 25316 3801 25344
rect 3712 25288 3740 25316
rect 3789 25313 3801 25316
rect 3835 25313 3847 25347
rect 3789 25307 3847 25313
rect 3970 25304 3976 25356
rect 4028 25304 4034 25356
rect 4153 25349 4211 25355
rect 4153 25346 4165 25349
rect 4152 25315 4165 25346
rect 4199 25315 4211 25349
rect 4321 25347 4379 25353
rect 4321 25344 4333 25347
rect 4152 25309 4211 25315
rect 4264 25316 4333 25344
rect 3237 25279 3295 25285
rect 3237 25245 3249 25279
rect 3283 25276 3295 25279
rect 3602 25276 3608 25288
rect 3283 25248 3608 25276
rect 3283 25245 3295 25248
rect 3237 25239 3295 25245
rect 3602 25236 3608 25248
rect 3660 25236 3666 25288
rect 3694 25236 3700 25288
rect 3752 25236 3758 25288
rect 4065 25279 4123 25285
rect 4065 25245 4077 25279
rect 4111 25245 4123 25279
rect 4065 25239 4123 25245
rect 4080 25208 4108 25239
rect 2056 25180 2452 25208
rect 3160 25180 4108 25208
rect 4152 25220 4180 25309
rect 4264 25276 4292 25316
rect 4321 25313 4333 25316
rect 4367 25313 4379 25347
rect 4601 25350 4629 25384
rect 4908 25384 6184 25412
rect 4693 25353 4751 25359
rect 4693 25350 4705 25353
rect 4601 25322 4705 25350
rect 4693 25319 4705 25322
rect 4739 25319 4751 25353
rect 4693 25313 4751 25319
rect 4321 25307 4379 25313
rect 4908 25288 4936 25384
rect 6178 25372 6184 25384
rect 6236 25372 6242 25424
rect 6730 25372 6736 25424
rect 6788 25412 6794 25424
rect 6932 25412 6960 25440
rect 6788 25384 6960 25412
rect 7300 25412 7328 25440
rect 8588 25412 8616 25440
rect 9585 25415 9643 25421
rect 9585 25412 9597 25415
rect 7300 25390 7880 25412
rect 7300 25384 7656 25390
rect 6788 25372 6794 25384
rect 5077 25347 5135 25353
rect 5077 25313 5089 25347
rect 5123 25313 5135 25347
rect 5077 25307 5135 25313
rect 4614 25276 4620 25288
rect 4264 25248 4620 25276
rect 4614 25236 4620 25248
rect 4672 25236 4678 25288
rect 4801 25279 4859 25285
rect 4801 25245 4813 25279
rect 4847 25276 4859 25279
rect 4890 25276 4896 25288
rect 4847 25248 4896 25276
rect 4847 25245 4859 25248
rect 4801 25239 4859 25245
rect 4890 25236 4896 25248
rect 4948 25236 4954 25288
rect 5092 25276 5120 25307
rect 5350 25304 5356 25356
rect 5408 25344 5414 25356
rect 5997 25347 6055 25353
rect 5997 25344 6009 25347
rect 5408 25316 6009 25344
rect 5408 25304 5414 25316
rect 5997 25313 6009 25316
rect 6043 25313 6055 25347
rect 5997 25307 6055 25313
rect 6270 25304 6276 25356
rect 6328 25304 6334 25356
rect 6638 25304 6644 25356
rect 6696 25304 6702 25356
rect 6932 25353 6960 25384
rect 6825 25347 6883 25353
rect 6825 25344 6837 25347
rect 6822 25334 6837 25344
rect 6794 25313 6837 25334
rect 6871 25313 6883 25347
rect 6794 25307 6883 25313
rect 6917 25347 6975 25353
rect 6917 25313 6929 25347
rect 6963 25313 6975 25347
rect 6917 25307 6975 25313
rect 6794 25306 6850 25307
rect 5629 25279 5687 25285
rect 5092 25248 5396 25276
rect 5368 25220 5396 25248
rect 5629 25245 5641 25279
rect 5675 25276 5687 25279
rect 6288 25276 6316 25304
rect 5675 25248 6316 25276
rect 5675 25245 5687 25248
rect 5629 25239 5687 25245
rect 6546 25236 6552 25288
rect 6604 25236 6610 25288
rect 4152 25180 4160 25220
rect 1394 25100 1400 25152
rect 1452 25140 1458 25152
rect 2317 25143 2375 25149
rect 2317 25140 2329 25143
rect 1452 25112 2329 25140
rect 1452 25100 1458 25112
rect 2317 25109 2329 25112
rect 2363 25109 2375 25143
rect 2424 25140 2452 25180
rect 4154 25168 4160 25180
rect 4212 25168 4218 25220
rect 5169 25211 5227 25217
rect 5169 25208 5181 25211
rect 4356 25180 5181 25208
rect 4356 25140 4384 25180
rect 5169 25177 5181 25180
rect 5215 25177 5227 25211
rect 5169 25171 5227 25177
rect 5350 25168 5356 25220
rect 5408 25168 5414 25220
rect 5537 25211 5595 25217
rect 5537 25177 5549 25211
rect 5583 25208 5595 25211
rect 5583 25180 6100 25208
rect 5583 25177 5595 25180
rect 5537 25171 5595 25177
rect 2424 25112 4384 25140
rect 2317 25103 2375 25109
rect 4430 25100 4436 25152
rect 4488 25100 4494 25152
rect 4982 25100 4988 25152
rect 5040 25100 5046 25152
rect 5813 25143 5871 25149
rect 5813 25109 5825 25143
rect 5859 25140 5871 25143
rect 5902 25140 5908 25152
rect 5859 25112 5908 25140
rect 5859 25109 5871 25112
rect 5813 25103 5871 25109
rect 5902 25100 5908 25112
rect 5960 25100 5966 25152
rect 6072 25140 6100 25180
rect 6178 25168 6184 25220
rect 6236 25168 6242 25220
rect 6564 25208 6592 25236
rect 6288 25180 6592 25208
rect 6794 25208 6822 25306
rect 7006 25304 7012 25356
rect 7064 25304 7070 25356
rect 7190 25304 7196 25356
rect 7248 25304 7254 25356
rect 7469 25347 7527 25353
rect 7469 25313 7481 25347
rect 7515 25344 7527 25347
rect 7558 25344 7564 25356
rect 7515 25316 7564 25344
rect 7515 25313 7527 25316
rect 7469 25307 7527 25313
rect 7558 25304 7564 25316
rect 7616 25304 7622 25356
rect 7650 25338 7656 25384
rect 7708 25384 7880 25390
rect 8588 25384 9597 25412
rect 7708 25338 7714 25384
rect 7742 25304 7748 25356
rect 7800 25304 7806 25356
rect 7852 25353 7880 25384
rect 9585 25381 9597 25384
rect 9631 25381 9643 25415
rect 9585 25375 9643 25381
rect 7837 25347 7895 25353
rect 7837 25313 7849 25347
rect 7883 25313 7895 25347
rect 7837 25307 7895 25313
rect 8021 25347 8079 25353
rect 8021 25313 8033 25347
rect 8067 25344 8079 25347
rect 8386 25344 8392 25356
rect 8067 25316 8392 25344
rect 8067 25313 8079 25316
rect 8021 25307 8079 25313
rect 8386 25304 8392 25316
rect 8444 25304 8450 25356
rect 8481 25347 8539 25353
rect 8481 25313 8493 25347
rect 8527 25344 8539 25347
rect 8570 25344 8576 25356
rect 8527 25316 8576 25344
rect 8527 25313 8539 25316
rect 8481 25307 8539 25313
rect 8570 25304 8576 25316
rect 8628 25304 8634 25356
rect 9122 25304 9128 25356
rect 9180 25304 9186 25356
rect 9217 25347 9275 25353
rect 9217 25313 9229 25347
rect 9263 25344 9275 25347
rect 10502 25344 10508 25356
rect 9263 25316 10508 25344
rect 9263 25313 9275 25316
rect 9217 25307 9275 25313
rect 10502 25304 10508 25316
rect 10560 25304 10566 25356
rect 7374 25236 7380 25288
rect 7432 25276 7438 25288
rect 7653 25279 7711 25285
rect 7653 25276 7665 25279
rect 7432 25248 7665 25276
rect 7432 25236 7438 25248
rect 7653 25245 7665 25248
rect 7699 25245 7711 25279
rect 7653 25239 7711 25245
rect 8665 25279 8723 25285
rect 8665 25245 8677 25279
rect 8711 25245 8723 25279
rect 8665 25239 8723 25245
rect 7285 25211 7343 25217
rect 7285 25208 7297 25211
rect 6794 25180 7297 25208
rect 6288 25140 6316 25180
rect 7285 25177 7297 25180
rect 7331 25208 7343 25211
rect 7926 25208 7932 25220
rect 7331 25180 7932 25208
rect 7331 25177 7343 25180
rect 7285 25171 7343 25177
rect 7926 25168 7932 25180
rect 7984 25168 7990 25220
rect 8018 25168 8024 25220
rect 8076 25208 8082 25220
rect 8680 25208 8708 25239
rect 8754 25236 8760 25288
rect 8812 25276 8818 25288
rect 9493 25279 9551 25285
rect 9493 25276 9505 25279
rect 8812 25248 9505 25276
rect 8812 25236 8818 25248
rect 9493 25245 9505 25248
rect 9539 25245 9551 25279
rect 9493 25239 9551 25245
rect 10137 25279 10195 25285
rect 10137 25245 10149 25279
rect 10183 25245 10195 25279
rect 10137 25239 10195 25245
rect 8076 25180 8708 25208
rect 8076 25168 8082 25180
rect 9122 25168 9128 25220
rect 9180 25208 9186 25220
rect 10042 25208 10048 25220
rect 9180 25180 10048 25208
rect 9180 25168 9186 25180
rect 10042 25168 10048 25180
rect 10100 25208 10106 25220
rect 10152 25208 10180 25239
rect 10100 25180 10180 25208
rect 10100 25168 10106 25180
rect 6072 25112 6316 25140
rect 7650 25100 7656 25152
rect 7708 25140 7714 25152
rect 8113 25143 8171 25149
rect 8113 25140 8125 25143
rect 7708 25112 8125 25140
rect 7708 25100 7714 25112
rect 8113 25109 8125 25112
rect 8159 25109 8171 25143
rect 8113 25103 8171 25109
rect 10781 25143 10839 25149
rect 10781 25109 10793 25143
rect 10827 25140 10839 25143
rect 11054 25140 11060 25152
rect 10827 25112 11060 25140
rect 10827 25109 10839 25112
rect 10781 25103 10839 25109
rect 11054 25100 11060 25112
rect 11112 25100 11118 25152
rect 552 25050 11132 25072
rect 552 24998 3662 25050
rect 3714 24998 3726 25050
rect 3778 24998 3790 25050
rect 3842 24998 3854 25050
rect 3906 24998 3918 25050
rect 3970 24998 10062 25050
rect 10114 24998 10126 25050
rect 10178 24998 10190 25050
rect 10242 24998 10254 25050
rect 10306 24998 10318 25050
rect 10370 24998 11132 25050
rect 552 24976 11132 24998
rect 1302 24896 1308 24948
rect 1360 24936 1366 24948
rect 3237 24939 3295 24945
rect 3237 24936 3249 24939
rect 1360 24908 3249 24936
rect 1360 24896 1366 24908
rect 3237 24905 3249 24908
rect 3283 24905 3295 24939
rect 3237 24899 3295 24905
rect 3418 24896 3424 24948
rect 3476 24936 3482 24948
rect 3970 24936 3976 24948
rect 3476 24908 3976 24936
rect 3476 24896 3482 24908
rect 3970 24896 3976 24908
rect 4028 24936 4034 24948
rect 4065 24939 4123 24945
rect 4065 24936 4077 24939
rect 4028 24908 4077 24936
rect 4028 24896 4034 24908
rect 4065 24905 4077 24908
rect 4111 24905 4123 24939
rect 4065 24899 4123 24905
rect 4154 24896 4160 24948
rect 4212 24936 4218 24948
rect 4798 24936 4804 24948
rect 4212 24908 4804 24936
rect 4212 24896 4218 24908
rect 4798 24896 4804 24908
rect 4856 24896 4862 24948
rect 5258 24936 5264 24948
rect 4908 24908 5264 24936
rect 1949 24871 2007 24877
rect 1949 24837 1961 24871
rect 1995 24868 2007 24871
rect 1995 24840 2728 24868
rect 1995 24837 2007 24840
rect 1949 24831 2007 24837
rect 1394 24760 1400 24812
rect 1452 24760 1458 24812
rect 1486 24760 1492 24812
rect 1544 24760 1550 24812
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24800 1731 24803
rect 2498 24800 2504 24812
rect 1719 24772 2504 24800
rect 1719 24769 1731 24772
rect 1673 24763 1731 24769
rect 2498 24760 2504 24772
rect 2556 24760 2562 24812
rect 1412 24732 1440 24760
rect 1765 24735 1823 24741
rect 1412 24704 1716 24732
rect 658 24624 664 24676
rect 716 24664 722 24676
rect 1486 24664 1492 24676
rect 716 24636 1492 24664
rect 716 24624 722 24636
rect 1486 24624 1492 24636
rect 1544 24624 1550 24676
rect 1688 24664 1716 24704
rect 1765 24701 1777 24735
rect 1811 24732 1823 24735
rect 2133 24735 2191 24741
rect 2133 24732 2145 24735
rect 1811 24704 2145 24732
rect 1811 24701 1823 24704
rect 1765 24695 1823 24701
rect 2133 24701 2145 24704
rect 2179 24732 2191 24735
rect 2222 24732 2228 24744
rect 2179 24704 2228 24732
rect 2179 24701 2191 24704
rect 2133 24695 2191 24701
rect 2222 24692 2228 24704
rect 2280 24692 2286 24744
rect 2406 24692 2412 24744
rect 2464 24692 2470 24744
rect 2700 24741 2728 24840
rect 2774 24828 2780 24880
rect 2832 24868 2838 24880
rect 4706 24868 4712 24880
rect 2832 24840 4712 24868
rect 2832 24828 2838 24840
rect 4706 24828 4712 24840
rect 4764 24828 4770 24880
rect 3513 24803 3571 24809
rect 3513 24769 3525 24803
rect 3559 24800 3571 24803
rect 4614 24800 4620 24812
rect 3559 24772 4620 24800
rect 3559 24769 3571 24772
rect 3513 24763 3571 24769
rect 4614 24760 4620 24772
rect 4672 24760 4678 24812
rect 4908 24800 4936 24908
rect 5258 24896 5264 24908
rect 5316 24936 5322 24948
rect 6454 24936 6460 24948
rect 5316 24908 6460 24936
rect 5316 24896 5322 24908
rect 6454 24896 6460 24908
rect 6512 24896 6518 24948
rect 7006 24896 7012 24948
rect 7064 24936 7070 24948
rect 8205 24939 8263 24945
rect 8205 24936 8217 24939
rect 7064 24908 8217 24936
rect 7064 24896 7070 24908
rect 8205 24905 8217 24908
rect 8251 24905 8263 24939
rect 8205 24899 8263 24905
rect 4982 24828 4988 24880
rect 5040 24828 5046 24880
rect 5534 24828 5540 24880
rect 5592 24868 5598 24880
rect 5592 24840 6040 24868
rect 5592 24828 5598 24840
rect 4724 24772 4936 24800
rect 5000 24800 5028 24828
rect 5718 24800 5724 24812
rect 5000 24772 5724 24800
rect 2593 24735 2651 24741
rect 2593 24701 2605 24735
rect 2639 24701 2651 24735
rect 2593 24695 2651 24701
rect 2685 24735 2743 24741
rect 2685 24701 2697 24735
rect 2731 24701 2743 24735
rect 2685 24695 2743 24701
rect 3237 24735 3295 24741
rect 3237 24701 3249 24735
rect 3283 24732 3295 24735
rect 3326 24732 3332 24744
rect 3283 24704 3332 24732
rect 3283 24701 3295 24704
rect 3237 24695 3295 24701
rect 2608 24664 2636 24695
rect 3326 24692 3332 24704
rect 3384 24692 3390 24744
rect 3418 24692 3424 24744
rect 3476 24732 3482 24744
rect 3476 24704 3648 24732
rect 3476 24692 3482 24704
rect 1688 24636 2636 24664
rect 2774 24624 2780 24676
rect 2832 24664 2838 24676
rect 2869 24667 2927 24673
rect 2869 24664 2881 24667
rect 2832 24636 2881 24664
rect 2832 24624 2838 24636
rect 2869 24633 2881 24636
rect 2915 24633 2927 24667
rect 3620 24664 3648 24704
rect 3694 24692 3700 24744
rect 3752 24692 3758 24744
rect 4062 24732 4068 24744
rect 3804 24704 4068 24732
rect 3804 24664 3832 24704
rect 4062 24692 4068 24704
rect 4120 24692 4126 24744
rect 4154 24692 4160 24744
rect 4212 24732 4218 24744
rect 4724 24741 4752 24772
rect 5718 24760 5724 24772
rect 5776 24760 5782 24812
rect 6012 24800 6040 24840
rect 6270 24828 6276 24880
rect 6328 24868 6334 24880
rect 7837 24871 7895 24877
rect 7837 24868 7849 24871
rect 6328 24840 7849 24868
rect 6328 24828 6334 24840
rect 7837 24837 7849 24840
rect 7883 24837 7895 24871
rect 8570 24868 8576 24880
rect 7837 24831 7895 24837
rect 8128 24840 8576 24868
rect 6012 24772 7604 24800
rect 4249 24735 4307 24741
rect 4249 24732 4261 24735
rect 4212 24704 4261 24732
rect 4212 24692 4218 24704
rect 4249 24701 4261 24704
rect 4295 24701 4307 24735
rect 4249 24695 4307 24701
rect 4709 24735 4767 24741
rect 4709 24701 4721 24735
rect 4755 24701 4767 24735
rect 4709 24695 4767 24701
rect 4798 24692 4804 24744
rect 4856 24692 4862 24744
rect 4985 24735 5043 24741
rect 4985 24701 4997 24735
rect 5031 24701 5043 24735
rect 4985 24695 5043 24701
rect 5169 24735 5227 24741
rect 5169 24701 5181 24735
rect 5215 24732 5227 24735
rect 5626 24732 5632 24744
rect 5215 24729 5488 24732
rect 5552 24729 5632 24732
rect 5215 24704 5632 24729
rect 5215 24701 5227 24704
rect 5460 24701 5580 24704
rect 5169 24695 5227 24701
rect 3620 24636 3832 24664
rect 2869 24627 2927 24633
rect 3878 24624 3884 24676
rect 3936 24664 3942 24676
rect 4525 24667 4583 24673
rect 4525 24664 4537 24667
rect 3936 24636 4537 24664
rect 3936 24624 3942 24636
rect 4525 24633 4537 24636
rect 4571 24633 4583 24667
rect 5000 24664 5028 24695
rect 5626 24692 5632 24704
rect 5684 24692 5690 24744
rect 6012 24741 6040 24772
rect 5905 24735 5963 24741
rect 5905 24701 5917 24735
rect 5951 24701 5963 24735
rect 5905 24695 5963 24701
rect 5997 24735 6055 24741
rect 5997 24701 6009 24735
rect 6043 24701 6055 24735
rect 6825 24735 6883 24741
rect 6825 24732 6837 24735
rect 5997 24695 6055 24701
rect 6288 24704 6837 24732
rect 5261 24667 5319 24673
rect 5261 24664 5273 24667
rect 5000 24636 5273 24664
rect 4525 24627 4583 24633
rect 5261 24633 5273 24636
rect 5307 24664 5319 24667
rect 5350 24664 5356 24676
rect 5307 24636 5356 24664
rect 5307 24633 5319 24636
rect 5261 24627 5319 24633
rect 5350 24624 5356 24636
rect 5408 24624 5414 24676
rect 5445 24667 5503 24673
rect 5445 24633 5457 24667
rect 5491 24664 5503 24667
rect 5718 24664 5724 24676
rect 5491 24636 5724 24664
rect 5491 24633 5503 24636
rect 5445 24627 5503 24633
rect 5718 24624 5724 24636
rect 5776 24624 5782 24676
rect 5920 24664 5948 24695
rect 6288 24676 6316 24704
rect 6825 24701 6837 24704
rect 6871 24701 6883 24735
rect 6825 24695 6883 24701
rect 7101 24735 7159 24741
rect 7101 24701 7113 24735
rect 7147 24701 7159 24735
rect 7101 24695 7159 24701
rect 6270 24664 6276 24676
rect 5920 24636 6276 24664
rect 6270 24624 6276 24636
rect 6328 24624 6334 24676
rect 7116 24664 7144 24695
rect 7190 24692 7196 24744
rect 7248 24692 7254 24744
rect 7282 24692 7288 24744
rect 7340 24732 7346 24744
rect 7377 24735 7435 24741
rect 7377 24732 7389 24735
rect 7340 24704 7389 24732
rect 7340 24692 7346 24704
rect 7377 24701 7389 24704
rect 7423 24701 7435 24735
rect 7377 24695 7435 24701
rect 7466 24692 7472 24744
rect 7524 24692 7530 24744
rect 7576 24741 7604 24772
rect 7561 24735 7619 24741
rect 7561 24701 7573 24735
rect 7607 24701 7619 24735
rect 7561 24695 7619 24701
rect 7650 24692 7656 24744
rect 7708 24732 7714 24744
rect 7834 24732 7840 24744
rect 7708 24704 7840 24732
rect 7708 24692 7714 24704
rect 7834 24692 7840 24704
rect 7892 24692 7898 24744
rect 7926 24692 7932 24744
rect 7984 24692 7990 24744
rect 8021 24735 8079 24741
rect 8021 24701 8033 24735
rect 8067 24732 8079 24735
rect 8128 24732 8156 24840
rect 8570 24828 8576 24840
rect 8628 24868 8634 24880
rect 8846 24868 8852 24880
rect 8628 24840 8852 24868
rect 8628 24828 8634 24840
rect 8846 24828 8852 24840
rect 8904 24828 8910 24880
rect 9674 24828 9680 24880
rect 9732 24868 9738 24880
rect 10226 24868 10232 24880
rect 9732 24840 10232 24868
rect 9732 24828 9738 24840
rect 10226 24828 10232 24840
rect 10284 24828 10290 24880
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 8757 24803 8815 24809
rect 8757 24800 8769 24803
rect 8444 24772 8769 24800
rect 8444 24760 8450 24772
rect 8757 24769 8769 24772
rect 8803 24769 8815 24803
rect 8757 24763 8815 24769
rect 10318 24760 10324 24812
rect 10376 24760 10382 24812
rect 10502 24760 10508 24812
rect 10560 24800 10566 24812
rect 10560 24772 10824 24800
rect 10560 24760 10566 24772
rect 8067 24704 8156 24732
rect 8205 24735 8263 24741
rect 8067 24701 8079 24704
rect 8021 24695 8079 24701
rect 8205 24701 8217 24735
rect 8251 24732 8263 24735
rect 9674 24732 9680 24744
rect 8251 24704 9680 24732
rect 8251 24701 8263 24704
rect 8205 24695 8263 24701
rect 9674 24692 9680 24704
rect 9732 24692 9738 24744
rect 10042 24692 10048 24744
rect 10100 24692 10106 24744
rect 10594 24692 10600 24744
rect 10652 24692 10658 24744
rect 10796 24741 10824 24772
rect 10781 24735 10839 24741
rect 10781 24701 10793 24735
rect 10827 24701 10839 24735
rect 10781 24695 10839 24701
rect 7116 24636 8156 24664
rect 8128 24608 8156 24636
rect 8386 24624 8392 24676
rect 8444 24624 8450 24676
rect 8478 24624 8484 24676
rect 8536 24664 8542 24676
rect 8573 24667 8631 24673
rect 8573 24664 8585 24667
rect 8536 24636 8585 24664
rect 8536 24624 8542 24636
rect 8573 24633 8585 24636
rect 8619 24633 8631 24667
rect 8573 24627 8631 24633
rect 8662 24624 8668 24676
rect 8720 24664 8726 24676
rect 9033 24667 9091 24673
rect 9033 24664 9045 24667
rect 8720 24636 9045 24664
rect 8720 24624 8726 24636
rect 9033 24633 9045 24636
rect 9079 24633 9091 24667
rect 9033 24627 9091 24633
rect 9214 24624 9220 24676
rect 9272 24624 9278 24676
rect 9582 24624 9588 24676
rect 9640 24664 9646 24676
rect 10134 24664 10140 24676
rect 9640 24636 10140 24664
rect 9640 24624 9646 24636
rect 10134 24624 10140 24636
rect 10192 24624 10198 24676
rect 10502 24624 10508 24676
rect 10560 24664 10566 24676
rect 10962 24664 10968 24676
rect 10560 24636 10968 24664
rect 10560 24624 10566 24636
rect 10962 24624 10968 24636
rect 11020 24624 11026 24676
rect 382 24556 388 24608
rect 440 24596 446 24608
rect 1305 24599 1363 24605
rect 1305 24596 1317 24599
rect 440 24568 1317 24596
rect 440 24556 446 24568
rect 1305 24565 1317 24568
rect 1351 24565 1363 24599
rect 1305 24559 1363 24565
rect 2317 24599 2375 24605
rect 2317 24565 2329 24599
rect 2363 24596 2375 24599
rect 2498 24596 2504 24608
rect 2363 24568 2504 24596
rect 2363 24565 2375 24568
rect 2317 24559 2375 24565
rect 2498 24556 2504 24568
rect 2556 24556 2562 24608
rect 2590 24556 2596 24608
rect 2648 24596 2654 24608
rect 4982 24596 4988 24608
rect 2648 24568 4988 24596
rect 2648 24556 2654 24568
rect 4982 24556 4988 24568
rect 5040 24556 5046 24608
rect 5074 24556 5080 24608
rect 5132 24556 5138 24608
rect 5626 24556 5632 24608
rect 5684 24596 5690 24608
rect 5994 24596 6000 24608
rect 5684 24568 6000 24596
rect 5684 24556 5690 24568
rect 5994 24556 6000 24568
rect 6052 24556 6058 24608
rect 6181 24599 6239 24605
rect 6181 24565 6193 24599
rect 6227 24596 6239 24599
rect 6546 24596 6552 24608
rect 6227 24568 6552 24596
rect 6227 24565 6239 24568
rect 6181 24559 6239 24565
rect 6546 24556 6552 24568
rect 6604 24556 6610 24608
rect 7374 24556 7380 24608
rect 7432 24596 7438 24608
rect 7650 24596 7656 24608
rect 7432 24568 7656 24596
rect 7432 24556 7438 24568
rect 7650 24556 7656 24568
rect 7708 24556 7714 24608
rect 8110 24556 8116 24608
rect 8168 24596 8174 24608
rect 8849 24599 8907 24605
rect 8849 24596 8861 24599
rect 8168 24568 8861 24596
rect 8168 24556 8174 24568
rect 8849 24565 8861 24568
rect 8895 24565 8907 24599
rect 8849 24559 8907 24565
rect 9306 24556 9312 24608
rect 9364 24596 9370 24608
rect 9401 24599 9459 24605
rect 9401 24596 9413 24599
rect 9364 24568 9413 24596
rect 9364 24556 9370 24568
rect 9401 24565 9413 24568
rect 9447 24565 9459 24599
rect 9401 24559 9459 24565
rect 9490 24556 9496 24608
rect 9548 24596 9554 24608
rect 10689 24599 10747 24605
rect 10689 24596 10701 24599
rect 9548 24568 10701 24596
rect 9548 24556 9554 24568
rect 10689 24565 10701 24568
rect 10735 24565 10747 24599
rect 10689 24559 10747 24565
rect 552 24506 11132 24528
rect 552 24454 4322 24506
rect 4374 24454 4386 24506
rect 4438 24454 4450 24506
rect 4502 24454 4514 24506
rect 4566 24454 4578 24506
rect 4630 24454 10722 24506
rect 10774 24454 10786 24506
rect 10838 24454 10850 24506
rect 10902 24454 10914 24506
rect 10966 24454 10978 24506
rect 11030 24454 11132 24506
rect 552 24432 11132 24454
rect 106 24352 112 24404
rect 164 24392 170 24404
rect 658 24392 664 24404
rect 164 24364 664 24392
rect 164 24352 170 24364
rect 658 24352 664 24364
rect 716 24352 722 24404
rect 1026 24352 1032 24404
rect 1084 24392 1090 24404
rect 1084 24364 2820 24392
rect 1084 24352 1090 24364
rect 1213 24327 1271 24333
rect 1213 24293 1225 24327
rect 1259 24324 1271 24327
rect 1394 24324 1400 24336
rect 1259 24296 1400 24324
rect 1259 24293 1271 24296
rect 1213 24287 1271 24293
rect 1394 24284 1400 24296
rect 1452 24284 1458 24336
rect 2792 24324 2820 24364
rect 3878 24352 3884 24404
rect 3936 24392 3942 24404
rect 4522 24392 4528 24404
rect 3936 24364 4528 24392
rect 3936 24352 3942 24364
rect 4522 24352 4528 24364
rect 4580 24352 4586 24404
rect 6273 24395 6331 24401
rect 5460 24364 6224 24392
rect 2792 24296 3096 24324
rect 1302 24216 1308 24268
rect 1360 24256 1366 24268
rect 1762 24256 1768 24268
rect 1360 24228 1768 24256
rect 1360 24216 1366 24228
rect 1762 24216 1768 24228
rect 1820 24216 1826 24268
rect 2041 24259 2099 24265
rect 2041 24225 2053 24259
rect 2087 24256 2099 24259
rect 2317 24259 2375 24265
rect 2317 24256 2329 24259
rect 2087 24228 2329 24256
rect 2087 24225 2099 24228
rect 2041 24219 2099 24225
rect 2317 24225 2329 24228
rect 2363 24225 2375 24259
rect 2317 24219 2375 24225
rect 2498 24216 2504 24268
rect 2556 24216 2562 24268
rect 2590 24216 2596 24268
rect 2648 24256 2654 24268
rect 3068 24265 3096 24296
rect 3326 24284 3332 24336
rect 3384 24324 3390 24336
rect 3973 24327 4031 24333
rect 3973 24324 3985 24327
rect 3384 24296 3985 24324
rect 3384 24284 3390 24296
rect 3973 24293 3985 24296
rect 4019 24293 4031 24327
rect 3973 24287 4031 24293
rect 4062 24284 4068 24336
rect 4120 24324 4126 24336
rect 4157 24327 4215 24333
rect 4157 24324 4169 24327
rect 4120 24296 4169 24324
rect 4120 24284 4126 24296
rect 4157 24293 4169 24296
rect 4203 24293 4215 24327
rect 4157 24287 4215 24293
rect 4617 24327 4675 24333
rect 4617 24293 4629 24327
rect 4663 24324 4675 24327
rect 4706 24324 4712 24336
rect 4663 24296 4712 24324
rect 4663 24293 4675 24296
rect 4617 24287 4675 24293
rect 4706 24284 4712 24296
rect 4764 24284 4770 24336
rect 5258 24284 5264 24336
rect 5316 24284 5322 24336
rect 5350 24284 5356 24336
rect 5408 24284 5414 24336
rect 5460 24333 5488 24364
rect 5460 24327 5529 24333
rect 5460 24296 5483 24327
rect 5471 24293 5483 24296
rect 5517 24293 5529 24327
rect 6196 24324 6224 24364
rect 6273 24361 6285 24395
rect 6319 24392 6331 24395
rect 6638 24392 6644 24404
rect 6319 24364 6644 24392
rect 6319 24361 6331 24364
rect 6273 24355 6331 24361
rect 6638 24352 6644 24364
rect 6696 24352 6702 24404
rect 6914 24352 6920 24404
rect 6972 24352 6978 24404
rect 7006 24352 7012 24404
rect 7064 24392 7070 24404
rect 7837 24395 7895 24401
rect 7837 24392 7849 24395
rect 7064 24364 7849 24392
rect 7064 24352 7070 24364
rect 7837 24361 7849 24364
rect 7883 24392 7895 24395
rect 7883 24364 8340 24392
rect 7883 24361 7895 24364
rect 7837 24355 7895 24361
rect 6362 24324 6368 24336
rect 6196 24296 6368 24324
rect 5471 24287 5529 24293
rect 6362 24284 6368 24296
rect 6420 24284 6426 24336
rect 7024 24302 8064 24324
rect 7024 24296 7288 24302
rect 2869 24259 2927 24265
rect 2869 24256 2881 24259
rect 2648 24228 2881 24256
rect 2648 24216 2654 24228
rect 2869 24225 2881 24228
rect 2915 24225 2927 24259
rect 2869 24219 2927 24225
rect 3053 24259 3111 24265
rect 3053 24225 3065 24259
rect 3099 24256 3111 24259
rect 3510 24256 3516 24268
rect 3099 24228 3516 24256
rect 3099 24225 3111 24228
rect 3053 24219 3111 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 4080 24256 4108 24284
rect 7024 24268 7052 24296
rect 3620 24228 4108 24256
rect 2222 24148 2228 24200
rect 2280 24148 2286 24200
rect 2777 24191 2835 24197
rect 2777 24157 2789 24191
rect 2823 24188 2835 24191
rect 2958 24188 2964 24200
rect 2823 24160 2964 24188
rect 2823 24157 2835 24160
rect 2777 24151 2835 24157
rect 2958 24148 2964 24160
rect 3016 24148 3022 24200
rect 3145 24191 3203 24197
rect 3145 24157 3157 24191
rect 3191 24188 3203 24191
rect 3326 24188 3332 24200
rect 3191 24160 3332 24188
rect 3191 24157 3203 24160
rect 3145 24151 3203 24157
rect 3326 24148 3332 24160
rect 3384 24148 3390 24200
rect 3620 24197 3648 24228
rect 4798 24216 4804 24268
rect 4856 24216 4862 24268
rect 5169 24259 5227 24265
rect 5169 24225 5181 24259
rect 5215 24256 5227 24259
rect 5215 24228 5322 24256
rect 5215 24225 5227 24228
rect 5169 24219 5227 24225
rect 3421 24191 3479 24197
rect 3421 24157 3433 24191
rect 3467 24157 3479 24191
rect 3421 24151 3479 24157
rect 3605 24191 3663 24197
rect 3605 24157 3617 24191
rect 3651 24157 3663 24191
rect 3605 24151 3663 24157
rect 842 24080 848 24132
rect 900 24120 906 24132
rect 900 24092 3004 24120
rect 900 24080 906 24092
rect 2590 24012 2596 24064
rect 2648 24052 2654 24064
rect 2685 24055 2743 24061
rect 2685 24052 2697 24055
rect 2648 24024 2697 24052
rect 2648 24012 2654 24024
rect 2685 24021 2697 24024
rect 2731 24021 2743 24055
rect 2976 24052 3004 24092
rect 3050 24080 3056 24132
rect 3108 24080 3114 24132
rect 3436 24120 3464 24151
rect 3694 24148 3700 24200
rect 3752 24188 3758 24200
rect 4062 24188 4068 24200
rect 3752 24160 4068 24188
rect 3752 24148 3758 24160
rect 4062 24148 4068 24160
rect 4120 24148 4126 24200
rect 4982 24188 4988 24200
rect 4264 24160 4988 24188
rect 3878 24120 3884 24132
rect 3436 24092 3884 24120
rect 3878 24080 3884 24092
rect 3936 24080 3942 24132
rect 3970 24080 3976 24132
rect 4028 24120 4034 24132
rect 4264 24120 4292 24160
rect 4982 24148 4988 24160
rect 5040 24148 5046 24200
rect 4028 24092 4292 24120
rect 4341 24123 4399 24129
rect 4028 24080 4034 24092
rect 4341 24089 4353 24123
rect 4387 24120 4399 24123
rect 4706 24120 4712 24132
rect 4387 24092 4712 24120
rect 4387 24089 4399 24092
rect 4341 24083 4399 24089
rect 4706 24080 4712 24092
rect 4764 24080 4770 24132
rect 5294 24120 5322 24228
rect 5368 24246 5949 24256
rect 5368 24228 6040 24246
rect 5368 24200 5396 24228
rect 5921 24218 6040 24228
rect 5350 24148 5356 24200
rect 5408 24148 5414 24200
rect 5629 24191 5687 24197
rect 5629 24157 5641 24191
rect 5675 24188 5687 24191
rect 6012 24188 6040 24218
rect 6178 24216 6184 24268
rect 6236 24216 6242 24268
rect 6546 24216 6552 24268
rect 6604 24256 6610 24268
rect 6825 24259 6883 24265
rect 6825 24256 6837 24259
rect 6604 24228 6837 24256
rect 6604 24216 6610 24228
rect 6825 24225 6837 24228
rect 6871 24225 6883 24259
rect 6825 24219 6883 24225
rect 7006 24216 7012 24268
rect 7064 24216 7070 24268
rect 7190 24216 7196 24268
rect 7248 24216 7254 24268
rect 7282 24250 7288 24296
rect 7340 24296 8064 24302
rect 7340 24250 7346 24296
rect 7377 24259 7435 24265
rect 7377 24225 7389 24259
rect 7423 24225 7435 24259
rect 7377 24219 7435 24225
rect 6086 24188 6092 24200
rect 5675 24160 5948 24188
rect 6012 24160 6092 24188
rect 5675 24157 5687 24160
rect 5629 24151 5687 24157
rect 5920 24132 5948 24160
rect 6086 24148 6092 24160
rect 6144 24148 6150 24200
rect 6362 24148 6368 24200
rect 6420 24148 6426 24200
rect 7282 24148 7288 24200
rect 7340 24188 7346 24200
rect 7392 24188 7420 24219
rect 7466 24216 7472 24268
rect 7524 24216 7530 24268
rect 8036 24265 8064 24296
rect 8312 24265 8340 24364
rect 8570 24352 8576 24404
rect 8628 24392 8634 24404
rect 9309 24395 9367 24401
rect 9309 24392 9321 24395
rect 8628 24364 9321 24392
rect 8628 24352 8634 24364
rect 9309 24361 9321 24364
rect 9355 24361 9367 24395
rect 9309 24355 9367 24361
rect 9858 24352 9864 24404
rect 9916 24392 9922 24404
rect 10137 24395 10195 24401
rect 10137 24392 10149 24395
rect 9916 24364 10149 24392
rect 9916 24352 9922 24364
rect 10137 24361 10149 24364
rect 10183 24361 10195 24395
rect 10137 24355 10195 24361
rect 10689 24395 10747 24401
rect 10689 24361 10701 24395
rect 10735 24392 10747 24395
rect 11238 24392 11244 24404
rect 10735 24364 11244 24392
rect 10735 24361 10747 24364
rect 10689 24355 10747 24361
rect 11238 24352 11244 24364
rect 11296 24352 11302 24404
rect 8938 24284 8944 24336
rect 8996 24284 9002 24336
rect 9030 24284 9036 24336
rect 9088 24284 9094 24336
rect 9766 24284 9772 24336
rect 9824 24324 9830 24336
rect 9824 24296 10824 24324
rect 9824 24284 9830 24296
rect 7653 24259 7711 24265
rect 7653 24225 7665 24259
rect 7699 24225 7711 24259
rect 7653 24219 7711 24225
rect 7745 24259 7803 24265
rect 7745 24225 7757 24259
rect 7791 24256 7803 24259
rect 8021 24259 8079 24265
rect 7791 24228 7972 24256
rect 7791 24225 7803 24228
rect 7745 24219 7803 24225
rect 7340 24160 7420 24188
rect 7668 24188 7696 24219
rect 7834 24188 7840 24200
rect 7668 24160 7840 24188
rect 7340 24148 7346 24160
rect 7834 24148 7840 24160
rect 7892 24148 7898 24200
rect 5813 24123 5871 24129
rect 5813 24120 5825 24123
rect 4804 24092 5212 24120
rect 5294 24092 5825 24120
rect 3602 24052 3608 24064
rect 2976 24024 3608 24052
rect 2685 24015 2743 24021
rect 3602 24012 3608 24024
rect 3660 24012 3666 24064
rect 4430 24012 4436 24064
rect 4488 24012 4494 24064
rect 4522 24012 4528 24064
rect 4580 24052 4586 24064
rect 4804 24052 4832 24092
rect 4580 24024 4832 24052
rect 4985 24055 5043 24061
rect 4580 24012 4586 24024
rect 4985 24021 4997 24055
rect 5031 24052 5043 24055
rect 5074 24052 5080 24064
rect 5031 24024 5080 24052
rect 5031 24021 5043 24024
rect 4985 24015 5043 24021
rect 5074 24012 5080 24024
rect 5132 24012 5138 24064
rect 5184 24052 5212 24092
rect 5813 24089 5825 24092
rect 5859 24089 5871 24123
rect 5813 24083 5871 24089
rect 5902 24080 5908 24132
rect 5960 24120 5966 24132
rect 6730 24120 6736 24132
rect 5960 24092 6736 24120
rect 5960 24080 5966 24092
rect 6730 24080 6736 24092
rect 6788 24120 6794 24132
rect 7944 24120 7972 24228
rect 8021 24225 8033 24259
rect 8067 24225 8079 24259
rect 8021 24219 8079 24225
rect 8297 24259 8355 24265
rect 8297 24225 8309 24259
rect 8343 24225 8355 24259
rect 8297 24219 8355 24225
rect 8665 24259 8723 24265
rect 8665 24225 8677 24259
rect 8711 24225 8723 24259
rect 8665 24219 8723 24225
rect 8205 24191 8263 24197
rect 8205 24188 8217 24191
rect 8128 24160 8217 24188
rect 8128 24132 8156 24160
rect 8205 24157 8217 24160
rect 8251 24157 8263 24191
rect 8680 24188 8708 24219
rect 8754 24216 8760 24268
rect 8812 24216 8818 24268
rect 9122 24216 9128 24268
rect 9180 24265 9186 24268
rect 9180 24259 9215 24265
rect 9203 24256 9215 24259
rect 9490 24256 9496 24268
rect 9203 24228 9496 24256
rect 9203 24225 9215 24228
rect 9180 24219 9215 24225
rect 9180 24216 9186 24219
rect 9490 24216 9496 24228
rect 9548 24216 9554 24268
rect 9582 24216 9588 24268
rect 9640 24256 9646 24268
rect 10229 24259 10287 24265
rect 10229 24256 10241 24259
rect 9640 24228 10241 24256
rect 9640 24216 9646 24228
rect 10229 24225 10241 24228
rect 10275 24225 10287 24259
rect 10229 24219 10287 24225
rect 10410 24216 10416 24268
rect 10468 24256 10474 24268
rect 10796 24265 10824 24296
rect 10597 24259 10655 24265
rect 10597 24256 10609 24259
rect 10468 24228 10609 24256
rect 10468 24216 10474 24228
rect 10597 24225 10609 24228
rect 10643 24225 10655 24259
rect 10597 24219 10655 24225
rect 10781 24259 10839 24265
rect 10781 24225 10793 24259
rect 10827 24225 10839 24259
rect 10781 24219 10839 24225
rect 8680 24160 9076 24188
rect 8205 24151 8263 24157
rect 9048 24132 9076 24160
rect 9306 24148 9312 24200
rect 9364 24188 9370 24200
rect 9677 24191 9735 24197
rect 9677 24188 9689 24191
rect 9364 24160 9689 24188
rect 9364 24148 9370 24160
rect 9677 24157 9689 24160
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 9769 24191 9827 24197
rect 9769 24157 9781 24191
rect 9815 24188 9827 24191
rect 9858 24188 9864 24200
rect 9815 24160 9864 24188
rect 9815 24157 9827 24160
rect 9769 24151 9827 24157
rect 9858 24148 9864 24160
rect 9916 24148 9922 24200
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 11238 24188 11244 24200
rect 10192 24160 11244 24188
rect 10192 24148 10198 24160
rect 11238 24148 11244 24160
rect 11296 24148 11302 24200
rect 6788 24092 7972 24120
rect 6788 24080 6794 24092
rect 8110 24080 8116 24132
rect 8168 24080 8174 24132
rect 8481 24123 8539 24129
rect 8481 24089 8493 24123
rect 8527 24120 8539 24123
rect 8846 24120 8852 24132
rect 8527 24092 8852 24120
rect 8527 24089 8539 24092
rect 8481 24083 8539 24089
rect 8846 24080 8852 24092
rect 8904 24080 8910 24132
rect 9030 24080 9036 24132
rect 9088 24080 9094 24132
rect 9232 24092 10456 24120
rect 9232 24064 9260 24092
rect 6362 24052 6368 24064
rect 5184 24024 6368 24052
rect 6362 24012 6368 24024
rect 6420 24052 6426 24064
rect 7282 24052 7288 24064
rect 6420 24024 7288 24052
rect 6420 24012 6426 24024
rect 7282 24012 7288 24024
rect 7340 24052 7346 24064
rect 8386 24052 8392 24064
rect 7340 24024 8392 24052
rect 7340 24012 7346 24024
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 9214 24012 9220 24064
rect 9272 24012 9278 24064
rect 9490 24012 9496 24064
rect 9548 24012 9554 24064
rect 9858 24012 9864 24064
rect 9916 24052 9922 24064
rect 10226 24052 10232 24064
rect 9916 24024 10232 24052
rect 9916 24012 9922 24024
rect 10226 24012 10232 24024
rect 10284 24012 10290 24064
rect 10428 24061 10456 24092
rect 10413 24055 10471 24061
rect 10413 24021 10425 24055
rect 10459 24052 10471 24055
rect 10594 24052 10600 24064
rect 10459 24024 10600 24052
rect 10459 24021 10471 24024
rect 10413 24015 10471 24021
rect 10594 24012 10600 24024
rect 10652 24012 10658 24064
rect 552 23962 11132 23984
rect 552 23910 3662 23962
rect 3714 23910 3726 23962
rect 3778 23910 3790 23962
rect 3842 23910 3854 23962
rect 3906 23910 3918 23962
rect 3970 23910 10062 23962
rect 10114 23910 10126 23962
rect 10178 23910 10190 23962
rect 10242 23910 10254 23962
rect 10306 23910 10318 23962
rect 10370 23910 11132 23962
rect 552 23888 11132 23910
rect 2406 23808 2412 23860
rect 2464 23848 2470 23860
rect 4157 23851 4215 23857
rect 4157 23848 4169 23851
rect 2464 23820 4169 23848
rect 2464 23808 2470 23820
rect 4157 23817 4169 23820
rect 4203 23817 4215 23851
rect 4157 23811 4215 23817
rect 5074 23808 5080 23860
rect 5132 23808 5138 23860
rect 5442 23808 5448 23860
rect 5500 23848 5506 23860
rect 5500 23820 6868 23848
rect 5500 23808 5506 23820
rect 2498 23740 2504 23792
rect 2556 23780 2562 23792
rect 2685 23783 2743 23789
rect 2556 23752 2655 23780
rect 2556 23740 2562 23752
rect 1762 23672 1768 23724
rect 1820 23672 1826 23724
rect 2317 23715 2375 23721
rect 2317 23712 2329 23715
rect 2056 23684 2329 23712
rect 2056 23653 2084 23684
rect 2317 23681 2329 23684
rect 2363 23681 2375 23715
rect 2317 23675 2375 23681
rect 2627 23712 2655 23752
rect 2685 23749 2697 23783
rect 2731 23780 2743 23783
rect 4709 23783 4767 23789
rect 4709 23780 4721 23783
rect 2731 23752 4721 23780
rect 2731 23749 2743 23752
rect 2685 23743 2743 23749
rect 4709 23749 4721 23752
rect 4755 23749 4767 23783
rect 4709 23743 4767 23749
rect 5350 23740 5356 23792
rect 5408 23780 5414 23792
rect 6546 23780 6552 23792
rect 5408 23752 6552 23780
rect 5408 23740 5414 23752
rect 6546 23740 6552 23752
rect 6604 23740 6610 23792
rect 6638 23740 6644 23792
rect 6696 23740 6702 23792
rect 3237 23715 3295 23721
rect 3237 23712 3249 23715
rect 2627 23684 3249 23712
rect 2041 23647 2099 23653
rect 2041 23613 2053 23647
rect 2087 23613 2099 23647
rect 2041 23607 2099 23613
rect 2222 23604 2228 23656
rect 2280 23604 2286 23656
rect 2501 23647 2559 23653
rect 2501 23613 2513 23647
rect 2547 23644 2559 23647
rect 2627 23644 2655 23684
rect 3237 23681 3249 23684
rect 3283 23681 3295 23715
rect 6457 23715 6515 23721
rect 6457 23712 6469 23715
rect 3237 23675 3295 23681
rect 3344 23684 4384 23712
rect 2547 23616 2655 23644
rect 2777 23647 2835 23653
rect 2547 23613 2559 23616
rect 2501 23607 2559 23613
rect 2777 23613 2789 23647
rect 2823 23644 2835 23647
rect 3050 23644 3056 23656
rect 2823 23616 3056 23644
rect 2823 23613 2835 23616
rect 2777 23607 2835 23613
rect 3050 23604 3056 23616
rect 3108 23644 3114 23656
rect 3344 23644 3372 23684
rect 3108 23616 3372 23644
rect 3421 23647 3479 23653
rect 3108 23604 3114 23616
rect 3421 23613 3433 23647
rect 3467 23613 3479 23647
rect 3421 23607 3479 23613
rect 1213 23579 1271 23585
rect 1213 23545 1225 23579
rect 1259 23576 1271 23579
rect 1394 23576 1400 23588
rect 1259 23548 1400 23576
rect 1259 23545 1271 23548
rect 1213 23539 1271 23545
rect 1394 23536 1400 23548
rect 1452 23536 1458 23588
rect 2314 23536 2320 23588
rect 2372 23576 2378 23588
rect 3436 23576 3464 23607
rect 3602 23604 3608 23656
rect 3660 23604 3666 23656
rect 3697 23647 3755 23653
rect 3697 23613 3709 23647
rect 3743 23613 3755 23647
rect 3697 23607 3755 23613
rect 2372 23548 3464 23576
rect 3712 23576 3740 23607
rect 4062 23604 4068 23656
rect 4120 23604 4126 23656
rect 4356 23653 4384 23684
rect 4632 23684 6469 23712
rect 4632 23653 4660 23684
rect 6457 23681 6469 23684
rect 6503 23681 6515 23715
rect 6656 23712 6684 23740
rect 6840 23721 6868 23820
rect 7466 23808 7472 23860
rect 7524 23848 7530 23860
rect 7561 23851 7619 23857
rect 7561 23848 7573 23851
rect 7524 23820 7573 23848
rect 7524 23808 7530 23820
rect 7561 23817 7573 23820
rect 7607 23817 7619 23851
rect 7561 23811 7619 23817
rect 7834 23808 7840 23860
rect 7892 23848 7898 23860
rect 7892 23820 8156 23848
rect 7892 23808 7898 23820
rect 7208 23752 8064 23780
rect 6457 23675 6515 23681
rect 6564 23684 6684 23712
rect 6825 23715 6883 23721
rect 6564 23656 6592 23684
rect 6825 23681 6837 23715
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 6917 23715 6975 23721
rect 6917 23681 6929 23715
rect 6963 23712 6975 23715
rect 7098 23712 7104 23724
rect 6963 23684 7104 23712
rect 6963 23681 6975 23684
rect 6917 23675 6975 23681
rect 7098 23672 7104 23684
rect 7156 23672 7162 23724
rect 4341 23647 4399 23653
rect 4341 23613 4353 23647
rect 4387 23613 4399 23647
rect 4341 23607 4399 23613
rect 4617 23647 4675 23653
rect 4617 23613 4629 23647
rect 4663 23613 4675 23647
rect 4617 23607 4675 23613
rect 4893 23647 4951 23653
rect 4893 23613 4905 23647
rect 4939 23644 4951 23647
rect 5074 23644 5080 23656
rect 4939 23616 5080 23644
rect 4939 23613 4951 23616
rect 4893 23607 4951 23613
rect 4430 23576 4436 23588
rect 3712 23548 4436 23576
rect 2372 23536 2378 23548
rect 2792 23520 2820 23548
rect 4430 23536 4436 23548
rect 4488 23576 4494 23588
rect 4525 23579 4583 23585
rect 4525 23576 4537 23579
rect 4488 23548 4537 23576
rect 4488 23536 4494 23548
rect 4525 23545 4537 23548
rect 4571 23576 4583 23579
rect 4908 23576 4936 23607
rect 5074 23604 5080 23616
rect 5132 23604 5138 23656
rect 5169 23647 5227 23653
rect 5169 23613 5181 23647
rect 5215 23613 5227 23647
rect 5169 23607 5227 23613
rect 4571 23548 4936 23576
rect 4571 23545 4583 23548
rect 4525 23539 4583 23545
rect 2774 23468 2780 23520
rect 2832 23468 2838 23520
rect 3786 23468 3792 23520
rect 3844 23508 3850 23520
rect 3973 23511 4031 23517
rect 3973 23508 3985 23511
rect 3844 23480 3985 23508
rect 3844 23468 3850 23480
rect 3973 23477 3985 23480
rect 4019 23477 4031 23511
rect 3973 23471 4031 23477
rect 4798 23468 4804 23520
rect 4856 23508 4862 23520
rect 5184 23508 5212 23607
rect 5258 23604 5264 23656
rect 5316 23604 5322 23656
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6161 23647 6219 23653
rect 6161 23644 6173 23647
rect 5921 23616 6173 23644
rect 5353 23579 5411 23585
rect 5353 23545 5365 23579
rect 5399 23576 5411 23579
rect 5718 23576 5724 23588
rect 5399 23548 5724 23576
rect 5399 23545 5411 23548
rect 5353 23539 5411 23545
rect 5718 23536 5724 23548
rect 5776 23536 5782 23588
rect 5921 23520 5949 23616
rect 6161 23613 6173 23616
rect 6207 23613 6219 23647
rect 6161 23607 6219 23613
rect 6365 23647 6423 23653
rect 6365 23613 6377 23647
rect 6411 23613 6423 23647
rect 6365 23607 6423 23613
rect 6079 23579 6137 23585
rect 6079 23545 6091 23579
rect 6125 23545 6137 23579
rect 6079 23539 6137 23545
rect 4856 23480 5212 23508
rect 4856 23468 4862 23480
rect 5442 23468 5448 23520
rect 5500 23508 5506 23520
rect 5626 23508 5632 23520
rect 5500 23480 5632 23508
rect 5500 23468 5506 23480
rect 5626 23468 5632 23480
rect 5684 23468 5690 23520
rect 5902 23468 5908 23520
rect 5960 23468 5966 23520
rect 6104 23508 6132 23539
rect 6270 23536 6276 23588
rect 6328 23536 6334 23588
rect 6380 23576 6408 23607
rect 6546 23604 6552 23656
rect 6604 23604 6610 23656
rect 6638 23604 6644 23656
rect 6696 23604 6702 23656
rect 6733 23647 6791 23653
rect 6733 23613 6745 23647
rect 6779 23644 6791 23647
rect 7208 23644 7236 23752
rect 7742 23672 7748 23724
rect 7800 23672 7806 23724
rect 6779 23616 7236 23644
rect 6779 23613 6791 23616
rect 6733 23607 6791 23613
rect 7282 23604 7288 23656
rect 7340 23604 7346 23656
rect 7377 23647 7435 23653
rect 7377 23613 7389 23647
rect 7423 23613 7435 23647
rect 7377 23607 7435 23613
rect 7635 23647 7693 23653
rect 7635 23613 7647 23647
rect 7681 23644 7693 23647
rect 7681 23616 7880 23644
rect 7681 23613 7693 23616
rect 7635 23607 7693 23613
rect 6914 23576 6920 23588
rect 6380 23548 6920 23576
rect 6914 23536 6920 23548
rect 6972 23576 6978 23588
rect 7101 23579 7159 23585
rect 7101 23576 7113 23579
rect 6972 23548 7113 23576
rect 6972 23536 6978 23548
rect 7101 23545 7113 23548
rect 7147 23545 7159 23579
rect 7101 23539 7159 23545
rect 7190 23536 7196 23588
rect 7248 23576 7254 23588
rect 7392 23576 7420 23607
rect 7852 23588 7880 23616
rect 7248 23548 7420 23576
rect 7248 23536 7254 23548
rect 7834 23536 7840 23588
rect 7892 23536 7898 23588
rect 7929 23579 7987 23585
rect 7929 23545 7941 23579
rect 7975 23545 7987 23579
rect 8036 23576 8064 23752
rect 8128 23712 8156 23820
rect 8202 23808 8208 23860
rect 8260 23808 8266 23860
rect 8386 23808 8392 23860
rect 8444 23808 8450 23860
rect 8496 23820 9352 23848
rect 8220 23780 8248 23808
rect 8496 23780 8524 23820
rect 8220 23752 8524 23780
rect 8662 23740 8668 23792
rect 8720 23740 8726 23792
rect 8754 23740 8760 23792
rect 8812 23780 8818 23792
rect 8938 23780 8944 23792
rect 8812 23752 8944 23780
rect 8812 23740 8818 23752
rect 8938 23740 8944 23752
rect 8996 23740 9002 23792
rect 9030 23740 9036 23792
rect 9088 23740 9094 23792
rect 9214 23740 9220 23792
rect 9272 23740 9278 23792
rect 9324 23780 9352 23820
rect 10134 23808 10140 23860
rect 10192 23848 10198 23860
rect 10321 23851 10379 23857
rect 10321 23848 10333 23851
rect 10192 23820 10333 23848
rect 10192 23808 10198 23820
rect 10321 23817 10333 23820
rect 10367 23848 10379 23851
rect 10410 23848 10416 23860
rect 10367 23820 10416 23848
rect 10367 23817 10379 23820
rect 10321 23811 10379 23817
rect 10410 23808 10416 23820
rect 10468 23808 10474 23860
rect 10597 23851 10655 23857
rect 10597 23817 10609 23851
rect 10643 23848 10655 23851
rect 11330 23848 11336 23860
rect 10643 23820 11336 23848
rect 10643 23817 10655 23820
rect 10597 23811 10655 23817
rect 11330 23808 11336 23820
rect 11388 23808 11394 23860
rect 9324 23752 10272 23780
rect 8680 23712 8708 23740
rect 9048 23712 9076 23740
rect 9232 23712 9260 23740
rect 8128 23684 8524 23712
rect 8110 23576 8116 23588
rect 8036 23548 8116 23576
rect 7929 23539 7987 23545
rect 6546 23508 6552 23520
rect 6104 23480 6552 23508
rect 6546 23468 6552 23480
rect 6604 23508 6610 23520
rect 7944 23508 7972 23539
rect 8110 23536 8116 23548
rect 8168 23536 8174 23588
rect 8496 23576 8524 23684
rect 8588 23684 8708 23712
rect 8864 23684 9076 23712
rect 9140 23684 9260 23712
rect 9401 23715 9459 23721
rect 8588 23653 8616 23684
rect 8573 23647 8631 23653
rect 8573 23613 8585 23647
rect 8619 23613 8631 23647
rect 8573 23607 8631 23613
rect 8665 23647 8723 23653
rect 8665 23613 8677 23647
rect 8711 23644 8723 23647
rect 8864 23644 8892 23684
rect 8711 23616 8892 23644
rect 8711 23613 8723 23616
rect 8665 23607 8723 23613
rect 8938 23604 8944 23656
rect 8996 23604 9002 23656
rect 9030 23604 9036 23656
rect 9088 23604 9094 23656
rect 9140 23653 9168 23684
rect 9401 23681 9413 23715
rect 9447 23712 9459 23715
rect 10134 23712 10140 23724
rect 9447 23684 9720 23712
rect 9447 23681 9459 23684
rect 9401 23675 9459 23681
rect 9125 23647 9183 23653
rect 9125 23613 9137 23647
rect 9171 23613 9183 23647
rect 9125 23607 9183 23613
rect 9214 23604 9220 23656
rect 9272 23604 9278 23656
rect 9493 23647 9551 23653
rect 9493 23613 9505 23647
rect 9539 23644 9551 23647
rect 9582 23644 9588 23656
rect 9539 23616 9588 23644
rect 9539 23613 9551 23616
rect 9493 23607 9551 23613
rect 9582 23604 9588 23616
rect 9640 23604 9646 23656
rect 8757 23579 8815 23585
rect 8757 23576 8769 23579
rect 8496 23548 8769 23576
rect 8757 23545 8769 23548
rect 8803 23545 8815 23579
rect 8956 23576 8984 23604
rect 8956 23548 9076 23576
rect 8757 23539 8815 23545
rect 6604 23480 7972 23508
rect 6604 23468 6610 23480
rect 8570 23468 8576 23520
rect 8628 23508 8634 23520
rect 8938 23508 8944 23520
rect 8628 23480 8944 23508
rect 8628 23468 8634 23480
rect 8938 23468 8944 23480
rect 8996 23468 9002 23520
rect 9048 23508 9076 23548
rect 9398 23536 9404 23588
rect 9456 23536 9462 23588
rect 9582 23508 9588 23520
rect 9048 23480 9588 23508
rect 9582 23468 9588 23480
rect 9640 23468 9646 23520
rect 9692 23517 9720 23684
rect 9876 23684 10140 23712
rect 9766 23604 9772 23656
rect 9824 23604 9830 23656
rect 9876 23653 9904 23684
rect 10134 23672 10140 23684
rect 10192 23672 10198 23724
rect 9861 23647 9919 23653
rect 9861 23613 9873 23647
rect 9907 23613 9919 23647
rect 9861 23607 9919 23613
rect 10042 23604 10048 23656
rect 10100 23604 10106 23656
rect 10244 23653 10272 23752
rect 11054 23672 11060 23724
rect 11112 23672 11118 23724
rect 10229 23647 10287 23653
rect 10229 23613 10241 23647
rect 10275 23613 10287 23647
rect 10229 23607 10287 23613
rect 10318 23604 10324 23656
rect 10376 23644 10382 23656
rect 10413 23647 10471 23653
rect 10413 23644 10425 23647
rect 10376 23616 10425 23644
rect 10376 23604 10382 23616
rect 10413 23613 10425 23616
rect 10459 23613 10471 23647
rect 10413 23607 10471 23613
rect 10505 23647 10563 23653
rect 10505 23613 10517 23647
rect 10551 23613 10563 23647
rect 10505 23607 10563 23613
rect 10689 23647 10747 23653
rect 10689 23613 10701 23647
rect 10735 23644 10747 23647
rect 11072 23644 11100 23672
rect 10735 23616 11100 23644
rect 10735 23613 10747 23616
rect 10689 23607 10747 23613
rect 9784 23576 9812 23604
rect 10520 23576 10548 23607
rect 9784 23548 10548 23576
rect 9677 23511 9735 23517
rect 9677 23477 9689 23511
rect 9723 23508 9735 23511
rect 9766 23508 9772 23520
rect 9723 23480 9772 23508
rect 9723 23477 9735 23480
rect 9677 23471 9735 23477
rect 9766 23468 9772 23480
rect 9824 23468 9830 23520
rect 9858 23468 9864 23520
rect 9916 23468 9922 23520
rect 10686 23468 10692 23520
rect 10744 23508 10750 23520
rect 11330 23508 11336 23520
rect 10744 23480 11336 23508
rect 10744 23468 10750 23480
rect 11330 23468 11336 23480
rect 11388 23468 11394 23520
rect 552 23418 11132 23440
rect 552 23366 4322 23418
rect 4374 23366 4386 23418
rect 4438 23366 4450 23418
rect 4502 23366 4514 23418
rect 4566 23366 4578 23418
rect 4630 23366 10722 23418
rect 10774 23366 10786 23418
rect 10838 23366 10850 23418
rect 10902 23366 10914 23418
rect 10966 23366 10978 23418
rect 11030 23366 11132 23418
rect 552 23344 11132 23366
rect 382 23264 388 23316
rect 440 23304 446 23316
rect 842 23304 848 23316
rect 440 23276 848 23304
rect 440 23264 446 23276
rect 842 23264 848 23276
rect 900 23264 906 23316
rect 1302 23264 1308 23316
rect 1360 23264 1366 23316
rect 1394 23264 1400 23316
rect 1452 23304 1458 23316
rect 1578 23304 1584 23316
rect 1452 23276 1584 23304
rect 1452 23264 1458 23276
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 2590 23264 2596 23316
rect 2648 23304 2654 23316
rect 5077 23307 5135 23313
rect 5077 23304 5089 23307
rect 2648 23276 5089 23304
rect 2648 23264 2654 23276
rect 5077 23273 5089 23276
rect 5123 23273 5135 23307
rect 5077 23267 5135 23273
rect 6270 23264 6276 23316
rect 6328 23264 6334 23316
rect 7006 23304 7012 23316
rect 6748 23276 7012 23304
rect 2777 23239 2835 23245
rect 2777 23236 2789 23239
rect 1504 23208 2789 23236
rect 474 23128 480 23180
rect 532 23168 538 23180
rect 1121 23171 1179 23177
rect 1121 23168 1133 23171
rect 532 23140 1133 23168
rect 532 23128 538 23140
rect 1121 23137 1133 23140
rect 1167 23168 1179 23171
rect 1210 23168 1216 23180
rect 1167 23140 1216 23168
rect 1167 23137 1179 23140
rect 1121 23131 1179 23137
rect 1210 23128 1216 23140
rect 1268 23128 1274 23180
rect 1504 23177 1532 23208
rect 2777 23205 2789 23208
rect 2823 23205 2835 23239
rect 2777 23199 2835 23205
rect 3326 23196 3332 23248
rect 3384 23236 3390 23248
rect 3384 23208 3924 23236
rect 3384 23196 3390 23208
rect 1489 23171 1547 23177
rect 1489 23137 1501 23171
rect 1535 23137 1547 23171
rect 1489 23131 1547 23137
rect 1949 23171 2007 23177
rect 1949 23137 1961 23171
rect 1995 23168 2007 23171
rect 2038 23168 2044 23180
rect 1995 23140 2044 23168
rect 1995 23137 2007 23140
rect 1949 23131 2007 23137
rect 2038 23128 2044 23140
rect 2096 23128 2102 23180
rect 2130 23128 2136 23180
rect 2188 23128 2194 23180
rect 2222 23128 2228 23180
rect 2280 23128 2286 23180
rect 2314 23128 2320 23180
rect 2372 23128 2378 23180
rect 2406 23128 2412 23180
rect 2464 23128 2470 23180
rect 2593 23171 2651 23177
rect 2593 23137 2605 23171
rect 2639 23137 2651 23171
rect 2593 23131 2651 23137
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23100 1731 23103
rect 1719 23072 1808 23100
rect 1719 23069 1731 23072
rect 1673 23063 1731 23069
rect 1780 22976 1808 23072
rect 1854 23060 1860 23112
rect 1912 23100 1918 23112
rect 2608 23100 2636 23131
rect 3418 23128 3424 23180
rect 3476 23128 3482 23180
rect 3786 23128 3792 23180
rect 3844 23128 3850 23180
rect 3896 23177 3924 23208
rect 4062 23196 4068 23248
rect 4120 23236 4126 23248
rect 4120 23208 4292 23236
rect 4120 23196 4126 23208
rect 4264 23177 4292 23208
rect 4982 23196 4988 23248
rect 5040 23236 5046 23248
rect 6288 23236 6316 23264
rect 5040 23208 6592 23236
rect 5040 23196 5046 23208
rect 3881 23171 3939 23177
rect 3881 23137 3893 23171
rect 3927 23137 3939 23171
rect 3881 23131 3939 23137
rect 4249 23171 4307 23177
rect 4249 23137 4261 23171
rect 4295 23168 4307 23171
rect 4614 23168 4620 23180
rect 4295 23140 4620 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 4706 23128 4712 23180
rect 4764 23128 4770 23180
rect 5074 23128 5080 23180
rect 5132 23168 5138 23180
rect 5261 23171 5319 23177
rect 5261 23168 5273 23171
rect 5132 23140 5273 23168
rect 5132 23128 5138 23140
rect 5261 23137 5273 23140
rect 5307 23137 5319 23171
rect 5261 23131 5319 23137
rect 5810 23128 5816 23180
rect 5868 23128 5874 23180
rect 5902 23128 5908 23180
rect 5960 23128 5966 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 6178 23128 6184 23180
rect 6236 23128 6242 23180
rect 6564 23177 6592 23208
rect 6748 23177 6776 23276
rect 7006 23264 7012 23276
rect 7064 23264 7070 23316
rect 7742 23264 7748 23316
rect 7800 23304 7806 23316
rect 7926 23304 7932 23316
rect 7800 23276 7932 23304
rect 7800 23264 7806 23276
rect 7926 23264 7932 23276
rect 7984 23264 7990 23316
rect 9030 23264 9036 23316
rect 9088 23304 9094 23316
rect 9125 23307 9183 23313
rect 9125 23304 9137 23307
rect 9088 23276 9137 23304
rect 9088 23264 9094 23276
rect 9125 23273 9137 23276
rect 9171 23273 9183 23307
rect 9125 23267 9183 23273
rect 9214 23264 9220 23316
rect 9272 23264 9278 23316
rect 10318 23264 10324 23316
rect 10376 23264 10382 23316
rect 7466 23236 7472 23248
rect 7024 23208 7472 23236
rect 6273 23171 6331 23177
rect 6273 23137 6285 23171
rect 6319 23137 6331 23171
rect 6273 23131 6331 23137
rect 6549 23171 6607 23177
rect 6549 23137 6561 23171
rect 6595 23137 6607 23171
rect 6549 23131 6607 23137
rect 6733 23171 6791 23177
rect 6733 23137 6745 23171
rect 6779 23137 6791 23171
rect 6733 23131 6791 23137
rect 1912 23072 2636 23100
rect 3804 23100 3832 23128
rect 4522 23100 4528 23112
rect 3804 23072 4528 23100
rect 1912 23060 1918 23072
rect 2240 23044 2268 23072
rect 4522 23060 4528 23072
rect 4580 23060 4586 23112
rect 4798 23060 4804 23112
rect 4856 23060 4862 23112
rect 5534 23060 5540 23112
rect 5592 23060 5598 23112
rect 6288 23100 6316 23131
rect 6822 23128 6828 23180
rect 6880 23128 6886 23180
rect 7024 23177 7052 23208
rect 7466 23196 7472 23208
rect 7524 23196 7530 23248
rect 7561 23239 7619 23245
rect 7561 23205 7573 23239
rect 7607 23236 7619 23239
rect 7607 23208 8156 23236
rect 7607 23205 7619 23208
rect 7561 23199 7619 23205
rect 7009 23171 7067 23177
rect 7009 23137 7021 23171
rect 7055 23137 7067 23171
rect 7009 23131 7067 23137
rect 7101 23171 7159 23177
rect 7101 23137 7113 23171
rect 7147 23168 7159 23171
rect 7282 23168 7288 23180
rect 7147 23140 7288 23168
rect 7147 23137 7159 23140
rect 7101 23131 7159 23137
rect 7282 23128 7288 23140
rect 7340 23128 7346 23180
rect 7377 23171 7435 23177
rect 7377 23137 7389 23171
rect 7423 23168 7435 23171
rect 7423 23140 7880 23168
rect 7423 23137 7435 23140
rect 7377 23131 7435 23137
rect 6914 23100 6920 23112
rect 6288 23072 6920 23100
rect 6914 23060 6920 23072
rect 6972 23060 6978 23112
rect 7193 23103 7251 23109
rect 7193 23069 7205 23103
rect 7239 23100 7251 23103
rect 7558 23100 7564 23112
rect 7239 23072 7564 23100
rect 7239 23069 7251 23072
rect 7193 23063 7251 23069
rect 7558 23060 7564 23072
rect 7616 23060 7622 23112
rect 7852 23100 7880 23140
rect 7926 23128 7932 23180
rect 7984 23128 7990 23180
rect 8128 23168 8156 23208
rect 8202 23196 8208 23248
rect 8260 23196 8266 23248
rect 10686 23236 10692 23248
rect 8404 23208 10692 23236
rect 8128 23140 8248 23168
rect 8220 23112 8248 23140
rect 7852 23072 8156 23100
rect 2222 22992 2228 23044
rect 2280 22992 2286 23044
rect 6270 22992 6276 23044
rect 6328 23032 6334 23044
rect 8021 23035 8079 23041
rect 8021 23032 8033 23035
rect 6328 23004 8033 23032
rect 6328 22992 6334 23004
rect 8021 23001 8033 23004
rect 8067 23001 8079 23035
rect 8128 23032 8156 23072
rect 8202 23060 8208 23112
rect 8260 23060 8266 23112
rect 8404 23032 8432 23208
rect 10686 23196 10692 23208
rect 10744 23196 10750 23248
rect 8478 23128 8484 23180
rect 8536 23128 8542 23180
rect 8570 23128 8576 23180
rect 8628 23168 8634 23180
rect 8665 23171 8723 23177
rect 8665 23168 8677 23171
rect 8628 23140 8677 23168
rect 8628 23128 8634 23140
rect 8665 23137 8677 23140
rect 8711 23137 8723 23171
rect 8665 23131 8723 23137
rect 8754 23128 8760 23180
rect 8812 23128 8818 23180
rect 8849 23171 8907 23177
rect 8849 23137 8861 23171
rect 8895 23168 8907 23171
rect 8895 23140 8984 23168
rect 8895 23137 8907 23140
rect 8849 23131 8907 23137
rect 8128 23004 8432 23032
rect 8956 23032 8984 23140
rect 9030 23128 9036 23180
rect 9088 23171 9094 23180
rect 9088 23168 9168 23171
rect 9088 23143 9444 23168
rect 9088 23128 9094 23143
rect 9140 23140 9444 23143
rect 9416 23100 9444 23140
rect 9582 23128 9588 23180
rect 9640 23128 9646 23180
rect 10134 23128 10140 23180
rect 10192 23128 10198 23180
rect 9493 23103 9551 23109
rect 9493 23100 9505 23103
rect 9416 23072 9505 23100
rect 9493 23069 9505 23072
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 9766 23060 9772 23112
rect 9824 23100 9830 23112
rect 9861 23103 9919 23109
rect 9861 23100 9873 23103
rect 9824 23072 9873 23100
rect 9824 23060 9830 23072
rect 9861 23069 9873 23072
rect 9907 23069 9919 23103
rect 9861 23063 9919 23069
rect 9784 23032 9812 23060
rect 8956 23004 9168 23032
rect 8021 22995 8079 23001
rect 934 22924 940 22976
rect 992 22924 998 22976
rect 1762 22924 1768 22976
rect 1820 22924 1826 22976
rect 1854 22924 1860 22976
rect 1912 22964 1918 22976
rect 2866 22964 2872 22976
rect 1912 22936 2872 22964
rect 1912 22924 1918 22936
rect 2866 22924 2872 22936
rect 2924 22924 2930 22976
rect 4065 22967 4123 22973
rect 4065 22933 4077 22967
rect 4111 22964 4123 22967
rect 5074 22964 5080 22976
rect 4111 22936 5080 22964
rect 4111 22933 4123 22936
rect 4065 22927 4123 22933
rect 5074 22924 5080 22936
rect 5132 22924 5138 22976
rect 5445 22967 5503 22973
rect 5445 22933 5457 22967
rect 5491 22964 5503 22967
rect 6457 22967 6515 22973
rect 6457 22964 6469 22967
rect 5491 22936 6469 22964
rect 5491 22933 5503 22936
rect 5445 22927 5503 22933
rect 6457 22933 6469 22936
rect 6503 22933 6515 22967
rect 6457 22927 6515 22933
rect 6546 22924 6552 22976
rect 6604 22964 6610 22976
rect 6641 22967 6699 22973
rect 6641 22964 6653 22967
rect 6604 22936 6653 22964
rect 6604 22924 6610 22936
rect 6641 22933 6653 22936
rect 6687 22964 6699 22967
rect 7282 22964 7288 22976
rect 6687 22936 7288 22964
rect 6687 22933 6699 22936
rect 6641 22927 6699 22933
rect 7282 22924 7288 22936
rect 7340 22924 7346 22976
rect 7558 22924 7564 22976
rect 7616 22964 7622 22976
rect 7745 22967 7803 22973
rect 7745 22964 7757 22967
rect 7616 22936 7757 22964
rect 7616 22924 7622 22936
rect 7745 22933 7757 22936
rect 7791 22964 7803 22967
rect 8478 22964 8484 22976
rect 7791 22936 8484 22964
rect 7791 22933 7803 22936
rect 7745 22927 7803 22933
rect 8478 22924 8484 22936
rect 8536 22924 8542 22976
rect 9140 22964 9168 23004
rect 9416 23004 9812 23032
rect 9953 23035 10011 23041
rect 9416 22964 9444 23004
rect 9953 23001 9965 23035
rect 9999 23032 10011 23035
rect 10778 23032 10784 23044
rect 9999 23004 10784 23032
rect 9999 23001 10011 23004
rect 9953 22995 10011 23001
rect 10778 22992 10784 23004
rect 10836 22992 10842 23044
rect 9140 22936 9444 22964
rect 9582 22924 9588 22976
rect 9640 22964 9646 22976
rect 10502 22964 10508 22976
rect 9640 22936 10508 22964
rect 9640 22924 9646 22936
rect 10502 22924 10508 22936
rect 10560 22924 10566 22976
rect 552 22874 11132 22896
rect 552 22822 3662 22874
rect 3714 22822 3726 22874
rect 3778 22822 3790 22874
rect 3842 22822 3854 22874
rect 3906 22822 3918 22874
rect 3970 22822 10062 22874
rect 10114 22822 10126 22874
rect 10178 22822 10190 22874
rect 10242 22822 10254 22874
rect 10306 22822 10318 22874
rect 10370 22822 11132 22874
rect 552 22800 11132 22822
rect 842 22720 848 22772
rect 900 22760 906 22772
rect 937 22763 995 22769
rect 937 22760 949 22763
rect 900 22732 949 22760
rect 900 22720 906 22732
rect 937 22729 949 22732
rect 983 22729 995 22763
rect 937 22723 995 22729
rect 1670 22720 1676 22772
rect 1728 22760 1734 22772
rect 2041 22763 2099 22769
rect 2041 22760 2053 22763
rect 1728 22732 2053 22760
rect 1728 22720 1734 22732
rect 2041 22729 2053 22732
rect 2087 22729 2099 22763
rect 2041 22723 2099 22729
rect 2225 22763 2283 22769
rect 2225 22729 2237 22763
rect 2271 22760 2283 22763
rect 2406 22760 2412 22772
rect 2271 22732 2412 22760
rect 2271 22729 2283 22732
rect 2225 22723 2283 22729
rect 2406 22720 2412 22732
rect 2464 22720 2470 22772
rect 3605 22763 3663 22769
rect 3605 22729 3617 22763
rect 3651 22729 3663 22763
rect 3605 22723 3663 22729
rect 4341 22763 4399 22769
rect 4341 22729 4353 22763
rect 4387 22760 4399 22763
rect 4430 22760 4436 22772
rect 4387 22732 4436 22760
rect 4387 22729 4399 22732
rect 4341 22723 4399 22729
rect 198 22652 204 22704
rect 256 22692 262 22704
rect 1302 22692 1308 22704
rect 256 22664 1308 22692
rect 256 22652 262 22664
rect 1302 22652 1308 22664
rect 1360 22692 1366 22704
rect 1360 22664 1808 22692
rect 1360 22652 1366 22664
rect 750 22584 756 22636
rect 808 22624 814 22636
rect 1213 22627 1271 22633
rect 1213 22624 1225 22627
rect 808 22596 1225 22624
rect 808 22584 814 22596
rect 1213 22593 1225 22596
rect 1259 22593 1271 22627
rect 1780 22624 1808 22664
rect 2590 22652 2596 22704
rect 2648 22692 2654 22704
rect 3050 22692 3056 22704
rect 2648 22664 3056 22692
rect 2648 22652 2654 22664
rect 3050 22652 3056 22664
rect 3108 22652 3114 22704
rect 2774 22624 2780 22636
rect 1780 22596 1900 22624
rect 1213 22587 1271 22593
rect 934 22516 940 22568
rect 992 22556 998 22568
rect 1121 22559 1179 22565
rect 1121 22556 1133 22559
rect 992 22528 1133 22556
rect 992 22516 998 22528
rect 1121 22525 1133 22528
rect 1167 22525 1179 22559
rect 1121 22519 1179 22525
rect 1670 22516 1676 22568
rect 1728 22516 1734 22568
rect 1762 22516 1768 22568
rect 1820 22516 1826 22568
rect 1872 22565 1900 22596
rect 2424 22596 2780 22624
rect 2424 22565 2452 22596
rect 2774 22584 2780 22596
rect 2832 22584 2838 22636
rect 3068 22565 3096 22652
rect 1857 22559 1915 22565
rect 1857 22525 1869 22559
rect 1903 22525 1915 22559
rect 1857 22519 1915 22525
rect 2409 22559 2467 22565
rect 2409 22525 2421 22559
rect 2455 22525 2467 22559
rect 2409 22519 2467 22525
rect 2685 22559 2743 22565
rect 2685 22525 2697 22559
rect 2731 22525 2743 22559
rect 2685 22519 2743 22525
rect 3053 22559 3111 22565
rect 3053 22525 3065 22559
rect 3099 22525 3111 22559
rect 3053 22519 3111 22525
rect 3237 22559 3295 22565
rect 3237 22525 3249 22559
rect 3283 22556 3295 22559
rect 3418 22556 3424 22568
rect 3283 22528 3424 22556
rect 3283 22525 3295 22528
rect 3237 22519 3295 22525
rect 1210 22448 1216 22500
rect 1268 22488 1274 22500
rect 2424 22488 2452 22519
rect 1268 22460 2452 22488
rect 1268 22448 1274 22460
rect 2700 22432 2728 22519
rect 3418 22516 3424 22528
rect 3476 22516 3482 22568
rect 3620 22556 3648 22723
rect 4430 22720 4436 22732
rect 4488 22720 4494 22772
rect 4801 22763 4859 22769
rect 4801 22729 4813 22763
rect 4847 22760 4859 22763
rect 4847 22732 5856 22760
rect 4847 22729 4859 22732
rect 4801 22723 4859 22729
rect 5169 22695 5227 22701
rect 5169 22661 5181 22695
rect 5215 22692 5227 22695
rect 5442 22692 5448 22704
rect 5215 22664 5448 22692
rect 5215 22661 5227 22664
rect 5169 22655 5227 22661
rect 5442 22652 5448 22664
rect 5500 22652 5506 22704
rect 5828 22692 5856 22732
rect 5902 22720 5908 22772
rect 5960 22720 5966 22772
rect 6178 22720 6184 22772
rect 6236 22760 6242 22772
rect 6365 22763 6423 22769
rect 6365 22760 6377 22763
rect 6236 22732 6377 22760
rect 6236 22720 6242 22732
rect 6365 22729 6377 22732
rect 6411 22729 6423 22763
rect 6365 22723 6423 22729
rect 6638 22720 6644 22772
rect 6696 22760 6702 22772
rect 6825 22763 6883 22769
rect 6825 22760 6837 22763
rect 6696 22732 6837 22760
rect 6696 22720 6702 22732
rect 6825 22729 6837 22732
rect 6871 22729 6883 22763
rect 6825 22723 6883 22729
rect 7098 22720 7104 22772
rect 7156 22760 7162 22772
rect 7653 22763 7711 22769
rect 7653 22760 7665 22763
rect 7156 22732 7665 22760
rect 7156 22720 7162 22732
rect 7653 22729 7665 22732
rect 7699 22729 7711 22763
rect 7653 22723 7711 22729
rect 8754 22720 8760 22772
rect 8812 22760 8818 22772
rect 9585 22763 9643 22769
rect 9585 22760 9597 22763
rect 8812 22732 9597 22760
rect 8812 22720 8818 22732
rect 9585 22729 9597 22732
rect 9631 22760 9643 22763
rect 10778 22760 10784 22772
rect 9631 22732 10784 22760
rect 9631 22729 9643 22732
rect 9585 22723 9643 22729
rect 10778 22720 10784 22732
rect 10836 22720 10842 22772
rect 7374 22692 7380 22704
rect 5828 22664 7380 22692
rect 7374 22652 7380 22664
rect 7432 22692 7438 22704
rect 7926 22692 7932 22704
rect 7432 22664 7932 22692
rect 7432 22652 7438 22664
rect 7926 22652 7932 22664
rect 7984 22652 7990 22704
rect 8665 22695 8723 22701
rect 8665 22661 8677 22695
rect 8711 22692 8723 22695
rect 9674 22692 9680 22704
rect 8711 22664 9680 22692
rect 8711 22661 8723 22664
rect 8665 22655 8723 22661
rect 9674 22652 9680 22664
rect 9732 22652 9738 22704
rect 10229 22695 10287 22701
rect 10229 22692 10241 22695
rect 10060 22664 10241 22692
rect 3694 22584 3700 22636
rect 3752 22624 3758 22636
rect 3752 22596 4289 22624
rect 3752 22584 3758 22596
rect 4154 22556 4160 22568
rect 3620 22528 4160 22556
rect 4154 22516 4160 22528
rect 4212 22516 4218 22568
rect 4261 22556 4289 22596
rect 4522 22584 4528 22636
rect 4580 22624 4586 22636
rect 4580 22596 5396 22624
rect 4580 22584 4586 22596
rect 5184 22565 5212 22596
rect 5368 22565 5396 22596
rect 5718 22584 5724 22636
rect 5776 22624 5782 22636
rect 5902 22624 5908 22636
rect 5776 22596 5908 22624
rect 5776 22584 5782 22596
rect 5902 22584 5908 22596
rect 5960 22584 5966 22636
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22624 7527 22627
rect 8021 22627 8079 22633
rect 8021 22624 8033 22627
rect 7515 22596 8033 22624
rect 7515 22593 7527 22596
rect 7469 22587 7527 22593
rect 8021 22593 8033 22596
rect 8067 22624 8079 22627
rect 8202 22624 8208 22636
rect 8067 22596 8208 22624
rect 8067 22593 8079 22596
rect 8021 22587 8079 22593
rect 8202 22584 8208 22596
rect 8260 22584 8266 22636
rect 8478 22584 8484 22636
rect 8536 22624 8542 22636
rect 9214 22624 9220 22636
rect 8536 22596 8984 22624
rect 8536 22584 8542 22596
rect 4985 22559 5043 22565
rect 4985 22556 4997 22559
rect 4261 22528 4997 22556
rect 4985 22525 4997 22528
rect 5031 22525 5043 22559
rect 4985 22519 5043 22525
rect 5169 22559 5227 22565
rect 5169 22525 5181 22559
rect 5215 22525 5227 22559
rect 5169 22519 5227 22525
rect 5353 22559 5411 22565
rect 5353 22525 5365 22559
rect 5399 22525 5411 22559
rect 5353 22519 5411 22525
rect 6089 22559 6147 22565
rect 6089 22525 6101 22559
rect 6135 22556 6147 22559
rect 6178 22556 6184 22568
rect 6135 22528 6184 22556
rect 6135 22525 6147 22528
rect 6089 22519 6147 22525
rect 6178 22516 6184 22528
rect 6236 22516 6242 22568
rect 6546 22516 6552 22568
rect 6604 22516 6610 22568
rect 7190 22556 7196 22568
rect 6656 22528 7196 22556
rect 3510 22448 3516 22500
rect 3568 22488 3574 22500
rect 3973 22491 4031 22497
rect 3973 22488 3985 22491
rect 3568 22460 3985 22488
rect 3568 22448 3574 22460
rect 3973 22457 3985 22460
rect 4019 22488 4031 22491
rect 4246 22488 4252 22500
rect 4019 22460 4252 22488
rect 4019 22457 4031 22460
rect 3973 22451 4031 22457
rect 4246 22448 4252 22460
rect 4304 22488 4310 22500
rect 4433 22491 4491 22497
rect 4433 22488 4445 22491
rect 4304 22460 4445 22488
rect 4304 22448 4310 22460
rect 4433 22457 4445 22460
rect 4479 22457 4491 22491
rect 4433 22451 4491 22457
rect 4614 22448 4620 22500
rect 4672 22448 4678 22500
rect 5442 22448 5448 22500
rect 5500 22488 5506 22500
rect 6273 22491 6331 22497
rect 5500 22460 5672 22488
rect 5500 22448 5506 22460
rect 2498 22380 2504 22432
rect 2556 22420 2562 22432
rect 2593 22423 2651 22429
rect 2593 22420 2605 22423
rect 2556 22392 2605 22420
rect 2556 22380 2562 22392
rect 2593 22389 2605 22392
rect 2639 22389 2651 22423
rect 2593 22383 2651 22389
rect 2682 22380 2688 22432
rect 2740 22380 2746 22432
rect 2866 22380 2872 22432
rect 2924 22380 2930 22432
rect 3326 22380 3332 22432
rect 3384 22420 3390 22432
rect 3605 22423 3663 22429
rect 3605 22420 3617 22423
rect 3384 22392 3617 22420
rect 3384 22380 3390 22392
rect 3605 22389 3617 22392
rect 3651 22389 3663 22423
rect 3605 22383 3663 22389
rect 3789 22423 3847 22429
rect 3789 22389 3801 22423
rect 3835 22420 3847 22423
rect 4062 22420 4068 22432
rect 3835 22392 4068 22420
rect 3835 22389 3847 22392
rect 3789 22383 3847 22389
rect 4062 22380 4068 22392
rect 4120 22420 4126 22432
rect 4338 22420 4344 22432
rect 4120 22392 4344 22420
rect 4120 22380 4126 22392
rect 4338 22380 4344 22392
rect 4396 22380 4402 22432
rect 4706 22380 4712 22432
rect 4764 22420 4770 22432
rect 4982 22420 4988 22432
rect 4764 22392 4988 22420
rect 4764 22380 4770 22392
rect 4982 22380 4988 22392
rect 5040 22380 5046 22432
rect 5258 22380 5264 22432
rect 5316 22420 5322 22432
rect 5537 22423 5595 22429
rect 5537 22420 5549 22423
rect 5316 22392 5549 22420
rect 5316 22380 5322 22392
rect 5537 22389 5549 22392
rect 5583 22389 5595 22423
rect 5644 22420 5672 22460
rect 6273 22457 6285 22491
rect 6319 22488 6331 22491
rect 6656 22488 6684 22528
rect 7190 22516 7196 22528
rect 7248 22556 7254 22568
rect 7248 22528 7788 22556
rect 7248 22516 7254 22528
rect 6319 22460 6684 22488
rect 6319 22457 6331 22460
rect 6273 22451 6331 22457
rect 6730 22448 6736 22500
rect 6788 22448 6794 22500
rect 7285 22491 7343 22497
rect 7285 22457 7297 22491
rect 7331 22488 7343 22491
rect 7650 22488 7656 22500
rect 7331 22460 7656 22488
rect 7331 22457 7343 22460
rect 7285 22451 7343 22457
rect 7650 22448 7656 22460
rect 7708 22448 7714 22500
rect 7760 22488 7788 22528
rect 7834 22516 7840 22568
rect 7892 22516 7898 22568
rect 7926 22516 7932 22568
rect 7984 22556 7990 22568
rect 8113 22559 8171 22565
rect 8113 22556 8125 22559
rect 7984 22528 8125 22556
rect 7984 22516 7990 22528
rect 8113 22525 8125 22528
rect 8159 22525 8171 22559
rect 8113 22519 8171 22525
rect 8389 22559 8447 22565
rect 8389 22525 8401 22559
rect 8435 22525 8447 22559
rect 8389 22519 8447 22525
rect 8404 22488 8432 22519
rect 8570 22516 8576 22568
rect 8628 22516 8634 22568
rect 8956 22565 8984 22596
rect 9048 22596 9220 22624
rect 9048 22565 9076 22596
rect 9214 22584 9220 22596
rect 9272 22584 9278 22636
rect 10060 22633 10088 22664
rect 10229 22661 10241 22664
rect 10275 22661 10287 22695
rect 10229 22655 10287 22661
rect 10045 22627 10103 22633
rect 10045 22593 10057 22627
rect 10091 22593 10103 22627
rect 10045 22587 10103 22593
rect 10502 22584 10508 22636
rect 10560 22584 10566 22636
rect 8941 22559 8999 22565
rect 8941 22525 8953 22559
rect 8987 22525 8999 22559
rect 8941 22519 8999 22525
rect 9033 22559 9091 22565
rect 9033 22525 9045 22559
rect 9079 22525 9091 22559
rect 9033 22519 9091 22525
rect 9122 22516 9128 22568
rect 9180 22516 9186 22568
rect 9309 22559 9367 22565
rect 9309 22556 9321 22559
rect 9232 22528 9321 22556
rect 7760 22460 8432 22488
rect 6546 22420 6552 22432
rect 5644 22392 6552 22420
rect 5537 22383 5595 22389
rect 6546 22380 6552 22392
rect 6604 22380 6610 22432
rect 6638 22380 6644 22432
rect 6696 22420 6702 22432
rect 7098 22420 7104 22432
rect 6696 22392 7104 22420
rect 6696 22380 6702 22392
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 7190 22380 7196 22432
rect 7248 22420 7254 22432
rect 7466 22420 7472 22432
rect 7248 22392 7472 22420
rect 7248 22380 7254 22392
rect 7466 22380 7472 22392
rect 7524 22380 7530 22432
rect 8478 22380 8484 22432
rect 8536 22380 8542 22432
rect 8938 22380 8944 22432
rect 8996 22420 9002 22432
rect 9232 22420 9260 22528
rect 9309 22525 9321 22528
rect 9355 22525 9367 22559
rect 9309 22519 9367 22525
rect 9953 22559 10011 22565
rect 9953 22525 9965 22559
rect 9999 22556 10011 22559
rect 10410 22556 10416 22568
rect 9999 22528 10416 22556
rect 9999 22525 10011 22528
rect 9953 22519 10011 22525
rect 10410 22516 10416 22528
rect 10468 22516 10474 22568
rect 10597 22559 10655 22565
rect 10597 22525 10609 22559
rect 10643 22556 10655 22559
rect 11330 22556 11336 22568
rect 10643 22528 11336 22556
rect 10643 22525 10655 22528
rect 10597 22519 10655 22525
rect 11330 22516 11336 22528
rect 11388 22516 11394 22568
rect 8996 22392 9260 22420
rect 8996 22380 9002 22392
rect 552 22330 11132 22352
rect 552 22278 4322 22330
rect 4374 22278 4386 22330
rect 4438 22278 4450 22330
rect 4502 22278 4514 22330
rect 4566 22278 4578 22330
rect 4630 22278 10722 22330
rect 10774 22278 10786 22330
rect 10838 22278 10850 22330
rect 10902 22278 10914 22330
rect 10966 22278 10978 22330
rect 11030 22278 11132 22330
rect 552 22256 11132 22278
rect 1854 22176 1860 22228
rect 1912 22176 1918 22228
rect 2314 22176 2320 22228
rect 2372 22176 2378 22228
rect 2869 22219 2927 22225
rect 2869 22216 2881 22219
rect 2608 22188 2881 22216
rect 1872 22148 1900 22176
rect 2608 22148 2636 22188
rect 2869 22185 2881 22188
rect 2915 22185 2927 22219
rect 2869 22179 2927 22185
rect 2958 22176 2964 22228
rect 3016 22216 3022 22228
rect 3326 22216 3332 22228
rect 3016 22188 3332 22216
rect 3016 22176 3022 22188
rect 3326 22176 3332 22188
rect 3384 22176 3390 22228
rect 3694 22176 3700 22228
rect 3752 22176 3758 22228
rect 4430 22176 4436 22228
rect 4488 22176 4494 22228
rect 4706 22176 4712 22228
rect 4764 22176 4770 22228
rect 5166 22176 5172 22228
rect 5224 22176 5230 22228
rect 5629 22219 5687 22225
rect 5369 22188 5580 22216
rect 3712 22148 3740 22176
rect 1872 22120 2636 22148
rect 3344 22120 3740 22148
rect 3344 22092 3372 22120
rect 4154 22108 4160 22160
rect 4212 22148 4218 22160
rect 4724 22148 4752 22176
rect 4801 22151 4859 22157
rect 4801 22148 4813 22151
rect 4212 22120 4568 22148
rect 4724 22120 4813 22148
rect 4212 22108 4218 22120
rect 1762 22040 1768 22092
rect 1820 22040 1826 22092
rect 1854 22040 1860 22092
rect 1912 22080 1918 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1912 22052 2053 22080
rect 1912 22040 1918 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 2501 22083 2559 22089
rect 2501 22049 2513 22083
rect 2547 22080 2559 22083
rect 2547 22052 2636 22080
rect 2547 22049 2559 22052
rect 2501 22043 2559 22049
rect 750 21972 756 22024
rect 808 22012 814 22024
rect 1213 22015 1271 22021
rect 1213 22012 1225 22015
rect 808 21984 1225 22012
rect 808 21972 814 21984
rect 1213 21981 1225 21984
rect 1259 21981 1271 22015
rect 1213 21975 1271 21981
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 22012 2283 22015
rect 2314 22012 2320 22024
rect 2271 21984 2320 22012
rect 2271 21981 2283 21984
rect 2225 21975 2283 21981
rect 2314 21972 2320 21984
rect 2372 21972 2378 22024
rect 2608 21876 2636 22052
rect 2682 22040 2688 22092
rect 2740 22040 2746 22092
rect 2777 22083 2835 22089
rect 2777 22049 2789 22083
rect 2823 22049 2835 22083
rect 2777 22043 2835 22049
rect 2792 21944 2820 22043
rect 2958 22040 2964 22092
rect 3016 22080 3022 22092
rect 3053 22083 3111 22089
rect 3053 22080 3065 22083
rect 3016 22052 3065 22080
rect 3016 22040 3022 22052
rect 3053 22049 3065 22052
rect 3099 22049 3111 22083
rect 3053 22043 3111 22049
rect 3145 22083 3203 22089
rect 3145 22049 3157 22083
rect 3191 22049 3203 22083
rect 3145 22043 3203 22049
rect 3160 22012 3188 22043
rect 3326 22040 3332 22092
rect 3384 22040 3390 22092
rect 3421 22083 3479 22089
rect 3421 22049 3433 22083
rect 3467 22080 3479 22083
rect 3467 22052 3648 22080
rect 3467 22049 3479 22052
rect 3421 22043 3479 22049
rect 3513 22015 3571 22021
rect 3513 22012 3525 22015
rect 3160 21984 3525 22012
rect 3513 21981 3525 21984
rect 3559 21981 3571 22015
rect 3513 21975 3571 21981
rect 3418 21944 3424 21956
rect 2792 21916 3424 21944
rect 3418 21904 3424 21916
rect 3476 21904 3482 21956
rect 3620 21944 3648 22052
rect 3694 22040 3700 22092
rect 3752 22040 3758 22092
rect 3786 22040 3792 22092
rect 3844 22040 3850 22092
rect 3878 22040 3884 22092
rect 3936 22040 3942 22092
rect 4062 22040 4068 22092
rect 4120 22040 4126 22092
rect 4246 22040 4252 22092
rect 4304 22040 4310 22092
rect 4540 22089 4568 22120
rect 4801 22117 4813 22120
rect 4847 22117 4859 22151
rect 5369 22148 5397 22188
rect 4801 22111 4859 22117
rect 5000 22120 5397 22148
rect 5000 22089 5028 22120
rect 5442 22108 5448 22160
rect 5500 22108 5506 22160
rect 5552 22148 5580 22188
rect 5629 22185 5641 22219
rect 5675 22216 5687 22219
rect 5810 22216 5816 22228
rect 5675 22188 5816 22216
rect 5675 22185 5687 22188
rect 5629 22179 5687 22185
rect 5810 22176 5816 22188
rect 5868 22176 5874 22228
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 6236 22188 6592 22216
rect 6236 22176 6242 22188
rect 6270 22148 6276 22160
rect 5552 22120 6276 22148
rect 4525 22083 4583 22089
rect 4525 22049 4537 22083
rect 4571 22049 4583 22083
rect 4985 22083 5043 22089
rect 4985 22080 4997 22083
rect 4525 22043 4583 22049
rect 4724 22052 4997 22080
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 22012 4031 22015
rect 4080 22012 4108 22040
rect 4724 22024 4752 22052
rect 4985 22049 4997 22052
rect 5031 22049 5043 22083
rect 4985 22043 5043 22049
rect 5077 22083 5135 22089
rect 5077 22049 5089 22083
rect 5123 22049 5135 22083
rect 5077 22043 5135 22049
rect 4338 22012 4344 22024
rect 4019 21984 4344 22012
rect 4019 21981 4031 21984
rect 3973 21975 4031 21981
rect 4338 21972 4344 21984
rect 4396 21972 4402 22024
rect 4706 21972 4712 22024
rect 4764 21972 4770 22024
rect 5092 21944 5120 22043
rect 5258 22040 5264 22092
rect 5316 22040 5322 22092
rect 5353 22083 5411 22089
rect 5353 22049 5365 22083
rect 5399 22080 5411 22083
rect 5460 22080 5488 22108
rect 5399 22052 5488 22080
rect 5399 22049 5411 22052
rect 5353 22043 5411 22049
rect 5442 21972 5448 22024
rect 5500 21972 5506 22024
rect 5552 22012 5580 22120
rect 6270 22108 6276 22120
rect 6328 22108 6334 22160
rect 6564 22148 6592 22188
rect 6638 22176 6644 22228
rect 6696 22216 6702 22228
rect 7926 22216 7932 22228
rect 6696 22188 7932 22216
rect 6696 22176 6702 22188
rect 7926 22176 7932 22188
rect 7984 22176 7990 22228
rect 8110 22176 8116 22228
rect 8168 22176 8174 22228
rect 8220 22188 8984 22216
rect 6914 22148 6920 22160
rect 6564 22120 6920 22148
rect 6914 22108 6920 22120
rect 6972 22108 6978 22160
rect 7006 22108 7012 22160
rect 7064 22148 7070 22160
rect 7561 22151 7619 22157
rect 7561 22148 7573 22151
rect 7064 22120 7573 22148
rect 7064 22108 7070 22120
rect 7561 22117 7573 22120
rect 7607 22117 7619 22151
rect 7561 22111 7619 22117
rect 5718 22040 5724 22092
rect 5776 22080 5782 22092
rect 6638 22080 6644 22092
rect 5776 22052 6644 22080
rect 5776 22040 5782 22052
rect 6638 22040 6644 22052
rect 6696 22040 6702 22092
rect 6730 22040 6736 22092
rect 6788 22080 6794 22092
rect 7653 22083 7711 22089
rect 7653 22080 7665 22083
rect 6788 22052 7665 22080
rect 6788 22040 6794 22052
rect 7653 22049 7665 22052
rect 7699 22049 7711 22083
rect 7653 22043 7711 22049
rect 7742 22040 7748 22092
rect 7800 22080 7806 22092
rect 8220 22080 8248 22188
rect 8386 22108 8392 22160
rect 8444 22108 8450 22160
rect 8481 22151 8539 22157
rect 8481 22117 8493 22151
rect 8527 22148 8539 22151
rect 8570 22148 8576 22160
rect 8527 22120 8576 22148
rect 8527 22117 8539 22120
rect 8481 22111 8539 22117
rect 8570 22108 8576 22120
rect 8628 22108 8634 22160
rect 8757 22105 8815 22111
rect 8846 22108 8852 22160
rect 8904 22108 8910 22160
rect 7800 22052 8248 22080
rect 8297 22083 8355 22089
rect 7800 22040 7806 22052
rect 8297 22049 8309 22083
rect 8343 22049 8355 22083
rect 8665 22083 8723 22089
rect 8665 22080 8677 22083
rect 8297 22043 8355 22049
rect 8588 22052 8677 22080
rect 5629 22015 5687 22021
rect 5629 22012 5641 22015
rect 5552 21984 5641 22012
rect 5629 21981 5641 21984
rect 5675 21981 5687 22015
rect 5902 22012 5908 22024
rect 5629 21975 5687 21981
rect 5736 21984 5908 22012
rect 5736 21944 5764 21984
rect 5902 21972 5908 21984
rect 5960 22012 5966 22024
rect 7834 22012 7840 22024
rect 5960 21984 7840 22012
rect 5960 21972 5966 21984
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 8202 21972 8208 22024
rect 8260 22012 8266 22024
rect 8312 22012 8340 22043
rect 8588 22024 8616 22052
rect 8665 22049 8677 22052
rect 8711 22049 8723 22083
rect 8757 22071 8769 22105
rect 8803 22080 8815 22105
rect 8864 22080 8892 22108
rect 8956 22089 8984 22188
rect 10410 22176 10416 22228
rect 10468 22176 10474 22228
rect 10318 22148 10324 22160
rect 9968 22120 10324 22148
rect 8803 22071 8892 22080
rect 8757 22065 8892 22071
rect 8772 22052 8892 22065
rect 8941 22083 8999 22089
rect 8665 22043 8723 22049
rect 8941 22049 8953 22083
rect 8987 22049 8999 22083
rect 8941 22043 8999 22049
rect 9125 22083 9183 22089
rect 9125 22049 9137 22083
rect 9171 22080 9183 22083
rect 9214 22080 9220 22092
rect 9171 22052 9220 22080
rect 9171 22049 9183 22052
rect 9125 22043 9183 22049
rect 9214 22040 9220 22052
rect 9272 22040 9278 22092
rect 9674 22040 9680 22092
rect 9732 22040 9738 22092
rect 9968 22089 9996 22120
rect 10318 22108 10324 22120
rect 10376 22148 10382 22160
rect 10686 22148 10692 22160
rect 10376 22120 10692 22148
rect 10376 22108 10382 22120
rect 10686 22108 10692 22120
rect 10744 22108 10750 22160
rect 9953 22083 10011 22089
rect 9953 22049 9965 22083
rect 9999 22049 10011 22083
rect 9953 22043 10011 22049
rect 10042 22040 10048 22092
rect 10100 22080 10106 22092
rect 10137 22083 10195 22089
rect 10137 22080 10149 22083
rect 10100 22052 10149 22080
rect 10100 22040 10106 22052
rect 10137 22049 10149 22052
rect 10183 22049 10195 22083
rect 10137 22043 10195 22049
rect 10410 22040 10416 22092
rect 10468 22040 10474 22092
rect 10597 22083 10655 22089
rect 10597 22049 10609 22083
rect 10643 22049 10655 22083
rect 10597 22043 10655 22049
rect 8260 21984 8340 22012
rect 8260 21972 8266 21984
rect 3620 21916 5028 21944
rect 5092 21916 5764 21944
rect 2866 21876 2872 21888
rect 2608 21848 2872 21876
rect 2866 21836 2872 21848
rect 2924 21836 2930 21888
rect 3326 21836 3332 21888
rect 3384 21836 3390 21888
rect 4246 21836 4252 21888
rect 4304 21876 4310 21888
rect 4617 21879 4675 21885
rect 4617 21876 4629 21879
rect 4304 21848 4629 21876
rect 4304 21836 4310 21848
rect 4617 21845 4629 21848
rect 4663 21845 4675 21879
rect 5000 21876 5028 21916
rect 6270 21904 6276 21956
rect 6328 21904 6334 21956
rect 7282 21944 7288 21956
rect 6840 21916 7288 21944
rect 6840 21876 6868 21916
rect 7282 21904 7288 21916
rect 7340 21904 7346 21956
rect 8312 21944 8340 21984
rect 8570 21972 8576 22024
rect 8628 21972 8634 22024
rect 8754 21972 8760 22024
rect 8812 22012 8818 22024
rect 8849 22015 8907 22021
rect 8849 22012 8861 22015
rect 8812 21984 8861 22012
rect 8812 21972 8818 21984
rect 8849 21981 8861 21984
rect 8895 21981 8907 22015
rect 8849 21975 8907 21981
rect 9398 21972 9404 22024
rect 9456 21972 9462 22024
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 22012 10379 22015
rect 10612 22012 10640 22043
rect 10367 21984 10640 22012
rect 10367 21981 10379 21984
rect 10321 21975 10379 21981
rect 10594 21944 10600 21956
rect 8312 21916 10600 21944
rect 10594 21904 10600 21916
rect 10652 21904 10658 21956
rect 5000 21848 6868 21876
rect 4617 21839 4675 21845
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 7837 21879 7895 21885
rect 7837 21876 7849 21879
rect 6972 21848 7849 21876
rect 6972 21836 6978 21848
rect 7837 21845 7849 21848
rect 7883 21845 7895 21879
rect 7837 21839 7895 21845
rect 7926 21836 7932 21888
rect 7984 21876 7990 21888
rect 9309 21879 9367 21885
rect 9309 21876 9321 21879
rect 7984 21848 9321 21876
rect 7984 21836 7990 21848
rect 9309 21845 9321 21848
rect 9355 21845 9367 21879
rect 9309 21839 9367 21845
rect 9493 21879 9551 21885
rect 9493 21845 9505 21879
rect 9539 21876 9551 21879
rect 9582 21876 9588 21888
rect 9539 21848 9588 21876
rect 9539 21845 9551 21848
rect 9493 21839 9551 21845
rect 9582 21836 9588 21848
rect 9640 21836 9646 21888
rect 9674 21836 9680 21888
rect 9732 21876 9738 21888
rect 9861 21879 9919 21885
rect 9861 21876 9873 21879
rect 9732 21848 9873 21876
rect 9732 21836 9738 21848
rect 9861 21845 9873 21848
rect 9907 21845 9919 21879
rect 9861 21839 9919 21845
rect 552 21786 11132 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 10062 21786
rect 10114 21734 10126 21786
rect 10178 21734 10190 21786
rect 10242 21734 10254 21786
rect 10306 21734 10318 21786
rect 10370 21734 11132 21786
rect 552 21712 11132 21734
rect 1026 21632 1032 21684
rect 1084 21632 1090 21684
rect 1489 21675 1547 21681
rect 1489 21641 1501 21675
rect 1535 21672 1547 21675
rect 1670 21672 1676 21684
rect 1535 21644 1676 21672
rect 1535 21641 1547 21644
rect 1489 21635 1547 21641
rect 1670 21632 1676 21644
rect 1728 21632 1734 21684
rect 3142 21632 3148 21684
rect 3200 21672 3206 21684
rect 3329 21675 3387 21681
rect 3329 21672 3341 21675
rect 3200 21644 3341 21672
rect 3200 21632 3206 21644
rect 3329 21641 3341 21644
rect 3375 21641 3387 21675
rect 3329 21635 3387 21641
rect 3418 21632 3424 21684
rect 3476 21672 3482 21684
rect 4338 21672 4344 21684
rect 3476 21644 4344 21672
rect 3476 21632 3482 21644
rect 4338 21632 4344 21644
rect 4396 21632 4402 21684
rect 4525 21675 4583 21681
rect 4525 21641 4537 21675
rect 4571 21641 4583 21675
rect 4525 21635 4583 21641
rect 2222 21564 2228 21616
rect 2280 21604 2286 21616
rect 2590 21604 2596 21616
rect 2280 21576 2596 21604
rect 2280 21564 2286 21576
rect 2590 21564 2596 21576
rect 2648 21604 2654 21616
rect 3605 21607 3663 21613
rect 3605 21604 3617 21607
rect 2648 21576 3617 21604
rect 2648 21564 2654 21576
rect 3605 21573 3617 21576
rect 3651 21604 3663 21607
rect 3786 21604 3792 21616
rect 3651 21576 3792 21604
rect 3651 21573 3663 21576
rect 3605 21567 3663 21573
rect 3786 21564 3792 21576
rect 3844 21564 3850 21616
rect 3970 21564 3976 21616
rect 4028 21604 4034 21616
rect 4430 21604 4436 21616
rect 4028 21576 4436 21604
rect 4028 21564 4034 21576
rect 4430 21564 4436 21576
rect 4488 21564 4494 21616
rect 4540 21604 4568 21635
rect 5166 21632 5172 21684
rect 5224 21672 5230 21684
rect 6365 21675 6423 21681
rect 6365 21672 6377 21675
rect 5224 21644 6377 21672
rect 5224 21632 5230 21644
rect 6365 21641 6377 21644
rect 6411 21641 6423 21675
rect 6546 21672 6552 21684
rect 6365 21635 6423 21641
rect 6472 21644 6552 21672
rect 5721 21607 5779 21613
rect 4540 21576 5212 21604
rect 5184 21548 5212 21576
rect 5276 21576 5580 21604
rect 2038 21536 2044 21548
rect 1872 21508 2044 21536
rect 1213 21471 1271 21477
rect 1213 21437 1225 21471
rect 1259 21468 1271 21471
rect 1302 21468 1308 21480
rect 1259 21440 1308 21468
rect 1259 21437 1271 21440
rect 1213 21431 1271 21437
rect 1302 21428 1308 21440
rect 1360 21428 1366 21480
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 1578 21468 1584 21480
rect 1443 21440 1584 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 1578 21428 1584 21440
rect 1636 21428 1642 21480
rect 1872 21477 1900 21508
rect 2038 21496 2044 21508
rect 2096 21536 2102 21548
rect 2406 21536 2412 21548
rect 2096 21508 2412 21536
rect 2096 21496 2102 21508
rect 2406 21496 2412 21508
rect 2464 21496 2470 21548
rect 4982 21536 4988 21548
rect 3436 21508 4988 21536
rect 1673 21471 1731 21477
rect 1673 21437 1685 21471
rect 1719 21437 1731 21471
rect 1673 21431 1731 21437
rect 1857 21471 1915 21477
rect 1857 21437 1869 21471
rect 1903 21437 1915 21471
rect 1857 21431 1915 21437
rect 1949 21471 2007 21477
rect 1949 21437 1961 21471
rect 1995 21468 2007 21471
rect 2593 21471 2651 21477
rect 2593 21468 2605 21471
rect 1995 21440 2605 21468
rect 1995 21437 2007 21440
rect 1949 21431 2007 21437
rect 2593 21437 2605 21440
rect 2639 21437 2651 21471
rect 2593 21431 2651 21437
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 2866 21468 2872 21480
rect 2823 21440 2872 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 1688 21400 1716 21431
rect 2866 21428 2872 21440
rect 2924 21428 2930 21480
rect 3053 21471 3111 21477
rect 3053 21437 3065 21471
rect 3099 21468 3111 21471
rect 3142 21468 3148 21480
rect 3099 21440 3148 21468
rect 3099 21437 3111 21440
rect 3053 21431 3111 21437
rect 3142 21428 3148 21440
rect 3200 21428 3206 21480
rect 3237 21471 3295 21477
rect 3237 21437 3249 21471
rect 3283 21468 3295 21471
rect 3326 21468 3332 21480
rect 3283 21440 3332 21468
rect 3283 21437 3295 21440
rect 3237 21431 3295 21437
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 3436 21477 3464 21508
rect 4982 21496 4988 21508
rect 5040 21496 5046 21548
rect 5166 21496 5172 21548
rect 5224 21496 5230 21548
rect 5276 21545 5304 21576
rect 5261 21539 5319 21545
rect 5261 21505 5273 21539
rect 5307 21505 5319 21539
rect 5261 21499 5319 21505
rect 5442 21496 5448 21548
rect 5500 21496 5506 21548
rect 5552 21536 5580 21576
rect 5721 21573 5733 21607
rect 5767 21604 5779 21607
rect 5902 21604 5908 21616
rect 5767 21576 5908 21604
rect 5767 21573 5779 21576
rect 5721 21567 5779 21573
rect 5902 21564 5908 21576
rect 5960 21564 5966 21616
rect 6181 21607 6239 21613
rect 6181 21573 6193 21607
rect 6227 21604 6239 21607
rect 6472 21604 6500 21644
rect 6546 21632 6552 21644
rect 6604 21672 6610 21684
rect 7466 21672 7472 21684
rect 6604 21644 7472 21672
rect 6604 21632 6610 21644
rect 7466 21632 7472 21644
rect 7524 21672 7530 21684
rect 7524 21644 8064 21672
rect 7524 21632 7530 21644
rect 7009 21607 7067 21613
rect 7009 21604 7021 21607
rect 6227 21576 6500 21604
rect 6656 21576 7021 21604
rect 6227 21573 6239 21576
rect 6181 21567 6239 21573
rect 6549 21539 6607 21545
rect 5552 21508 6390 21536
rect 3421 21471 3479 21477
rect 3421 21437 3433 21471
rect 3467 21437 3479 21471
rect 3421 21431 3479 21437
rect 3602 21428 3608 21480
rect 3660 21468 3666 21480
rect 3970 21468 3976 21480
rect 3660 21440 3976 21468
rect 3660 21428 3666 21440
rect 3970 21428 3976 21440
rect 4028 21428 4034 21480
rect 4249 21471 4307 21477
rect 4249 21437 4261 21471
rect 4295 21468 4307 21471
rect 4338 21468 4344 21480
rect 4295 21440 4344 21468
rect 4295 21437 4307 21440
rect 4249 21431 4307 21437
rect 4338 21428 4344 21440
rect 4396 21428 4402 21480
rect 4798 21428 4804 21480
rect 4856 21468 4862 21480
rect 5626 21468 5632 21480
rect 4856 21440 5632 21468
rect 4856 21428 4862 21440
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 5718 21428 5724 21480
rect 5776 21468 5782 21480
rect 5906 21471 5964 21477
rect 5906 21470 5918 21471
rect 5828 21468 5918 21470
rect 5776 21442 5918 21468
rect 5776 21440 5856 21442
rect 5776 21428 5782 21440
rect 5906 21437 5918 21442
rect 5952 21437 5964 21471
rect 5906 21431 5964 21437
rect 5994 21428 6000 21480
rect 6052 21468 6058 21480
rect 6178 21468 6184 21480
rect 6052 21440 6184 21468
rect 6052 21428 6058 21440
rect 6178 21428 6184 21440
rect 6236 21428 6242 21480
rect 6270 21428 6276 21480
rect 6328 21428 6334 21480
rect 2409 21403 2467 21409
rect 2409 21400 2421 21403
rect 1688 21372 2421 21400
rect 2409 21369 2421 21372
rect 2455 21400 2467 21403
rect 2498 21400 2504 21412
rect 2455 21372 2504 21400
rect 2455 21369 2467 21372
rect 2409 21363 2467 21369
rect 2498 21360 2504 21372
rect 2556 21360 2562 21412
rect 2682 21360 2688 21412
rect 2740 21400 2746 21412
rect 2961 21403 3019 21409
rect 2961 21400 2973 21403
rect 2740 21372 2973 21400
rect 2740 21360 2746 21372
rect 2961 21369 2973 21372
rect 3007 21400 3019 21403
rect 3878 21400 3884 21412
rect 3007 21372 3884 21400
rect 3007 21369 3019 21372
rect 2961 21363 3019 21369
rect 3878 21360 3884 21372
rect 3936 21360 3942 21412
rect 4062 21360 4068 21412
rect 4120 21400 4126 21412
rect 4709 21403 4767 21409
rect 4709 21400 4721 21403
rect 4120 21372 4721 21400
rect 4120 21360 4126 21372
rect 4709 21369 4721 21372
rect 4755 21400 4767 21403
rect 5810 21400 5816 21412
rect 4755 21372 5816 21400
rect 4755 21369 4767 21372
rect 4709 21363 4767 21369
rect 5810 21360 5816 21372
rect 5868 21360 5874 21412
rect 6362 21400 6390 21508
rect 6549 21505 6561 21539
rect 6595 21536 6607 21539
rect 6656 21536 6684 21576
rect 7009 21573 7021 21576
rect 7055 21573 7067 21607
rect 7009 21567 7067 21573
rect 7098 21564 7104 21616
rect 7156 21604 7162 21616
rect 7282 21604 7288 21616
rect 7156 21576 7288 21604
rect 7156 21564 7162 21576
rect 7282 21564 7288 21576
rect 7340 21564 7346 21616
rect 7926 21604 7932 21616
rect 7576 21576 7932 21604
rect 6595 21508 6684 21536
rect 6595 21505 6607 21508
rect 6549 21499 6607 21505
rect 6730 21496 6736 21548
rect 6788 21496 6794 21548
rect 6825 21539 6883 21545
rect 6825 21505 6837 21539
rect 6871 21536 6883 21539
rect 7576 21536 7604 21576
rect 7926 21564 7932 21576
rect 7984 21564 7990 21616
rect 8036 21604 8064 21644
rect 8570 21632 8576 21684
rect 8628 21672 8634 21684
rect 8849 21675 8907 21681
rect 8849 21672 8861 21675
rect 8628 21644 8861 21672
rect 8628 21632 8634 21644
rect 8849 21641 8861 21644
rect 8895 21641 8907 21675
rect 8849 21635 8907 21641
rect 8938 21632 8944 21684
rect 8996 21672 9002 21684
rect 9214 21672 9220 21684
rect 8996 21644 9220 21672
rect 8996 21632 9002 21644
rect 9214 21632 9220 21644
rect 9272 21632 9278 21684
rect 9861 21675 9919 21681
rect 9861 21641 9873 21675
rect 9907 21672 9919 21675
rect 10410 21672 10416 21684
rect 9907 21644 10416 21672
rect 9907 21641 9919 21644
rect 9861 21635 9919 21641
rect 10410 21632 10416 21644
rect 10468 21632 10474 21684
rect 9585 21607 9643 21613
rect 9585 21604 9597 21607
rect 8036 21576 9597 21604
rect 9585 21573 9597 21576
rect 9631 21573 9643 21607
rect 9585 21567 9643 21573
rect 6871 21508 7604 21536
rect 7653 21539 7711 21545
rect 6871 21505 6883 21508
rect 6825 21499 6883 21505
rect 7653 21505 7665 21539
rect 7699 21536 7711 21539
rect 7742 21536 7748 21548
rect 7699 21508 7748 21536
rect 7699 21505 7711 21508
rect 7653 21499 7711 21505
rect 7742 21496 7748 21508
rect 7800 21496 7806 21548
rect 8662 21496 8668 21548
rect 8720 21536 8726 21548
rect 8938 21536 8944 21548
rect 8720 21508 8944 21536
rect 8720 21496 8726 21508
rect 8938 21496 8944 21508
rect 8996 21496 9002 21548
rect 9306 21496 9312 21548
rect 9364 21536 9370 21548
rect 9364 21508 9444 21536
rect 9364 21496 9370 21508
rect 6638 21428 6644 21480
rect 6696 21428 6702 21480
rect 7190 21468 7196 21480
rect 6748 21440 7196 21468
rect 6748 21400 6776 21440
rect 7190 21428 7196 21440
rect 7248 21468 7254 21480
rect 7377 21471 7435 21477
rect 7377 21468 7389 21471
rect 7248 21440 7389 21468
rect 7248 21428 7254 21440
rect 7377 21437 7389 21440
rect 7423 21437 7435 21471
rect 7377 21431 7435 21437
rect 7926 21428 7932 21480
rect 7984 21468 7990 21480
rect 8205 21471 8263 21477
rect 8205 21468 8217 21471
rect 7984 21440 8217 21468
rect 7984 21428 7990 21440
rect 8205 21437 8217 21440
rect 8251 21437 8263 21471
rect 8205 21431 8263 21437
rect 8386 21428 8392 21480
rect 8444 21428 8450 21480
rect 8478 21428 8484 21480
rect 8536 21468 8542 21480
rect 9416 21477 9444 21508
rect 9222 21471 9280 21477
rect 9222 21468 9234 21471
rect 8536 21440 9234 21468
rect 8536 21428 8542 21440
rect 9222 21437 9234 21440
rect 9268 21437 9280 21471
rect 9222 21431 9280 21437
rect 9401 21471 9459 21477
rect 9401 21437 9413 21471
rect 9447 21437 9459 21471
rect 9401 21431 9459 21437
rect 9582 21428 9588 21480
rect 9640 21428 9646 21480
rect 9769 21471 9827 21477
rect 9769 21437 9781 21471
rect 9815 21437 9827 21471
rect 9769 21431 9827 21437
rect 6362 21372 6776 21400
rect 7006 21360 7012 21412
rect 7064 21400 7070 21412
rect 7558 21400 7564 21412
rect 7064 21372 7564 21400
rect 7064 21360 7070 21372
rect 7558 21360 7564 21372
rect 7616 21400 7622 21412
rect 8021 21403 8079 21409
rect 8021 21400 8033 21403
rect 7616 21372 8033 21400
rect 7616 21360 7622 21372
rect 8021 21369 8033 21372
rect 8067 21369 8079 21403
rect 8021 21363 8079 21369
rect 8754 21360 8760 21412
rect 8812 21400 8818 21412
rect 8849 21403 8907 21409
rect 8849 21400 8861 21403
rect 8812 21372 8861 21400
rect 8812 21360 8818 21372
rect 8849 21369 8861 21372
rect 8895 21369 8907 21403
rect 8849 21363 8907 21369
rect 8938 21360 8944 21412
rect 8996 21400 9002 21412
rect 9033 21403 9091 21409
rect 9033 21400 9045 21403
rect 8996 21372 9045 21400
rect 8996 21360 9002 21372
rect 9033 21369 9045 21372
rect 9079 21369 9091 21403
rect 9033 21363 9091 21369
rect 9125 21403 9183 21409
rect 9125 21369 9137 21403
rect 9171 21400 9183 21403
rect 9600 21400 9628 21428
rect 9171 21372 9628 21400
rect 9784 21400 9812 21431
rect 9950 21428 9956 21480
rect 10008 21428 10014 21480
rect 10134 21400 10140 21412
rect 9784 21372 10140 21400
rect 9171 21369 9183 21372
rect 9125 21363 9183 21369
rect 10134 21360 10140 21372
rect 10192 21400 10198 21412
rect 10686 21400 10692 21412
rect 10192 21372 10692 21400
rect 10192 21360 10198 21372
rect 10686 21360 10692 21372
rect 10744 21360 10750 21412
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 2133 21335 2191 21341
rect 2133 21332 2145 21335
rect 1452 21304 2145 21332
rect 1452 21292 1458 21304
rect 2133 21301 2145 21304
rect 2179 21332 2191 21335
rect 2222 21332 2228 21344
rect 2179 21304 2228 21332
rect 2179 21301 2191 21304
rect 2133 21295 2191 21301
rect 2222 21292 2228 21304
rect 2280 21292 2286 21344
rect 2314 21292 2320 21344
rect 2372 21332 2378 21344
rect 3050 21332 3056 21344
rect 2372 21304 3056 21332
rect 2372 21292 2378 21304
rect 3050 21292 3056 21304
rect 3108 21292 3114 21344
rect 3694 21292 3700 21344
rect 3752 21332 3758 21344
rect 4341 21335 4399 21341
rect 4341 21332 4353 21335
rect 3752 21304 4353 21332
rect 3752 21292 3758 21304
rect 4341 21301 4353 21304
rect 4387 21301 4399 21335
rect 4341 21295 4399 21301
rect 4509 21335 4567 21341
rect 4509 21301 4521 21335
rect 4555 21332 4567 21335
rect 4801 21335 4859 21341
rect 4801 21332 4813 21335
rect 4555 21304 4813 21332
rect 4555 21301 4567 21304
rect 4509 21295 4567 21301
rect 4801 21301 4813 21304
rect 4847 21301 4859 21335
rect 4801 21295 4859 21301
rect 5169 21335 5227 21341
rect 5169 21301 5181 21335
rect 5215 21332 5227 21335
rect 7469 21335 7527 21341
rect 7469 21332 7481 21335
rect 5215 21304 7481 21332
rect 5215 21301 5227 21304
rect 5169 21295 5227 21301
rect 7469 21301 7481 21304
rect 7515 21332 7527 21335
rect 7650 21332 7656 21344
rect 7515 21304 7656 21332
rect 7515 21301 7527 21304
rect 7469 21295 7527 21301
rect 7650 21292 7656 21304
rect 7708 21292 7714 21344
rect 7834 21292 7840 21344
rect 7892 21292 7898 21344
rect 8570 21292 8576 21344
rect 8628 21292 8634 21344
rect 9582 21292 9588 21344
rect 9640 21332 9646 21344
rect 11238 21332 11244 21344
rect 9640 21304 11244 21332
rect 9640 21292 9646 21304
rect 11238 21292 11244 21304
rect 11296 21292 11302 21344
rect 552 21242 11132 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 10722 21242
rect 10774 21190 10786 21242
rect 10838 21190 10850 21242
rect 10902 21190 10914 21242
rect 10966 21190 10978 21242
rect 11030 21190 11132 21242
rect 552 21168 11132 21190
rect 1302 21088 1308 21140
rect 1360 21088 1366 21140
rect 1854 21088 1860 21140
rect 1912 21088 1918 21140
rect 2130 21088 2136 21140
rect 2188 21128 2194 21140
rect 2498 21128 2504 21140
rect 2188 21100 2504 21128
rect 2188 21088 2194 21100
rect 2498 21088 2504 21100
rect 2556 21128 2562 21140
rect 2556 21100 4384 21128
rect 2556 21088 2562 21100
rect 3234 21060 3240 21072
rect 1780 21032 3240 21060
rect 1394 20952 1400 21004
rect 1452 20992 1458 21004
rect 1489 20995 1547 21001
rect 1489 20992 1501 20995
rect 1452 20964 1501 20992
rect 1452 20952 1458 20964
rect 1489 20961 1501 20964
rect 1535 20961 1547 20995
rect 1489 20955 1547 20961
rect 1670 20952 1676 21004
rect 1728 20952 1734 21004
rect 1780 21001 1808 21032
rect 3234 21020 3240 21032
rect 3292 21020 3298 21072
rect 3326 21020 3332 21072
rect 3384 21020 3390 21072
rect 3786 21020 3792 21072
rect 3844 21060 3850 21072
rect 3844 21032 4200 21060
rect 3844 21020 3850 21032
rect 1765 20995 1823 21001
rect 1765 20961 1777 20995
rect 1811 20961 1823 20995
rect 1765 20955 1823 20961
rect 2038 20952 2044 21004
rect 2096 20952 2102 21004
rect 2314 20952 2320 21004
rect 2372 20952 2378 21004
rect 2498 20952 2504 21004
rect 2556 20992 2562 21004
rect 2593 20995 2651 21001
rect 2593 20992 2605 20995
rect 2556 20964 2605 20992
rect 2556 20952 2562 20964
rect 2593 20961 2605 20964
rect 2639 20961 2651 20995
rect 2593 20955 2651 20961
rect 2682 20952 2688 21004
rect 2740 20992 2746 21004
rect 2777 20995 2835 21001
rect 2777 20992 2789 20995
rect 2740 20964 2789 20992
rect 2740 20952 2746 20964
rect 2777 20961 2789 20964
rect 2823 20961 2835 20995
rect 2777 20955 2835 20961
rect 3142 20952 3148 21004
rect 3200 20952 3206 21004
rect 3418 20952 3424 21004
rect 3476 20992 3482 21004
rect 3602 20992 3608 21004
rect 3476 20964 3608 20992
rect 3476 20952 3482 20964
rect 3602 20952 3608 20964
rect 3660 20952 3666 21004
rect 3694 20952 3700 21004
rect 3752 20952 3758 21004
rect 3878 20952 3884 21004
rect 3936 20952 3942 21004
rect 4062 20952 4068 21004
rect 4120 20952 4126 21004
rect 4172 21001 4200 21032
rect 4356 21001 4384 21100
rect 4706 21088 4712 21140
rect 4764 21128 4770 21140
rect 7006 21128 7012 21140
rect 4764 21100 5028 21128
rect 4764 21088 4770 21100
rect 4798 21020 4804 21072
rect 4856 21020 4862 21072
rect 5000 21069 5028 21100
rect 5644 21100 7012 21128
rect 4985 21063 5043 21069
rect 4985 21029 4997 21063
rect 5031 21060 5043 21063
rect 5534 21060 5540 21072
rect 5031 21032 5540 21060
rect 5031 21029 5043 21032
rect 4985 21023 5043 21029
rect 5534 21020 5540 21032
rect 5592 21020 5598 21072
rect 4157 20995 4215 21001
rect 4157 20961 4169 20995
rect 4203 20961 4215 20995
rect 4157 20955 4215 20961
rect 4341 20995 4399 21001
rect 4341 20961 4353 20995
rect 4387 20961 4399 20995
rect 4341 20955 4399 20961
rect 4890 20952 4896 21004
rect 4948 20992 4954 21004
rect 5077 20995 5135 21001
rect 5077 20992 5089 20995
rect 4948 20964 5089 20992
rect 4948 20952 4954 20964
rect 5077 20961 5089 20964
rect 5123 20961 5135 20995
rect 5077 20955 5135 20961
rect 5261 20995 5319 21001
rect 5261 20961 5273 20995
rect 5307 20992 5319 20995
rect 5442 20992 5448 21004
rect 5307 20964 5448 20992
rect 5307 20961 5319 20964
rect 5261 20955 5319 20961
rect 5442 20952 5448 20964
rect 5500 20952 5506 21004
rect 5644 21001 5672 21100
rect 5813 21063 5871 21069
rect 5813 21029 5825 21063
rect 5859 21060 5871 21063
rect 6362 21060 6368 21072
rect 5859 21032 6368 21060
rect 5859 21029 5871 21032
rect 5813 21023 5871 21029
rect 6362 21020 6368 21032
rect 6420 21020 6426 21072
rect 6492 21060 6520 21100
rect 7006 21088 7012 21100
rect 7064 21088 7070 21140
rect 7101 21131 7159 21137
rect 7101 21097 7113 21131
rect 7147 21128 7159 21131
rect 7742 21128 7748 21140
rect 7147 21100 7748 21128
rect 7147 21097 7159 21100
rect 7101 21091 7159 21097
rect 7742 21088 7748 21100
rect 7800 21088 7806 21140
rect 9858 21088 9864 21140
rect 9916 21128 9922 21140
rect 10137 21131 10195 21137
rect 10137 21128 10149 21131
rect 9916 21100 10149 21128
rect 9916 21088 9922 21100
rect 10137 21097 10149 21100
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 10502 21088 10508 21140
rect 10560 21128 10566 21140
rect 11238 21128 11244 21140
rect 10560 21100 11244 21128
rect 10560 21088 10566 21100
rect 11238 21088 11244 21100
rect 11296 21088 11302 21140
rect 6492 21032 6592 21060
rect 5629 20995 5687 21001
rect 5629 20961 5641 20995
rect 5675 20961 5687 20995
rect 5629 20955 5687 20961
rect 5718 20952 5724 21004
rect 5776 20992 5782 21004
rect 5994 20992 6000 21004
rect 5776 20964 6000 20992
rect 5776 20952 5782 20964
rect 5994 20952 6000 20964
rect 6052 20952 6058 21004
rect 6564 21001 6592 21032
rect 6730 21020 6736 21072
rect 6788 21060 6794 21072
rect 8570 21060 8576 21072
rect 6788 21032 8576 21060
rect 6788 21020 6794 21032
rect 6181 20995 6239 21001
rect 6181 20961 6193 20995
rect 6227 20992 6239 20995
rect 6273 20995 6331 21001
rect 6273 20992 6285 20995
rect 6227 20964 6285 20992
rect 6227 20961 6239 20964
rect 6181 20955 6239 20961
rect 6273 20961 6285 20964
rect 6319 20961 6331 20995
rect 6273 20955 6331 20961
rect 6457 20995 6515 21001
rect 6457 20961 6469 20995
rect 6503 20961 6515 20995
rect 6457 20955 6515 20961
rect 6549 20995 6607 21001
rect 6549 20961 6561 20995
rect 6595 20961 6607 20995
rect 6549 20955 6607 20961
rect 6825 20995 6883 21001
rect 6825 20961 6837 20995
rect 6871 20992 6883 20995
rect 6871 20990 7052 20992
rect 6871 20964 7063 20990
rect 6871 20961 6883 20964
rect 7024 20962 7063 20964
rect 6825 20955 6883 20961
rect 2869 20927 2927 20933
rect 2869 20893 2881 20927
rect 2915 20893 2927 20927
rect 2869 20887 2927 20893
rect 2225 20859 2283 20865
rect 2225 20825 2237 20859
rect 2271 20856 2283 20859
rect 2884 20856 2912 20887
rect 2958 20884 2964 20936
rect 3016 20884 3022 20936
rect 3896 20924 3924 20952
rect 4246 20924 4252 20936
rect 3896 20896 4252 20924
rect 4246 20884 4252 20896
rect 4304 20884 4310 20936
rect 5350 20884 5356 20936
rect 5408 20884 5414 20936
rect 3142 20856 3148 20868
rect 2271 20828 2853 20856
rect 2884 20828 3148 20856
rect 2271 20825 2283 20828
rect 2225 20819 2283 20825
rect 1578 20748 1584 20800
rect 1636 20788 1642 20800
rect 2409 20791 2467 20797
rect 2409 20788 2421 20791
rect 1636 20760 2421 20788
rect 1636 20748 1642 20760
rect 2409 20757 2421 20760
rect 2455 20757 2467 20791
rect 2825 20788 2853 20828
rect 3142 20816 3148 20828
rect 3200 20816 3206 20868
rect 3326 20816 3332 20868
rect 3384 20856 3390 20868
rect 3789 20859 3847 20865
rect 3384 20828 3556 20856
rect 3384 20816 3390 20828
rect 3421 20791 3479 20797
rect 3421 20788 3433 20791
rect 2825 20760 3433 20788
rect 2409 20751 2467 20757
rect 3421 20757 3433 20760
rect 3467 20757 3479 20791
rect 3528 20788 3556 20828
rect 3789 20825 3801 20859
rect 3835 20856 3847 20859
rect 5261 20859 5319 20865
rect 5261 20856 5273 20859
rect 3835 20828 5273 20856
rect 3835 20825 3847 20828
rect 3789 20819 3847 20825
rect 5261 20825 5273 20828
rect 5307 20825 5319 20859
rect 5261 20819 5319 20825
rect 5442 20816 5448 20868
rect 5500 20816 5506 20868
rect 6472 20856 6500 20955
rect 6641 20927 6699 20933
rect 6641 20893 6653 20927
rect 6687 20924 6699 20927
rect 6914 20924 6920 20936
rect 6687 20896 6920 20924
rect 6687 20893 6699 20896
rect 6641 20887 6699 20893
rect 6730 20856 6736 20868
rect 6472 20828 6736 20856
rect 6730 20816 6736 20828
rect 6788 20816 6794 20868
rect 4525 20791 4583 20797
rect 4525 20788 4537 20791
rect 3528 20760 4537 20788
rect 3421 20751 3479 20757
rect 4525 20757 4537 20760
rect 4571 20757 4583 20791
rect 4525 20751 4583 20757
rect 4617 20791 4675 20797
rect 4617 20757 4629 20791
rect 4663 20788 4675 20791
rect 4706 20788 4712 20800
rect 4663 20760 4712 20788
rect 4663 20757 4675 20760
rect 4617 20751 4675 20757
rect 4706 20748 4712 20760
rect 4764 20748 4770 20800
rect 5537 20791 5595 20797
rect 5537 20757 5549 20791
rect 5583 20788 5595 20791
rect 6831 20788 6859 20896
rect 6914 20884 6920 20896
rect 6972 20884 6978 20936
rect 7035 20924 7063 20962
rect 7282 20952 7288 21004
rect 7340 20952 7346 21004
rect 7466 20952 7472 21004
rect 7524 20952 7530 21004
rect 7668 21001 7696 21032
rect 8570 21020 8576 21032
rect 8628 21020 8634 21072
rect 9122 21020 9128 21072
rect 9180 21060 9186 21072
rect 9180 21032 10272 21060
rect 9180 21020 9186 21032
rect 7653 20995 7711 21001
rect 7653 20961 7665 20995
rect 7699 20961 7711 20995
rect 7653 20955 7711 20961
rect 7834 20952 7840 21004
rect 7892 20952 7898 21004
rect 9217 20995 9275 21001
rect 9217 20961 9229 20995
rect 9263 20961 9275 20995
rect 9217 20955 9275 20961
rect 7190 20924 7196 20936
rect 7035 20896 7196 20924
rect 7190 20884 7196 20896
rect 7248 20924 7254 20936
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 7248 20896 7573 20924
rect 7248 20884 7254 20896
rect 7561 20893 7573 20896
rect 7607 20924 7619 20927
rect 8018 20924 8024 20936
rect 7607 20896 8024 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 8018 20884 8024 20896
rect 8076 20884 8082 20936
rect 8846 20884 8852 20936
rect 8904 20884 8910 20936
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20924 8999 20927
rect 9122 20924 9128 20936
rect 8987 20896 9128 20924
rect 8987 20893 8999 20896
rect 8941 20887 8999 20893
rect 9122 20884 9128 20896
rect 9180 20884 9186 20936
rect 8386 20816 8392 20868
rect 8444 20856 8450 20868
rect 8757 20859 8815 20865
rect 8757 20856 8769 20859
rect 8444 20828 8769 20856
rect 8444 20816 8450 20828
rect 8757 20825 8769 20828
rect 8803 20825 8815 20859
rect 9232 20856 9260 20955
rect 9324 20924 9352 21032
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 10244 21001 10272 21032
rect 9493 20995 9551 21001
rect 9493 20992 9505 20995
rect 9456 20964 9505 20992
rect 9456 20952 9462 20964
rect 9493 20961 9505 20964
rect 9539 20992 9551 20995
rect 9953 20995 10011 21001
rect 9953 20992 9965 20995
rect 9539 20964 9965 20992
rect 9539 20961 9551 20964
rect 9493 20955 9551 20961
rect 9953 20961 9965 20964
rect 9999 20961 10011 20995
rect 9953 20955 10011 20961
rect 10229 20995 10287 21001
rect 10229 20961 10241 20995
rect 10275 20961 10287 20995
rect 10229 20955 10287 20961
rect 9585 20927 9643 20933
rect 9585 20924 9597 20927
rect 9324 20896 9597 20924
rect 9585 20893 9597 20896
rect 9631 20893 9643 20927
rect 9585 20887 9643 20893
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20893 9735 20927
rect 9677 20887 9735 20893
rect 9769 20927 9827 20933
rect 9769 20893 9781 20927
rect 9815 20924 9827 20927
rect 10042 20924 10048 20936
rect 9815 20896 10048 20924
rect 9815 20893 9827 20896
rect 9769 20887 9827 20893
rect 9692 20856 9720 20887
rect 10042 20884 10048 20896
rect 10100 20884 10106 20936
rect 9858 20856 9864 20868
rect 9232 20828 9628 20856
rect 9692 20828 9864 20856
rect 8757 20819 8815 20825
rect 5583 20760 6859 20788
rect 7009 20791 7067 20797
rect 5583 20757 5595 20760
rect 5537 20751 5595 20757
rect 7009 20757 7021 20791
rect 7055 20788 7067 20791
rect 7098 20788 7104 20800
rect 7055 20760 7104 20788
rect 7055 20757 7067 20760
rect 7009 20751 7067 20757
rect 7098 20748 7104 20760
rect 7156 20748 7162 20800
rect 9125 20791 9183 20797
rect 9125 20757 9137 20791
rect 9171 20788 9183 20791
rect 9309 20791 9367 20797
rect 9309 20788 9321 20791
rect 9171 20760 9321 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 9309 20757 9321 20760
rect 9355 20757 9367 20791
rect 9600 20788 9628 20828
rect 9858 20816 9864 20828
rect 9916 20816 9922 20868
rect 9674 20788 9680 20800
rect 9600 20760 9680 20788
rect 9309 20751 9367 20757
rect 9674 20748 9680 20760
rect 9732 20788 9738 20800
rect 9953 20791 10011 20797
rect 9953 20788 9965 20791
rect 9732 20760 9965 20788
rect 9732 20748 9738 20760
rect 9953 20757 9965 20760
rect 9999 20757 10011 20791
rect 9953 20751 10011 20757
rect 552 20698 11132 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 10062 20698
rect 10114 20646 10126 20698
rect 10178 20646 10190 20698
rect 10242 20646 10254 20698
rect 10306 20646 10318 20698
rect 10370 20646 11132 20698
rect 552 20624 11132 20646
rect 2590 20544 2596 20596
rect 2648 20584 2654 20596
rect 2685 20587 2743 20593
rect 2685 20584 2697 20587
rect 2648 20556 2697 20584
rect 2648 20544 2654 20556
rect 2685 20553 2697 20556
rect 2731 20553 2743 20587
rect 2685 20547 2743 20553
rect 3510 20544 3516 20596
rect 3568 20584 3574 20596
rect 5445 20587 5503 20593
rect 5445 20584 5457 20587
rect 3568 20556 5457 20584
rect 3568 20544 3574 20556
rect 5445 20553 5457 20556
rect 5491 20553 5503 20587
rect 5445 20547 5503 20553
rect 5537 20587 5595 20593
rect 5537 20553 5549 20587
rect 5583 20584 5595 20587
rect 5994 20584 6000 20596
rect 5583 20556 6000 20584
rect 5583 20553 5595 20556
rect 5537 20547 5595 20553
rect 5994 20544 6000 20556
rect 6052 20584 6058 20596
rect 6546 20584 6552 20596
rect 6052 20556 6552 20584
rect 6052 20544 6058 20556
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 7469 20587 7527 20593
rect 7469 20584 7481 20587
rect 6972 20556 7481 20584
rect 6972 20544 6978 20556
rect 7469 20553 7481 20556
rect 7515 20553 7527 20587
rect 7469 20547 7527 20553
rect 7650 20544 7656 20596
rect 7708 20544 7714 20596
rect 9398 20544 9404 20596
rect 9456 20544 9462 20596
rect 1670 20476 1676 20528
rect 1728 20516 1734 20528
rect 3237 20519 3295 20525
rect 3237 20516 3249 20519
rect 1728 20488 3249 20516
rect 1728 20476 1734 20488
rect 3237 20485 3249 20488
rect 3283 20485 3295 20519
rect 3237 20479 3295 20485
rect 3418 20476 3424 20528
rect 3476 20476 3482 20528
rect 4157 20519 4215 20525
rect 4157 20485 4169 20519
rect 4203 20516 4215 20519
rect 4246 20516 4252 20528
rect 4203 20488 4252 20516
rect 4203 20485 4215 20488
rect 4157 20479 4215 20485
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 5718 20476 5724 20528
rect 5776 20516 5782 20528
rect 5776 20488 7696 20516
rect 5776 20476 5782 20488
rect 1213 20451 1271 20457
rect 1213 20417 1225 20451
rect 1259 20448 1271 20451
rect 1394 20448 1400 20460
rect 1259 20420 1400 20448
rect 1259 20417 1271 20420
rect 1213 20411 1271 20417
rect 1394 20408 1400 20420
rect 1452 20408 1458 20460
rect 1578 20408 1584 20460
rect 1636 20448 1642 20460
rect 1765 20451 1823 20457
rect 1765 20448 1777 20451
rect 1636 20420 1777 20448
rect 1636 20408 1642 20420
rect 1765 20417 1777 20420
rect 1811 20417 1823 20451
rect 3436 20448 3464 20476
rect 4617 20451 4675 20457
rect 3436 20420 4552 20448
rect 1765 20411 1823 20417
rect 2038 20340 2044 20392
rect 2096 20340 2102 20392
rect 2222 20340 2228 20392
rect 2280 20340 2286 20392
rect 2498 20340 2504 20392
rect 2556 20340 2562 20392
rect 2774 20340 2780 20392
rect 2832 20340 2838 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 2876 20352 3433 20380
rect 1210 20272 1216 20324
rect 1268 20312 1274 20324
rect 2876 20312 2904 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 3694 20340 3700 20392
rect 3752 20340 3758 20392
rect 4062 20340 4068 20392
rect 4120 20340 4126 20392
rect 4246 20340 4252 20392
rect 4304 20380 4310 20392
rect 4341 20383 4399 20389
rect 4341 20380 4353 20383
rect 4304 20352 4353 20380
rect 4304 20340 4310 20352
rect 4341 20349 4353 20352
rect 4387 20349 4399 20383
rect 4341 20343 4399 20349
rect 4433 20383 4491 20389
rect 4433 20349 4445 20383
rect 4479 20349 4491 20383
rect 4433 20343 4491 20349
rect 1268 20284 2904 20312
rect 1268 20272 1274 20284
rect 3326 20272 3332 20324
rect 3384 20312 3390 20324
rect 3605 20315 3663 20321
rect 3605 20312 3617 20315
rect 3384 20284 3617 20312
rect 3384 20272 3390 20284
rect 3605 20281 3617 20284
rect 3651 20281 3663 20315
rect 3605 20275 3663 20281
rect 3970 20272 3976 20324
rect 4028 20312 4034 20324
rect 4448 20312 4476 20343
rect 4028 20284 4476 20312
rect 4524 20312 4552 20420
rect 4617 20417 4629 20451
rect 4663 20448 4675 20451
rect 5353 20451 5411 20457
rect 5353 20448 5365 20451
rect 4663 20420 5365 20448
rect 4663 20417 4675 20420
rect 4617 20411 4675 20417
rect 5353 20417 5365 20420
rect 5399 20417 5411 20451
rect 6457 20451 6515 20457
rect 5353 20411 5411 20417
rect 5644 20420 6040 20448
rect 4798 20340 4804 20392
rect 4856 20380 4862 20392
rect 4893 20383 4951 20389
rect 4893 20380 4905 20383
rect 4856 20352 4905 20380
rect 4856 20340 4862 20352
rect 4893 20349 4905 20352
rect 4939 20349 4951 20383
rect 4893 20343 4951 20349
rect 4982 20340 4988 20392
rect 5040 20340 5046 20392
rect 5077 20383 5135 20389
rect 5077 20349 5089 20383
rect 5123 20349 5135 20383
rect 5077 20343 5135 20349
rect 5092 20312 5120 20343
rect 5166 20340 5172 20392
rect 5224 20340 5230 20392
rect 5644 20389 5672 20420
rect 5629 20383 5687 20389
rect 5629 20349 5641 20383
rect 5675 20349 5687 20383
rect 5629 20343 5687 20349
rect 5810 20340 5816 20392
rect 5868 20340 5874 20392
rect 5828 20312 5856 20340
rect 4524 20284 4844 20312
rect 5092 20284 5856 20312
rect 4028 20272 4034 20284
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 2317 20247 2375 20253
rect 2317 20244 2329 20247
rect 1820 20216 2329 20244
rect 1820 20204 1826 20216
rect 2317 20213 2329 20216
rect 2363 20213 2375 20247
rect 2317 20207 2375 20213
rect 3510 20204 3516 20256
rect 3568 20244 3574 20256
rect 4709 20247 4767 20253
rect 4709 20244 4721 20247
rect 3568 20216 4721 20244
rect 3568 20204 3574 20216
rect 4709 20213 4721 20216
rect 4755 20213 4767 20247
rect 4816 20244 4844 20284
rect 5718 20244 5724 20256
rect 4816 20216 5724 20244
rect 4709 20207 4767 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 5810 20204 5816 20256
rect 5868 20204 5874 20256
rect 6012 20244 6040 20420
rect 6457 20417 6469 20451
rect 6503 20448 6515 20451
rect 6546 20448 6552 20460
rect 6503 20420 6552 20448
rect 6503 20417 6515 20420
rect 6457 20411 6515 20417
rect 6546 20408 6552 20420
rect 6604 20408 6610 20460
rect 6825 20451 6883 20457
rect 6825 20417 6837 20451
rect 6871 20448 6883 20451
rect 7098 20448 7104 20460
rect 6871 20420 7104 20448
rect 6871 20417 6883 20420
rect 6825 20411 6883 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 7668 20389 7696 20488
rect 9140 20488 10364 20516
rect 7837 20451 7895 20457
rect 7837 20417 7849 20451
rect 7883 20448 7895 20451
rect 9033 20451 9091 20457
rect 9033 20448 9045 20451
rect 7883 20420 9045 20448
rect 7883 20417 7895 20420
rect 7837 20411 7895 20417
rect 9033 20417 9045 20420
rect 9079 20417 9091 20451
rect 9033 20411 9091 20417
rect 6181 20383 6239 20389
rect 6181 20349 6193 20383
rect 6227 20380 6239 20383
rect 7653 20383 7711 20389
rect 6227 20352 7052 20380
rect 6227 20349 6239 20352
rect 6181 20343 6239 20349
rect 6086 20272 6092 20324
rect 6144 20312 6150 20324
rect 6273 20315 6331 20321
rect 6273 20312 6285 20315
rect 6144 20284 6285 20312
rect 6144 20272 6150 20284
rect 6273 20281 6285 20284
rect 6319 20312 6331 20315
rect 6917 20315 6975 20321
rect 6917 20312 6929 20315
rect 6319 20284 6929 20312
rect 6319 20281 6331 20284
rect 6273 20275 6331 20281
rect 6917 20281 6929 20284
rect 6963 20281 6975 20315
rect 6917 20275 6975 20281
rect 6822 20244 6828 20256
rect 6012 20216 6828 20244
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7024 20253 7052 20352
rect 7653 20349 7665 20383
rect 7699 20349 7711 20383
rect 7653 20343 7711 20349
rect 8478 20340 8484 20392
rect 8536 20340 8542 20392
rect 8570 20340 8576 20392
rect 8628 20380 8634 20392
rect 9140 20389 9168 20488
rect 9490 20408 9496 20460
rect 9548 20448 9554 20460
rect 10336 20457 10364 20488
rect 9677 20451 9735 20457
rect 9677 20448 9689 20451
rect 9548 20420 9689 20448
rect 9548 20408 9554 20420
rect 9677 20417 9689 20420
rect 9723 20417 9735 20451
rect 9677 20411 9735 20417
rect 10321 20451 10379 20457
rect 10321 20417 10333 20451
rect 10367 20448 10379 20451
rect 10502 20448 10508 20460
rect 10367 20420 10508 20448
rect 10367 20417 10379 20420
rect 10321 20411 10379 20417
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 8941 20383 8999 20389
rect 8941 20380 8953 20383
rect 8628 20352 8953 20380
rect 8628 20340 8634 20352
rect 8941 20349 8953 20352
rect 8987 20349 8999 20383
rect 8941 20343 8999 20349
rect 9125 20383 9183 20389
rect 9125 20349 9137 20383
rect 9171 20349 9183 20383
rect 9125 20343 9183 20349
rect 9766 20340 9772 20392
rect 9824 20340 9830 20392
rect 10413 20383 10471 20389
rect 10413 20349 10425 20383
rect 10459 20380 10471 20383
rect 11330 20380 11336 20392
rect 10459 20352 11336 20380
rect 10459 20349 10471 20352
rect 10413 20343 10471 20349
rect 7929 20315 7987 20321
rect 7929 20312 7941 20315
rect 7392 20284 7941 20312
rect 7009 20247 7067 20253
rect 7009 20213 7021 20247
rect 7055 20244 7067 20247
rect 7282 20244 7288 20256
rect 7055 20216 7288 20244
rect 7055 20213 7067 20216
rect 7009 20207 7067 20213
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 7392 20253 7420 20284
rect 7929 20281 7941 20284
rect 7975 20281 7987 20315
rect 7929 20275 7987 20281
rect 8018 20272 8024 20324
rect 8076 20312 8082 20324
rect 10428 20312 10456 20343
rect 11330 20340 11336 20352
rect 11388 20340 11394 20392
rect 8076 20284 10456 20312
rect 8076 20272 8082 20284
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20213 7435 20247
rect 7377 20207 7435 20213
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 8573 20247 8631 20253
rect 8573 20244 8585 20247
rect 7524 20216 8585 20244
rect 7524 20204 7530 20216
rect 8573 20213 8585 20216
rect 8619 20213 8631 20247
rect 8573 20207 8631 20213
rect 9766 20204 9772 20256
rect 9824 20244 9830 20256
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 9824 20216 10057 20244
rect 9824 20204 9830 20216
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 10045 20207 10103 20213
rect 552 20154 11132 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 10722 20154
rect 10774 20102 10786 20154
rect 10838 20102 10850 20154
rect 10902 20102 10914 20154
rect 10966 20102 10978 20154
rect 11030 20102 11132 20154
rect 552 20080 11132 20102
rect 1946 20000 1952 20052
rect 2004 20040 2010 20052
rect 2593 20043 2651 20049
rect 2593 20040 2605 20043
rect 2004 20012 2605 20040
rect 2004 20000 2010 20012
rect 2593 20009 2605 20012
rect 2639 20009 2651 20043
rect 2593 20003 2651 20009
rect 3145 20043 3203 20049
rect 3145 20009 3157 20043
rect 3191 20040 3203 20043
rect 3234 20040 3240 20052
rect 3191 20012 3240 20040
rect 3191 20009 3203 20012
rect 3145 20003 3203 20009
rect 3234 20000 3240 20012
rect 3292 20000 3298 20052
rect 3326 20000 3332 20052
rect 3384 20040 3390 20052
rect 3513 20043 3571 20049
rect 3513 20040 3525 20043
rect 3384 20012 3525 20040
rect 3384 20000 3390 20012
rect 3513 20009 3525 20012
rect 3559 20040 3571 20043
rect 3694 20040 3700 20052
rect 3559 20012 3700 20040
rect 3559 20009 3571 20012
rect 3513 20003 3571 20009
rect 3694 20000 3700 20012
rect 3752 20000 3758 20052
rect 4522 20040 4528 20052
rect 4264 20012 4528 20040
rect 1670 19932 1676 19984
rect 1728 19972 1734 19984
rect 2498 19972 2504 19984
rect 1728 19944 2504 19972
rect 1728 19932 1734 19944
rect 2498 19932 2504 19944
rect 2556 19932 2562 19984
rect 2866 19972 2872 19984
rect 2608 19944 2872 19972
rect 2608 19916 2636 19944
rect 2866 19932 2872 19944
rect 2924 19972 2930 19984
rect 2924 19944 3372 19972
rect 2924 19932 2930 19944
rect 1578 19864 1584 19916
rect 1636 19904 1642 19916
rect 1765 19907 1823 19913
rect 1765 19904 1777 19907
rect 1636 19876 1777 19904
rect 1636 19864 1642 19876
rect 1765 19873 1777 19876
rect 1811 19873 1823 19907
rect 1765 19867 1823 19873
rect 2041 19907 2099 19913
rect 2041 19873 2053 19907
rect 2087 19904 2099 19907
rect 2314 19904 2320 19916
rect 2087 19876 2320 19904
rect 2087 19873 2099 19876
rect 2041 19867 2099 19873
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 2590 19864 2596 19916
rect 2648 19864 2654 19916
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 3142 19904 3148 19916
rect 2832 19876 3148 19904
rect 2832 19864 2838 19876
rect 3142 19864 3148 19876
rect 3200 19864 3206 19916
rect 3344 19913 3372 19944
rect 3970 19932 3976 19984
rect 4028 19972 4034 19984
rect 4264 19972 4292 20012
rect 4522 20000 4528 20012
rect 4580 20000 4586 20052
rect 4798 20000 4804 20052
rect 4856 20000 4862 20052
rect 5166 20000 5172 20052
rect 5224 20000 5230 20052
rect 5261 20043 5319 20049
rect 5261 20009 5273 20043
rect 5307 20040 5319 20043
rect 5626 20040 5632 20052
rect 5307 20012 5632 20040
rect 5307 20009 5319 20012
rect 5261 20003 5319 20009
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 4028 19944 4292 19972
rect 4028 19932 4034 19944
rect 3329 19907 3387 19913
rect 3329 19873 3341 19907
rect 3375 19873 3387 19907
rect 3329 19867 3387 19873
rect 3605 19907 3663 19913
rect 3605 19873 3617 19907
rect 3651 19904 3663 19907
rect 3881 19907 3939 19913
rect 3651 19876 3832 19904
rect 3651 19873 3663 19876
rect 3605 19867 3663 19873
rect 1210 19796 1216 19848
rect 1268 19796 1274 19848
rect 2222 19796 2228 19848
rect 2280 19796 2286 19848
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19836 3111 19839
rect 3234 19836 3240 19848
rect 3099 19808 3240 19836
rect 3099 19805 3111 19808
rect 3053 19799 3111 19805
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 2406 19728 2412 19780
rect 2464 19768 2470 19780
rect 2961 19771 3019 19777
rect 2961 19768 2973 19771
rect 2464 19740 2973 19768
rect 2464 19728 2470 19740
rect 2961 19737 2973 19740
rect 3007 19768 3019 19771
rect 3697 19771 3755 19777
rect 3697 19768 3709 19771
rect 3007 19740 3709 19768
rect 3007 19737 3019 19740
rect 2961 19731 3019 19737
rect 3697 19737 3709 19740
rect 3743 19737 3755 19771
rect 3697 19731 3755 19737
rect 1026 19660 1032 19712
rect 1084 19700 1090 19712
rect 2682 19700 2688 19712
rect 1084 19672 2688 19700
rect 1084 19660 1090 19672
rect 2682 19660 2688 19672
rect 2740 19660 2746 19712
rect 3804 19700 3832 19876
rect 3881 19873 3893 19907
rect 3927 19873 3939 19907
rect 3881 19867 3939 19873
rect 3896 19768 3924 19867
rect 4154 19864 4160 19916
rect 4212 19864 4218 19916
rect 4264 19913 4292 19944
rect 4617 19975 4675 19981
rect 4617 19941 4629 19975
rect 4663 19972 4675 19975
rect 5184 19972 5212 20000
rect 6086 19972 6092 19984
rect 4663 19944 5212 19972
rect 5828 19944 6092 19972
rect 4663 19941 4675 19944
rect 4617 19935 4675 19941
rect 4249 19907 4307 19913
rect 4249 19873 4261 19907
rect 4295 19873 4307 19907
rect 4249 19867 4307 19873
rect 4430 19864 4436 19916
rect 4488 19864 4494 19916
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19904 4583 19907
rect 4709 19907 4767 19913
rect 4571 19876 4660 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 4062 19796 4068 19848
rect 4120 19796 4126 19848
rect 4246 19768 4252 19780
rect 3896 19740 4252 19768
rect 4246 19728 4252 19740
rect 4304 19728 4310 19780
rect 4632 19768 4660 19876
rect 4709 19873 4721 19907
rect 4755 19873 4767 19907
rect 4709 19867 4767 19873
rect 5169 19907 5227 19913
rect 5169 19873 5181 19907
rect 5215 19904 5227 19907
rect 5828 19904 5856 19944
rect 6086 19932 6092 19944
rect 6144 19932 6150 19984
rect 6546 19932 6552 19984
rect 6604 19932 6610 19984
rect 7745 19975 7803 19981
rect 6656 19944 7420 19972
rect 5215 19876 5856 19904
rect 5215 19873 5227 19876
rect 5169 19867 5227 19873
rect 4724 19836 4752 19867
rect 5902 19864 5908 19916
rect 5960 19904 5966 19916
rect 6273 19907 6331 19913
rect 6273 19904 6285 19907
rect 5960 19876 6285 19904
rect 5960 19864 5966 19876
rect 6273 19873 6285 19876
rect 6319 19873 6331 19907
rect 6273 19867 6331 19873
rect 6365 19907 6423 19913
rect 6365 19873 6377 19907
rect 6411 19904 6423 19907
rect 6656 19904 6684 19944
rect 6411 19876 6684 19904
rect 6733 19907 6791 19913
rect 6411 19873 6423 19876
rect 6365 19867 6423 19873
rect 6733 19873 6745 19907
rect 6779 19873 6791 19907
rect 6733 19867 6791 19873
rect 5442 19836 5448 19848
rect 4724 19808 5448 19836
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 6089 19839 6147 19845
rect 6089 19805 6101 19839
rect 6135 19805 6147 19839
rect 6089 19799 6147 19805
rect 4890 19768 4896 19780
rect 4632 19740 4896 19768
rect 4890 19728 4896 19740
rect 4948 19728 4954 19780
rect 5905 19703 5963 19709
rect 5905 19700 5917 19703
rect 3804 19672 5917 19700
rect 5905 19669 5917 19672
rect 5951 19669 5963 19703
rect 6104 19700 6132 19799
rect 6178 19796 6184 19848
rect 6236 19796 6242 19848
rect 6748 19768 6776 19867
rect 6822 19864 6828 19916
rect 6880 19904 6886 19916
rect 7098 19904 7104 19916
rect 6880 19876 7104 19904
rect 6880 19864 6886 19876
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 7190 19864 7196 19916
rect 7248 19904 7254 19916
rect 7285 19907 7343 19913
rect 7285 19904 7297 19907
rect 7248 19876 7297 19904
rect 7248 19864 7254 19876
rect 7285 19873 7297 19876
rect 7331 19873 7343 19907
rect 7392 19904 7420 19944
rect 7745 19941 7757 19975
rect 7791 19972 7803 19975
rect 7926 19972 7932 19984
rect 7791 19944 7932 19972
rect 7791 19941 7803 19944
rect 7745 19935 7803 19941
rect 7926 19932 7932 19944
rect 7984 19932 7990 19984
rect 8662 19972 8668 19984
rect 8404 19944 8668 19972
rect 8205 19907 8263 19913
rect 8205 19904 8217 19907
rect 7392 19876 8217 19904
rect 7285 19867 7343 19873
rect 8205 19873 8217 19876
rect 8251 19873 8263 19907
rect 8205 19867 8263 19873
rect 8294 19864 8300 19916
rect 8352 19904 8358 19916
rect 8404 19913 8432 19944
rect 8662 19932 8668 19944
rect 8720 19932 8726 19984
rect 9677 19975 9735 19981
rect 9677 19941 9689 19975
rect 9723 19972 9735 19975
rect 9766 19972 9772 19984
rect 9723 19944 9772 19972
rect 9723 19941 9735 19944
rect 9677 19935 9735 19941
rect 9766 19932 9772 19944
rect 9824 19932 9830 19984
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 8352 19876 8401 19904
rect 8352 19864 8358 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 8941 19907 8999 19913
rect 8941 19873 8953 19907
rect 8987 19904 8999 19907
rect 9030 19904 9036 19916
rect 8987 19876 9036 19904
rect 8987 19873 8999 19876
rect 8941 19867 8999 19873
rect 9030 19864 9036 19876
rect 9088 19864 9094 19916
rect 9122 19864 9128 19916
rect 9180 19864 9186 19916
rect 6914 19796 6920 19848
rect 6972 19796 6978 19848
rect 7006 19796 7012 19848
rect 7064 19836 7070 19848
rect 7466 19836 7472 19848
rect 7064 19808 7472 19836
rect 7064 19796 7070 19808
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 7742 19796 7748 19848
rect 7800 19836 7806 19848
rect 7837 19839 7895 19845
rect 7837 19836 7849 19839
rect 7800 19808 7849 19836
rect 7800 19796 7806 19808
rect 7837 19805 7849 19808
rect 7883 19805 7895 19839
rect 7837 19799 7895 19805
rect 8021 19839 8079 19845
rect 8021 19805 8033 19839
rect 8067 19836 8079 19839
rect 8573 19839 8631 19845
rect 8573 19836 8585 19839
rect 8067 19808 8585 19836
rect 8067 19805 8079 19808
rect 8021 19799 8079 19805
rect 8573 19805 8585 19808
rect 8619 19805 8631 19839
rect 8573 19799 8631 19805
rect 8665 19839 8723 19845
rect 8665 19805 8677 19839
rect 8711 19805 8723 19839
rect 8665 19799 8723 19805
rect 6822 19768 6828 19780
rect 6748 19740 6828 19768
rect 6822 19728 6828 19740
rect 6880 19728 6886 19780
rect 7377 19771 7435 19777
rect 7377 19768 7389 19771
rect 6932 19740 7389 19768
rect 6932 19700 6960 19740
rect 7377 19737 7389 19740
rect 7423 19737 7435 19771
rect 7377 19731 7435 19737
rect 6104 19672 6960 19700
rect 5905 19663 5963 19669
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 7466 19700 7472 19712
rect 7340 19672 7472 19700
rect 7340 19660 7346 19672
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 7926 19660 7932 19712
rect 7984 19700 7990 19712
rect 8036 19700 8064 19799
rect 8386 19728 8392 19780
rect 8444 19768 8450 19780
rect 8680 19768 8708 19799
rect 8444 19740 8708 19768
rect 8444 19728 8450 19740
rect 9490 19728 9496 19780
rect 9548 19768 9554 19780
rect 9953 19771 10011 19777
rect 9953 19768 9965 19771
rect 9548 19740 9965 19768
rect 9548 19728 9554 19740
rect 9953 19737 9965 19740
rect 9999 19737 10011 19771
rect 9953 19731 10011 19737
rect 7984 19672 8064 19700
rect 7984 19660 7990 19672
rect 8846 19660 8852 19712
rect 8904 19700 8910 19712
rect 8941 19703 8999 19709
rect 8941 19700 8953 19703
rect 8904 19672 8953 19700
rect 8904 19660 8910 19672
rect 8941 19669 8953 19672
rect 8987 19669 8999 19703
rect 8941 19663 8999 19669
rect 10137 19703 10195 19709
rect 10137 19669 10149 19703
rect 10183 19700 10195 19703
rect 10410 19700 10416 19712
rect 10183 19672 10416 19700
rect 10183 19669 10195 19672
rect 10137 19663 10195 19669
rect 10410 19660 10416 19672
rect 10468 19660 10474 19712
rect 552 19610 11132 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 10062 19610
rect 10114 19558 10126 19610
rect 10178 19558 10190 19610
rect 10242 19558 10254 19610
rect 10306 19558 10318 19610
rect 10370 19558 11132 19610
rect 552 19536 11132 19558
rect 2038 19456 2044 19508
rect 2096 19496 2102 19508
rect 2317 19499 2375 19505
rect 2317 19496 2329 19499
rect 2096 19468 2329 19496
rect 2096 19456 2102 19468
rect 2317 19465 2329 19468
rect 2363 19465 2375 19499
rect 2317 19459 2375 19465
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 3050 19496 3056 19508
rect 2832 19468 3056 19496
rect 2832 19456 2838 19468
rect 3050 19456 3056 19468
rect 3108 19456 3114 19508
rect 3510 19456 3516 19508
rect 3568 19496 3574 19508
rect 3973 19499 4031 19505
rect 3973 19496 3985 19499
rect 3568 19468 3985 19496
rect 3568 19456 3574 19468
rect 3973 19465 3985 19468
rect 4019 19465 4031 19499
rect 3973 19459 4031 19465
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 4430 19496 4436 19508
rect 4120 19468 4436 19496
rect 4120 19456 4126 19468
rect 4430 19456 4436 19468
rect 4488 19456 4494 19508
rect 5810 19496 5816 19508
rect 5092 19468 5816 19496
rect 198 19388 204 19440
rect 256 19428 262 19440
rect 566 19428 572 19440
rect 256 19400 572 19428
rect 256 19388 262 19400
rect 566 19388 572 19400
rect 624 19388 630 19440
rect 1118 19388 1124 19440
rect 1176 19428 1182 19440
rect 1176 19400 2452 19428
rect 1176 19388 1182 19400
rect 1136 19360 1164 19388
rect 1044 19332 1164 19360
rect 1213 19363 1271 19369
rect 566 19252 572 19304
rect 624 19292 630 19304
rect 1044 19301 1072 19332
rect 1213 19329 1225 19363
rect 1259 19360 1271 19363
rect 1486 19360 1492 19372
rect 1259 19332 1492 19360
rect 1259 19329 1271 19332
rect 1213 19323 1271 19329
rect 1486 19320 1492 19332
rect 1544 19320 1550 19372
rect 1029 19295 1087 19301
rect 1029 19292 1041 19295
rect 624 19264 1041 19292
rect 624 19252 630 19264
rect 1029 19261 1041 19264
rect 1075 19261 1087 19295
rect 1029 19255 1087 19261
rect 1118 19252 1124 19304
rect 1176 19252 1182 19304
rect 1302 19252 1308 19304
rect 1360 19292 1366 19304
rect 1765 19295 1823 19301
rect 1765 19292 1777 19295
rect 1360 19264 1777 19292
rect 1360 19252 1366 19264
rect 1765 19261 1777 19264
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19261 2099 19295
rect 2041 19255 2099 19261
rect 842 19184 848 19236
rect 900 19184 906 19236
rect 952 19196 1164 19224
rect 952 19165 980 19196
rect 943 19159 1001 19165
rect 943 19125 955 19159
rect 989 19125 1001 19159
rect 1136 19156 1164 19196
rect 2056 19156 2084 19255
rect 2222 19252 2228 19304
rect 2280 19252 2286 19304
rect 1136 19128 2084 19156
rect 2424 19156 2452 19400
rect 2682 19388 2688 19440
rect 2740 19428 2746 19440
rect 3605 19431 3663 19437
rect 3605 19428 3617 19431
rect 2740 19400 3617 19428
rect 2740 19388 2746 19400
rect 3605 19397 3617 19400
rect 3651 19397 3663 19431
rect 3605 19391 3663 19397
rect 3694 19388 3700 19440
rect 3752 19428 3758 19440
rect 4522 19428 4528 19440
rect 3752 19400 4528 19428
rect 3752 19388 3758 19400
rect 4522 19388 4528 19400
rect 4580 19388 4586 19440
rect 2590 19320 2596 19372
rect 2648 19360 2654 19372
rect 2777 19363 2835 19369
rect 2777 19360 2789 19363
rect 2648 19332 2789 19360
rect 2648 19320 2654 19332
rect 2777 19329 2789 19332
rect 2823 19329 2835 19363
rect 2777 19323 2835 19329
rect 3234 19320 3240 19372
rect 3292 19320 3298 19372
rect 3326 19320 3332 19372
rect 3384 19360 3390 19372
rect 4706 19360 4712 19372
rect 3384 19332 4712 19360
rect 3384 19320 3390 19332
rect 2498 19252 2504 19304
rect 2556 19252 2562 19304
rect 2685 19295 2743 19301
rect 2685 19261 2697 19295
rect 2731 19261 2743 19295
rect 2685 19255 2743 19261
rect 2700 19224 2728 19255
rect 3418 19252 3424 19304
rect 3476 19252 3482 19304
rect 3513 19295 3571 19301
rect 3513 19261 3525 19295
rect 3559 19292 3571 19295
rect 3694 19292 3700 19304
rect 3559 19264 3700 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 3694 19252 3700 19264
rect 3752 19252 3758 19304
rect 3804 19301 3832 19332
rect 4706 19320 4712 19332
rect 4764 19360 4770 19372
rect 5092 19369 5120 19468
rect 5810 19456 5816 19468
rect 5868 19456 5874 19508
rect 5994 19456 6000 19508
rect 6052 19496 6058 19508
rect 6733 19499 6791 19505
rect 6733 19496 6745 19499
rect 6052 19468 6745 19496
rect 6052 19456 6058 19468
rect 6733 19465 6745 19468
rect 6779 19496 6791 19499
rect 7282 19496 7288 19508
rect 6779 19468 7288 19496
rect 6779 19465 6791 19468
rect 6733 19459 6791 19465
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 7653 19499 7711 19505
rect 7653 19465 7665 19499
rect 7699 19496 7711 19499
rect 7926 19496 7932 19508
rect 7699 19468 7932 19496
rect 7699 19465 7711 19468
rect 7653 19459 7711 19465
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 8570 19456 8576 19508
rect 8628 19456 8634 19508
rect 8662 19456 8668 19508
rect 8720 19456 8726 19508
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 9732 19468 10241 19496
rect 9732 19456 9738 19468
rect 10229 19465 10241 19468
rect 10275 19465 10287 19499
rect 10229 19459 10287 19465
rect 6273 19431 6331 19437
rect 6273 19428 6285 19431
rect 5460 19400 6285 19428
rect 5460 19369 5488 19400
rect 6273 19397 6285 19400
rect 6319 19397 6331 19431
rect 7374 19428 7380 19440
rect 6273 19391 6331 19397
rect 6748 19400 7380 19428
rect 5077 19363 5135 19369
rect 4764 19332 4936 19360
rect 4764 19320 4770 19332
rect 3789 19295 3847 19301
rect 3789 19261 3801 19295
rect 3835 19261 3847 19295
rect 3789 19255 3847 19261
rect 3970 19252 3976 19304
rect 4028 19292 4034 19304
rect 4065 19295 4123 19301
rect 4065 19292 4077 19295
rect 4028 19264 4077 19292
rect 4028 19252 4034 19264
rect 4065 19261 4077 19264
rect 4111 19261 4123 19295
rect 4801 19295 4859 19301
rect 4801 19292 4813 19295
rect 4065 19255 4123 19261
rect 4172 19264 4813 19292
rect 4172 19224 4200 19264
rect 4801 19261 4813 19264
rect 4847 19261 4859 19295
rect 4801 19255 4859 19261
rect 2700 19196 4200 19224
rect 4341 19227 4399 19233
rect 4341 19193 4353 19227
rect 4387 19193 4399 19227
rect 4341 19187 4399 19193
rect 3050 19156 3056 19168
rect 2424 19128 3056 19156
rect 943 19119 1001 19125
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3237 19159 3295 19165
rect 3237 19125 3249 19159
rect 3283 19156 3295 19159
rect 3326 19156 3332 19168
rect 3283 19128 3332 19156
rect 3283 19125 3295 19128
rect 3237 19119 3295 19125
rect 3326 19116 3332 19128
rect 3384 19116 3390 19168
rect 3510 19116 3516 19168
rect 3568 19156 3574 19168
rect 4157 19159 4215 19165
rect 4157 19156 4169 19159
rect 3568 19128 4169 19156
rect 3568 19116 3574 19128
rect 4157 19125 4169 19128
rect 4203 19125 4215 19159
rect 4356 19156 4384 19187
rect 4522 19184 4528 19236
rect 4580 19184 4586 19236
rect 4908 19224 4936 19332
rect 5077 19329 5089 19363
rect 5123 19329 5135 19363
rect 5077 19323 5135 19329
rect 5169 19363 5227 19369
rect 5169 19329 5181 19363
rect 5215 19360 5227 19363
rect 5445 19363 5503 19369
rect 5215 19332 5396 19360
rect 5215 19329 5227 19332
rect 5169 19323 5227 19329
rect 4982 19252 4988 19304
rect 5040 19252 5046 19304
rect 5261 19295 5319 19301
rect 5261 19261 5273 19295
rect 5307 19261 5319 19295
rect 5261 19255 5319 19261
rect 5276 19224 5304 19255
rect 4908 19196 5304 19224
rect 5368 19224 5396 19332
rect 5445 19329 5457 19363
rect 5491 19329 5503 19363
rect 5445 19323 5503 19329
rect 5534 19320 5540 19372
rect 5592 19360 5598 19372
rect 5813 19363 5871 19369
rect 5813 19360 5825 19363
rect 5592 19332 5825 19360
rect 5592 19320 5598 19332
rect 5813 19329 5825 19332
rect 5859 19329 5871 19363
rect 6748 19360 6776 19400
rect 7374 19388 7380 19400
rect 7432 19428 7438 19440
rect 8588 19428 8616 19456
rect 7432 19400 8616 19428
rect 7432 19388 7438 19400
rect 9122 19388 9128 19440
rect 9180 19388 9186 19440
rect 9692 19400 10548 19428
rect 7193 19363 7251 19369
rect 7193 19360 7205 19363
rect 5813 19323 5871 19329
rect 6104 19332 6776 19360
rect 6840 19332 7205 19360
rect 5626 19252 5632 19304
rect 5684 19252 5690 19304
rect 5721 19295 5779 19301
rect 5721 19261 5733 19295
rect 5767 19292 5779 19295
rect 5767 19264 5948 19292
rect 5767 19261 5779 19264
rect 5721 19255 5779 19261
rect 5813 19227 5871 19233
rect 5813 19224 5825 19227
rect 5368 19196 5825 19224
rect 5813 19193 5825 19196
rect 5859 19193 5871 19227
rect 5813 19187 5871 19193
rect 5074 19156 5080 19168
rect 4356 19128 5080 19156
rect 4157 19119 4215 19125
rect 5074 19116 5080 19128
rect 5132 19116 5138 19168
rect 5442 19116 5448 19168
rect 5500 19116 5506 19168
rect 5920 19156 5948 19264
rect 5994 19252 6000 19304
rect 6052 19252 6058 19304
rect 6104 19301 6132 19332
rect 6840 19304 6868 19332
rect 7193 19329 7205 19332
rect 7239 19360 7251 19363
rect 7742 19360 7748 19372
rect 7239 19332 7748 19360
rect 7239 19329 7251 19332
rect 7193 19323 7251 19329
rect 7742 19320 7748 19332
rect 7800 19320 7806 19372
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 9140 19360 9168 19388
rect 8628 19332 9260 19360
rect 8628 19320 8634 19332
rect 6089 19295 6147 19301
rect 6089 19261 6101 19295
rect 6135 19261 6147 19295
rect 6089 19255 6147 19261
rect 6454 19252 6460 19304
rect 6512 19252 6518 19304
rect 6549 19295 6607 19301
rect 6549 19261 6561 19295
rect 6595 19261 6607 19295
rect 6549 19255 6607 19261
rect 6270 19184 6276 19236
rect 6328 19224 6334 19236
rect 6564 19224 6592 19255
rect 6822 19252 6828 19304
rect 6880 19252 6886 19304
rect 6914 19252 6920 19304
rect 6972 19252 6978 19304
rect 7098 19252 7104 19304
rect 7156 19252 7162 19304
rect 7282 19252 7288 19304
rect 7340 19252 7346 19304
rect 7469 19295 7527 19301
rect 7469 19261 7481 19295
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 8021 19295 8079 19301
rect 8021 19261 8033 19295
rect 8067 19292 8079 19295
rect 8110 19292 8116 19304
rect 8067 19264 8116 19292
rect 8067 19261 8079 19264
rect 8021 19255 8079 19261
rect 6328 19196 6592 19224
rect 7484 19224 7512 19255
rect 8110 19252 8116 19264
rect 8168 19252 8174 19304
rect 8846 19252 8852 19304
rect 8904 19252 8910 19304
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19261 8999 19295
rect 8941 19255 8999 19261
rect 8478 19224 8484 19236
rect 7484 19196 8484 19224
rect 6328 19184 6334 19196
rect 7484 19156 7512 19196
rect 8478 19184 8484 19196
rect 8536 19184 8542 19236
rect 8956 19224 8984 19255
rect 9122 19252 9128 19304
rect 9180 19252 9186 19304
rect 9232 19301 9260 19332
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 9306 19252 9312 19304
rect 9364 19292 9370 19304
rect 9493 19295 9551 19301
rect 9493 19292 9505 19295
rect 9364 19264 9505 19292
rect 9364 19252 9370 19264
rect 9493 19261 9505 19264
rect 9539 19292 9551 19295
rect 9692 19292 9720 19400
rect 10321 19363 10379 19369
rect 10321 19360 10333 19363
rect 9968 19332 10333 19360
rect 9539 19264 9720 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 9766 19252 9772 19304
rect 9824 19252 9830 19304
rect 9968 19301 9996 19332
rect 10321 19329 10333 19332
rect 10367 19360 10379 19363
rect 10410 19360 10416 19372
rect 10367 19332 10416 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10410 19320 10416 19332
rect 10468 19320 10474 19372
rect 9965 19295 10023 19301
rect 9965 19261 9977 19295
rect 10011 19261 10023 19295
rect 10520 19292 10548 19400
rect 10597 19295 10655 19301
rect 10597 19292 10609 19295
rect 10520 19264 10609 19292
rect 9965 19255 10023 19261
rect 10597 19261 10609 19264
rect 10643 19261 10655 19295
rect 10597 19255 10655 19261
rect 8956 19196 10088 19224
rect 5920 19128 7512 19156
rect 7837 19159 7895 19165
rect 7837 19125 7849 19159
rect 7883 19156 7895 19159
rect 7926 19156 7932 19168
rect 7883 19128 7932 19156
rect 7883 19125 7895 19128
rect 7837 19119 7895 19125
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 8846 19116 8852 19168
rect 8904 19156 8910 19168
rect 9030 19156 9036 19168
rect 8904 19128 9036 19156
rect 8904 19116 8910 19128
rect 9030 19116 9036 19128
rect 9088 19156 9094 19168
rect 9309 19159 9367 19165
rect 9309 19156 9321 19159
rect 9088 19128 9321 19156
rect 9088 19116 9094 19128
rect 9309 19125 9321 19128
rect 9355 19125 9367 19159
rect 9309 19119 9367 19125
rect 9398 19116 9404 19168
rect 9456 19156 9462 19168
rect 9766 19156 9772 19168
rect 9456 19128 9772 19156
rect 9456 19116 9462 19128
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 10060 19165 10088 19196
rect 10045 19159 10103 19165
rect 10045 19125 10057 19159
rect 10091 19125 10103 19159
rect 10045 19119 10103 19125
rect 552 19066 11132 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 10722 19066
rect 10774 19014 10786 19066
rect 10838 19014 10850 19066
rect 10902 19014 10914 19066
rect 10966 19014 10978 19066
rect 11030 19014 11132 19066
rect 552 18992 11132 19014
rect 934 18912 940 18964
rect 992 18952 998 18964
rect 1486 18952 1492 18964
rect 992 18924 1492 18952
rect 992 18912 998 18924
rect 1486 18912 1492 18924
rect 1544 18912 1550 18964
rect 2130 18912 2136 18964
rect 2188 18952 2194 18964
rect 3237 18955 3295 18961
rect 3237 18952 3249 18955
rect 2188 18924 3249 18952
rect 2188 18912 2194 18924
rect 3237 18921 3249 18924
rect 3283 18921 3295 18955
rect 3237 18915 3295 18921
rect 4062 18912 4068 18964
rect 4120 18912 4126 18964
rect 4338 18912 4344 18964
rect 4396 18952 4402 18964
rect 5258 18952 5264 18964
rect 4396 18924 5264 18952
rect 4396 18912 4402 18924
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 5442 18912 5448 18964
rect 5500 18952 5506 18964
rect 6270 18952 6276 18964
rect 5500 18924 6276 18952
rect 5500 18912 5506 18924
rect 6270 18912 6276 18924
rect 6328 18912 6334 18964
rect 6914 18912 6920 18964
rect 6972 18912 6978 18964
rect 8389 18955 8447 18961
rect 8389 18921 8401 18955
rect 8435 18921 8447 18955
rect 8389 18915 8447 18921
rect 10321 18955 10379 18961
rect 10321 18921 10333 18955
rect 10367 18952 10379 18955
rect 10410 18952 10416 18964
rect 10367 18924 10416 18952
rect 10367 18921 10379 18924
rect 10321 18915 10379 18921
rect 566 18844 572 18896
rect 624 18884 630 18896
rect 845 18887 903 18893
rect 845 18884 857 18887
rect 624 18856 857 18884
rect 624 18844 630 18856
rect 845 18853 857 18856
rect 891 18853 903 18887
rect 2866 18884 2872 18896
rect 845 18847 903 18853
rect 1136 18856 2872 18884
rect 1136 18825 1164 18856
rect 2866 18844 2872 18856
rect 2924 18844 2930 18896
rect 4985 18887 5043 18893
rect 4985 18884 4997 18887
rect 3160 18856 4997 18884
rect 1029 18819 1087 18825
rect 1029 18785 1041 18819
rect 1075 18785 1087 18819
rect 1029 18779 1087 18785
rect 1121 18819 1179 18825
rect 1121 18785 1133 18819
rect 1167 18785 1179 18819
rect 1121 18779 1179 18785
rect 1213 18819 1271 18825
rect 1213 18785 1225 18819
rect 1259 18816 1271 18819
rect 1394 18816 1400 18828
rect 1259 18788 1400 18816
rect 1259 18785 1271 18788
rect 1213 18779 1271 18785
rect 1044 18748 1072 18779
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 1762 18776 1768 18828
rect 1820 18776 1826 18828
rect 2038 18776 2044 18828
rect 2096 18776 2102 18828
rect 2314 18776 2320 18828
rect 2372 18776 2378 18828
rect 2498 18776 2504 18828
rect 2556 18776 2562 18828
rect 2682 18776 2688 18828
rect 2740 18776 2746 18828
rect 3050 18776 3056 18828
rect 3108 18776 3114 18828
rect 2130 18748 2136 18760
rect 1044 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 2222 18708 2228 18760
rect 2280 18708 2286 18760
rect 2590 18708 2596 18760
rect 2648 18748 2654 18760
rect 2777 18751 2835 18757
rect 2777 18748 2789 18751
rect 2648 18720 2789 18748
rect 2648 18708 2654 18720
rect 2777 18717 2789 18720
rect 2823 18717 2835 18751
rect 2777 18711 2835 18717
rect 1578 18640 1584 18692
rect 1636 18680 1642 18692
rect 2608 18680 2636 18708
rect 3160 18680 3188 18856
rect 4985 18853 4997 18856
rect 5031 18853 5043 18887
rect 5718 18884 5724 18896
rect 4985 18847 5043 18853
rect 5506 18856 5724 18884
rect 3329 18819 3387 18825
rect 3329 18785 3341 18819
rect 3375 18816 3387 18819
rect 3510 18816 3516 18828
rect 3375 18788 3516 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 3510 18776 3516 18788
rect 3568 18776 3574 18828
rect 3697 18819 3755 18825
rect 3697 18785 3709 18819
rect 3743 18785 3755 18819
rect 3697 18779 3755 18785
rect 3712 18748 3740 18779
rect 3878 18776 3884 18828
rect 3936 18776 3942 18828
rect 4157 18819 4215 18825
rect 4157 18785 4169 18819
rect 4203 18785 4215 18819
rect 4157 18779 4215 18785
rect 4172 18748 4200 18779
rect 4338 18776 4344 18828
rect 4396 18776 4402 18828
rect 4893 18819 4951 18825
rect 4893 18816 4905 18819
rect 4804 18788 4905 18816
rect 3712 18720 4200 18748
rect 1636 18652 2636 18680
rect 2691 18652 3188 18680
rect 1636 18640 1642 18652
rect 842 18572 848 18624
rect 900 18572 906 18624
rect 2314 18572 2320 18624
rect 2372 18612 2378 18624
rect 2691 18612 2719 18652
rect 3418 18640 3424 18692
rect 3476 18680 3482 18692
rect 4172 18680 4200 18720
rect 4246 18708 4252 18760
rect 4304 18748 4310 18760
rect 4804 18748 4832 18788
rect 4893 18785 4905 18788
rect 4939 18785 4951 18819
rect 4893 18779 4951 18785
rect 5074 18776 5080 18828
rect 5132 18776 5138 18828
rect 5261 18819 5319 18825
rect 5261 18785 5273 18819
rect 5307 18816 5319 18819
rect 5506 18816 5534 18856
rect 5718 18844 5724 18856
rect 5776 18844 5782 18896
rect 5994 18844 6000 18896
rect 6052 18884 6058 18896
rect 6825 18887 6883 18893
rect 6052 18856 6776 18884
rect 6052 18844 6058 18856
rect 5307 18788 5534 18816
rect 5307 18785 5319 18788
rect 5261 18779 5319 18785
rect 6086 18776 6092 18828
rect 6144 18776 6150 18828
rect 6181 18819 6239 18825
rect 6181 18785 6193 18819
rect 6227 18785 6239 18819
rect 6181 18779 6239 18785
rect 4304 18720 4832 18748
rect 4985 18751 5043 18757
rect 4304 18708 4310 18720
rect 4985 18717 4997 18751
rect 5031 18748 5043 18751
rect 5092 18748 5120 18776
rect 5031 18720 5120 18748
rect 5031 18717 5043 18720
rect 4985 18711 5043 18717
rect 5902 18708 5908 18760
rect 5960 18708 5966 18760
rect 6196 18748 6224 18779
rect 6362 18776 6368 18828
rect 6420 18816 6426 18828
rect 6457 18819 6515 18825
rect 6457 18816 6469 18819
rect 6420 18788 6469 18816
rect 6420 18776 6426 18788
rect 6457 18785 6469 18788
rect 6503 18785 6515 18819
rect 6457 18779 6515 18785
rect 6546 18776 6552 18828
rect 6604 18816 6610 18828
rect 6641 18819 6699 18825
rect 6641 18816 6653 18819
rect 6604 18788 6653 18816
rect 6604 18776 6610 18788
rect 6641 18785 6653 18788
rect 6687 18785 6699 18819
rect 6748 18816 6776 18856
rect 6825 18853 6837 18887
rect 6871 18884 6883 18887
rect 7190 18884 7196 18896
rect 6871 18856 7196 18884
rect 6871 18853 6883 18856
rect 6825 18847 6883 18853
rect 7190 18844 7196 18856
rect 7248 18844 7254 18896
rect 7282 18844 7288 18896
rect 7340 18844 7346 18896
rect 7101 18819 7159 18825
rect 6748 18788 7063 18816
rect 6641 18779 6699 18785
rect 6914 18748 6920 18760
rect 6196 18720 6920 18748
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 7035 18748 7063 18788
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 7558 18816 7564 18828
rect 7147 18788 7564 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7800 18788 8033 18816
rect 7800 18776 7806 18788
rect 8021 18785 8033 18788
rect 8067 18816 8079 18819
rect 8404 18816 8432 18915
rect 10410 18912 10416 18924
rect 10468 18952 10474 18964
rect 10597 18955 10655 18961
rect 10597 18952 10609 18955
rect 10468 18924 10609 18952
rect 10468 18912 10474 18924
rect 10597 18921 10609 18924
rect 10643 18921 10655 18955
rect 10597 18915 10655 18921
rect 9401 18887 9459 18893
rect 9401 18853 9413 18887
rect 9447 18884 9459 18887
rect 9582 18884 9588 18896
rect 9447 18856 9588 18884
rect 9447 18853 9459 18856
rect 9401 18847 9459 18853
rect 9582 18844 9588 18856
rect 9640 18844 9646 18896
rect 10689 18887 10747 18893
rect 10689 18853 10701 18887
rect 10735 18884 10747 18887
rect 11238 18884 11244 18896
rect 10735 18856 11244 18884
rect 10735 18853 10747 18856
rect 10689 18847 10747 18853
rect 11238 18844 11244 18856
rect 11296 18844 11302 18896
rect 8662 18816 8668 18828
rect 8067 18788 8340 18816
rect 8404 18788 8668 18816
rect 8067 18785 8079 18788
rect 8021 18779 8079 18785
rect 7929 18751 7987 18757
rect 7929 18748 7941 18751
rect 7035 18720 7941 18748
rect 7929 18717 7941 18720
rect 7975 18748 7987 18751
rect 8110 18748 8116 18760
rect 7975 18720 8116 18748
rect 7975 18717 7987 18720
rect 7929 18711 7987 18717
rect 8110 18708 8116 18720
rect 8168 18708 8174 18760
rect 4525 18683 4583 18689
rect 3476 18652 4108 18680
rect 4172 18652 4289 18680
rect 3476 18640 3482 18652
rect 2372 18584 2719 18612
rect 2372 18572 2378 18584
rect 2866 18572 2872 18624
rect 2924 18572 2930 18624
rect 3050 18572 3056 18624
rect 3108 18612 3114 18624
rect 3602 18612 3608 18624
rect 3108 18584 3608 18612
rect 3108 18572 3114 18584
rect 3602 18572 3608 18584
rect 3660 18612 3666 18624
rect 3970 18612 3976 18624
rect 3660 18584 3976 18612
rect 3660 18572 3666 18584
rect 3970 18572 3976 18584
rect 4028 18572 4034 18624
rect 4080 18612 4108 18652
rect 4154 18612 4160 18624
rect 4080 18584 4160 18612
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 4261 18612 4289 18652
rect 4525 18649 4537 18683
rect 4571 18680 4583 18683
rect 4614 18680 4620 18692
rect 4571 18652 4620 18680
rect 4571 18649 4583 18652
rect 4525 18643 4583 18649
rect 4614 18640 4620 18652
rect 4672 18640 4678 18692
rect 4706 18640 4712 18692
rect 4764 18640 4770 18692
rect 5074 18640 5080 18692
rect 5132 18680 5138 18692
rect 5169 18683 5227 18689
rect 5169 18680 5181 18683
rect 5132 18652 5181 18680
rect 5132 18640 5138 18652
rect 5169 18649 5181 18652
rect 5215 18649 5227 18683
rect 6362 18680 6368 18692
rect 5169 18643 5227 18649
rect 5276 18652 6368 18680
rect 5276 18612 5304 18652
rect 6362 18640 6368 18652
rect 6420 18640 6426 18692
rect 6546 18640 6552 18692
rect 6604 18680 6610 18692
rect 7282 18680 7288 18692
rect 6604 18652 7288 18680
rect 6604 18640 6610 18652
rect 7282 18640 7288 18652
rect 7340 18640 7346 18692
rect 8312 18680 8340 18788
rect 8662 18776 8668 18788
rect 8720 18816 8726 18828
rect 8941 18819 8999 18825
rect 8941 18816 8953 18819
rect 8720 18788 8953 18816
rect 8720 18776 8726 18788
rect 8941 18785 8953 18788
rect 8987 18785 8999 18819
rect 9953 18819 10011 18825
rect 9953 18816 9965 18819
rect 8941 18779 8999 18785
rect 9048 18788 9965 18816
rect 9048 18760 9076 18788
rect 9953 18785 9965 18788
rect 9999 18785 10011 18819
rect 9953 18779 10011 18785
rect 10137 18819 10195 18825
rect 10137 18785 10149 18819
rect 10183 18785 10195 18819
rect 10137 18779 10195 18785
rect 10413 18819 10471 18825
rect 10413 18785 10425 18819
rect 10459 18816 10471 18819
rect 10502 18816 10508 18828
rect 10459 18788 10508 18816
rect 10459 18785 10471 18788
rect 10413 18779 10471 18785
rect 9030 18708 9036 18760
rect 9088 18708 9094 18760
rect 9306 18708 9312 18760
rect 9364 18708 9370 18760
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18748 9919 18751
rect 10152 18748 10180 18779
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 9907 18720 10180 18748
rect 9907 18717 9919 18720
rect 9861 18711 9919 18717
rect 9490 18680 9496 18692
rect 8312 18652 9496 18680
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 9674 18640 9680 18692
rect 9732 18640 9738 18692
rect 4261 18584 5304 18612
rect 5994 18572 6000 18624
rect 6052 18572 6058 18624
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 6730 18612 6736 18624
rect 6144 18584 6736 18612
rect 6144 18572 6150 18584
rect 6730 18572 6736 18584
rect 6788 18612 6794 18624
rect 7098 18612 7104 18624
rect 6788 18584 7104 18612
rect 6788 18572 6794 18584
rect 7098 18572 7104 18584
rect 7156 18572 7162 18624
rect 552 18522 11132 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 10062 18522
rect 10114 18470 10126 18522
rect 10178 18470 10190 18522
rect 10242 18470 10254 18522
rect 10306 18470 10318 18522
rect 10370 18470 11132 18522
rect 552 18448 11132 18470
rect 2038 18368 2044 18420
rect 2096 18368 2102 18420
rect 5166 18408 5172 18420
rect 3344 18380 5172 18408
rect 1397 18343 1455 18349
rect 1397 18309 1409 18343
rect 1443 18340 1455 18343
rect 3344 18340 3372 18380
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 5350 18368 5356 18420
rect 5408 18368 5414 18420
rect 5534 18368 5540 18420
rect 5592 18368 5598 18420
rect 5718 18368 5724 18420
rect 5776 18408 5782 18420
rect 5813 18411 5871 18417
rect 5813 18408 5825 18411
rect 5776 18380 5825 18408
rect 5776 18368 5782 18380
rect 5813 18377 5825 18380
rect 5859 18377 5871 18411
rect 6546 18408 6552 18420
rect 5813 18371 5871 18377
rect 6196 18380 6552 18408
rect 1443 18312 3372 18340
rect 1443 18309 1455 18312
rect 1397 18303 1455 18309
rect 3418 18300 3424 18352
rect 3476 18340 3482 18352
rect 3881 18343 3939 18349
rect 3881 18340 3893 18343
rect 3476 18312 3893 18340
rect 3476 18300 3482 18312
rect 3881 18309 3893 18312
rect 3927 18309 3939 18343
rect 3881 18303 3939 18309
rect 1118 18232 1124 18284
rect 1176 18272 1182 18284
rect 2133 18275 2191 18281
rect 2133 18272 2145 18275
rect 1176 18244 2145 18272
rect 1176 18232 1182 18244
rect 2133 18241 2145 18244
rect 2179 18241 2191 18275
rect 2133 18235 2191 18241
rect 2314 18232 2320 18284
rect 2372 18232 2378 18284
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18272 2467 18275
rect 3789 18275 3847 18281
rect 3789 18272 3801 18275
rect 2455 18244 3801 18272
rect 2455 18241 2467 18244
rect 2409 18235 2467 18241
rect 3789 18241 3801 18244
rect 3835 18241 3847 18275
rect 3789 18235 3847 18241
rect 1213 18207 1271 18213
rect 1213 18173 1225 18207
rect 1259 18204 1271 18207
rect 1489 18207 1547 18213
rect 1259 18176 1440 18204
rect 1259 18173 1271 18176
rect 1213 18167 1271 18173
rect 1412 18148 1440 18176
rect 1489 18173 1501 18207
rect 1535 18204 1547 18207
rect 1578 18204 1584 18216
rect 1535 18176 1584 18204
rect 1535 18173 1547 18176
rect 1489 18167 1547 18173
rect 1578 18164 1584 18176
rect 1636 18164 1642 18216
rect 1670 18164 1676 18216
rect 1728 18164 1734 18216
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18204 1915 18207
rect 2866 18204 2872 18216
rect 1903 18176 2872 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 1394 18096 1400 18148
rect 1452 18136 1458 18148
rect 1872 18136 1900 18167
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 3234 18164 3240 18216
rect 3292 18164 3298 18216
rect 3326 18164 3332 18216
rect 3384 18164 3390 18216
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18173 3571 18207
rect 3513 18167 3571 18173
rect 3605 18207 3663 18213
rect 3605 18173 3617 18207
rect 3651 18204 3663 18207
rect 3896 18204 3924 18303
rect 3970 18300 3976 18352
rect 4028 18340 4034 18352
rect 5368 18340 5396 18368
rect 5445 18343 5503 18349
rect 5445 18340 5457 18343
rect 4028 18312 4660 18340
rect 5368 18312 5457 18340
rect 4028 18300 4034 18312
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 4338 18272 4344 18284
rect 4212 18244 4344 18272
rect 4212 18232 4218 18244
rect 4338 18232 4344 18244
rect 4396 18232 4402 18284
rect 4522 18232 4528 18284
rect 4580 18232 4586 18284
rect 4632 18272 4660 18312
rect 5445 18309 5457 18312
rect 5491 18309 5503 18343
rect 5994 18340 6000 18352
rect 5445 18303 5503 18309
rect 5644 18312 6000 18340
rect 5537 18275 5595 18281
rect 4632 18244 5488 18272
rect 3651 18176 3924 18204
rect 3651 18173 3663 18176
rect 3605 18167 3663 18173
rect 1452 18108 1900 18136
rect 2777 18139 2835 18145
rect 1452 18096 1458 18108
rect 2777 18105 2789 18139
rect 2823 18136 2835 18139
rect 2958 18136 2964 18148
rect 2823 18108 2964 18136
rect 2823 18105 2835 18108
rect 2777 18099 2835 18105
rect 2958 18096 2964 18108
rect 3016 18096 3022 18148
rect 3528 18136 3556 18167
rect 3970 18164 3976 18216
rect 4028 18204 4034 18216
rect 4065 18207 4123 18213
rect 4065 18204 4077 18207
rect 4028 18176 4077 18204
rect 4028 18164 4034 18176
rect 4065 18173 4077 18176
rect 4111 18173 4123 18207
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 4065 18167 4123 18173
rect 4172 18176 4261 18204
rect 3786 18136 3792 18148
rect 3528 18108 3792 18136
rect 3786 18096 3792 18108
rect 3844 18096 3850 18148
rect 1029 18071 1087 18077
rect 1029 18037 1041 18071
rect 1075 18068 1087 18071
rect 1946 18068 1952 18080
rect 1075 18040 1952 18068
rect 1075 18037 1087 18040
rect 1029 18031 1087 18037
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 3694 18028 3700 18080
rect 3752 18068 3758 18080
rect 4172 18068 4200 18176
rect 4249 18173 4261 18176
rect 4295 18173 4307 18207
rect 4249 18167 4307 18173
rect 4433 18207 4491 18213
rect 4433 18173 4445 18207
rect 4479 18204 4491 18207
rect 4524 18204 4552 18232
rect 4479 18176 4552 18204
rect 4893 18207 4951 18213
rect 4617 18185 4675 18191
rect 4479 18173 4491 18176
rect 4433 18167 4491 18173
rect 4617 18151 4629 18185
rect 4663 18151 4675 18185
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 5074 18204 5080 18216
rect 4939 18176 5080 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5166 18164 5172 18216
rect 5224 18204 5230 18216
rect 5353 18207 5411 18213
rect 5353 18204 5365 18207
rect 5224 18176 5365 18204
rect 5224 18164 5230 18176
rect 5353 18173 5365 18176
rect 5399 18173 5411 18207
rect 5353 18167 5411 18173
rect 4617 18148 4675 18151
rect 4614 18096 4620 18148
rect 4672 18096 4678 18148
rect 4709 18139 4767 18145
rect 4709 18105 4721 18139
rect 4755 18105 4767 18139
rect 4709 18099 4767 18105
rect 3752 18040 4200 18068
rect 3752 18028 3758 18040
rect 4430 18028 4436 18080
rect 4488 18068 4494 18080
rect 4724 18068 4752 18099
rect 4488 18040 4752 18068
rect 4488 18028 4494 18040
rect 5074 18028 5080 18080
rect 5132 18028 5138 18080
rect 5460 18068 5488 18244
rect 5537 18241 5549 18275
rect 5583 18272 5595 18275
rect 5644 18272 5672 18312
rect 5994 18300 6000 18312
rect 6052 18300 6058 18352
rect 5583 18244 5672 18272
rect 5583 18241 5595 18244
rect 5537 18235 5595 18241
rect 5718 18232 5724 18284
rect 5776 18232 5782 18284
rect 5810 18232 5816 18284
rect 5868 18272 5874 18284
rect 5868 18244 6040 18272
rect 5868 18232 5874 18244
rect 6012 18214 6040 18244
rect 6012 18207 6132 18214
rect 6196 18213 6224 18380
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 6822 18300 6828 18352
rect 6880 18340 6886 18352
rect 7558 18340 7564 18352
rect 6880 18312 7564 18340
rect 6880 18300 6886 18312
rect 7558 18300 7564 18312
rect 7616 18300 7622 18352
rect 7650 18300 7656 18352
rect 7708 18340 7714 18352
rect 7708 18312 7880 18340
rect 7708 18300 7714 18312
rect 6546 18232 6552 18284
rect 6604 18272 6610 18284
rect 6604 18244 7696 18272
rect 6604 18232 6610 18244
rect 7668 18216 7696 18244
rect 7742 18232 7748 18284
rect 7800 18232 7806 18284
rect 6012 18186 6081 18207
rect 6069 18173 6081 18186
rect 6115 18176 6132 18207
rect 6181 18207 6239 18213
rect 6115 18173 6127 18176
rect 6069 18167 6127 18173
rect 6181 18173 6193 18207
rect 6227 18173 6239 18207
rect 6181 18167 6239 18173
rect 6273 18207 6331 18213
rect 6273 18173 6285 18207
rect 6319 18173 6331 18207
rect 6273 18167 6331 18173
rect 6457 18207 6515 18213
rect 6457 18173 6469 18207
rect 6503 18173 6515 18207
rect 6457 18167 6515 18173
rect 6288 18136 6316 18167
rect 6362 18136 6368 18148
rect 6288 18108 6368 18136
rect 6362 18096 6368 18108
rect 6420 18096 6426 18148
rect 6472 18068 6500 18167
rect 7282 18164 7288 18216
rect 7340 18164 7346 18216
rect 7469 18207 7527 18213
rect 7469 18173 7481 18207
rect 7515 18173 7527 18207
rect 7469 18167 7527 18173
rect 7561 18207 7619 18213
rect 7561 18173 7573 18207
rect 7607 18173 7619 18207
rect 7561 18167 7619 18173
rect 6546 18096 6552 18148
rect 6604 18136 6610 18148
rect 6641 18139 6699 18145
rect 6641 18136 6653 18139
rect 6604 18108 6653 18136
rect 6604 18096 6610 18108
rect 6641 18105 6653 18108
rect 6687 18105 6699 18139
rect 6641 18099 6699 18105
rect 5460 18040 6500 18068
rect 6914 18028 6920 18080
rect 6972 18028 6978 18080
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 7101 18071 7159 18077
rect 7101 18068 7113 18071
rect 7064 18040 7113 18068
rect 7064 18028 7070 18040
rect 7101 18037 7113 18040
rect 7147 18037 7159 18071
rect 7101 18031 7159 18037
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 7484 18068 7512 18167
rect 7576 18136 7604 18167
rect 7650 18164 7656 18216
rect 7708 18164 7714 18216
rect 7852 18213 7880 18312
rect 9030 18300 9036 18352
rect 9088 18300 9094 18352
rect 9582 18340 9588 18352
rect 9324 18312 9588 18340
rect 8018 18232 8024 18284
rect 8076 18232 8082 18284
rect 8662 18232 8668 18284
rect 8720 18232 8726 18284
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 8036 18136 8064 18232
rect 8386 18164 8392 18216
rect 8444 18204 8450 18216
rect 9324 18213 9352 18312
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 9398 18232 9404 18284
rect 9456 18272 9462 18284
rect 10321 18275 10379 18281
rect 10321 18272 10333 18275
rect 9456 18244 10333 18272
rect 9456 18232 9462 18244
rect 10321 18241 10333 18244
rect 10367 18272 10379 18275
rect 10502 18272 10508 18284
rect 10367 18244 10508 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 10502 18232 10508 18244
rect 10560 18232 10566 18284
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 8444 18176 9321 18204
rect 8444 18164 8450 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 9493 18207 9551 18213
rect 9493 18173 9505 18207
rect 9539 18204 9551 18207
rect 9674 18204 9680 18216
rect 9539 18176 9680 18204
rect 9539 18173 9551 18176
rect 9493 18167 9551 18173
rect 7576 18108 8064 18136
rect 8478 18096 8484 18148
rect 8536 18136 8542 18148
rect 9508 18136 9536 18167
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 8536 18108 9536 18136
rect 8536 18096 8542 18108
rect 7340 18040 7512 18068
rect 9125 18071 9183 18077
rect 7340 18028 7346 18040
rect 9125 18037 9137 18071
rect 9171 18068 9183 18071
rect 9214 18068 9220 18080
rect 9171 18040 9220 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 552 17978 11132 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 10722 17978
rect 10774 17926 10786 17978
rect 10838 17926 10850 17978
rect 10902 17926 10914 17978
rect 10966 17926 10978 17978
rect 11030 17926 11132 17978
rect 552 17904 11132 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 3697 17867 3755 17873
rect 3697 17864 3709 17867
rect 1728 17836 3709 17864
rect 1728 17824 1734 17836
rect 3697 17833 3709 17836
rect 3743 17833 3755 17867
rect 3697 17827 3755 17833
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4338 17864 4344 17876
rect 4120 17836 4344 17864
rect 4120 17824 4126 17836
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 5074 17824 5080 17876
rect 5132 17824 5138 17876
rect 5813 17867 5871 17873
rect 5813 17833 5825 17867
rect 5859 17864 5871 17867
rect 5902 17864 5908 17876
rect 5859 17836 5908 17864
rect 5859 17833 5871 17836
rect 5813 17827 5871 17833
rect 5902 17824 5908 17836
rect 5960 17824 5966 17876
rect 6730 17824 6736 17876
rect 6788 17824 6794 17876
rect 6932 17836 7696 17864
rect 842 17756 848 17808
rect 900 17796 906 17808
rect 4522 17796 4528 17808
rect 900 17768 2636 17796
rect 900 17756 906 17768
rect 1302 17688 1308 17740
rect 1360 17688 1366 17740
rect 1872 17737 1900 17768
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17697 1639 17731
rect 1581 17691 1639 17697
rect 1857 17731 1915 17737
rect 1857 17697 1869 17731
rect 1903 17697 1915 17731
rect 1857 17691 1915 17697
rect 382 17620 388 17672
rect 440 17660 446 17672
rect 842 17660 848 17672
rect 440 17632 848 17660
rect 440 17620 446 17632
rect 842 17620 848 17632
rect 900 17620 906 17672
rect 1118 17484 1124 17536
rect 1176 17484 1182 17536
rect 1320 17524 1348 17688
rect 1596 17660 1624 17691
rect 2130 17688 2136 17740
rect 2188 17688 2194 17740
rect 2608 17737 2636 17768
rect 2700 17768 3096 17796
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17728 2375 17731
rect 2593 17731 2651 17737
rect 2363 17700 2544 17728
rect 2363 17697 2375 17700
rect 2317 17691 2375 17697
rect 2516 17672 2544 17700
rect 2593 17697 2605 17731
rect 2639 17697 2651 17731
rect 2593 17691 2651 17697
rect 2222 17660 2228 17672
rect 1596 17632 2228 17660
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 2498 17620 2504 17672
rect 2556 17660 2562 17672
rect 2700 17660 2728 17768
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 3068 17737 3096 17768
rect 3620 17768 4528 17796
rect 2869 17731 2927 17737
rect 2869 17728 2881 17731
rect 2832 17700 2881 17728
rect 2832 17688 2838 17700
rect 2869 17697 2881 17700
rect 2915 17697 2927 17731
rect 2869 17691 2927 17697
rect 3053 17731 3111 17737
rect 3053 17697 3065 17731
rect 3099 17728 3111 17731
rect 3329 17731 3387 17737
rect 3329 17728 3341 17731
rect 3099 17700 3341 17728
rect 3099 17697 3111 17700
rect 3053 17691 3111 17697
rect 3329 17697 3341 17700
rect 3375 17697 3387 17731
rect 3329 17691 3387 17697
rect 3510 17688 3516 17740
rect 3568 17688 3574 17740
rect 3620 17737 3648 17768
rect 4522 17756 4528 17768
rect 4580 17756 4586 17808
rect 5092 17796 5120 17824
rect 6546 17796 6552 17808
rect 5000 17768 5120 17796
rect 6012 17768 6552 17796
rect 3605 17731 3663 17737
rect 3605 17697 3617 17731
rect 3651 17697 3663 17731
rect 3605 17691 3663 17697
rect 3878 17688 3884 17740
rect 3936 17688 3942 17740
rect 4246 17688 4252 17740
rect 4304 17728 4310 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 4304 17700 4445 17728
rect 4304 17688 4310 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4614 17728 4620 17740
rect 4433 17691 4491 17697
rect 4540 17700 4620 17728
rect 2556 17632 2728 17660
rect 3528 17660 3556 17688
rect 3896 17660 3924 17688
rect 3528 17632 3924 17660
rect 2556 17620 2562 17632
rect 4062 17620 4068 17672
rect 4120 17620 4126 17672
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17660 4215 17663
rect 4203 17632 4476 17660
rect 4203 17629 4215 17632
rect 4157 17623 4215 17629
rect 4448 17604 4476 17632
rect 1489 17595 1547 17601
rect 1489 17561 1501 17595
rect 1535 17592 1547 17595
rect 1673 17595 1731 17601
rect 1673 17592 1685 17595
rect 1535 17564 1685 17592
rect 1535 17561 1547 17564
rect 1489 17555 1547 17561
rect 1673 17561 1685 17564
rect 1719 17561 1731 17595
rect 1673 17555 1731 17561
rect 1854 17552 1860 17604
rect 1912 17592 1918 17604
rect 2682 17592 2688 17604
rect 1912 17564 2688 17592
rect 1912 17552 1918 17564
rect 2682 17552 2688 17564
rect 2740 17552 2746 17604
rect 2866 17552 2872 17604
rect 2924 17592 2930 17604
rect 3050 17592 3056 17604
rect 2924 17564 3056 17592
rect 2924 17552 2930 17564
rect 3050 17552 3056 17564
rect 3108 17552 3114 17604
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 4249 17595 4307 17601
rect 4249 17592 4261 17595
rect 3568 17564 4261 17592
rect 3568 17552 3574 17564
rect 4249 17561 4261 17564
rect 4295 17561 4307 17595
rect 4249 17555 4307 17561
rect 4430 17552 4436 17604
rect 4488 17552 4494 17604
rect 4540 17592 4568 17700
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 4798 17688 4804 17740
rect 4856 17688 4862 17740
rect 5000 17737 5028 17768
rect 4985 17731 5043 17737
rect 4985 17697 4997 17731
rect 5031 17697 5043 17731
rect 4985 17691 5043 17697
rect 5074 17688 5080 17740
rect 5132 17688 5138 17740
rect 5258 17688 5264 17740
rect 5316 17688 5322 17740
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17728 5411 17731
rect 5442 17728 5448 17740
rect 5399 17700 5448 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 5626 17688 5632 17740
rect 5684 17688 5690 17740
rect 5902 17688 5908 17740
rect 5960 17728 5966 17740
rect 6012 17737 6040 17768
rect 6546 17756 6552 17768
rect 6604 17756 6610 17808
rect 6748 17796 6776 17824
rect 6656 17768 6776 17796
rect 5997 17731 6055 17737
rect 5997 17728 6009 17731
rect 5960 17700 6009 17728
rect 5960 17688 5966 17700
rect 5997 17697 6009 17700
rect 6043 17697 6055 17731
rect 5997 17691 6055 17697
rect 6089 17731 6147 17737
rect 6089 17697 6101 17731
rect 6135 17728 6147 17731
rect 6270 17728 6276 17740
rect 6135 17700 6276 17728
rect 6135 17697 6147 17700
rect 6089 17691 6147 17697
rect 6270 17688 6276 17700
rect 6328 17688 6334 17740
rect 6365 17731 6423 17737
rect 6365 17730 6377 17731
rect 6362 17697 6377 17730
rect 6411 17697 6423 17731
rect 6362 17691 6423 17697
rect 4706 17620 4712 17672
rect 4764 17620 4770 17672
rect 6362 17660 6390 17691
rect 6454 17688 6460 17740
rect 6512 17688 6518 17740
rect 6656 17737 6684 17768
rect 6641 17731 6699 17737
rect 6641 17697 6653 17731
rect 6687 17697 6699 17731
rect 6932 17728 6960 17836
rect 7374 17796 7380 17808
rect 7024 17768 7380 17796
rect 7024 17737 7052 17768
rect 7374 17756 7380 17768
rect 7432 17796 7438 17808
rect 7668 17796 7696 17836
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 8021 17867 8079 17873
rect 8021 17864 8033 17867
rect 7800 17836 8033 17864
rect 7800 17824 7806 17836
rect 8021 17833 8033 17836
rect 8067 17833 8079 17867
rect 8662 17864 8668 17876
rect 8021 17827 8079 17833
rect 8128 17836 8668 17864
rect 7432 17768 7604 17796
rect 7668 17768 7880 17796
rect 7432 17756 7438 17768
rect 6641 17691 6699 17697
rect 6748 17700 6960 17728
rect 7009 17731 7067 17737
rect 6546 17660 6552 17672
rect 6362 17632 6552 17660
rect 6546 17620 6552 17632
rect 6604 17660 6610 17672
rect 6748 17669 6776 17700
rect 7009 17697 7021 17731
rect 7055 17697 7067 17731
rect 7009 17691 7067 17697
rect 7190 17688 7196 17740
rect 7248 17688 7254 17740
rect 7576 17737 7604 17768
rect 7285 17731 7343 17737
rect 7285 17697 7297 17731
rect 7331 17697 7343 17731
rect 7285 17691 7343 17697
rect 7469 17731 7527 17737
rect 7469 17697 7481 17731
rect 7515 17697 7527 17731
rect 7469 17691 7527 17697
rect 7564 17731 7622 17737
rect 7564 17697 7576 17731
rect 7610 17697 7622 17731
rect 7564 17691 7622 17697
rect 6733 17663 6791 17669
rect 6733 17660 6745 17663
rect 6604 17632 6745 17660
rect 6604 17620 6610 17632
rect 6733 17629 6745 17632
rect 6779 17629 6791 17663
rect 6733 17623 6791 17629
rect 6822 17620 6828 17672
rect 6880 17620 6886 17672
rect 7300 17604 7328 17691
rect 5537 17595 5595 17601
rect 4540 17564 5120 17592
rect 1578 17524 1584 17536
rect 1320 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 2038 17484 2044 17536
rect 2096 17524 2102 17536
rect 2409 17527 2467 17533
rect 2409 17524 2421 17527
rect 2096 17496 2421 17524
rect 2096 17484 2102 17496
rect 2409 17493 2421 17496
rect 2455 17493 2467 17527
rect 2409 17487 2467 17493
rect 2498 17484 2504 17536
rect 2556 17524 2562 17536
rect 3145 17527 3203 17533
rect 3145 17524 3157 17527
rect 2556 17496 3157 17524
rect 2556 17484 2562 17496
rect 3145 17493 3157 17496
rect 3191 17493 3203 17527
rect 3145 17487 3203 17493
rect 3418 17484 3424 17536
rect 3476 17524 3482 17536
rect 3694 17524 3700 17536
rect 3476 17496 3700 17524
rect 3476 17484 3482 17496
rect 3694 17484 3700 17496
rect 3752 17524 3758 17536
rect 4798 17524 4804 17536
rect 3752 17496 4804 17524
rect 3752 17484 3758 17496
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 5092 17524 5120 17564
rect 5537 17561 5549 17595
rect 5583 17592 5595 17595
rect 5583 17564 5856 17592
rect 5583 17561 5595 17564
rect 5537 17555 5595 17561
rect 5552 17524 5580 17555
rect 5092 17496 5580 17524
rect 5828 17524 5856 17564
rect 6270 17552 6276 17604
rect 6328 17592 6334 17604
rect 6328 17564 6960 17592
rect 6328 17552 6334 17564
rect 6822 17524 6828 17536
rect 5828 17496 6828 17524
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 6932 17524 6960 17564
rect 7282 17552 7288 17604
rect 7340 17552 7346 17604
rect 7472 17524 7500 17691
rect 7650 17688 7656 17740
rect 7708 17688 7714 17740
rect 7852 17737 7880 17768
rect 7837 17731 7895 17737
rect 7837 17697 7849 17731
rect 7883 17697 7895 17731
rect 7837 17691 7895 17697
rect 8018 17688 8024 17740
rect 8076 17728 8082 17740
rect 8128 17728 8156 17836
rect 8662 17824 8668 17836
rect 8720 17824 8726 17876
rect 9674 17864 9680 17876
rect 9048 17836 9680 17864
rect 8386 17756 8392 17808
rect 8444 17796 8450 17808
rect 8570 17796 8576 17808
rect 8444 17768 8576 17796
rect 8444 17756 8450 17768
rect 8570 17756 8576 17768
rect 8628 17756 8634 17808
rect 8680 17796 8708 17824
rect 9048 17805 9076 17836
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 9033 17799 9091 17805
rect 8680 17768 8800 17796
rect 8076 17700 8156 17728
rect 8297 17731 8355 17737
rect 8076 17688 8082 17700
rect 8297 17697 8309 17731
rect 8343 17697 8355 17731
rect 8297 17691 8355 17697
rect 8312 17660 8340 17691
rect 8478 17688 8484 17740
rect 8536 17688 8542 17740
rect 8662 17688 8668 17740
rect 8720 17688 8726 17740
rect 8772 17737 8800 17768
rect 9033 17765 9045 17799
rect 9079 17765 9091 17799
rect 9033 17759 9091 17765
rect 8757 17731 8815 17737
rect 8757 17697 8769 17731
rect 8803 17697 8815 17731
rect 8757 17691 8815 17697
rect 9398 17688 9404 17740
rect 9456 17688 9462 17740
rect 9858 17688 9864 17740
rect 9916 17728 9922 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9916 17700 10057 17728
rect 9916 17688 9922 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 9122 17660 9128 17672
rect 8312 17632 9128 17660
rect 9122 17620 9128 17632
rect 9180 17660 9186 17672
rect 9585 17663 9643 17669
rect 9180 17632 9444 17660
rect 9180 17620 9186 17632
rect 9416 17604 9444 17632
rect 9585 17629 9597 17663
rect 9631 17660 9643 17663
rect 9674 17660 9680 17672
rect 9631 17632 9680 17660
rect 9631 17629 9643 17632
rect 9585 17623 9643 17629
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 8294 17552 8300 17604
rect 8352 17592 8358 17604
rect 9030 17592 9036 17604
rect 8352 17564 9036 17592
rect 8352 17552 8358 17564
rect 9030 17552 9036 17564
rect 9088 17552 9094 17604
rect 9398 17552 9404 17604
rect 9456 17552 9462 17604
rect 9490 17552 9496 17604
rect 9548 17592 9554 17604
rect 9861 17595 9919 17601
rect 9861 17592 9873 17595
rect 9548 17564 9873 17592
rect 9548 17552 9554 17564
rect 9861 17561 9873 17564
rect 9907 17561 9919 17595
rect 9861 17555 9919 17561
rect 6932 17496 7500 17524
rect 7558 17484 7564 17536
rect 7616 17524 7622 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7616 17496 8125 17524
rect 7616 17484 7622 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8113 17487 8171 17493
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 9125 17527 9183 17533
rect 9125 17524 9137 17527
rect 8444 17496 9137 17524
rect 8444 17484 8450 17496
rect 9125 17493 9137 17496
rect 9171 17493 9183 17527
rect 9125 17487 9183 17493
rect 552 17434 11132 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 10062 17434
rect 10114 17382 10126 17434
rect 10178 17382 10190 17434
rect 10242 17382 10254 17434
rect 10306 17382 10318 17434
rect 10370 17382 11132 17434
rect 552 17360 11132 17382
rect 2130 17280 2136 17332
rect 2188 17320 2194 17332
rect 2317 17323 2375 17329
rect 2317 17320 2329 17323
rect 2188 17292 2329 17320
rect 2188 17280 2194 17292
rect 2317 17289 2329 17292
rect 2363 17289 2375 17323
rect 3605 17323 3663 17329
rect 3605 17320 3617 17323
rect 2317 17283 2375 17289
rect 2424 17292 3617 17320
rect 106 17212 112 17264
rect 164 17252 170 17264
rect 2424 17252 2452 17292
rect 3605 17289 3617 17292
rect 3651 17289 3663 17323
rect 3605 17283 3663 17289
rect 3804 17292 4016 17320
rect 3050 17252 3056 17264
rect 164 17224 2452 17252
rect 2608 17224 3056 17252
rect 164 17212 170 17224
rect 1762 17144 1768 17196
rect 1820 17144 1826 17196
rect 1946 17076 1952 17128
rect 2004 17116 2010 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 2004 17088 2053 17116
rect 2004 17076 2010 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 2222 17076 2228 17128
rect 2280 17076 2286 17128
rect 2608 17125 2636 17224
rect 3050 17212 3056 17224
rect 3108 17212 3114 17264
rect 3142 17212 3148 17264
rect 3200 17252 3206 17264
rect 3329 17255 3387 17261
rect 3329 17252 3341 17255
rect 3200 17224 3341 17252
rect 3200 17212 3206 17224
rect 3329 17221 3341 17224
rect 3375 17221 3387 17255
rect 3329 17215 3387 17221
rect 3418 17184 3424 17196
rect 2700 17156 3424 17184
rect 2700 17125 2728 17156
rect 3418 17144 3424 17156
rect 3476 17144 3482 17196
rect 3513 17187 3571 17193
rect 3513 17153 3525 17187
rect 3559 17184 3571 17187
rect 3804 17184 3832 17292
rect 3988 17252 4016 17292
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 4120 17292 5641 17320
rect 4120 17280 4126 17292
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 5629 17283 5687 17289
rect 6822 17280 6828 17332
rect 6880 17320 6886 17332
rect 7650 17320 7656 17332
rect 6880 17292 7656 17320
rect 6880 17280 6886 17292
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 10410 17320 10416 17332
rect 8864 17292 10416 17320
rect 5074 17252 5080 17264
rect 3988 17224 5080 17252
rect 5074 17212 5080 17224
rect 5132 17212 5138 17264
rect 5810 17212 5816 17264
rect 5868 17252 5874 17264
rect 5868 17224 6868 17252
rect 5868 17212 5874 17224
rect 6840 17196 6868 17224
rect 3559 17156 3832 17184
rect 3559 17153 3571 17156
rect 3513 17147 3571 17153
rect 3970 17144 3976 17196
rect 4028 17184 4034 17196
rect 4028 17156 5580 17184
rect 4028 17144 4034 17156
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17085 2651 17119
rect 2593 17079 2651 17085
rect 2685 17119 2743 17125
rect 2685 17085 2697 17119
rect 2731 17085 2743 17119
rect 2685 17079 2743 17085
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17085 2835 17119
rect 2777 17079 2835 17085
rect 658 17008 664 17060
rect 716 17048 722 17060
rect 1213 17051 1271 17057
rect 1213 17048 1225 17051
rect 716 17020 1225 17048
rect 716 17008 722 17020
rect 1213 17017 1225 17020
rect 1259 17017 1271 17051
rect 1213 17011 1271 17017
rect 2590 16940 2596 16992
rect 2648 16980 2654 16992
rect 2792 16980 2820 17079
rect 2958 17076 2964 17128
rect 3016 17076 3022 17128
rect 3237 17119 3295 17125
rect 3237 17085 3249 17119
rect 3283 17085 3295 17119
rect 3237 17079 3295 17085
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17085 3847 17119
rect 3789 17079 3847 17085
rect 3252 17048 3280 17079
rect 3694 17048 3700 17060
rect 3252 17020 3700 17048
rect 3694 17008 3700 17020
rect 3752 17008 3758 17060
rect 3804 17048 3832 17079
rect 3878 17076 3884 17128
rect 3936 17076 3942 17128
rect 4062 17076 4068 17128
rect 4120 17076 4126 17128
rect 4172 17125 4200 17156
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17085 4215 17119
rect 4157 17079 4215 17085
rect 4338 17076 4344 17128
rect 4396 17116 4402 17128
rect 4433 17119 4491 17125
rect 4433 17116 4445 17119
rect 4396 17088 4445 17116
rect 4396 17076 4402 17088
rect 4433 17085 4445 17088
rect 4479 17085 4491 17119
rect 4433 17079 4491 17085
rect 4614 17076 4620 17128
rect 4672 17076 4678 17128
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17085 4767 17119
rect 4709 17079 4767 17085
rect 3804 17020 4292 17048
rect 2648 16952 2820 16980
rect 3513 16983 3571 16989
rect 2648 16940 2654 16952
rect 3513 16949 3525 16983
rect 3559 16980 3571 16983
rect 3878 16980 3884 16992
rect 3559 16952 3884 16980
rect 3559 16949 3571 16952
rect 3513 16943 3571 16949
rect 3878 16940 3884 16952
rect 3936 16940 3942 16992
rect 4264 16989 4292 17020
rect 4522 17008 4528 17060
rect 4580 17048 4586 17060
rect 4724 17048 4752 17079
rect 4798 17076 4804 17128
rect 4856 17076 4862 17128
rect 4985 17119 5043 17125
rect 4985 17085 4997 17119
rect 5031 17116 5043 17119
rect 5445 17119 5503 17125
rect 5445 17116 5457 17119
rect 5031 17088 5457 17116
rect 5031 17085 5043 17088
rect 4985 17079 5043 17085
rect 5445 17085 5457 17088
rect 5491 17085 5503 17119
rect 5445 17079 5503 17085
rect 4580 17020 4752 17048
rect 4580 17008 4586 17020
rect 5074 17008 5080 17060
rect 5132 17008 5138 17060
rect 5261 17051 5319 17057
rect 5261 17017 5273 17051
rect 5307 17048 5319 17051
rect 5307 17020 5488 17048
rect 5307 17017 5319 17020
rect 5261 17011 5319 17017
rect 5460 16992 5488 17020
rect 4249 16983 4307 16989
rect 4249 16949 4261 16983
rect 4295 16980 4307 16983
rect 5166 16980 5172 16992
rect 4295 16952 5172 16980
rect 4295 16949 4307 16952
rect 4249 16943 4307 16949
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 5442 16940 5448 16992
rect 5500 16940 5506 16992
rect 5552 16980 5580 17156
rect 5718 17144 5724 17196
rect 5776 17144 5782 17196
rect 5994 17184 6000 17196
rect 5828 17156 6000 17184
rect 5736 17048 5764 17144
rect 5828 17125 5856 17156
rect 5994 17144 6000 17156
rect 6052 17144 6058 17196
rect 6822 17144 6828 17196
rect 6880 17144 6886 17196
rect 7009 17187 7067 17193
rect 7009 17153 7021 17187
rect 7055 17184 7067 17187
rect 7190 17184 7196 17196
rect 7055 17156 7196 17184
rect 7055 17153 7067 17156
rect 7009 17147 7067 17153
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 8018 17184 8024 17196
rect 7392 17156 8024 17184
rect 7392 17128 7420 17156
rect 8018 17144 8024 17156
rect 8076 17144 8082 17196
rect 8202 17144 8208 17196
rect 8260 17144 8266 17196
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17085 5871 17119
rect 5813 17079 5871 17085
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17085 5963 17119
rect 5905 17079 5963 17085
rect 5920 17048 5948 17079
rect 6086 17076 6092 17128
rect 6144 17076 6150 17128
rect 6181 17119 6239 17125
rect 6181 17085 6193 17119
rect 6227 17085 6239 17119
rect 6181 17079 6239 17085
rect 6196 17048 6224 17079
rect 7374 17076 7380 17128
rect 7432 17076 7438 17128
rect 7558 17076 7564 17128
rect 7616 17076 7622 17128
rect 7653 17119 7711 17125
rect 7653 17085 7665 17119
rect 7699 17085 7711 17119
rect 7653 17079 7711 17085
rect 5736 17020 5948 17048
rect 6012 17020 6224 17048
rect 6012 16980 6040 17020
rect 6270 17008 6276 17060
rect 6328 17048 6334 17060
rect 6733 17051 6791 17057
rect 6733 17048 6745 17051
rect 6328 17020 6745 17048
rect 6328 17008 6334 17020
rect 6733 17017 6745 17020
rect 6779 17048 6791 17051
rect 7668 17048 7696 17079
rect 7742 17076 7748 17128
rect 7800 17076 7806 17128
rect 7926 17076 7932 17128
rect 7984 17076 7990 17128
rect 8220 17048 8248 17144
rect 8864 17116 8892 17292
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 9030 17144 9036 17196
rect 9088 17184 9094 17196
rect 9401 17187 9459 17193
rect 9401 17184 9413 17187
rect 9088 17156 9413 17184
rect 9088 17144 9094 17156
rect 9401 17153 9413 17156
rect 9447 17153 9459 17187
rect 9401 17147 9459 17153
rect 8941 17119 8999 17125
rect 8941 17116 8953 17119
rect 8864 17088 8953 17116
rect 8941 17085 8953 17088
rect 8987 17085 8999 17119
rect 9950 17116 9956 17128
rect 8941 17079 8999 17085
rect 9038 17088 9956 17116
rect 8478 17048 8484 17060
rect 6779 17020 8248 17048
rect 8312 17020 8484 17048
rect 6779 17017 6791 17020
rect 6733 17011 6791 17017
rect 5552 16952 6040 16980
rect 6086 16940 6092 16992
rect 6144 16980 6150 16992
rect 6365 16983 6423 16989
rect 6365 16980 6377 16983
rect 6144 16952 6377 16980
rect 6144 16940 6150 16952
rect 6365 16949 6377 16952
rect 6411 16949 6423 16983
rect 6365 16943 6423 16949
rect 7193 16983 7251 16989
rect 7193 16949 7205 16983
rect 7239 16980 7251 16983
rect 7742 16980 7748 16992
rect 7239 16952 7748 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7742 16940 7748 16952
rect 7800 16940 7806 16992
rect 8018 16940 8024 16992
rect 8076 16980 8082 16992
rect 8312 16980 8340 17020
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 8849 17051 8907 17057
rect 8849 17017 8861 17051
rect 8895 17048 8907 17051
rect 9038 17048 9066 17088
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 8895 17020 9066 17048
rect 9125 17051 9183 17057
rect 8895 17017 8907 17020
rect 8849 17011 8907 17017
rect 9125 17017 9137 17051
rect 9171 17048 9183 17051
rect 9490 17048 9496 17060
rect 9171 17020 9496 17048
rect 9171 17017 9183 17020
rect 9125 17011 9183 17017
rect 9490 17008 9496 17020
rect 9548 17008 9554 17060
rect 9674 17057 9680 17060
rect 9668 17011 9680 17057
rect 9674 17008 9680 17011
rect 9732 17008 9738 17060
rect 10226 17048 10232 17060
rect 9784 17020 10232 17048
rect 8076 16952 8340 16980
rect 8076 16940 8082 16952
rect 8386 16940 8392 16992
rect 8444 16980 8450 16992
rect 8573 16983 8631 16989
rect 8573 16980 8585 16983
rect 8444 16952 8585 16980
rect 8444 16940 8450 16952
rect 8573 16949 8585 16952
rect 8619 16949 8631 16983
rect 8573 16943 8631 16949
rect 8757 16983 8815 16989
rect 8757 16949 8769 16983
rect 8803 16980 8815 16983
rect 9784 16980 9812 17020
rect 10226 17008 10232 17020
rect 10284 17008 10290 17060
rect 8803 16952 9812 16980
rect 8803 16949 8815 16952
rect 8757 16943 8815 16949
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 9916 16952 10793 16980
rect 9916 16940 9922 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 10781 16943 10839 16949
rect 552 16890 11132 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 10722 16890
rect 10774 16838 10786 16890
rect 10838 16838 10850 16890
rect 10902 16838 10914 16890
rect 10966 16838 10978 16890
rect 11030 16838 11132 16890
rect 552 16816 11132 16838
rect 4982 16736 4988 16788
rect 5040 16736 5046 16788
rect 5718 16736 5724 16788
rect 5776 16776 5782 16788
rect 5813 16779 5871 16785
rect 5813 16776 5825 16779
rect 5776 16748 5825 16776
rect 5776 16736 5782 16748
rect 5813 16745 5825 16748
rect 5859 16745 5871 16779
rect 5813 16739 5871 16745
rect 6454 16736 6460 16788
rect 6512 16736 6518 16788
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 6880 16748 7144 16776
rect 6880 16736 6886 16748
rect 3050 16668 3056 16720
rect 3108 16708 3114 16720
rect 4430 16708 4436 16720
rect 3108 16680 4436 16708
rect 3108 16668 3114 16680
rect 4430 16668 4436 16680
rect 4488 16708 4494 16720
rect 7006 16708 7012 16720
rect 4488 16680 6224 16708
rect 4488 16668 4494 16680
rect 1578 16600 1584 16652
rect 1636 16640 1642 16652
rect 1765 16643 1823 16649
rect 1765 16640 1777 16643
rect 1636 16612 1777 16640
rect 1636 16600 1642 16612
rect 1765 16609 1777 16612
rect 1811 16609 1823 16643
rect 1765 16603 1823 16609
rect 2038 16600 2044 16652
rect 2096 16600 2102 16652
rect 2593 16643 2651 16649
rect 2593 16609 2605 16643
rect 2639 16640 2651 16643
rect 2958 16640 2964 16652
rect 2639 16612 2964 16640
rect 2639 16609 2651 16612
rect 2593 16603 2651 16609
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3329 16643 3387 16649
rect 3329 16609 3341 16643
rect 3375 16609 3387 16643
rect 3329 16603 3387 16609
rect 382 16532 388 16584
rect 440 16572 446 16584
rect 1213 16575 1271 16581
rect 1213 16572 1225 16575
rect 440 16544 1225 16572
rect 440 16532 446 16544
rect 1213 16541 1225 16544
rect 1259 16541 1271 16575
rect 1213 16535 1271 16541
rect 1946 16532 1952 16584
rect 2004 16572 2010 16584
rect 2222 16572 2228 16584
rect 2004 16544 2228 16572
rect 2004 16532 2010 16544
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16572 2467 16575
rect 2774 16572 2780 16584
rect 2455 16544 2780 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 2866 16532 2872 16584
rect 2924 16532 2930 16584
rect 3344 16572 3372 16603
rect 3418 16600 3424 16652
rect 3476 16640 3482 16652
rect 4157 16643 4215 16649
rect 4157 16640 4169 16643
rect 3476 16612 4169 16640
rect 3476 16600 3482 16612
rect 4157 16609 4169 16612
rect 4203 16640 4215 16643
rect 5077 16643 5135 16649
rect 5077 16640 5089 16643
rect 4203 16612 5089 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 5077 16609 5089 16612
rect 5123 16640 5135 16643
rect 5810 16640 5816 16652
rect 5123 16612 5816 16640
rect 5123 16609 5135 16612
rect 5077 16603 5135 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 5994 16600 6000 16652
rect 6052 16600 6058 16652
rect 6086 16600 6092 16652
rect 6144 16600 6150 16652
rect 6196 16649 6224 16680
rect 6288 16680 7012 16708
rect 6288 16649 6316 16680
rect 7006 16668 7012 16680
rect 7064 16668 7070 16720
rect 7116 16717 7144 16748
rect 7282 16736 7288 16788
rect 7340 16736 7346 16788
rect 7834 16736 7840 16788
rect 7892 16776 7898 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 7892 16748 8217 16776
rect 7892 16736 7898 16748
rect 8205 16745 8217 16748
rect 8251 16745 8263 16779
rect 8205 16739 8263 16745
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 8763 16779 8821 16785
rect 8763 16776 8775 16779
rect 8720 16748 8775 16776
rect 8720 16736 8726 16748
rect 8763 16745 8775 16748
rect 8809 16745 8821 16779
rect 8763 16739 8821 16745
rect 8849 16779 8907 16785
rect 8849 16745 8861 16779
rect 8895 16776 8907 16779
rect 9585 16779 9643 16785
rect 8895 16748 9536 16776
rect 8895 16745 8907 16748
rect 8849 16739 8907 16745
rect 7101 16711 7159 16717
rect 7101 16677 7113 16711
rect 7147 16677 7159 16711
rect 7101 16671 7159 16677
rect 7466 16668 7472 16720
rect 7524 16708 7530 16720
rect 7561 16711 7619 16717
rect 7561 16708 7573 16711
rect 7524 16680 7573 16708
rect 7524 16668 7530 16680
rect 7561 16677 7573 16680
rect 7607 16677 7619 16711
rect 7561 16671 7619 16677
rect 7742 16668 7748 16720
rect 7800 16668 7806 16720
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 8389 16711 8447 16717
rect 8389 16708 8401 16711
rect 8352 16680 8401 16708
rect 8352 16668 8358 16680
rect 8389 16677 8401 16680
rect 8435 16677 8447 16711
rect 8389 16671 8447 16677
rect 9401 16711 9459 16717
rect 9401 16677 9413 16711
rect 9447 16677 9459 16711
rect 9508 16708 9536 16748
rect 9585 16745 9597 16779
rect 9631 16776 9643 16779
rect 9766 16776 9772 16788
rect 9631 16748 9772 16776
rect 9631 16745 9643 16748
rect 9585 16739 9643 16745
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 10413 16779 10471 16785
rect 10413 16745 10425 16779
rect 10459 16776 10471 16779
rect 10502 16776 10508 16788
rect 10459 16748 10508 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 10502 16736 10508 16748
rect 10560 16736 10566 16788
rect 10226 16708 10232 16720
rect 9508 16680 9812 16708
rect 9401 16671 9459 16677
rect 6181 16643 6239 16649
rect 6181 16609 6193 16643
rect 6227 16609 6239 16643
rect 6181 16603 6239 16609
rect 6273 16643 6331 16649
rect 6273 16609 6285 16643
rect 6319 16609 6331 16643
rect 6273 16603 6331 16609
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16640 6699 16643
rect 6730 16640 6736 16652
rect 6687 16612 6736 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 6822 16600 6828 16652
rect 6880 16640 6886 16652
rect 6917 16643 6975 16649
rect 6917 16640 6929 16643
rect 6880 16612 6929 16640
rect 6880 16600 6886 16612
rect 6917 16609 6929 16612
rect 6963 16609 6975 16643
rect 6917 16603 6975 16609
rect 7926 16600 7932 16652
rect 7984 16640 7990 16652
rect 8113 16643 8171 16649
rect 8113 16640 8125 16643
rect 7984 16612 8125 16640
rect 7984 16600 7990 16612
rect 8113 16609 8125 16612
rect 8159 16609 8171 16643
rect 8665 16643 8723 16649
rect 8665 16640 8677 16643
rect 8113 16603 8171 16609
rect 8496 16612 8677 16640
rect 3344 16544 3464 16572
rect 3436 16504 3464 16544
rect 3510 16532 3516 16584
rect 3568 16532 3574 16584
rect 3878 16532 3884 16584
rect 3936 16532 3942 16584
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 4111 16544 5028 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 4080 16504 4108 16535
rect 5000 16516 5028 16544
rect 5166 16532 5172 16584
rect 5224 16532 5230 16584
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 7377 16575 7435 16581
rect 7377 16572 7389 16575
rect 6604 16544 7389 16572
rect 6604 16532 6610 16544
rect 7377 16541 7389 16544
rect 7423 16541 7435 16575
rect 8496 16572 8524 16612
rect 8665 16609 8677 16612
rect 8711 16609 8723 16643
rect 8665 16603 8723 16609
rect 8938 16600 8944 16652
rect 8996 16600 9002 16652
rect 9033 16643 9091 16649
rect 9033 16609 9045 16643
rect 9079 16640 9091 16643
rect 9122 16640 9128 16652
rect 9079 16612 9128 16640
rect 9079 16609 9091 16612
rect 9033 16603 9091 16609
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 9416 16640 9444 16671
rect 9416 16630 9674 16640
rect 9416 16612 9720 16630
rect 9646 16602 9720 16612
rect 7377 16535 7435 16541
rect 8404 16544 8524 16572
rect 3436 16476 4108 16504
rect 3528 16448 3556 16476
rect 4982 16464 4988 16516
rect 5040 16504 5046 16516
rect 6270 16504 6276 16516
rect 5040 16476 6276 16504
rect 5040 16464 5046 16476
rect 6270 16464 6276 16476
rect 6328 16464 6334 16516
rect 8404 16513 8432 16544
rect 9692 16513 9720 16602
rect 8389 16507 8447 16513
rect 8389 16473 8401 16507
rect 8435 16473 8447 16507
rect 8389 16467 8447 16473
rect 9677 16507 9735 16513
rect 9677 16473 9689 16507
rect 9723 16473 9735 16507
rect 9784 16504 9812 16680
rect 9876 16680 10232 16708
rect 9876 16649 9904 16680
rect 10226 16668 10232 16680
rect 10284 16708 10290 16720
rect 11054 16708 11060 16720
rect 10284 16680 11060 16708
rect 10284 16668 10290 16680
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 9861 16643 9919 16649
rect 9861 16609 9873 16643
rect 9907 16609 9919 16643
rect 9861 16603 9919 16609
rect 9950 16600 9956 16652
rect 10008 16640 10014 16652
rect 10321 16643 10379 16649
rect 10321 16640 10333 16643
rect 10008 16612 10333 16640
rect 10008 16600 10014 16612
rect 10321 16609 10333 16612
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 11330 16640 11336 16652
rect 10551 16612 11336 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 10045 16575 10103 16581
rect 10045 16541 10057 16575
rect 10091 16541 10103 16575
rect 10045 16535 10103 16541
rect 9950 16504 9956 16516
rect 9784 16476 9956 16504
rect 9677 16467 9735 16473
rect 9950 16464 9956 16476
rect 10008 16464 10014 16516
rect 10060 16504 10088 16535
rect 10134 16532 10140 16584
rect 10192 16532 10198 16584
rect 10318 16504 10324 16516
rect 10060 16476 10324 16504
rect 10318 16464 10324 16476
rect 10376 16504 10382 16516
rect 11054 16504 11060 16516
rect 10376 16476 11060 16504
rect 10376 16464 10382 16476
rect 11054 16464 11060 16476
rect 11112 16464 11118 16516
rect 2774 16396 2780 16448
rect 2832 16396 2838 16448
rect 2958 16396 2964 16448
rect 3016 16396 3022 16448
rect 3510 16396 3516 16448
rect 3568 16396 3574 16448
rect 4246 16396 4252 16448
rect 4304 16436 4310 16448
rect 4525 16439 4583 16445
rect 4525 16436 4537 16439
rect 4304 16408 4537 16436
rect 4304 16396 4310 16408
rect 4525 16405 4537 16408
rect 4571 16405 4583 16439
rect 4525 16399 4583 16405
rect 4617 16439 4675 16445
rect 4617 16405 4629 16439
rect 4663 16436 4675 16439
rect 4798 16436 4804 16448
rect 4663 16408 4804 16436
rect 4663 16405 4675 16408
rect 4617 16399 4675 16405
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 9398 16396 9404 16448
rect 9456 16396 9462 16448
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 10134 16436 10140 16448
rect 9548 16408 10140 16436
rect 9548 16396 9554 16408
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 552 16346 11132 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 10062 16346
rect 10114 16294 10126 16346
rect 10178 16294 10190 16346
rect 10242 16294 10254 16346
rect 10306 16294 10318 16346
rect 10370 16294 11132 16346
rect 552 16272 11132 16294
rect 934 16192 940 16244
rect 992 16232 998 16244
rect 1121 16235 1179 16241
rect 1121 16232 1133 16235
rect 992 16204 1133 16232
rect 992 16192 998 16204
rect 1121 16201 1133 16204
rect 1167 16201 1179 16235
rect 1121 16195 1179 16201
rect 2406 16192 2412 16244
rect 2464 16192 2470 16244
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 4065 16235 4123 16241
rect 4065 16232 4077 16235
rect 2832 16204 4077 16232
rect 2832 16192 2838 16204
rect 4065 16201 4077 16204
rect 4111 16201 4123 16235
rect 4065 16195 4123 16201
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 6822 16232 6828 16244
rect 6420 16204 6828 16232
rect 6420 16192 6426 16204
rect 6822 16192 6828 16204
rect 6880 16192 6886 16244
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 8389 16235 8447 16241
rect 8389 16232 8401 16235
rect 7616 16204 8401 16232
rect 7616 16192 7622 16204
rect 8389 16201 8401 16204
rect 8435 16201 8447 16235
rect 8389 16195 8447 16201
rect 8662 16192 8668 16244
rect 8720 16232 8726 16244
rect 8846 16232 8852 16244
rect 8720 16204 8852 16232
rect 8720 16192 8726 16204
rect 8846 16192 8852 16204
rect 8904 16232 8910 16244
rect 9217 16235 9275 16241
rect 9217 16232 9229 16235
rect 8904 16204 9229 16232
rect 8904 16192 8910 16204
rect 9217 16201 9229 16204
rect 9263 16201 9275 16235
rect 9217 16195 9275 16201
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 10045 16235 10103 16241
rect 10045 16232 10057 16235
rect 10008 16204 10057 16232
rect 10008 16192 10014 16204
rect 10045 16201 10057 16204
rect 10091 16201 10103 16235
rect 10045 16195 10103 16201
rect 3050 16164 3056 16176
rect 2700 16136 3056 16164
rect 1581 16099 1639 16105
rect 1581 16096 1593 16099
rect 1320 16068 1593 16096
rect 1320 16037 1348 16068
rect 1581 16065 1593 16068
rect 1627 16065 1639 16099
rect 2498 16096 2504 16108
rect 1581 16059 1639 16065
rect 2056 16068 2504 16096
rect 1305 16031 1363 16037
rect 1305 15997 1317 16031
rect 1351 15997 1363 16031
rect 1305 15991 1363 15997
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 16028 1547 16031
rect 1670 16028 1676 16040
rect 1535 16000 1676 16028
rect 1535 15997 1547 16000
rect 1489 15991 1547 15997
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 16028 1823 16031
rect 1946 16028 1952 16040
rect 1811 16000 1952 16028
rect 1811 15997 1823 16000
rect 1765 15991 1823 15997
rect 1946 15988 1952 16000
rect 2004 15988 2010 16040
rect 2056 16037 2084 16068
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 2700 16037 2728 16136
rect 3050 16124 3056 16136
rect 3108 16124 3114 16176
rect 3237 16167 3295 16173
rect 3237 16133 3249 16167
rect 3283 16133 3295 16167
rect 5442 16164 5448 16176
rect 3237 16127 3295 16133
rect 4356 16136 5448 16164
rect 3252 16096 3280 16127
rect 2884 16068 3280 16096
rect 2884 16037 2912 16068
rect 3418 16056 3424 16108
rect 3476 16096 3482 16108
rect 3697 16099 3755 16105
rect 3697 16096 3709 16099
rect 3476 16068 3709 16096
rect 3476 16056 3482 16068
rect 3697 16065 3709 16068
rect 3743 16065 3755 16099
rect 3697 16059 3755 16065
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16065 3847 16099
rect 3789 16059 3847 16065
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 2685 16031 2743 16037
rect 2685 15997 2697 16031
rect 2731 15997 2743 16031
rect 2685 15991 2743 15997
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 15997 2835 16031
rect 2777 15991 2835 15997
rect 2869 16031 2927 16037
rect 2869 15997 2881 16031
rect 2915 15997 2927 16031
rect 2869 15991 2927 15997
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 16028 3111 16031
rect 3142 16028 3148 16040
rect 3099 16000 3148 16028
rect 3099 15997 3111 16000
rect 3053 15991 3111 15997
rect 2498 15920 2504 15972
rect 2556 15960 2562 15972
rect 2792 15960 2820 15991
rect 3142 15988 3148 16000
rect 3200 15988 3206 16040
rect 3510 15988 3516 16040
rect 3568 16028 3574 16040
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 3568 16000 3617 16028
rect 3568 15988 3574 16000
rect 3605 15997 3617 16000
rect 3651 15997 3663 16031
rect 3605 15991 3663 15997
rect 3804 15960 3832 16059
rect 4246 16056 4252 16108
rect 4304 16056 4310 16108
rect 4356 16105 4384 16136
rect 5442 16124 5448 16136
rect 5500 16124 5506 16176
rect 9033 16167 9091 16173
rect 9033 16164 9045 16167
rect 8680 16136 9045 16164
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 4430 16056 4436 16108
rect 4488 16056 4494 16108
rect 8680 16105 8708 16136
rect 9033 16133 9045 16136
rect 9079 16133 9091 16167
rect 9033 16127 9091 16133
rect 4525 16099 4583 16105
rect 4525 16065 4537 16099
rect 4571 16096 4583 16099
rect 4801 16099 4859 16105
rect 4801 16096 4813 16099
rect 4571 16068 4813 16096
rect 4571 16065 4583 16068
rect 4525 16059 4583 16065
rect 4801 16065 4813 16068
rect 4847 16065 4859 16099
rect 4801 16059 4859 16065
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16065 8723 16099
rect 9306 16096 9312 16108
rect 8665 16059 8723 16065
rect 8772 16068 9312 16096
rect 4706 15988 4712 16040
rect 4764 15988 4770 16040
rect 4890 15988 4896 16040
rect 4948 15988 4954 16040
rect 8570 15988 8576 16040
rect 8628 15988 8634 16040
rect 8772 16037 8800 16068
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 9398 16056 9404 16108
rect 9456 16096 9462 16108
rect 9456 16068 9720 16096
rect 9456 16056 9462 16068
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 2556 15932 2820 15960
rect 3252 15932 3832 15960
rect 2556 15920 2562 15932
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 1949 15895 2007 15901
rect 1949 15892 1961 15895
rect 1452 15864 1961 15892
rect 1452 15852 1458 15864
rect 1949 15861 1961 15864
rect 1995 15861 2007 15895
rect 1949 15855 2007 15861
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 3252 15892 3280 15932
rect 6270 15920 6276 15972
rect 6328 15960 6334 15972
rect 8772 15960 8800 15991
rect 8846 15988 8852 16040
rect 8904 15988 8910 16040
rect 9214 15988 9220 16040
rect 9272 15988 9278 16040
rect 9692 16037 9720 16068
rect 9585 16031 9643 16037
rect 9585 15997 9597 16031
rect 9631 15997 9643 16031
rect 9585 15991 9643 15997
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 6328 15932 8800 15960
rect 9600 15960 9628 15991
rect 9766 15960 9772 15972
rect 9600 15932 9772 15960
rect 6328 15920 6334 15932
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 9861 15963 9919 15969
rect 9861 15929 9873 15963
rect 9907 15929 9919 15963
rect 9861 15923 9919 15929
rect 2372 15864 3280 15892
rect 2372 15852 2378 15864
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 9876 15892 9904 15923
rect 9364 15864 9904 15892
rect 9364 15852 9370 15864
rect 552 15802 11132 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 10722 15802
rect 10774 15750 10786 15802
rect 10838 15750 10850 15802
rect 10902 15750 10914 15802
rect 10966 15750 10978 15802
rect 11030 15750 11132 15802
rect 552 15728 11132 15750
rect 2409 15691 2467 15697
rect 2409 15657 2421 15691
rect 2455 15688 2467 15691
rect 2498 15688 2504 15700
rect 2455 15660 2504 15688
rect 2455 15657 2467 15660
rect 2409 15651 2467 15657
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 2869 15691 2927 15697
rect 2869 15657 2881 15691
rect 2915 15688 2927 15691
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 2915 15660 3341 15688
rect 2915 15657 2927 15660
rect 2869 15651 2927 15657
rect 3329 15657 3341 15660
rect 3375 15657 3387 15691
rect 3329 15651 3387 15657
rect 4062 15648 4068 15700
rect 4120 15688 4126 15700
rect 4341 15691 4399 15697
rect 4341 15688 4353 15691
rect 4120 15660 4353 15688
rect 4120 15648 4126 15660
rect 4341 15657 4353 15660
rect 4387 15657 4399 15691
rect 4341 15651 4399 15657
rect 6178 15648 6184 15700
rect 6236 15648 6242 15700
rect 6822 15688 6828 15700
rect 6472 15660 6828 15688
rect 1946 15580 1952 15632
rect 2004 15620 2010 15632
rect 3605 15623 3663 15629
rect 2004 15592 3096 15620
rect 2004 15580 2010 15592
rect 2130 15512 2136 15564
rect 2188 15512 2194 15564
rect 2682 15512 2688 15564
rect 2740 15512 2746 15564
rect 2958 15512 2964 15564
rect 3016 15512 3022 15564
rect 3068 15561 3096 15592
rect 3605 15589 3617 15623
rect 3651 15620 3663 15623
rect 4154 15620 4160 15632
rect 3651 15592 4160 15620
rect 3651 15589 3663 15592
rect 3605 15583 3663 15589
rect 4154 15580 4160 15592
rect 4212 15620 4218 15632
rect 4982 15620 4988 15632
rect 4212 15592 4988 15620
rect 4212 15580 4218 15592
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 6472 15629 6500 15660
rect 6822 15648 6828 15660
rect 6880 15688 6886 15700
rect 7098 15688 7104 15700
rect 6880 15660 7104 15688
rect 6880 15648 6886 15660
rect 7098 15648 7104 15660
rect 7156 15688 7162 15700
rect 7650 15688 7656 15700
rect 7156 15660 7656 15688
rect 7156 15648 7162 15660
rect 7650 15648 7656 15660
rect 7708 15648 7714 15700
rect 7745 15691 7803 15697
rect 7745 15657 7757 15691
rect 7791 15688 7803 15691
rect 8386 15688 8392 15700
rect 7791 15660 8392 15688
rect 7791 15657 7803 15660
rect 7745 15651 7803 15657
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 8570 15648 8576 15700
rect 8628 15648 8634 15700
rect 9125 15691 9183 15697
rect 9125 15657 9137 15691
rect 9171 15688 9183 15691
rect 9306 15688 9312 15700
rect 9171 15660 9312 15688
rect 9171 15657 9183 15660
rect 9125 15651 9183 15657
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 9490 15648 9496 15700
rect 9548 15648 9554 15700
rect 10229 15691 10287 15697
rect 10229 15688 10241 15691
rect 9692 15660 10241 15688
rect 6457 15623 6515 15629
rect 6457 15589 6469 15623
rect 6503 15589 6515 15623
rect 6457 15583 6515 15589
rect 7466 15580 7472 15632
rect 7524 15620 7530 15632
rect 8588 15620 8616 15648
rect 9508 15620 9536 15648
rect 9692 15629 9720 15660
rect 10229 15657 10241 15660
rect 10275 15657 10287 15691
rect 10229 15651 10287 15657
rect 7524 15592 8616 15620
rect 8770 15592 9536 15620
rect 9677 15623 9735 15629
rect 7524 15580 7530 15592
rect 3053 15555 3111 15561
rect 3053 15521 3065 15555
rect 3099 15521 3111 15555
rect 3053 15515 3111 15521
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15521 3295 15555
rect 3237 15515 3295 15521
rect 3513 15555 3571 15561
rect 3513 15521 3525 15555
rect 3559 15521 3571 15555
rect 3513 15515 3571 15521
rect 2406 15444 2412 15496
rect 2464 15444 2470 15496
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 2590 15484 2596 15496
rect 2547 15456 2596 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 2866 15444 2872 15496
rect 2924 15484 2930 15496
rect 3252 15484 3280 15515
rect 2924 15456 3280 15484
rect 2924 15444 2930 15456
rect 1762 15376 1768 15428
rect 1820 15416 1826 15428
rect 3053 15419 3111 15425
rect 3053 15416 3065 15419
rect 1820 15388 3065 15416
rect 1820 15376 1826 15388
rect 3053 15385 3065 15388
rect 3099 15385 3111 15419
rect 3528 15416 3556 15515
rect 3694 15512 3700 15564
rect 3752 15512 3758 15564
rect 3881 15555 3939 15561
rect 3881 15521 3893 15555
rect 3927 15521 3939 15555
rect 3881 15515 3939 15521
rect 3973 15555 4031 15561
rect 3973 15521 3985 15555
rect 4019 15552 4031 15555
rect 4525 15555 4583 15561
rect 4525 15552 4537 15555
rect 4019 15524 4537 15552
rect 4019 15521 4031 15524
rect 3973 15515 4031 15521
rect 4525 15521 4537 15524
rect 4571 15521 4583 15555
rect 4525 15515 4583 15521
rect 3896 15484 3924 15515
rect 4062 15484 4068 15496
rect 3896 15456 4068 15484
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 4540 15484 4568 15515
rect 4798 15512 4804 15564
rect 4856 15512 4862 15564
rect 6270 15512 6276 15564
rect 6328 15552 6334 15564
rect 6365 15555 6423 15561
rect 6365 15552 6377 15555
rect 6328 15524 6377 15552
rect 6328 15512 6334 15524
rect 6365 15521 6377 15524
rect 6411 15521 6423 15555
rect 6365 15515 6423 15521
rect 6546 15512 6552 15564
rect 6604 15512 6610 15564
rect 6730 15512 6736 15564
rect 6788 15512 6794 15564
rect 6825 15555 6883 15561
rect 6825 15521 6837 15555
rect 6871 15552 6883 15555
rect 7190 15552 7196 15564
rect 6871 15524 7196 15552
rect 6871 15521 6883 15524
rect 6825 15515 6883 15521
rect 5810 15484 5816 15496
rect 4540 15456 5816 15484
rect 5810 15444 5816 15456
rect 5868 15484 5874 15496
rect 6840 15484 6868 15515
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 7340 15524 7389 15552
rect 7340 15512 7346 15524
rect 7377 15521 7389 15524
rect 7423 15521 7435 15555
rect 7377 15515 7435 15521
rect 7834 15512 7840 15564
rect 7892 15512 7898 15564
rect 8021 15555 8079 15561
rect 8021 15521 8033 15555
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 8113 15555 8171 15561
rect 8113 15521 8125 15555
rect 8159 15552 8171 15555
rect 8202 15552 8208 15564
rect 8159 15524 8208 15552
rect 8159 15521 8171 15524
rect 8113 15515 8171 15521
rect 5868 15456 6868 15484
rect 7469 15487 7527 15493
rect 5868 15444 5874 15456
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 8036 15484 8064 15515
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8386 15512 8392 15564
rect 8444 15512 8450 15564
rect 8662 15512 8668 15564
rect 8720 15512 8726 15564
rect 8770 15484 8798 15592
rect 9677 15589 9689 15623
rect 9723 15589 9735 15623
rect 9677 15583 9735 15589
rect 9766 15580 9772 15632
rect 9824 15620 9830 15632
rect 10381 15623 10439 15629
rect 10381 15620 10393 15623
rect 9824 15592 10393 15620
rect 9824 15580 9830 15592
rect 10381 15589 10393 15592
rect 10427 15589 10439 15623
rect 10381 15583 10439 15589
rect 10597 15623 10655 15629
rect 10597 15589 10609 15623
rect 10643 15620 10655 15623
rect 10686 15620 10692 15632
rect 10643 15592 10692 15620
rect 10643 15589 10655 15592
rect 10597 15583 10655 15589
rect 10686 15580 10692 15592
rect 10744 15580 10750 15632
rect 8849 15555 8907 15561
rect 8849 15521 8861 15555
rect 8895 15521 8907 15555
rect 8849 15515 8907 15521
rect 8941 15555 8999 15561
rect 8941 15521 8953 15555
rect 8987 15552 8999 15555
rect 9217 15555 9275 15561
rect 8987 15524 9168 15552
rect 8987 15521 8999 15524
rect 8941 15515 8999 15521
rect 7515 15456 7880 15484
rect 8036 15456 8798 15484
rect 8864 15484 8892 15515
rect 9140 15484 9168 15524
rect 9217 15521 9229 15555
rect 9263 15552 9275 15555
rect 9306 15552 9312 15564
rect 9263 15524 9312 15552
rect 9263 15521 9275 15524
rect 9217 15515 9275 15521
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 9490 15512 9496 15564
rect 9548 15512 9554 15564
rect 9950 15512 9956 15564
rect 10008 15512 10014 15564
rect 9582 15484 9588 15496
rect 8864 15456 9076 15484
rect 9140 15456 9588 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 4338 15416 4344 15428
rect 3528 15388 4344 15416
rect 3053 15379 3111 15385
rect 4338 15376 4344 15388
rect 4396 15376 4402 15428
rect 4614 15376 4620 15428
rect 4672 15376 4678 15428
rect 4709 15419 4767 15425
rect 4709 15385 4721 15419
rect 4755 15416 4767 15419
rect 4798 15416 4804 15428
rect 4755 15388 4804 15416
rect 4755 15385 4767 15388
rect 4709 15379 4767 15385
rect 4798 15376 4804 15388
rect 4856 15376 4862 15428
rect 2038 15308 2044 15360
rect 2096 15348 2102 15360
rect 2225 15351 2283 15357
rect 2225 15348 2237 15351
rect 2096 15320 2237 15348
rect 2096 15308 2102 15320
rect 2225 15317 2237 15320
rect 2271 15317 2283 15351
rect 2225 15311 2283 15317
rect 2958 15308 2964 15360
rect 3016 15348 3022 15360
rect 3326 15348 3332 15360
rect 3016 15320 3332 15348
rect 3016 15308 3022 15320
rect 3326 15308 3332 15320
rect 3384 15308 3390 15360
rect 7852 15357 7880 15456
rect 8770 15416 8798 15456
rect 8846 15416 8852 15428
rect 8770 15388 8852 15416
rect 8846 15376 8852 15388
rect 8904 15376 8910 15428
rect 8938 15376 8944 15428
rect 8996 15376 9002 15428
rect 9048 15416 9076 15456
rect 9214 15416 9220 15428
rect 9048 15388 9220 15416
rect 9214 15376 9220 15388
rect 9272 15376 9278 15428
rect 7837 15351 7895 15357
rect 7837 15317 7849 15351
rect 7883 15348 7895 15351
rect 8202 15348 8208 15360
rect 7883 15320 8208 15348
rect 7883 15317 7895 15320
rect 7837 15311 7895 15317
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 8570 15308 8576 15360
rect 8628 15348 8634 15360
rect 9324 15348 9352 15456
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 10137 15487 10195 15493
rect 10137 15453 10149 15487
rect 10183 15484 10195 15487
rect 10183 15456 10456 15484
rect 10183 15453 10195 15456
rect 10137 15447 10195 15453
rect 8628 15320 9352 15348
rect 8628 15308 8634 15320
rect 9398 15308 9404 15360
rect 9456 15348 9462 15360
rect 10428 15357 10456 15456
rect 9769 15351 9827 15357
rect 9769 15348 9781 15351
rect 9456 15320 9781 15348
rect 9456 15308 9462 15320
rect 9769 15317 9781 15320
rect 9815 15317 9827 15351
rect 9769 15311 9827 15317
rect 10413 15351 10471 15357
rect 10413 15317 10425 15351
rect 10459 15348 10471 15351
rect 10594 15348 10600 15360
rect 10459 15320 10600 15348
rect 10459 15317 10471 15320
rect 10413 15311 10471 15317
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 552 15258 11132 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 10062 15258
rect 10114 15206 10126 15258
rect 10178 15206 10190 15258
rect 10242 15206 10254 15258
rect 10306 15206 10318 15258
rect 10370 15206 11132 15258
rect 552 15184 11132 15206
rect 2222 15104 2228 15156
rect 2280 15104 2286 15156
rect 2314 15104 2320 15156
rect 2372 15144 2378 15156
rect 4154 15144 4160 15156
rect 2372 15116 4160 15144
rect 2372 15104 2378 15116
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 4614 15104 4620 15156
rect 4672 15144 4678 15156
rect 5169 15147 5227 15153
rect 5169 15144 5181 15147
rect 4672 15116 5181 15144
rect 4672 15104 4678 15116
rect 5169 15113 5181 15116
rect 5215 15113 5227 15147
rect 5169 15107 5227 15113
rect 5353 15147 5411 15153
rect 5353 15113 5365 15147
rect 5399 15113 5411 15147
rect 5353 15107 5411 15113
rect 1486 15036 1492 15088
rect 1544 15076 1550 15088
rect 1544 15048 2636 15076
rect 1544 15036 1550 15048
rect 1213 15011 1271 15017
rect 1213 14977 1225 15011
rect 1259 15008 1271 15011
rect 1857 15011 1915 15017
rect 1857 15008 1869 15011
rect 1259 14980 1869 15008
rect 1259 14977 1271 14980
rect 1213 14971 1271 14977
rect 1857 14977 1869 14980
rect 1903 14977 1915 15011
rect 1857 14971 1915 14977
rect 2130 14968 2136 15020
rect 2188 15008 2194 15020
rect 2188 14980 2452 15008
rect 2188 14968 2194 14980
rect 2424 14952 2452 14980
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1578 14940 1584 14952
rect 1443 14912 1584 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1578 14900 1584 14912
rect 1636 14900 1642 14952
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14909 1731 14943
rect 1673 14903 1731 14909
rect 1688 14872 1716 14903
rect 1762 14900 1768 14952
rect 1820 14900 1826 14952
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 2317 14943 2375 14949
rect 2317 14940 2329 14943
rect 2087 14912 2329 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 2317 14909 2329 14912
rect 2363 14909 2375 14943
rect 2317 14903 2375 14909
rect 2406 14900 2412 14952
rect 2464 14940 2470 14952
rect 2501 14943 2559 14949
rect 2501 14940 2513 14943
rect 2464 14912 2513 14940
rect 2464 14900 2470 14912
rect 2501 14909 2513 14912
rect 2547 14909 2559 14943
rect 2501 14903 2559 14909
rect 1946 14872 1952 14884
rect 1688 14844 1952 14872
rect 1946 14832 1952 14844
rect 2004 14832 2010 14884
rect 2608 14872 2636 15048
rect 2682 15036 2688 15088
rect 2740 15076 2746 15088
rect 2740 15048 3096 15076
rect 2740 15036 2746 15048
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 15008 2835 15011
rect 2823 14980 3004 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 2682 14900 2688 14952
rect 2740 14900 2746 14952
rect 2866 14900 2872 14952
rect 2924 14900 2930 14952
rect 2884 14872 2912 14900
rect 2608 14844 2912 14872
rect 198 14764 204 14816
rect 256 14804 262 14816
rect 1486 14804 1492 14816
rect 256 14776 1492 14804
rect 256 14764 262 14776
rect 1486 14764 1492 14776
rect 1544 14804 1550 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 1544 14776 1593 14804
rect 1544 14764 1550 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 1581 14767 1639 14773
rect 1670 14764 1676 14816
rect 1728 14804 1734 14816
rect 2682 14804 2688 14816
rect 1728 14776 2688 14804
rect 1728 14764 1734 14776
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 2866 14764 2872 14816
rect 2924 14804 2930 14816
rect 2976 14804 3004 14980
rect 3068 14949 3096 15048
rect 3142 15036 3148 15088
rect 3200 15076 3206 15088
rect 3789 15079 3847 15085
rect 3789 15076 3801 15079
rect 3200 15048 3801 15076
rect 3200 15036 3206 15048
rect 3789 15045 3801 15048
rect 3835 15045 3847 15079
rect 3789 15039 3847 15045
rect 4893 15079 4951 15085
rect 4893 15045 4905 15079
rect 4939 15076 4951 15079
rect 5368 15076 5396 15107
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 6457 15147 6515 15153
rect 6457 15144 6469 15147
rect 6144 15116 6469 15144
rect 6144 15104 6150 15116
rect 6457 15113 6469 15116
rect 6503 15113 6515 15147
rect 6457 15107 6515 15113
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 7064 15116 8064 15144
rect 7064 15104 7070 15116
rect 4939 15048 5396 15076
rect 4939 15045 4951 15048
rect 4893 15039 4951 15045
rect 3694 14968 3700 15020
rect 3752 15008 3758 15020
rect 4908 15008 4936 15039
rect 5534 15036 5540 15088
rect 5592 15076 5598 15088
rect 8036 15076 8064 15116
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 8168 15116 8677 15144
rect 8168 15104 8174 15116
rect 8665 15113 8677 15116
rect 8711 15113 8723 15147
rect 8665 15107 8723 15113
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 8849 15147 8907 15153
rect 8849 15144 8861 15147
rect 8812 15116 8861 15144
rect 8812 15104 8818 15116
rect 8849 15113 8861 15116
rect 8895 15113 8907 15147
rect 8849 15107 8907 15113
rect 8938 15104 8944 15156
rect 8996 15144 9002 15156
rect 9398 15144 9404 15156
rect 8996 15116 9404 15144
rect 8996 15104 9002 15116
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 10008 15116 10149 15144
rect 10008 15104 10014 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 8570 15076 8576 15088
rect 5592 15048 7972 15076
rect 8036 15048 8576 15076
rect 5592 15036 5598 15048
rect 3752 14980 4936 15008
rect 3752 14968 3758 14980
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14940 3111 14943
rect 3970 14940 3976 14952
rect 3099 14912 3976 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 4080 14949 4108 14980
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 6178 15008 6184 15020
rect 5408 14980 6184 15008
rect 5408 14968 5414 14980
rect 6178 14968 6184 14980
rect 6236 15008 6242 15020
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6236 14980 6653 15008
rect 6236 14968 6242 14980
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 7466 14968 7472 15020
rect 7524 14968 7530 15020
rect 7561 15011 7619 15017
rect 7561 14977 7573 15011
rect 7607 15008 7619 15011
rect 7742 15008 7748 15020
rect 7607 14980 7748 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 7742 14968 7748 14980
rect 7800 15008 7806 15020
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 7800 14980 7849 15008
rect 7800 14968 7806 14980
rect 7837 14977 7849 14980
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 4065 14943 4123 14949
rect 4065 14909 4077 14943
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14940 4675 14943
rect 4706 14940 4712 14952
rect 4663 14912 4712 14940
rect 4663 14909 4675 14912
rect 4617 14903 4675 14909
rect 4706 14900 4712 14912
rect 4764 14900 4770 14952
rect 4890 14900 4896 14952
rect 4948 14900 4954 14952
rect 5074 14900 5080 14952
rect 5132 14900 5138 14952
rect 5810 14900 5816 14952
rect 5868 14900 5874 14952
rect 5902 14900 5908 14952
rect 5960 14900 5966 14952
rect 6270 14940 6276 14952
rect 6012 14912 6276 14940
rect 3326 14832 3332 14884
rect 3384 14832 3390 14884
rect 3418 14832 3424 14884
rect 3476 14872 3482 14884
rect 3513 14875 3571 14881
rect 3513 14872 3525 14875
rect 3476 14844 3525 14872
rect 3476 14832 3482 14844
rect 3513 14841 3525 14844
rect 3559 14841 3571 14875
rect 3513 14835 3571 14841
rect 3789 14875 3847 14881
rect 3789 14841 3801 14875
rect 3835 14872 3847 14875
rect 3878 14872 3884 14884
rect 3835 14844 3884 14872
rect 3835 14841 3847 14844
rect 3789 14835 3847 14841
rect 3878 14832 3884 14844
rect 3936 14832 3942 14884
rect 4338 14832 4344 14884
rect 4396 14872 4402 14884
rect 5537 14875 5595 14881
rect 5537 14872 5549 14875
rect 4396 14844 5549 14872
rect 4396 14832 4402 14844
rect 5537 14841 5549 14844
rect 5583 14872 5595 14875
rect 6012 14872 6040 14912
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 6733 14943 6791 14949
rect 6733 14940 6745 14943
rect 6512 14912 6745 14940
rect 6512 14900 6518 14912
rect 6733 14909 6745 14912
rect 6779 14909 6791 14943
rect 7098 14940 7104 14952
rect 6733 14903 6791 14909
rect 6932 14912 7104 14940
rect 6932 14884 6960 14912
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 7374 14900 7380 14952
rect 7432 14900 7438 14952
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 7944 14940 7972 15048
rect 8570 15036 8576 15048
rect 8628 15036 8634 15088
rect 9125 15079 9183 15085
rect 9125 15076 9137 15079
rect 8673 15048 9137 15076
rect 8673 15020 8701 15048
rect 9125 15045 9137 15048
rect 9171 15045 9183 15079
rect 9125 15039 9183 15045
rect 9217 15079 9275 15085
rect 9217 15045 9229 15079
rect 9263 15076 9275 15079
rect 9582 15076 9588 15088
rect 9263 15048 9588 15076
rect 9263 15045 9275 15048
rect 9217 15039 9275 15045
rect 9582 15036 9588 15048
rect 9640 15036 9646 15088
rect 8662 15008 8668 15020
rect 8496 14980 8668 15008
rect 7699 14912 7972 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 8202 14900 8208 14952
rect 8260 14900 8266 14952
rect 8496 14949 8524 14980
rect 8662 14968 8668 14980
rect 8720 14968 8726 15020
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 15008 8815 15011
rect 8938 15008 8944 15020
rect 8803 14980 8944 15008
rect 8803 14977 8815 14980
rect 8757 14971 8815 14977
rect 8938 14968 8944 14980
rect 8996 15008 9002 15020
rect 9398 15016 9404 15020
rect 9324 15008 9404 15016
rect 8996 14980 9066 15008
rect 8996 14968 9002 14980
rect 9038 14949 9066 14980
rect 9248 14988 9404 15008
rect 9248 14980 9352 14988
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14909 8539 14943
rect 8481 14903 8539 14909
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14909 9091 14943
rect 9248 14940 9276 14980
rect 9398 14968 9404 14988
rect 9456 14968 9462 15020
rect 9953 15011 10011 15017
rect 9953 14977 9965 15011
rect 9999 15008 10011 15011
rect 10226 15008 10232 15020
rect 9999 14980 10232 15008
rect 9999 14977 10011 14980
rect 9953 14971 10011 14977
rect 10226 14968 10232 14980
rect 10284 15008 10290 15020
rect 10284 14980 10456 15008
rect 10284 14968 10290 14980
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 9248 14912 9321 14940
rect 9033 14903 9091 14909
rect 9309 14909 9321 14912
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 9861 14943 9919 14949
rect 9861 14909 9873 14943
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 5583 14844 6040 14872
rect 5583 14841 5595 14844
rect 5537 14835 5595 14841
rect 6086 14832 6092 14884
rect 6144 14832 6150 14884
rect 6181 14875 6239 14881
rect 6181 14841 6193 14875
rect 6227 14872 6239 14875
rect 6914 14872 6920 14884
rect 6227 14844 6920 14872
rect 6227 14841 6239 14844
rect 6181 14835 6239 14841
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7282 14872 7288 14884
rect 7116 14844 7288 14872
rect 2924 14776 3004 14804
rect 3697 14807 3755 14813
rect 2924 14764 2930 14776
rect 3697 14773 3709 14807
rect 3743 14804 3755 14807
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 3743 14776 3985 14804
rect 3743 14773 3755 14776
rect 3697 14767 3755 14773
rect 3973 14773 3985 14776
rect 4019 14804 4031 14807
rect 4154 14804 4160 14816
rect 4019 14776 4160 14804
rect 4019 14773 4031 14776
rect 3973 14767 4031 14773
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 5350 14813 5356 14816
rect 5337 14807 5356 14813
rect 5337 14773 5349 14807
rect 5337 14767 5356 14773
rect 5350 14764 5356 14767
rect 5408 14764 5414 14816
rect 7116 14813 7144 14844
rect 7282 14832 7288 14844
rect 7340 14872 7346 14884
rect 8021 14875 8079 14881
rect 8021 14872 8033 14875
rect 7340 14844 8033 14872
rect 7340 14832 7346 14844
rect 8021 14841 8033 14844
rect 8067 14841 8079 14875
rect 8588 14872 8616 14903
rect 8754 14872 8760 14884
rect 8588 14844 8760 14872
rect 8021 14835 8079 14841
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 9876 14872 9904 14903
rect 10318 14900 10324 14952
rect 10376 14900 10382 14952
rect 10428 14949 10456 14980
rect 10413 14943 10471 14949
rect 10413 14909 10425 14943
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 10686 14940 10692 14952
rect 10551 14912 10692 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 10520 14872 10548 14903
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 9416 14844 10548 14872
rect 7101 14807 7159 14813
rect 7101 14773 7113 14807
rect 7147 14773 7159 14807
rect 7101 14767 7159 14773
rect 7190 14764 7196 14816
rect 7248 14764 7254 14816
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9416 14804 9444 14844
rect 10428 14816 10456 14844
rect 8996 14776 9444 14804
rect 9493 14807 9551 14813
rect 8996 14764 9002 14776
rect 9493 14773 9505 14807
rect 9539 14804 9551 14807
rect 10318 14804 10324 14816
rect 9539 14776 10324 14804
rect 9539 14773 9551 14776
rect 9493 14767 9551 14773
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 10410 14764 10416 14816
rect 10468 14764 10474 14816
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 10689 14807 10747 14813
rect 10689 14804 10701 14807
rect 10652 14776 10701 14804
rect 10652 14764 10658 14776
rect 10689 14773 10701 14776
rect 10735 14773 10747 14807
rect 10689 14767 10747 14773
rect 552 14714 11132 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 10722 14714
rect 10774 14662 10786 14714
rect 10838 14662 10850 14714
rect 10902 14662 10914 14714
rect 10966 14662 10978 14714
rect 11030 14662 11132 14714
rect 552 14640 11132 14662
rect 1762 14560 1768 14612
rect 1820 14600 1826 14612
rect 1857 14603 1915 14609
rect 1857 14600 1869 14603
rect 1820 14572 1869 14600
rect 1820 14560 1826 14572
rect 1857 14569 1869 14572
rect 1903 14569 1915 14603
rect 1857 14563 1915 14569
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2130 14600 2136 14612
rect 2004 14572 2136 14600
rect 2004 14560 2010 14572
rect 2130 14560 2136 14572
rect 2188 14560 2194 14612
rect 2590 14560 2596 14612
rect 2648 14560 2654 14612
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 2961 14603 3019 14609
rect 2961 14600 2973 14603
rect 2740 14572 2973 14600
rect 2740 14560 2746 14572
rect 2961 14569 2973 14572
rect 3007 14569 3019 14603
rect 2961 14563 3019 14569
rect 3053 14603 3111 14609
rect 3053 14569 3065 14603
rect 3099 14600 3111 14603
rect 3234 14600 3240 14612
rect 3099 14572 3240 14600
rect 3099 14569 3111 14572
rect 3053 14563 3111 14569
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 3510 14560 3516 14612
rect 3568 14600 3574 14612
rect 4338 14600 4344 14612
rect 3568 14572 4344 14600
rect 3568 14560 3574 14572
rect 4338 14560 4344 14572
rect 4396 14560 4402 14612
rect 5261 14603 5319 14609
rect 5261 14569 5273 14603
rect 5307 14600 5319 14603
rect 5350 14600 5356 14612
rect 5307 14572 5356 14600
rect 5307 14569 5319 14572
rect 5261 14563 5319 14569
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 5442 14560 5448 14612
rect 5500 14600 5506 14612
rect 6365 14603 6423 14609
rect 5500 14572 6132 14600
rect 5500 14560 5506 14572
rect 2608 14532 2636 14560
rect 3970 14532 3976 14544
rect 2332 14504 2636 14532
rect 3252 14504 3464 14532
rect 1486 14424 1492 14476
rect 1544 14424 1550 14476
rect 2332 14473 2360 14504
rect 3252 14476 3280 14504
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14433 2375 14467
rect 2317 14427 2375 14433
rect 2498 14424 2504 14476
rect 2556 14424 2562 14476
rect 2590 14424 2596 14476
rect 2648 14424 2654 14476
rect 2685 14467 2743 14473
rect 2685 14433 2697 14467
rect 2731 14464 2743 14467
rect 3142 14464 3148 14476
rect 2731 14436 3148 14464
rect 2731 14433 2743 14436
rect 2685 14427 2743 14433
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 3234 14424 3240 14476
rect 3292 14424 3298 14476
rect 3436 14473 3464 14504
rect 3804 14504 3976 14532
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 3421 14467 3479 14473
rect 3421 14433 3433 14467
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 1394 14356 1400 14408
rect 1452 14356 1458 14408
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 3344 14396 3372 14427
rect 3510 14424 3516 14476
rect 3568 14424 3574 14476
rect 3691 14467 3749 14473
rect 3691 14433 3703 14467
rect 3737 14462 3749 14467
rect 3804 14462 3832 14504
rect 3970 14492 3976 14504
rect 4028 14492 4034 14544
rect 5074 14532 5080 14544
rect 5000 14504 5080 14532
rect 3737 14434 3832 14462
rect 3737 14433 3749 14434
rect 3691 14427 3749 14433
rect 4154 14424 4160 14476
rect 4212 14424 4218 14476
rect 4706 14424 4712 14476
rect 4764 14424 4770 14476
rect 5000 14473 5028 14504
rect 5074 14492 5080 14504
rect 5132 14532 5138 14544
rect 5537 14535 5595 14541
rect 5537 14532 5549 14535
rect 5132 14504 5549 14532
rect 5132 14492 5138 14504
rect 5537 14501 5549 14504
rect 5583 14501 5595 14535
rect 6104 14532 6132 14572
rect 6365 14569 6377 14603
rect 6411 14600 6423 14603
rect 7374 14600 7380 14612
rect 6411 14572 7380 14600
rect 6411 14569 6423 14572
rect 6365 14563 6423 14569
rect 7374 14560 7380 14572
rect 7432 14600 7438 14612
rect 7432 14572 7604 14600
rect 7432 14560 7438 14572
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 6104 14504 6469 14532
rect 5537 14495 5595 14501
rect 6457 14501 6469 14504
rect 6503 14501 6515 14535
rect 6457 14495 6515 14501
rect 6638 14492 6644 14544
rect 6696 14492 6702 14544
rect 7190 14532 7196 14544
rect 6840 14504 7196 14532
rect 4985 14467 5043 14473
rect 4985 14433 4997 14467
rect 5031 14433 5043 14467
rect 4985 14427 5043 14433
rect 5445 14467 5503 14473
rect 5445 14433 5457 14467
rect 5491 14433 5503 14467
rect 5445 14427 5503 14433
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14439 5764 14467
rect 5675 14433 5687 14439
rect 5629 14427 5687 14433
rect 2464 14368 3464 14396
rect 2464 14356 2470 14368
rect 3436 14328 3464 14368
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3936 14368 3985 14396
rect 3936 14356 3942 14368
rect 3973 14365 3985 14368
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14396 4123 14399
rect 4249 14399 4307 14405
rect 4111 14368 4200 14396
rect 4111 14365 4123 14368
rect 4065 14359 4123 14365
rect 4172 14340 4200 14368
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 5350 14396 5356 14408
rect 4295 14368 5356 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 3436 14300 3924 14328
rect 2590 14220 2596 14272
rect 2648 14260 2654 14272
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 2648 14232 3801 14260
rect 2648 14220 2654 14232
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 3896 14260 3924 14300
rect 4154 14288 4160 14340
rect 4212 14288 4218 14340
rect 4264 14260 4292 14359
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 3896 14232 4292 14260
rect 3789 14223 3847 14229
rect 4890 14220 4896 14272
rect 4948 14260 4954 14272
rect 5074 14260 5080 14272
rect 4948 14232 5080 14260
rect 4948 14220 4954 14232
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 5350 14220 5356 14272
rect 5408 14260 5414 14272
rect 5460 14260 5488 14427
rect 5736 14396 5764 14439
rect 5810 14424 5816 14476
rect 5868 14464 5874 14476
rect 6022 14467 6080 14473
rect 6022 14464 6034 14467
rect 5868 14462 5948 14464
rect 6012 14462 6034 14464
rect 5868 14436 6034 14462
rect 5868 14424 5874 14436
rect 5920 14434 6034 14436
rect 6022 14433 6034 14434
rect 6068 14433 6080 14467
rect 6022 14427 6080 14433
rect 6549 14467 6607 14473
rect 6549 14433 6561 14467
rect 6595 14464 6607 14467
rect 6656 14464 6684 14492
rect 6840 14473 6868 14504
rect 7190 14492 7196 14504
rect 7248 14492 7254 14544
rect 7466 14492 7472 14544
rect 7524 14492 7530 14544
rect 7576 14541 7604 14572
rect 7742 14560 7748 14612
rect 7800 14560 7806 14612
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8662 14609 8668 14612
rect 8021 14603 8079 14609
rect 8021 14600 8033 14603
rect 7892 14572 8033 14600
rect 7892 14560 7898 14572
rect 8021 14569 8033 14572
rect 8067 14569 8079 14603
rect 8658 14600 8668 14609
rect 8623 14572 8668 14600
rect 8021 14563 8079 14569
rect 8658 14563 8668 14572
rect 8662 14560 8668 14563
rect 8720 14560 8726 14612
rect 9217 14603 9275 14609
rect 9217 14600 9229 14603
rect 8864 14572 9229 14600
rect 7561 14535 7619 14541
rect 7561 14501 7573 14535
rect 7607 14501 7619 14535
rect 7561 14495 7619 14501
rect 7650 14492 7656 14544
rect 7708 14532 7714 14544
rect 8864 14541 8892 14572
rect 9217 14569 9229 14572
rect 9263 14600 9275 14603
rect 9766 14600 9772 14612
rect 9263 14572 9772 14600
rect 9263 14569 9275 14572
rect 9217 14563 9275 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 10226 14560 10232 14612
rect 10284 14560 10290 14612
rect 10410 14560 10416 14612
rect 10468 14560 10474 14612
rect 8849 14535 8907 14541
rect 7708 14504 7972 14532
rect 7708 14492 7714 14504
rect 6595 14436 6684 14464
rect 6825 14467 6883 14473
rect 6595 14433 6607 14436
rect 6549 14427 6607 14433
rect 6825 14433 6837 14467
rect 6871 14433 6883 14467
rect 6825 14427 6883 14433
rect 6917 14467 6975 14473
rect 6917 14433 6929 14467
rect 6963 14464 6975 14467
rect 7374 14464 7380 14476
rect 6963 14436 7380 14464
rect 6963 14433 6975 14436
rect 6917 14427 6975 14433
rect 7374 14424 7380 14436
rect 7432 14424 7438 14476
rect 7484 14464 7512 14492
rect 7944 14473 7972 14504
rect 8849 14501 8861 14535
rect 8895 14501 8907 14535
rect 8849 14495 8907 14501
rect 8938 14492 8944 14544
rect 8996 14532 9002 14544
rect 9033 14535 9091 14541
rect 9033 14532 9045 14535
rect 8996 14504 9045 14532
rect 8996 14492 9002 14504
rect 9033 14501 9045 14504
rect 9079 14501 9091 14535
rect 10594 14532 10600 14544
rect 9033 14495 9091 14501
rect 9140 14504 10600 14532
rect 7837 14467 7895 14473
rect 7837 14464 7849 14467
rect 7484 14436 7849 14464
rect 7837 14433 7849 14436
rect 7883 14433 7895 14467
rect 7837 14427 7895 14433
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14433 7987 14467
rect 7929 14427 7987 14433
rect 8113 14467 8171 14473
rect 8113 14433 8125 14467
rect 8159 14464 8171 14467
rect 8297 14467 8355 14473
rect 8297 14464 8309 14467
rect 8159 14436 8309 14464
rect 8159 14433 8171 14436
rect 8113 14427 8171 14433
rect 8297 14433 8309 14436
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 8386 14424 8392 14476
rect 8444 14424 8450 14476
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14433 8539 14467
rect 8481 14427 8539 14433
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 8619 14436 8708 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 5905 14399 5963 14405
rect 5905 14396 5917 14399
rect 5736 14368 5917 14396
rect 5905 14365 5917 14368
rect 5951 14396 5963 14399
rect 6270 14396 6276 14408
rect 5951 14368 6276 14396
rect 5951 14365 5963 14368
rect 5905 14359 5963 14365
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 6638 14356 6644 14408
rect 6696 14356 6702 14408
rect 7009 14399 7067 14405
rect 7009 14365 7021 14399
rect 7055 14396 7067 14399
rect 7055 14368 7236 14396
rect 7055 14365 7067 14368
rect 7009 14359 7067 14365
rect 5994 14288 6000 14340
rect 6052 14328 6058 14340
rect 7101 14331 7159 14337
rect 7101 14328 7113 14331
rect 6052 14300 7113 14328
rect 6052 14288 6058 14300
rect 7101 14297 7113 14300
rect 7147 14297 7159 14331
rect 7101 14291 7159 14297
rect 7208 14272 7236 14368
rect 7282 14356 7288 14408
rect 7340 14396 7346 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 7340 14368 7481 14396
rect 7340 14356 7346 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 8496 14396 8524 14427
rect 7469 14359 7527 14365
rect 8128 14368 8524 14396
rect 8128 14340 8156 14368
rect 7374 14288 7380 14340
rect 7432 14328 7438 14340
rect 7561 14331 7619 14337
rect 7561 14328 7573 14331
rect 7432 14300 7573 14328
rect 7432 14288 7438 14300
rect 7561 14297 7573 14300
rect 7607 14297 7619 14331
rect 7561 14291 7619 14297
rect 8110 14288 8116 14340
rect 8168 14288 8174 14340
rect 8680 14328 8708 14436
rect 8754 14424 8760 14476
rect 8812 14424 8818 14476
rect 9140 14473 9168 14504
rect 10594 14492 10600 14504
rect 10652 14492 10658 14544
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14433 9183 14467
rect 9585 14467 9643 14473
rect 9585 14464 9597 14467
rect 9125 14427 9183 14433
rect 9232 14436 9597 14464
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 9232 14396 9260 14436
rect 9585 14433 9597 14436
rect 9631 14433 9643 14467
rect 9585 14427 9643 14433
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 9861 14467 9919 14473
rect 9861 14464 9873 14467
rect 9824 14436 9873 14464
rect 9824 14424 9830 14436
rect 9861 14433 9873 14436
rect 9907 14433 9919 14467
rect 9861 14427 9919 14433
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14433 10103 14467
rect 10045 14427 10103 14433
rect 8904 14368 9260 14396
rect 8904 14356 8910 14368
rect 9398 14356 9404 14408
rect 9456 14396 9462 14408
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 9456 14368 9505 14396
rect 9456 14356 9462 14368
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 10060 14396 10088 14427
rect 10318 14424 10324 14476
rect 10376 14424 10382 14476
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 11054 14464 11060 14476
rect 10551 14436 11060 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10520 14396 10548 14427
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 10594 14396 10600 14408
rect 10060 14368 10600 14396
rect 10060 14328 10088 14368
rect 10594 14356 10600 14368
rect 10652 14356 10658 14408
rect 8680 14300 10088 14328
rect 10318 14288 10324 14340
rect 10376 14328 10382 14340
rect 11146 14328 11152 14340
rect 10376 14300 11152 14328
rect 10376 14288 10382 14300
rect 11146 14288 11152 14300
rect 11204 14288 11210 14340
rect 5810 14260 5816 14272
rect 5408 14232 5816 14260
rect 5408 14220 5414 14232
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 7190 14220 7196 14272
rect 7248 14220 7254 14272
rect 8570 14220 8576 14272
rect 8628 14260 8634 14272
rect 8849 14263 8907 14269
rect 8849 14260 8861 14263
rect 8628 14232 8861 14260
rect 8628 14220 8634 14232
rect 8849 14229 8861 14232
rect 8895 14260 8907 14263
rect 9490 14260 9496 14272
rect 8895 14232 9496 14260
rect 8895 14229 8907 14232
rect 8849 14223 8907 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 10336 14260 10364 14288
rect 9824 14232 10364 14260
rect 9824 14220 9830 14232
rect 552 14170 11132 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 10062 14170
rect 10114 14118 10126 14170
rect 10178 14118 10190 14170
rect 10242 14118 10254 14170
rect 10306 14118 10318 14170
rect 10370 14118 11132 14170
rect 552 14096 11132 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1489 14059 1547 14065
rect 1489 14056 1501 14059
rect 1452 14028 1501 14056
rect 1452 14016 1458 14028
rect 1489 14025 1501 14028
rect 1535 14025 1547 14059
rect 1489 14019 1547 14025
rect 2409 14059 2467 14065
rect 2409 14025 2421 14059
rect 2455 14056 2467 14059
rect 3418 14056 3424 14068
rect 2455 14028 3424 14056
rect 2455 14025 2467 14028
rect 2409 14019 2467 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 3789 14059 3847 14065
rect 3789 14025 3801 14059
rect 3835 14056 3847 14059
rect 4706 14056 4712 14068
rect 3835 14028 4712 14056
rect 3835 14025 3847 14028
rect 3789 14019 3847 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 6270 14016 6276 14068
rect 6328 14056 6334 14068
rect 6457 14059 6515 14065
rect 6457 14056 6469 14059
rect 6328 14028 6469 14056
rect 6328 14016 6334 14028
rect 6457 14025 6469 14028
rect 6503 14025 6515 14059
rect 6457 14019 6515 14025
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8846 14056 8852 14068
rect 8536 14028 8852 14056
rect 8536 14016 8542 14028
rect 8846 14016 8852 14028
rect 8904 14016 8910 14068
rect 9769 14059 9827 14065
rect 9769 14056 9781 14059
rect 9248 14028 9781 14056
rect 2777 13991 2835 13997
rect 2777 13957 2789 13991
rect 2823 13957 2835 13991
rect 2777 13951 2835 13957
rect 1213 13923 1271 13929
rect 1213 13889 1225 13923
rect 1259 13920 1271 13923
rect 1394 13920 1400 13932
rect 1259 13892 1400 13920
rect 1259 13889 1271 13892
rect 1213 13883 1271 13889
rect 1394 13880 1400 13892
rect 1452 13920 1458 13932
rect 1670 13920 1676 13932
rect 1452 13892 1676 13920
rect 1452 13880 1458 13892
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 2038 13880 2044 13932
rect 2096 13880 2102 13932
rect 2590 13880 2596 13932
rect 2648 13920 2654 13932
rect 2792 13920 2820 13951
rect 3234 13948 3240 14000
rect 3292 13988 3298 14000
rect 3694 13988 3700 14000
rect 3292 13960 3700 13988
rect 3292 13948 3298 13960
rect 3694 13948 3700 13960
rect 3752 13948 3758 14000
rect 4249 13991 4307 13997
rect 4249 13957 4261 13991
rect 4295 13988 4307 13991
rect 4338 13988 4344 14000
rect 4295 13960 4344 13988
rect 4295 13957 4307 13960
rect 4249 13951 4307 13957
rect 4338 13948 4344 13960
rect 4396 13988 4402 14000
rect 4890 13988 4896 14000
rect 4396 13960 4896 13988
rect 4396 13948 4402 13960
rect 4890 13948 4896 13960
rect 4948 13948 4954 14000
rect 5169 13991 5227 13997
rect 5169 13957 5181 13991
rect 5215 13988 5227 13991
rect 5350 13988 5356 14000
rect 5215 13960 5356 13988
rect 5215 13957 5227 13960
rect 5169 13951 5227 13957
rect 5350 13948 5356 13960
rect 5408 13948 5414 14000
rect 5442 13948 5448 14000
rect 5500 13988 5506 14000
rect 7006 13988 7012 14000
rect 5500 13960 7012 13988
rect 5500 13948 5506 13960
rect 7006 13948 7012 13960
rect 7064 13948 7070 14000
rect 8754 13948 8760 14000
rect 8812 13988 8818 14000
rect 8938 13988 8944 14000
rect 8812 13960 8944 13988
rect 8812 13948 8818 13960
rect 8938 13948 8944 13960
rect 8996 13948 9002 14000
rect 2648 13892 2820 13920
rect 3605 13923 3663 13929
rect 2648 13880 2654 13892
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 3712 13920 3740 13948
rect 4709 13923 4767 13929
rect 4709 13920 4721 13923
rect 3712 13892 4721 13920
rect 3605 13883 3663 13889
rect 4709 13889 4721 13892
rect 4755 13889 4767 13923
rect 4709 13883 4767 13889
rect 1118 13812 1124 13864
rect 1176 13812 1182 13864
rect 1946 13812 1952 13864
rect 2004 13852 2010 13864
rect 2133 13855 2191 13861
rect 2133 13852 2145 13855
rect 2004 13824 2145 13852
rect 2004 13812 2010 13824
rect 2133 13821 2145 13824
rect 2179 13852 2191 13855
rect 2314 13852 2320 13864
rect 2179 13824 2320 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 3513 13855 3571 13861
rect 3513 13852 3525 13855
rect 3476 13824 3525 13852
rect 3476 13812 3482 13824
rect 3513 13821 3525 13824
rect 3559 13821 3571 13855
rect 3513 13815 3571 13821
rect 3620 13852 3648 13883
rect 7374 13880 7380 13932
rect 7432 13920 7438 13932
rect 8110 13920 8116 13932
rect 7432 13892 8116 13920
rect 7432 13880 7438 13892
rect 8110 13880 8116 13892
rect 8168 13920 8174 13932
rect 9248 13920 9276 14028
rect 9769 14025 9781 14028
rect 9815 14056 9827 14059
rect 11330 14056 11336 14068
rect 9815 14028 11336 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 9582 13948 9588 14000
rect 9640 13948 9646 14000
rect 8168 13892 9276 13920
rect 9401 13923 9459 13929
rect 8168 13880 8174 13892
rect 9401 13889 9413 13923
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 3878 13852 3884 13864
rect 3620 13824 3884 13852
rect 2222 13744 2228 13796
rect 2280 13784 2286 13796
rect 3053 13787 3111 13793
rect 3053 13784 3065 13787
rect 2280 13756 3065 13784
rect 2280 13744 2286 13756
rect 3053 13753 3065 13756
rect 3099 13784 3111 13787
rect 3142 13784 3148 13796
rect 3099 13756 3148 13784
rect 3099 13753 3111 13756
rect 3053 13747 3111 13753
rect 3142 13744 3148 13756
rect 3200 13744 3206 13796
rect 3326 13744 3332 13796
rect 3384 13784 3390 13796
rect 3620 13784 3648 13824
rect 3878 13812 3884 13824
rect 3936 13812 3942 13864
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4801 13855 4859 13861
rect 4801 13852 4813 13855
rect 4212 13824 4813 13852
rect 4212 13812 4218 13824
rect 4801 13821 4813 13824
rect 4847 13852 4859 13855
rect 5626 13852 5632 13864
rect 4847 13824 5632 13852
rect 4847 13821 4859 13824
rect 4801 13815 4859 13821
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 6178 13812 6184 13864
rect 6236 13812 6242 13864
rect 6457 13855 6515 13861
rect 6457 13821 6469 13855
rect 6503 13852 6515 13855
rect 7190 13852 7196 13864
rect 6503 13824 7196 13852
rect 6503 13821 6515 13824
rect 6457 13815 6515 13821
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 9309 13855 9367 13861
rect 9309 13852 9321 13855
rect 8536 13824 9321 13852
rect 8536 13812 8542 13824
rect 9309 13821 9321 13824
rect 9355 13821 9367 13855
rect 9309 13815 9367 13821
rect 3384 13756 3648 13784
rect 4525 13787 4583 13793
rect 3384 13744 3390 13756
rect 4525 13753 4537 13787
rect 4571 13784 4583 13787
rect 4706 13784 4712 13796
rect 4571 13756 4712 13784
rect 4571 13753 4583 13756
rect 4525 13747 4583 13753
rect 4706 13744 4712 13756
rect 4764 13784 4770 13796
rect 4982 13784 4988 13796
rect 4764 13756 4988 13784
rect 4764 13744 4770 13756
rect 4982 13744 4988 13756
rect 5040 13744 5046 13796
rect 6086 13744 6092 13796
rect 6144 13784 6150 13796
rect 7098 13784 7104 13796
rect 6144 13756 7104 13784
rect 6144 13744 6150 13756
rect 7098 13744 7104 13756
rect 7156 13744 7162 13796
rect 9214 13744 9220 13796
rect 9272 13784 9278 13796
rect 9416 13784 9444 13883
rect 9272 13756 9444 13784
rect 9272 13744 9278 13756
rect 9490 13744 9496 13796
rect 9548 13784 9554 13796
rect 9737 13787 9795 13793
rect 9737 13784 9749 13787
rect 9548 13756 9749 13784
rect 9548 13744 9554 13756
rect 9737 13753 9749 13756
rect 9783 13753 9795 13787
rect 9737 13747 9795 13753
rect 9953 13787 10011 13793
rect 9953 13753 9965 13787
rect 9999 13784 10011 13787
rect 10594 13784 10600 13796
rect 9999 13756 10600 13784
rect 9999 13753 10011 13756
rect 9953 13747 10011 13753
rect 10594 13744 10600 13756
rect 10652 13744 10658 13796
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 2593 13719 2651 13725
rect 2593 13716 2605 13719
rect 1820 13688 2605 13716
rect 1820 13676 1826 13688
rect 2593 13685 2605 13688
rect 2639 13685 2651 13719
rect 2593 13679 2651 13685
rect 4062 13676 4068 13728
rect 4120 13676 4126 13728
rect 6273 13719 6331 13725
rect 6273 13685 6285 13719
rect 6319 13716 6331 13719
rect 6454 13716 6460 13728
rect 6319 13688 6460 13716
rect 6319 13685 6331 13688
rect 6273 13679 6331 13685
rect 6454 13676 6460 13688
rect 6512 13716 6518 13728
rect 8754 13716 8760 13728
rect 6512 13688 8760 13716
rect 6512 13676 6518 13688
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 552 13626 11132 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 10722 13626
rect 10774 13574 10786 13626
rect 10838 13574 10850 13626
rect 10902 13574 10914 13626
rect 10966 13574 10978 13626
rect 11030 13574 11132 13626
rect 552 13552 11132 13574
rect 1486 13472 1492 13524
rect 1544 13512 1550 13524
rect 1581 13515 1639 13521
rect 1581 13512 1593 13515
rect 1544 13484 1593 13512
rect 1544 13472 1550 13484
rect 1581 13481 1593 13484
rect 1627 13481 1639 13515
rect 1581 13475 1639 13481
rect 1946 13472 1952 13524
rect 2004 13472 2010 13524
rect 2682 13472 2688 13524
rect 2740 13512 2746 13524
rect 2740 13484 3464 13512
rect 2740 13472 2746 13484
rect 2314 13404 2320 13456
rect 2372 13404 2378 13456
rect 1762 13336 1768 13388
rect 1820 13336 1826 13388
rect 2038 13336 2044 13388
rect 2096 13336 2102 13388
rect 2332 13376 2360 13404
rect 2593 13379 2651 13385
rect 2593 13376 2605 13379
rect 2332 13348 2605 13376
rect 2593 13345 2605 13348
rect 2639 13345 2651 13379
rect 2593 13339 2651 13345
rect 2866 13336 2872 13388
rect 2924 13336 2930 13388
rect 3145 13379 3203 13385
rect 3145 13345 3157 13379
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 2056 13240 2084 13336
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13308 2375 13311
rect 2884 13308 2912 13336
rect 2363 13280 2912 13308
rect 2363 13277 2375 13280
rect 2317 13271 2375 13277
rect 2409 13243 2467 13249
rect 2409 13240 2421 13243
rect 2056 13212 2421 13240
rect 2409 13209 2421 13212
rect 2455 13209 2467 13243
rect 3160 13240 3188 13339
rect 3234 13336 3240 13388
rect 3292 13336 3298 13388
rect 3436 13385 3464 13484
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 4120 13484 4292 13512
rect 4120 13472 4126 13484
rect 3694 13404 3700 13456
rect 3752 13444 3758 13456
rect 4154 13444 4160 13456
rect 3752 13416 4016 13444
rect 3752 13404 3758 13416
rect 3421 13379 3479 13385
rect 3421 13345 3433 13379
rect 3467 13345 3479 13379
rect 3421 13339 3479 13345
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13345 3571 13379
rect 3513 13339 3571 13345
rect 3605 13379 3663 13385
rect 3605 13345 3617 13379
rect 3651 13345 3663 13379
rect 3605 13339 3663 13345
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 3528 13308 3556 13339
rect 3384 13280 3556 13308
rect 3620 13308 3648 13339
rect 3786 13336 3792 13388
rect 3844 13336 3850 13388
rect 3988 13385 4016 13416
rect 4080 13416 4160 13444
rect 4080 13385 4108 13416
rect 4154 13404 4160 13416
rect 4212 13404 4218 13456
rect 4264 13453 4292 13484
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 4890 13512 4896 13524
rect 4580 13484 4896 13512
rect 4580 13472 4586 13484
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 6089 13515 6147 13521
rect 6089 13481 6101 13515
rect 6135 13512 6147 13515
rect 7926 13512 7932 13524
rect 6135 13484 7932 13512
rect 6135 13481 6147 13484
rect 6089 13475 6147 13481
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 9214 13512 9220 13524
rect 8404 13484 9220 13512
rect 4249 13447 4307 13453
rect 4249 13413 4261 13447
rect 4295 13413 4307 13447
rect 7006 13444 7012 13456
rect 4249 13407 4307 13413
rect 5000 13416 7012 13444
rect 3973 13379 4031 13385
rect 3973 13345 3985 13379
rect 4019 13345 4031 13379
rect 3973 13339 4031 13345
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13345 4123 13379
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 4065 13339 4123 13345
rect 4172 13348 4445 13376
rect 3988 13308 4016 13339
rect 4172 13320 4200 13348
rect 4433 13345 4445 13348
rect 4479 13345 4491 13379
rect 4433 13339 4491 13345
rect 4614 13336 4620 13388
rect 4672 13336 4678 13388
rect 4890 13336 4896 13388
rect 4948 13336 4954 13388
rect 4154 13308 4160 13320
rect 3620 13280 3832 13308
rect 3988 13280 4160 13308
rect 3384 13268 3390 13280
rect 3804 13240 3832 13280
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 5000 13308 5028 13416
rect 7006 13404 7012 13416
rect 7064 13404 7070 13456
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13376 5135 13379
rect 6362 13376 6368 13388
rect 5123 13348 6368 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 4396 13280 5028 13308
rect 4396 13268 4402 13280
rect 3160 13212 3832 13240
rect 2409 13203 2467 13209
rect 2774 13132 2780 13184
rect 2832 13132 2838 13184
rect 2958 13132 2964 13184
rect 3016 13132 3022 13184
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 3697 13175 3755 13181
rect 3697 13172 3709 13175
rect 3384 13144 3709 13172
rect 3384 13132 3390 13144
rect 3697 13141 3709 13144
rect 3743 13141 3755 13175
rect 3804 13172 3832 13212
rect 3878 13200 3884 13252
rect 3936 13240 3942 13252
rect 4249 13243 4307 13249
rect 4249 13240 4261 13243
rect 3936 13212 4261 13240
rect 3936 13200 3942 13212
rect 4249 13209 4261 13212
rect 4295 13209 4307 13243
rect 5092 13240 5120 13339
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 6546 13336 6552 13388
rect 6604 13376 6610 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 6604 13348 6745 13376
rect 6604 13336 6610 13348
rect 6733 13345 6745 13348
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 7561 13379 7619 13385
rect 7561 13376 7573 13379
rect 6972 13348 7573 13376
rect 6972 13336 6978 13348
rect 7561 13345 7573 13348
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 7926 13336 7932 13388
rect 7984 13336 7990 13388
rect 8110 13336 8116 13388
rect 8168 13336 8174 13388
rect 8404 13385 8432 13484
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 8665 13447 8723 13453
rect 8665 13413 8677 13447
rect 8711 13444 8723 13447
rect 9582 13444 9588 13456
rect 8711 13416 9588 13444
rect 8711 13413 8723 13416
rect 8665 13407 8723 13413
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 8478 13336 8484 13388
rect 8536 13336 8542 13388
rect 9401 13379 9459 13385
rect 9401 13345 9413 13379
rect 9447 13376 9459 13379
rect 9858 13376 9864 13388
rect 9447 13348 9864 13376
rect 9447 13345 9459 13348
rect 9401 13339 9459 13345
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 6822 13268 6828 13320
rect 6880 13268 6886 13320
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 8128 13308 8156 13336
rect 7064 13280 8156 13308
rect 7064 13268 7070 13280
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9582 13308 9588 13320
rect 9272 13280 9588 13308
rect 9272 13268 9278 13280
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 4249 13203 4307 13209
rect 4356 13212 5120 13240
rect 6840 13240 6868 13268
rect 7282 13240 7288 13252
rect 6840 13212 7288 13240
rect 4356 13172 4384 13212
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 3804 13144 4384 13172
rect 4801 13175 4859 13181
rect 3697 13135 3755 13141
rect 4801 13141 4813 13175
rect 4847 13172 4859 13175
rect 4890 13172 4896 13184
rect 4847 13144 4896 13172
rect 4847 13141 4859 13144
rect 4801 13135 4859 13141
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 4982 13132 4988 13184
rect 5040 13132 5046 13184
rect 7650 13132 7656 13184
rect 7708 13132 7714 13184
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8665 13175 8723 13181
rect 8665 13172 8677 13175
rect 8076 13144 8677 13172
rect 8076 13132 8082 13144
rect 8665 13141 8677 13144
rect 8711 13141 8723 13175
rect 8665 13135 8723 13141
rect 9217 13175 9275 13181
rect 9217 13141 9229 13175
rect 9263 13172 9275 13175
rect 9490 13172 9496 13184
rect 9263 13144 9496 13172
rect 9263 13141 9275 13144
rect 9217 13135 9275 13141
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 552 13082 11132 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 10062 13082
rect 10114 13030 10126 13082
rect 10178 13030 10190 13082
rect 10242 13030 10254 13082
rect 10306 13030 10318 13082
rect 10370 13030 11132 13082
rect 552 13008 11132 13030
rect 2590 12968 2596 12980
rect 1872 12940 2596 12968
rect 1872 12900 1900 12940
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 3053 12971 3111 12977
rect 3053 12937 3065 12971
rect 3099 12968 3111 12971
rect 3142 12968 3148 12980
rect 3099 12940 3148 12968
rect 3099 12937 3111 12940
rect 3053 12931 3111 12937
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 3697 12971 3755 12977
rect 3697 12968 3709 12971
rect 3568 12940 3709 12968
rect 3568 12928 3574 12940
rect 3697 12937 3709 12940
rect 3743 12937 3755 12971
rect 3697 12931 3755 12937
rect 9122 12928 9128 12980
rect 9180 12928 9186 12980
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 10008 12940 10333 12968
rect 10008 12928 10014 12940
rect 10321 12937 10333 12940
rect 10367 12937 10379 12971
rect 10321 12931 10379 12937
rect 1228 12872 1900 12900
rect 14 12724 20 12776
rect 72 12764 78 12776
rect 1228 12773 1256 12872
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 5261 12903 5319 12909
rect 5261 12900 5273 12903
rect 4672 12872 5273 12900
rect 4672 12860 4678 12872
rect 5261 12869 5273 12872
rect 5307 12869 5319 12903
rect 5261 12863 5319 12869
rect 2038 12792 2044 12844
rect 2096 12792 2102 12844
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 1213 12767 1271 12773
rect 1213 12764 1225 12767
rect 72 12736 1225 12764
rect 72 12724 78 12736
rect 1213 12733 1225 12736
rect 1259 12733 1271 12767
rect 1213 12727 1271 12733
rect 1302 12724 1308 12776
rect 1360 12764 1366 12776
rect 1673 12767 1731 12773
rect 1673 12764 1685 12767
rect 1360 12736 1685 12764
rect 1360 12724 1366 12736
rect 1673 12733 1685 12736
rect 1719 12764 1731 12767
rect 2222 12764 2228 12776
rect 1719 12736 2228 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 2516 12764 2544 12795
rect 2774 12792 2780 12844
rect 2832 12832 2838 12844
rect 3881 12835 3939 12841
rect 2832 12804 3556 12832
rect 2832 12792 2838 12804
rect 2516 12736 2820 12764
rect 2682 12656 2688 12708
rect 2740 12656 2746 12708
rect 2406 12588 2412 12640
rect 2464 12628 2470 12640
rect 2593 12631 2651 12637
rect 2593 12628 2605 12631
rect 2464 12600 2605 12628
rect 2464 12588 2470 12600
rect 2593 12597 2605 12600
rect 2639 12597 2651 12631
rect 2792 12628 2820 12736
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3528 12773 3556 12804
rect 3881 12801 3893 12835
rect 3927 12832 3939 12835
rect 4154 12832 4160 12844
rect 3927 12804 4160 12832
rect 3927 12801 3939 12804
rect 3881 12795 3939 12801
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 4706 12792 4712 12844
rect 4764 12792 4770 12844
rect 5276 12832 5304 12863
rect 5350 12860 5356 12912
rect 5408 12900 5414 12912
rect 8662 12900 8668 12912
rect 5408 12872 8668 12900
rect 5408 12860 5414 12872
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 8941 12903 8999 12909
rect 8941 12869 8953 12903
rect 8987 12900 8999 12903
rect 9306 12900 9312 12912
rect 8987 12872 9312 12900
rect 8987 12869 8999 12872
rect 8941 12863 8999 12869
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 5276 12804 7328 12832
rect 3237 12767 3295 12773
rect 3237 12764 3249 12767
rect 3200 12736 3249 12764
rect 3200 12724 3206 12736
rect 3237 12733 3249 12736
rect 3283 12733 3295 12767
rect 3237 12727 3295 12733
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12733 3571 12767
rect 4522 12764 4528 12776
rect 3513 12727 3571 12733
rect 4172 12736 4528 12764
rect 4172 12708 4200 12736
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 5442 12764 5448 12776
rect 5092 12736 5448 12764
rect 5092 12708 5120 12736
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5994 12724 6000 12776
rect 6052 12724 6058 12776
rect 6086 12724 6092 12776
rect 6144 12724 6150 12776
rect 6178 12724 6184 12776
rect 6236 12764 6242 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6236 12736 6653 12764
rect 6236 12724 6242 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 2866 12656 2872 12708
rect 2924 12696 2930 12708
rect 3694 12696 3700 12708
rect 2924 12668 3700 12696
rect 2924 12656 2930 12668
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 4154 12656 4160 12708
rect 4212 12656 4218 12708
rect 5074 12656 5080 12708
rect 5132 12656 5138 12708
rect 5718 12656 5724 12708
rect 5776 12696 5782 12708
rect 6104 12696 6132 12724
rect 5776 12668 6132 12696
rect 6656 12696 6684 12727
rect 6932 12696 6960 12727
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 7064 12736 7113 12764
rect 7064 12724 7070 12736
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 6656 12668 6960 12696
rect 5776 12656 5782 12668
rect 7190 12656 7196 12708
rect 7248 12656 7254 12708
rect 7300 12705 7328 12804
rect 8018 12792 8024 12844
rect 8076 12832 8082 12844
rect 8481 12835 8539 12841
rect 8481 12832 8493 12835
rect 8076 12804 8493 12832
rect 8076 12792 8082 12804
rect 8481 12801 8493 12804
rect 8527 12801 8539 12835
rect 8680 12832 8708 12860
rect 9493 12835 9551 12841
rect 9493 12832 9505 12835
rect 8680 12804 9505 12832
rect 8481 12795 8539 12801
rect 9493 12801 9505 12804
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 9674 12832 9680 12844
rect 9631 12804 9680 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12764 7619 12767
rect 7650 12764 7656 12776
rect 7607 12736 7656 12764
rect 7607 12733 7619 12736
rect 7561 12727 7619 12733
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 7742 12724 7748 12776
rect 7800 12724 7806 12776
rect 7834 12724 7840 12776
rect 7892 12724 7898 12776
rect 7926 12724 7932 12776
rect 7984 12724 7990 12776
rect 8110 12724 8116 12776
rect 8168 12724 8174 12776
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 7285 12699 7343 12705
rect 7285 12665 7297 12699
rect 7331 12696 7343 12699
rect 8021 12699 8079 12705
rect 7331 12668 7880 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 7852 12640 7880 12668
rect 8021 12665 8033 12699
rect 8067 12696 8079 12699
rect 8588 12696 8616 12727
rect 9306 12724 9312 12776
rect 9364 12724 9370 12776
rect 9398 12724 9404 12776
rect 9456 12724 9462 12776
rect 9508 12764 9536 12795
rect 9674 12792 9680 12804
rect 9732 12832 9738 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9732 12804 9873 12832
rect 9732 12792 9738 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12832 10103 12835
rect 10505 12835 10563 12841
rect 10505 12832 10517 12835
rect 10091 12804 10517 12832
rect 10091 12801 10103 12804
rect 10045 12795 10103 12801
rect 10505 12801 10517 12804
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 9953 12767 10011 12773
rect 9953 12764 9965 12767
rect 9508 12736 9965 12764
rect 9953 12733 9965 12736
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 10134 12724 10140 12776
rect 10192 12724 10198 12776
rect 10410 12724 10416 12776
rect 10468 12724 10474 12776
rect 10594 12724 10600 12776
rect 10652 12724 10658 12776
rect 8067 12668 8616 12696
rect 8067 12665 8079 12668
rect 8021 12659 8079 12665
rect 9674 12656 9680 12708
rect 9732 12696 9738 12708
rect 10318 12696 10324 12708
rect 9732 12668 10324 12696
rect 9732 12656 9738 12668
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 3329 12631 3387 12637
rect 3329 12628 3341 12631
rect 2792 12600 3341 12628
rect 2593 12591 2651 12597
rect 3329 12597 3341 12600
rect 3375 12628 3387 12631
rect 3418 12628 3424 12640
rect 3375 12600 3424 12628
rect 3375 12597 3387 12600
rect 3329 12591 3387 12597
rect 3418 12588 3424 12600
rect 3476 12628 3482 12640
rect 3786 12628 3792 12640
rect 3476 12600 3792 12628
rect 3476 12588 3482 12600
rect 3786 12588 3792 12600
rect 3844 12588 3850 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7377 12631 7435 12637
rect 7377 12628 7389 12631
rect 7156 12600 7389 12628
rect 7156 12588 7162 12600
rect 7377 12597 7389 12600
rect 7423 12597 7435 12631
rect 7377 12591 7435 12597
rect 7466 12588 7472 12640
rect 7524 12628 7530 12640
rect 7650 12628 7656 12640
rect 7524 12600 7656 12628
rect 7524 12588 7530 12600
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 7834 12588 7840 12640
rect 7892 12588 7898 12640
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 9490 12628 9496 12640
rect 8536 12600 9496 12628
rect 8536 12588 8542 12600
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 552 12538 11132 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 10722 12538
rect 10774 12486 10786 12538
rect 10838 12486 10850 12538
rect 10902 12486 10914 12538
rect 10966 12486 10978 12538
rect 11030 12486 11132 12538
rect 552 12464 11132 12486
rect 1578 12384 1584 12436
rect 1636 12424 1642 12436
rect 1636 12396 2452 12424
rect 1636 12384 1642 12396
rect 2222 12316 2228 12368
rect 2280 12316 2286 12368
rect 1581 12291 1639 12297
rect 1581 12257 1593 12291
rect 1627 12288 1639 12291
rect 1670 12288 1676 12300
rect 1627 12260 1676 12288
rect 1627 12257 1639 12260
rect 1581 12251 1639 12257
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 1762 12248 1768 12300
rect 1820 12288 1826 12300
rect 2424 12297 2452 12396
rect 2682 12384 2688 12436
rect 2740 12384 2746 12436
rect 2869 12427 2927 12433
rect 2869 12393 2881 12427
rect 2915 12424 2927 12427
rect 3050 12424 3056 12436
rect 2915 12396 3056 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 4062 12384 4068 12436
rect 4120 12384 4126 12436
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4982 12424 4988 12436
rect 4295 12396 4988 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4982 12384 4988 12396
rect 5040 12384 5046 12436
rect 5350 12384 5356 12436
rect 5408 12384 5414 12436
rect 6549 12427 6607 12433
rect 6104 12396 6408 12424
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 3421 12359 3479 12365
rect 3421 12356 3433 12359
rect 2556 12328 3433 12356
rect 2556 12316 2562 12328
rect 3421 12325 3433 12328
rect 3467 12325 3479 12359
rect 4801 12359 4859 12365
rect 4801 12356 4813 12359
rect 3421 12319 3479 12325
rect 4261 12328 4813 12356
rect 1949 12291 2007 12297
rect 1949 12288 1961 12291
rect 1820 12260 1961 12288
rect 1820 12248 1826 12260
rect 1949 12257 1961 12260
rect 1995 12257 2007 12291
rect 1949 12251 2007 12257
rect 2409 12291 2467 12297
rect 2409 12257 2421 12291
rect 2455 12288 2467 12291
rect 2682 12288 2688 12300
rect 2455 12260 2688 12288
rect 2455 12257 2467 12260
rect 2409 12251 2467 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 2866 12291 2924 12297
rect 2866 12288 2878 12291
rect 2832 12260 2878 12288
rect 2832 12248 2838 12260
rect 2866 12257 2878 12260
rect 2912 12288 2924 12291
rect 3605 12291 3663 12297
rect 3605 12288 3617 12291
rect 2912 12260 3617 12288
rect 2912 12257 2924 12260
rect 2866 12251 2924 12257
rect 3605 12257 3617 12260
rect 3651 12257 3663 12291
rect 3605 12251 3663 12257
rect 3786 12248 3792 12300
rect 3844 12248 3850 12300
rect 3881 12291 3939 12297
rect 3881 12257 3893 12291
rect 3927 12288 3939 12291
rect 4062 12288 4068 12300
rect 3927 12260 4068 12288
rect 3927 12257 3939 12260
rect 3881 12251 3939 12257
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4261 12297 4289 12328
rect 4801 12325 4813 12328
rect 4847 12356 4859 12359
rect 4890 12356 4896 12368
rect 4847 12328 4896 12356
rect 4847 12325 4859 12328
rect 4801 12319 4859 12325
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 5368 12356 5396 12384
rect 5000 12328 5396 12356
rect 5000 12297 5028 12328
rect 5534 12316 5540 12368
rect 5592 12356 5598 12368
rect 6104 12365 6132 12396
rect 6089 12359 6147 12365
rect 6089 12356 6101 12359
rect 5592 12328 6101 12356
rect 5592 12316 5598 12328
rect 6089 12325 6101 12328
rect 6135 12325 6147 12359
rect 6380 12356 6408 12396
rect 6549 12393 6561 12427
rect 6595 12424 6607 12427
rect 6730 12424 6736 12436
rect 6595 12396 6736 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 8478 12424 8484 12436
rect 7484 12396 8484 12424
rect 7190 12356 7196 12368
rect 6380 12328 7196 12356
rect 6089 12319 6147 12325
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 4246 12291 4304 12297
rect 4246 12257 4258 12291
rect 4292 12257 4304 12291
rect 4985 12291 5043 12297
rect 4985 12288 4997 12291
rect 4246 12251 4304 12257
rect 4356 12260 4997 12288
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 2958 12220 2964 12232
rect 2271 12192 2964 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 3326 12180 3332 12232
rect 3384 12180 3390 12232
rect 3804 12220 3832 12248
rect 4356 12220 4384 12260
rect 4985 12257 4997 12260
rect 5031 12257 5043 12291
rect 4985 12251 5043 12257
rect 5077 12291 5135 12297
rect 5077 12257 5089 12291
rect 5123 12257 5135 12291
rect 5077 12251 5135 12257
rect 3804 12192 4384 12220
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 4890 12220 4896 12232
rect 4755 12192 4896 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 1946 12112 1952 12164
rect 2004 12152 2010 12164
rect 2682 12152 2688 12164
rect 2004 12124 2688 12152
rect 2004 12112 2010 12124
rect 2682 12112 2688 12124
rect 2740 12112 2746 12164
rect 4798 12112 4804 12164
rect 4856 12112 4862 12164
rect 4982 12112 4988 12164
rect 5040 12152 5046 12164
rect 5092 12152 5120 12251
rect 5166 12248 5172 12300
rect 5224 12248 5230 12300
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 5445 12291 5503 12297
rect 5445 12288 5457 12291
rect 5408 12260 5457 12288
rect 5408 12248 5414 12260
rect 5445 12257 5457 12260
rect 5491 12257 5503 12291
rect 5445 12251 5503 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 6288 12220 6316 12251
rect 6362 12248 6368 12300
rect 6420 12248 6426 12300
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 7098 12288 7104 12300
rect 6779 12260 7104 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 7098 12248 7104 12260
rect 7156 12248 7162 12300
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12288 7343 12291
rect 7374 12288 7380 12300
rect 7331 12260 7380 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7484 12297 7512 12396
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 9493 12427 9551 12433
rect 9493 12424 9505 12427
rect 9364 12396 9505 12424
rect 9364 12384 9370 12396
rect 9493 12393 9505 12396
rect 9539 12393 9551 12427
rect 9493 12387 9551 12393
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10192 12396 10241 12424
rect 10192 12384 10198 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 7926 12356 7932 12368
rect 7760 12328 7932 12356
rect 7760 12297 7788 12328
rect 7926 12316 7932 12328
rect 7984 12356 7990 12368
rect 8297 12359 8355 12365
rect 8297 12356 8309 12359
rect 7984 12328 8309 12356
rect 7984 12316 7990 12328
rect 8297 12325 8309 12328
rect 8343 12325 8355 12359
rect 8849 12359 8907 12365
rect 8849 12356 8861 12359
rect 8297 12319 8355 12325
rect 8404 12328 8861 12356
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12257 7803 12291
rect 7745 12251 7803 12257
rect 8018 12248 8024 12300
rect 8076 12248 8082 12300
rect 8110 12248 8116 12300
rect 8168 12288 8174 12300
rect 8205 12291 8263 12297
rect 8205 12288 8217 12291
rect 8168 12260 8217 12288
rect 8168 12248 8174 12260
rect 8205 12257 8217 12260
rect 8251 12288 8263 12291
rect 8404 12288 8432 12328
rect 8849 12325 8861 12328
rect 8895 12325 8907 12359
rect 8849 12319 8907 12325
rect 10594 12316 10600 12368
rect 10652 12316 10658 12368
rect 8251 12260 8432 12288
rect 8251 12257 8263 12260
rect 8205 12251 8263 12257
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 8757 12291 8815 12297
rect 8757 12288 8769 12291
rect 8536 12260 8769 12288
rect 8536 12248 8542 12260
rect 8757 12257 8769 12260
rect 8803 12257 8815 12291
rect 8757 12251 8815 12257
rect 8941 12291 8999 12297
rect 8941 12257 8953 12291
rect 8987 12257 8999 12291
rect 8941 12251 8999 12257
rect 6454 12220 6460 12232
rect 6288 12192 6460 12220
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 7006 12180 7012 12232
rect 7064 12180 7070 12232
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 8956 12220 8984 12251
rect 9122 12248 9128 12300
rect 9180 12248 9186 12300
rect 9306 12248 9312 12300
rect 9364 12248 9370 12300
rect 9766 12248 9772 12300
rect 9824 12248 9830 12300
rect 10410 12248 10416 12300
rect 10468 12248 10474 12300
rect 9214 12220 9220 12232
rect 8956 12192 9220 12220
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12220 9919 12223
rect 10502 12220 10508 12232
rect 9907 12192 10508 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 5040 12124 5120 12152
rect 5169 12155 5227 12161
rect 5040 12112 5046 12124
rect 5169 12121 5181 12155
rect 5215 12152 5227 12155
rect 5258 12152 5264 12164
rect 5215 12124 5264 12152
rect 5215 12121 5227 12124
rect 5169 12115 5227 12121
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 6638 12112 6644 12164
rect 6696 12152 6702 12164
rect 7561 12155 7619 12161
rect 7561 12152 7573 12155
rect 6696 12124 7573 12152
rect 6696 12112 6702 12124
rect 7561 12121 7573 12124
rect 7607 12121 7619 12155
rect 7561 12115 7619 12121
rect 10137 12155 10195 12161
rect 10137 12121 10149 12155
rect 10183 12152 10195 12155
rect 10594 12152 10600 12164
rect 10183 12124 10600 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10594 12112 10600 12124
rect 10652 12112 10658 12164
rect 1397 12087 1455 12093
rect 1397 12053 1409 12087
rect 1443 12084 1455 12087
rect 1486 12084 1492 12096
rect 1443 12056 1492 12084
rect 1443 12053 1455 12056
rect 1397 12047 1455 12053
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 2038 12044 2044 12096
rect 2096 12044 2102 12096
rect 2314 12044 2320 12096
rect 2372 12084 2378 12096
rect 2501 12087 2559 12093
rect 2501 12084 2513 12087
rect 2372 12056 2513 12084
rect 2372 12044 2378 12056
rect 2501 12053 2513 12056
rect 2547 12053 2559 12087
rect 2501 12047 2559 12053
rect 3234 12044 3240 12096
rect 3292 12044 3298 12096
rect 4617 12087 4675 12093
rect 4617 12053 4629 12087
rect 4663 12084 4675 12087
rect 4706 12084 4712 12096
rect 4663 12056 4712 12084
rect 4663 12053 4675 12056
rect 4617 12047 4675 12053
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 6089 12087 6147 12093
rect 6089 12053 6101 12087
rect 6135 12084 6147 12087
rect 6178 12084 6184 12096
rect 6135 12056 6184 12084
rect 6135 12053 6147 12056
rect 6089 12047 6147 12053
rect 6178 12044 6184 12056
rect 6236 12044 6242 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6788 12056 6929 12084
rect 6788 12044 6794 12056
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 6917 12047 6975 12053
rect 7377 12087 7435 12093
rect 7377 12053 7389 12087
rect 7423 12084 7435 12087
rect 8110 12084 8116 12096
rect 7423 12056 8116 12084
rect 7423 12053 7435 12056
rect 7377 12047 7435 12053
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 552 11994 11132 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 10062 11994
rect 10114 11942 10126 11994
rect 10178 11942 10190 11994
rect 10242 11942 10254 11994
rect 10306 11942 10318 11994
rect 10370 11942 11132 11994
rect 552 11920 11132 11942
rect 2590 11840 2596 11892
rect 2648 11840 2654 11892
rect 3234 11840 3240 11892
rect 3292 11840 3298 11892
rect 3326 11840 3332 11892
rect 3384 11880 3390 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3384 11852 3801 11880
rect 3384 11840 3390 11852
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 5902 11840 5908 11892
rect 5960 11880 5966 11892
rect 6181 11883 6239 11889
rect 6181 11880 6193 11883
rect 5960 11852 6193 11880
rect 5960 11840 5966 11852
rect 6181 11849 6193 11852
rect 6227 11849 6239 11883
rect 6181 11843 6239 11849
rect 6730 11840 6736 11892
rect 6788 11840 6794 11892
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7285 11883 7343 11889
rect 7285 11880 7297 11883
rect 7064 11852 7297 11880
rect 7064 11840 7070 11852
rect 7285 11849 7297 11852
rect 7331 11849 7343 11883
rect 7285 11843 7343 11849
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 8849 11883 8907 11889
rect 8168 11852 8708 11880
rect 8168 11840 8174 11852
rect 7668 11784 8432 11812
rect 1394 11704 1400 11756
rect 1452 11744 1458 11756
rect 1452 11716 2084 11744
rect 1452 11704 1458 11716
rect 1578 11636 1584 11688
rect 1636 11636 1642 11688
rect 1946 11636 1952 11688
rect 2004 11636 2010 11688
rect 2056 11676 2084 11716
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 2372 11716 4844 11744
rect 2372 11704 2378 11716
rect 2498 11676 2504 11688
rect 2056 11648 2504 11676
rect 2498 11636 2504 11648
rect 2556 11676 2562 11688
rect 2593 11679 2651 11685
rect 2593 11676 2605 11679
rect 2556 11648 2605 11676
rect 2556 11636 2562 11648
rect 2593 11645 2605 11648
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 2774 11636 2780 11688
rect 2832 11636 2838 11688
rect 3436 11685 3464 11716
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11645 3479 11679
rect 3421 11639 3479 11645
rect 3510 11636 3516 11688
rect 3568 11676 3574 11688
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 3568 11648 3709 11676
rect 3568 11636 3574 11648
rect 3697 11645 3709 11648
rect 3743 11676 3755 11679
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3743 11648 3801 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 3789 11639 3847 11645
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11645 4031 11679
rect 3973 11639 4031 11645
rect 3988 11608 4016 11639
rect 4816 11620 4844 11716
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 5905 11679 5963 11685
rect 5905 11676 5917 11679
rect 5684 11648 5917 11676
rect 5684 11636 5690 11648
rect 5905 11645 5917 11648
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 6178 11636 6184 11688
rect 6236 11636 6242 11688
rect 6914 11636 6920 11688
rect 6972 11636 6978 11688
rect 7190 11636 7196 11688
rect 7248 11676 7254 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 7248 11648 7297 11676
rect 7248 11636 7254 11648
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 7466 11636 7472 11688
rect 7524 11636 7530 11688
rect 7668 11685 7696 11784
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 7852 11716 7941 11744
rect 7852 11685 7880 11716
rect 7929 11713 7941 11716
rect 7975 11744 7987 11747
rect 8018 11744 8024 11756
rect 7975 11716 8024 11744
rect 7975 11713 7987 11716
rect 7929 11707 7987 11713
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8404 11744 8432 11784
rect 8478 11744 8484 11756
rect 8220 11716 8340 11744
rect 8404 11716 8484 11744
rect 8220 11685 8248 11716
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11645 7711 11679
rect 7653 11639 7711 11645
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11645 7895 11679
rect 8186 11679 8248 11685
rect 8186 11676 8198 11679
rect 7837 11639 7895 11645
rect 8128 11648 8198 11676
rect 3620 11580 4016 11608
rect 3620 11552 3648 11580
rect 4798 11568 4804 11620
rect 4856 11608 4862 11620
rect 6932 11608 6960 11636
rect 4856 11580 6960 11608
rect 7101 11611 7159 11617
rect 4856 11568 4862 11580
rect 7101 11577 7113 11611
rect 7147 11608 7159 11611
rect 7484 11608 7512 11636
rect 7147 11580 7512 11608
rect 7745 11611 7803 11617
rect 7147 11577 7159 11580
rect 7101 11571 7159 11577
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 8128 11608 8156 11648
rect 8186 11645 8198 11648
rect 8232 11648 8248 11679
rect 8312 11676 8340 11716
rect 8478 11704 8484 11716
rect 8536 11704 8542 11756
rect 8680 11753 8708 11852
rect 8849 11849 8861 11883
rect 8895 11880 8907 11883
rect 9122 11880 9128 11892
rect 8895 11852 9128 11880
rect 8895 11849 8907 11852
rect 8849 11843 8907 11849
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 10229 11883 10287 11889
rect 10229 11849 10241 11883
rect 10275 11880 10287 11883
rect 10502 11880 10508 11892
rect 10275 11852 10508 11880
rect 10275 11849 10287 11852
rect 10229 11843 10287 11849
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8904 11716 9045 11744
rect 8904 11704 8910 11716
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 9033 11707 9091 11713
rect 9140 11716 9597 11744
rect 8573 11679 8631 11685
rect 8573 11676 8585 11679
rect 8312 11648 8585 11676
rect 8232 11645 8244 11648
rect 8186 11639 8244 11645
rect 8573 11645 8585 11648
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 9140 11608 9168 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 10134 11744 10140 11756
rect 9824 11716 10140 11744
rect 9824 11704 9830 11716
rect 10134 11704 10140 11716
rect 10192 11744 10198 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 10192 11716 10333 11744
rect 10192 11704 10198 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 9493 11679 9551 11685
rect 9493 11676 9505 11679
rect 9232 11648 9505 11676
rect 9232 11617 9260 11648
rect 9493 11645 9505 11648
rect 9539 11645 9551 11679
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 9493 11639 9551 11645
rect 9600 11648 9689 11676
rect 9600 11620 9628 11648
rect 9677 11645 9689 11648
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 10042 11636 10048 11688
rect 10100 11636 10106 11688
rect 10594 11636 10600 11688
rect 10652 11676 10658 11688
rect 11054 11676 11060 11688
rect 10652 11648 11060 11676
rect 10652 11636 10658 11648
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 7791 11580 8156 11608
rect 8312 11580 9168 11608
rect 9217 11611 9275 11617
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 1394 11500 1400 11552
rect 1452 11500 1458 11552
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 1765 11543 1823 11549
rect 1765 11540 1777 11543
rect 1636 11512 1777 11540
rect 1636 11500 1642 11512
rect 1765 11509 1777 11512
rect 1811 11509 1823 11543
rect 1765 11503 1823 11509
rect 3602 11500 3608 11552
rect 3660 11500 3666 11552
rect 5997 11543 6055 11549
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 6178 11540 6184 11552
rect 6043 11512 6184 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 7374 11500 7380 11552
rect 7432 11540 7438 11552
rect 7929 11543 7987 11549
rect 7929 11540 7941 11543
rect 7432 11512 7941 11540
rect 7432 11500 7438 11512
rect 7929 11509 7941 11512
rect 7975 11509 7987 11543
rect 7929 11503 7987 11509
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8312 11540 8340 11580
rect 9217 11577 9229 11611
rect 9263 11577 9275 11611
rect 9217 11571 9275 11577
rect 9401 11611 9459 11617
rect 9401 11577 9413 11611
rect 9447 11608 9459 11611
rect 9582 11608 9588 11620
rect 9447 11580 9588 11608
rect 9447 11577 9459 11580
rect 9401 11571 9459 11577
rect 8076 11512 8340 11540
rect 8076 11500 8082 11512
rect 8662 11500 8668 11552
rect 8720 11540 8726 11552
rect 9232 11540 9260 11571
rect 9582 11568 9588 11580
rect 9640 11608 9646 11620
rect 10413 11611 10471 11617
rect 10413 11608 10425 11611
rect 9640 11580 10425 11608
rect 9640 11568 9646 11580
rect 10413 11577 10425 11580
rect 10459 11577 10471 11611
rect 10413 11571 10471 11577
rect 8720 11512 9260 11540
rect 8720 11500 8726 11512
rect 9858 11500 9864 11552
rect 9916 11500 9922 11552
rect 10781 11543 10839 11549
rect 10781 11509 10793 11543
rect 10827 11540 10839 11543
rect 10827 11512 11192 11540
rect 10827 11509 10839 11512
rect 10781 11503 10839 11509
rect 552 11450 11132 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 10722 11450
rect 10774 11398 10786 11450
rect 10838 11398 10850 11450
rect 10902 11398 10914 11450
rect 10966 11398 10978 11450
rect 11030 11398 11132 11450
rect 552 11376 11132 11398
rect 1762 11296 1768 11348
rect 1820 11296 1826 11348
rect 2038 11296 2044 11348
rect 2096 11336 2102 11348
rect 3053 11339 3111 11345
rect 3053 11336 3065 11339
rect 2096 11308 3065 11336
rect 2096 11296 2102 11308
rect 3053 11305 3065 11308
rect 3099 11305 3111 11339
rect 3053 11299 3111 11305
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4246 11336 4252 11348
rect 4120 11308 4252 11336
rect 4120 11296 4126 11308
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 4706 11296 4712 11348
rect 4764 11296 4770 11348
rect 4890 11296 4896 11348
rect 4948 11296 4954 11348
rect 5810 11336 5816 11348
rect 5368 11308 5816 11336
rect 1946 11268 1952 11280
rect 1688 11240 1952 11268
rect 1688 11209 1716 11240
rect 1946 11228 1952 11240
rect 2004 11268 2010 11280
rect 2685 11271 2743 11277
rect 2685 11268 2697 11271
rect 2004 11240 2697 11268
rect 2004 11228 2010 11240
rect 2685 11237 2697 11240
rect 2731 11237 2743 11271
rect 2685 11231 2743 11237
rect 4264 11240 4844 11268
rect 4264 11212 4292 11240
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11169 1731 11203
rect 1673 11163 1731 11169
rect 1854 11160 1860 11212
rect 1912 11160 1918 11212
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11200 2191 11203
rect 2314 11200 2320 11212
rect 2179 11172 2320 11200
rect 2179 11169 2191 11172
rect 2133 11163 2191 11169
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 2593 11203 2651 11209
rect 2593 11200 2605 11203
rect 2424 11172 2605 11200
rect 2222 11092 2228 11144
rect 2280 11092 2286 11144
rect 1854 11024 1860 11076
rect 1912 11064 1918 11076
rect 2424 11064 2452 11172
rect 2593 11169 2605 11172
rect 2639 11169 2651 11203
rect 2593 11163 2651 11169
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11169 2927 11203
rect 2869 11163 2927 11169
rect 2884 11132 2912 11163
rect 3418 11160 3424 11212
rect 3476 11200 3482 11212
rect 3970 11200 3976 11212
rect 3476 11172 3976 11200
rect 3476 11160 3482 11172
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 4246 11160 4252 11212
rect 4304 11160 4310 11212
rect 4338 11160 4344 11212
rect 4396 11160 4402 11212
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 4706 11200 4712 11212
rect 4571 11172 4712 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 4816 11209 4844 11240
rect 4807 11203 4865 11209
rect 4807 11169 4819 11203
rect 4853 11169 4865 11203
rect 4807 11163 4865 11169
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 4356 11132 4384 11160
rect 5000 11132 5028 11163
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5368 11209 5396 11308
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 6178 11296 6184 11348
rect 6236 11296 6242 11348
rect 9398 11296 9404 11348
rect 9456 11296 9462 11348
rect 10042 11296 10048 11348
rect 10100 11296 10106 11348
rect 10134 11296 10140 11348
rect 10192 11296 10198 11348
rect 5445 11271 5503 11277
rect 5445 11237 5457 11271
rect 5491 11268 5503 11271
rect 5491 11240 5948 11268
rect 5491 11237 5503 11240
rect 5445 11231 5503 11237
rect 5920 11212 5948 11240
rect 8846 11228 8852 11280
rect 8904 11268 8910 11280
rect 9490 11268 9496 11280
rect 8904 11240 9496 11268
rect 8904 11228 8910 11240
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 10060 11268 10088 11296
rect 10060 11240 10180 11268
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 5316 11172 5365 11200
rect 5316 11160 5322 11172
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 5675 11172 5764 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5736 11132 5764 11172
rect 5810 11160 5816 11212
rect 5868 11160 5874 11212
rect 5902 11160 5908 11212
rect 5960 11200 5966 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5960 11172 6009 11200
rect 5960 11160 5966 11172
rect 5997 11169 6009 11172
rect 6043 11169 6055 11203
rect 5997 11163 6055 11169
rect 6454 11160 6460 11212
rect 6512 11200 6518 11212
rect 6549 11203 6607 11209
rect 6549 11200 6561 11203
rect 6512 11172 6561 11200
rect 6512 11160 6518 11172
rect 6549 11169 6561 11172
rect 6595 11169 6607 11203
rect 6549 11163 6607 11169
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 8665 11203 8723 11209
rect 8665 11200 8677 11203
rect 8628 11172 8677 11200
rect 8628 11160 8634 11172
rect 8665 11169 8677 11172
rect 8711 11169 8723 11203
rect 8665 11163 8723 11169
rect 8754 11160 8760 11212
rect 8812 11200 8818 11212
rect 8938 11200 8944 11212
rect 8812 11172 8944 11200
rect 8812 11160 8818 11172
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 9217 11203 9275 11209
rect 9217 11200 9229 11203
rect 9180 11172 9229 11200
rect 9180 11160 9186 11172
rect 9217 11169 9229 11172
rect 9263 11169 9275 11203
rect 9217 11163 9275 11169
rect 9398 11160 9404 11212
rect 9456 11160 9462 11212
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 10152 11209 10180 11240
rect 9861 11203 9919 11209
rect 9861 11200 9873 11203
rect 9640 11172 9873 11200
rect 9640 11160 9646 11172
rect 9861 11169 9873 11172
rect 9907 11169 9919 11203
rect 9861 11163 9919 11169
rect 10045 11203 10103 11209
rect 10045 11169 10057 11203
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 11164 11200 11192 11512
rect 10367 11172 11192 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 2884 11104 3740 11132
rect 4356 11104 5028 11132
rect 5092 11104 5764 11132
rect 1912 11036 2452 11064
rect 2501 11067 2559 11073
rect 1912 11024 1918 11036
rect 2501 11033 2513 11067
rect 2547 11064 2559 11067
rect 3602 11064 3608 11076
rect 2547 11036 3608 11064
rect 2547 11033 2559 11036
rect 2501 11027 2559 11033
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 3712 11064 3740 11104
rect 5092 11064 5120 11104
rect 3712 11036 5120 11064
rect 5626 11024 5632 11076
rect 5684 11024 5690 11076
rect 5736 11064 5764 11104
rect 6638 11092 6644 11144
rect 6696 11092 6702 11144
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 7190 11132 7196 11144
rect 6963 11104 7196 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 10060 11132 10088 11163
rect 10594 11132 10600 11144
rect 9824 11104 10600 11132
rect 9824 11092 9830 11104
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 7834 11064 7840 11076
rect 5736 11036 7840 11064
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 7926 11024 7932 11076
rect 7984 11064 7990 11076
rect 8481 11067 8539 11073
rect 8481 11064 8493 11067
rect 7984 11036 8493 11064
rect 7984 11024 7990 11036
rect 8481 11033 8493 11036
rect 8527 11033 8539 11067
rect 8481 11027 8539 11033
rect 552 10906 11132 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 10062 10906
rect 10114 10854 10126 10906
rect 10178 10854 10190 10906
rect 10242 10854 10254 10906
rect 10306 10854 10318 10906
rect 10370 10854 11132 10906
rect 552 10832 11132 10854
rect 1857 10795 1915 10801
rect 1857 10761 1869 10795
rect 1903 10792 1915 10795
rect 1946 10792 1952 10804
rect 1903 10764 1952 10792
rect 1903 10761 1915 10764
rect 1857 10755 1915 10761
rect 1946 10752 1952 10764
rect 2004 10752 2010 10804
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 2280 10764 2513 10792
rect 2280 10752 2286 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 2501 10755 2559 10761
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 6270 10792 6276 10804
rect 5500 10764 6276 10792
rect 5500 10752 5506 10764
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 6365 10795 6423 10801
rect 6365 10761 6377 10795
rect 6411 10792 6423 10795
rect 6638 10792 6644 10804
rect 6411 10764 6644 10792
rect 6411 10761 6423 10764
rect 6365 10755 6423 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 7561 10795 7619 10801
rect 7561 10792 7573 10795
rect 7524 10764 7573 10792
rect 7524 10752 7530 10764
rect 7561 10761 7573 10764
rect 7607 10761 7619 10795
rect 7561 10755 7619 10761
rect 3234 10684 3240 10736
rect 3292 10724 3298 10736
rect 4154 10724 4160 10736
rect 3292 10696 4160 10724
rect 3292 10684 3298 10696
rect 4154 10684 4160 10696
rect 4212 10684 4218 10736
rect 4249 10727 4307 10733
rect 4249 10693 4261 10727
rect 4295 10724 4307 10727
rect 4338 10724 4344 10736
rect 4295 10696 4344 10724
rect 4295 10693 4307 10696
rect 4249 10687 4307 10693
rect 4338 10684 4344 10696
rect 4396 10684 4402 10736
rect 4985 10727 5043 10733
rect 4985 10693 4997 10727
rect 5031 10693 5043 10727
rect 5718 10724 5724 10736
rect 4985 10687 5043 10693
rect 5276 10696 5724 10724
rect 1213 10659 1271 10665
rect 1213 10625 1225 10659
rect 1259 10656 1271 10659
rect 1765 10659 1823 10665
rect 1259 10628 1716 10656
rect 1259 10625 1271 10628
rect 1213 10619 1271 10625
rect 1118 10548 1124 10600
rect 1176 10548 1182 10600
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 1397 10591 1455 10597
rect 1397 10588 1409 10591
rect 1360 10560 1409 10588
rect 1360 10548 1366 10560
rect 1397 10557 1409 10560
rect 1443 10557 1455 10591
rect 1688 10588 1716 10628
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 1811 10628 2636 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 2041 10591 2099 10597
rect 2041 10588 2053 10591
rect 1688 10560 2053 10588
rect 1397 10551 1455 10557
rect 2041 10557 2053 10560
rect 2087 10557 2099 10591
rect 2041 10551 2099 10557
rect 1136 10452 1164 10548
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10489 1639 10523
rect 2056 10520 2084 10551
rect 2314 10548 2320 10600
rect 2372 10548 2378 10600
rect 2608 10597 2636 10628
rect 3970 10616 3976 10668
rect 4028 10616 4034 10668
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10557 2467 10591
rect 2409 10551 2467 10557
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10557 2651 10591
rect 2593 10551 2651 10557
rect 2424 10520 2452 10551
rect 3786 10548 3792 10600
rect 3844 10588 3850 10600
rect 3881 10591 3939 10597
rect 3881 10588 3893 10591
rect 3844 10560 3893 10588
rect 3844 10548 3850 10560
rect 3881 10557 3893 10560
rect 3927 10588 3939 10591
rect 5000 10588 5028 10687
rect 5276 10597 5304 10696
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10724 5871 10727
rect 6454 10724 6460 10736
rect 5859 10696 6460 10724
rect 5859 10693 5871 10696
rect 5813 10687 5871 10693
rect 6454 10684 6460 10696
rect 6512 10724 6518 10736
rect 6512 10696 6684 10724
rect 6512 10684 6518 10696
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10656 5595 10659
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 5583 10628 5764 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 3927 10560 5028 10588
rect 5261 10591 5319 10597
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 5442 10548 5448 10600
rect 5500 10548 5506 10600
rect 5626 10548 5632 10600
rect 5684 10548 5690 10600
rect 5736 10597 5764 10628
rect 5920 10628 6561 10656
rect 5920 10597 5948 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10557 6239 10591
rect 6181 10551 6239 10557
rect 6457 10591 6515 10597
rect 6457 10557 6469 10591
rect 6503 10588 6515 10591
rect 6656 10588 6684 10696
rect 7190 10684 7196 10736
rect 7248 10724 7254 10736
rect 7926 10724 7932 10736
rect 7248 10696 7932 10724
rect 7248 10684 7254 10696
rect 7926 10684 7932 10696
rect 7984 10684 7990 10736
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 6503 10560 6684 10588
rect 6831 10628 7849 10656
rect 6503 10557 6515 10560
rect 6457 10551 6515 10557
rect 2056 10492 2452 10520
rect 1581 10483 1639 10489
rect 1596 10452 1624 10483
rect 4706 10480 4712 10532
rect 4764 10520 4770 10532
rect 4985 10523 5043 10529
rect 4985 10520 4997 10523
rect 4764 10492 4997 10520
rect 4764 10480 4770 10492
rect 4985 10489 4997 10492
rect 5031 10489 5043 10523
rect 4985 10483 5043 10489
rect 5169 10523 5227 10529
rect 5169 10489 5181 10523
rect 5215 10520 5227 10523
rect 5460 10520 5488 10548
rect 5215 10492 5488 10520
rect 5736 10520 5764 10551
rect 6196 10520 6224 10551
rect 5736 10492 6224 10520
rect 5215 10489 5227 10492
rect 5169 10483 5227 10489
rect 6270 10480 6276 10532
rect 6328 10520 6334 10532
rect 6733 10523 6791 10529
rect 6733 10520 6745 10523
rect 6328 10492 6745 10520
rect 6328 10480 6334 10492
rect 6733 10489 6745 10492
rect 6779 10489 6791 10523
rect 6733 10483 6791 10489
rect 3326 10452 3332 10464
rect 1136 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 5997 10455 6055 10461
rect 5997 10452 6009 10455
rect 5500 10424 6009 10452
rect 5500 10412 5506 10424
rect 5997 10421 6009 10424
rect 6043 10421 6055 10455
rect 5997 10415 6055 10421
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 6831 10452 6859 10628
rect 6914 10548 6920 10600
rect 6972 10548 6978 10600
rect 7190 10548 7196 10600
rect 7248 10548 7254 10600
rect 7668 10597 7696 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 8260 10628 9168 10656
rect 8260 10616 8266 10628
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10588 7435 10591
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 7423 10560 7481 10588
rect 7423 10557 7435 10560
rect 7377 10551 7435 10557
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 7760 10520 7788 10551
rect 7926 10548 7932 10600
rect 7984 10548 7990 10600
rect 8846 10548 8852 10600
rect 8904 10588 8910 10600
rect 9140 10597 9168 10628
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 8904 10560 8953 10588
rect 8904 10548 8910 10560
rect 8941 10557 8953 10560
rect 8987 10557 8999 10591
rect 8941 10551 8999 10557
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9306 10588 9312 10600
rect 9171 10560 9312 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9306 10548 9312 10560
rect 9364 10588 9370 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 9364 10560 9597 10588
rect 9364 10548 9370 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 9766 10548 9772 10600
rect 9824 10548 9830 10600
rect 7064 10492 7788 10520
rect 7064 10480 7070 10492
rect 6420 10424 6859 10452
rect 6420 10412 6426 10424
rect 8938 10412 8944 10464
rect 8996 10412 9002 10464
rect 9769 10455 9827 10461
rect 9769 10421 9781 10455
rect 9815 10452 9827 10455
rect 10594 10452 10600 10464
rect 9815 10424 10600 10452
rect 9815 10421 9827 10424
rect 9769 10415 9827 10421
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 552 10362 11132 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 10722 10362
rect 10774 10310 10786 10362
rect 10838 10310 10850 10362
rect 10902 10310 10914 10362
rect 10966 10310 10978 10362
rect 11030 10310 11132 10362
rect 552 10288 11132 10310
rect 1302 10208 1308 10260
rect 1360 10248 1366 10260
rect 1762 10248 1768 10260
rect 1360 10220 1768 10248
rect 1360 10208 1366 10220
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 2314 10208 2320 10260
rect 2372 10248 2378 10260
rect 3329 10251 3387 10257
rect 3329 10248 3341 10251
rect 2372 10220 3341 10248
rect 2372 10208 2378 10220
rect 3329 10217 3341 10220
rect 3375 10217 3387 10251
rect 3329 10211 3387 10217
rect 5258 10208 5264 10260
rect 5316 10208 5322 10260
rect 5537 10251 5595 10257
rect 5537 10217 5549 10251
rect 5583 10248 5595 10251
rect 5583 10220 6500 10248
rect 5583 10217 5595 10220
rect 5537 10211 5595 10217
rect 3145 10183 3203 10189
rect 3145 10149 3157 10183
rect 3191 10180 3203 10183
rect 5353 10183 5411 10189
rect 3191 10152 4384 10180
rect 3191 10149 3203 10152
rect 3145 10143 3203 10149
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1857 10115 1915 10121
rect 1857 10112 1869 10115
rect 1443 10084 1869 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1857 10081 1869 10084
rect 1903 10081 1915 10115
rect 1857 10075 1915 10081
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 2682 10112 2688 10124
rect 2087 10084 2688 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 2866 10072 2872 10124
rect 2924 10112 2930 10124
rect 3528 10121 3556 10152
rect 3053 10115 3111 10121
rect 3053 10112 3065 10115
rect 2924 10084 3065 10112
rect 2924 10072 2930 10084
rect 3053 10081 3065 10084
rect 3099 10081 3111 10115
rect 3053 10075 3111 10081
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10081 3295 10115
rect 3237 10075 3295 10081
rect 3513 10115 3571 10121
rect 3513 10081 3525 10115
rect 3559 10081 3571 10115
rect 3513 10075 3571 10081
rect 1486 10004 1492 10056
rect 1544 10004 1550 10056
rect 2314 10004 2320 10056
rect 2372 10004 2378 10056
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 3252 10044 3280 10075
rect 3786 10072 3792 10124
rect 3844 10072 3850 10124
rect 3878 10072 3884 10124
rect 3936 10072 3942 10124
rect 4356 10121 4384 10152
rect 5353 10149 5365 10183
rect 5399 10180 5411 10183
rect 5994 10180 6000 10192
rect 5399 10152 6000 10180
rect 5399 10149 5411 10152
rect 5353 10143 5411 10149
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 4341 10115 4399 10121
rect 4341 10081 4353 10115
rect 4387 10081 4399 10115
rect 4341 10075 4399 10081
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 4080 10044 4108 10075
rect 4154 10044 4160 10056
rect 2832 10016 4160 10044
rect 2832 10004 2838 10016
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10044 4307 10047
rect 4540 10044 4568 10075
rect 4890 10072 4896 10124
rect 4948 10072 4954 10124
rect 5442 10112 5448 10124
rect 5000 10084 5448 10112
rect 5000 10056 5028 10084
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 5675 10084 6132 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 4295 10016 4568 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 4982 10004 4988 10056
rect 5040 10004 5046 10056
rect 3697 9979 3755 9985
rect 3697 9945 3709 9979
rect 3743 9976 3755 9979
rect 3970 9976 3976 9988
rect 3743 9948 3976 9976
rect 3743 9945 3755 9948
rect 3697 9939 3755 9945
rect 3970 9936 3976 9948
rect 4028 9976 4034 9988
rect 4433 9979 4491 9985
rect 4433 9976 4445 9979
rect 4028 9948 4445 9976
rect 4028 9936 4034 9948
rect 4433 9945 4445 9948
rect 4479 9945 4491 9979
rect 4433 9939 4491 9945
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 5353 9979 5411 9985
rect 5353 9976 5365 9979
rect 4764 9948 5365 9976
rect 4764 9936 4770 9948
rect 5353 9945 5365 9948
rect 5399 9945 5411 9979
rect 5353 9939 5411 9945
rect 1670 9868 1676 9920
rect 1728 9868 1734 9920
rect 2225 9911 2283 9917
rect 2225 9877 2237 9911
rect 2271 9908 2283 9911
rect 2590 9908 2596 9920
rect 2271 9880 2596 9908
rect 2271 9877 2283 9880
rect 2225 9871 2283 9877
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 5368 9908 5396 9939
rect 5902 9936 5908 9988
rect 5960 9976 5966 9988
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 5960 9948 6009 9976
rect 5960 9936 5966 9948
rect 5997 9945 6009 9948
rect 6043 9945 6055 9979
rect 6104 9976 6132 10084
rect 6178 10072 6184 10124
rect 6236 10072 6242 10124
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 6328 10084 6377 10112
rect 6328 10072 6334 10084
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 6472 10112 6500 10220
rect 7006 10208 7012 10260
rect 7064 10208 7070 10260
rect 7282 10208 7288 10260
rect 7340 10208 7346 10260
rect 9217 10251 9275 10257
rect 9217 10217 9229 10251
rect 9263 10248 9275 10251
rect 9398 10248 9404 10260
rect 9263 10220 9404 10248
rect 9263 10217 9275 10220
rect 9217 10211 9275 10217
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 10410 10208 10416 10260
rect 10468 10208 10474 10260
rect 7300 10180 7328 10208
rect 7469 10183 7527 10189
rect 7469 10180 7481 10183
rect 7300 10152 7481 10180
rect 7469 10149 7481 10152
rect 7515 10149 7527 10183
rect 7469 10143 7527 10149
rect 9490 10140 9496 10192
rect 9548 10180 9554 10192
rect 9548 10152 9628 10180
rect 9548 10140 9554 10152
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 6472 10084 6653 10112
rect 6365 10075 6423 10081
rect 6641 10081 6653 10084
rect 6687 10112 6699 10115
rect 6730 10112 6736 10124
rect 6687 10084 6736 10112
rect 6687 10081 6699 10084
rect 6641 10075 6699 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 6871 10084 7113 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 7248 10084 7297 10112
rect 7248 10072 7254 10084
rect 7285 10081 7297 10084
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 8846 10072 8852 10124
rect 8904 10072 8910 10124
rect 9600 10121 9628 10152
rect 10152 10152 10548 10180
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10081 9643 10115
rect 9585 10075 9643 10081
rect 8938 10004 8944 10056
rect 8996 10004 9002 10056
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10044 9551 10047
rect 9674 10044 9680 10056
rect 9539 10016 9680 10044
rect 9539 10013 9551 10016
rect 9493 10007 9551 10013
rect 6362 9976 6368 9988
rect 6104 9948 6368 9976
rect 5997 9939 6055 9945
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 8662 9936 8668 9988
rect 8720 9976 8726 9988
rect 9508 9976 9536 10007
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 10045 10047 10103 10053
rect 10045 10044 10057 10047
rect 9824 10016 10057 10044
rect 9824 10004 9830 10016
rect 10045 10013 10057 10016
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 8720 9948 9536 9976
rect 8720 9936 8726 9948
rect 9950 9936 9956 9988
rect 10008 9976 10014 9988
rect 10152 9976 10180 10152
rect 10520 10121 10548 10152
rect 10594 10140 10600 10192
rect 10652 10140 10658 10192
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10081 10563 10115
rect 10612 10112 10640 10140
rect 10689 10115 10747 10121
rect 10689 10112 10701 10115
rect 10612 10084 10701 10112
rect 10505 10075 10563 10081
rect 10689 10081 10701 10084
rect 10735 10081 10747 10115
rect 10689 10075 10747 10081
rect 10244 10044 10272 10075
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 10244 10016 10609 10044
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 10008 9948 10180 9976
rect 10008 9936 10014 9948
rect 6178 9908 6184 9920
rect 5368 9880 6184 9908
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 552 9818 11132 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 10062 9818
rect 10114 9766 10126 9818
rect 10178 9766 10190 9818
rect 10242 9766 10254 9818
rect 10306 9766 10318 9818
rect 10370 9766 11132 9818
rect 552 9744 11132 9766
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 5169 9707 5227 9713
rect 5169 9704 5181 9707
rect 4948 9676 5181 9704
rect 4948 9664 4954 9676
rect 5169 9673 5181 9676
rect 5215 9673 5227 9707
rect 5169 9667 5227 9673
rect 6181 9707 6239 9713
rect 6181 9673 6193 9707
rect 6227 9704 6239 9707
rect 6270 9704 6276 9716
rect 6227 9676 6276 9704
rect 6227 9673 6239 9676
rect 6181 9667 6239 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6362 9664 6368 9716
rect 6420 9664 6426 9716
rect 6730 9664 6736 9716
rect 6788 9664 6794 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 8941 9707 8999 9713
rect 8941 9704 8953 9707
rect 8904 9676 8953 9704
rect 8904 9664 8910 9676
rect 8941 9673 8953 9676
rect 8987 9673 8999 9707
rect 8941 9667 8999 9673
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 1949 9639 2007 9645
rect 1949 9636 1961 9639
rect 1912 9608 1961 9636
rect 1912 9596 1918 9608
rect 1949 9605 1961 9608
rect 1995 9605 2007 9639
rect 1949 9599 2007 9605
rect 2593 9639 2651 9645
rect 2593 9605 2605 9639
rect 2639 9636 2651 9639
rect 3510 9636 3516 9648
rect 2639 9608 3516 9636
rect 2639 9605 2651 9608
rect 2593 9599 2651 9605
rect 3510 9596 3516 9608
rect 3568 9596 3574 9648
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 4341 9639 4399 9645
rect 4341 9636 4353 9639
rect 4304 9608 4353 9636
rect 4304 9596 4310 9608
rect 4341 9605 4353 9608
rect 4387 9605 4399 9639
rect 4341 9599 4399 9605
rect 5074 9596 5080 9648
rect 5132 9636 5138 9648
rect 5350 9636 5356 9648
rect 5132 9608 5356 9636
rect 5132 9596 5138 9608
rect 5350 9596 5356 9608
rect 5408 9596 5414 9648
rect 5994 9596 6000 9648
rect 6052 9596 6058 9648
rect 1670 9528 1676 9580
rect 1728 9528 1734 9580
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4632 9540 5396 9568
rect 1302 9460 1308 9512
rect 1360 9500 1366 9512
rect 1581 9503 1639 9509
rect 1581 9500 1593 9503
rect 1360 9472 1593 9500
rect 1360 9460 1366 9472
rect 1581 9469 1593 9472
rect 1627 9469 1639 9503
rect 1581 9463 1639 9469
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9469 2283 9503
rect 2332 9500 2360 9531
rect 2590 9500 2596 9512
rect 2332 9472 2596 9500
rect 2225 9463 2283 9469
rect 2240 9432 2268 9463
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 2682 9460 2688 9512
rect 2740 9460 2746 9512
rect 2866 9460 2872 9512
rect 2924 9460 2930 9512
rect 3970 9460 3976 9512
rect 4028 9460 4034 9512
rect 4080 9500 4108 9531
rect 4632 9509 4660 9540
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4080 9472 4445 9500
rect 2314 9432 2320 9444
rect 2240 9404 2320 9432
rect 2314 9392 2320 9404
rect 2372 9432 2378 9444
rect 2777 9435 2835 9441
rect 2777 9432 2789 9435
rect 2372 9404 2789 9432
rect 2372 9392 2378 9404
rect 2777 9401 2789 9404
rect 2823 9401 2835 9435
rect 2777 9395 2835 9401
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4080 9432 4108 9472
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9500 4675 9503
rect 4706 9500 4712 9512
rect 4663 9472 4712 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9500 4951 9503
rect 4982 9500 4988 9512
rect 4939 9472 4988 9500
rect 4939 9469 4951 9472
rect 4893 9463 4951 9469
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5368 9509 5396 9540
rect 5718 9528 5724 9580
rect 5776 9528 5782 9580
rect 7282 9568 7288 9580
rect 6656 9540 7288 9568
rect 6656 9512 6684 9540
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 8956 9568 8984 9667
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 9953 9707 10011 9713
rect 9953 9704 9965 9707
rect 9824 9676 9965 9704
rect 9824 9664 9830 9676
rect 9953 9673 9965 9676
rect 9999 9673 10011 9707
rect 9953 9667 10011 9673
rect 9490 9636 9496 9648
rect 9416 9608 9496 9636
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 8956 9540 9229 9568
rect 9217 9537 9229 9540
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 9416 9577 9444 9608
rect 9490 9596 9496 9608
rect 9548 9596 9554 9648
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 5132 9472 5181 9500
rect 5132 9460 5138 9472
rect 5169 9469 5181 9472
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 5500 9472 5641 9500
rect 5500 9460 5506 9472
rect 5629 9469 5641 9472
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 3936 9404 4108 9432
rect 3936 9392 3942 9404
rect 5644 9364 5672 9463
rect 6638 9460 6644 9512
rect 6696 9460 6702 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 7190 9500 7196 9512
rect 6871 9472 7196 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 7190 9460 7196 9472
rect 7248 9500 7254 9512
rect 8478 9500 8484 9512
rect 7248 9472 8484 9500
rect 7248 9460 7254 9472
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 8570 9460 8576 9512
rect 8628 9460 8634 9512
rect 9490 9460 9496 9512
rect 9548 9460 9554 9512
rect 9950 9460 9956 9512
rect 10008 9500 10014 9512
rect 10137 9503 10195 9509
rect 10137 9500 10149 9503
rect 10008 9472 10149 9500
rect 10008 9460 10014 9472
rect 10137 9469 10149 9472
rect 10183 9469 10195 9503
rect 10137 9463 10195 9469
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9500 10379 9503
rect 10594 9500 10600 9512
rect 10367 9472 10600 9500
rect 10367 9469 10379 9472
rect 10321 9463 10379 9469
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 5994 9392 6000 9444
rect 6052 9432 6058 9444
rect 6333 9435 6391 9441
rect 6333 9432 6345 9435
rect 6052 9404 6345 9432
rect 6052 9392 6058 9404
rect 6333 9401 6345 9404
rect 6379 9401 6391 9435
rect 6333 9395 6391 9401
rect 6549 9435 6607 9441
rect 6549 9401 6561 9435
rect 6595 9432 6607 9435
rect 6730 9432 6736 9444
rect 6595 9404 6736 9432
rect 6595 9401 6607 9404
rect 6549 9395 6607 9401
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 8588 9432 8616 9460
rect 10502 9432 10508 9444
rect 8588 9404 10508 9432
rect 10502 9392 10508 9404
rect 10560 9392 10566 9444
rect 7190 9364 7196 9376
rect 5644 9336 7196 9364
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 8938 9364 8944 9376
rect 7892 9336 8944 9364
rect 7892 9324 7898 9336
rect 8938 9324 8944 9336
rect 8996 9364 9002 9376
rect 9033 9367 9091 9373
rect 9033 9364 9045 9367
rect 8996 9336 9045 9364
rect 8996 9324 9002 9336
rect 9033 9333 9045 9336
rect 9079 9333 9091 9367
rect 9033 9327 9091 9333
rect 552 9274 11132 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 10722 9274
rect 10774 9222 10786 9274
rect 10838 9222 10850 9274
rect 10902 9222 10914 9274
rect 10966 9222 10978 9274
rect 11030 9222 11132 9274
rect 552 9200 11132 9222
rect 1302 9120 1308 9172
rect 1360 9120 1366 9172
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 2866 9160 2872 9172
rect 2363 9132 2872 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 3970 9120 3976 9172
rect 4028 9160 4034 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 4028 9132 4077 9160
rect 4028 9120 4034 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4154 9120 4160 9172
rect 4212 9120 4218 9172
rect 4706 9120 4712 9172
rect 4764 9120 4770 9172
rect 4893 9163 4951 9169
rect 4893 9129 4905 9163
rect 4939 9160 4951 9163
rect 5074 9160 5080 9172
rect 4939 9132 5080 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7650 9160 7656 9172
rect 7331 9132 7656 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9490 9160 9496 9172
rect 9171 9132 9496 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 2133 9095 2191 9101
rect 2133 9092 2145 9095
rect 1688 9064 2145 9092
rect 1688 9033 1716 9064
rect 2133 9061 2145 9064
rect 2179 9061 2191 9095
rect 2133 9055 2191 9061
rect 2501 9095 2559 9101
rect 2501 9061 2513 9095
rect 2547 9092 2559 9095
rect 2682 9092 2688 9104
rect 2547 9064 2688 9092
rect 2547 9061 2559 9064
rect 2501 9055 2559 9061
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 8993 1731 9027
rect 1673 8987 1731 8993
rect 1946 8984 1952 9036
rect 2004 8984 2010 9036
rect 2148 9024 2176 9055
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 3329 9095 3387 9101
rect 3329 9061 3341 9095
rect 3375 9092 3387 9095
rect 3375 9064 3740 9092
rect 3375 9061 3387 9064
rect 3329 9055 3387 9061
rect 2314 9024 2320 9036
rect 2148 8996 2320 9024
rect 2314 8984 2320 8996
rect 2372 9024 2378 9036
rect 2409 9027 2467 9033
rect 2409 9024 2421 9027
rect 2372 8996 2421 9024
rect 2372 8984 2378 8996
rect 2409 8993 2421 8996
rect 2455 8993 2467 9027
rect 2409 8987 2467 8993
rect 2593 9027 2651 9033
rect 2593 8993 2605 9027
rect 2639 8993 2651 9027
rect 2593 8987 2651 8993
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1394 8956 1400 8968
rect 992 8928 1400 8956
rect 992 8916 998 8928
rect 1394 8916 1400 8928
rect 1452 8956 1458 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1452 8928 1593 8956
rect 1452 8916 1458 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1964 8956 1992 8984
rect 2608 8956 2636 8987
rect 3234 8984 3240 9036
rect 3292 8984 3298 9036
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 9024 3479 9027
rect 3510 9024 3516 9036
rect 3467 8996 3516 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 1964 8928 2636 8956
rect 1581 8919 1639 8925
rect 3326 8916 3332 8968
rect 3384 8956 3390 8968
rect 3436 8956 3464 8987
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 3712 9033 3740 9064
rect 3697 9027 3755 9033
rect 3697 8993 3709 9027
rect 3743 8993 3755 9027
rect 3697 8987 3755 8993
rect 3384 8928 3464 8956
rect 3712 8956 3740 8987
rect 3878 8984 3884 9036
rect 3936 8984 3942 9036
rect 3988 9033 4016 9120
rect 4172 9092 4200 9120
rect 8294 9092 8300 9104
rect 4172 9064 4384 9092
rect 3973 9027 4031 9033
rect 3973 8993 3985 9027
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 4080 8956 4108 8987
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4356 9033 4384 9064
rect 4540 9064 5028 9092
rect 4540 9033 4568 9064
rect 5000 9033 5028 9064
rect 8266 9052 8300 9092
rect 8352 9092 8358 9104
rect 8352 9064 9066 9092
rect 8352 9052 8358 9064
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 4212 8996 4261 9024
rect 4212 8984 4218 8996
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 4525 9027 4583 9033
rect 4525 8993 4537 9027
rect 4571 8993 4583 9027
rect 4525 8987 4583 8993
rect 4801 9027 4859 9033
rect 4801 8993 4813 9027
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 5074 9024 5080 9036
rect 5031 8996 5080 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 3712 8928 4108 8956
rect 4356 8956 4384 8987
rect 4816 8956 4844 8987
rect 5074 8984 5080 8996
rect 5132 9024 5138 9036
rect 6086 9024 6092 9036
rect 5132 8996 6092 9024
rect 5132 8984 5138 8996
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 7469 9027 7527 9033
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 8266 9024 8294 9052
rect 7515 8996 8294 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 8662 8984 8668 9036
rect 8720 9024 8726 9036
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 8720 8996 8953 9024
rect 8720 8984 8726 8996
rect 8941 8993 8953 8996
rect 8987 8993 8999 9027
rect 9038 9024 9066 9064
rect 9214 9052 9220 9104
rect 9272 9052 9278 9104
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 9038 8996 9413 9024
rect 8941 8987 8999 8993
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 4356 8928 6132 8956
rect 3384 8916 3390 8928
rect 6104 8900 6132 8928
rect 7742 8916 7748 8968
rect 7800 8916 7806 8968
rect 8018 8916 8024 8968
rect 8076 8916 8082 8968
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 2590 8848 2596 8900
rect 2648 8888 2654 8900
rect 3513 8891 3571 8897
rect 3513 8888 3525 8891
rect 2648 8860 3525 8888
rect 2648 8848 2654 8860
rect 3513 8857 3525 8860
rect 3559 8857 3571 8891
rect 3513 8851 3571 8857
rect 6086 8848 6092 8900
rect 6144 8848 6150 8900
rect 8128 8888 8156 8919
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 8294 8916 8300 8968
rect 8352 8916 8358 8968
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8536 8928 8769 8956
rect 8536 8916 8542 8928
rect 8757 8925 8769 8928
rect 8803 8925 8815 8959
rect 8956 8956 8984 8987
rect 9490 8956 9496 8968
rect 8956 8928 9496 8956
rect 8757 8919 8815 8925
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8956 9735 8959
rect 10594 8956 10600 8968
rect 9723 8928 10600 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 8570 8888 8576 8900
rect 8128 8860 8576 8888
rect 8570 8848 8576 8860
rect 8628 8848 8634 8900
rect 7653 8823 7711 8829
rect 7653 8789 7665 8823
rect 7699 8820 7711 8823
rect 7837 8823 7895 8829
rect 7837 8820 7849 8823
rect 7699 8792 7849 8820
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 7837 8789 7849 8792
rect 7883 8789 7895 8823
rect 7837 8783 7895 8789
rect 7926 8780 7932 8832
rect 7984 8820 7990 8832
rect 8294 8820 8300 8832
rect 7984 8792 8300 8820
rect 7984 8780 7990 8792
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 9582 8780 9588 8832
rect 9640 8780 9646 8832
rect 552 8730 11132 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 10062 8730
rect 10114 8678 10126 8730
rect 10178 8678 10190 8730
rect 10242 8678 10254 8730
rect 10306 8678 10318 8730
rect 10370 8678 11132 8730
rect 552 8656 11132 8678
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 7800 8588 8401 8616
rect 7800 8576 7806 8588
rect 8389 8585 8401 8588
rect 8435 8585 8447 8619
rect 8389 8579 8447 8585
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 8849 8619 8907 8625
rect 8849 8616 8861 8619
rect 8628 8588 8861 8616
rect 8628 8576 8634 8588
rect 8849 8585 8861 8588
rect 8895 8585 8907 8619
rect 8849 8579 8907 8585
rect 9582 8576 9588 8628
rect 9640 8576 9646 8628
rect 10594 8576 10600 8628
rect 10652 8576 10658 8628
rect 2041 8551 2099 8557
rect 2041 8517 2053 8551
rect 2087 8548 2099 8551
rect 2130 8548 2136 8560
rect 2087 8520 2136 8548
rect 2087 8517 2099 8520
rect 2041 8511 2099 8517
rect 2130 8508 2136 8520
rect 2188 8508 2194 8560
rect 8018 8508 8024 8560
rect 8076 8548 8082 8560
rect 8205 8551 8263 8557
rect 8205 8548 8217 8551
rect 8076 8520 8217 8548
rect 8076 8508 8082 8520
rect 8205 8517 8217 8520
rect 8251 8517 8263 8551
rect 8205 8511 8263 8517
rect 1578 8440 1584 8492
rect 1636 8440 1642 8492
rect 7374 8440 7380 8492
rect 7432 8440 7438 8492
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 7699 8452 8156 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 3510 8372 3516 8424
rect 3568 8412 3574 8424
rect 7285 8415 7343 8421
rect 3568 8384 4016 8412
rect 3568 8372 3574 8384
rect 3988 8353 4016 8384
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7926 8412 7932 8424
rect 7331 8384 7932 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 3789 8347 3847 8353
rect 3789 8313 3801 8347
rect 3835 8313 3847 8347
rect 3789 8307 3847 8313
rect 3973 8347 4031 8353
rect 3973 8313 3985 8347
rect 4019 8344 4031 8347
rect 4154 8344 4160 8356
rect 4019 8316 4160 8344
rect 4019 8313 4031 8316
rect 3973 8307 4031 8313
rect 3234 8236 3240 8288
rect 3292 8276 3298 8288
rect 3510 8276 3516 8288
rect 3292 8248 3516 8276
rect 3292 8236 3298 8248
rect 3510 8236 3516 8248
rect 3568 8276 3574 8288
rect 3804 8276 3832 8307
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 7834 8304 7840 8356
rect 7892 8304 7898 8356
rect 8021 8347 8079 8353
rect 8021 8313 8033 8347
rect 8067 8313 8079 8347
rect 8128 8344 8156 8452
rect 8220 8412 8248 8511
rect 9398 8508 9404 8560
rect 9456 8548 9462 8560
rect 10410 8548 10416 8560
rect 9456 8520 10416 8548
rect 9456 8508 9462 8520
rect 10410 8508 10416 8520
rect 10468 8508 10474 8560
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 8846 8480 8852 8492
rect 8352 8452 8852 8480
rect 8352 8440 8358 8452
rect 8846 8440 8852 8452
rect 8904 8480 8910 8492
rect 10505 8483 10563 8489
rect 10505 8480 10517 8483
rect 8904 8452 9812 8480
rect 8904 8440 8910 8452
rect 8665 8415 8723 8421
rect 8665 8412 8677 8415
rect 8220 8384 8677 8412
rect 8665 8381 8677 8384
rect 8711 8381 8723 8415
rect 8665 8375 8723 8381
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8202 8344 8208 8356
rect 8128 8316 8208 8344
rect 8021 8307 8079 8313
rect 3568 8248 3832 8276
rect 8036 8276 8064 8307
rect 8202 8304 8208 8316
rect 8260 8344 8266 8356
rect 8389 8347 8447 8353
rect 8389 8344 8401 8347
rect 8260 8316 8401 8344
rect 8260 8304 8266 8316
rect 8389 8313 8401 8316
rect 8435 8313 8447 8347
rect 8389 8307 8447 8313
rect 8570 8304 8576 8356
rect 8628 8304 8634 8356
rect 8294 8276 8300 8288
rect 8036 8248 8300 8276
rect 3568 8236 3574 8248
rect 8294 8236 8300 8248
rect 8352 8276 8358 8288
rect 8772 8276 8800 8375
rect 8938 8372 8944 8424
rect 8996 8372 9002 8424
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 9398 8412 9404 8424
rect 9355 8384 9404 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 9490 8372 9496 8424
rect 9548 8372 9554 8424
rect 9784 8421 9812 8452
rect 9968 8452 10517 8480
rect 9968 8421 9996 8452
rect 10505 8449 10517 8452
rect 10551 8480 10563 8483
rect 10551 8452 10824 8480
rect 10551 8449 10563 8452
rect 10505 8443 10563 8449
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8381 10011 8415
rect 9953 8375 10011 8381
rect 10042 8372 10048 8424
rect 10100 8412 10106 8424
rect 10796 8421 10824 8452
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 10100 8384 10609 8412
rect 10100 8372 10106 8384
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8381 10839 8415
rect 10781 8375 10839 8381
rect 10134 8304 10140 8356
rect 10192 8304 10198 8356
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8313 10379 8347
rect 10321 8307 10379 8313
rect 8352 8248 8800 8276
rect 8352 8236 8358 8248
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9309 8279 9367 8285
rect 9309 8276 9321 8279
rect 9180 8248 9321 8276
rect 9180 8236 9186 8248
rect 9309 8245 9321 8248
rect 9355 8245 9367 8279
rect 9309 8239 9367 8245
rect 9398 8236 9404 8288
rect 9456 8276 9462 8288
rect 10336 8276 10364 8307
rect 9456 8248 10364 8276
rect 9456 8236 9462 8248
rect 552 8186 11132 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 10722 8186
rect 10774 8134 10786 8186
rect 10838 8134 10850 8186
rect 10902 8134 10914 8186
rect 10966 8134 10978 8186
rect 11030 8134 11132 8186
rect 552 8112 11132 8134
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2498 8072 2504 8084
rect 2188 8044 2504 8072
rect 2188 8032 2194 8044
rect 2498 8032 2504 8044
rect 2556 8072 2562 8084
rect 2593 8075 2651 8081
rect 2593 8072 2605 8075
rect 2556 8044 2605 8072
rect 2556 8032 2562 8044
rect 2593 8041 2605 8044
rect 2639 8041 2651 8075
rect 2593 8035 2651 8041
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 8386 8072 8392 8084
rect 6604 8044 8392 8072
rect 6604 8032 6610 8044
rect 8386 8032 8392 8044
rect 8444 8072 8450 8084
rect 9401 8075 9459 8081
rect 8444 8044 9352 8072
rect 8444 8032 8450 8044
rect 6273 8007 6331 8013
rect 6273 7973 6285 8007
rect 6319 8004 6331 8007
rect 7101 8007 7159 8013
rect 7101 8004 7113 8007
rect 6319 7976 7113 8004
rect 6319 7973 6331 7976
rect 6273 7967 6331 7973
rect 7101 7973 7113 7976
rect 7147 8004 7159 8007
rect 7147 7976 7880 8004
rect 7147 7973 7159 7976
rect 7101 7967 7159 7973
rect 1394 7896 1400 7948
rect 1452 7936 1458 7948
rect 1581 7939 1639 7945
rect 1581 7936 1593 7939
rect 1452 7908 1593 7936
rect 1452 7896 1458 7908
rect 1581 7905 1593 7908
rect 1627 7905 1639 7939
rect 1581 7899 1639 7905
rect 1596 7868 1624 7899
rect 1946 7896 1952 7948
rect 2004 7936 2010 7948
rect 3142 7936 3148 7948
rect 2004 7908 3148 7936
rect 2004 7896 2010 7908
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 6454 7896 6460 7948
rect 6512 7896 6518 7948
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 6604 7908 6653 7936
rect 6604 7896 6610 7908
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7936 7251 7939
rect 7374 7936 7380 7948
rect 7239 7908 7380 7936
rect 7239 7905 7251 7908
rect 7193 7899 7251 7905
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 7469 7899 7527 7905
rect 2498 7868 2504 7880
rect 1596 7840 2504 7868
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7484 7868 7512 7899
rect 7650 7896 7656 7948
rect 7708 7896 7714 7948
rect 7742 7896 7748 7948
rect 7800 7896 7806 7948
rect 7852 7936 7880 7976
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 8481 8007 8539 8013
rect 8481 8004 8493 8007
rect 7984 7976 8493 8004
rect 7984 7964 7990 7976
rect 8481 7973 8493 7976
rect 8527 7973 8539 8007
rect 8481 7967 8539 7973
rect 8757 8007 8815 8013
rect 8757 7973 8769 8007
rect 8803 8004 8815 8007
rect 9033 8007 9091 8013
rect 9033 8004 9045 8007
rect 8803 7976 9045 8004
rect 8803 7973 8815 7976
rect 8757 7967 8815 7973
rect 9033 7973 9045 7976
rect 9079 8004 9091 8007
rect 9122 8004 9128 8016
rect 9079 7976 9128 8004
rect 9079 7973 9091 7976
rect 9033 7967 9091 7973
rect 9122 7964 9128 7976
rect 9180 7964 9186 8016
rect 9233 8007 9291 8013
rect 9233 8004 9245 8007
rect 9232 7973 9245 8004
rect 9279 7973 9291 8007
rect 9324 8004 9352 8044
rect 9401 8041 9413 8075
rect 9447 8072 9459 8075
rect 10134 8072 10140 8084
rect 9447 8044 10140 8072
rect 9447 8041 9459 8044
rect 9401 8035 9459 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 9324 7976 10640 8004
rect 9232 7967 9291 7973
rect 7852 7908 8248 7936
rect 7558 7868 7564 7880
rect 6788 7840 7420 7868
rect 7484 7840 7564 7868
rect 6788 7828 6794 7840
rect 6914 7692 6920 7744
rect 6972 7692 6978 7744
rect 7282 7692 7288 7744
rect 7340 7692 7346 7744
rect 7392 7732 7420 7840
rect 7558 7828 7564 7840
rect 7616 7868 7622 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7616 7840 7849 7868
rect 7616 7828 7622 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 8113 7803 8171 7809
rect 8113 7800 8125 7803
rect 7708 7772 8125 7800
rect 7708 7760 7714 7772
rect 8113 7769 8125 7772
rect 8159 7769 8171 7803
rect 8220 7800 8248 7908
rect 8386 7896 8392 7948
rect 8444 7896 8450 7948
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7905 8631 7939
rect 8573 7899 8631 7905
rect 8665 7939 8723 7945
rect 8665 7905 8677 7939
rect 8711 7905 8723 7939
rect 8665 7899 8723 7905
rect 8294 7828 8300 7880
rect 8352 7828 8358 7880
rect 8588 7800 8616 7899
rect 8220 7772 8616 7800
rect 8113 7763 8171 7769
rect 8386 7732 8392 7744
rect 7392 7704 8392 7732
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8680 7732 8708 7899
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 9232 7936 9260 7967
rect 8996 7908 9260 7936
rect 8996 7896 9002 7908
rect 9674 7896 9680 7948
rect 9732 7896 9738 7948
rect 10336 7945 10364 7976
rect 10321 7939 10379 7945
rect 10321 7905 10333 7939
rect 10367 7905 10379 7939
rect 10321 7899 10379 7905
rect 10410 7896 10416 7948
rect 10468 7896 10474 7948
rect 10612 7945 10640 7976
rect 10597 7939 10655 7945
rect 10597 7905 10609 7939
rect 10643 7905 10655 7939
rect 10597 7899 10655 7905
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7868 9827 7871
rect 9858 7868 9864 7880
rect 9815 7840 9864 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 10008 7840 10149 7868
rect 10008 7828 10014 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10428 7868 10456 7896
rect 10796 7868 10824 7899
rect 10428 7840 10824 7868
rect 10137 7831 10195 7837
rect 8941 7803 8999 7809
rect 8941 7769 8953 7803
rect 8987 7800 8999 7803
rect 9398 7800 9404 7812
rect 8987 7772 9404 7800
rect 8987 7769 8999 7772
rect 8941 7763 8999 7769
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 10042 7760 10048 7812
rect 10100 7760 10106 7812
rect 9217 7735 9275 7741
rect 9217 7732 9229 7735
rect 8680 7704 9229 7732
rect 9217 7701 9229 7704
rect 9263 7732 9275 7735
rect 9766 7732 9772 7744
rect 9263 7704 9772 7732
rect 9263 7701 9275 7704
rect 9217 7695 9275 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 10502 7692 10508 7744
rect 10560 7732 10566 7744
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 10560 7704 10609 7732
rect 10560 7692 10566 7704
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10597 7695 10655 7701
rect 552 7642 11132 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 10062 7642
rect 10114 7590 10126 7642
rect 10178 7590 10190 7642
rect 10242 7590 10254 7642
rect 10306 7590 10318 7642
rect 10370 7590 11132 7642
rect 552 7568 11132 7590
rect 1029 7531 1087 7537
rect 1029 7497 1041 7531
rect 1075 7528 1087 7531
rect 1578 7528 1584 7540
rect 1075 7500 1584 7528
rect 1075 7497 1087 7500
rect 1029 7491 1087 7497
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2130 7528 2136 7540
rect 1688 7500 2136 7528
rect 937 7463 995 7469
rect 937 7429 949 7463
rect 983 7460 995 7463
rect 1394 7460 1400 7472
rect 983 7432 1400 7460
rect 983 7429 995 7432
rect 937 7423 995 7429
rect 1394 7420 1400 7432
rect 1452 7420 1458 7472
rect 1121 7395 1179 7401
rect 1121 7361 1133 7395
rect 1167 7361 1179 7395
rect 1121 7355 1179 7361
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7392 1547 7395
rect 1578 7392 1584 7404
rect 1535 7364 1584 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 845 7327 903 7333
rect 845 7293 857 7327
rect 891 7293 903 7327
rect 845 7287 903 7293
rect 860 7188 888 7287
rect 1136 7256 1164 7355
rect 1578 7352 1584 7364
rect 1636 7352 1642 7404
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 1688 7324 1716 7500
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 3142 7528 3148 7540
rect 2915 7500 3148 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 4120 7500 5365 7528
rect 4120 7488 4126 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5353 7491 5411 7497
rect 6730 7488 6736 7540
rect 6788 7488 6794 7540
rect 7374 7528 7380 7540
rect 6831 7500 7380 7528
rect 1765 7463 1823 7469
rect 1765 7429 1777 7463
rect 1811 7429 1823 7463
rect 1765 7423 1823 7429
rect 1780 7392 1808 7423
rect 2406 7420 2412 7472
rect 2464 7420 2470 7472
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 6831 7460 6859 7500
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 7558 7488 7564 7540
rect 7616 7488 7622 7540
rect 7650 7488 7656 7540
rect 7708 7488 7714 7540
rect 8938 7488 8944 7540
rect 8996 7528 9002 7540
rect 9033 7531 9091 7537
rect 9033 7528 9045 7531
rect 8996 7500 9045 7528
rect 8996 7488 9002 7500
rect 9033 7497 9045 7500
rect 9079 7497 9091 7531
rect 9033 7491 9091 7497
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 9732 7500 10517 7528
rect 9732 7488 9738 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 10505 7491 10563 7497
rect 5592 7432 6859 7460
rect 5592 7420 5598 7432
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1780 7364 1961 7392
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2832 7364 2973 7392
rect 2832 7352 2838 7364
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5859 7364 6009 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 5997 7361 6009 7364
rect 6043 7361 6055 7395
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 5997 7355 6055 7361
rect 6196 7364 7021 7392
rect 6196 7336 6224 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7558 7392 7564 7404
rect 7009 7355 7067 7361
rect 7116 7364 7564 7392
rect 1443 7296 1716 7324
rect 2041 7327 2099 7333
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 2041 7293 2053 7327
rect 2087 7324 2099 7327
rect 2406 7324 2412 7336
rect 2087 7296 2412 7324
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 2406 7284 2412 7296
rect 2464 7324 2470 7336
rect 2685 7327 2743 7333
rect 2685 7324 2697 7327
rect 2464 7296 2697 7324
rect 2464 7284 2470 7296
rect 2685 7293 2697 7296
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 2924 7296 3433 7324
rect 2924 7284 2930 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 3605 7327 3663 7333
rect 3605 7324 3617 7327
rect 3568 7296 3617 7324
rect 3568 7284 3574 7296
rect 3605 7293 3617 7296
rect 3651 7324 3663 7327
rect 3878 7324 3884 7336
rect 3651 7296 3884 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 4304 7296 4629 7324
rect 4304 7284 4310 7296
rect 4617 7293 4629 7296
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7324 4859 7327
rect 5074 7324 5080 7336
rect 4847 7296 5080 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 5534 7284 5540 7336
rect 5592 7284 5598 7336
rect 5718 7284 5724 7336
rect 5776 7284 5782 7336
rect 5902 7284 5908 7336
rect 5960 7284 5966 7336
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 2222 7256 2228 7268
rect 1136 7228 2228 7256
rect 2222 7216 2228 7228
rect 2280 7216 2286 7268
rect 5810 7216 5816 7268
rect 5868 7256 5874 7268
rect 6104 7256 6132 7287
rect 6178 7284 6184 7336
rect 6236 7284 6242 7336
rect 6362 7284 6368 7336
rect 6420 7284 6426 7336
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6604 7296 6653 7324
rect 6604 7284 6610 7296
rect 6641 7293 6653 7296
rect 6687 7293 6699 7327
rect 6816 7329 6874 7335
rect 7116 7333 7144 7364
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 8754 7392 8760 7404
rect 8036 7364 8760 7392
rect 6816 7326 6828 7329
rect 6641 7287 6699 7293
rect 6748 7298 6828 7326
rect 6748 7268 6776 7298
rect 6816 7295 6828 7298
rect 6862 7295 6874 7329
rect 6816 7289 6874 7295
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 5868 7228 6132 7256
rect 5868 7216 5874 7228
rect 6454 7216 6460 7268
rect 6512 7256 6518 7268
rect 6730 7256 6736 7268
rect 6512 7228 6736 7256
rect 6512 7216 6518 7228
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 1578 7188 1584 7200
rect 860 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1854 7148 1860 7200
rect 1912 7188 1918 7200
rect 2501 7191 2559 7197
rect 2501 7188 2513 7191
rect 1912 7160 2513 7188
rect 1912 7148 1918 7160
rect 2501 7157 2513 7160
rect 2547 7157 2559 7191
rect 2501 7151 2559 7157
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 3789 7191 3847 7197
rect 3789 7188 3801 7191
rect 3568 7160 3801 7188
rect 3568 7148 3574 7160
rect 3789 7157 3801 7160
rect 3835 7157 3847 7191
rect 3789 7151 3847 7157
rect 4709 7191 4767 7197
rect 4709 7157 4721 7191
rect 4755 7188 4767 7191
rect 4982 7188 4988 7200
rect 4755 7160 4988 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 6270 7148 6276 7200
rect 6328 7148 6334 7200
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 6932 7188 6960 7287
rect 6604 7160 6960 7188
rect 6604 7148 6610 7160
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7116 7188 7144 7287
rect 7190 7284 7196 7336
rect 7248 7324 7254 7336
rect 8036 7333 8064 7364
rect 8754 7352 8760 7364
rect 8812 7392 8818 7404
rect 9214 7392 9220 7404
rect 8812 7364 9220 7392
rect 8812 7352 8818 7364
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 9600 7364 10548 7392
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 7248 7296 7297 7324
rect 7248 7284 7254 7296
rect 7285 7293 7297 7296
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 7423 7296 8033 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 8021 7293 8033 7296
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 7300 7256 7328 7287
rect 8478 7284 8484 7336
rect 8536 7324 8542 7336
rect 9122 7324 9128 7336
rect 8536 7296 9128 7324
rect 8536 7284 8542 7296
rect 9122 7284 9128 7296
rect 9180 7324 9186 7336
rect 9600 7333 9628 7364
rect 10520 7336 10548 7364
rect 9309 7327 9367 7333
rect 9309 7324 9321 7327
rect 9180 7296 9321 7324
rect 9180 7284 9186 7296
rect 9309 7293 9321 7296
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7324 9827 7327
rect 9858 7324 9864 7336
rect 9815 7296 9864 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 9858 7284 9864 7296
rect 9916 7284 9922 7336
rect 9950 7284 9956 7336
rect 10008 7324 10014 7336
rect 10045 7327 10103 7333
rect 10045 7324 10057 7327
rect 10008 7296 10057 7324
rect 10008 7284 10014 7296
rect 10045 7293 10057 7296
rect 10091 7324 10103 7327
rect 10321 7327 10379 7333
rect 10321 7324 10333 7327
rect 10091 7296 10333 7324
rect 10091 7293 10103 7296
rect 10045 7287 10103 7293
rect 10321 7293 10333 7296
rect 10367 7293 10379 7327
rect 10321 7287 10379 7293
rect 10502 7284 10508 7336
rect 10560 7284 10566 7336
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7300 7228 7849 7256
rect 7837 7225 7849 7228
rect 7883 7256 7895 7259
rect 8754 7256 8760 7268
rect 7883 7228 8760 7256
rect 7883 7225 7895 7228
rect 7837 7219 7895 7225
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 7064 7160 7144 7188
rect 7064 7148 7070 7160
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 9916 7160 10241 7188
rect 9916 7148 9922 7160
rect 10229 7157 10241 7160
rect 10275 7157 10287 7191
rect 10229 7151 10287 7157
rect 552 7098 11132 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 10722 7098
rect 10774 7046 10786 7098
rect 10838 7046 10850 7098
rect 10902 7046 10914 7098
rect 10966 7046 10978 7098
rect 11030 7046 11132 7098
rect 552 7024 11132 7046
rect 2222 6944 2228 6996
rect 2280 6944 2286 6996
rect 3878 6984 3884 6996
rect 2976 6956 3884 6984
rect 1946 6916 1952 6928
rect 1596 6888 1952 6916
rect 1213 6851 1271 6857
rect 1213 6817 1225 6851
rect 1259 6817 1271 6851
rect 1596 6848 1624 6888
rect 1946 6876 1952 6888
rect 2004 6916 2010 6928
rect 2004 6888 2176 6916
rect 2004 6876 2010 6888
rect 1213 6811 1271 6817
rect 1320 6820 1624 6848
rect 1228 6644 1256 6811
rect 1320 6789 1348 6820
rect 1670 6808 1676 6860
rect 1728 6808 1734 6860
rect 1854 6808 1860 6860
rect 1912 6808 1918 6860
rect 2148 6857 2176 6888
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6817 2099 6851
rect 2041 6811 2099 6817
rect 2133 6851 2191 6857
rect 2133 6817 2145 6851
rect 2179 6817 2191 6851
rect 2133 6811 2191 6817
rect 1305 6783 1363 6789
rect 1305 6749 1317 6783
rect 1351 6749 1363 6783
rect 1305 6743 1363 6749
rect 1486 6740 1492 6792
rect 1544 6780 1550 6792
rect 1581 6783 1639 6789
rect 1581 6780 1593 6783
rect 1544 6752 1593 6780
rect 1544 6740 1550 6752
rect 1581 6749 1593 6752
rect 1627 6749 1639 6783
rect 2056 6780 2084 6811
rect 2222 6808 2228 6860
rect 2280 6808 2286 6860
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2498 6848 2504 6860
rect 2455 6820 2504 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2682 6808 2688 6860
rect 2740 6808 2746 6860
rect 2777 6851 2835 6857
rect 2777 6817 2789 6851
rect 2823 6848 2835 6851
rect 2866 6848 2872 6860
rect 2823 6820 2872 6848
rect 2823 6817 2835 6820
rect 2777 6811 2835 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 2976 6857 3004 6956
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 5629 6987 5687 6993
rect 5629 6953 5641 6987
rect 5675 6984 5687 6987
rect 5902 6984 5908 6996
rect 5675 6956 5908 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 6917 6987 6975 6993
rect 6917 6953 6929 6987
rect 6963 6984 6975 6987
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 6963 6956 7941 6984
rect 6963 6953 6975 6956
rect 6917 6947 6975 6953
rect 7929 6953 7941 6956
rect 7975 6984 7987 6987
rect 8202 6984 8208 6996
rect 7975 6956 8208 6984
rect 7975 6953 7987 6956
rect 7929 6947 7987 6953
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 9180 6956 9413 6984
rect 9180 6944 9186 6956
rect 9401 6953 9413 6956
rect 9447 6984 9459 6987
rect 9582 6984 9588 6996
rect 9447 6956 9588 6984
rect 9447 6953 9459 6956
rect 9401 6947 9459 6953
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 7466 6916 7472 6928
rect 3804 6888 4200 6916
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6817 3019 6851
rect 2961 6811 3019 6817
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3804 6848 3832 6888
rect 3292 6820 3832 6848
rect 3881 6851 3939 6857
rect 3292 6808 3298 6820
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 4062 6848 4068 6860
rect 3927 6820 4068 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4172 6848 4200 6888
rect 7300 6888 7472 6916
rect 4341 6851 4399 6857
rect 4341 6848 4353 6851
rect 4172 6820 4353 6848
rect 4341 6817 4353 6820
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6848 4583 6851
rect 4706 6848 4712 6860
rect 4571 6820 4712 6848
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6817 4859 6851
rect 4801 6811 4859 6817
rect 2240 6780 2268 6808
rect 2700 6780 2728 6808
rect 2056 6752 2728 6780
rect 1581 6743 1639 6749
rect 3142 6740 3148 6792
rect 3200 6740 3206 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3620 6752 3801 6780
rect 1394 6672 1400 6724
rect 1452 6712 1458 6724
rect 3620 6721 3648 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 4816 6780 4844 6811
rect 4982 6808 4988 6860
rect 5040 6808 5046 6860
rect 5258 6808 5264 6860
rect 5316 6808 5322 6860
rect 5997 6851 6055 6857
rect 5997 6817 6009 6851
rect 6043 6848 6055 6851
rect 6178 6848 6184 6860
rect 6043 6820 6184 6848
rect 6043 6817 6055 6820
rect 5997 6811 6055 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6270 6808 6276 6860
rect 6328 6848 6334 6860
rect 6549 6851 6607 6857
rect 6549 6848 6561 6851
rect 6328 6820 6561 6848
rect 6328 6808 6334 6820
rect 6549 6817 6561 6820
rect 6595 6817 6607 6851
rect 6914 6848 6920 6860
rect 6549 6811 6607 6817
rect 6656 6820 6920 6848
rect 6656 6789 6684 6820
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7193 6851 7251 6857
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 7300 6848 7328 6888
rect 7466 6876 7472 6888
rect 7524 6876 7530 6928
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7239 6820 7328 6848
rect 7392 6820 7757 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 5353 6783 5411 6789
rect 5353 6780 5365 6783
rect 4816 6752 5365 6780
rect 3789 6743 3847 6749
rect 5353 6749 5365 6752
rect 5399 6780 5411 6783
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5399 6752 5825 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 6641 6783 6699 6789
rect 6641 6780 6653 6783
rect 5813 6743 5871 6749
rect 6196 6752 6653 6780
rect 2501 6715 2559 6721
rect 2501 6712 2513 6715
rect 1452 6684 2513 6712
rect 1452 6672 1458 6684
rect 2501 6681 2513 6684
rect 2547 6681 2559 6715
rect 2501 6675 2559 6681
rect 3605 6715 3663 6721
rect 3605 6681 3617 6715
rect 3651 6681 3663 6715
rect 3605 6675 3663 6681
rect 4249 6715 4307 6721
rect 4249 6681 4261 6715
rect 4295 6712 4307 6715
rect 5166 6712 5172 6724
rect 4295 6684 5172 6712
rect 4295 6681 4307 6684
rect 4249 6675 4307 6681
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 6196 6721 6224 6752
rect 6641 6749 6653 6752
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6880 6752 7021 6780
rect 6880 6740 6886 6752
rect 7009 6749 7021 6752
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 6181 6715 6239 6721
rect 6181 6681 6193 6715
rect 6227 6681 6239 6715
rect 7392 6712 7420 6820
rect 7745 6817 7757 6820
rect 7791 6848 7803 6851
rect 7791 6820 7880 6848
rect 7791 6817 7803 6820
rect 7745 6811 7803 6817
rect 7469 6783 7527 6789
rect 7469 6749 7481 6783
rect 7515 6780 7527 6783
rect 7852 6780 7880 6820
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 8113 6851 8171 6857
rect 8113 6848 8125 6851
rect 8076 6820 8125 6848
rect 8076 6808 8082 6820
rect 8113 6817 8125 6820
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 8260 6820 8309 6848
rect 8260 6808 8266 6820
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9272 6820 9321 6848
rect 9272 6808 9278 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 9548 6820 9597 6848
rect 9548 6808 9554 6820
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 8846 6780 8852 6792
rect 7515 6752 7788 6780
rect 7852 6752 8852 6780
rect 7515 6749 7527 6752
rect 7469 6743 7527 6749
rect 6181 6675 6239 6681
rect 7208 6684 7420 6712
rect 1486 6644 1492 6656
rect 1228 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6644 3019 6647
rect 3418 6644 3424 6656
rect 3007 6616 3424 6644
rect 3007 6613 3019 6616
rect 2961 6607 3019 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 4614 6644 4620 6656
rect 3936 6616 4620 6644
rect 3936 6604 3942 6616
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6822 6644 6828 6656
rect 5592 6616 6828 6644
rect 5592 6604 5598 6616
rect 6822 6604 6828 6616
rect 6880 6644 6886 6656
rect 7208 6644 7236 6684
rect 6880 6616 7236 6644
rect 7377 6647 7435 6653
rect 6880 6604 6886 6616
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 7561 6647 7619 6653
rect 7561 6644 7573 6647
rect 7423 6616 7573 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7561 6613 7573 6616
rect 7607 6613 7619 6647
rect 7760 6644 7788 6752
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 8113 6647 8171 6653
rect 8113 6644 8125 6647
rect 7760 6616 8125 6644
rect 7561 6607 7619 6613
rect 8113 6613 8125 6616
rect 8159 6613 8171 6647
rect 8113 6607 8171 6613
rect 9766 6604 9772 6656
rect 9824 6604 9830 6656
rect 552 6554 11132 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 10062 6554
rect 10114 6502 10126 6554
rect 10178 6502 10190 6554
rect 10242 6502 10254 6554
rect 10306 6502 10318 6554
rect 10370 6502 11132 6554
rect 552 6480 11132 6502
rect 2406 6400 2412 6452
rect 2464 6400 2470 6452
rect 3510 6400 3516 6452
rect 3568 6440 3574 6452
rect 3697 6443 3755 6449
rect 3697 6440 3709 6443
rect 3568 6412 3709 6440
rect 3568 6400 3574 6412
rect 3697 6409 3709 6412
rect 3743 6409 3755 6443
rect 3697 6403 3755 6409
rect 3421 6375 3479 6381
rect 3421 6372 3433 6375
rect 2746 6344 3433 6372
rect 1394 6196 1400 6248
rect 1452 6236 1458 6248
rect 2038 6236 2044 6248
rect 1452 6208 2044 6236
rect 1452 6196 1458 6208
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 2130 6196 2136 6248
rect 2188 6196 2194 6248
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2746 6236 2774 6344
rect 3421 6341 3433 6344
rect 3467 6341 3479 6375
rect 3421 6335 3479 6341
rect 2271 6208 2774 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 1946 6128 1952 6180
rect 2004 6168 2010 6180
rect 2240 6168 2268 6199
rect 3234 6196 3240 6248
rect 3292 6196 3298 6248
rect 3418 6196 3424 6248
rect 3476 6196 3482 6248
rect 3712 6236 3740 6403
rect 4706 6400 4712 6452
rect 4764 6400 4770 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5258 6440 5264 6452
rect 5031 6412 5264 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5353 6443 5411 6449
rect 5353 6409 5365 6443
rect 5399 6440 5411 6443
rect 5718 6440 5724 6452
rect 5399 6412 5724 6440
rect 5399 6409 5411 6412
rect 5353 6403 5411 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 6362 6400 6368 6452
rect 6420 6400 6426 6452
rect 7098 6400 7104 6452
rect 7156 6400 7162 6452
rect 3786 6332 3792 6384
rect 3844 6332 3850 6384
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 4304 6276 4353 6304
rect 4304 6264 4310 6276
rect 4341 6273 4353 6276
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 3789 6239 3847 6245
rect 3789 6236 3801 6239
rect 3712 6208 3801 6236
rect 3789 6205 3801 6208
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 4525 6239 4583 6245
rect 4525 6205 4537 6239
rect 4571 6205 4583 6239
rect 4724 6236 4752 6400
rect 7282 6372 7288 6384
rect 6932 6344 7288 6372
rect 6932 6304 6960 6344
rect 7282 6332 7288 6344
rect 7340 6332 7346 6384
rect 6840 6276 6960 6304
rect 7009 6307 7067 6313
rect 4801 6239 4859 6245
rect 4801 6236 4813 6239
rect 4724 6208 4813 6236
rect 4525 6199 4583 6205
rect 4801 6205 4813 6208
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 2004 6140 2268 6168
rect 3436 6168 3464 6196
rect 3988 6168 4016 6199
rect 3436 6140 4016 6168
rect 4540 6168 4568 6199
rect 4982 6196 4988 6248
rect 5040 6196 5046 6248
rect 5534 6196 5540 6248
rect 5592 6196 5598 6248
rect 5810 6196 5816 6248
rect 5868 6196 5874 6248
rect 6454 6196 6460 6248
rect 6512 6196 6518 6248
rect 6840 6245 6868 6276
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7374 6304 7380 6316
rect 7055 6276 7380 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 7524 6276 8984 6304
rect 7524 6264 7530 6276
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 5074 6168 5080 6180
rect 4540 6140 5080 6168
rect 2004 6128 2010 6140
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 5721 6171 5779 6177
rect 5721 6137 5733 6171
rect 5767 6168 5779 6171
rect 5902 6168 5908 6180
rect 5767 6140 5908 6168
rect 5767 6137 5779 6140
rect 5721 6131 5779 6137
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 5997 6171 6055 6177
rect 5997 6137 6009 6171
rect 6043 6168 6055 6171
rect 6086 6168 6092 6180
rect 6043 6140 6092 6168
rect 6043 6137 6055 6140
rect 5997 6131 6055 6137
rect 6086 6128 6092 6140
rect 6144 6128 6150 6180
rect 6181 6171 6239 6177
rect 6181 6137 6193 6171
rect 6227 6168 6239 6171
rect 6546 6168 6552 6180
rect 6227 6140 6552 6168
rect 6227 6137 6239 6140
rect 6181 6131 6239 6137
rect 6546 6128 6552 6140
rect 6604 6128 6610 6180
rect 6656 6168 6684 6199
rect 6914 6196 6920 6248
rect 6972 6196 6978 6248
rect 7190 6196 7196 6248
rect 7248 6196 7254 6248
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 8110 6236 8116 6248
rect 7331 6208 8116 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8956 6245 8984 6276
rect 8941 6239 8999 6245
rect 8941 6205 8953 6239
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 9122 6196 9128 6248
rect 9180 6196 9186 6248
rect 9217 6239 9275 6245
rect 9217 6205 9229 6239
rect 9263 6236 9275 6239
rect 10410 6236 10416 6248
rect 9263 6208 10416 6236
rect 9263 6205 9275 6208
rect 9217 6199 9275 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 7098 6168 7104 6180
rect 6656 6140 7104 6168
rect 7098 6128 7104 6140
rect 7156 6128 7162 6180
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6100 1823 6103
rect 2406 6100 2412 6112
rect 1811 6072 2412 6100
rect 1811 6069 1823 6072
rect 1765 6063 1823 6069
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 3016 6072 8769 6100
rect 3016 6060 3022 6072
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8757 6063 8815 6069
rect 552 6010 11132 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 10722 6010
rect 10774 5958 10786 6010
rect 10838 5958 10850 6010
rect 10902 5958 10914 6010
rect 10966 5958 10978 6010
rect 11030 5958 11132 6010
rect 552 5936 11132 5958
rect 1305 5899 1363 5905
rect 1305 5865 1317 5899
rect 1351 5896 1363 5899
rect 2406 5896 2412 5908
rect 1351 5868 2412 5896
rect 1351 5865 1363 5868
rect 1305 5859 1363 5865
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5896 2743 5899
rect 3050 5896 3056 5908
rect 2731 5868 3056 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 7248 5868 7481 5896
rect 7248 5856 7254 5868
rect 7469 5865 7481 5868
rect 7515 5865 7527 5899
rect 7469 5859 7527 5865
rect 8110 5856 8116 5908
rect 8168 5856 8174 5908
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 9309 5899 9367 5905
rect 9309 5896 9321 5899
rect 9180 5868 9321 5896
rect 9180 5856 9186 5868
rect 9309 5865 9321 5868
rect 9355 5865 9367 5899
rect 9309 5859 9367 5865
rect 10410 5856 10416 5908
rect 10468 5856 10474 5908
rect 2869 5831 2927 5837
rect 2869 5828 2881 5831
rect 1688 5800 2881 5828
rect 1213 5763 1271 5769
rect 1213 5729 1225 5763
rect 1259 5729 1271 5763
rect 1213 5723 1271 5729
rect 1228 5692 1256 5723
rect 1394 5720 1400 5772
rect 1452 5720 1458 5772
rect 1688 5769 1716 5800
rect 2869 5797 2881 5800
rect 2915 5797 2927 5831
rect 2869 5791 2927 5797
rect 5074 5788 5080 5840
rect 5132 5828 5138 5840
rect 5132 5800 6592 5828
rect 5132 5788 5138 5800
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 2317 5763 2375 5769
rect 2317 5760 2329 5763
rect 1912 5732 2329 5760
rect 1912 5720 1918 5732
rect 2317 5729 2329 5732
rect 2363 5729 2375 5763
rect 2317 5723 2375 5729
rect 2406 5720 2412 5772
rect 2464 5760 2470 5772
rect 2777 5763 2835 5769
rect 2777 5760 2789 5763
rect 2464 5732 2789 5760
rect 2464 5720 2470 5732
rect 2777 5729 2789 5732
rect 2823 5729 2835 5763
rect 2777 5723 2835 5729
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5729 3019 5763
rect 2961 5723 3019 5729
rect 1486 5692 1492 5704
rect 1228 5664 1492 5692
rect 1486 5652 1492 5664
rect 1544 5652 1550 5704
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5692 1823 5695
rect 1946 5692 1952 5704
rect 1811 5664 1952 5692
rect 1811 5661 1823 5664
rect 1765 5655 1823 5661
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 2225 5695 2283 5701
rect 2225 5692 2237 5695
rect 2056 5664 2237 5692
rect 2056 5633 2084 5664
rect 2225 5661 2237 5664
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2041 5627 2099 5633
rect 2041 5593 2053 5627
rect 2087 5593 2099 5627
rect 2041 5587 2099 5593
rect 2130 5584 2136 5636
rect 2188 5624 2194 5636
rect 2976 5624 3004 5723
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 5868 5732 6193 5760
rect 5868 5720 5874 5732
rect 6181 5729 6193 5732
rect 6227 5729 6239 5763
rect 6181 5723 6239 5729
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 5592 5664 6285 5692
rect 5592 5652 5598 5664
rect 6273 5661 6285 5664
rect 6319 5692 6331 5695
rect 6454 5692 6460 5704
rect 6319 5664 6460 5692
rect 6319 5661 6331 5664
rect 6273 5655 6331 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 2188 5596 3004 5624
rect 2188 5584 2194 5596
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 5902 5624 5908 5636
rect 5408 5596 5908 5624
rect 5408 5584 5414 5596
rect 5902 5584 5908 5596
rect 5960 5584 5966 5636
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 5813 5559 5871 5565
rect 5813 5556 5825 5559
rect 5776 5528 5825 5556
rect 5776 5516 5782 5528
rect 5813 5525 5825 5528
rect 5859 5525 5871 5559
rect 6564 5556 6592 5800
rect 6822 5788 6828 5840
rect 6880 5828 6886 5840
rect 6880 5800 7696 5828
rect 6880 5788 6886 5800
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 7282 5760 7288 5772
rect 7055 5732 7288 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7668 5769 7696 5800
rect 7944 5800 8248 5828
rect 7653 5763 7711 5769
rect 7653 5729 7665 5763
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 7834 5720 7840 5772
rect 7892 5720 7898 5772
rect 7944 5769 7972 5800
rect 8220 5769 8248 5800
rect 8846 5788 8852 5840
rect 8904 5828 8910 5840
rect 9677 5831 9735 5837
rect 8904 5800 9536 5828
rect 8904 5788 8910 5800
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5729 7987 5763
rect 7929 5723 7987 5729
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 8938 5760 8944 5772
rect 8251 5732 8944 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7852 5692 7880 5720
rect 8036 5692 8064 5723
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 9508 5769 9536 5800
rect 9677 5797 9689 5831
rect 9723 5828 9735 5831
rect 10229 5831 10287 5837
rect 10229 5828 10241 5831
rect 9723 5800 10241 5828
rect 9723 5797 9735 5800
rect 9677 5791 9735 5797
rect 10229 5797 10241 5800
rect 10275 5828 10287 5831
rect 10275 5800 10548 5828
rect 10275 5797 10287 5800
rect 10229 5791 10287 5797
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 9769 5763 9827 5769
rect 9769 5760 9781 5763
rect 9640 5732 9781 5760
rect 9640 5720 9646 5732
rect 9769 5729 9781 5732
rect 9815 5760 9827 5763
rect 9815 5732 9996 5760
rect 9815 5729 9827 5732
rect 9769 5723 9827 5729
rect 7852 5664 8064 5692
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9968 5692 9996 5732
rect 10042 5720 10048 5772
rect 10100 5720 10106 5772
rect 10520 5769 10548 5800
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 10505 5763 10563 5769
rect 10505 5729 10517 5763
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5729 10655 5763
rect 10597 5723 10655 5729
rect 10336 5692 10364 5723
rect 9968 5664 10364 5692
rect 9861 5655 9919 5661
rect 7377 5627 7435 5633
rect 7377 5593 7389 5627
rect 7423 5624 7435 5627
rect 8018 5624 8024 5636
rect 7423 5596 8024 5624
rect 7423 5593 7435 5596
rect 7377 5587 7435 5593
rect 8018 5584 8024 5596
rect 8076 5584 8082 5636
rect 8570 5556 8576 5568
rect 6564 5528 8576 5556
rect 5813 5519 5871 5525
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 9876 5556 9904 5655
rect 10410 5652 10416 5704
rect 10468 5692 10474 5704
rect 10612 5692 10640 5723
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 10744 5732 10793 5760
rect 10744 5720 10750 5732
rect 10781 5729 10793 5732
rect 10827 5729 10839 5763
rect 10781 5723 10839 5729
rect 10468 5664 10640 5692
rect 10468 5652 10474 5664
rect 9456 5528 9904 5556
rect 9456 5516 9462 5528
rect 10686 5516 10692 5568
rect 10744 5516 10750 5568
rect 552 5466 11132 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 10062 5466
rect 10114 5414 10126 5466
rect 10178 5414 10190 5466
rect 10242 5414 10254 5466
rect 10306 5414 10318 5466
rect 10370 5414 11132 5466
rect 552 5392 11132 5414
rect 2130 5312 2136 5364
rect 2188 5312 2194 5364
rect 6914 5312 6920 5364
rect 6972 5312 6978 5364
rect 7009 5355 7067 5361
rect 7009 5321 7021 5355
rect 7055 5352 7067 5355
rect 7098 5352 7104 5364
rect 7055 5324 7104 5352
rect 7055 5321 7067 5324
rect 7009 5315 7067 5321
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 8478 5312 8484 5364
rect 8536 5352 8542 5364
rect 9398 5352 9404 5364
rect 8536 5324 9404 5352
rect 8536 5312 8542 5324
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 3789 5287 3847 5293
rect 3789 5253 3801 5287
rect 3835 5284 3847 5287
rect 4062 5284 4068 5296
rect 3835 5256 4068 5284
rect 3835 5253 3847 5256
rect 3789 5247 3847 5253
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 5810 5244 5816 5296
rect 5868 5244 5874 5296
rect 9582 5244 9588 5296
rect 9640 5244 9646 5296
rect 10597 5287 10655 5293
rect 10597 5284 10609 5287
rect 9876 5256 10609 5284
rect 9876 5228 9904 5256
rect 10597 5253 10609 5256
rect 10643 5253 10655 5287
rect 10597 5247 10655 5253
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 1728 5188 2452 5216
rect 1728 5176 1734 5188
rect 1486 5108 1492 5160
rect 1544 5148 1550 5160
rect 2424 5157 2452 5188
rect 3510 5176 3516 5228
rect 3568 5176 3574 5228
rect 5092 5188 5488 5216
rect 2409 5151 2467 5157
rect 1544 5120 1992 5148
rect 1544 5108 1550 5120
rect 1394 5040 1400 5092
rect 1452 5080 1458 5092
rect 1762 5080 1768 5092
rect 1452 5052 1768 5080
rect 1452 5040 1458 5052
rect 1762 5040 1768 5052
rect 1820 5040 1826 5092
rect 1964 5089 1992 5120
rect 2409 5117 2421 5151
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 1949 5083 2007 5089
rect 1949 5049 1961 5083
rect 1995 5080 2007 5083
rect 2038 5080 2044 5092
rect 1995 5052 2044 5080
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 2038 5040 2044 5052
rect 2096 5080 2102 5092
rect 2516 5080 2544 5111
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 5092 5157 5120 5188
rect 5460 5160 5488 5188
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 8757 5219 8815 5225
rect 6696 5188 8432 5216
rect 6696 5176 6702 5188
rect 3421 5151 3479 5157
rect 3421 5148 3433 5151
rect 3200 5120 3433 5148
rect 3200 5108 3206 5120
rect 3421 5117 3433 5120
rect 3467 5148 3479 5151
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 3467 5120 4905 5148
rect 3467 5117 3479 5120
rect 3421 5111 3479 5117
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 5350 5108 5356 5160
rect 5408 5108 5414 5160
rect 5442 5108 5448 5160
rect 5500 5108 5506 5160
rect 5568 5151 5626 5157
rect 5568 5148 5580 5151
rect 5552 5117 5580 5148
rect 5614 5117 5626 5151
rect 5552 5111 5626 5117
rect 2096 5052 2544 5080
rect 5261 5083 5319 5089
rect 2096 5040 2102 5052
rect 5261 5049 5273 5083
rect 5307 5080 5319 5083
rect 5552 5080 5580 5111
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6273 5151 6331 5157
rect 6273 5148 6285 5151
rect 6052 5120 6285 5148
rect 6052 5108 6058 5120
rect 6273 5117 6285 5120
rect 6319 5117 6331 5151
rect 6273 5111 6331 5117
rect 6546 5108 6552 5160
rect 6604 5108 6610 5160
rect 7208 5157 7236 5188
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 7282 5108 7288 5160
rect 7340 5108 7346 5160
rect 7852 5157 7880 5188
rect 8404 5157 8432 5188
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 8803 5188 9076 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 9048 5157 9076 5188
rect 9858 5176 9864 5228
rect 9916 5176 9922 5228
rect 10686 5216 10692 5228
rect 9968 5188 10692 5216
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5117 7895 5151
rect 7837 5111 7895 5117
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5117 8079 5151
rect 8021 5111 8079 5117
rect 8389 5151 8447 5157
rect 8389 5117 8401 5151
rect 8435 5117 8447 5151
rect 8389 5111 8447 5117
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5148 9275 5151
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 9263 5120 9321 5148
rect 9263 5117 9275 5120
rect 9217 5111 9275 5117
rect 9309 5117 9321 5120
rect 9355 5148 9367 5151
rect 9398 5148 9404 5160
rect 9355 5120 9404 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 5905 5083 5963 5089
rect 5905 5080 5917 5083
rect 5307 5052 5917 5080
rect 5307 5049 5319 5052
rect 5261 5043 5319 5049
rect 5905 5049 5917 5052
rect 5951 5049 5963 5083
rect 5905 5043 5963 5049
rect 6089 5083 6147 5089
rect 6089 5049 6101 5083
rect 6135 5049 6147 5083
rect 6564 5080 6592 5108
rect 7300 5080 7328 5108
rect 8036 5080 8064 5111
rect 8573 5083 8631 5089
rect 8573 5080 8585 5083
rect 6564 5052 7328 5080
rect 7852 5052 8585 5080
rect 6089 5043 6147 5049
rect 2222 4972 2228 5024
rect 2280 4972 2286 5024
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 6104 5012 6132 5043
rect 5408 4984 6132 5012
rect 5408 4972 5414 4984
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 7190 5012 7196 5024
rect 6788 4984 7196 5012
rect 6788 4972 6794 4984
rect 7190 4972 7196 4984
rect 7248 5012 7254 5024
rect 7852 5012 7880 5052
rect 8573 5049 8585 5052
rect 8619 5049 8631 5083
rect 8573 5043 8631 5049
rect 7248 4984 7880 5012
rect 7248 4972 7254 4984
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8662 5012 8668 5024
rect 7984 4984 8668 5012
rect 7984 4972 7990 4984
rect 8662 4972 8668 4984
rect 8720 5012 8726 5024
rect 8864 5012 8892 5111
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 9766 5148 9772 5160
rect 9539 5120 9772 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 9968 5157 9996 5188
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 9953 5151 10011 5157
rect 9953 5117 9965 5151
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 10410 5108 10416 5160
rect 10468 5108 10474 5160
rect 8720 4984 8892 5012
rect 8720 4972 8726 4984
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 9548 4984 10241 5012
rect 9548 4972 9554 4984
rect 10229 4981 10241 4984
rect 10275 4981 10287 5015
rect 10229 4975 10287 4981
rect 552 4922 11132 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 10722 4922
rect 10774 4870 10786 4922
rect 10838 4870 10850 4922
rect 10902 4870 10914 4922
rect 10966 4870 10978 4922
rect 11030 4870 11132 4922
rect 552 4848 11132 4870
rect 1394 4808 1400 4820
rect 1136 4780 1400 4808
rect 1136 4681 1164 4780
rect 1394 4768 1400 4780
rect 1452 4768 1458 4820
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 2777 4811 2835 4817
rect 2777 4808 2789 4811
rect 2087 4780 2789 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 2222 4740 2228 4752
rect 1228 4712 2228 4740
rect 1228 4681 1256 4712
rect 2222 4700 2228 4712
rect 2280 4700 2286 4752
rect 1120 4675 1178 4681
rect 1120 4641 1132 4675
rect 1166 4641 1178 4675
rect 1120 4635 1178 4641
rect 1213 4675 1271 4681
rect 1213 4641 1225 4675
rect 1259 4641 1271 4675
rect 1213 4635 1271 4641
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4641 1547 4675
rect 1489 4635 1547 4641
rect 845 4607 903 4613
rect 845 4573 857 4607
rect 891 4604 903 4607
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 891 4576 1409 4604
rect 891 4573 903 4576
rect 845 4567 903 4573
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1504 4604 1532 4635
rect 1946 4632 1952 4684
rect 2004 4632 2010 4684
rect 2314 4632 2320 4684
rect 2372 4632 2378 4684
rect 2424 4604 2452 4780
rect 2777 4777 2789 4780
rect 2823 4777 2835 4811
rect 2777 4771 2835 4777
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 3697 4811 3755 4817
rect 3697 4808 3709 4811
rect 3568 4780 3709 4808
rect 3568 4768 3574 4780
rect 3697 4777 3709 4780
rect 3743 4777 3755 4811
rect 3697 4771 3755 4777
rect 5353 4811 5411 4817
rect 5353 4777 5365 4811
rect 5399 4808 5411 4811
rect 5442 4808 5448 4820
rect 5399 4780 5448 4808
rect 5399 4777 5411 4780
rect 5353 4771 5411 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 7834 4768 7840 4820
rect 7892 4768 7898 4820
rect 8297 4811 8355 4817
rect 8297 4808 8309 4811
rect 8220 4780 8309 4808
rect 4157 4743 4215 4749
rect 2976 4712 3372 4740
rect 2976 4681 3004 4712
rect 3344 4681 3372 4712
rect 4157 4709 4169 4743
rect 4203 4740 4215 4743
rect 4522 4740 4528 4752
rect 4203 4712 4528 4740
rect 4203 4709 4215 4712
rect 4157 4703 4215 4709
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4641 2559 4675
rect 2501 4635 2559 4641
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 2961 4675 3019 4681
rect 2961 4672 2973 4675
rect 2731 4644 2973 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 2961 4641 2973 4644
rect 3007 4641 3019 4675
rect 2961 4635 3019 4641
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 3329 4675 3387 4681
rect 3329 4641 3341 4675
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 3483 4675 3541 4681
rect 3483 4641 3495 4675
rect 3529 4672 3541 4675
rect 3789 4675 3847 4681
rect 3789 4672 3801 4675
rect 3529 4644 3801 4672
rect 3529 4641 3556 4644
rect 3483 4635 3556 4641
rect 3789 4641 3801 4644
rect 3835 4641 3847 4675
rect 3789 4635 3847 4641
rect 3973 4675 4031 4681
rect 3973 4641 3985 4675
rect 4019 4641 4031 4675
rect 3973 4635 4031 4641
rect 1504 4576 2452 4604
rect 1397 4567 1455 4573
rect 1854 4496 1860 4548
rect 1912 4496 1918 4548
rect 2516 4536 2544 4635
rect 3252 4604 3280 4635
rect 3528 4604 3556 4635
rect 3252 4576 3556 4604
rect 2516 4508 2774 4536
rect 1578 4428 1584 4480
rect 1636 4468 1642 4480
rect 2225 4471 2283 4477
rect 2225 4468 2237 4471
rect 1636 4440 2237 4468
rect 1636 4428 1642 4440
rect 2225 4437 2237 4440
rect 2271 4437 2283 4471
rect 2746 4468 2774 4508
rect 2958 4496 2964 4548
rect 3016 4536 3022 4548
rect 3988 4536 4016 4635
rect 3016 4508 4016 4536
rect 3016 4496 3022 4508
rect 4172 4468 4200 4703
rect 4522 4700 4528 4712
rect 4580 4740 4586 4752
rect 4890 4740 4896 4752
rect 4580 4712 4896 4740
rect 4580 4700 4586 4712
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 8220 4749 8248 4780
rect 8297 4777 8309 4780
rect 8343 4777 8355 4811
rect 8297 4771 8355 4777
rect 8938 4768 8944 4820
rect 8996 4768 9002 4820
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 9732 4780 9904 4808
rect 9732 4768 9738 4780
rect 8205 4743 8263 4749
rect 8205 4709 8217 4743
rect 8251 4709 8263 4743
rect 8449 4743 8507 4749
rect 8449 4740 8461 4743
rect 8205 4703 8263 4709
rect 8312 4712 8461 4740
rect 4246 4632 4252 4684
rect 4304 4672 4310 4684
rect 4706 4672 4712 4684
rect 4304 4644 4712 4672
rect 4304 4632 4310 4644
rect 4706 4632 4712 4644
rect 4764 4672 4770 4684
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4764 4644 4997 4672
rect 4764 4632 4770 4644
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 4985 4635 5043 4641
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4672 5227 4675
rect 5994 4672 6000 4684
rect 5215 4644 6000 4672
rect 5215 4641 5227 4644
rect 5169 4635 5227 4641
rect 5000 4604 5028 4635
rect 5994 4632 6000 4644
rect 6052 4672 6058 4684
rect 6052 4644 7236 4672
rect 6052 4632 6058 4644
rect 5442 4604 5448 4616
rect 5000 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 7208 4613 7236 4644
rect 7282 4632 7288 4684
rect 7340 4632 7346 4684
rect 8018 4632 8024 4684
rect 8076 4632 8082 4684
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7653 4539 7711 4545
rect 7653 4505 7665 4539
rect 7699 4536 7711 4539
rect 7834 4536 7840 4548
rect 7699 4508 7840 4536
rect 7699 4505 7711 4508
rect 7653 4499 7711 4505
rect 7834 4496 7840 4508
rect 7892 4536 7898 4548
rect 8312 4536 8340 4712
rect 8449 4709 8461 4712
rect 8495 4709 8507 4743
rect 8449 4703 8507 4709
rect 8662 4700 8668 4752
rect 8720 4700 8726 4752
rect 9398 4700 9404 4752
rect 9456 4740 9462 4752
rect 9585 4743 9643 4749
rect 9585 4740 9597 4743
rect 9456 4712 9597 4740
rect 9456 4700 9462 4712
rect 9585 4709 9597 4712
rect 9631 4709 9643 4743
rect 9585 4703 9643 4709
rect 9766 4700 9772 4752
rect 9824 4700 9830 4752
rect 9876 4740 9904 4780
rect 9950 4768 9956 4820
rect 10008 4768 10014 4820
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 10468 4780 10609 4808
rect 10468 4768 10474 4780
rect 10597 4777 10609 4780
rect 10643 4777 10655 4811
rect 10597 4771 10655 4777
rect 10229 4743 10287 4749
rect 10229 4740 10241 4743
rect 9876 4712 10241 4740
rect 10229 4709 10241 4712
rect 10275 4740 10287 4743
rect 10275 4712 10732 4740
rect 10275 4709 10287 4712
rect 10229 4703 10287 4709
rect 9306 4632 9312 4684
rect 9364 4632 9370 4684
rect 10704 4681 10732 4712
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 10091 4644 10517 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10505 4641 10517 4644
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4641 10747 4675
rect 10689 4635 10747 4641
rect 9214 4564 9220 4616
rect 9272 4604 9278 4616
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 9272 4576 9413 4604
rect 9272 4564 9278 4576
rect 9401 4573 9413 4576
rect 9447 4604 9459 4607
rect 9490 4604 9496 4616
rect 9447 4576 9496 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 10060 4536 10088 4635
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4604 10471 4607
rect 10594 4604 10600 4616
rect 10459 4576 10600 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 7892 4508 8340 4536
rect 8404 4508 10088 4536
rect 7892 4496 7898 4508
rect 2746 4440 4200 4468
rect 2225 4431 2283 4437
rect 6086 4428 6092 4480
rect 6144 4468 6150 4480
rect 7558 4468 7564 4480
rect 6144 4440 7564 4468
rect 6144 4428 6150 4440
rect 7558 4428 7564 4440
rect 7616 4468 7622 4480
rect 8404 4468 8432 4508
rect 7616 4440 8432 4468
rect 7616 4428 7622 4440
rect 8478 4428 8484 4480
rect 8536 4428 8542 4480
rect 8570 4428 8576 4480
rect 8628 4468 8634 4480
rect 9766 4468 9772 4480
rect 8628 4440 9772 4468
rect 8628 4428 8634 4440
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 552 4378 11132 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 10062 4378
rect 10114 4326 10126 4378
rect 10178 4326 10190 4378
rect 10242 4326 10254 4378
rect 10306 4326 10318 4378
rect 10370 4326 11132 4378
rect 552 4304 11132 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 1946 4264 1952 4276
rect 1452 4236 1952 4264
rect 1452 4224 1458 4236
rect 1946 4224 1952 4236
rect 2004 4224 2010 4276
rect 3326 4224 3332 4276
rect 3384 4264 3390 4276
rect 3973 4267 4031 4273
rect 3973 4264 3985 4267
rect 3384 4236 3985 4264
rect 3384 4224 3390 4236
rect 3973 4233 3985 4236
rect 4019 4233 4031 4267
rect 3973 4227 4031 4233
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 5718 4264 5724 4276
rect 4580 4236 5724 4264
rect 4580 4224 4586 4236
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 7190 4224 7196 4276
rect 7248 4264 7254 4276
rect 8665 4267 8723 4273
rect 7248 4236 8616 4264
rect 7248 4224 7254 4236
rect 2314 4156 2320 4208
rect 2372 4196 2378 4208
rect 2498 4196 2504 4208
rect 2372 4168 2504 4196
rect 2372 4156 2378 4168
rect 2498 4156 2504 4168
rect 2556 4196 2562 4208
rect 2958 4196 2964 4208
rect 2556 4168 2964 4196
rect 2556 4156 2562 4168
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 2133 4131 2191 4137
rect 2133 4128 2145 4131
rect 1820 4100 2145 4128
rect 1820 4088 1826 4100
rect 2133 4097 2145 4100
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2406 4088 2412 4140
rect 2464 4088 2470 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4097 2651 4131
rect 2792 4128 2820 4168
rect 2958 4156 2964 4168
rect 3016 4156 3022 4208
rect 3053 4199 3111 4205
rect 3053 4165 3065 4199
rect 3099 4196 3111 4199
rect 3789 4199 3847 4205
rect 3099 4168 3464 4196
rect 3099 4165 3111 4168
rect 3053 4159 3111 4165
rect 2593 4091 2651 4097
rect 2700 4100 2820 4128
rect 1946 4020 1952 4072
rect 2004 4060 2010 4072
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 2004 4032 2053 4060
rect 2004 4020 2010 4032
rect 2041 4029 2053 4032
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3961 1639 3995
rect 1581 3955 1639 3961
rect 1596 3924 1624 3955
rect 1670 3952 1676 4004
rect 1728 3992 1734 4004
rect 1765 3995 1823 4001
rect 1765 3992 1777 3995
rect 1728 3964 1777 3992
rect 1728 3952 1734 3964
rect 1765 3961 1777 3964
rect 1811 3992 1823 3995
rect 2608 3992 2636 4091
rect 2700 4069 2728 4100
rect 3436 4069 3464 4168
rect 3789 4165 3801 4199
rect 3835 4196 3847 4199
rect 3835 4168 4200 4196
rect 3835 4165 3847 4168
rect 3789 4159 3847 4165
rect 3510 4088 3516 4140
rect 3568 4088 3574 4140
rect 4172 4137 4200 4168
rect 4246 4156 4252 4208
rect 4304 4196 4310 4208
rect 5169 4199 5227 4205
rect 5169 4196 5181 4199
rect 4304 4168 5181 4196
rect 4304 4156 4310 4168
rect 5169 4165 5181 4168
rect 5215 4165 5227 4199
rect 6917 4199 6975 4205
rect 6917 4196 6929 4199
rect 5169 4159 5227 4165
rect 5460 4168 6929 4196
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4128 4859 4131
rect 5460 4128 5488 4168
rect 6917 4165 6929 4168
rect 6963 4165 6975 4199
rect 6917 4159 6975 4165
rect 7837 4199 7895 4205
rect 7837 4165 7849 4199
rect 7883 4196 7895 4199
rect 8018 4196 8024 4208
rect 7883 4168 8024 4196
rect 7883 4165 7895 4168
rect 7837 4159 7895 4165
rect 4847 4100 4936 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4029 2743 4063
rect 2685 4023 2743 4029
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4029 3479 4063
rect 3421 4023 3479 4029
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 1811 3964 2636 3992
rect 4264 3992 4292 4023
rect 4522 4020 4528 4072
rect 4580 4020 4586 4072
rect 4706 4020 4712 4072
rect 4764 4020 4770 4072
rect 4801 3995 4859 4001
rect 4801 3992 4813 3995
rect 4264 3964 4813 3992
rect 1811 3961 1823 3964
rect 1765 3955 1823 3961
rect 4801 3961 4813 3964
rect 4847 3961 4859 3995
rect 4801 3955 4859 3961
rect 2038 3924 2044 3936
rect 1596 3896 2044 3924
rect 2038 3884 2044 3896
rect 2096 3924 2102 3936
rect 2590 3924 2596 3936
rect 2096 3896 2596 3924
rect 2096 3884 2102 3896
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 4706 3884 4712 3936
rect 4764 3924 4770 3936
rect 4908 3924 4936 4100
rect 5092 4100 5488 4128
rect 5092 4072 5120 4100
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 7852 4128 7880 4159
rect 8018 4156 8024 4168
rect 8076 4156 8082 4208
rect 8478 4196 8484 4208
rect 8404 4168 8484 4196
rect 5592 4100 6859 4128
rect 5592 4088 5598 4100
rect 4982 4020 4988 4072
rect 5040 4020 5046 4072
rect 5074 4020 5080 4072
rect 5132 4020 5138 4072
rect 5350 4020 5356 4072
rect 5408 4020 5414 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4029 5687 4063
rect 5629 4023 5687 4029
rect 5258 3952 5264 4004
rect 5316 3992 5322 4004
rect 5644 3992 5672 4023
rect 5718 4020 5724 4072
rect 5776 4020 5782 4072
rect 5994 4020 6000 4072
rect 6052 4060 6058 4072
rect 6641 4063 6699 4069
rect 6641 4060 6653 4063
rect 6052 4032 6653 4060
rect 6052 4020 6058 4032
rect 6641 4029 6653 4032
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 5316 3964 5672 3992
rect 5905 3995 5963 4001
rect 5316 3952 5322 3964
rect 5905 3961 5917 3995
rect 5951 3961 5963 3995
rect 5905 3955 5963 3961
rect 4764 3896 4936 3924
rect 4764 3884 4770 3896
rect 5442 3884 5448 3936
rect 5500 3924 5506 3936
rect 5920 3924 5948 3955
rect 5500 3896 5948 3924
rect 5500 3884 5506 3896
rect 6086 3884 6092 3936
rect 6144 3884 6150 3936
rect 6730 3884 6736 3936
rect 6788 3884 6794 3936
rect 6831 3924 6859 4100
rect 6932 4100 7880 4128
rect 6932 4069 6960 4100
rect 6917 4063 6975 4069
rect 6917 4029 6929 4063
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8021 4063 8079 4069
rect 8021 4060 8033 4063
rect 7984 4032 8033 4060
rect 7984 4020 7990 4032
rect 8021 4029 8033 4032
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4060 8171 4063
rect 8404 4060 8432 4168
rect 8478 4156 8484 4168
rect 8536 4156 8542 4208
rect 8588 4196 8616 4236
rect 8665 4233 8677 4267
rect 8711 4264 8723 4267
rect 9306 4264 9312 4276
rect 8711 4236 9312 4264
rect 8711 4233 8723 4236
rect 8665 4227 8723 4233
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 8588 4168 9688 4196
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 8496 4100 9505 4128
rect 8496 4069 8524 4100
rect 8956 4069 8984 4100
rect 9493 4097 9505 4100
rect 9539 4097 9551 4131
rect 9660 4128 9688 4168
rect 9858 4128 9864 4140
rect 9660 4100 9864 4128
rect 9493 4091 9551 4097
rect 9858 4088 9864 4100
rect 9916 4128 9922 4140
rect 9916 4100 10180 4128
rect 9916 4088 9922 4100
rect 8159 4032 8432 4060
rect 8481 4063 8539 4069
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 8481 4029 8493 4063
rect 8527 4029 8539 4063
rect 8481 4023 8539 4029
rect 8665 4063 8723 4069
rect 8665 4029 8677 4063
rect 8711 4029 8723 4063
rect 8665 4023 8723 4029
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 8680 3992 8708 4023
rect 9214 4020 9220 4072
rect 9272 4020 9278 4072
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4029 9459 4063
rect 9401 4023 9459 4029
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 9766 4060 9772 4072
rect 9723 4032 9772 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 9416 3992 9444 4023
rect 9766 4020 9772 4032
rect 9824 4060 9830 4072
rect 10152 4069 10180 4100
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9824 4032 9965 4060
rect 9824 4020 9830 4032
rect 9953 4029 9965 4032
rect 9999 4029 10011 4063
rect 9953 4023 10011 4029
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4029 10195 4063
rect 10137 4023 10195 4029
rect 10045 3995 10103 4001
rect 10045 3992 10057 3995
rect 8680 3964 10057 3992
rect 10045 3961 10057 3964
rect 10091 3961 10103 3995
rect 10045 3955 10103 3961
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 6831 3896 8769 3924
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 8757 3887 8815 3893
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 9674 3924 9680 3936
rect 8904 3896 9680 3924
rect 8904 3884 8910 3896
rect 9674 3884 9680 3896
rect 9732 3924 9738 3936
rect 10594 3924 10600 3936
rect 9732 3896 10600 3924
rect 9732 3884 9738 3896
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 552 3834 11132 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 10722 3834
rect 10774 3782 10786 3834
rect 10838 3782 10850 3834
rect 10902 3782 10914 3834
rect 10966 3782 10978 3834
rect 11030 3782 11132 3834
rect 552 3760 11132 3782
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 3697 3723 3755 3729
rect 3697 3720 3709 3723
rect 3568 3692 3709 3720
rect 3568 3680 3574 3692
rect 3697 3689 3709 3692
rect 3743 3689 3755 3723
rect 6086 3720 6092 3732
rect 3697 3683 3755 3689
rect 4448 3692 6092 3720
rect 2393 3655 2451 3661
rect 2393 3621 2405 3655
rect 2439 3652 2451 3655
rect 2439 3621 2452 3652
rect 2393 3615 2452 3621
rect 2424 3584 2452 3615
rect 2590 3612 2596 3664
rect 2648 3612 2654 3664
rect 2332 3556 2452 3584
rect 3329 3587 3387 3593
rect 2332 3528 2360 3556
rect 3329 3553 3341 3587
rect 3375 3584 3387 3587
rect 4246 3584 4252 3596
rect 3375 3556 4252 3584
rect 3375 3553 3387 3556
rect 3329 3547 3387 3553
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4448 3584 4476 3692
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 8294 3720 8300 3732
rect 6236 3692 8300 3720
rect 6236 3680 6242 3692
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 9122 3720 9128 3732
rect 9048 3692 9128 3720
rect 4706 3652 4712 3664
rect 4540 3624 4712 3652
rect 4540 3593 4568 3624
rect 4706 3612 4712 3624
rect 4764 3612 4770 3664
rect 5350 3612 5356 3664
rect 5408 3652 5414 3664
rect 6549 3655 6607 3661
rect 6549 3652 6561 3655
rect 5408 3624 6561 3652
rect 5408 3612 5414 3624
rect 6549 3621 6561 3624
rect 6595 3621 6607 3655
rect 8110 3652 8116 3664
rect 6549 3615 6607 3621
rect 8036 3624 8116 3652
rect 4387 3556 4476 3584
rect 4525 3587 4583 3593
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4525 3553 4537 3587
rect 4571 3553 4583 3587
rect 4525 3547 4583 3553
rect 4614 3544 4620 3596
rect 4672 3544 4678 3596
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3553 4859 3587
rect 4801 3547 4859 3553
rect 2314 3476 2320 3528
rect 2372 3476 2378 3528
rect 2406 3476 2412 3528
rect 2464 3516 2470 3528
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 2464 3488 3249 3516
rect 2464 3476 2470 3488
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 4816 3448 4844 3547
rect 5258 3544 5264 3596
rect 5316 3544 5322 3596
rect 6178 3544 6184 3596
rect 6236 3544 6242 3596
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3553 6515 3587
rect 6457 3547 6515 3553
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5534 3516 5540 3528
rect 5399 3488 5540 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 5675 3488 6101 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 6089 3485 6101 3488
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 6472 3516 6500 3547
rect 6638 3544 6644 3596
rect 6696 3544 6702 3596
rect 7558 3544 7564 3596
rect 7616 3584 7622 3596
rect 8036 3593 8064 3624
rect 8110 3612 8116 3624
rect 8168 3652 8174 3664
rect 9048 3661 9076 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 8168 3624 9045 3652
rect 8168 3612 8174 3624
rect 9033 3621 9045 3624
rect 9079 3621 9091 3655
rect 9033 3615 9091 3621
rect 8021 3587 8079 3593
rect 7616 3556 7880 3584
rect 7616 3544 7622 3556
rect 6730 3516 6736 3528
rect 6472 3488 6736 3516
rect 6472 3448 6500 3488
rect 6730 3476 6736 3488
rect 6788 3516 6794 3528
rect 7282 3516 7288 3528
rect 6788 3488 7288 3516
rect 6788 3476 6794 3488
rect 7282 3476 7288 3488
rect 7340 3516 7346 3528
rect 7852 3516 7880 3556
rect 8021 3553 8033 3587
rect 8067 3553 8079 3587
rect 8021 3547 8079 3553
rect 8294 3544 8300 3596
rect 8352 3544 8358 3596
rect 8846 3584 8852 3596
rect 8496 3556 8852 3584
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7340 3488 7788 3516
rect 7852 3488 8217 3516
rect 7340 3476 7346 3488
rect 7760 3460 7788 3488
rect 8205 3485 8217 3488
rect 8251 3516 8263 3519
rect 8496 3516 8524 3556
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3584 9551 3587
rect 9582 3584 9588 3596
rect 9539 3556 9588 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 9140 3516 9168 3547
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 8251 3488 8524 3516
rect 8588 3488 9168 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 4816 3420 6500 3448
rect 7742 3408 7748 3460
rect 7800 3448 7806 3460
rect 8481 3451 8539 3457
rect 8481 3448 8493 3451
rect 7800 3420 8493 3448
rect 7800 3408 7806 3420
rect 8481 3417 8493 3420
rect 8527 3417 8539 3451
rect 8481 3411 8539 3417
rect 2222 3340 2228 3392
rect 2280 3340 2286 3392
rect 2409 3383 2467 3389
rect 2409 3349 2421 3383
rect 2455 3380 2467 3383
rect 2498 3380 2504 3392
rect 2455 3352 2504 3380
rect 2455 3349 2467 3352
rect 2409 3343 2467 3349
rect 2498 3340 2504 3352
rect 2556 3340 2562 3392
rect 4430 3340 4436 3392
rect 4488 3340 4494 3392
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 5718 3380 5724 3392
rect 5031 3352 5724 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 5902 3340 5908 3392
rect 5960 3340 5966 3392
rect 7282 3340 7288 3392
rect 7340 3380 7346 3392
rect 7837 3383 7895 3389
rect 7837 3380 7849 3383
rect 7340 3352 7849 3380
rect 7340 3340 7346 3352
rect 7837 3349 7849 3352
rect 7883 3380 7895 3383
rect 7926 3380 7932 3392
rect 7883 3352 7932 3380
rect 7883 3349 7895 3352
rect 7837 3343 7895 3349
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8588 3380 8616 3488
rect 8076 3352 8616 3380
rect 8665 3383 8723 3389
rect 8076 3340 8082 3352
rect 8665 3349 8677 3383
rect 8711 3380 8723 3383
rect 8754 3380 8760 3392
rect 8711 3352 8760 3380
rect 8711 3349 8723 3352
rect 8665 3343 8723 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9122 3380 9128 3392
rect 8904 3352 9128 3380
rect 8904 3340 8910 3352
rect 9122 3340 9128 3352
rect 9180 3380 9186 3392
rect 9309 3383 9367 3389
rect 9309 3380 9321 3383
rect 9180 3352 9321 3380
rect 9180 3340 9186 3352
rect 9309 3349 9321 3352
rect 9355 3349 9367 3383
rect 9309 3343 9367 3349
rect 9677 3383 9735 3389
rect 9677 3349 9689 3383
rect 9723 3380 9735 3383
rect 10502 3380 10508 3392
rect 9723 3352 10508 3380
rect 9723 3349 9735 3352
rect 9677 3343 9735 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 552 3290 11132 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 10062 3290
rect 10114 3238 10126 3290
rect 10178 3238 10190 3290
rect 10242 3238 10254 3290
rect 10306 3238 10318 3290
rect 10370 3238 11132 3290
rect 552 3216 11132 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 3602 3176 3608 3188
rect 2915 3148 3608 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 6178 3176 6184 3188
rect 5675 3148 6184 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 7190 3136 7196 3188
rect 7248 3136 7254 3188
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8294 3176 8300 3188
rect 8159 3148 8300 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 8938 3176 8944 3188
rect 8803 3148 8944 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 10413 3179 10471 3185
rect 10413 3176 10425 3179
rect 9732 3148 10425 3176
rect 9732 3136 9738 3148
rect 10413 3145 10425 3148
rect 10459 3145 10471 3179
rect 10413 3139 10471 3145
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 10689 3179 10747 3185
rect 10689 3176 10701 3179
rect 10652 3148 10701 3176
rect 10652 3136 10658 3148
rect 10689 3145 10701 3148
rect 10735 3145 10747 3179
rect 10689 3139 10747 3145
rect 2222 3068 2228 3120
rect 2280 3108 2286 3120
rect 2501 3111 2559 3117
rect 2501 3108 2513 3111
rect 2280 3080 2513 3108
rect 2280 3068 2286 3080
rect 2501 3077 2513 3080
rect 2547 3077 2559 3111
rect 3421 3111 3479 3117
rect 3421 3108 3433 3111
rect 2501 3071 2559 3077
rect 2746 3080 3433 3108
rect 1026 3000 1032 3052
rect 1084 3000 1090 3052
rect 1044 2972 1072 3000
rect 1044 2944 1624 2972
rect 1296 2907 1354 2913
rect 1296 2873 1308 2907
rect 1342 2904 1354 2907
rect 1596 2904 1624 2944
rect 2498 2932 2504 2984
rect 2556 2972 2562 2984
rect 2746 2972 2774 3080
rect 3421 3077 3433 3080
rect 3467 3077 3479 3111
rect 3421 3071 3479 3077
rect 5258 3068 5264 3120
rect 5316 3108 5322 3120
rect 5813 3111 5871 3117
rect 5813 3108 5825 3111
rect 5316 3080 5825 3108
rect 5316 3068 5322 3080
rect 5813 3077 5825 3080
rect 5859 3077 5871 3111
rect 5813 3071 5871 3077
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 4982 3040 4988 3052
rect 4488 3012 4988 3040
rect 4488 3000 4494 3012
rect 4982 3000 4988 3012
rect 5040 3040 5046 3052
rect 5169 3043 5227 3049
rect 5169 3040 5181 3043
rect 5040 3012 5181 3040
rect 5040 3000 5046 3012
rect 5169 3009 5181 3012
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 5408 3012 5948 3040
rect 5408 3000 5414 3012
rect 2556 2944 2774 2972
rect 2556 2932 2562 2944
rect 2866 2932 2872 2984
rect 2924 2972 2930 2984
rect 3050 2972 3056 2984
rect 2924 2944 3056 2972
rect 2924 2932 2930 2944
rect 3050 2932 3056 2944
rect 3108 2972 3114 2984
rect 3237 2975 3295 2981
rect 3237 2972 3249 2975
rect 3108 2944 3249 2972
rect 3108 2932 3114 2944
rect 3237 2941 3249 2944
rect 3283 2941 3295 2975
rect 3237 2935 3295 2941
rect 5074 2932 5080 2984
rect 5132 2972 5138 2984
rect 5261 2975 5319 2981
rect 5261 2972 5273 2975
rect 5132 2944 5273 2972
rect 5132 2932 5138 2944
rect 5261 2941 5273 2944
rect 5307 2941 5319 2975
rect 5261 2935 5319 2941
rect 5718 2932 5724 2984
rect 5776 2932 5782 2984
rect 5920 2981 5948 3012
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 5905 2975 5963 2981
rect 5905 2941 5917 2975
rect 5951 2941 5963 2975
rect 5905 2935 5963 2941
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 7984 2944 8401 2972
rect 7984 2932 7990 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 10502 2932 10508 2984
rect 10560 2932 10566 2984
rect 2958 2904 2964 2916
rect 1342 2876 1532 2904
rect 1596 2876 2964 2904
rect 1342 2873 1354 2876
rect 1296 2867 1354 2873
rect 1504 2836 1532 2876
rect 2958 2864 2964 2876
rect 3016 2864 3022 2916
rect 4614 2864 4620 2916
rect 4672 2904 4678 2916
rect 4890 2904 4896 2916
rect 4672 2876 4896 2904
rect 4672 2864 4678 2876
rect 4890 2864 4896 2876
rect 4948 2904 4954 2916
rect 6638 2904 6644 2916
rect 4948 2876 6644 2904
rect 4948 2864 4954 2876
rect 6638 2864 6644 2876
rect 6696 2864 6702 2916
rect 7177 2907 7235 2913
rect 7177 2873 7189 2907
rect 7223 2904 7235 2907
rect 7282 2904 7288 2916
rect 7223 2876 7288 2904
rect 7223 2873 7235 2876
rect 7177 2867 7235 2873
rect 7282 2864 7288 2876
rect 7340 2864 7346 2916
rect 7377 2907 7435 2913
rect 7377 2873 7389 2907
rect 7423 2904 7435 2907
rect 7742 2904 7748 2916
rect 7423 2876 7748 2904
rect 7423 2873 7435 2876
rect 7377 2867 7435 2873
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 7834 2864 7840 2916
rect 7892 2864 7898 2916
rect 8754 2864 8760 2916
rect 8812 2864 8818 2916
rect 9278 2907 9336 2913
rect 9278 2904 9290 2907
rect 8956 2876 9290 2904
rect 1578 2836 1584 2848
rect 1504 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 2130 2836 2136 2848
rect 1728 2808 2136 2836
rect 1728 2796 1734 2808
rect 2130 2796 2136 2808
rect 2188 2836 2194 2848
rect 2409 2839 2467 2845
rect 2409 2836 2421 2839
rect 2188 2808 2421 2836
rect 2188 2796 2194 2808
rect 2409 2805 2421 2808
rect 2455 2805 2467 2839
rect 2409 2799 2467 2805
rect 2866 2796 2872 2848
rect 2924 2796 2930 2848
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 3142 2836 3148 2848
rect 3099 2808 3148 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 7006 2796 7012 2848
rect 7064 2796 7070 2848
rect 8956 2845 8984 2876
rect 9278 2873 9290 2876
rect 9324 2873 9336 2907
rect 9278 2867 9336 2873
rect 8941 2839 8999 2845
rect 8941 2805 8953 2839
rect 8987 2805 8999 2839
rect 8941 2799 8999 2805
rect 552 2746 11132 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 10722 2746
rect 10774 2694 10786 2746
rect 10838 2694 10850 2746
rect 10902 2694 10914 2746
rect 10966 2694 10978 2746
rect 11030 2694 11132 2746
rect 552 2672 11132 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 2866 2592 2872 2644
rect 2924 2632 2930 2644
rect 3237 2635 3295 2641
rect 3237 2632 3249 2635
rect 2924 2604 3249 2632
rect 2924 2592 2930 2604
rect 3237 2601 3249 2604
rect 3283 2601 3295 2635
rect 3237 2595 3295 2601
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 7892 2604 7941 2632
rect 7892 2592 7898 2604
rect 7929 2601 7941 2604
rect 7975 2601 7987 2635
rect 7929 2595 7987 2601
rect 8018 2592 8024 2644
rect 8076 2592 8082 2644
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8938 2632 8944 2644
rect 8352 2604 8944 2632
rect 8352 2592 8358 2604
rect 8938 2592 8944 2604
rect 8996 2632 9002 2644
rect 8996 2604 9904 2632
rect 8996 2592 9002 2604
rect 1121 2567 1179 2573
rect 1121 2533 1133 2567
rect 1167 2564 1179 2567
rect 1489 2567 1547 2573
rect 1167 2536 1440 2564
rect 1167 2533 1179 2536
rect 1121 2527 1179 2533
rect 1412 2508 1440 2536
rect 1489 2533 1501 2567
rect 1535 2564 1547 2567
rect 1765 2567 1823 2573
rect 1765 2564 1777 2567
rect 1535 2536 1777 2564
rect 1535 2533 1547 2536
rect 1489 2527 1547 2533
rect 1765 2533 1777 2536
rect 1811 2533 1823 2567
rect 1765 2527 1823 2533
rect 2225 2567 2283 2573
rect 2225 2533 2237 2567
rect 2271 2564 2283 2567
rect 2314 2564 2320 2576
rect 2271 2536 2320 2564
rect 2271 2533 2283 2536
rect 2225 2527 2283 2533
rect 2314 2524 2320 2536
rect 2372 2564 2378 2576
rect 2372 2536 3464 2564
rect 2372 2524 2378 2536
rect 1305 2499 1363 2505
rect 1305 2465 1317 2499
rect 1351 2465 1363 2499
rect 1305 2459 1363 2465
rect 1320 2428 1348 2459
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 2130 2496 2136 2508
rect 1452 2468 2136 2496
rect 1452 2456 1458 2468
rect 2130 2456 2136 2468
rect 2188 2456 2194 2508
rect 2409 2499 2467 2505
rect 2409 2465 2421 2499
rect 2455 2496 2467 2499
rect 2498 2496 2504 2508
rect 2455 2468 2504 2496
rect 2455 2465 2467 2468
rect 2409 2459 2467 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 2590 2456 2596 2508
rect 2648 2496 2654 2508
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2648 2468 2789 2496
rect 2648 2456 2654 2468
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 2961 2499 3019 2505
rect 2961 2465 2973 2499
rect 3007 2496 3019 2499
rect 3234 2496 3240 2508
rect 3007 2468 3240 2496
rect 3007 2465 3019 2468
rect 2961 2459 3019 2465
rect 3234 2456 3240 2468
rect 3292 2456 3298 2508
rect 3436 2505 3464 2536
rect 3510 2524 3516 2576
rect 3568 2564 3574 2576
rect 3789 2567 3847 2573
rect 3789 2564 3801 2567
rect 3568 2536 3801 2564
rect 3568 2524 3574 2536
rect 3789 2533 3801 2536
rect 3835 2533 3847 2567
rect 9030 2564 9036 2576
rect 3789 2527 3847 2533
rect 6564 2536 9036 2564
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2465 3479 2499
rect 3421 2459 3479 2465
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 5166 2496 5172 2508
rect 4387 2468 5172 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 6564 2505 6592 2536
rect 9030 2524 9036 2536
rect 9088 2564 9094 2576
rect 9088 2536 9444 2564
rect 9088 2524 9094 2536
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2465 6607 2499
rect 6549 2459 6607 2465
rect 6816 2499 6874 2505
rect 6816 2465 6828 2499
rect 6862 2496 6874 2499
rect 7098 2496 7104 2508
rect 6862 2468 7104 2496
rect 6862 2465 6874 2468
rect 6816 2459 6874 2465
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 9416 2505 9444 2536
rect 9490 2524 9496 2576
rect 9548 2564 9554 2576
rect 9876 2573 9904 2604
rect 9645 2567 9703 2573
rect 9645 2564 9657 2567
rect 9548 2536 9657 2564
rect 9548 2524 9554 2536
rect 9645 2533 9657 2536
rect 9691 2533 9703 2567
rect 9645 2527 9703 2533
rect 9861 2567 9919 2573
rect 9861 2533 9873 2567
rect 9907 2533 9919 2567
rect 9861 2527 9919 2533
rect 9145 2499 9203 2505
rect 9145 2465 9157 2499
rect 9191 2496 9203 2499
rect 9401 2499 9459 2505
rect 9191 2468 9352 2496
rect 9191 2465 9203 2468
rect 9145 2459 9203 2465
rect 1486 2428 1492 2440
rect 1320 2400 1492 2428
rect 1486 2388 1492 2400
rect 1544 2388 1550 2440
rect 2038 2388 2044 2440
rect 2096 2428 2102 2440
rect 2516 2428 2544 2456
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2096 2400 2881 2428
rect 2096 2388 2102 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3326 2428 3332 2440
rect 3099 2400 3332 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3326 2388 3332 2400
rect 3384 2388 3390 2440
rect 9324 2428 9352 2468
rect 9401 2465 9413 2499
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 9324 2400 9536 2428
rect 1578 2320 1584 2372
rect 1636 2360 1642 2372
rect 2133 2363 2191 2369
rect 2133 2360 2145 2363
rect 1636 2332 2145 2360
rect 1636 2320 1642 2332
rect 2133 2329 2145 2332
rect 2179 2329 2191 2363
rect 2774 2360 2780 2372
rect 2133 2323 2191 2329
rect 2516 2332 2780 2360
rect 1765 2295 1823 2301
rect 1765 2261 1777 2295
rect 1811 2292 1823 2295
rect 2516 2292 2544 2332
rect 2774 2320 2780 2332
rect 2832 2360 2838 2372
rect 3602 2360 3608 2372
rect 2832 2332 3608 2360
rect 2832 2320 2838 2332
rect 3602 2320 3608 2332
rect 3660 2360 3666 2372
rect 9508 2369 9536 2400
rect 9493 2363 9551 2369
rect 3660 2332 4292 2360
rect 3660 2320 3666 2332
rect 1811 2264 2544 2292
rect 2593 2295 2651 2301
rect 1811 2261 1823 2264
rect 1765 2255 1823 2261
rect 2593 2261 2605 2295
rect 2639 2292 2651 2295
rect 3418 2292 3424 2304
rect 2639 2264 3424 2292
rect 2639 2261 2651 2264
rect 2593 2255 2651 2261
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 3804 2301 3832 2332
rect 3789 2295 3847 2301
rect 3789 2261 3801 2295
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 3973 2295 4031 2301
rect 3973 2261 3985 2295
rect 4019 2292 4031 2295
rect 4062 2292 4068 2304
rect 4019 2264 4068 2292
rect 4019 2261 4031 2264
rect 3973 2255 4031 2261
rect 4062 2252 4068 2264
rect 4120 2252 4126 2304
rect 4154 2252 4160 2304
rect 4212 2252 4218 2304
rect 4264 2292 4292 2332
rect 9493 2329 9505 2363
rect 9539 2329 9551 2363
rect 9493 2323 9551 2329
rect 6914 2292 6920 2304
rect 4264 2264 6920 2292
rect 6914 2252 6920 2264
rect 6972 2292 6978 2304
rect 8294 2292 8300 2304
rect 6972 2264 8300 2292
rect 6972 2252 6978 2264
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 8754 2252 8760 2304
rect 8812 2292 8818 2304
rect 9677 2295 9735 2301
rect 9677 2292 9689 2295
rect 8812 2264 9689 2292
rect 8812 2252 8818 2264
rect 9677 2261 9689 2264
rect 9723 2261 9735 2295
rect 9677 2255 9735 2261
rect 552 2202 11132 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 10062 2202
rect 10114 2150 10126 2202
rect 10178 2150 10190 2202
rect 10242 2150 10254 2202
rect 10306 2150 10318 2202
rect 10370 2150 11132 2202
rect 552 2128 11132 2150
rect 1578 2048 1584 2100
rect 1636 2048 1642 2100
rect 3510 2048 3516 2100
rect 3568 2088 3574 2100
rect 3697 2091 3755 2097
rect 3697 2088 3709 2091
rect 3568 2060 3709 2088
rect 3568 2048 3574 2060
rect 3697 2057 3709 2060
rect 3743 2057 3755 2091
rect 3697 2051 3755 2057
rect 3804 2060 4752 2088
rect 3602 2020 3608 2032
rect 3068 1992 3608 2020
rect 1213 1955 1271 1961
rect 1213 1921 1225 1955
rect 1259 1952 1271 1955
rect 1486 1952 1492 1964
rect 1259 1924 1492 1952
rect 1259 1921 1271 1924
rect 1213 1915 1271 1921
rect 1486 1912 1492 1924
rect 1544 1912 1550 1964
rect 1394 1844 1400 1896
rect 1452 1844 1458 1896
rect 2958 1844 2964 1896
rect 3016 1884 3022 1896
rect 3068 1893 3096 1992
rect 3602 1980 3608 1992
rect 3660 1980 3666 2032
rect 3326 1912 3332 1964
rect 3384 1952 3390 1964
rect 3804 1952 3832 2060
rect 4724 2020 4752 2060
rect 5166 2048 5172 2100
rect 5224 2048 5230 2100
rect 6914 2048 6920 2100
rect 6972 2048 6978 2100
rect 7098 2048 7104 2100
rect 7156 2048 7162 2100
rect 8110 2088 8116 2100
rect 7484 2060 8116 2088
rect 6549 2023 6607 2029
rect 6549 2020 6561 2023
rect 4724 1992 6561 2020
rect 6549 1989 6561 1992
rect 6595 2020 6607 2023
rect 7006 2020 7012 2032
rect 6595 1992 7012 2020
rect 6595 1989 6607 1992
rect 6549 1983 6607 1989
rect 7006 1980 7012 1992
rect 7064 1980 7070 2032
rect 7484 1961 7512 2060
rect 8110 2048 8116 2060
rect 8168 2048 8174 2100
rect 8754 2048 8760 2100
rect 8812 2048 8818 2100
rect 8941 2091 8999 2097
rect 8941 2057 8953 2091
rect 8987 2088 8999 2091
rect 9858 2088 9864 2100
rect 8987 2060 9864 2088
rect 8987 2057 8999 2060
rect 8941 2051 8999 2057
rect 9858 2048 9864 2060
rect 9916 2048 9922 2100
rect 8021 2023 8079 2029
rect 8021 1989 8033 2023
rect 8067 2020 8079 2023
rect 9490 2020 9496 2032
rect 8067 1992 9496 2020
rect 8067 1989 8079 1992
rect 8021 1983 8079 1989
rect 9490 1980 9496 1992
rect 9548 1980 9554 2032
rect 3384 1924 3832 1952
rect 7469 1955 7527 1961
rect 3384 1912 3390 1924
rect 7469 1921 7481 1955
rect 7515 1921 7527 1955
rect 7469 1915 7527 1921
rect 7558 1912 7564 1964
rect 7616 1912 7622 1964
rect 7742 1912 7748 1964
rect 7800 1912 7806 1964
rect 7852 1924 8156 1952
rect 3053 1887 3111 1893
rect 3053 1884 3065 1887
rect 3016 1856 3065 1884
rect 3016 1844 3022 1856
rect 3053 1853 3065 1856
rect 3099 1853 3111 1887
rect 3053 1847 3111 1853
rect 2808 1819 2866 1825
rect 2808 1785 2820 1819
rect 2854 1816 2866 1819
rect 3142 1816 3148 1828
rect 2854 1788 3148 1816
rect 2854 1785 2866 1788
rect 2808 1779 2866 1785
rect 3142 1776 3148 1788
rect 3200 1776 3206 1828
rect 3344 1825 3372 1912
rect 3602 1844 3608 1896
rect 3660 1884 3666 1896
rect 3789 1887 3847 1893
rect 3789 1884 3801 1887
rect 3660 1856 3801 1884
rect 3660 1844 3666 1856
rect 3789 1853 3801 1856
rect 3835 1884 3847 1887
rect 3835 1856 4200 1884
rect 3835 1853 3847 1856
rect 3789 1847 3847 1853
rect 3329 1819 3387 1825
rect 3329 1785 3341 1819
rect 3375 1785 3387 1819
rect 3329 1779 3387 1785
rect 3510 1776 3516 1828
rect 3568 1776 3574 1828
rect 4062 1825 4068 1828
rect 4056 1816 4068 1825
rect 4023 1788 4068 1816
rect 4056 1779 4068 1788
rect 4062 1776 4068 1779
rect 4120 1776 4126 1828
rect 4172 1816 4200 1856
rect 7190 1844 7196 1896
rect 7248 1884 7254 1896
rect 7653 1887 7711 1893
rect 7653 1884 7665 1887
rect 7248 1856 7665 1884
rect 7248 1844 7254 1856
rect 7653 1853 7665 1856
rect 7699 1884 7711 1887
rect 7852 1884 7880 1924
rect 7699 1856 7880 1884
rect 7699 1853 7711 1856
rect 7653 1847 7711 1853
rect 7926 1844 7932 1896
rect 7984 1844 7990 1896
rect 8128 1893 8156 1924
rect 8113 1887 8171 1893
rect 8113 1853 8125 1887
rect 8159 1884 8171 1887
rect 8573 1887 8631 1893
rect 8573 1884 8585 1887
rect 8159 1856 8585 1884
rect 8159 1853 8171 1856
rect 8113 1847 8171 1853
rect 8573 1853 8585 1856
rect 8619 1853 8631 1887
rect 8573 1847 8631 1853
rect 9033 1887 9091 1893
rect 9033 1853 9045 1887
rect 9079 1884 9091 1887
rect 9122 1884 9128 1896
rect 9079 1856 9128 1884
rect 9079 1853 9091 1856
rect 9033 1847 9091 1853
rect 9122 1844 9128 1856
rect 9180 1844 9186 1896
rect 4246 1816 4252 1828
rect 4172 1788 4252 1816
rect 4246 1776 4252 1788
rect 4304 1776 4310 1828
rect 6917 1819 6975 1825
rect 6917 1785 6929 1819
rect 6963 1816 6975 1819
rect 7944 1816 7972 1844
rect 8389 1819 8447 1825
rect 8389 1816 8401 1819
rect 6963 1788 7328 1816
rect 7944 1788 8401 1816
rect 6963 1785 6975 1788
rect 6917 1779 6975 1785
rect 1673 1751 1731 1757
rect 1673 1717 1685 1751
rect 1719 1748 1731 1751
rect 2590 1748 2596 1760
rect 1719 1720 2596 1748
rect 1719 1717 1731 1720
rect 1673 1711 1731 1717
rect 2590 1708 2596 1720
rect 2648 1708 2654 1760
rect 3234 1708 3240 1760
rect 3292 1748 3298 1760
rect 3528 1748 3556 1776
rect 7300 1757 7328 1788
rect 8389 1785 8401 1788
rect 8435 1785 8447 1819
rect 8389 1779 8447 1785
rect 3292 1720 3556 1748
rect 7285 1751 7343 1757
rect 3292 1708 3298 1720
rect 7285 1717 7297 1751
rect 7331 1717 7343 1751
rect 7285 1711 7343 1717
rect 552 1658 11132 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 10722 1658
rect 10774 1606 10786 1658
rect 10838 1606 10850 1658
rect 10902 1606 10914 1658
rect 10966 1606 10978 1658
rect 11030 1606 11132 1658
rect 552 1584 11132 1606
rect 2314 1504 2320 1556
rect 2372 1544 2378 1556
rect 2777 1547 2835 1553
rect 2777 1544 2789 1547
rect 2372 1516 2789 1544
rect 2372 1504 2378 1516
rect 2777 1513 2789 1516
rect 2823 1513 2835 1547
rect 2777 1507 2835 1513
rect 2869 1547 2927 1553
rect 2869 1513 2881 1547
rect 2915 1544 2927 1547
rect 2958 1544 2964 1556
rect 2915 1516 2964 1544
rect 2915 1513 2927 1516
rect 2869 1507 2927 1513
rect 2958 1504 2964 1516
rect 3016 1504 3022 1556
rect 2225 1479 2283 1485
rect 2225 1445 2237 1479
rect 2271 1476 2283 1479
rect 3050 1476 3056 1488
rect 2271 1448 3056 1476
rect 2271 1445 2283 1448
rect 2225 1439 2283 1445
rect 3050 1436 3056 1448
rect 3108 1436 3114 1488
rect 3326 1476 3332 1488
rect 3160 1448 3332 1476
rect 2038 1368 2044 1420
rect 2096 1408 2102 1420
rect 2133 1411 2191 1417
rect 2133 1408 2145 1411
rect 2096 1380 2145 1408
rect 2096 1368 2102 1380
rect 2133 1377 2145 1380
rect 2179 1377 2191 1411
rect 2133 1371 2191 1377
rect 2314 1368 2320 1420
rect 2372 1368 2378 1420
rect 2593 1411 2651 1417
rect 2593 1377 2605 1411
rect 2639 1408 2651 1411
rect 3160 1408 3188 1448
rect 3326 1436 3332 1448
rect 3384 1436 3390 1488
rect 3510 1436 3516 1488
rect 3568 1476 3574 1488
rect 3568 1448 4108 1476
rect 3568 1436 3574 1448
rect 2639 1380 3188 1408
rect 2639 1377 2651 1380
rect 2593 1371 2651 1377
rect 3234 1368 3240 1420
rect 3292 1408 3298 1420
rect 3982 1411 4040 1417
rect 3982 1408 3994 1411
rect 3292 1380 3994 1408
rect 3292 1368 3298 1380
rect 3982 1377 3994 1380
rect 4028 1377 4040 1411
rect 4080 1408 4108 1448
rect 4154 1436 4160 1488
rect 4212 1476 4218 1488
rect 4525 1479 4583 1485
rect 4525 1476 4537 1479
rect 4212 1448 4537 1476
rect 4212 1436 4218 1448
rect 4525 1445 4537 1448
rect 4571 1445 4583 1479
rect 4525 1439 4583 1445
rect 4080 1380 4384 1408
rect 3982 1371 4040 1377
rect 1946 1300 1952 1352
rect 2004 1340 2010 1352
rect 2409 1343 2467 1349
rect 2409 1340 2421 1343
rect 2004 1312 2421 1340
rect 2004 1300 2010 1312
rect 2409 1309 2421 1312
rect 2455 1309 2467 1343
rect 2409 1303 2467 1309
rect 2424 1204 2452 1303
rect 4246 1300 4252 1352
rect 4304 1300 4310 1352
rect 4356 1349 4384 1380
rect 4341 1343 4399 1349
rect 4341 1309 4353 1343
rect 4387 1340 4399 1343
rect 4798 1340 4804 1352
rect 4387 1312 4804 1340
rect 4387 1309 4399 1312
rect 4341 1303 4399 1309
rect 4798 1300 4804 1312
rect 4856 1300 4862 1352
rect 3510 1204 3516 1216
rect 2424 1176 3516 1204
rect 3510 1164 3516 1176
rect 3568 1164 3574 1216
rect 552 1114 11132 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 10062 1114
rect 10114 1062 10126 1114
rect 10178 1062 10190 1114
rect 10242 1062 10254 1114
rect 10306 1062 10318 1114
rect 10370 1062 11132 1114
rect 552 1040 11132 1062
rect 3234 960 3240 1012
rect 3292 960 3298 1012
rect 3418 960 3424 1012
rect 3476 960 3482 1012
rect 2774 756 2780 808
rect 2832 796 2838 808
rect 2832 768 3648 796
rect 2832 756 2838 768
rect 3050 688 3056 740
rect 3108 728 3114 740
rect 3620 737 3648 768
rect 3389 731 3447 737
rect 3389 728 3401 731
rect 3108 700 3401 728
rect 3108 688 3114 700
rect 3389 697 3401 700
rect 3435 697 3447 731
rect 3389 691 3447 697
rect 3605 731 3663 737
rect 3605 697 3617 731
rect 3651 697 3663 731
rect 3605 691 3663 697
rect 552 570 11132 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 10722 570
rect 10774 518 10786 570
rect 10838 518 10850 570
rect 10902 518 10914 570
rect 10966 518 10978 570
rect 11030 518 11132 570
rect 552 496 11132 518
<< via1 >>
rect 5816 43596 5868 43648
rect 10508 43596 10560 43648
rect 4322 42950 4374 43002
rect 4386 42950 4438 43002
rect 4450 42950 4502 43002
rect 4514 42950 4566 43002
rect 4578 42950 4630 43002
rect 10722 42950 10774 43002
rect 10786 42950 10838 43002
rect 10850 42950 10902 43002
rect 10914 42950 10966 43002
rect 10978 42950 11030 43002
rect 1768 42891 1820 42900
rect 1768 42857 1777 42891
rect 1777 42857 1811 42891
rect 1811 42857 1820 42891
rect 1768 42848 1820 42857
rect 2136 42848 2188 42900
rect 5632 42780 5684 42832
rect 6644 42780 6696 42832
rect 2320 42712 2372 42764
rect 3056 42755 3108 42764
rect 3056 42721 3065 42755
rect 3065 42721 3099 42755
rect 3099 42721 3108 42755
rect 3056 42712 3108 42721
rect 3884 42712 3936 42764
rect 2044 42687 2096 42696
rect 2044 42653 2053 42687
rect 2053 42653 2087 42687
rect 2087 42653 2096 42687
rect 2044 42644 2096 42653
rect 1584 42508 1636 42560
rect 2136 42576 2188 42628
rect 4252 42687 4304 42696
rect 4252 42653 4261 42687
rect 4261 42653 4295 42687
rect 4295 42653 4304 42687
rect 4252 42644 4304 42653
rect 4712 42644 4764 42696
rect 6184 42755 6236 42764
rect 6184 42721 6193 42755
rect 6193 42721 6227 42755
rect 6227 42721 6236 42755
rect 6184 42712 6236 42721
rect 7196 42712 7248 42764
rect 8392 42755 8444 42764
rect 8392 42721 8401 42755
rect 8401 42721 8435 42755
rect 8435 42721 8444 42755
rect 8392 42712 8444 42721
rect 8484 42712 8536 42764
rect 8668 42755 8720 42764
rect 8668 42721 8677 42755
rect 8677 42721 8711 42755
rect 8711 42721 8720 42755
rect 8668 42712 8720 42721
rect 8852 42712 8904 42764
rect 10324 42780 10376 42832
rect 9220 42755 9272 42764
rect 9220 42721 9229 42755
rect 9229 42721 9263 42755
rect 9263 42721 9272 42755
rect 9220 42712 9272 42721
rect 10508 42780 10560 42832
rect 4344 42576 4396 42628
rect 4804 42576 4856 42628
rect 5816 42619 5868 42628
rect 5816 42585 5825 42619
rect 5825 42585 5859 42619
rect 5859 42585 5868 42619
rect 5816 42576 5868 42585
rect 6184 42576 6236 42628
rect 7012 42644 7064 42696
rect 7748 42644 7800 42696
rect 10600 42712 10652 42764
rect 7656 42576 7708 42628
rect 9772 42576 9824 42628
rect 2504 42508 2556 42560
rect 4896 42551 4948 42560
rect 4896 42517 4905 42551
rect 4905 42517 4939 42551
rect 4939 42517 4948 42551
rect 4896 42508 4948 42517
rect 5356 42508 5408 42560
rect 9036 42508 9088 42560
rect 3662 42406 3714 42458
rect 3726 42406 3778 42458
rect 3790 42406 3842 42458
rect 3854 42406 3906 42458
rect 3918 42406 3970 42458
rect 10062 42406 10114 42458
rect 10126 42406 10178 42458
rect 10190 42406 10242 42458
rect 10254 42406 10306 42458
rect 10318 42406 10370 42458
rect 6552 42304 6604 42356
rect 8392 42304 8444 42356
rect 8668 42304 8720 42356
rect 9128 42304 9180 42356
rect 2964 42168 3016 42220
rect 6092 42211 6144 42220
rect 6092 42177 6101 42211
rect 6101 42177 6135 42211
rect 6135 42177 6144 42211
rect 6092 42168 6144 42177
rect 10508 42236 10560 42288
rect 7656 42168 7708 42220
rect 8116 42168 8168 42220
rect 1216 42143 1268 42152
rect 1216 42109 1225 42143
rect 1225 42109 1259 42143
rect 1259 42109 1268 42143
rect 1216 42100 1268 42109
rect 1400 42100 1452 42152
rect 1584 42143 1636 42152
rect 1584 42109 1618 42143
rect 1618 42109 1636 42143
rect 1584 42100 1636 42109
rect 2872 42100 2924 42152
rect 3700 42100 3752 42152
rect 4160 42032 4212 42084
rect 4896 42032 4948 42084
rect 572 41964 624 42016
rect 2780 41964 2832 42016
rect 3056 41964 3108 42016
rect 4344 41964 4396 42016
rect 5080 42007 5132 42016
rect 5080 41973 5089 42007
rect 5089 41973 5123 42007
rect 5123 41973 5132 42007
rect 5080 41964 5132 41973
rect 6000 42100 6052 42152
rect 5724 42032 5776 42084
rect 7380 42143 7432 42152
rect 7380 42109 7389 42143
rect 7389 42109 7423 42143
rect 7423 42109 7432 42143
rect 7380 42100 7432 42109
rect 8392 42143 8444 42152
rect 8392 42109 8401 42143
rect 8401 42109 8435 42143
rect 8435 42109 8444 42143
rect 8392 42100 8444 42109
rect 9680 42168 9732 42220
rect 10600 42211 10652 42220
rect 10600 42177 10609 42211
rect 10609 42177 10643 42211
rect 10643 42177 10652 42211
rect 10600 42168 10652 42177
rect 7564 42032 7616 42084
rect 7748 42075 7800 42084
rect 7748 42041 7757 42075
rect 7757 42041 7791 42075
rect 7791 42041 7800 42075
rect 7748 42032 7800 42041
rect 6460 41964 6512 42016
rect 8208 42007 8260 42016
rect 8208 41973 8217 42007
rect 8217 41973 8251 42007
rect 8251 41973 8260 42007
rect 8208 41964 8260 41973
rect 8668 42075 8720 42084
rect 8668 42041 8702 42075
rect 8702 42041 8720 42075
rect 8668 42032 8720 42041
rect 9772 41964 9824 42016
rect 9956 42007 10008 42016
rect 9956 41973 9965 42007
rect 9965 41973 9999 42007
rect 9999 41973 10008 42007
rect 9956 41964 10008 41973
rect 4322 41862 4374 41914
rect 4386 41862 4438 41914
rect 4450 41862 4502 41914
rect 4514 41862 4566 41914
rect 4578 41862 4630 41914
rect 10722 41862 10774 41914
rect 10786 41862 10838 41914
rect 10850 41862 10902 41914
rect 10914 41862 10966 41914
rect 10978 41862 11030 41914
rect 1124 41624 1176 41676
rect 1400 41692 1452 41744
rect 2228 41692 2280 41744
rect 3700 41760 3752 41812
rect 3332 41692 3384 41744
rect 756 41556 808 41608
rect 3240 41667 3292 41676
rect 3240 41633 3249 41667
rect 3249 41633 3283 41667
rect 3283 41633 3292 41667
rect 3240 41624 3292 41633
rect 3700 41667 3752 41676
rect 3700 41633 3709 41667
rect 3709 41633 3743 41667
rect 3743 41633 3752 41667
rect 3700 41624 3752 41633
rect 5356 41692 5408 41744
rect 8116 41760 8168 41812
rect 8392 41760 8444 41812
rect 9772 41760 9824 41812
rect 10692 41760 10744 41812
rect 6644 41692 6696 41744
rect 7656 41692 7708 41744
rect 5172 41624 5224 41676
rect 5724 41624 5776 41676
rect 6000 41667 6052 41676
rect 6000 41633 6009 41667
rect 6009 41633 6043 41667
rect 6043 41633 6052 41667
rect 6000 41624 6052 41633
rect 7380 41667 7432 41676
rect 7380 41633 7389 41667
rect 7389 41633 7423 41667
rect 7423 41633 7432 41667
rect 7380 41624 7432 41633
rect 7840 41624 7892 41676
rect 9036 41692 9088 41744
rect 9496 41692 9548 41744
rect 8392 41667 8444 41676
rect 8392 41633 8401 41667
rect 8401 41633 8435 41667
rect 8435 41633 8444 41667
rect 8392 41624 8444 41633
rect 9220 41624 9272 41676
rect 9772 41667 9824 41676
rect 11060 41692 11112 41744
rect 9772 41633 9790 41667
rect 9790 41633 9824 41667
rect 9772 41624 9824 41633
rect 10600 41667 10652 41676
rect 10600 41633 10609 41667
rect 10609 41633 10643 41667
rect 10643 41633 10652 41667
rect 10600 41624 10652 41633
rect 1032 41463 1084 41472
rect 1032 41429 1041 41463
rect 1041 41429 1075 41463
rect 1075 41429 1084 41463
rect 1032 41420 1084 41429
rect 1584 41420 1636 41472
rect 3424 41420 3476 41472
rect 6460 41488 6512 41540
rect 4804 41420 4856 41472
rect 5908 41463 5960 41472
rect 5908 41429 5917 41463
rect 5917 41429 5951 41463
rect 5951 41429 5960 41463
rect 5908 41420 5960 41429
rect 7656 41420 7708 41472
rect 8760 41488 8812 41540
rect 8576 41463 8628 41472
rect 8576 41429 8585 41463
rect 8585 41429 8619 41463
rect 8619 41429 8628 41463
rect 8576 41420 8628 41429
rect 9864 41420 9916 41472
rect 3662 41318 3714 41370
rect 3726 41318 3778 41370
rect 3790 41318 3842 41370
rect 3854 41318 3906 41370
rect 3918 41318 3970 41370
rect 10062 41318 10114 41370
rect 10126 41318 10178 41370
rect 10190 41318 10242 41370
rect 10254 41318 10306 41370
rect 10318 41318 10370 41370
rect 4712 41216 4764 41268
rect 204 41148 256 41200
rect 1492 41148 1544 41200
rect 1676 41148 1728 41200
rect 2688 41148 2740 41200
rect 4896 41148 4948 41200
rect 8484 41216 8536 41268
rect 8852 41216 8904 41268
rect 9036 41216 9088 41268
rect 9680 41216 9732 41268
rect 6736 41148 6788 41200
rect 3516 41080 3568 41132
rect 6092 41123 6144 41132
rect 6092 41089 6101 41123
rect 6101 41089 6135 41123
rect 6135 41089 6144 41123
rect 6092 41080 6144 41089
rect 8576 41148 8628 41200
rect 1584 41055 1636 41064
rect 1584 41021 1593 41055
rect 1593 41021 1627 41055
rect 1627 41021 1636 41055
rect 1584 41012 1636 41021
rect 2228 41012 2280 41064
rect 2780 41012 2832 41064
rect 4988 41012 5040 41064
rect 5908 41055 5960 41064
rect 5908 41021 5917 41055
rect 5917 41021 5951 41055
rect 5951 41021 5960 41055
rect 5908 41012 5960 41021
rect 8300 41012 8352 41064
rect 8392 41012 8444 41064
rect 8576 41055 8628 41064
rect 8576 41021 8585 41055
rect 8585 41021 8619 41055
rect 8619 41021 8628 41055
rect 8576 41012 8628 41021
rect 8760 41055 8812 41064
rect 8760 41021 8769 41055
rect 8769 41021 8803 41055
rect 8803 41021 8812 41055
rect 8760 41012 8812 41021
rect 8852 41055 8904 41064
rect 8852 41021 8861 41055
rect 8861 41021 8895 41055
rect 8895 41021 8904 41055
rect 8852 41012 8904 41021
rect 9220 41012 9272 41064
rect 9404 41012 9456 41064
rect 388 40876 440 40928
rect 664 40876 716 40928
rect 1492 40944 1544 40996
rect 1768 40944 1820 40996
rect 2044 40876 2096 40928
rect 4068 40944 4120 40996
rect 7932 40987 7984 40996
rect 7932 40953 7950 40987
rect 7950 40953 7984 40987
rect 7932 40944 7984 40953
rect 10140 40944 10192 40996
rect 4896 40876 4948 40928
rect 4988 40876 5040 40928
rect 5172 40876 5224 40928
rect 5264 40919 5316 40928
rect 5264 40885 5273 40919
rect 5273 40885 5307 40919
rect 5307 40885 5316 40919
rect 5264 40876 5316 40885
rect 5356 40876 5408 40928
rect 6552 40876 6604 40928
rect 6644 40919 6696 40928
rect 6644 40885 6653 40919
rect 6653 40885 6687 40919
rect 6687 40885 6696 40919
rect 6644 40876 6696 40885
rect 10324 40876 10376 40928
rect 10692 40919 10744 40928
rect 10692 40885 10701 40919
rect 10701 40885 10735 40919
rect 10735 40885 10744 40919
rect 10692 40876 10744 40885
rect 4322 40774 4374 40826
rect 4386 40774 4438 40826
rect 4450 40774 4502 40826
rect 4514 40774 4566 40826
rect 4578 40774 4630 40826
rect 10722 40774 10774 40826
rect 10786 40774 10838 40826
rect 10850 40774 10902 40826
rect 10914 40774 10966 40826
rect 10978 40774 11030 40826
rect 664 40672 716 40724
rect 3240 40672 3292 40724
rect 5080 40672 5132 40724
rect 6092 40672 6144 40724
rect 6552 40672 6604 40724
rect 7840 40672 7892 40724
rect 7932 40715 7984 40724
rect 7932 40681 7941 40715
rect 7941 40681 7975 40715
rect 7975 40681 7984 40715
rect 7932 40672 7984 40681
rect 1308 40536 1360 40588
rect 1492 40579 1544 40588
rect 1492 40545 1501 40579
rect 1501 40545 1535 40579
rect 1535 40545 1544 40579
rect 1492 40536 1544 40545
rect 1676 40536 1728 40588
rect 3240 40536 3292 40588
rect 1400 40468 1452 40520
rect 3516 40468 3568 40520
rect 4988 40536 5040 40588
rect 5080 40536 5132 40588
rect 6184 40604 6236 40656
rect 8484 40672 8536 40724
rect 8668 40672 8720 40724
rect 8944 40672 8996 40724
rect 9404 40672 9456 40724
rect 10140 40715 10192 40724
rect 10140 40681 10149 40715
rect 10149 40681 10183 40715
rect 10183 40681 10192 40715
rect 10140 40672 10192 40681
rect 8392 40647 8444 40656
rect 8392 40613 8401 40647
rect 8401 40613 8435 40647
rect 8435 40613 8444 40647
rect 8392 40604 8444 40613
rect 6736 40536 6788 40588
rect 8300 40536 8352 40588
rect 8484 40536 8536 40588
rect 8668 40579 8720 40588
rect 8668 40545 8677 40579
rect 8677 40545 8711 40579
rect 8711 40545 8720 40579
rect 8668 40536 8720 40545
rect 8944 40579 8996 40588
rect 8944 40545 8978 40579
rect 8978 40545 8996 40579
rect 8944 40536 8996 40545
rect 9128 40604 9180 40656
rect 10140 40536 10192 40588
rect 4528 40511 4580 40520
rect 4528 40477 4537 40511
rect 4537 40477 4571 40511
rect 4571 40477 4580 40511
rect 4528 40468 4580 40477
rect 4804 40468 4856 40520
rect 4896 40511 4948 40520
rect 4896 40477 4905 40511
rect 4905 40477 4939 40511
rect 4939 40477 4948 40511
rect 4896 40468 4948 40477
rect 5816 40468 5868 40520
rect 2596 40400 2648 40452
rect 2872 40400 2924 40452
rect 5632 40400 5684 40452
rect 940 40375 992 40384
rect 940 40341 949 40375
rect 949 40341 983 40375
rect 983 40341 992 40375
rect 940 40332 992 40341
rect 1308 40375 1360 40384
rect 1308 40341 1317 40375
rect 1317 40341 1351 40375
rect 1351 40341 1360 40375
rect 1308 40332 1360 40341
rect 1860 40332 1912 40384
rect 3056 40332 3108 40384
rect 4620 40332 4672 40384
rect 8392 40468 8444 40520
rect 9680 40468 9732 40520
rect 10324 40536 10376 40588
rect 10692 40536 10744 40588
rect 10416 40400 10468 40452
rect 8024 40332 8076 40384
rect 8576 40332 8628 40384
rect 9036 40332 9088 40384
rect 9588 40332 9640 40384
rect 10140 40332 10192 40384
rect 10508 40332 10560 40384
rect 3662 40230 3714 40282
rect 3726 40230 3778 40282
rect 3790 40230 3842 40282
rect 3854 40230 3906 40282
rect 3918 40230 3970 40282
rect 10062 40230 10114 40282
rect 10126 40230 10178 40282
rect 10190 40230 10242 40282
rect 10254 40230 10306 40282
rect 10318 40230 10370 40282
rect 2596 40128 2648 40180
rect 3056 40128 3108 40180
rect 3700 40128 3752 40180
rect 4068 40128 4120 40180
rect 4896 40128 4948 40180
rect 8208 40128 8260 40180
rect 8300 40128 8352 40180
rect 8852 40128 8904 40180
rect 9404 40128 9456 40180
rect 2044 40060 2096 40112
rect 3240 40060 3292 40112
rect 1584 39924 1636 39976
rect 1860 39967 1912 39976
rect 1860 39933 1869 39967
rect 1869 39933 1903 39967
rect 1903 39933 1912 39967
rect 1860 39924 1912 39933
rect 1952 39967 2004 39976
rect 1952 39933 1961 39967
rect 1961 39933 1995 39967
rect 1995 39933 2004 39967
rect 1952 39924 2004 39933
rect 2044 39967 2096 39976
rect 2044 39933 2053 39967
rect 2053 39933 2087 39967
rect 2087 39933 2096 39967
rect 2044 39924 2096 39933
rect 2320 39967 2372 39976
rect 2320 39933 2329 39967
rect 2329 39933 2363 39967
rect 2363 39933 2372 39967
rect 2320 39924 2372 39933
rect 2872 40035 2924 40044
rect 2872 40001 2881 40035
rect 2881 40001 2915 40035
rect 2915 40001 2924 40035
rect 2872 39992 2924 40001
rect 3424 40035 3476 40044
rect 3424 40001 3433 40035
rect 3433 40001 3467 40035
rect 3467 40001 3476 40035
rect 3424 39992 3476 40001
rect 3332 39924 3384 39976
rect 4620 40035 4672 40044
rect 4620 40001 4629 40035
rect 4629 40001 4663 40035
rect 4663 40001 4672 40035
rect 4620 39992 4672 40001
rect 8024 40060 8076 40112
rect 2688 39856 2740 39908
rect 2964 39856 3016 39908
rect 3056 39856 3108 39908
rect 5172 39967 5224 39976
rect 5172 39933 5181 39967
rect 5181 39933 5215 39967
rect 5215 39933 5224 39967
rect 5172 39924 5224 39933
rect 5448 39967 5500 39976
rect 5448 39933 5457 39967
rect 5457 39933 5491 39967
rect 5491 39933 5500 39967
rect 5448 39924 5500 39933
rect 8576 39992 8628 40044
rect 11244 40060 11296 40112
rect 4528 39788 4580 39840
rect 4712 39788 4764 39840
rect 5080 39899 5132 39908
rect 5080 39865 5089 39899
rect 5089 39865 5123 39899
rect 5123 39865 5132 39899
rect 5080 39856 5132 39865
rect 7840 39924 7892 39976
rect 8392 39967 8444 39976
rect 8392 39933 8401 39967
rect 8401 39933 8435 39967
rect 8435 39933 8444 39967
rect 8392 39924 8444 39933
rect 10048 40035 10100 40044
rect 10048 40001 10057 40035
rect 10057 40001 10091 40035
rect 10091 40001 10100 40035
rect 10048 39992 10100 40001
rect 11060 39992 11112 40044
rect 5356 39831 5408 39840
rect 5356 39797 5365 39831
rect 5365 39797 5399 39831
rect 5399 39797 5408 39831
rect 5356 39788 5408 39797
rect 5540 39831 5592 39840
rect 5540 39797 5549 39831
rect 5549 39797 5583 39831
rect 5583 39797 5592 39831
rect 5540 39788 5592 39797
rect 6460 39856 6512 39908
rect 6644 39856 6696 39908
rect 8668 39899 8720 39908
rect 8668 39865 8677 39899
rect 8677 39865 8711 39899
rect 8711 39865 8720 39899
rect 8668 39856 8720 39865
rect 8760 39899 8812 39908
rect 8760 39865 8769 39899
rect 8769 39865 8803 39899
rect 8803 39865 8812 39899
rect 8760 39856 8812 39865
rect 7012 39788 7064 39840
rect 7104 39788 7156 39840
rect 8116 39831 8168 39840
rect 8116 39797 8125 39831
rect 8125 39797 8159 39831
rect 8159 39797 8168 39831
rect 8116 39788 8168 39797
rect 8484 39831 8536 39840
rect 8484 39797 8493 39831
rect 8493 39797 8527 39831
rect 8527 39797 8536 39831
rect 8484 39788 8536 39797
rect 8576 39788 8628 39840
rect 8944 39788 8996 39840
rect 9864 39856 9916 39908
rect 10600 39924 10652 39976
rect 10416 39899 10468 39908
rect 10416 39865 10425 39899
rect 10425 39865 10459 39899
rect 10459 39865 10468 39899
rect 10416 39856 10468 39865
rect 10692 39899 10744 39908
rect 10692 39865 10701 39899
rect 10701 39865 10735 39899
rect 10735 39865 10744 39899
rect 10692 39856 10744 39865
rect 11152 39856 11204 39908
rect 9956 39831 10008 39840
rect 9956 39797 9965 39831
rect 9965 39797 9999 39831
rect 9999 39797 10008 39831
rect 9956 39788 10008 39797
rect 10232 39788 10284 39840
rect 4322 39686 4374 39738
rect 4386 39686 4438 39738
rect 4450 39686 4502 39738
rect 4514 39686 4566 39738
rect 4578 39686 4630 39738
rect 10722 39686 10774 39738
rect 10786 39686 10838 39738
rect 10850 39686 10902 39738
rect 10914 39686 10966 39738
rect 10978 39686 11030 39738
rect 1584 39584 1636 39636
rect 1676 39627 1728 39636
rect 1676 39593 1685 39627
rect 1685 39593 1719 39627
rect 1719 39593 1728 39627
rect 1676 39584 1728 39593
rect 4160 39627 4212 39636
rect 4160 39593 4169 39627
rect 4169 39593 4203 39627
rect 4203 39593 4212 39627
rect 4160 39584 4212 39593
rect 4712 39584 4764 39636
rect 6552 39584 6604 39636
rect 6644 39627 6696 39636
rect 6644 39593 6653 39627
rect 6653 39593 6687 39627
rect 6687 39593 6696 39627
rect 6644 39584 6696 39593
rect 7104 39627 7156 39636
rect 7104 39593 7113 39627
rect 7113 39593 7147 39627
rect 7147 39593 7156 39627
rect 7104 39584 7156 39593
rect 7380 39584 7432 39636
rect 8944 39584 8996 39636
rect 9588 39584 9640 39636
rect 1952 39516 2004 39568
rect 2044 39516 2096 39568
rect 3148 39516 3200 39568
rect 3608 39516 3660 39568
rect 5448 39516 5500 39568
rect 572 39448 624 39500
rect 1584 39491 1636 39500
rect 1584 39457 1593 39491
rect 1593 39457 1627 39491
rect 1627 39457 1636 39491
rect 1584 39448 1636 39457
rect 2412 39491 2464 39500
rect 2412 39457 2446 39491
rect 2446 39457 2464 39491
rect 2412 39448 2464 39457
rect 1492 39380 1544 39432
rect 1676 39312 1728 39364
rect 1124 39287 1176 39296
rect 1124 39253 1133 39287
rect 1133 39253 1167 39287
rect 1167 39253 1176 39287
rect 1124 39244 1176 39253
rect 1860 39287 1912 39296
rect 1860 39253 1869 39287
rect 1869 39253 1903 39287
rect 1903 39253 1912 39287
rect 1860 39244 1912 39253
rect 3332 39244 3384 39296
rect 5080 39448 5132 39500
rect 4068 39380 4120 39432
rect 4804 39423 4856 39432
rect 4804 39389 4813 39423
rect 4813 39389 4847 39423
rect 4847 39389 4856 39423
rect 4804 39380 4856 39389
rect 4896 39380 4948 39432
rect 5264 39380 5316 39432
rect 5632 39423 5684 39432
rect 5632 39389 5641 39423
rect 5641 39389 5675 39423
rect 5675 39389 5684 39423
rect 5632 39380 5684 39389
rect 5816 39491 5868 39500
rect 5816 39457 5825 39491
rect 5825 39457 5859 39491
rect 5859 39457 5868 39491
rect 5816 39448 5868 39457
rect 9772 39584 9824 39636
rect 11060 39584 11112 39636
rect 6092 39448 6144 39500
rect 6460 39491 6512 39500
rect 6460 39457 6469 39491
rect 6469 39457 6503 39491
rect 6503 39457 6512 39491
rect 6460 39448 6512 39457
rect 7104 39448 7156 39500
rect 7472 39491 7524 39500
rect 7472 39457 7481 39491
rect 7481 39457 7515 39491
rect 7515 39457 7524 39491
rect 7472 39448 7524 39457
rect 7564 39448 7616 39500
rect 7748 39448 7800 39500
rect 7196 39380 7248 39432
rect 7288 39423 7340 39432
rect 7288 39389 7297 39423
rect 7297 39389 7331 39423
rect 7331 39389 7340 39423
rect 7288 39380 7340 39389
rect 6920 39312 6972 39364
rect 5724 39244 5776 39296
rect 8208 39448 8260 39500
rect 8944 39491 8996 39500
rect 8944 39457 8953 39491
rect 8953 39457 8987 39491
rect 8987 39457 8996 39491
rect 8944 39448 8996 39457
rect 9036 39448 9088 39500
rect 9956 39448 10008 39500
rect 8484 39380 8536 39432
rect 9404 39423 9456 39432
rect 9404 39389 9413 39423
rect 9413 39389 9447 39423
rect 9447 39389 9456 39423
rect 9404 39380 9456 39389
rect 8668 39287 8720 39296
rect 8668 39253 8677 39287
rect 8677 39253 8711 39287
rect 8711 39253 8720 39287
rect 8668 39244 8720 39253
rect 8852 39244 8904 39296
rect 9680 39244 9732 39296
rect 10048 39244 10100 39296
rect 3662 39142 3714 39194
rect 3726 39142 3778 39194
rect 3790 39142 3842 39194
rect 3854 39142 3906 39194
rect 3918 39142 3970 39194
rect 10062 39142 10114 39194
rect 10126 39142 10178 39194
rect 10190 39142 10242 39194
rect 10254 39142 10306 39194
rect 10318 39142 10370 39194
rect 664 39040 716 39092
rect 1860 39040 1912 39092
rect 3700 39040 3752 39092
rect 5080 39040 5132 39092
rect 5724 39083 5776 39092
rect 5724 39049 5733 39083
rect 5733 39049 5767 39083
rect 5767 39049 5776 39083
rect 5724 39040 5776 39049
rect 5908 39040 5960 39092
rect 6828 39083 6880 39092
rect 6828 39049 6837 39083
rect 6837 39049 6871 39083
rect 6871 39049 6880 39083
rect 6828 39040 6880 39049
rect 7288 39040 7340 39092
rect 8300 39040 8352 39092
rect 8392 39040 8444 39092
rect 1400 39015 1452 39024
rect 1400 38981 1409 39015
rect 1409 38981 1443 39015
rect 1443 38981 1452 39015
rect 1400 38972 1452 38981
rect 3056 39015 3108 39024
rect 3056 38981 3065 39015
rect 3065 38981 3099 39015
rect 3099 38981 3108 39015
rect 3056 38972 3108 38981
rect 5632 38972 5684 39024
rect 6644 38972 6696 39024
rect 6736 38972 6788 39024
rect 1308 38904 1360 38956
rect 1492 38904 1544 38956
rect 8208 38972 8260 39024
rect 1032 38879 1084 38888
rect 1032 38845 1041 38879
rect 1041 38845 1075 38879
rect 1075 38845 1084 38879
rect 1032 38836 1084 38845
rect 7196 38904 7248 38956
rect 8392 38904 8444 38956
rect 1124 38811 1176 38820
rect 1124 38777 1133 38811
rect 1133 38777 1167 38811
rect 1167 38777 1176 38811
rect 1124 38768 1176 38777
rect 1676 38700 1728 38752
rect 3884 38836 3936 38888
rect 4160 38768 4212 38820
rect 5908 38836 5960 38888
rect 6736 38836 6788 38888
rect 7288 38836 7340 38888
rect 6828 38768 6880 38820
rect 7472 38879 7524 38888
rect 7472 38845 7481 38879
rect 7481 38845 7515 38879
rect 7515 38845 7524 38879
rect 7472 38836 7524 38845
rect 7564 38836 7616 38888
rect 7748 38879 7800 38888
rect 7748 38845 7757 38879
rect 7757 38845 7791 38879
rect 7791 38845 7800 38879
rect 7748 38836 7800 38845
rect 7932 38879 7984 38888
rect 7932 38845 7941 38879
rect 7941 38845 7975 38879
rect 7975 38845 7984 38879
rect 7932 38836 7984 38845
rect 8208 38836 8260 38888
rect 8300 38836 8352 38888
rect 9588 39040 9640 39092
rect 9772 39083 9824 39092
rect 9772 39049 9781 39083
rect 9781 39049 9815 39083
rect 9815 39049 9824 39083
rect 9772 39040 9824 39049
rect 8944 38972 8996 39024
rect 9956 38972 10008 39024
rect 8852 38879 8904 38888
rect 8852 38845 8861 38879
rect 8861 38845 8895 38879
rect 8895 38845 8904 38879
rect 8852 38836 8904 38845
rect 8944 38879 8996 38888
rect 8944 38845 8953 38879
rect 8953 38845 8987 38879
rect 8987 38845 8996 38879
rect 8944 38836 8996 38845
rect 9588 38904 9640 38956
rect 9864 38836 9916 38888
rect 10140 38879 10192 38888
rect 10140 38845 10149 38879
rect 10149 38845 10183 38879
rect 10183 38845 10192 38879
rect 10140 38836 10192 38845
rect 9680 38768 9732 38820
rect 5908 38743 5960 38752
rect 5908 38709 5917 38743
rect 5917 38709 5951 38743
rect 5951 38709 5960 38743
rect 5908 38700 5960 38709
rect 7104 38700 7156 38752
rect 8300 38700 8352 38752
rect 8484 38700 8536 38752
rect 8668 38700 8720 38752
rect 9312 38700 9364 38752
rect 10232 38743 10284 38752
rect 10232 38709 10241 38743
rect 10241 38709 10275 38743
rect 10275 38709 10284 38743
rect 10232 38700 10284 38709
rect 10416 38700 10468 38752
rect 4322 38598 4374 38650
rect 4386 38598 4438 38650
rect 4450 38598 4502 38650
rect 4514 38598 4566 38650
rect 4578 38598 4630 38650
rect 10722 38598 10774 38650
rect 10786 38598 10838 38650
rect 10850 38598 10902 38650
rect 10914 38598 10966 38650
rect 10978 38598 11030 38650
rect 756 38496 808 38548
rect 1768 38539 1820 38548
rect 1768 38505 1777 38539
rect 1777 38505 1811 38539
rect 1811 38505 1820 38539
rect 1768 38496 1820 38505
rect 1308 38360 1360 38412
rect 2412 38496 2464 38548
rect 3792 38496 3844 38548
rect 5356 38496 5408 38548
rect 2320 38428 2372 38480
rect 3240 38428 3292 38480
rect 3700 38471 3752 38480
rect 3700 38437 3709 38471
rect 3709 38437 3743 38471
rect 3743 38437 3752 38471
rect 3700 38428 3752 38437
rect 4068 38428 4120 38480
rect 5908 38496 5960 38548
rect 7472 38496 7524 38548
rect 7748 38496 7800 38548
rect 1952 38360 2004 38412
rect 388 38224 440 38276
rect 1492 38292 1544 38344
rect 3516 38360 3568 38412
rect 3792 38403 3844 38412
rect 3792 38369 3801 38403
rect 3801 38369 3835 38403
rect 3835 38369 3844 38403
rect 3792 38360 3844 38369
rect 4712 38360 4764 38412
rect 5632 38360 5684 38412
rect 7012 38360 7064 38412
rect 7380 38428 7432 38480
rect 8300 38428 8352 38480
rect 8944 38496 8996 38548
rect 9220 38496 9272 38548
rect 9864 38496 9916 38548
rect 7288 38360 7340 38412
rect 1124 38199 1176 38208
rect 1124 38165 1133 38199
rect 1133 38165 1167 38199
rect 1167 38165 1176 38199
rect 1124 38156 1176 38165
rect 1676 38224 1728 38276
rect 2964 38224 3016 38276
rect 4436 38224 4488 38276
rect 6276 38292 6328 38344
rect 6920 38335 6972 38344
rect 6920 38301 6929 38335
rect 6929 38301 6963 38335
rect 6963 38301 6972 38335
rect 6920 38292 6972 38301
rect 7104 38224 7156 38276
rect 7748 38403 7800 38412
rect 7748 38369 7757 38403
rect 7757 38369 7791 38403
rect 7791 38369 7800 38403
rect 7748 38360 7800 38369
rect 8024 38403 8076 38412
rect 8024 38369 8033 38403
rect 8033 38369 8067 38403
rect 8067 38369 8076 38403
rect 8024 38360 8076 38369
rect 8392 38403 8444 38412
rect 8392 38369 8401 38403
rect 8401 38369 8435 38403
rect 8435 38369 8444 38403
rect 8392 38360 8444 38369
rect 8944 38360 8996 38412
rect 9680 38428 9732 38480
rect 9312 38292 9364 38344
rect 9128 38224 9180 38276
rect 10508 38403 10560 38412
rect 10508 38369 10517 38403
rect 10517 38369 10551 38403
rect 10551 38369 10560 38403
rect 10508 38360 10560 38369
rect 10048 38292 10100 38344
rect 10508 38224 10560 38276
rect 2504 38156 2556 38208
rect 3516 38156 3568 38208
rect 4160 38156 4212 38208
rect 6736 38156 6788 38208
rect 7288 38156 7340 38208
rect 7472 38156 7524 38208
rect 7656 38156 7708 38208
rect 8116 38156 8168 38208
rect 9220 38156 9272 38208
rect 9772 38156 9824 38208
rect 9956 38199 10008 38208
rect 9956 38165 9965 38199
rect 9965 38165 9999 38199
rect 9999 38165 10008 38199
rect 9956 38156 10008 38165
rect 10232 38156 10284 38208
rect 10324 38156 10376 38208
rect 11060 38156 11112 38208
rect 3662 38054 3714 38106
rect 3726 38054 3778 38106
rect 3790 38054 3842 38106
rect 3854 38054 3906 38106
rect 3918 38054 3970 38106
rect 10062 38054 10114 38106
rect 10126 38054 10178 38106
rect 10190 38054 10242 38106
rect 10254 38054 10306 38106
rect 10318 38054 10370 38106
rect 848 37952 900 38004
rect 2136 37995 2188 38004
rect 2136 37961 2145 37995
rect 2145 37961 2179 37995
rect 2179 37961 2188 37995
rect 2136 37952 2188 37961
rect 2504 37995 2556 38004
rect 2504 37961 2513 37995
rect 2513 37961 2547 37995
rect 2547 37961 2556 37995
rect 2504 37952 2556 37961
rect 2964 37995 3016 38004
rect 2964 37961 2973 37995
rect 2973 37961 3007 37995
rect 3007 37961 3016 37995
rect 2964 37952 3016 37961
rect 3056 37952 3108 38004
rect 3332 37952 3384 38004
rect 3884 37952 3936 38004
rect 5632 37952 5684 38004
rect 1124 37884 1176 37936
rect 2412 37884 2464 37936
rect 3976 37884 4028 37936
rect 7564 37952 7616 38004
rect 3332 37816 3384 37868
rect 4804 37859 4856 37868
rect 4804 37825 4813 37859
rect 4813 37825 4847 37859
rect 4847 37825 4856 37859
rect 4804 37816 4856 37825
rect 6276 37816 6328 37868
rect 7748 37884 7800 37936
rect 7932 37952 7984 38004
rect 9128 37952 9180 38004
rect 9588 37995 9640 38004
rect 9588 37961 9597 37995
rect 9597 37961 9631 37995
rect 9631 37961 9640 37995
rect 9588 37952 9640 37961
rect 8116 37884 8168 37936
rect 7104 37816 7156 37868
rect 8576 37816 8628 37868
rect 112 37748 164 37800
rect 1584 37791 1636 37800
rect 1584 37757 1593 37791
rect 1593 37757 1627 37791
rect 1627 37757 1636 37791
rect 1584 37748 1636 37757
rect 1952 37791 2004 37800
rect 1952 37757 1961 37791
rect 1961 37757 1995 37791
rect 1995 37757 2004 37791
rect 1952 37748 2004 37757
rect 2320 37791 2372 37800
rect 2320 37757 2329 37791
rect 2329 37757 2363 37791
rect 2363 37757 2372 37791
rect 2320 37748 2372 37757
rect 1860 37680 1912 37732
rect 2136 37680 2188 37732
rect 3608 37791 3660 37800
rect 3608 37757 3617 37791
rect 3617 37757 3651 37791
rect 3651 37757 3660 37791
rect 3608 37748 3660 37757
rect 4252 37748 4304 37800
rect 4712 37748 4764 37800
rect 5448 37748 5500 37800
rect 5540 37791 5592 37800
rect 5540 37757 5549 37791
rect 5549 37757 5583 37791
rect 5583 37757 5592 37791
rect 5540 37748 5592 37757
rect 6092 37748 6144 37800
rect 6736 37791 6788 37800
rect 6736 37757 6745 37791
rect 6745 37757 6779 37791
rect 6779 37757 6788 37791
rect 6736 37748 6788 37757
rect 6828 37748 6880 37800
rect 2504 37680 2556 37732
rect 6184 37680 6236 37732
rect 6276 37680 6328 37732
rect 8392 37748 8444 37800
rect 1124 37612 1176 37664
rect 1676 37612 1728 37664
rect 3056 37612 3108 37664
rect 4252 37655 4304 37664
rect 4252 37621 4261 37655
rect 4261 37621 4295 37655
rect 4295 37621 4304 37655
rect 4252 37612 4304 37621
rect 4712 37655 4764 37664
rect 4712 37621 4721 37655
rect 4721 37621 4755 37655
rect 4755 37621 4764 37655
rect 4712 37612 4764 37621
rect 6736 37612 6788 37664
rect 10508 37884 10560 37936
rect 9864 37816 9916 37868
rect 9128 37791 9180 37800
rect 9128 37757 9137 37791
rect 9137 37757 9171 37791
rect 9171 37757 9180 37791
rect 9128 37748 9180 37757
rect 9404 37791 9456 37800
rect 9404 37757 9429 37791
rect 9429 37757 9456 37791
rect 9404 37748 9456 37757
rect 9956 37748 10008 37800
rect 10508 37748 10560 37800
rect 9864 37723 9916 37732
rect 9864 37689 9873 37723
rect 9873 37689 9907 37723
rect 9907 37689 9916 37723
rect 9864 37680 9916 37689
rect 10416 37680 10468 37732
rect 8668 37612 8720 37664
rect 8760 37612 8812 37664
rect 9312 37612 9364 37664
rect 9404 37612 9456 37664
rect 4322 37510 4374 37562
rect 4386 37510 4438 37562
rect 4450 37510 4502 37562
rect 4514 37510 4566 37562
rect 4578 37510 4630 37562
rect 10722 37510 10774 37562
rect 10786 37510 10838 37562
rect 10850 37510 10902 37562
rect 10914 37510 10966 37562
rect 10978 37510 11030 37562
rect 1032 37408 1084 37460
rect 3332 37408 3384 37460
rect 5816 37408 5868 37460
rect 6184 37408 6236 37460
rect 6920 37408 6972 37460
rect 7840 37408 7892 37460
rect 8208 37451 8260 37460
rect 8208 37417 8217 37451
rect 8217 37417 8251 37451
rect 8251 37417 8260 37451
rect 8208 37408 8260 37417
rect 8760 37408 8812 37460
rect 9128 37408 9180 37460
rect 1584 37340 1636 37392
rect 3424 37340 3476 37392
rect 1124 37315 1176 37324
rect 1124 37281 1133 37315
rect 1133 37281 1167 37315
rect 1167 37281 1176 37315
rect 1124 37272 1176 37281
rect 1492 37272 1544 37324
rect 1676 37315 1728 37324
rect 1676 37281 1710 37315
rect 1710 37281 1728 37315
rect 1676 37272 1728 37281
rect 2872 37272 2924 37324
rect 6092 37340 6144 37392
rect 7196 37340 7248 37392
rect 3884 37315 3936 37324
rect 3884 37281 3893 37315
rect 3893 37281 3927 37315
rect 3927 37281 3936 37315
rect 3884 37272 3936 37281
rect 3976 37315 4028 37324
rect 3976 37281 3985 37315
rect 3985 37281 4019 37315
rect 4019 37281 4028 37315
rect 3976 37272 4028 37281
rect 4160 37315 4212 37324
rect 4160 37281 4169 37315
rect 4169 37281 4203 37315
rect 4203 37281 4212 37315
rect 4160 37272 4212 37281
rect 5172 37272 5224 37324
rect 5264 37315 5316 37324
rect 5264 37281 5273 37315
rect 5273 37281 5307 37315
rect 5307 37281 5316 37315
rect 5264 37272 5316 37281
rect 5356 37315 5408 37324
rect 5356 37281 5365 37315
rect 5365 37281 5399 37315
rect 5399 37281 5408 37315
rect 5356 37272 5408 37281
rect 5448 37315 5500 37324
rect 5448 37281 5457 37315
rect 5457 37281 5491 37315
rect 5491 37281 5500 37315
rect 5448 37272 5500 37281
rect 5632 37315 5684 37324
rect 5632 37281 5641 37315
rect 5641 37281 5675 37315
rect 5675 37281 5684 37315
rect 5632 37272 5684 37281
rect 2688 37204 2740 37256
rect 3424 37247 3476 37256
rect 3424 37213 3433 37247
rect 3433 37213 3467 37247
rect 3467 37213 3476 37247
rect 3424 37204 3476 37213
rect 4804 37247 4856 37256
rect 4804 37213 4813 37247
rect 4813 37213 4847 37247
rect 4847 37213 4856 37247
rect 4804 37204 4856 37213
rect 5080 37204 5132 37256
rect 1768 37068 1820 37120
rect 5540 37136 5592 37188
rect 6276 37315 6328 37324
rect 6276 37281 6285 37315
rect 6285 37281 6319 37315
rect 6319 37281 6328 37315
rect 6276 37272 6328 37281
rect 6644 37272 6696 37324
rect 7380 37272 7432 37324
rect 7656 37315 7708 37324
rect 7656 37281 7665 37315
rect 7665 37281 7699 37315
rect 7699 37281 7708 37315
rect 7656 37272 7708 37281
rect 9220 37340 9272 37392
rect 6552 37204 6604 37256
rect 6920 37204 6972 37256
rect 7012 37136 7064 37188
rect 7380 37136 7432 37188
rect 8024 37204 8076 37256
rect 8392 37272 8444 37324
rect 8852 37272 8904 37324
rect 11060 37272 11112 37324
rect 4620 37068 4672 37120
rect 6460 37068 6512 37120
rect 8116 37136 8168 37188
rect 8300 37068 8352 37120
rect 8944 37136 8996 37188
rect 10508 37068 10560 37120
rect 3662 36966 3714 37018
rect 3726 36966 3778 37018
rect 3790 36966 3842 37018
rect 3854 36966 3906 37018
rect 3918 36966 3970 37018
rect 10062 36966 10114 37018
rect 10126 36966 10178 37018
rect 10190 36966 10242 37018
rect 10254 36966 10306 37018
rect 10318 36966 10370 37018
rect 1124 36864 1176 36916
rect 4712 36864 4764 36916
rect 1400 36728 1452 36780
rect 3332 36771 3384 36780
rect 3332 36737 3341 36771
rect 3341 36737 3375 36771
rect 3375 36737 3384 36771
rect 3332 36728 3384 36737
rect 1032 36660 1084 36712
rect 1768 36660 1820 36712
rect 4068 36660 4120 36712
rect 4252 36703 4304 36712
rect 4252 36669 4286 36703
rect 4286 36669 4304 36703
rect 4252 36660 4304 36669
rect 1308 36592 1360 36644
rect 2872 36635 2924 36644
rect 2872 36601 2881 36635
rect 2881 36601 2915 36635
rect 2915 36601 2924 36635
rect 2872 36592 2924 36601
rect 3516 36592 3568 36644
rect 5356 36660 5408 36712
rect 5908 36728 5960 36780
rect 5816 36703 5868 36712
rect 5816 36669 5825 36703
rect 5825 36669 5859 36703
rect 5859 36669 5868 36703
rect 5816 36660 5868 36669
rect 9128 36864 9180 36916
rect 9864 36864 9916 36916
rect 10324 36907 10376 36916
rect 10324 36873 10333 36907
rect 10333 36873 10367 36907
rect 10367 36873 10376 36907
rect 10324 36864 10376 36873
rect 7380 36796 7432 36848
rect 7932 36796 7984 36848
rect 9680 36796 9732 36848
rect 6092 36728 6144 36780
rect 6184 36703 6236 36712
rect 6184 36669 6193 36703
rect 6193 36669 6227 36703
rect 6227 36669 6236 36703
rect 6184 36660 6236 36669
rect 6552 36703 6604 36712
rect 6552 36669 6561 36703
rect 6561 36669 6595 36703
rect 6595 36669 6604 36703
rect 6552 36660 6604 36669
rect 7196 36660 7248 36712
rect 6644 36592 6696 36644
rect 7104 36592 7156 36644
rect 7932 36703 7984 36712
rect 7932 36669 7941 36703
rect 7941 36669 7975 36703
rect 7975 36669 7984 36703
rect 7932 36660 7984 36669
rect 10600 36796 10652 36848
rect 8392 36703 8444 36712
rect 8392 36669 8401 36703
rect 8401 36669 8435 36703
rect 8435 36669 8444 36703
rect 8392 36660 8444 36669
rect 8760 36660 8812 36712
rect 8668 36635 8720 36644
rect 8668 36601 8677 36635
rect 8677 36601 8711 36635
rect 8711 36601 8720 36635
rect 8668 36592 8720 36601
rect 9128 36703 9180 36712
rect 9128 36669 9137 36703
rect 9137 36669 9171 36703
rect 9171 36669 9180 36703
rect 9128 36660 9180 36669
rect 9312 36660 9364 36712
rect 3884 36567 3936 36576
rect 3884 36533 3893 36567
rect 3893 36533 3927 36567
rect 3927 36533 3936 36567
rect 3884 36524 3936 36533
rect 6920 36524 6972 36576
rect 7564 36524 7616 36576
rect 7748 36524 7800 36576
rect 8208 36567 8260 36576
rect 8208 36533 8217 36567
rect 8217 36533 8251 36567
rect 8251 36533 8260 36567
rect 8208 36524 8260 36533
rect 8300 36524 8352 36576
rect 9864 36635 9916 36644
rect 9864 36601 9873 36635
rect 9873 36601 9907 36635
rect 9907 36601 9916 36635
rect 9864 36592 9916 36601
rect 10140 36660 10192 36712
rect 11244 36728 11296 36780
rect 10692 36660 10744 36712
rect 10508 36635 10560 36644
rect 10508 36601 10517 36635
rect 10517 36601 10551 36635
rect 10551 36601 10560 36635
rect 10508 36592 10560 36601
rect 9220 36567 9272 36576
rect 9220 36533 9229 36567
rect 9229 36533 9263 36567
rect 9263 36533 9272 36567
rect 9220 36524 9272 36533
rect 9496 36524 9548 36576
rect 9680 36567 9732 36576
rect 9680 36533 9689 36567
rect 9689 36533 9723 36567
rect 9723 36533 9732 36567
rect 9680 36524 9732 36533
rect 9956 36524 10008 36576
rect 4322 36422 4374 36474
rect 4386 36422 4438 36474
rect 4450 36422 4502 36474
rect 4514 36422 4566 36474
rect 4578 36422 4630 36474
rect 10722 36422 10774 36474
rect 10786 36422 10838 36474
rect 10850 36422 10902 36474
rect 10914 36422 10966 36474
rect 10978 36422 11030 36474
rect 2688 36320 2740 36372
rect 1400 36252 1452 36304
rect 1768 36252 1820 36304
rect 3792 36363 3844 36372
rect 3792 36329 3801 36363
rect 3801 36329 3835 36363
rect 3835 36329 3844 36363
rect 3792 36320 3844 36329
rect 5172 36320 5224 36372
rect 6184 36320 6236 36372
rect 6552 36320 6604 36372
rect 7932 36320 7984 36372
rect 8392 36320 8444 36372
rect 9128 36363 9180 36372
rect 9128 36329 9153 36363
rect 9153 36329 9180 36363
rect 9128 36320 9180 36329
rect 10324 36320 10376 36372
rect 3424 36252 3476 36304
rect 1124 36184 1176 36236
rect 2872 36227 2924 36236
rect 2872 36193 2881 36227
rect 2881 36193 2915 36227
rect 2915 36193 2924 36227
rect 2872 36184 2924 36193
rect 3148 36184 3200 36236
rect 2228 36116 2280 36168
rect 3516 36184 3568 36236
rect 3884 36252 3936 36304
rect 1032 35980 1084 36032
rect 3148 35980 3200 36032
rect 4068 36184 4120 36236
rect 5540 36184 5592 36236
rect 6276 36252 6328 36304
rect 4896 35980 4948 36032
rect 5356 35980 5408 36032
rect 6092 36184 6144 36236
rect 6276 36159 6328 36168
rect 6276 36125 6285 36159
rect 6285 36125 6319 36159
rect 6319 36125 6328 36159
rect 6276 36116 6328 36125
rect 6460 36116 6512 36168
rect 7748 36184 7800 36236
rect 8116 36227 8168 36236
rect 8116 36193 8125 36227
rect 8125 36193 8159 36227
rect 8159 36193 8168 36227
rect 8116 36184 8168 36193
rect 8944 36295 8996 36304
rect 8944 36261 8953 36295
rect 8953 36261 8987 36295
rect 8987 36261 8996 36295
rect 8944 36252 8996 36261
rect 8484 36184 8536 36236
rect 8668 36227 8720 36236
rect 8668 36193 8677 36227
rect 8677 36193 8711 36227
rect 8711 36193 8720 36227
rect 8668 36184 8720 36193
rect 9128 36184 9180 36236
rect 9404 36227 9456 36236
rect 9404 36193 9413 36227
rect 9413 36193 9447 36227
rect 9447 36193 9456 36227
rect 9404 36184 9456 36193
rect 9496 36184 9548 36236
rect 9956 36184 10008 36236
rect 6920 35980 6972 36032
rect 7104 35980 7156 36032
rect 7472 35980 7524 36032
rect 8392 35980 8444 36032
rect 8668 35980 8720 36032
rect 9036 35980 9088 36032
rect 9680 35980 9732 36032
rect 3662 35878 3714 35930
rect 3726 35878 3778 35930
rect 3790 35878 3842 35930
rect 3854 35878 3906 35930
rect 3918 35878 3970 35930
rect 10062 35878 10114 35930
rect 10126 35878 10178 35930
rect 10190 35878 10242 35930
rect 10254 35878 10306 35930
rect 10318 35878 10370 35930
rect 3884 35776 3936 35828
rect 3976 35776 4028 35828
rect 5448 35776 5500 35828
rect 7288 35776 7340 35828
rect 7840 35776 7892 35828
rect 8760 35819 8812 35828
rect 8760 35785 8769 35819
rect 8769 35785 8803 35819
rect 8803 35785 8812 35819
rect 8760 35776 8812 35785
rect 9220 35776 9272 35828
rect 4068 35708 4120 35760
rect 1308 35572 1360 35624
rect 1492 35683 1544 35692
rect 1492 35649 1501 35683
rect 1501 35649 1535 35683
rect 1535 35649 1544 35683
rect 1492 35640 1544 35649
rect 4252 35640 4304 35692
rect 6644 35708 6696 35760
rect 1584 35572 1636 35624
rect 3976 35572 4028 35624
rect 4160 35572 4212 35624
rect 5172 35572 5224 35624
rect 6184 35572 6236 35624
rect 3056 35504 3108 35556
rect 1768 35436 1820 35488
rect 3148 35436 3200 35488
rect 6552 35547 6604 35556
rect 6552 35513 6561 35547
rect 6561 35513 6595 35547
rect 6595 35513 6604 35547
rect 6552 35504 6604 35513
rect 8300 35640 8352 35692
rect 9036 35640 9088 35692
rect 9220 35683 9272 35692
rect 9220 35649 9229 35683
rect 9229 35649 9263 35683
rect 9263 35649 9272 35683
rect 9220 35640 9272 35649
rect 8576 35615 8628 35624
rect 8576 35581 8585 35615
rect 8585 35581 8619 35615
rect 8619 35581 8628 35615
rect 8576 35572 8628 35581
rect 8944 35615 8996 35624
rect 8944 35581 8953 35615
rect 8953 35581 8987 35615
rect 8987 35581 8996 35615
rect 8944 35572 8996 35581
rect 9680 35572 9732 35624
rect 4804 35436 4856 35488
rect 4988 35436 5040 35488
rect 5172 35436 5224 35488
rect 5816 35479 5868 35488
rect 5816 35445 5825 35479
rect 5825 35445 5859 35479
rect 5859 35445 5868 35479
rect 5816 35436 5868 35445
rect 6000 35436 6052 35488
rect 8208 35436 8260 35488
rect 9496 35436 9548 35488
rect 9588 35479 9640 35488
rect 9588 35445 9597 35479
rect 9597 35445 9631 35479
rect 9631 35445 9640 35479
rect 9588 35436 9640 35445
rect 9772 35479 9824 35488
rect 9772 35445 9781 35479
rect 9781 35445 9815 35479
rect 9815 35445 9824 35479
rect 9772 35436 9824 35445
rect 10416 35436 10468 35488
rect 4322 35334 4374 35386
rect 4386 35334 4438 35386
rect 4450 35334 4502 35386
rect 4514 35334 4566 35386
rect 4578 35334 4630 35386
rect 10722 35334 10774 35386
rect 10786 35334 10838 35386
rect 10850 35334 10902 35386
rect 10914 35334 10966 35386
rect 10978 35334 11030 35386
rect 2780 35232 2832 35284
rect 572 35164 624 35216
rect 4252 35232 4304 35284
rect 5816 35232 5868 35284
rect 6460 35275 6512 35284
rect 6460 35241 6469 35275
rect 6469 35241 6503 35275
rect 6503 35241 6512 35275
rect 6460 35232 6512 35241
rect 6920 35232 6972 35284
rect 8024 35232 8076 35284
rect 8668 35275 8720 35284
rect 8668 35241 8677 35275
rect 8677 35241 8711 35275
rect 8711 35241 8720 35275
rect 8668 35232 8720 35241
rect 9036 35232 9088 35284
rect 3332 35164 3384 35216
rect 3424 35164 3476 35216
rect 5632 35164 5684 35216
rect 1124 35096 1176 35148
rect 1584 35139 1636 35148
rect 1584 35105 1593 35139
rect 1593 35105 1627 35139
rect 1627 35105 1636 35139
rect 1584 35096 1636 35105
rect 1768 35096 1820 35148
rect 2504 35096 2556 35148
rect 2872 35139 2924 35148
rect 2872 35105 2881 35139
rect 2881 35105 2915 35139
rect 2915 35105 2924 35139
rect 2872 35096 2924 35105
rect 3056 35139 3108 35148
rect 3056 35105 3065 35139
rect 3065 35105 3099 35139
rect 3099 35105 3108 35139
rect 3056 35096 3108 35105
rect 3148 35139 3200 35148
rect 3148 35105 3157 35139
rect 3157 35105 3191 35139
rect 3191 35105 3200 35139
rect 3148 35096 3200 35105
rect 3976 35096 4028 35148
rect 1860 35028 1912 35080
rect 2228 35071 2280 35080
rect 2228 35037 2237 35071
rect 2237 35037 2271 35071
rect 2271 35037 2280 35071
rect 2228 35028 2280 35037
rect 2320 35071 2372 35080
rect 2320 35037 2329 35071
rect 2329 35037 2363 35071
rect 2363 35037 2372 35071
rect 2320 35028 2372 35037
rect 3424 35028 3476 35080
rect 5264 35096 5316 35148
rect 5448 35096 5500 35148
rect 6368 35164 6420 35216
rect 7196 35164 7248 35216
rect 9128 35164 9180 35216
rect 9772 35164 9824 35216
rect 6000 35139 6052 35148
rect 6000 35105 6009 35139
rect 6009 35105 6043 35139
rect 6043 35105 6052 35139
rect 6000 35096 6052 35105
rect 6644 35096 6696 35148
rect 6828 35139 6880 35148
rect 6828 35105 6837 35139
rect 6837 35105 6871 35139
rect 6871 35105 6880 35139
rect 6828 35096 6880 35105
rect 7380 35139 7432 35148
rect 7380 35105 7389 35139
rect 7389 35105 7423 35139
rect 7423 35105 7432 35139
rect 7380 35096 7432 35105
rect 7472 35096 7524 35148
rect 8208 35096 8260 35148
rect 8300 35139 8352 35148
rect 8300 35105 8309 35139
rect 8309 35105 8343 35139
rect 8343 35105 8352 35139
rect 8300 35096 8352 35105
rect 4344 35028 4396 35080
rect 4988 35071 5040 35080
rect 4988 35037 4997 35071
rect 4997 35037 5031 35071
rect 5031 35037 5040 35071
rect 4988 35028 5040 35037
rect 5080 35071 5132 35080
rect 5080 35037 5089 35071
rect 5089 35037 5123 35071
rect 5123 35037 5132 35071
rect 5080 35028 5132 35037
rect 6184 35071 6236 35080
rect 6184 35037 6193 35071
rect 6193 35037 6227 35071
rect 6227 35037 6236 35071
rect 6184 35028 6236 35037
rect 6552 35028 6604 35080
rect 7748 35028 7800 35080
rect 1124 34935 1176 34944
rect 1124 34901 1133 34935
rect 1133 34901 1167 34935
rect 1167 34901 1176 34935
rect 1124 34892 1176 34901
rect 2596 34892 2648 34944
rect 5172 34960 5224 35012
rect 5356 34892 5408 34944
rect 6000 34960 6052 35012
rect 8208 34960 8260 35012
rect 8852 35096 8904 35148
rect 8944 35139 8996 35148
rect 8944 35105 8953 35139
rect 8953 35105 8987 35139
rect 8987 35105 8996 35139
rect 8944 35096 8996 35105
rect 8760 35028 8812 35080
rect 9312 34960 9364 35012
rect 8024 34892 8076 34944
rect 10416 34892 10468 34944
rect 10508 34892 10560 34944
rect 3662 34790 3714 34842
rect 3726 34790 3778 34842
rect 3790 34790 3842 34842
rect 3854 34790 3906 34842
rect 3918 34790 3970 34842
rect 10062 34790 10114 34842
rect 10126 34790 10178 34842
rect 10190 34790 10242 34842
rect 10254 34790 10306 34842
rect 10318 34790 10370 34842
rect 1308 34731 1360 34740
rect 1308 34697 1317 34731
rect 1317 34697 1351 34731
rect 1351 34697 1360 34731
rect 1308 34688 1360 34697
rect 2320 34688 2372 34740
rect 2688 34688 2740 34740
rect 3608 34688 3660 34740
rect 4344 34688 4396 34740
rect 2872 34620 2924 34672
rect 204 34484 256 34536
rect 480 34484 532 34536
rect 2596 34484 2648 34536
rect 2964 34552 3016 34604
rect 3976 34595 4028 34604
rect 3976 34561 3985 34595
rect 3985 34561 4019 34595
rect 4019 34561 4028 34595
rect 3976 34552 4028 34561
rect 4252 34552 4304 34604
rect 3056 34484 3108 34536
rect 3424 34484 3476 34536
rect 3792 34527 3844 34536
rect 3792 34493 3801 34527
rect 3801 34493 3835 34527
rect 3835 34493 3844 34527
rect 3792 34484 3844 34493
rect 4068 34527 4120 34536
rect 4068 34493 4077 34527
rect 4077 34493 4111 34527
rect 4111 34493 4120 34527
rect 4068 34484 4120 34493
rect 3148 34416 3200 34468
rect 3516 34459 3568 34468
rect 3516 34425 3525 34459
rect 3525 34425 3559 34459
rect 3559 34425 3568 34459
rect 3516 34416 3568 34425
rect 4620 34620 4672 34672
rect 4620 34484 4672 34536
rect 4988 34688 5040 34740
rect 5172 34731 5224 34740
rect 5172 34697 5181 34731
rect 5181 34697 5215 34731
rect 5215 34697 5224 34731
rect 5172 34688 5224 34697
rect 5264 34688 5316 34740
rect 8944 34688 8996 34740
rect 9312 34688 9364 34740
rect 6184 34620 6236 34672
rect 4804 34527 4856 34536
rect 4804 34493 4813 34527
rect 4813 34493 4847 34527
rect 4847 34493 4856 34527
rect 4804 34484 4856 34493
rect 5356 34484 5408 34536
rect 6276 34527 6328 34536
rect 6276 34493 6285 34527
rect 6285 34493 6319 34527
rect 6319 34493 6328 34527
rect 6276 34484 6328 34493
rect 8392 34620 8444 34672
rect 9956 34620 10008 34672
rect 11060 34620 11112 34672
rect 6644 34527 6696 34536
rect 6644 34493 6653 34527
rect 6653 34493 6687 34527
rect 6687 34493 6696 34527
rect 6644 34484 6696 34493
rect 6920 34527 6972 34536
rect 6920 34493 6929 34527
rect 6929 34493 6963 34527
rect 6963 34493 6972 34527
rect 6920 34484 6972 34493
rect 7288 34484 7340 34536
rect 7380 34484 7432 34536
rect 5264 34416 5316 34468
rect 10416 34552 10468 34604
rect 7840 34484 7892 34536
rect 8024 34527 8076 34536
rect 8024 34493 8033 34527
rect 8033 34493 8067 34527
rect 8067 34493 8076 34527
rect 8024 34484 8076 34493
rect 8116 34484 8168 34536
rect 8392 34527 8444 34536
rect 8392 34493 8401 34527
rect 8401 34493 8435 34527
rect 8435 34493 8444 34527
rect 8392 34484 8444 34493
rect 8576 34527 8628 34536
rect 8576 34493 8585 34527
rect 8585 34493 8619 34527
rect 8619 34493 8628 34527
rect 8576 34484 8628 34493
rect 8668 34527 8720 34536
rect 8668 34493 8677 34527
rect 8677 34493 8711 34527
rect 8711 34493 8720 34527
rect 8668 34484 8720 34493
rect 940 34391 992 34400
rect 940 34357 949 34391
rect 949 34357 983 34391
rect 983 34357 992 34391
rect 940 34348 992 34357
rect 2780 34348 2832 34400
rect 4896 34348 4948 34400
rect 5448 34348 5500 34400
rect 5632 34348 5684 34400
rect 6552 34348 6604 34400
rect 8392 34348 8444 34400
rect 8760 34416 8812 34468
rect 10140 34484 10192 34536
rect 10324 34527 10376 34536
rect 10324 34493 10333 34527
rect 10333 34493 10367 34527
rect 10367 34493 10376 34527
rect 10324 34484 10376 34493
rect 10600 34527 10652 34536
rect 10600 34493 10609 34527
rect 10609 34493 10643 34527
rect 10643 34493 10652 34527
rect 10600 34484 10652 34493
rect 10968 34484 11020 34536
rect 9404 34416 9456 34468
rect 10416 34416 10468 34468
rect 10232 34348 10284 34400
rect 10600 34348 10652 34400
rect 4322 34246 4374 34298
rect 4386 34246 4438 34298
rect 4450 34246 4502 34298
rect 4514 34246 4566 34298
rect 4578 34246 4630 34298
rect 10722 34246 10774 34298
rect 10786 34246 10838 34298
rect 10850 34246 10902 34298
rect 10914 34246 10966 34298
rect 10978 34246 11030 34298
rect 1032 34076 1084 34128
rect 1952 34008 2004 34060
rect 1308 33983 1360 33992
rect 1308 33949 1317 33983
rect 1317 33949 1351 33983
rect 1351 33949 1360 33983
rect 1308 33940 1360 33949
rect 2504 34076 2556 34128
rect 3424 34051 3476 34060
rect 3424 34017 3458 34051
rect 3458 34017 3476 34051
rect 3424 34008 3476 34017
rect 1584 33804 1636 33856
rect 2504 33804 2556 33856
rect 2964 33804 3016 33856
rect 3148 33983 3200 33992
rect 3148 33949 3157 33983
rect 3157 33949 3191 33983
rect 3191 33949 3200 33983
rect 3148 33940 3200 33949
rect 4528 33915 4580 33924
rect 4528 33881 4537 33915
rect 4537 33881 4571 33915
rect 4571 33881 4580 33915
rect 4528 33872 4580 33881
rect 4896 34051 4948 34060
rect 4896 34017 4905 34051
rect 4905 34017 4939 34051
rect 4939 34017 4948 34051
rect 4896 34008 4948 34017
rect 5356 34144 5408 34196
rect 6276 34144 6328 34196
rect 5172 34051 5224 34060
rect 5172 34017 5181 34051
rect 5181 34017 5215 34051
rect 5215 34017 5224 34051
rect 5172 34008 5224 34017
rect 5264 34008 5316 34060
rect 5632 34051 5684 34060
rect 5632 34017 5641 34051
rect 5641 34017 5675 34051
rect 5675 34017 5684 34051
rect 5632 34008 5684 34017
rect 5816 34008 5868 34060
rect 7104 34008 7156 34060
rect 8668 34076 8720 34128
rect 8852 34187 8904 34196
rect 8852 34153 8861 34187
rect 8861 34153 8895 34187
rect 8895 34153 8904 34187
rect 8852 34144 8904 34153
rect 8944 34144 8996 34196
rect 9404 34144 9456 34196
rect 9588 34187 9640 34196
rect 9588 34153 9597 34187
rect 9597 34153 9631 34187
rect 9631 34153 9640 34187
rect 9588 34144 9640 34153
rect 10600 34144 10652 34196
rect 7380 34008 7432 34060
rect 7840 34051 7892 34060
rect 7840 34017 7849 34051
rect 7849 34017 7883 34051
rect 7883 34017 7892 34051
rect 7840 34008 7892 34017
rect 6092 33940 6144 33992
rect 8484 34008 8536 34060
rect 8760 34008 8812 34060
rect 8944 34051 8996 34060
rect 8944 34017 8953 34051
rect 8953 34017 8987 34051
rect 8987 34017 8996 34051
rect 8944 34008 8996 34017
rect 9036 34008 9088 34060
rect 9772 34008 9824 34060
rect 10324 34008 10376 34060
rect 8208 33983 8260 33992
rect 8208 33949 8217 33983
rect 8217 33949 8251 33983
rect 8251 33949 8260 33983
rect 8208 33940 8260 33949
rect 5724 33872 5776 33924
rect 8852 33940 8904 33992
rect 6000 33804 6052 33856
rect 6828 33804 6880 33856
rect 6920 33804 6972 33856
rect 7656 33804 7708 33856
rect 8208 33847 8260 33856
rect 8208 33813 8217 33847
rect 8217 33813 8251 33847
rect 8251 33813 8260 33847
rect 8208 33804 8260 33813
rect 9312 33872 9364 33924
rect 10140 33872 10192 33924
rect 10692 33872 10744 33924
rect 8760 33804 8812 33856
rect 10232 33847 10284 33856
rect 10232 33813 10241 33847
rect 10241 33813 10275 33847
rect 10275 33813 10284 33847
rect 10232 33804 10284 33813
rect 10416 33804 10468 33856
rect 3662 33702 3714 33754
rect 3726 33702 3778 33754
rect 3790 33702 3842 33754
rect 3854 33702 3906 33754
rect 3918 33702 3970 33754
rect 10062 33702 10114 33754
rect 10126 33702 10178 33754
rect 10190 33702 10242 33754
rect 10254 33702 10306 33754
rect 10318 33702 10370 33754
rect 1952 33643 2004 33652
rect 1952 33609 1961 33643
rect 1961 33609 1995 33643
rect 1995 33609 2004 33643
rect 1952 33600 2004 33609
rect 3424 33600 3476 33652
rect 5540 33600 5592 33652
rect 2320 33532 2372 33584
rect 6920 33600 6972 33652
rect 7656 33600 7708 33652
rect 8300 33600 8352 33652
rect 8668 33600 8720 33652
rect 9312 33600 9364 33652
rect 1952 33464 2004 33516
rect 2228 33464 2280 33516
rect 5816 33507 5868 33516
rect 5816 33473 5844 33507
rect 5844 33473 5868 33507
rect 5816 33464 5868 33473
rect 1124 33439 1176 33448
rect 1124 33405 1133 33439
rect 1133 33405 1167 33439
rect 1167 33405 1176 33439
rect 1124 33396 1176 33405
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 3056 33439 3108 33448
rect 3056 33405 3065 33439
rect 3065 33405 3099 33439
rect 3099 33405 3108 33439
rect 3056 33396 3108 33405
rect 4252 33396 4304 33448
rect 5080 33439 5132 33448
rect 5080 33405 5089 33439
rect 5089 33405 5123 33439
rect 5123 33405 5132 33439
rect 5080 33396 5132 33405
rect 5540 33439 5592 33448
rect 5540 33405 5549 33439
rect 5549 33405 5583 33439
rect 5583 33405 5592 33439
rect 5540 33396 5592 33405
rect 5724 33439 5776 33448
rect 5724 33405 5733 33439
rect 5733 33405 5767 33439
rect 5767 33405 5776 33439
rect 5724 33396 5776 33405
rect 6276 33439 6328 33448
rect 6276 33405 6285 33439
rect 6285 33405 6319 33439
rect 6319 33405 6328 33439
rect 6276 33396 6328 33405
rect 6368 33439 6420 33448
rect 6368 33405 6377 33439
rect 6377 33405 6411 33439
rect 6411 33405 6420 33439
rect 6368 33396 6420 33405
rect 6552 33439 6604 33448
rect 6552 33405 6565 33439
rect 6565 33405 6604 33439
rect 6552 33396 6604 33405
rect 7104 33396 7156 33448
rect 7840 33439 7892 33448
rect 7840 33405 7849 33439
rect 7849 33405 7883 33439
rect 7883 33405 7892 33439
rect 7840 33396 7892 33405
rect 7932 33396 7984 33448
rect 6000 33371 6052 33380
rect 6000 33337 6009 33371
rect 6009 33337 6043 33371
rect 6043 33337 6052 33371
rect 6000 33328 6052 33337
rect 848 33260 900 33312
rect 2044 33260 2096 33312
rect 2504 33260 2556 33312
rect 2964 33303 3016 33312
rect 2964 33269 2973 33303
rect 2973 33269 3007 33303
rect 3007 33269 3016 33303
rect 2964 33260 3016 33269
rect 3976 33303 4028 33312
rect 3976 33269 3985 33303
rect 3985 33269 4019 33303
rect 4019 33269 4028 33303
rect 3976 33260 4028 33269
rect 4528 33260 4580 33312
rect 5172 33260 5224 33312
rect 7380 33328 7432 33380
rect 8300 33398 8352 33450
rect 8392 33439 8444 33448
rect 8392 33405 8401 33439
rect 8401 33405 8435 33439
rect 8435 33405 8444 33439
rect 8392 33396 8444 33405
rect 9220 33532 9272 33584
rect 6368 33260 6420 33312
rect 7104 33260 7156 33312
rect 7656 33260 7708 33312
rect 7840 33260 7892 33312
rect 8576 33328 8628 33380
rect 10692 33600 10744 33652
rect 9864 33532 9916 33584
rect 10416 33532 10468 33584
rect 9312 33328 9364 33380
rect 9036 33303 9088 33312
rect 9036 33269 9045 33303
rect 9045 33269 9079 33303
rect 9079 33269 9088 33303
rect 9036 33260 9088 33269
rect 9220 33260 9272 33312
rect 9772 33464 9824 33516
rect 9588 33396 9640 33448
rect 10140 33439 10192 33448
rect 10140 33405 10149 33439
rect 10149 33405 10183 33439
rect 10183 33405 10192 33439
rect 10140 33396 10192 33405
rect 10416 33439 10468 33448
rect 10416 33405 10425 33439
rect 10425 33405 10459 33439
rect 10459 33405 10468 33439
rect 10416 33396 10468 33405
rect 9772 33303 9824 33312
rect 9772 33269 9781 33303
rect 9781 33269 9815 33303
rect 9815 33269 9824 33303
rect 9772 33260 9824 33269
rect 10416 33260 10468 33312
rect 11244 33260 11296 33312
rect 4322 33158 4374 33210
rect 4386 33158 4438 33210
rect 4450 33158 4502 33210
rect 4514 33158 4566 33210
rect 4578 33158 4630 33210
rect 10722 33158 10774 33210
rect 10786 33158 10838 33210
rect 10850 33158 10902 33210
rect 10914 33158 10966 33210
rect 10978 33158 11030 33210
rect 848 33056 900 33108
rect 4344 33056 4396 33108
rect 1124 32963 1176 32972
rect 1124 32929 1133 32963
rect 1133 32929 1167 32963
rect 1167 32929 1176 32963
rect 1124 32920 1176 32929
rect 1492 32920 1544 32972
rect 1584 32963 1636 32972
rect 1584 32929 1593 32963
rect 1593 32929 1627 32963
rect 1627 32929 1636 32963
rect 1584 32920 1636 32929
rect 2044 32920 2096 32972
rect 2136 32963 2188 32972
rect 2136 32929 2145 32963
rect 2145 32929 2179 32963
rect 2179 32929 2188 32963
rect 2136 32920 2188 32929
rect 2688 32963 2740 32972
rect 2688 32929 2697 32963
rect 2697 32929 2731 32963
rect 2731 32929 2740 32963
rect 2688 32920 2740 32929
rect 1400 32852 1452 32904
rect 5816 32988 5868 33040
rect 3056 32920 3108 32972
rect 1768 32784 1820 32836
rect 2964 32784 3016 32836
rect 3516 32920 3568 32972
rect 3700 32963 3752 32972
rect 3700 32929 3709 32963
rect 3709 32929 3743 32963
rect 3743 32929 3752 32963
rect 3700 32920 3752 32929
rect 4252 32963 4304 32972
rect 4252 32929 4261 32963
rect 4261 32929 4295 32963
rect 4295 32929 4304 32963
rect 4252 32920 4304 32929
rect 4344 32963 4396 32972
rect 4344 32929 4353 32963
rect 4353 32929 4387 32963
rect 4387 32929 4396 32963
rect 4344 32920 4396 32929
rect 4896 32920 4948 32972
rect 5540 32963 5592 32972
rect 5540 32929 5549 32963
rect 5549 32929 5583 32963
rect 5583 32929 5592 32963
rect 5540 32920 5592 32929
rect 5908 32963 5960 32972
rect 5908 32929 5917 32963
rect 5917 32929 5951 32963
rect 5951 32929 5960 32963
rect 5908 32920 5960 32929
rect 6736 33056 6788 33108
rect 6828 33056 6880 33108
rect 7564 32988 7616 33040
rect 8024 32988 8076 33040
rect 5632 32852 5684 32904
rect 5724 32852 5776 32904
rect 6828 32963 6880 32972
rect 6828 32929 6837 32963
rect 6837 32929 6871 32963
rect 6871 32929 6880 32963
rect 6828 32920 6880 32929
rect 7012 32963 7064 32972
rect 7012 32929 7021 32963
rect 7021 32929 7055 32963
rect 7055 32929 7064 32963
rect 7012 32920 7064 32929
rect 7472 32963 7524 32972
rect 7472 32929 7481 32963
rect 7481 32929 7515 32963
rect 7515 32929 7524 32963
rect 7472 32920 7524 32929
rect 6368 32852 6420 32904
rect 2044 32716 2096 32768
rect 2412 32716 2464 32768
rect 2504 32759 2556 32768
rect 2504 32725 2513 32759
rect 2513 32725 2547 32759
rect 2547 32725 2556 32759
rect 2504 32716 2556 32725
rect 2688 32716 2740 32768
rect 4620 32784 4672 32836
rect 6000 32827 6052 32836
rect 6000 32793 6009 32827
rect 6009 32793 6043 32827
rect 6043 32793 6052 32827
rect 6000 32784 6052 32793
rect 4068 32759 4120 32768
rect 4068 32725 4077 32759
rect 4077 32725 4111 32759
rect 4111 32725 4120 32759
rect 4068 32716 4120 32725
rect 4988 32716 5040 32768
rect 5080 32759 5132 32768
rect 5080 32725 5089 32759
rect 5089 32725 5123 32759
rect 5123 32725 5132 32759
rect 5080 32716 5132 32725
rect 5908 32716 5960 32768
rect 6552 32784 6604 32836
rect 6736 32895 6788 32904
rect 6736 32861 6745 32895
rect 6745 32861 6779 32895
rect 6779 32861 6788 32895
rect 6736 32852 6788 32861
rect 7932 32895 7984 32904
rect 7932 32861 7941 32895
rect 7941 32861 7975 32895
rect 7975 32861 7984 32895
rect 7932 32852 7984 32861
rect 8024 32895 8076 32904
rect 8024 32861 8033 32895
rect 8033 32861 8067 32895
rect 8067 32861 8076 32895
rect 8024 32852 8076 32861
rect 8852 33099 8904 33108
rect 8852 33065 8861 33099
rect 8861 33065 8895 33099
rect 8895 33065 8904 33099
rect 8852 33056 8904 33065
rect 8300 32988 8352 33040
rect 9680 33056 9732 33108
rect 10600 33056 10652 33108
rect 10876 33056 10928 33108
rect 9036 33031 9088 33040
rect 9036 32997 9045 33031
rect 9045 32997 9079 33031
rect 9079 32997 9088 33031
rect 9036 32988 9088 32997
rect 9956 32988 10008 33040
rect 8392 32963 8444 32972
rect 8392 32929 8401 32963
rect 8401 32929 8435 32963
rect 8435 32929 8444 32963
rect 8392 32920 8444 32929
rect 8300 32852 8352 32904
rect 8668 32963 8720 32972
rect 8668 32929 8677 32963
rect 8677 32929 8711 32963
rect 8711 32929 8720 32963
rect 8668 32920 8720 32929
rect 8760 32963 8812 32972
rect 8760 32929 8769 32963
rect 8769 32929 8803 32963
rect 8803 32929 8812 32963
rect 8760 32920 8812 32929
rect 7380 32784 7432 32836
rect 9680 32920 9732 32972
rect 11336 32988 11388 33040
rect 10508 32895 10560 32904
rect 10508 32861 10517 32895
rect 10517 32861 10551 32895
rect 10551 32861 10560 32895
rect 10508 32852 10560 32861
rect 10784 32784 10836 32836
rect 6736 32716 6788 32768
rect 6920 32716 6972 32768
rect 7104 32759 7156 32768
rect 7104 32725 7113 32759
rect 7113 32725 7147 32759
rect 7147 32725 7156 32759
rect 7104 32716 7156 32725
rect 7288 32716 7340 32768
rect 7840 32716 7892 32768
rect 8576 32716 8628 32768
rect 3662 32614 3714 32666
rect 3726 32614 3778 32666
rect 3790 32614 3842 32666
rect 3854 32614 3906 32666
rect 3918 32614 3970 32666
rect 10062 32614 10114 32666
rect 10126 32614 10178 32666
rect 10190 32614 10242 32666
rect 10254 32614 10306 32666
rect 10318 32614 10370 32666
rect 1952 32512 2004 32564
rect 3516 32512 3568 32564
rect 5908 32512 5960 32564
rect 6092 32555 6144 32564
rect 6092 32521 6101 32555
rect 6101 32521 6135 32555
rect 6135 32521 6144 32555
rect 6092 32512 6144 32521
rect 6920 32512 6972 32564
rect 7104 32555 7156 32564
rect 7104 32521 7113 32555
rect 7113 32521 7147 32555
rect 7147 32521 7156 32555
rect 7104 32512 7156 32521
rect 7840 32512 7892 32564
rect 8208 32512 8260 32564
rect 10508 32512 10560 32564
rect 10876 32512 10928 32564
rect 2412 32444 2464 32496
rect 3240 32444 3292 32496
rect 3700 32444 3752 32496
rect 5540 32444 5592 32496
rect 5816 32376 5868 32428
rect 2320 32308 2372 32360
rect 1308 32240 1360 32292
rect 2688 32308 2740 32360
rect 2872 32351 2924 32360
rect 2872 32317 2881 32351
rect 2881 32317 2915 32351
rect 2915 32317 2924 32351
rect 2872 32308 2924 32317
rect 3240 32308 3292 32360
rect 3884 32308 3936 32360
rect 5264 32351 5316 32360
rect 5264 32317 5273 32351
rect 5273 32317 5307 32351
rect 5307 32317 5316 32351
rect 5264 32308 5316 32317
rect 5448 32308 5500 32360
rect 2504 32283 2556 32292
rect 2504 32249 2513 32283
rect 2513 32249 2547 32283
rect 2547 32249 2556 32283
rect 2504 32240 2556 32249
rect 20 32172 72 32224
rect 1584 32172 1636 32224
rect 2688 32172 2740 32224
rect 3516 32215 3568 32224
rect 3516 32181 3525 32215
rect 3525 32181 3559 32215
rect 3559 32181 3568 32215
rect 3516 32172 3568 32181
rect 4804 32240 4856 32292
rect 5816 32240 5868 32292
rect 6460 32444 6512 32496
rect 6184 32376 6236 32428
rect 8024 32444 8076 32496
rect 6276 32308 6328 32360
rect 7380 32419 7432 32428
rect 7380 32385 7389 32419
rect 7389 32385 7423 32419
rect 7423 32385 7432 32419
rect 7380 32376 7432 32385
rect 6552 32351 6604 32360
rect 6552 32317 6561 32351
rect 6561 32317 6595 32351
rect 6595 32317 6604 32351
rect 6552 32308 6604 32317
rect 7196 32308 7248 32360
rect 7472 32351 7524 32360
rect 7472 32317 7481 32351
rect 7481 32317 7515 32351
rect 7515 32317 7524 32351
rect 7472 32308 7524 32317
rect 6184 32240 6236 32292
rect 7012 32283 7064 32292
rect 7012 32249 7021 32283
rect 7021 32249 7055 32283
rect 7055 32249 7064 32283
rect 7012 32240 7064 32249
rect 4436 32172 4488 32224
rect 5356 32172 5408 32224
rect 5540 32172 5592 32224
rect 8300 32308 8352 32360
rect 8668 32444 8720 32496
rect 9036 32444 9088 32496
rect 9588 32444 9640 32496
rect 9496 32376 9548 32428
rect 10784 32419 10836 32428
rect 10784 32385 10793 32419
rect 10793 32385 10827 32419
rect 10827 32385 10836 32419
rect 10784 32376 10836 32385
rect 8208 32240 8260 32292
rect 8392 32240 8444 32292
rect 8668 32308 8720 32360
rect 8944 32351 8996 32360
rect 8944 32317 8953 32351
rect 8953 32317 8987 32351
rect 8987 32317 8996 32351
rect 8944 32308 8996 32317
rect 8852 32240 8904 32292
rect 9312 32308 9364 32360
rect 9588 32308 9640 32360
rect 7932 32172 7984 32224
rect 9128 32240 9180 32292
rect 9772 32240 9824 32292
rect 4322 32070 4374 32122
rect 4386 32070 4438 32122
rect 4450 32070 4502 32122
rect 4514 32070 4566 32122
rect 4578 32070 4630 32122
rect 10722 32070 10774 32122
rect 10786 32070 10838 32122
rect 10850 32070 10902 32122
rect 10914 32070 10966 32122
rect 10978 32070 11030 32122
rect 388 31968 440 32020
rect 1400 31900 1452 31952
rect 1032 31832 1084 31884
rect 1952 31832 2004 31884
rect 2228 31832 2280 31884
rect 3240 31900 3292 31952
rect 3792 32011 3844 32020
rect 3792 31977 3801 32011
rect 3801 31977 3835 32011
rect 3835 31977 3844 32011
rect 3792 31968 3844 31977
rect 4712 31968 4764 32020
rect 2688 31875 2740 31884
rect 2688 31841 2722 31875
rect 2722 31841 2740 31875
rect 2688 31832 2740 31841
rect 4436 31832 4488 31884
rect 5540 31968 5592 32020
rect 5724 31900 5776 31952
rect 5816 31943 5868 31952
rect 5816 31909 5825 31943
rect 5825 31909 5859 31943
rect 5859 31909 5868 31943
rect 5816 31900 5868 31909
rect 6092 31900 6144 31952
rect 2136 31764 2188 31816
rect 940 31628 992 31680
rect 2412 31628 2464 31680
rect 3700 31628 3752 31680
rect 5264 31696 5316 31748
rect 5816 31764 5868 31816
rect 5540 31696 5592 31748
rect 6092 31764 6144 31816
rect 6828 31968 6880 32020
rect 7564 31968 7616 32020
rect 7840 31968 7892 32020
rect 6736 31900 6788 31952
rect 8300 31968 8352 32020
rect 9312 31968 9364 32020
rect 10140 31968 10192 32020
rect 10416 31968 10468 32020
rect 6828 31875 6880 31884
rect 6828 31841 6837 31875
rect 6837 31841 6871 31875
rect 6871 31841 6880 31875
rect 6828 31832 6880 31841
rect 7380 31875 7432 31884
rect 7380 31841 7389 31875
rect 7389 31841 7423 31875
rect 7423 31841 7432 31875
rect 7380 31832 7432 31841
rect 6368 31807 6420 31816
rect 6368 31773 6377 31807
rect 6377 31773 6411 31807
rect 6411 31773 6420 31807
rect 6368 31764 6420 31773
rect 6736 31764 6788 31816
rect 7104 31764 7156 31816
rect 7564 31832 7616 31884
rect 8944 31943 8996 31952
rect 8944 31909 8953 31943
rect 8953 31909 8987 31943
rect 8987 31909 8996 31943
rect 8944 31900 8996 31909
rect 9496 31943 9548 31952
rect 9496 31909 9505 31943
rect 9505 31909 9539 31943
rect 9539 31909 9548 31943
rect 9496 31900 9548 31909
rect 9956 31900 10008 31952
rect 9036 31832 9088 31884
rect 9128 31875 9180 31884
rect 9128 31841 9137 31875
rect 9137 31841 9171 31875
rect 9171 31841 9180 31875
rect 9128 31832 9180 31841
rect 5172 31628 5224 31680
rect 6184 31696 6236 31748
rect 7196 31696 7248 31748
rect 8852 31764 8904 31816
rect 9128 31696 9180 31748
rect 10508 31875 10560 31884
rect 10508 31841 10517 31875
rect 10517 31841 10551 31875
rect 10551 31841 10560 31875
rect 10508 31832 10560 31841
rect 9496 31764 9548 31816
rect 6736 31671 6788 31680
rect 6736 31637 6745 31671
rect 6745 31637 6779 31671
rect 6779 31637 6788 31671
rect 6736 31628 6788 31637
rect 6920 31628 6972 31680
rect 7564 31628 7616 31680
rect 8208 31628 8260 31680
rect 8668 31628 8720 31680
rect 9956 31807 10008 31816
rect 9956 31773 9965 31807
rect 9965 31773 9999 31807
rect 9999 31773 10008 31807
rect 9956 31764 10008 31773
rect 10048 31807 10100 31816
rect 10048 31773 10057 31807
rect 10057 31773 10091 31807
rect 10091 31773 10100 31807
rect 10048 31764 10100 31773
rect 10140 31807 10192 31816
rect 10140 31773 10149 31807
rect 10149 31773 10183 31807
rect 10183 31773 10192 31807
rect 10140 31764 10192 31773
rect 9680 31671 9732 31680
rect 9680 31637 9689 31671
rect 9689 31637 9723 31671
rect 9723 31637 9732 31671
rect 9680 31628 9732 31637
rect 3662 31526 3714 31578
rect 3726 31526 3778 31578
rect 3790 31526 3842 31578
rect 3854 31526 3906 31578
rect 3918 31526 3970 31578
rect 10062 31526 10114 31578
rect 10126 31526 10178 31578
rect 10190 31526 10242 31578
rect 10254 31526 10306 31578
rect 10318 31526 10370 31578
rect 848 31424 900 31476
rect 2872 31424 2924 31476
rect 3148 31424 3200 31476
rect 5632 31467 5684 31476
rect 5632 31433 5641 31467
rect 5641 31433 5675 31467
rect 5675 31433 5684 31467
rect 5632 31424 5684 31433
rect 5908 31424 5960 31476
rect 6552 31467 6604 31476
rect 6552 31433 6561 31467
rect 6561 31433 6595 31467
rect 6595 31433 6604 31467
rect 6552 31424 6604 31433
rect 2780 31356 2832 31408
rect 1308 31220 1360 31272
rect 1584 31263 1636 31272
rect 1584 31229 1593 31263
rect 1593 31229 1627 31263
rect 1627 31229 1636 31263
rect 1584 31220 1636 31229
rect 1952 31288 2004 31340
rect 4252 31356 4304 31408
rect 4896 31356 4948 31408
rect 6368 31356 6420 31408
rect 6736 31356 6788 31408
rect 7380 31424 7432 31476
rect 7564 31424 7616 31476
rect 8392 31424 8444 31476
rect 9404 31424 9456 31476
rect 7840 31356 7892 31408
rect 8576 31356 8628 31408
rect 2228 31220 2280 31272
rect 3056 31288 3108 31340
rect 5264 31331 5316 31340
rect 5264 31297 5273 31331
rect 5273 31297 5307 31331
rect 5307 31297 5316 31331
rect 5264 31288 5316 31297
rect 5540 31288 5592 31340
rect 6460 31288 6512 31340
rect 2320 31195 2372 31204
rect 2320 31161 2329 31195
rect 2329 31161 2363 31195
rect 2363 31161 2372 31195
rect 2320 31152 2372 31161
rect 1400 31127 1452 31136
rect 1400 31093 1409 31127
rect 1409 31093 1443 31127
rect 1443 31093 1452 31127
rect 1400 31084 1452 31093
rect 1768 31127 1820 31136
rect 1768 31093 1777 31127
rect 1777 31093 1811 31127
rect 1811 31093 1820 31127
rect 1768 31084 1820 31093
rect 2044 31084 2096 31136
rect 2872 31152 2924 31204
rect 2596 31084 2648 31136
rect 3240 31263 3292 31272
rect 3240 31229 3249 31263
rect 3249 31229 3283 31263
rect 3283 31229 3292 31263
rect 3240 31220 3292 31229
rect 4068 31220 4120 31272
rect 4988 31263 5040 31272
rect 4988 31229 4997 31263
rect 4997 31229 5031 31263
rect 5031 31229 5040 31263
rect 4988 31220 5040 31229
rect 6092 31220 6144 31272
rect 6184 31263 6236 31272
rect 6184 31229 6193 31263
rect 6193 31229 6227 31263
rect 6227 31229 6236 31263
rect 6184 31220 6236 31229
rect 6276 31220 6328 31272
rect 6644 31263 6696 31272
rect 6644 31229 6653 31263
rect 6653 31229 6687 31263
rect 6687 31229 6696 31263
rect 6644 31220 6696 31229
rect 7656 31288 7708 31340
rect 5356 31152 5408 31204
rect 5540 31152 5592 31204
rect 3240 31084 3292 31136
rect 4252 31084 4304 31136
rect 4620 31084 4672 31136
rect 5632 31084 5684 31136
rect 5908 31195 5960 31204
rect 5908 31161 5917 31195
rect 5917 31161 5951 31195
rect 5951 31161 5960 31195
rect 5908 31152 5960 31161
rect 6460 31152 6512 31204
rect 7380 31127 7432 31136
rect 7380 31093 7389 31127
rect 7389 31093 7423 31127
rect 7423 31093 7432 31127
rect 7380 31084 7432 31093
rect 8116 31220 8168 31272
rect 8392 31152 8444 31204
rect 8576 31195 8628 31204
rect 8576 31161 8585 31195
rect 8585 31161 8619 31195
rect 8619 31161 8628 31195
rect 8576 31152 8628 31161
rect 9864 31263 9916 31272
rect 9864 31229 9882 31263
rect 9882 31229 9916 31263
rect 9864 31220 9916 31229
rect 10508 31220 10560 31272
rect 10600 31152 10652 31204
rect 8208 31127 8260 31136
rect 8208 31093 8217 31127
rect 8217 31093 8251 31127
rect 8251 31093 8260 31127
rect 8208 31084 8260 31093
rect 8300 31084 8352 31136
rect 8852 31084 8904 31136
rect 9956 31084 10008 31136
rect 4322 30982 4374 31034
rect 4386 30982 4438 31034
rect 4450 30982 4502 31034
rect 4514 30982 4566 31034
rect 4578 30982 4630 31034
rect 10722 30982 10774 31034
rect 10786 30982 10838 31034
rect 10850 30982 10902 31034
rect 10914 30982 10966 31034
rect 10978 30982 11030 31034
rect 1032 30923 1084 30932
rect 1032 30889 1041 30923
rect 1041 30889 1075 30923
rect 1075 30889 1084 30923
rect 1032 30880 1084 30889
rect 1308 30812 1360 30864
rect 1952 30880 2004 30932
rect 2964 30880 3016 30932
rect 3332 30923 3384 30932
rect 3332 30889 3359 30923
rect 3359 30889 3384 30923
rect 3332 30880 3384 30889
rect 4160 30880 4212 30932
rect 4436 30880 4488 30932
rect 5724 30880 5776 30932
rect 6460 30880 6512 30932
rect 6644 30880 6696 30932
rect 6736 30880 6788 30932
rect 7380 30880 7432 30932
rect 8944 30880 8996 30932
rect 1492 30744 1544 30796
rect 1952 30787 2004 30796
rect 1952 30753 1961 30787
rect 1961 30753 1995 30787
rect 1995 30753 2004 30787
rect 1952 30744 2004 30753
rect 2044 30787 2096 30796
rect 2044 30753 2053 30787
rect 2053 30753 2087 30787
rect 2087 30753 2096 30787
rect 2044 30744 2096 30753
rect 1032 30676 1084 30728
rect 2596 30744 2648 30796
rect 2688 30744 2740 30796
rect 3424 30812 3476 30864
rect 3516 30855 3568 30864
rect 3516 30821 3525 30855
rect 3525 30821 3559 30855
rect 3559 30821 3568 30855
rect 3516 30812 3568 30821
rect 4252 30812 4304 30864
rect 5356 30787 5408 30796
rect 5356 30753 5365 30787
rect 5365 30753 5399 30787
rect 5399 30753 5408 30787
rect 5356 30744 5408 30753
rect 5540 30744 5592 30796
rect 5816 30787 5868 30796
rect 5816 30753 5825 30787
rect 5825 30753 5859 30787
rect 5859 30753 5868 30787
rect 5816 30744 5868 30753
rect 2228 30676 2280 30728
rect 3516 30676 3568 30728
rect 1584 30608 1636 30660
rect 2780 30608 2832 30660
rect 1400 30540 1452 30592
rect 1676 30540 1728 30592
rect 1768 30540 1820 30592
rect 2964 30583 3016 30592
rect 2964 30549 2973 30583
rect 2973 30549 3007 30583
rect 3007 30549 3016 30583
rect 2964 30540 3016 30549
rect 4896 30676 4948 30728
rect 4988 30676 5040 30728
rect 6276 30676 6328 30728
rect 7288 30812 7340 30864
rect 3976 30608 4028 30660
rect 4344 30608 4396 30660
rect 5632 30608 5684 30660
rect 7564 30787 7616 30796
rect 7564 30753 7573 30787
rect 7573 30753 7607 30787
rect 7607 30753 7616 30787
rect 7564 30744 7616 30753
rect 7748 30812 7800 30864
rect 8116 30744 8168 30796
rect 8300 30787 8352 30796
rect 8300 30753 8309 30787
rect 8309 30753 8343 30787
rect 8343 30753 8352 30787
rect 8300 30744 8352 30753
rect 9680 30812 9732 30864
rect 7104 30719 7156 30728
rect 7104 30685 7113 30719
rect 7113 30685 7147 30719
rect 7147 30685 7156 30719
rect 7104 30676 7156 30685
rect 9772 30676 9824 30728
rect 7564 30608 7616 30660
rect 4252 30540 4304 30592
rect 4804 30540 4856 30592
rect 6184 30583 6236 30592
rect 6184 30549 6193 30583
rect 6193 30549 6227 30583
rect 6227 30549 6236 30583
rect 6184 30540 6236 30549
rect 6552 30540 6604 30592
rect 7472 30540 7524 30592
rect 8392 30540 8444 30592
rect 8944 30540 8996 30592
rect 9404 30540 9456 30592
rect 10508 30540 10560 30592
rect 3662 30438 3714 30490
rect 3726 30438 3778 30490
rect 3790 30438 3842 30490
rect 3854 30438 3906 30490
rect 3918 30438 3970 30490
rect 10062 30438 10114 30490
rect 10126 30438 10178 30490
rect 10190 30438 10242 30490
rect 10254 30438 10306 30490
rect 10318 30438 10370 30490
rect 20 30336 72 30388
rect 388 30336 440 30388
rect 1492 30379 1544 30388
rect 1492 30345 1501 30379
rect 1501 30345 1535 30379
rect 1535 30345 1544 30379
rect 1492 30336 1544 30345
rect 2872 30336 2924 30388
rect 3240 30336 3292 30388
rect 1308 30268 1360 30320
rect 848 30200 900 30252
rect 4344 30336 4396 30388
rect 5080 30336 5132 30388
rect 5264 30336 5316 30388
rect 5816 30336 5868 30388
rect 6092 30336 6144 30388
rect 4252 30268 4304 30320
rect 2044 30132 2096 30184
rect 2228 30175 2280 30184
rect 2228 30141 2237 30175
rect 2237 30141 2271 30175
rect 2271 30141 2280 30175
rect 2228 30132 2280 30141
rect 1584 30064 1636 30116
rect 2228 29996 2280 30048
rect 2964 30132 3016 30184
rect 3148 30064 3200 30116
rect 3332 30132 3384 30184
rect 3424 30175 3476 30184
rect 3424 30141 3433 30175
rect 3433 30141 3467 30175
rect 3467 30141 3476 30175
rect 3424 30132 3476 30141
rect 3884 30132 3936 30184
rect 4436 30132 4488 30184
rect 5540 30268 5592 30320
rect 6460 30336 6512 30388
rect 7196 30336 7248 30388
rect 8300 30336 8352 30388
rect 9588 30336 9640 30388
rect 6552 30268 6604 30320
rect 6920 30268 6972 30320
rect 4804 30200 4856 30252
rect 5080 30200 5132 30252
rect 5356 30200 5408 30252
rect 4896 30175 4948 30184
rect 4896 30141 4905 30175
rect 4905 30141 4939 30175
rect 4939 30141 4948 30175
rect 4896 30132 4948 30141
rect 5724 30132 5776 30184
rect 5908 30132 5960 30184
rect 6092 30175 6144 30184
rect 6092 30141 6101 30175
rect 6101 30141 6135 30175
rect 6135 30141 6144 30175
rect 6092 30132 6144 30141
rect 6184 30132 6236 30184
rect 6552 30132 6604 30184
rect 4712 30064 4764 30116
rect 4804 30064 4856 30116
rect 5172 30064 5224 30116
rect 4252 29996 4304 30048
rect 5540 29996 5592 30048
rect 6920 30175 6972 30184
rect 6920 30141 6929 30175
rect 6929 30141 6963 30175
rect 6963 30141 6972 30175
rect 6920 30132 6972 30141
rect 7196 30200 7248 30252
rect 8208 30268 8260 30320
rect 8668 30200 8720 30252
rect 8852 30200 8904 30252
rect 7932 30175 7984 30184
rect 7932 30141 7941 30175
rect 7941 30141 7975 30175
rect 7975 30141 7984 30175
rect 7932 30132 7984 30141
rect 8208 30175 8260 30184
rect 8208 30141 8217 30175
rect 8217 30141 8251 30175
rect 8251 30141 8260 30175
rect 8208 30132 8260 30141
rect 9128 30132 9180 30184
rect 7472 29996 7524 30048
rect 7748 29996 7800 30048
rect 8300 30064 8352 30116
rect 8484 30064 8536 30116
rect 9220 30064 9272 30116
rect 10232 30039 10284 30048
rect 10232 30005 10241 30039
rect 10241 30005 10275 30039
rect 10275 30005 10284 30039
rect 10232 29996 10284 30005
rect 11336 29996 11388 30048
rect 4322 29894 4374 29946
rect 4386 29894 4438 29946
rect 4450 29894 4502 29946
rect 4514 29894 4566 29946
rect 4578 29894 4630 29946
rect 10722 29894 10774 29946
rect 10786 29894 10838 29946
rect 10850 29894 10902 29946
rect 10914 29894 10966 29946
rect 10978 29894 11030 29946
rect 2228 29792 2280 29844
rect 2596 29792 2648 29844
rect 2872 29792 2924 29844
rect 3424 29767 3476 29776
rect 3424 29733 3433 29767
rect 3433 29733 3467 29767
rect 3467 29733 3476 29767
rect 3424 29724 3476 29733
rect 4068 29724 4120 29776
rect 4804 29792 4856 29844
rect 4344 29724 4396 29776
rect 5448 29792 5500 29844
rect 5632 29792 5684 29844
rect 1676 29699 1728 29708
rect 1676 29665 1685 29699
rect 1685 29665 1719 29699
rect 1719 29665 1728 29699
rect 1676 29656 1728 29665
rect 1768 29699 1820 29708
rect 1768 29665 1777 29699
rect 1777 29665 1811 29699
rect 1811 29665 1820 29699
rect 1768 29656 1820 29665
rect 1860 29699 1912 29708
rect 1860 29665 1869 29699
rect 1869 29665 1903 29699
rect 1903 29665 1912 29699
rect 1860 29656 1912 29665
rect 1216 29631 1268 29640
rect 1216 29597 1225 29631
rect 1225 29597 1259 29631
rect 1259 29597 1268 29631
rect 1216 29588 1268 29597
rect 2228 29656 2280 29708
rect 1676 29520 1728 29572
rect 20 29452 72 29504
rect 2136 29631 2188 29640
rect 2136 29597 2145 29631
rect 2145 29597 2179 29631
rect 2179 29597 2188 29631
rect 2136 29588 2188 29597
rect 2320 29588 2372 29640
rect 2872 29699 2924 29708
rect 2872 29665 2881 29699
rect 2881 29665 2915 29699
rect 2915 29665 2924 29699
rect 2872 29656 2924 29665
rect 3332 29656 3384 29708
rect 4896 29656 4948 29708
rect 5356 29656 5408 29708
rect 5632 29699 5684 29708
rect 5632 29665 5641 29699
rect 5641 29665 5675 29699
rect 5675 29665 5684 29699
rect 5632 29656 5684 29665
rect 3148 29588 3200 29640
rect 4712 29631 4764 29640
rect 4712 29597 4721 29631
rect 4721 29597 4755 29631
rect 4755 29597 4764 29631
rect 4712 29588 4764 29597
rect 6092 29792 6144 29844
rect 7104 29792 7156 29844
rect 8208 29792 8260 29844
rect 8576 29792 8628 29844
rect 9312 29792 9364 29844
rect 11244 29792 11296 29844
rect 6368 29656 6420 29708
rect 6460 29699 6512 29708
rect 6460 29665 6469 29699
rect 6469 29665 6503 29699
rect 6503 29665 6512 29699
rect 6460 29656 6512 29665
rect 6552 29656 6604 29708
rect 6736 29656 6788 29708
rect 7472 29699 7524 29708
rect 7472 29665 7481 29699
rect 7481 29665 7515 29699
rect 7515 29665 7524 29699
rect 7472 29656 7524 29665
rect 7656 29656 7708 29708
rect 7840 29699 7892 29708
rect 7840 29665 7849 29699
rect 7849 29665 7883 29699
rect 7883 29665 7892 29699
rect 7840 29656 7892 29665
rect 6644 29520 6696 29572
rect 7472 29520 7524 29572
rect 7748 29631 7800 29640
rect 7748 29597 7757 29631
rect 7757 29597 7791 29631
rect 7791 29597 7800 29631
rect 7748 29588 7800 29597
rect 8668 29656 8720 29708
rect 9404 29724 9456 29776
rect 9956 29724 10008 29776
rect 10232 29724 10284 29776
rect 8944 29588 8996 29640
rect 8576 29520 8628 29572
rect 10692 29588 10744 29640
rect 2320 29452 2372 29504
rect 2688 29452 2740 29504
rect 2964 29452 3016 29504
rect 4988 29452 5040 29504
rect 5080 29452 5132 29504
rect 5724 29452 5776 29504
rect 6092 29452 6144 29504
rect 6368 29452 6420 29504
rect 6828 29452 6880 29504
rect 7104 29452 7156 29504
rect 7196 29495 7248 29504
rect 7196 29461 7205 29495
rect 7205 29461 7239 29495
rect 7239 29461 7248 29495
rect 7196 29452 7248 29461
rect 9404 29452 9456 29504
rect 9588 29452 9640 29504
rect 9680 29452 9732 29504
rect 10508 29520 10560 29572
rect 10416 29452 10468 29504
rect 3662 29350 3714 29402
rect 3726 29350 3778 29402
rect 3790 29350 3842 29402
rect 3854 29350 3906 29402
rect 3918 29350 3970 29402
rect 10062 29350 10114 29402
rect 10126 29350 10178 29402
rect 10190 29350 10242 29402
rect 10254 29350 10306 29402
rect 10318 29350 10370 29402
rect 388 29112 440 29164
rect 1124 29248 1176 29300
rect 1952 29248 2004 29300
rect 6460 29248 6512 29300
rect 6828 29248 6880 29300
rect 6920 29291 6972 29300
rect 6920 29257 6929 29291
rect 6929 29257 6963 29291
rect 6963 29257 6972 29291
rect 6920 29248 6972 29257
rect 7104 29248 7156 29300
rect 1400 29180 1452 29232
rect 1492 29180 1544 29232
rect 2136 29180 2188 29232
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 848 29019 900 29028
rect 848 28985 857 29019
rect 857 28985 891 29019
rect 891 28985 900 29019
rect 848 28976 900 28985
rect 1032 29087 1084 29096
rect 1032 29053 1041 29087
rect 1041 29053 1075 29087
rect 1075 29053 1084 29087
rect 1032 29044 1084 29053
rect 1124 29087 1176 29096
rect 1124 29053 1133 29087
rect 1133 29053 1167 29087
rect 1167 29053 1176 29087
rect 1124 29044 1176 29053
rect 3056 29180 3108 29232
rect 4620 29180 4672 29232
rect 5080 29223 5132 29232
rect 5080 29189 5089 29223
rect 5089 29189 5123 29223
rect 5123 29189 5132 29223
rect 5080 29180 5132 29189
rect 1216 29019 1268 29028
rect 1216 28985 1225 29019
rect 1225 28985 1259 29019
rect 1259 28985 1268 29019
rect 1216 28976 1268 28985
rect 2872 29047 2873 29074
rect 2873 29047 2907 29074
rect 2907 29047 2924 29074
rect 2872 29022 2924 29047
rect 1032 28908 1084 28960
rect 1308 28908 1360 28960
rect 2228 28908 2280 28960
rect 2872 28951 2924 28960
rect 2872 28917 2881 28951
rect 2881 28917 2915 28951
rect 2915 28917 2924 28951
rect 2872 28908 2924 28917
rect 3148 29112 3200 29164
rect 5632 29112 5684 29164
rect 4068 29044 4120 29096
rect 5540 29044 5592 29096
rect 5816 29087 5868 29096
rect 5816 29053 5825 29087
rect 5825 29053 5859 29087
rect 5859 29053 5868 29087
rect 5816 29044 5868 29053
rect 3240 28976 3292 29028
rect 3332 28976 3384 29028
rect 3884 28908 3936 28960
rect 4344 28908 4396 28960
rect 4804 28908 4856 28960
rect 4896 28951 4948 28960
rect 4896 28917 4905 28951
rect 4905 28917 4939 28951
rect 4939 28917 4948 28951
rect 4896 28908 4948 28917
rect 5448 28976 5500 29028
rect 5080 28908 5132 28960
rect 5816 28908 5868 28960
rect 7288 29180 7340 29232
rect 6184 29044 6236 29096
rect 6736 29044 6788 29096
rect 7104 29087 7156 29096
rect 7104 29053 7113 29087
rect 7113 29053 7147 29087
rect 7147 29053 7156 29087
rect 7104 29044 7156 29053
rect 7196 29044 7248 29096
rect 8208 29291 8260 29300
rect 8208 29257 8217 29291
rect 8217 29257 8251 29291
rect 8251 29257 8260 29291
rect 8208 29248 8260 29257
rect 8392 29180 8444 29232
rect 8576 29180 8628 29232
rect 9128 29291 9180 29300
rect 9128 29257 9137 29291
rect 9137 29257 9171 29291
rect 9171 29257 9180 29291
rect 9128 29248 9180 29257
rect 8024 29112 8076 29164
rect 9588 29248 9640 29300
rect 6184 28908 6236 28960
rect 6460 28976 6512 29028
rect 7748 29019 7800 29028
rect 7748 28985 7757 29019
rect 7757 28985 7791 29019
rect 7791 28985 7800 29019
rect 7748 28976 7800 28985
rect 8024 28976 8076 29028
rect 8576 29044 8628 29096
rect 8760 29044 8812 29096
rect 8392 28976 8444 29028
rect 9220 28976 9272 29028
rect 9128 28951 9180 28960
rect 9128 28917 9137 28951
rect 9137 28917 9171 28951
rect 9171 28917 9180 28951
rect 9128 28908 9180 28917
rect 10140 28908 10192 28960
rect 10692 28908 10744 28960
rect 388 28772 440 28824
rect 4322 28806 4374 28858
rect 4386 28806 4438 28858
rect 4450 28806 4502 28858
rect 4514 28806 4566 28858
rect 4578 28806 4630 28858
rect 10722 28806 10774 28858
rect 10786 28806 10838 28858
rect 10850 28806 10902 28858
rect 10914 28806 10966 28858
rect 10978 28806 11030 28858
rect 1952 28704 2004 28756
rect 2228 28704 2280 28756
rect 2964 28704 3016 28756
rect 112 28636 164 28688
rect 1308 28636 1360 28688
rect 3332 28704 3384 28756
rect 4068 28747 4120 28756
rect 4068 28713 4077 28747
rect 4077 28713 4111 28747
rect 4111 28713 4120 28747
rect 4068 28704 4120 28713
rect 6276 28704 6328 28756
rect 6920 28704 6972 28756
rect 9128 28704 9180 28756
rect 848 28611 900 28620
rect 848 28577 857 28611
rect 857 28577 891 28611
rect 891 28577 900 28611
rect 848 28568 900 28577
rect 1952 28568 2004 28620
rect 112 28500 164 28552
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 940 28432 992 28484
rect 1584 28432 1636 28484
rect 1308 28364 1360 28416
rect 2136 28568 2188 28620
rect 2136 28432 2188 28484
rect 2872 28611 2924 28620
rect 2872 28577 2881 28611
rect 2881 28577 2915 28611
rect 2915 28577 2924 28611
rect 2872 28568 2924 28577
rect 3332 28568 3384 28620
rect 2228 28364 2280 28416
rect 2412 28407 2464 28416
rect 2412 28373 2421 28407
rect 2421 28373 2455 28407
rect 2455 28373 2464 28407
rect 2412 28364 2464 28373
rect 3240 28500 3292 28552
rect 3608 28611 3660 28620
rect 3608 28577 3617 28611
rect 3617 28577 3651 28611
rect 3651 28577 3660 28611
rect 3608 28568 3660 28577
rect 4896 28636 4948 28688
rect 4252 28568 4304 28620
rect 4620 28611 4672 28620
rect 4620 28577 4629 28611
rect 4629 28577 4663 28611
rect 4663 28577 4672 28611
rect 4620 28568 4672 28577
rect 2780 28432 2832 28484
rect 4252 28475 4304 28484
rect 4252 28441 4261 28475
rect 4261 28441 4295 28475
rect 4295 28441 4304 28475
rect 4252 28432 4304 28441
rect 4436 28500 4488 28552
rect 4988 28500 5040 28552
rect 5448 28611 5500 28620
rect 5448 28577 5457 28611
rect 5457 28577 5491 28611
rect 5491 28577 5500 28611
rect 5448 28568 5500 28577
rect 5816 28636 5868 28688
rect 6368 28611 6420 28620
rect 6368 28577 6377 28611
rect 6377 28577 6411 28611
rect 6411 28577 6420 28611
rect 6368 28568 6420 28577
rect 6460 28611 6512 28620
rect 6460 28577 6469 28611
rect 6469 28577 6503 28611
rect 6503 28577 6512 28611
rect 6460 28568 6512 28577
rect 6552 28568 6604 28620
rect 7012 28568 7064 28620
rect 7196 28679 7248 28688
rect 7196 28645 7205 28679
rect 7205 28645 7239 28679
rect 7239 28645 7248 28679
rect 7196 28636 7248 28645
rect 9404 28679 9456 28688
rect 9404 28645 9413 28679
rect 9413 28645 9447 28679
rect 9447 28645 9456 28679
rect 9404 28636 9456 28645
rect 9496 28636 9548 28688
rect 7656 28568 7708 28620
rect 2964 28364 3016 28416
rect 3608 28364 3660 28416
rect 3884 28364 3936 28416
rect 4344 28364 4396 28416
rect 4528 28364 4580 28416
rect 5448 28364 5500 28416
rect 7380 28407 7432 28416
rect 7380 28373 7389 28407
rect 7389 28373 7423 28407
rect 7423 28373 7432 28407
rect 7380 28364 7432 28373
rect 7656 28364 7708 28416
rect 8208 28611 8260 28620
rect 8208 28577 8217 28611
rect 8217 28577 8251 28611
rect 8251 28577 8260 28611
rect 8208 28568 8260 28577
rect 8392 28611 8444 28620
rect 8392 28577 8401 28611
rect 8401 28577 8435 28611
rect 8435 28577 8444 28611
rect 8392 28568 8444 28577
rect 8576 28568 8628 28620
rect 8944 28611 8996 28620
rect 8944 28577 8953 28611
rect 8953 28577 8987 28611
rect 8987 28577 8996 28611
rect 8944 28568 8996 28577
rect 9128 28568 9180 28620
rect 9956 28568 10008 28620
rect 10416 28568 10468 28620
rect 9312 28500 9364 28552
rect 9404 28500 9456 28552
rect 11336 28500 11388 28552
rect 8300 28432 8352 28484
rect 8760 28432 8812 28484
rect 9312 28364 9364 28416
rect 9496 28407 9548 28416
rect 9496 28373 9505 28407
rect 9505 28373 9539 28407
rect 9539 28373 9548 28407
rect 9496 28364 9548 28373
rect 10508 28432 10560 28484
rect 3662 28262 3714 28314
rect 3726 28262 3778 28314
rect 3790 28262 3842 28314
rect 3854 28262 3906 28314
rect 3918 28262 3970 28314
rect 10062 28262 10114 28314
rect 10126 28262 10178 28314
rect 10190 28262 10242 28314
rect 10254 28262 10306 28314
rect 10318 28262 10370 28314
rect 1860 28160 1912 28212
rect 848 28135 900 28144
rect 848 28101 857 28135
rect 857 28101 891 28135
rect 891 28101 900 28135
rect 3056 28160 3108 28212
rect 3148 28160 3200 28212
rect 3608 28203 3660 28212
rect 3608 28169 3617 28203
rect 3617 28169 3651 28203
rect 3651 28169 3660 28203
rect 3608 28160 3660 28169
rect 3884 28160 3936 28212
rect 4436 28160 4488 28212
rect 9496 28160 9548 28212
rect 10140 28160 10192 28212
rect 848 28092 900 28101
rect 112 27956 164 28008
rect 1492 28024 1544 28076
rect 2228 28024 2280 28076
rect 1124 27999 1176 28008
rect 1124 27965 1133 27999
rect 1133 27965 1167 27999
rect 1167 27965 1176 27999
rect 1124 27956 1176 27965
rect 1400 27999 1452 28008
rect 1400 27965 1409 27999
rect 1409 27965 1443 27999
rect 1443 27965 1452 27999
rect 1400 27956 1452 27965
rect 1860 27956 1912 28008
rect 848 27820 900 27872
rect 1584 27888 1636 27940
rect 2136 27820 2188 27872
rect 2596 28024 2648 28076
rect 3148 28024 3200 28076
rect 4068 28092 4120 28144
rect 6184 28092 6236 28144
rect 8208 28092 8260 28144
rect 3700 28067 3752 28076
rect 3700 28033 3709 28067
rect 3709 28033 3743 28067
rect 3743 28033 3752 28067
rect 3700 28024 3752 28033
rect 3792 28067 3844 28076
rect 3792 28033 3801 28067
rect 3801 28033 3835 28067
rect 3835 28033 3844 28067
rect 3792 28024 3844 28033
rect 4804 28024 4856 28076
rect 7012 28024 7064 28076
rect 2688 27888 2740 27940
rect 2780 27820 2832 27872
rect 3516 27956 3568 28008
rect 4344 27956 4396 28008
rect 4712 27956 4764 28008
rect 4896 27999 4948 28008
rect 4896 27965 4905 27999
rect 4905 27965 4939 27999
rect 4939 27965 4948 27999
rect 4896 27956 4948 27965
rect 4804 27888 4856 27940
rect 4528 27820 4580 27872
rect 5080 27820 5132 27872
rect 5632 27888 5684 27940
rect 6184 27956 6236 28008
rect 6000 27888 6052 27940
rect 5908 27820 5960 27872
rect 6552 27999 6604 28008
rect 6552 27965 6561 27999
rect 6561 27965 6595 27999
rect 6595 27965 6604 27999
rect 6552 27956 6604 27965
rect 6736 27956 6788 28008
rect 8208 27999 8260 28008
rect 8208 27965 8217 27999
rect 8217 27965 8251 27999
rect 8251 27965 8260 27999
rect 8208 27956 8260 27965
rect 11060 28092 11112 28144
rect 8944 28024 8996 28076
rect 9404 28067 9456 28076
rect 9404 28033 9413 28067
rect 9413 28033 9447 28067
rect 9447 28033 9456 28067
rect 9404 28024 9456 28033
rect 9496 28067 9548 28076
rect 9496 28033 9505 28067
rect 9505 28033 9539 28067
rect 9539 28033 9548 28067
rect 9496 28024 9548 28033
rect 9772 28024 9824 28076
rect 9956 28024 10008 28076
rect 10600 28067 10652 28076
rect 10600 28033 10609 28067
rect 10609 28033 10643 28067
rect 10643 28033 10652 28067
rect 10600 28024 10652 28033
rect 9128 27956 9180 28008
rect 10416 27956 10468 28008
rect 6920 27888 6972 27940
rect 7104 27888 7156 27940
rect 7472 27820 7524 27872
rect 8116 27888 8168 27940
rect 9312 27888 9364 27940
rect 9496 27888 9548 27940
rect 9772 27888 9824 27940
rect 10048 27888 10100 27940
rect 8300 27820 8352 27872
rect 9220 27820 9272 27872
rect 4322 27718 4374 27770
rect 4386 27718 4438 27770
rect 4450 27718 4502 27770
rect 4514 27718 4566 27770
rect 4578 27718 4630 27770
rect 10722 27718 10774 27770
rect 10786 27718 10838 27770
rect 10850 27718 10902 27770
rect 10914 27718 10966 27770
rect 10978 27718 11030 27770
rect 1400 27616 1452 27668
rect 1768 27548 1820 27600
rect 1952 27616 2004 27668
rect 4068 27616 4120 27668
rect 2780 27548 2832 27600
rect 3792 27548 3844 27600
rect 4252 27548 4304 27600
rect 4620 27548 4672 27600
rect 4988 27548 5040 27600
rect 5448 27548 5500 27600
rect 5724 27616 5776 27668
rect 20 27480 72 27532
rect 1584 27412 1636 27464
rect 940 27344 992 27396
rect 1860 27523 1912 27532
rect 1860 27489 1869 27523
rect 1869 27489 1903 27523
rect 1903 27489 1912 27523
rect 1860 27480 1912 27489
rect 2044 27480 2096 27532
rect 2412 27480 2464 27532
rect 2688 27523 2740 27532
rect 2688 27489 2697 27523
rect 2697 27489 2731 27523
rect 2731 27489 2740 27523
rect 2688 27480 2740 27489
rect 1768 27412 1820 27464
rect 3976 27480 4028 27532
rect 4712 27480 4764 27532
rect 3240 27412 3292 27464
rect 3056 27344 3108 27396
rect 3516 27455 3568 27464
rect 3516 27421 3525 27455
rect 3525 27421 3559 27455
rect 3559 27421 3568 27455
rect 3516 27412 3568 27421
rect 5080 27480 5132 27532
rect 5356 27480 5408 27532
rect 5724 27480 5776 27532
rect 6000 27548 6052 27600
rect 6736 27591 6788 27600
rect 6736 27557 6745 27591
rect 6745 27557 6779 27591
rect 6779 27557 6788 27591
rect 6736 27548 6788 27557
rect 7380 27548 7432 27600
rect 8944 27616 8996 27668
rect 848 27319 900 27328
rect 848 27285 857 27319
rect 857 27285 891 27319
rect 891 27285 900 27319
rect 848 27276 900 27285
rect 1124 27276 1176 27328
rect 1216 27276 1268 27328
rect 1676 27276 1728 27328
rect 2596 27276 2648 27328
rect 2780 27276 2832 27328
rect 3240 27276 3292 27328
rect 5448 27412 5500 27464
rect 6276 27480 6328 27532
rect 7196 27480 7248 27532
rect 7656 27480 7708 27532
rect 4160 27276 4212 27328
rect 5264 27344 5316 27396
rect 5356 27344 5408 27396
rect 6920 27412 6972 27464
rect 8024 27412 8076 27464
rect 8576 27412 8628 27464
rect 9128 27480 9180 27532
rect 9680 27548 9732 27600
rect 11244 27548 11296 27600
rect 4988 27276 5040 27328
rect 5816 27276 5868 27328
rect 8300 27344 8352 27396
rect 8760 27344 8812 27396
rect 8944 27344 8996 27396
rect 6184 27276 6236 27328
rect 7656 27319 7708 27328
rect 7656 27285 7665 27319
rect 7665 27285 7699 27319
rect 7699 27285 7708 27319
rect 7656 27276 7708 27285
rect 8116 27276 8168 27328
rect 9496 27276 9548 27328
rect 10692 27276 10744 27328
rect 3662 27174 3714 27226
rect 3726 27174 3778 27226
rect 3790 27174 3842 27226
rect 3854 27174 3906 27226
rect 3918 27174 3970 27226
rect 10062 27174 10114 27226
rect 10126 27174 10178 27226
rect 10190 27174 10242 27226
rect 10254 27174 10306 27226
rect 10318 27174 10370 27226
rect 1216 27072 1268 27124
rect 2688 27072 2740 27124
rect 2780 27072 2832 27124
rect 3424 27072 3476 27124
rect 4252 27072 4304 27124
rect 4712 27072 4764 27124
rect 6920 27072 6972 27124
rect 7196 27072 7248 27124
rect 7288 27072 7340 27124
rect 7472 27072 7524 27124
rect 10140 27072 10192 27124
rect 848 26936 900 26988
rect 1032 26732 1084 26784
rect 1308 26868 1360 26920
rect 1860 26936 1912 26988
rect 2412 26936 2464 26988
rect 4068 27004 4120 27056
rect 2596 26979 2648 26988
rect 2596 26945 2605 26979
rect 2605 26945 2639 26979
rect 2639 26945 2648 26979
rect 2596 26936 2648 26945
rect 3516 26936 3568 26988
rect 4528 26936 4580 26988
rect 7380 27004 7432 27056
rect 8024 27004 8076 27056
rect 1768 26800 1820 26852
rect 2412 26800 2464 26852
rect 3608 26911 3660 26920
rect 3608 26877 3617 26911
rect 3617 26877 3651 26911
rect 3651 26877 3660 26911
rect 3608 26868 3660 26877
rect 4068 26911 4120 26920
rect 4068 26877 4077 26911
rect 4077 26877 4111 26911
rect 4111 26877 4120 26911
rect 4068 26868 4120 26877
rect 4344 26911 4396 26920
rect 4344 26877 4353 26911
rect 4353 26877 4387 26911
rect 4387 26877 4396 26911
rect 4344 26868 4396 26877
rect 1216 26732 1268 26784
rect 2504 26732 2556 26784
rect 3700 26800 3752 26852
rect 5540 26868 5592 26920
rect 6368 26936 6420 26988
rect 6460 26868 6512 26920
rect 6736 26868 6788 26920
rect 7748 26936 7800 26988
rect 8944 26936 8996 26988
rect 9312 26936 9364 26988
rect 6920 26911 6972 26920
rect 6920 26877 6929 26911
rect 6929 26877 6963 26911
rect 6963 26877 6972 26911
rect 6920 26868 6972 26877
rect 7104 26868 7156 26920
rect 7196 26911 7248 26920
rect 7196 26877 7205 26911
rect 7205 26877 7239 26911
rect 7239 26877 7248 26911
rect 7196 26868 7248 26877
rect 8024 26868 8076 26920
rect 8300 26868 8352 26920
rect 8576 26868 8628 26920
rect 8852 26911 8904 26920
rect 8852 26877 8861 26911
rect 8861 26877 8895 26911
rect 8895 26877 8904 26911
rect 8852 26868 8904 26877
rect 9036 26911 9088 26920
rect 9036 26877 9045 26911
rect 9045 26877 9079 26911
rect 9079 26877 9088 26911
rect 9036 26868 9088 26877
rect 9128 26911 9180 26920
rect 9128 26877 9137 26911
rect 9137 26877 9171 26911
rect 9171 26877 9180 26911
rect 9128 26868 9180 26877
rect 4712 26800 4764 26852
rect 4896 26843 4948 26852
rect 4896 26809 4905 26843
rect 4905 26809 4939 26843
rect 4939 26809 4948 26843
rect 4896 26800 4948 26809
rect 5080 26800 5132 26852
rect 4620 26732 4672 26784
rect 6000 26843 6052 26852
rect 6000 26809 6009 26843
rect 6009 26809 6043 26843
rect 6043 26809 6052 26843
rect 6000 26800 6052 26809
rect 6276 26800 6328 26852
rect 7656 26843 7708 26852
rect 7656 26809 7665 26843
rect 7665 26809 7699 26843
rect 7699 26809 7708 26843
rect 7656 26800 7708 26809
rect 7748 26800 7800 26852
rect 8208 26800 8260 26852
rect 5632 26732 5684 26784
rect 6368 26732 6420 26784
rect 6644 26775 6696 26784
rect 6644 26741 6653 26775
rect 6653 26741 6687 26775
rect 6687 26741 6696 26775
rect 6644 26732 6696 26741
rect 6736 26732 6788 26784
rect 7196 26732 7248 26784
rect 7288 26775 7340 26784
rect 7288 26741 7297 26775
rect 7297 26741 7331 26775
rect 7331 26741 7340 26775
rect 7288 26732 7340 26741
rect 9128 26732 9180 26784
rect 9680 26868 9732 26920
rect 10508 26843 10560 26852
rect 10508 26809 10526 26843
rect 10526 26809 10560 26843
rect 10508 26800 10560 26809
rect 11336 26732 11388 26784
rect 4322 26630 4374 26682
rect 4386 26630 4438 26682
rect 4450 26630 4502 26682
rect 4514 26630 4566 26682
rect 4578 26630 4630 26682
rect 10722 26630 10774 26682
rect 10786 26630 10838 26682
rect 10850 26630 10902 26682
rect 10914 26630 10966 26682
rect 10978 26630 11030 26682
rect 1124 26528 1176 26580
rect 1676 26528 1728 26580
rect 2044 26571 2096 26580
rect 2044 26537 2053 26571
rect 2053 26537 2087 26571
rect 2087 26537 2096 26571
rect 2044 26528 2096 26537
rect 2780 26528 2832 26580
rect 3700 26528 3752 26580
rect 4068 26528 4120 26580
rect 4620 26528 4672 26580
rect 4712 26528 4764 26580
rect 5264 26528 5316 26580
rect 5356 26528 5408 26580
rect 5540 26528 5592 26580
rect 6000 26528 6052 26580
rect 7748 26528 7800 26580
rect 9036 26528 9088 26580
rect 9312 26528 9364 26580
rect 4528 26460 4580 26512
rect 5632 26460 5684 26512
rect 6368 26460 6420 26512
rect 848 26435 900 26444
rect 848 26401 857 26435
rect 857 26401 891 26435
rect 891 26401 900 26435
rect 848 26392 900 26401
rect 1032 26435 1084 26444
rect 1032 26401 1041 26435
rect 1041 26401 1075 26435
rect 1075 26401 1084 26435
rect 1032 26392 1084 26401
rect 1400 26435 1452 26444
rect 1400 26401 1409 26435
rect 1409 26401 1443 26435
rect 1443 26401 1452 26435
rect 1400 26392 1452 26401
rect 1676 26435 1728 26444
rect 1676 26401 1685 26435
rect 1685 26401 1719 26435
rect 1719 26401 1728 26435
rect 1676 26392 1728 26401
rect 1952 26435 2004 26444
rect 1952 26401 1961 26435
rect 1961 26401 1995 26435
rect 1995 26401 2004 26435
rect 1952 26392 2004 26401
rect 2044 26392 2096 26444
rect 2228 26435 2280 26444
rect 2228 26401 2237 26435
rect 2237 26401 2271 26435
rect 2271 26401 2280 26435
rect 2228 26392 2280 26401
rect 2504 26435 2556 26444
rect 2504 26401 2513 26435
rect 2513 26401 2547 26435
rect 2547 26401 2556 26435
rect 2504 26392 2556 26401
rect 2412 26324 2464 26376
rect 1400 26256 1452 26308
rect 2136 26256 2188 26308
rect 2228 26256 2280 26308
rect 4712 26392 4764 26444
rect 5080 26435 5132 26444
rect 5080 26401 5089 26435
rect 5089 26401 5123 26435
rect 5123 26401 5132 26435
rect 5080 26392 5132 26401
rect 5356 26435 5408 26444
rect 5356 26401 5365 26435
rect 5365 26401 5399 26435
rect 5399 26401 5408 26435
rect 5356 26392 5408 26401
rect 3056 26324 3108 26376
rect 6092 26392 6144 26444
rect 6276 26392 6328 26444
rect 7012 26503 7064 26512
rect 7012 26469 7021 26503
rect 7021 26469 7055 26503
rect 7055 26469 7064 26503
rect 7012 26460 7064 26469
rect 6644 26435 6696 26444
rect 6644 26401 6653 26435
rect 6653 26401 6687 26435
rect 6687 26401 6696 26435
rect 6644 26392 6696 26401
rect 7196 26435 7248 26444
rect 7196 26401 7205 26435
rect 7205 26401 7239 26435
rect 7239 26401 7248 26435
rect 7196 26392 7248 26401
rect 7564 26392 7616 26444
rect 8668 26460 8720 26512
rect 9588 26460 9640 26512
rect 5540 26324 5592 26376
rect 1124 26188 1176 26240
rect 1492 26231 1544 26240
rect 1492 26197 1501 26231
rect 1501 26197 1535 26231
rect 1535 26197 1544 26231
rect 1492 26188 1544 26197
rect 1952 26188 2004 26240
rect 2320 26188 2372 26240
rect 2688 26188 2740 26240
rect 3608 26231 3660 26240
rect 3608 26197 3617 26231
rect 3617 26197 3651 26231
rect 3651 26197 3660 26231
rect 3608 26188 3660 26197
rect 3792 26256 3844 26308
rect 6736 26324 6788 26376
rect 6276 26256 6328 26308
rect 6460 26256 6512 26308
rect 8116 26392 8168 26444
rect 8300 26392 8352 26444
rect 9036 26392 9088 26444
rect 9312 26435 9364 26444
rect 9312 26401 9321 26435
rect 9321 26401 9355 26435
rect 9355 26401 9364 26435
rect 9312 26392 9364 26401
rect 5540 26231 5592 26240
rect 5540 26197 5549 26231
rect 5549 26197 5583 26231
rect 5583 26197 5592 26231
rect 5540 26188 5592 26197
rect 6368 26188 6420 26240
rect 7196 26188 7248 26240
rect 7472 26188 7524 26240
rect 8576 26256 8628 26308
rect 9220 26256 9272 26308
rect 9312 26188 9364 26240
rect 10140 26392 10192 26444
rect 11244 26392 11296 26444
rect 9956 26256 10008 26308
rect 10048 26188 10100 26240
rect 10508 26188 10560 26240
rect 3662 26086 3714 26138
rect 3726 26086 3778 26138
rect 3790 26086 3842 26138
rect 3854 26086 3906 26138
rect 3918 26086 3970 26138
rect 10062 26086 10114 26138
rect 10126 26086 10178 26138
rect 10190 26086 10242 26138
rect 10254 26086 10306 26138
rect 10318 26086 10370 26138
rect 1400 25984 1452 26036
rect 2320 25984 2372 26036
rect 3516 25984 3568 26036
rect 1584 25916 1636 25968
rect 1400 25848 1452 25900
rect 1492 25848 1544 25900
rect 2504 25916 2556 25968
rect 2596 25916 2648 25968
rect 3056 25916 3108 25968
rect 3240 25959 3292 25968
rect 3240 25925 3249 25959
rect 3249 25925 3283 25959
rect 3283 25925 3292 25959
rect 3240 25916 3292 25925
rect 1308 25780 1360 25832
rect 848 25712 900 25764
rect 2228 25823 2280 25832
rect 2228 25789 2237 25823
rect 2237 25789 2271 25823
rect 2271 25789 2280 25823
rect 2228 25780 2280 25789
rect 2320 25780 2372 25832
rect 2504 25823 2556 25832
rect 2504 25789 2513 25823
rect 2513 25789 2547 25823
rect 2547 25789 2556 25823
rect 2504 25780 2556 25789
rect 2596 25823 2648 25832
rect 2596 25789 2624 25823
rect 2624 25789 2648 25823
rect 2596 25780 2648 25789
rect 3424 25848 3476 25900
rect 3608 25848 3660 25900
rect 1584 25644 1636 25696
rect 1768 25644 1820 25696
rect 2964 25780 3016 25832
rect 3884 25916 3936 25968
rect 4252 25984 4304 26036
rect 4988 25916 5040 25968
rect 5724 25916 5776 25968
rect 6644 25984 6696 26036
rect 6736 25984 6788 26036
rect 7012 25984 7064 26036
rect 6184 25916 6236 25968
rect 5908 25848 5960 25900
rect 6736 25848 6788 25900
rect 3056 25644 3108 25696
rect 3240 25644 3292 25696
rect 3792 25823 3844 25832
rect 3792 25789 3801 25823
rect 3801 25789 3835 25823
rect 3835 25789 3844 25823
rect 3792 25780 3844 25789
rect 3884 25780 3936 25832
rect 4436 25712 4488 25764
rect 3884 25644 3936 25696
rect 4712 25780 4764 25832
rect 4988 25823 5040 25832
rect 4988 25789 4997 25823
rect 4997 25789 5031 25823
rect 5031 25789 5040 25823
rect 4988 25780 5040 25789
rect 4896 25712 4948 25764
rect 4804 25644 4856 25696
rect 5724 25780 5776 25832
rect 6092 25823 6144 25832
rect 6092 25789 6101 25823
rect 6101 25789 6135 25823
rect 6135 25789 6144 25823
rect 6092 25780 6144 25789
rect 6552 25780 6604 25832
rect 6644 25780 6696 25832
rect 8208 25984 8260 26036
rect 8300 25984 8352 26036
rect 9588 25984 9640 26036
rect 7564 25916 7616 25968
rect 7288 25848 7340 25900
rect 9036 25916 9088 25968
rect 10048 25916 10100 25968
rect 7196 25823 7248 25832
rect 7196 25789 7205 25823
rect 7205 25789 7239 25823
rect 7239 25789 7248 25823
rect 7196 25780 7248 25789
rect 7380 25712 7432 25764
rect 5724 25644 5776 25696
rect 6552 25687 6604 25696
rect 6552 25653 6561 25687
rect 6561 25653 6595 25687
rect 6595 25653 6604 25687
rect 6552 25644 6604 25653
rect 6736 25644 6788 25696
rect 7288 25644 7340 25696
rect 7564 25823 7616 25832
rect 7564 25789 7573 25823
rect 7573 25789 7607 25823
rect 7607 25789 7616 25823
rect 8392 25848 8444 25900
rect 7564 25780 7616 25789
rect 7840 25823 7892 25832
rect 7840 25789 7849 25823
rect 7849 25789 7883 25823
rect 7883 25789 7892 25823
rect 7840 25780 7892 25789
rect 8484 25823 8536 25832
rect 8484 25789 8493 25823
rect 8493 25789 8527 25823
rect 8527 25789 8536 25823
rect 8484 25780 8536 25789
rect 10508 25823 10560 25832
rect 10508 25789 10517 25823
rect 10517 25789 10551 25823
rect 10551 25789 10560 25823
rect 10508 25780 10560 25789
rect 10600 25780 10652 25832
rect 8024 25687 8076 25696
rect 8024 25653 8033 25687
rect 8033 25653 8067 25687
rect 8067 25653 8076 25687
rect 8024 25644 8076 25653
rect 9036 25644 9088 25696
rect 4322 25542 4374 25594
rect 4386 25542 4438 25594
rect 4450 25542 4502 25594
rect 4514 25542 4566 25594
rect 4578 25542 4630 25594
rect 10722 25542 10774 25594
rect 10786 25542 10838 25594
rect 10850 25542 10902 25594
rect 10914 25542 10966 25594
rect 10978 25542 11030 25594
rect 2504 25440 2556 25492
rect 2964 25440 3016 25492
rect 1584 25372 1636 25424
rect 940 25304 992 25356
rect 1492 25304 1544 25356
rect 1124 25279 1176 25288
rect 1124 25245 1133 25279
rect 1133 25245 1167 25279
rect 1167 25245 1176 25279
rect 1124 25236 1176 25245
rect 1216 25279 1268 25288
rect 1216 25245 1225 25279
rect 1225 25245 1259 25279
rect 1259 25245 1268 25279
rect 1216 25236 1268 25245
rect 848 25168 900 25220
rect 1584 25168 1636 25220
rect 2228 25347 2280 25356
rect 2228 25313 2237 25347
rect 2237 25313 2271 25347
rect 2271 25313 2280 25347
rect 2228 25304 2280 25313
rect 2412 25372 2464 25424
rect 2780 25372 2832 25424
rect 2964 25304 3016 25356
rect 3056 25347 3108 25356
rect 3056 25313 3065 25347
rect 3065 25313 3099 25347
rect 3099 25313 3108 25347
rect 3056 25304 3108 25313
rect 2136 25236 2188 25288
rect 2780 25279 2832 25288
rect 2780 25245 2789 25279
rect 2789 25245 2823 25279
rect 2823 25245 2832 25279
rect 2780 25236 2832 25245
rect 3700 25372 3752 25424
rect 4620 25483 4672 25492
rect 4620 25449 4629 25483
rect 4629 25449 4663 25483
rect 4663 25449 4672 25483
rect 4620 25440 4672 25449
rect 4804 25483 4856 25492
rect 4804 25449 4813 25483
rect 4813 25449 4847 25483
rect 4847 25449 4856 25483
rect 4804 25440 4856 25449
rect 5540 25440 5592 25492
rect 6920 25440 6972 25492
rect 7288 25440 7340 25492
rect 7656 25440 7708 25492
rect 8484 25440 8536 25492
rect 8576 25483 8628 25492
rect 8576 25449 8585 25483
rect 8585 25449 8619 25483
rect 8619 25449 8628 25483
rect 8576 25440 8628 25449
rect 8852 25440 8904 25492
rect 9496 25440 9548 25492
rect 9772 25440 9824 25492
rect 3424 25347 3476 25356
rect 3424 25313 3433 25347
rect 3433 25313 3467 25347
rect 3467 25313 3476 25347
rect 3424 25304 3476 25313
rect 3976 25347 4028 25356
rect 3976 25313 3985 25347
rect 3985 25313 4019 25347
rect 4019 25313 4028 25347
rect 3976 25304 4028 25313
rect 3608 25236 3660 25288
rect 3700 25236 3752 25288
rect 6184 25372 6236 25424
rect 6736 25372 6788 25424
rect 4620 25236 4672 25288
rect 4896 25236 4948 25288
rect 5356 25347 5408 25356
rect 5356 25313 5365 25347
rect 5365 25313 5399 25347
rect 5399 25313 5408 25347
rect 5356 25304 5408 25313
rect 6276 25347 6328 25356
rect 6276 25313 6285 25347
rect 6285 25313 6319 25347
rect 6319 25313 6328 25347
rect 6276 25304 6328 25313
rect 6644 25347 6696 25356
rect 6644 25313 6653 25347
rect 6653 25313 6687 25347
rect 6687 25313 6696 25347
rect 6644 25304 6696 25313
rect 6552 25236 6604 25288
rect 1400 25100 1452 25152
rect 4160 25168 4212 25220
rect 5356 25168 5408 25220
rect 4436 25143 4488 25152
rect 4436 25109 4445 25143
rect 4445 25109 4479 25143
rect 4479 25109 4488 25143
rect 4436 25100 4488 25109
rect 4988 25143 5040 25152
rect 4988 25109 4997 25143
rect 4997 25109 5031 25143
rect 5031 25109 5040 25143
rect 4988 25100 5040 25109
rect 5908 25100 5960 25152
rect 6184 25211 6236 25220
rect 6184 25177 6193 25211
rect 6193 25177 6227 25211
rect 6227 25177 6236 25211
rect 6184 25168 6236 25177
rect 7012 25347 7064 25356
rect 7012 25313 7021 25347
rect 7021 25313 7055 25347
rect 7055 25313 7064 25347
rect 7012 25304 7064 25313
rect 7196 25347 7248 25356
rect 7196 25313 7205 25347
rect 7205 25313 7239 25347
rect 7239 25313 7248 25347
rect 7196 25304 7248 25313
rect 7564 25304 7616 25356
rect 7656 25338 7708 25390
rect 7748 25347 7800 25356
rect 7748 25313 7757 25347
rect 7757 25313 7791 25347
rect 7791 25313 7800 25347
rect 7748 25304 7800 25313
rect 8392 25304 8444 25356
rect 8576 25304 8628 25356
rect 9128 25347 9180 25356
rect 9128 25313 9137 25347
rect 9137 25313 9171 25347
rect 9171 25313 9180 25347
rect 9128 25304 9180 25313
rect 10508 25304 10560 25356
rect 7380 25236 7432 25288
rect 7932 25168 7984 25220
rect 8024 25168 8076 25220
rect 8760 25236 8812 25288
rect 9128 25168 9180 25220
rect 10048 25168 10100 25220
rect 7656 25100 7708 25152
rect 11060 25100 11112 25152
rect 3662 24998 3714 25050
rect 3726 24998 3778 25050
rect 3790 24998 3842 25050
rect 3854 24998 3906 25050
rect 3918 24998 3970 25050
rect 10062 24998 10114 25050
rect 10126 24998 10178 25050
rect 10190 24998 10242 25050
rect 10254 24998 10306 25050
rect 10318 24998 10370 25050
rect 1308 24896 1360 24948
rect 3424 24896 3476 24948
rect 3976 24896 4028 24948
rect 4160 24896 4212 24948
rect 4804 24896 4856 24948
rect 1400 24760 1452 24812
rect 1492 24803 1544 24812
rect 1492 24769 1501 24803
rect 1501 24769 1535 24803
rect 1535 24769 1544 24803
rect 1492 24760 1544 24769
rect 2504 24760 2556 24812
rect 664 24624 716 24676
rect 1492 24624 1544 24676
rect 2228 24692 2280 24744
rect 2412 24735 2464 24744
rect 2412 24701 2421 24735
rect 2421 24701 2455 24735
rect 2455 24701 2464 24735
rect 2412 24692 2464 24701
rect 2780 24828 2832 24880
rect 4712 24828 4764 24880
rect 4620 24760 4672 24812
rect 5264 24896 5316 24948
rect 6460 24896 6512 24948
rect 7012 24896 7064 24948
rect 4988 24828 5040 24880
rect 5540 24828 5592 24880
rect 3332 24692 3384 24744
rect 3424 24735 3476 24744
rect 3424 24701 3433 24735
rect 3433 24701 3467 24735
rect 3467 24701 3476 24735
rect 3424 24692 3476 24701
rect 2780 24624 2832 24676
rect 3700 24735 3752 24744
rect 3700 24701 3709 24735
rect 3709 24701 3743 24735
rect 3743 24701 3752 24735
rect 3700 24692 3752 24701
rect 4068 24692 4120 24744
rect 4160 24692 4212 24744
rect 5724 24760 5776 24812
rect 6276 24828 6328 24880
rect 4804 24735 4856 24744
rect 4804 24701 4813 24735
rect 4813 24701 4847 24735
rect 4847 24701 4856 24735
rect 4804 24692 4856 24701
rect 3884 24667 3936 24676
rect 3884 24633 3893 24667
rect 3893 24633 3927 24667
rect 3927 24633 3936 24667
rect 3884 24624 3936 24633
rect 5632 24692 5684 24744
rect 5356 24624 5408 24676
rect 5724 24624 5776 24676
rect 6276 24624 6328 24676
rect 7196 24735 7248 24744
rect 7196 24701 7205 24735
rect 7205 24701 7239 24735
rect 7239 24701 7248 24735
rect 7196 24692 7248 24701
rect 7288 24692 7340 24744
rect 7472 24735 7524 24744
rect 7472 24701 7481 24735
rect 7481 24701 7515 24735
rect 7515 24701 7524 24735
rect 7472 24692 7524 24701
rect 7656 24692 7708 24744
rect 7840 24692 7892 24744
rect 7932 24735 7984 24744
rect 7932 24701 7941 24735
rect 7941 24701 7975 24735
rect 7975 24701 7984 24735
rect 7932 24692 7984 24701
rect 8576 24828 8628 24880
rect 8852 24828 8904 24880
rect 9680 24828 9732 24880
rect 10232 24828 10284 24880
rect 8392 24760 8444 24812
rect 10324 24803 10376 24812
rect 10324 24769 10333 24803
rect 10333 24769 10367 24803
rect 10367 24769 10376 24803
rect 10324 24760 10376 24769
rect 10508 24760 10560 24812
rect 9680 24692 9732 24744
rect 10048 24735 10100 24744
rect 10048 24701 10057 24735
rect 10057 24701 10091 24735
rect 10091 24701 10100 24735
rect 10048 24692 10100 24701
rect 10600 24735 10652 24744
rect 10600 24701 10609 24735
rect 10609 24701 10643 24735
rect 10643 24701 10652 24735
rect 10600 24692 10652 24701
rect 8392 24667 8444 24676
rect 8392 24633 8401 24667
rect 8401 24633 8435 24667
rect 8435 24633 8444 24667
rect 8392 24624 8444 24633
rect 8484 24624 8536 24676
rect 8668 24624 8720 24676
rect 9220 24667 9272 24676
rect 9220 24633 9229 24667
rect 9229 24633 9263 24667
rect 9263 24633 9272 24667
rect 9220 24624 9272 24633
rect 9588 24624 9640 24676
rect 10140 24624 10192 24676
rect 10508 24624 10560 24676
rect 10968 24624 11020 24676
rect 388 24556 440 24608
rect 2504 24556 2556 24608
rect 2596 24556 2648 24608
rect 4988 24556 5040 24608
rect 5080 24599 5132 24608
rect 5080 24565 5089 24599
rect 5089 24565 5123 24599
rect 5123 24565 5132 24599
rect 5080 24556 5132 24565
rect 5632 24599 5684 24608
rect 5632 24565 5641 24599
rect 5641 24565 5675 24599
rect 5675 24565 5684 24599
rect 5632 24556 5684 24565
rect 6000 24556 6052 24608
rect 6552 24556 6604 24608
rect 7380 24556 7432 24608
rect 7656 24556 7708 24608
rect 8116 24556 8168 24608
rect 9312 24556 9364 24608
rect 9496 24556 9548 24608
rect 4322 24454 4374 24506
rect 4386 24454 4438 24506
rect 4450 24454 4502 24506
rect 4514 24454 4566 24506
rect 4578 24454 4630 24506
rect 10722 24454 10774 24506
rect 10786 24454 10838 24506
rect 10850 24454 10902 24506
rect 10914 24454 10966 24506
rect 10978 24454 11030 24506
rect 112 24352 164 24404
rect 664 24352 716 24404
rect 1032 24352 1084 24404
rect 1400 24284 1452 24336
rect 3884 24352 3936 24404
rect 4528 24352 4580 24404
rect 1308 24216 1360 24268
rect 1768 24259 1820 24268
rect 1768 24225 1777 24259
rect 1777 24225 1811 24259
rect 1811 24225 1820 24259
rect 1768 24216 1820 24225
rect 2504 24259 2556 24268
rect 2504 24225 2513 24259
rect 2513 24225 2547 24259
rect 2547 24225 2556 24259
rect 2504 24216 2556 24225
rect 2596 24216 2648 24268
rect 3332 24284 3384 24336
rect 4068 24284 4120 24336
rect 4712 24284 4764 24336
rect 5264 24327 5316 24336
rect 5264 24293 5273 24327
rect 5273 24293 5307 24327
rect 5307 24293 5316 24327
rect 5264 24284 5316 24293
rect 5356 24327 5408 24336
rect 5356 24293 5365 24327
rect 5365 24293 5399 24327
rect 5399 24293 5408 24327
rect 5356 24284 5408 24293
rect 6644 24352 6696 24404
rect 6920 24395 6972 24404
rect 6920 24361 6929 24395
rect 6929 24361 6963 24395
rect 6963 24361 6972 24395
rect 6920 24352 6972 24361
rect 7012 24352 7064 24404
rect 6368 24284 6420 24336
rect 3516 24216 3568 24268
rect 2228 24191 2280 24200
rect 2228 24157 2237 24191
rect 2237 24157 2271 24191
rect 2271 24157 2280 24191
rect 2228 24148 2280 24157
rect 2964 24148 3016 24200
rect 3332 24148 3384 24200
rect 4804 24259 4856 24268
rect 4804 24225 4813 24259
rect 4813 24225 4847 24259
rect 4847 24225 4856 24259
rect 4804 24216 4856 24225
rect 848 24080 900 24132
rect 2596 24012 2648 24064
rect 3056 24123 3108 24132
rect 3056 24089 3065 24123
rect 3065 24089 3099 24123
rect 3099 24089 3108 24123
rect 3056 24080 3108 24089
rect 3700 24191 3752 24200
rect 3700 24157 3709 24191
rect 3709 24157 3743 24191
rect 3743 24157 3752 24191
rect 3700 24148 3752 24157
rect 4068 24148 4120 24200
rect 3884 24080 3936 24132
rect 3976 24080 4028 24132
rect 4988 24148 5040 24200
rect 4712 24080 4764 24132
rect 5356 24148 5408 24200
rect 6184 24259 6236 24268
rect 6184 24225 6193 24259
rect 6193 24225 6227 24259
rect 6227 24225 6236 24259
rect 6184 24216 6236 24225
rect 6552 24216 6604 24268
rect 7012 24216 7064 24268
rect 7196 24259 7248 24268
rect 7196 24225 7205 24259
rect 7205 24225 7239 24259
rect 7239 24225 7248 24259
rect 7196 24216 7248 24225
rect 7288 24250 7340 24302
rect 6092 24148 6144 24200
rect 6368 24191 6420 24200
rect 6368 24157 6377 24191
rect 6377 24157 6411 24191
rect 6411 24157 6420 24191
rect 6368 24148 6420 24157
rect 7288 24148 7340 24200
rect 7472 24259 7524 24268
rect 7472 24225 7481 24259
rect 7481 24225 7515 24259
rect 7515 24225 7524 24259
rect 7472 24216 7524 24225
rect 8576 24352 8628 24404
rect 9864 24352 9916 24404
rect 11244 24352 11296 24404
rect 8944 24327 8996 24336
rect 8944 24293 8953 24327
rect 8953 24293 8987 24327
rect 8987 24293 8996 24327
rect 8944 24284 8996 24293
rect 9036 24327 9088 24336
rect 9036 24293 9045 24327
rect 9045 24293 9079 24327
rect 9079 24293 9088 24327
rect 9036 24284 9088 24293
rect 9772 24284 9824 24336
rect 7840 24148 7892 24200
rect 3608 24012 3660 24064
rect 4436 24055 4488 24064
rect 4436 24021 4445 24055
rect 4445 24021 4479 24055
rect 4479 24021 4488 24055
rect 4436 24012 4488 24021
rect 4528 24012 4580 24064
rect 5080 24012 5132 24064
rect 5908 24080 5960 24132
rect 6736 24080 6788 24132
rect 8760 24259 8812 24268
rect 8760 24225 8769 24259
rect 8769 24225 8803 24259
rect 8803 24225 8812 24259
rect 8760 24216 8812 24225
rect 9128 24259 9180 24268
rect 9128 24225 9169 24259
rect 9169 24225 9180 24259
rect 9128 24216 9180 24225
rect 9496 24216 9548 24268
rect 9588 24216 9640 24268
rect 10416 24216 10468 24268
rect 9312 24148 9364 24200
rect 9864 24148 9916 24200
rect 10140 24148 10192 24200
rect 11244 24148 11296 24200
rect 8116 24080 8168 24132
rect 8852 24080 8904 24132
rect 9036 24080 9088 24132
rect 6368 24012 6420 24064
rect 7288 24012 7340 24064
rect 8392 24012 8444 24064
rect 9220 24012 9272 24064
rect 9496 24055 9548 24064
rect 9496 24021 9505 24055
rect 9505 24021 9539 24055
rect 9539 24021 9548 24055
rect 9496 24012 9548 24021
rect 9864 24012 9916 24064
rect 10232 24012 10284 24064
rect 10600 24012 10652 24064
rect 3662 23910 3714 23962
rect 3726 23910 3778 23962
rect 3790 23910 3842 23962
rect 3854 23910 3906 23962
rect 3918 23910 3970 23962
rect 10062 23910 10114 23962
rect 10126 23910 10178 23962
rect 10190 23910 10242 23962
rect 10254 23910 10306 23962
rect 10318 23910 10370 23962
rect 2412 23808 2464 23860
rect 5080 23851 5132 23860
rect 5080 23817 5089 23851
rect 5089 23817 5123 23851
rect 5123 23817 5132 23851
rect 5080 23808 5132 23817
rect 5448 23808 5500 23860
rect 2504 23740 2556 23792
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 5356 23740 5408 23792
rect 6552 23740 6604 23792
rect 6644 23740 6696 23792
rect 2228 23647 2280 23656
rect 2228 23613 2237 23647
rect 2237 23613 2271 23647
rect 2271 23613 2280 23647
rect 2228 23604 2280 23613
rect 3056 23604 3108 23656
rect 1400 23536 1452 23588
rect 2320 23536 2372 23588
rect 3608 23647 3660 23656
rect 3608 23613 3617 23647
rect 3617 23613 3651 23647
rect 3651 23613 3660 23647
rect 3608 23604 3660 23613
rect 4068 23647 4120 23656
rect 4068 23613 4077 23647
rect 4077 23613 4111 23647
rect 4111 23613 4120 23647
rect 4068 23604 4120 23613
rect 7472 23808 7524 23860
rect 7840 23808 7892 23860
rect 7104 23672 7156 23724
rect 4436 23536 4488 23588
rect 5080 23604 5132 23656
rect 2780 23468 2832 23520
rect 3792 23468 3844 23520
rect 4804 23468 4856 23520
rect 5264 23647 5316 23656
rect 5264 23613 5273 23647
rect 5273 23613 5307 23647
rect 5307 23613 5316 23647
rect 5264 23604 5316 23613
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 5724 23536 5776 23588
rect 5448 23468 5500 23520
rect 5632 23468 5684 23520
rect 5908 23468 5960 23520
rect 6276 23579 6328 23588
rect 6276 23545 6285 23579
rect 6285 23545 6319 23579
rect 6319 23545 6328 23579
rect 6276 23536 6328 23545
rect 6552 23604 6604 23656
rect 6644 23647 6696 23656
rect 6644 23613 6653 23647
rect 6653 23613 6687 23647
rect 6687 23613 6696 23647
rect 6644 23604 6696 23613
rect 7748 23715 7800 23724
rect 7748 23681 7757 23715
rect 7757 23681 7791 23715
rect 7791 23681 7800 23715
rect 7748 23672 7800 23681
rect 7288 23647 7340 23656
rect 7288 23613 7297 23647
rect 7297 23613 7331 23647
rect 7331 23613 7340 23647
rect 7288 23604 7340 23613
rect 6920 23536 6972 23588
rect 7196 23536 7248 23588
rect 7840 23536 7892 23588
rect 8208 23808 8260 23860
rect 8392 23851 8444 23860
rect 8392 23817 8401 23851
rect 8401 23817 8435 23851
rect 8435 23817 8444 23851
rect 8392 23808 8444 23817
rect 8668 23740 8720 23792
rect 8760 23740 8812 23792
rect 8944 23740 8996 23792
rect 9036 23740 9088 23792
rect 9220 23740 9272 23792
rect 10140 23808 10192 23860
rect 10416 23808 10468 23860
rect 11336 23808 11388 23860
rect 6552 23468 6604 23520
rect 8116 23536 8168 23588
rect 8944 23647 8996 23656
rect 8944 23613 8953 23647
rect 8953 23613 8987 23647
rect 8987 23613 8996 23647
rect 8944 23604 8996 23613
rect 9036 23647 9088 23656
rect 9036 23613 9045 23647
rect 9045 23613 9079 23647
rect 9079 23613 9088 23647
rect 9036 23604 9088 23613
rect 9220 23647 9272 23656
rect 9220 23613 9229 23647
rect 9229 23613 9263 23647
rect 9263 23613 9272 23647
rect 9220 23604 9272 23613
rect 9588 23604 9640 23656
rect 8576 23468 8628 23520
rect 8944 23468 8996 23520
rect 9404 23579 9456 23588
rect 9404 23545 9413 23579
rect 9413 23545 9447 23579
rect 9447 23545 9456 23579
rect 9404 23536 9456 23545
rect 9588 23468 9640 23520
rect 9772 23604 9824 23656
rect 10140 23672 10192 23724
rect 10048 23647 10100 23656
rect 10048 23613 10057 23647
rect 10057 23613 10091 23647
rect 10091 23613 10100 23647
rect 10048 23604 10100 23613
rect 11060 23672 11112 23724
rect 10324 23604 10376 23656
rect 9772 23468 9824 23520
rect 9864 23511 9916 23520
rect 9864 23477 9873 23511
rect 9873 23477 9907 23511
rect 9907 23477 9916 23511
rect 9864 23468 9916 23477
rect 10692 23468 10744 23520
rect 11336 23468 11388 23520
rect 4322 23366 4374 23418
rect 4386 23366 4438 23418
rect 4450 23366 4502 23418
rect 4514 23366 4566 23418
rect 4578 23366 4630 23418
rect 10722 23366 10774 23418
rect 10786 23366 10838 23418
rect 10850 23366 10902 23418
rect 10914 23366 10966 23418
rect 10978 23366 11030 23418
rect 388 23264 440 23316
rect 848 23264 900 23316
rect 1308 23307 1360 23316
rect 1308 23273 1317 23307
rect 1317 23273 1351 23307
rect 1351 23273 1360 23307
rect 1308 23264 1360 23273
rect 1400 23264 1452 23316
rect 1584 23264 1636 23316
rect 2596 23264 2648 23316
rect 6276 23264 6328 23316
rect 480 23128 532 23180
rect 1216 23128 1268 23180
rect 3332 23196 3384 23248
rect 2044 23128 2096 23180
rect 2136 23171 2188 23180
rect 2136 23137 2145 23171
rect 2145 23137 2179 23171
rect 2179 23137 2188 23171
rect 2136 23128 2188 23137
rect 2228 23171 2280 23180
rect 2228 23137 2237 23171
rect 2237 23137 2271 23171
rect 2271 23137 2280 23171
rect 2228 23128 2280 23137
rect 2320 23171 2372 23180
rect 2320 23137 2329 23171
rect 2329 23137 2363 23171
rect 2363 23137 2372 23171
rect 2320 23128 2372 23137
rect 2412 23171 2464 23180
rect 2412 23137 2421 23171
rect 2421 23137 2455 23171
rect 2455 23137 2464 23171
rect 2412 23128 2464 23137
rect 1860 23060 1912 23112
rect 3424 23171 3476 23180
rect 3424 23137 3433 23171
rect 3433 23137 3467 23171
rect 3467 23137 3476 23171
rect 3424 23128 3476 23137
rect 3792 23171 3844 23180
rect 3792 23137 3801 23171
rect 3801 23137 3835 23171
rect 3835 23137 3844 23171
rect 3792 23128 3844 23137
rect 4068 23196 4120 23248
rect 4988 23196 5040 23248
rect 4620 23128 4672 23180
rect 4712 23171 4764 23180
rect 4712 23137 4721 23171
rect 4721 23137 4755 23171
rect 4755 23137 4764 23171
rect 4712 23128 4764 23137
rect 5080 23128 5132 23180
rect 5816 23171 5868 23180
rect 5816 23137 5825 23171
rect 5825 23137 5859 23171
rect 5859 23137 5868 23171
rect 5816 23128 5868 23137
rect 5908 23171 5960 23180
rect 5908 23137 5917 23171
rect 5917 23137 5951 23171
rect 5951 23137 5960 23171
rect 5908 23128 5960 23137
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 6184 23171 6236 23180
rect 6184 23137 6193 23171
rect 6193 23137 6227 23171
rect 6227 23137 6236 23171
rect 6184 23128 6236 23137
rect 7012 23264 7064 23316
rect 7748 23264 7800 23316
rect 7932 23264 7984 23316
rect 9036 23264 9088 23316
rect 9220 23307 9272 23316
rect 9220 23273 9229 23307
rect 9229 23273 9263 23307
rect 9263 23273 9272 23307
rect 9220 23264 9272 23273
rect 10324 23307 10376 23316
rect 10324 23273 10333 23307
rect 10333 23273 10367 23307
rect 10367 23273 10376 23307
rect 10324 23264 10376 23273
rect 4528 23060 4580 23112
rect 4804 23103 4856 23112
rect 4804 23069 4813 23103
rect 4813 23069 4847 23103
rect 4847 23069 4856 23103
rect 4804 23060 4856 23069
rect 5540 23103 5592 23112
rect 5540 23069 5549 23103
rect 5549 23069 5583 23103
rect 5583 23069 5592 23103
rect 5540 23060 5592 23069
rect 6828 23171 6880 23180
rect 6828 23137 6837 23171
rect 6837 23137 6871 23171
rect 6871 23137 6880 23171
rect 6828 23128 6880 23137
rect 7472 23196 7524 23248
rect 7288 23128 7340 23180
rect 6920 23060 6972 23112
rect 7564 23060 7616 23112
rect 7932 23171 7984 23180
rect 7932 23137 7941 23171
rect 7941 23137 7975 23171
rect 7975 23137 7984 23171
rect 7932 23128 7984 23137
rect 8208 23239 8260 23248
rect 8208 23205 8217 23239
rect 8217 23205 8251 23239
rect 8251 23205 8260 23239
rect 8208 23196 8260 23205
rect 2228 22992 2280 23044
rect 6276 22992 6328 23044
rect 8208 23060 8260 23112
rect 10692 23196 10744 23248
rect 8484 23171 8536 23180
rect 8484 23137 8493 23171
rect 8493 23137 8527 23171
rect 8527 23137 8536 23171
rect 8484 23128 8536 23137
rect 8576 23128 8628 23180
rect 8760 23171 8812 23180
rect 8760 23137 8769 23171
rect 8769 23137 8803 23171
rect 8803 23137 8812 23171
rect 8760 23128 8812 23137
rect 9036 23128 9088 23180
rect 9588 23171 9640 23180
rect 9588 23137 9597 23171
rect 9597 23137 9631 23171
rect 9631 23137 9640 23171
rect 9588 23128 9640 23137
rect 10140 23171 10192 23180
rect 10140 23137 10149 23171
rect 10149 23137 10183 23171
rect 10183 23137 10192 23171
rect 10140 23128 10192 23137
rect 9772 23060 9824 23112
rect 940 22967 992 22976
rect 940 22933 949 22967
rect 949 22933 983 22967
rect 983 22933 992 22967
rect 940 22924 992 22933
rect 1768 22967 1820 22976
rect 1768 22933 1777 22967
rect 1777 22933 1811 22967
rect 1811 22933 1820 22967
rect 1768 22924 1820 22933
rect 1860 22924 1912 22976
rect 2872 22924 2924 22976
rect 5080 22924 5132 22976
rect 6552 22924 6604 22976
rect 7288 22924 7340 22976
rect 7564 22924 7616 22976
rect 8484 22924 8536 22976
rect 10784 22992 10836 23044
rect 9588 22924 9640 22976
rect 10508 22924 10560 22976
rect 3662 22822 3714 22874
rect 3726 22822 3778 22874
rect 3790 22822 3842 22874
rect 3854 22822 3906 22874
rect 3918 22822 3970 22874
rect 10062 22822 10114 22874
rect 10126 22822 10178 22874
rect 10190 22822 10242 22874
rect 10254 22822 10306 22874
rect 10318 22822 10370 22874
rect 848 22720 900 22772
rect 1676 22720 1728 22772
rect 2412 22720 2464 22772
rect 204 22652 256 22704
rect 1308 22652 1360 22704
rect 756 22584 808 22636
rect 2596 22652 2648 22704
rect 3056 22652 3108 22704
rect 940 22516 992 22568
rect 1676 22559 1728 22568
rect 1676 22525 1685 22559
rect 1685 22525 1719 22559
rect 1719 22525 1728 22559
rect 1676 22516 1728 22525
rect 1768 22559 1820 22568
rect 1768 22525 1777 22559
rect 1777 22525 1811 22559
rect 1811 22525 1820 22559
rect 1768 22516 1820 22525
rect 2780 22584 2832 22636
rect 1216 22448 1268 22500
rect 3424 22516 3476 22568
rect 4436 22720 4488 22772
rect 5448 22652 5500 22704
rect 5908 22763 5960 22772
rect 5908 22729 5917 22763
rect 5917 22729 5951 22763
rect 5951 22729 5960 22763
rect 5908 22720 5960 22729
rect 6184 22720 6236 22772
rect 6644 22720 6696 22772
rect 7104 22720 7156 22772
rect 8760 22720 8812 22772
rect 10784 22720 10836 22772
rect 7380 22652 7432 22704
rect 7932 22652 7984 22704
rect 9680 22652 9732 22704
rect 3700 22584 3752 22636
rect 4160 22559 4212 22568
rect 4160 22525 4169 22559
rect 4169 22525 4203 22559
rect 4203 22525 4212 22559
rect 4160 22516 4212 22525
rect 4528 22584 4580 22636
rect 5724 22584 5776 22636
rect 5908 22584 5960 22636
rect 8208 22584 8260 22636
rect 8484 22584 8536 22636
rect 6184 22516 6236 22568
rect 6552 22559 6604 22568
rect 6552 22525 6561 22559
rect 6561 22525 6595 22559
rect 6595 22525 6604 22559
rect 6552 22516 6604 22525
rect 3516 22448 3568 22500
rect 4252 22448 4304 22500
rect 4620 22491 4672 22500
rect 4620 22457 4629 22491
rect 4629 22457 4663 22491
rect 4663 22457 4672 22491
rect 4620 22448 4672 22457
rect 5448 22448 5500 22500
rect 2504 22380 2556 22432
rect 2688 22380 2740 22432
rect 2872 22423 2924 22432
rect 2872 22389 2881 22423
rect 2881 22389 2915 22423
rect 2915 22389 2924 22423
rect 2872 22380 2924 22389
rect 3332 22380 3384 22432
rect 4068 22380 4120 22432
rect 4344 22380 4396 22432
rect 4712 22380 4764 22432
rect 4988 22380 5040 22432
rect 5264 22380 5316 22432
rect 7196 22516 7248 22568
rect 6736 22491 6788 22500
rect 6736 22457 6745 22491
rect 6745 22457 6779 22491
rect 6779 22457 6788 22491
rect 6736 22448 6788 22457
rect 7656 22448 7708 22500
rect 7840 22559 7892 22568
rect 7840 22525 7849 22559
rect 7849 22525 7883 22559
rect 7883 22525 7892 22559
rect 7840 22516 7892 22525
rect 7932 22516 7984 22568
rect 8576 22559 8628 22568
rect 8576 22525 8585 22559
rect 8585 22525 8619 22559
rect 8619 22525 8628 22559
rect 8576 22516 8628 22525
rect 9220 22584 9272 22636
rect 10508 22627 10560 22636
rect 10508 22593 10517 22627
rect 10517 22593 10551 22627
rect 10551 22593 10560 22627
rect 10508 22584 10560 22593
rect 9128 22559 9180 22568
rect 9128 22525 9137 22559
rect 9137 22525 9171 22559
rect 9171 22525 9180 22559
rect 9128 22516 9180 22525
rect 6552 22380 6604 22432
rect 6644 22380 6696 22432
rect 7104 22380 7156 22432
rect 7196 22423 7248 22432
rect 7196 22389 7205 22423
rect 7205 22389 7239 22423
rect 7239 22389 7248 22423
rect 7196 22380 7248 22389
rect 7472 22380 7524 22432
rect 8484 22423 8536 22432
rect 8484 22389 8493 22423
rect 8493 22389 8527 22423
rect 8527 22389 8536 22423
rect 8484 22380 8536 22389
rect 8944 22380 8996 22432
rect 10416 22516 10468 22568
rect 11336 22516 11388 22568
rect 4322 22278 4374 22330
rect 4386 22278 4438 22330
rect 4450 22278 4502 22330
rect 4514 22278 4566 22330
rect 4578 22278 4630 22330
rect 10722 22278 10774 22330
rect 10786 22278 10838 22330
rect 10850 22278 10902 22330
rect 10914 22278 10966 22330
rect 10978 22278 11030 22330
rect 1860 22176 1912 22228
rect 2320 22219 2372 22228
rect 2320 22185 2329 22219
rect 2329 22185 2363 22219
rect 2363 22185 2372 22219
rect 2320 22176 2372 22185
rect 2964 22176 3016 22228
rect 3332 22176 3384 22228
rect 3700 22176 3752 22228
rect 4436 22219 4488 22228
rect 4436 22185 4445 22219
rect 4445 22185 4479 22219
rect 4479 22185 4488 22219
rect 4436 22176 4488 22185
rect 4712 22176 4764 22228
rect 5172 22219 5224 22228
rect 5172 22185 5181 22219
rect 5181 22185 5215 22219
rect 5215 22185 5224 22219
rect 5172 22176 5224 22185
rect 4160 22108 4212 22160
rect 1768 22083 1820 22092
rect 1768 22049 1777 22083
rect 1777 22049 1811 22083
rect 1811 22049 1820 22083
rect 1768 22040 1820 22049
rect 1860 22040 1912 22092
rect 756 21972 808 22024
rect 2320 21972 2372 22024
rect 2688 22083 2740 22092
rect 2688 22049 2697 22083
rect 2697 22049 2731 22083
rect 2731 22049 2740 22083
rect 2688 22040 2740 22049
rect 2964 22040 3016 22092
rect 3332 22040 3384 22092
rect 3424 21904 3476 21956
rect 3700 22083 3752 22092
rect 3700 22049 3709 22083
rect 3709 22049 3743 22083
rect 3743 22049 3752 22083
rect 3700 22040 3752 22049
rect 3792 22083 3844 22092
rect 3792 22049 3801 22083
rect 3801 22049 3835 22083
rect 3835 22049 3844 22083
rect 3792 22040 3844 22049
rect 3884 22083 3936 22092
rect 3884 22049 3893 22083
rect 3893 22049 3927 22083
rect 3927 22049 3936 22083
rect 3884 22040 3936 22049
rect 4068 22040 4120 22092
rect 4252 22083 4304 22092
rect 4252 22049 4261 22083
rect 4261 22049 4295 22083
rect 4295 22049 4304 22083
rect 4252 22040 4304 22049
rect 5448 22108 5500 22160
rect 5816 22176 5868 22228
rect 6184 22176 6236 22228
rect 4344 21972 4396 22024
rect 4712 21972 4764 22024
rect 5264 22083 5316 22092
rect 5264 22049 5273 22083
rect 5273 22049 5307 22083
rect 5307 22049 5316 22083
rect 5264 22040 5316 22049
rect 5448 22015 5500 22024
rect 5448 21981 5457 22015
rect 5457 21981 5491 22015
rect 5491 21981 5500 22015
rect 5448 21972 5500 21981
rect 6276 22108 6328 22160
rect 6644 22176 6696 22228
rect 7932 22176 7984 22228
rect 8116 22219 8168 22228
rect 8116 22185 8125 22219
rect 8125 22185 8159 22219
rect 8159 22185 8168 22219
rect 8116 22176 8168 22185
rect 6920 22108 6972 22160
rect 7012 22108 7064 22160
rect 5724 22040 5776 22092
rect 6644 22040 6696 22092
rect 6736 22040 6788 22092
rect 7748 22040 7800 22092
rect 8392 22151 8444 22160
rect 8392 22117 8401 22151
rect 8401 22117 8435 22151
rect 8435 22117 8444 22151
rect 8392 22108 8444 22117
rect 8576 22108 8628 22160
rect 8852 22108 8904 22160
rect 5908 21972 5960 22024
rect 7840 21972 7892 22024
rect 8208 21972 8260 22024
rect 10416 22219 10468 22228
rect 10416 22185 10425 22219
rect 10425 22185 10459 22219
rect 10459 22185 10468 22219
rect 10416 22176 10468 22185
rect 9220 22040 9272 22092
rect 9680 22083 9732 22092
rect 9680 22049 9689 22083
rect 9689 22049 9723 22083
rect 9723 22049 9732 22083
rect 9680 22040 9732 22049
rect 10324 22108 10376 22160
rect 10692 22108 10744 22160
rect 10048 22040 10100 22092
rect 10416 22083 10468 22092
rect 10416 22049 10425 22083
rect 10425 22049 10459 22083
rect 10459 22049 10468 22083
rect 10416 22040 10468 22049
rect 2872 21836 2924 21888
rect 3332 21879 3384 21888
rect 3332 21845 3341 21879
rect 3341 21845 3375 21879
rect 3375 21845 3384 21879
rect 3332 21836 3384 21845
rect 4252 21836 4304 21888
rect 6276 21947 6328 21956
rect 6276 21913 6285 21947
rect 6285 21913 6319 21947
rect 6319 21913 6328 21947
rect 6276 21904 6328 21913
rect 7288 21904 7340 21956
rect 8576 21972 8628 22024
rect 8760 21972 8812 22024
rect 9404 22015 9456 22024
rect 9404 21981 9413 22015
rect 9413 21981 9447 22015
rect 9447 21981 9456 22015
rect 9404 21972 9456 21981
rect 10600 21904 10652 21956
rect 6920 21836 6972 21888
rect 7932 21836 7984 21888
rect 9588 21836 9640 21888
rect 9680 21836 9732 21888
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 10062 21734 10114 21786
rect 10126 21734 10178 21786
rect 10190 21734 10242 21786
rect 10254 21734 10306 21786
rect 10318 21734 10370 21786
rect 1032 21675 1084 21684
rect 1032 21641 1041 21675
rect 1041 21641 1075 21675
rect 1075 21641 1084 21675
rect 1032 21632 1084 21641
rect 1676 21632 1728 21684
rect 3148 21632 3200 21684
rect 3424 21632 3476 21684
rect 4344 21632 4396 21684
rect 2228 21564 2280 21616
rect 2596 21564 2648 21616
rect 3792 21564 3844 21616
rect 3976 21564 4028 21616
rect 4436 21564 4488 21616
rect 5172 21632 5224 21684
rect 1308 21428 1360 21480
rect 1584 21428 1636 21480
rect 2044 21496 2096 21548
rect 2412 21496 2464 21548
rect 2872 21428 2924 21480
rect 3148 21428 3200 21480
rect 3332 21428 3384 21480
rect 4988 21496 5040 21548
rect 5172 21496 5224 21548
rect 5448 21539 5500 21548
rect 5448 21505 5457 21539
rect 5457 21505 5491 21539
rect 5491 21505 5500 21539
rect 5448 21496 5500 21505
rect 5908 21564 5960 21616
rect 6552 21632 6604 21684
rect 7472 21632 7524 21684
rect 3608 21471 3660 21480
rect 3608 21437 3617 21471
rect 3617 21437 3651 21471
rect 3651 21437 3660 21471
rect 3608 21428 3660 21437
rect 3976 21428 4028 21480
rect 4344 21428 4396 21480
rect 4804 21428 4856 21480
rect 5632 21428 5684 21480
rect 5724 21428 5776 21480
rect 6000 21471 6052 21480
rect 6000 21437 6009 21471
rect 6009 21437 6043 21471
rect 6043 21437 6052 21471
rect 6000 21428 6052 21437
rect 6184 21428 6236 21480
rect 6276 21471 6328 21480
rect 6276 21437 6285 21471
rect 6285 21437 6319 21471
rect 6319 21437 6328 21471
rect 6276 21428 6328 21437
rect 2504 21360 2556 21412
rect 2688 21360 2740 21412
rect 3884 21360 3936 21412
rect 4068 21360 4120 21412
rect 5816 21360 5868 21412
rect 7104 21564 7156 21616
rect 7288 21564 7340 21616
rect 6736 21539 6788 21548
rect 6736 21505 6745 21539
rect 6745 21505 6779 21539
rect 6779 21505 6788 21539
rect 6736 21496 6788 21505
rect 7932 21564 7984 21616
rect 8576 21632 8628 21684
rect 8944 21632 8996 21684
rect 9220 21632 9272 21684
rect 10416 21632 10468 21684
rect 7748 21496 7800 21548
rect 8668 21496 8720 21548
rect 8944 21496 8996 21548
rect 9312 21496 9364 21548
rect 6644 21471 6696 21480
rect 6644 21437 6653 21471
rect 6653 21437 6687 21471
rect 6687 21437 6696 21471
rect 6644 21428 6696 21437
rect 7196 21428 7248 21480
rect 7932 21428 7984 21480
rect 8392 21471 8444 21480
rect 8392 21437 8401 21471
rect 8401 21437 8435 21471
rect 8435 21437 8444 21471
rect 8392 21428 8444 21437
rect 8484 21428 8536 21480
rect 9588 21428 9640 21480
rect 7012 21360 7064 21412
rect 7564 21360 7616 21412
rect 8760 21360 8812 21412
rect 8944 21360 8996 21412
rect 9956 21471 10008 21480
rect 9956 21437 9965 21471
rect 9965 21437 9999 21471
rect 9999 21437 10008 21471
rect 9956 21428 10008 21437
rect 10140 21360 10192 21412
rect 10692 21360 10744 21412
rect 1400 21292 1452 21344
rect 2228 21292 2280 21344
rect 2320 21292 2372 21344
rect 3056 21292 3108 21344
rect 3700 21292 3752 21344
rect 7656 21292 7708 21344
rect 7840 21335 7892 21344
rect 7840 21301 7849 21335
rect 7849 21301 7883 21335
rect 7883 21301 7892 21335
rect 7840 21292 7892 21301
rect 8576 21335 8628 21344
rect 8576 21301 8585 21335
rect 8585 21301 8619 21335
rect 8619 21301 8628 21335
rect 8576 21292 8628 21301
rect 9588 21292 9640 21344
rect 11244 21292 11296 21344
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 10722 21190 10774 21242
rect 10786 21190 10838 21242
rect 10850 21190 10902 21242
rect 10914 21190 10966 21242
rect 10978 21190 11030 21242
rect 1308 21131 1360 21140
rect 1308 21097 1317 21131
rect 1317 21097 1351 21131
rect 1351 21097 1360 21131
rect 1308 21088 1360 21097
rect 1860 21131 1912 21140
rect 1860 21097 1869 21131
rect 1869 21097 1903 21131
rect 1903 21097 1912 21131
rect 1860 21088 1912 21097
rect 2136 21088 2188 21140
rect 2504 21088 2556 21140
rect 1400 20952 1452 21004
rect 1676 20995 1728 21004
rect 1676 20961 1685 20995
rect 1685 20961 1719 20995
rect 1719 20961 1728 20995
rect 1676 20952 1728 20961
rect 3240 21020 3292 21072
rect 3332 21063 3384 21072
rect 3332 21029 3341 21063
rect 3341 21029 3375 21063
rect 3375 21029 3384 21063
rect 3332 21020 3384 21029
rect 3792 21020 3844 21072
rect 2044 20995 2096 21004
rect 2044 20961 2053 20995
rect 2053 20961 2087 20995
rect 2087 20961 2096 20995
rect 2044 20952 2096 20961
rect 2320 20995 2372 21004
rect 2320 20961 2329 20995
rect 2329 20961 2363 20995
rect 2363 20961 2372 20995
rect 2320 20952 2372 20961
rect 2504 20952 2556 21004
rect 2688 20952 2740 21004
rect 3148 20995 3200 21004
rect 3148 20961 3157 20995
rect 3157 20961 3191 20995
rect 3191 20961 3200 20995
rect 3148 20952 3200 20961
rect 3424 20952 3476 21004
rect 3608 20995 3660 21004
rect 3608 20961 3617 20995
rect 3617 20961 3651 20995
rect 3651 20961 3660 20995
rect 3608 20952 3660 20961
rect 3700 20995 3752 21004
rect 3700 20961 3709 20995
rect 3709 20961 3743 20995
rect 3743 20961 3752 20995
rect 3700 20952 3752 20961
rect 3884 20995 3936 21004
rect 3884 20961 3893 20995
rect 3893 20961 3927 20995
rect 3927 20961 3936 20995
rect 3884 20952 3936 20961
rect 4068 20995 4120 21004
rect 4068 20961 4077 20995
rect 4077 20961 4111 20995
rect 4111 20961 4120 20995
rect 4068 20952 4120 20961
rect 4712 21088 4764 21140
rect 4804 21063 4856 21072
rect 4804 21029 4813 21063
rect 4813 21029 4847 21063
rect 4847 21029 4856 21063
rect 4804 21020 4856 21029
rect 5540 21020 5592 21072
rect 4896 20952 4948 21004
rect 5448 20952 5500 21004
rect 6368 21020 6420 21072
rect 7012 21088 7064 21140
rect 7748 21088 7800 21140
rect 9864 21088 9916 21140
rect 10508 21088 10560 21140
rect 11244 21088 11296 21140
rect 5724 20952 5776 21004
rect 6000 20995 6052 21004
rect 6000 20961 6009 20995
rect 6009 20961 6043 20995
rect 6043 20961 6052 20995
rect 6000 20952 6052 20961
rect 6736 21020 6788 21072
rect 2964 20927 3016 20936
rect 2964 20893 2973 20927
rect 2973 20893 3007 20927
rect 3007 20893 3016 20927
rect 2964 20884 3016 20893
rect 4252 20884 4304 20936
rect 5356 20927 5408 20936
rect 5356 20893 5365 20927
rect 5365 20893 5399 20927
rect 5399 20893 5408 20927
rect 5356 20884 5408 20893
rect 1584 20748 1636 20800
rect 3148 20816 3200 20868
rect 3332 20816 3384 20868
rect 5448 20859 5500 20868
rect 5448 20825 5457 20859
rect 5457 20825 5491 20859
rect 5491 20825 5500 20859
rect 5448 20816 5500 20825
rect 6736 20816 6788 20868
rect 4712 20748 4764 20800
rect 6920 20884 6972 20936
rect 7288 20995 7340 21004
rect 7288 20961 7297 20995
rect 7297 20961 7331 20995
rect 7331 20961 7340 20995
rect 7288 20952 7340 20961
rect 7472 20995 7524 21004
rect 7472 20961 7481 20995
rect 7481 20961 7515 20995
rect 7515 20961 7524 20995
rect 7472 20952 7524 20961
rect 8576 21020 8628 21072
rect 9128 21020 9180 21072
rect 7840 20995 7892 21004
rect 7840 20961 7849 20995
rect 7849 20961 7883 20995
rect 7883 20961 7892 20995
rect 7840 20952 7892 20961
rect 7196 20884 7248 20936
rect 8024 20884 8076 20936
rect 8852 20927 8904 20936
rect 8852 20893 8861 20927
rect 8861 20893 8895 20927
rect 8895 20893 8904 20927
rect 8852 20884 8904 20893
rect 9128 20884 9180 20936
rect 8392 20816 8444 20868
rect 9404 20952 9456 21004
rect 10048 20884 10100 20936
rect 7104 20748 7156 20800
rect 9864 20816 9916 20868
rect 9680 20748 9732 20800
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 10062 20646 10114 20698
rect 10126 20646 10178 20698
rect 10190 20646 10242 20698
rect 10254 20646 10306 20698
rect 10318 20646 10370 20698
rect 2596 20544 2648 20596
rect 3516 20544 3568 20596
rect 6000 20544 6052 20596
rect 6552 20544 6604 20596
rect 6920 20544 6972 20596
rect 7656 20587 7708 20596
rect 7656 20553 7665 20587
rect 7665 20553 7699 20587
rect 7699 20553 7708 20587
rect 7656 20544 7708 20553
rect 9404 20587 9456 20596
rect 9404 20553 9413 20587
rect 9413 20553 9447 20587
rect 9447 20553 9456 20587
rect 9404 20544 9456 20553
rect 1676 20476 1728 20528
rect 3424 20476 3476 20528
rect 4252 20476 4304 20528
rect 5724 20476 5776 20528
rect 1400 20408 1452 20460
rect 1584 20408 1636 20460
rect 2044 20383 2096 20392
rect 2044 20349 2053 20383
rect 2053 20349 2087 20383
rect 2087 20349 2096 20383
rect 2044 20340 2096 20349
rect 2228 20383 2280 20392
rect 2228 20349 2237 20383
rect 2237 20349 2271 20383
rect 2271 20349 2280 20383
rect 2228 20340 2280 20349
rect 2504 20383 2556 20392
rect 2504 20349 2513 20383
rect 2513 20349 2547 20383
rect 2547 20349 2556 20383
rect 2504 20340 2556 20349
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 1216 20272 1268 20324
rect 3700 20383 3752 20392
rect 3700 20349 3709 20383
rect 3709 20349 3743 20383
rect 3743 20349 3752 20383
rect 3700 20340 3752 20349
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 4252 20340 4304 20392
rect 3332 20272 3384 20324
rect 3976 20272 4028 20324
rect 4804 20340 4856 20392
rect 4988 20383 5040 20392
rect 4988 20349 4997 20383
rect 4997 20349 5031 20383
rect 5031 20349 5040 20383
rect 4988 20340 5040 20349
rect 5172 20383 5224 20392
rect 5172 20349 5181 20383
rect 5181 20349 5215 20383
rect 5215 20349 5224 20383
rect 5172 20340 5224 20349
rect 5816 20340 5868 20392
rect 1768 20204 1820 20256
rect 3516 20204 3568 20256
rect 5724 20204 5776 20256
rect 5816 20247 5868 20256
rect 5816 20213 5825 20247
rect 5825 20213 5859 20247
rect 5859 20213 5868 20247
rect 5816 20204 5868 20213
rect 6552 20408 6604 20460
rect 7104 20408 7156 20460
rect 6092 20272 6144 20324
rect 6828 20204 6880 20256
rect 8484 20383 8536 20392
rect 8484 20349 8493 20383
rect 8493 20349 8527 20383
rect 8527 20349 8536 20383
rect 8484 20340 8536 20349
rect 8576 20340 8628 20392
rect 9496 20408 9548 20460
rect 10508 20408 10560 20460
rect 9772 20383 9824 20392
rect 9772 20349 9781 20383
rect 9781 20349 9815 20383
rect 9815 20349 9824 20383
rect 9772 20340 9824 20349
rect 7288 20204 7340 20256
rect 8024 20272 8076 20324
rect 11336 20340 11388 20392
rect 7472 20204 7524 20256
rect 9772 20204 9824 20256
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 10722 20102 10774 20154
rect 10786 20102 10838 20154
rect 10850 20102 10902 20154
rect 10914 20102 10966 20154
rect 10978 20102 11030 20154
rect 1952 20000 2004 20052
rect 3240 20000 3292 20052
rect 3332 20000 3384 20052
rect 3700 20000 3752 20052
rect 1676 19932 1728 19984
rect 2504 19932 2556 19984
rect 2872 19932 2924 19984
rect 1584 19864 1636 19916
rect 2320 19864 2372 19916
rect 2596 19864 2648 19916
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 3148 19864 3200 19916
rect 3976 19932 4028 19984
rect 4528 20000 4580 20052
rect 4804 20043 4856 20052
rect 4804 20009 4813 20043
rect 4813 20009 4847 20043
rect 4847 20009 4856 20043
rect 4804 20000 4856 20009
rect 5172 20000 5224 20052
rect 5632 20000 5684 20052
rect 1216 19839 1268 19848
rect 1216 19805 1225 19839
rect 1225 19805 1259 19839
rect 1259 19805 1268 19839
rect 1216 19796 1268 19805
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 3240 19796 3292 19848
rect 2412 19728 2464 19780
rect 1032 19660 1084 19712
rect 2688 19660 2740 19712
rect 4160 19907 4212 19916
rect 4160 19873 4169 19907
rect 4169 19873 4203 19907
rect 4203 19873 4212 19907
rect 4160 19864 4212 19873
rect 4436 19907 4488 19916
rect 4436 19873 4445 19907
rect 4445 19873 4479 19907
rect 4479 19873 4488 19907
rect 4436 19864 4488 19873
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 4252 19728 4304 19780
rect 6092 19932 6144 19984
rect 6552 19975 6604 19984
rect 6552 19941 6561 19975
rect 6561 19941 6595 19975
rect 6595 19941 6604 19975
rect 6552 19932 6604 19941
rect 5908 19864 5960 19916
rect 5448 19839 5500 19848
rect 5448 19805 5457 19839
rect 5457 19805 5491 19839
rect 5491 19805 5500 19839
rect 5448 19796 5500 19805
rect 4896 19728 4948 19780
rect 6184 19839 6236 19848
rect 6184 19805 6193 19839
rect 6193 19805 6227 19839
rect 6227 19805 6236 19839
rect 6184 19796 6236 19805
rect 6828 19864 6880 19916
rect 7104 19907 7156 19916
rect 7104 19873 7113 19907
rect 7113 19873 7147 19907
rect 7147 19873 7156 19907
rect 7104 19864 7156 19873
rect 7196 19864 7248 19916
rect 7932 19932 7984 19984
rect 8300 19864 8352 19916
rect 8668 19932 8720 19984
rect 9772 19932 9824 19984
rect 9036 19864 9088 19916
rect 9128 19907 9180 19916
rect 9128 19873 9137 19907
rect 9137 19873 9171 19907
rect 9171 19873 9180 19907
rect 9128 19864 9180 19873
rect 6920 19839 6972 19848
rect 6920 19805 6929 19839
rect 6929 19805 6963 19839
rect 6963 19805 6972 19839
rect 6920 19796 6972 19805
rect 7012 19839 7064 19848
rect 7012 19805 7021 19839
rect 7021 19805 7055 19839
rect 7055 19805 7064 19839
rect 7012 19796 7064 19805
rect 7472 19796 7524 19848
rect 7748 19796 7800 19848
rect 6828 19728 6880 19780
rect 7288 19660 7340 19712
rect 7472 19660 7524 19712
rect 7932 19660 7984 19712
rect 8392 19728 8444 19780
rect 9496 19728 9548 19780
rect 8852 19660 8904 19712
rect 10416 19660 10468 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 10062 19558 10114 19610
rect 10126 19558 10178 19610
rect 10190 19558 10242 19610
rect 10254 19558 10306 19610
rect 10318 19558 10370 19610
rect 2044 19456 2096 19508
rect 2780 19456 2832 19508
rect 3056 19456 3108 19508
rect 3516 19456 3568 19508
rect 4068 19456 4120 19508
rect 4436 19456 4488 19508
rect 204 19388 256 19440
rect 572 19388 624 19440
rect 1124 19388 1176 19440
rect 572 19252 624 19304
rect 1492 19320 1544 19372
rect 1124 19295 1176 19304
rect 1124 19261 1133 19295
rect 1133 19261 1167 19295
rect 1167 19261 1176 19295
rect 1124 19252 1176 19261
rect 1308 19252 1360 19304
rect 848 19227 900 19236
rect 848 19193 857 19227
rect 857 19193 891 19227
rect 891 19193 900 19227
rect 848 19184 900 19193
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 2688 19388 2740 19440
rect 3700 19388 3752 19440
rect 4528 19388 4580 19440
rect 2596 19320 2648 19372
rect 3240 19363 3292 19372
rect 3240 19329 3249 19363
rect 3249 19329 3283 19363
rect 3283 19329 3292 19363
rect 3240 19320 3292 19329
rect 3332 19320 3384 19372
rect 2504 19295 2556 19304
rect 2504 19261 2513 19295
rect 2513 19261 2547 19295
rect 2547 19261 2556 19295
rect 2504 19252 2556 19261
rect 3424 19295 3476 19304
rect 3424 19261 3433 19295
rect 3433 19261 3467 19295
rect 3467 19261 3476 19295
rect 3424 19252 3476 19261
rect 3700 19252 3752 19304
rect 4712 19320 4764 19372
rect 5816 19456 5868 19508
rect 6000 19456 6052 19508
rect 7288 19456 7340 19508
rect 7932 19456 7984 19508
rect 8576 19456 8628 19508
rect 8668 19499 8720 19508
rect 8668 19465 8677 19499
rect 8677 19465 8711 19499
rect 8711 19465 8720 19499
rect 8668 19456 8720 19465
rect 9680 19456 9732 19508
rect 3976 19252 4028 19304
rect 3056 19116 3108 19168
rect 3332 19116 3384 19168
rect 3516 19116 3568 19168
rect 4528 19227 4580 19236
rect 4528 19193 4537 19227
rect 4537 19193 4571 19227
rect 4571 19193 4580 19227
rect 4528 19184 4580 19193
rect 4988 19295 5040 19304
rect 4988 19261 4997 19295
rect 4997 19261 5031 19295
rect 5031 19261 5040 19295
rect 4988 19252 5040 19261
rect 5540 19320 5592 19372
rect 7380 19388 7432 19440
rect 9128 19388 9180 19440
rect 5632 19295 5684 19304
rect 5632 19261 5641 19295
rect 5641 19261 5675 19295
rect 5675 19261 5684 19295
rect 5632 19252 5684 19261
rect 5080 19116 5132 19168
rect 5448 19159 5500 19168
rect 5448 19125 5457 19159
rect 5457 19125 5491 19159
rect 5491 19125 5500 19159
rect 5448 19116 5500 19125
rect 6000 19295 6052 19304
rect 6000 19261 6009 19295
rect 6009 19261 6043 19295
rect 6043 19261 6052 19295
rect 6000 19252 6052 19261
rect 7748 19320 7800 19372
rect 8576 19320 8628 19372
rect 6460 19295 6512 19304
rect 6460 19261 6469 19295
rect 6469 19261 6503 19295
rect 6503 19261 6512 19295
rect 6460 19252 6512 19261
rect 6276 19184 6328 19236
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 6920 19295 6972 19304
rect 6920 19261 6929 19295
rect 6929 19261 6963 19295
rect 6963 19261 6972 19295
rect 6920 19252 6972 19261
rect 7104 19295 7156 19304
rect 7104 19261 7113 19295
rect 7113 19261 7147 19295
rect 7147 19261 7156 19295
rect 7104 19252 7156 19261
rect 7288 19295 7340 19304
rect 7288 19261 7297 19295
rect 7297 19261 7331 19295
rect 7331 19261 7340 19295
rect 7288 19252 7340 19261
rect 8116 19252 8168 19304
rect 8852 19295 8904 19304
rect 8852 19261 8861 19295
rect 8861 19261 8895 19295
rect 8895 19261 8904 19295
rect 8852 19252 8904 19261
rect 8484 19184 8536 19236
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 9312 19252 9364 19304
rect 9772 19295 9824 19304
rect 9772 19261 9781 19295
rect 9781 19261 9815 19295
rect 9815 19261 9824 19295
rect 9772 19252 9824 19261
rect 10416 19320 10468 19372
rect 7932 19116 7984 19168
rect 8852 19116 8904 19168
rect 9036 19116 9088 19168
rect 9404 19116 9456 19168
rect 9772 19116 9824 19168
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 10722 19014 10774 19066
rect 10786 19014 10838 19066
rect 10850 19014 10902 19066
rect 10914 19014 10966 19066
rect 10978 19014 11030 19066
rect 940 18912 992 18964
rect 1492 18912 1544 18964
rect 2136 18912 2188 18964
rect 4068 18955 4120 18964
rect 4068 18921 4077 18955
rect 4077 18921 4111 18955
rect 4111 18921 4120 18955
rect 4068 18912 4120 18921
rect 4344 18912 4396 18964
rect 5264 18912 5316 18964
rect 5448 18912 5500 18964
rect 6276 18912 6328 18964
rect 6920 18955 6972 18964
rect 6920 18921 6929 18955
rect 6929 18921 6963 18955
rect 6963 18921 6972 18955
rect 6920 18912 6972 18921
rect 572 18844 624 18896
rect 2872 18844 2924 18896
rect 1400 18776 1452 18828
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 2044 18819 2096 18828
rect 2044 18785 2053 18819
rect 2053 18785 2087 18819
rect 2087 18785 2096 18819
rect 2044 18776 2096 18785
rect 2320 18819 2372 18828
rect 2320 18785 2329 18819
rect 2329 18785 2363 18819
rect 2363 18785 2372 18819
rect 2320 18776 2372 18785
rect 2504 18819 2556 18828
rect 2504 18785 2513 18819
rect 2513 18785 2547 18819
rect 2547 18785 2556 18819
rect 2504 18776 2556 18785
rect 2688 18819 2740 18828
rect 2688 18785 2697 18819
rect 2697 18785 2731 18819
rect 2731 18785 2740 18819
rect 2688 18776 2740 18785
rect 3056 18819 3108 18828
rect 3056 18785 3065 18819
rect 3065 18785 3099 18819
rect 3099 18785 3108 18819
rect 3056 18776 3108 18785
rect 2136 18708 2188 18760
rect 2228 18751 2280 18760
rect 2228 18717 2237 18751
rect 2237 18717 2271 18751
rect 2271 18717 2280 18751
rect 2228 18708 2280 18717
rect 2596 18708 2648 18760
rect 1584 18640 1636 18692
rect 3516 18776 3568 18828
rect 3884 18819 3936 18828
rect 3884 18785 3893 18819
rect 3893 18785 3927 18819
rect 3927 18785 3936 18819
rect 3884 18776 3936 18785
rect 4344 18819 4396 18828
rect 4344 18785 4353 18819
rect 4353 18785 4387 18819
rect 4387 18785 4396 18819
rect 4344 18776 4396 18785
rect 848 18615 900 18624
rect 848 18581 857 18615
rect 857 18581 891 18615
rect 891 18581 900 18615
rect 848 18572 900 18581
rect 2320 18572 2372 18624
rect 3424 18640 3476 18692
rect 4252 18708 4304 18760
rect 5080 18776 5132 18828
rect 5724 18844 5776 18896
rect 6000 18844 6052 18896
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 5908 18751 5960 18760
rect 5908 18717 5917 18751
rect 5917 18717 5951 18751
rect 5951 18717 5960 18751
rect 5908 18708 5960 18717
rect 6368 18776 6420 18828
rect 6552 18776 6604 18828
rect 7196 18844 7248 18896
rect 7288 18887 7340 18896
rect 7288 18853 7297 18887
rect 7297 18853 7331 18887
rect 7331 18853 7340 18887
rect 7288 18844 7340 18853
rect 6920 18708 6972 18760
rect 7564 18776 7616 18828
rect 7748 18776 7800 18828
rect 10416 18912 10468 18964
rect 9588 18844 9640 18896
rect 11244 18844 11296 18896
rect 8116 18708 8168 18760
rect 2872 18615 2924 18624
rect 2872 18581 2881 18615
rect 2881 18581 2915 18615
rect 2915 18581 2924 18615
rect 2872 18572 2924 18581
rect 3056 18572 3108 18624
rect 3608 18572 3660 18624
rect 3976 18572 4028 18624
rect 4160 18572 4212 18624
rect 4620 18640 4672 18692
rect 4712 18683 4764 18692
rect 4712 18649 4721 18683
rect 4721 18649 4755 18683
rect 4755 18649 4764 18683
rect 4712 18640 4764 18649
rect 5080 18640 5132 18692
rect 6368 18640 6420 18692
rect 6552 18640 6604 18692
rect 7288 18640 7340 18692
rect 8668 18776 8720 18828
rect 9036 18751 9088 18760
rect 9036 18717 9045 18751
rect 9045 18717 9079 18751
rect 9079 18717 9088 18751
rect 9036 18708 9088 18717
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 10508 18776 10560 18828
rect 9496 18640 9548 18692
rect 9680 18683 9732 18692
rect 9680 18649 9689 18683
rect 9689 18649 9723 18683
rect 9723 18649 9732 18683
rect 9680 18640 9732 18649
rect 6000 18615 6052 18624
rect 6000 18581 6009 18615
rect 6009 18581 6043 18615
rect 6043 18581 6052 18615
rect 6000 18572 6052 18581
rect 6092 18572 6144 18624
rect 6736 18572 6788 18624
rect 7104 18572 7156 18624
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 10062 18470 10114 18522
rect 10126 18470 10178 18522
rect 10190 18470 10242 18522
rect 10254 18470 10306 18522
rect 10318 18470 10370 18522
rect 2044 18411 2096 18420
rect 2044 18377 2053 18411
rect 2053 18377 2087 18411
rect 2087 18377 2096 18411
rect 2044 18368 2096 18377
rect 5172 18368 5224 18420
rect 5356 18368 5408 18420
rect 5540 18411 5592 18420
rect 5540 18377 5549 18411
rect 5549 18377 5583 18411
rect 5583 18377 5592 18411
rect 5540 18368 5592 18377
rect 5724 18368 5776 18420
rect 3424 18300 3476 18352
rect 1124 18232 1176 18284
rect 2320 18275 2372 18284
rect 2320 18241 2329 18275
rect 2329 18241 2363 18275
rect 2363 18241 2372 18275
rect 2320 18232 2372 18241
rect 1584 18207 1636 18216
rect 1584 18173 1593 18207
rect 1593 18173 1627 18207
rect 1627 18173 1636 18207
rect 1584 18164 1636 18173
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 1400 18096 1452 18148
rect 2872 18164 2924 18216
rect 3240 18207 3292 18216
rect 3240 18173 3249 18207
rect 3249 18173 3283 18207
rect 3283 18173 3292 18207
rect 3240 18164 3292 18173
rect 3332 18207 3384 18216
rect 3332 18173 3341 18207
rect 3341 18173 3375 18207
rect 3375 18173 3384 18207
rect 3332 18164 3384 18173
rect 3976 18300 4028 18352
rect 4160 18232 4212 18284
rect 4344 18275 4396 18284
rect 4344 18241 4353 18275
rect 4353 18241 4387 18275
rect 4387 18241 4396 18275
rect 4344 18232 4396 18241
rect 4528 18232 4580 18284
rect 2964 18096 3016 18148
rect 3976 18164 4028 18216
rect 3792 18096 3844 18148
rect 1952 18028 2004 18080
rect 3700 18028 3752 18080
rect 5080 18164 5132 18216
rect 5172 18164 5224 18216
rect 4620 18096 4672 18148
rect 4436 18028 4488 18080
rect 5080 18071 5132 18080
rect 5080 18037 5089 18071
rect 5089 18037 5123 18071
rect 5123 18037 5132 18071
rect 5080 18028 5132 18037
rect 6000 18300 6052 18352
rect 5724 18275 5776 18284
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 5724 18232 5776 18241
rect 5816 18232 5868 18284
rect 6552 18368 6604 18420
rect 6828 18300 6880 18352
rect 7564 18300 7616 18352
rect 7656 18300 7708 18352
rect 6552 18232 6604 18284
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 6368 18096 6420 18148
rect 7288 18207 7340 18216
rect 7288 18173 7297 18207
rect 7297 18173 7331 18207
rect 7331 18173 7340 18207
rect 7288 18164 7340 18173
rect 6552 18096 6604 18148
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 7012 18028 7064 18080
rect 7288 18028 7340 18080
rect 7656 18207 7708 18216
rect 7656 18173 7665 18207
rect 7665 18173 7699 18207
rect 7699 18173 7708 18207
rect 7656 18164 7708 18173
rect 9036 18343 9088 18352
rect 9036 18309 9045 18343
rect 9045 18309 9079 18343
rect 9079 18309 9088 18343
rect 9036 18300 9088 18309
rect 8024 18232 8076 18284
rect 8668 18275 8720 18284
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 8668 18232 8720 18241
rect 8392 18164 8444 18216
rect 9588 18300 9640 18352
rect 9404 18232 9456 18284
rect 10508 18232 10560 18284
rect 8484 18096 8536 18148
rect 9680 18164 9732 18216
rect 9220 18028 9272 18080
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 10722 17926 10774 17978
rect 10786 17926 10838 17978
rect 10850 17926 10902 17978
rect 10914 17926 10966 17978
rect 10978 17926 11030 17978
rect 1676 17824 1728 17876
rect 4068 17824 4120 17876
rect 4344 17824 4396 17876
rect 5080 17824 5132 17876
rect 5908 17824 5960 17876
rect 6736 17824 6788 17876
rect 848 17756 900 17808
rect 1308 17731 1360 17740
rect 1308 17697 1317 17731
rect 1317 17697 1351 17731
rect 1351 17697 1360 17731
rect 1308 17688 1360 17697
rect 388 17620 440 17672
rect 848 17620 900 17672
rect 1124 17527 1176 17536
rect 1124 17493 1133 17527
rect 1133 17493 1167 17527
rect 1167 17493 1176 17527
rect 1124 17484 1176 17493
rect 2136 17731 2188 17740
rect 2136 17697 2145 17731
rect 2145 17697 2179 17731
rect 2179 17697 2188 17731
rect 2136 17688 2188 17697
rect 2228 17620 2280 17672
rect 2504 17620 2556 17672
rect 2780 17688 2832 17740
rect 3516 17731 3568 17740
rect 3516 17697 3525 17731
rect 3525 17697 3559 17731
rect 3559 17697 3568 17731
rect 3516 17688 3568 17697
rect 4528 17756 4580 17808
rect 3884 17731 3936 17740
rect 3884 17697 3893 17731
rect 3893 17697 3927 17731
rect 3927 17697 3936 17731
rect 3884 17688 3936 17697
rect 4252 17688 4304 17740
rect 4620 17731 4672 17740
rect 4068 17663 4120 17672
rect 4068 17629 4077 17663
rect 4077 17629 4111 17663
rect 4111 17629 4120 17663
rect 4068 17620 4120 17629
rect 1860 17552 1912 17604
rect 2688 17552 2740 17604
rect 2872 17552 2924 17604
rect 3056 17552 3108 17604
rect 3516 17552 3568 17604
rect 4436 17552 4488 17604
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 4804 17731 4856 17740
rect 4804 17697 4813 17731
rect 4813 17697 4847 17731
rect 4847 17697 4856 17731
rect 4804 17688 4856 17697
rect 5080 17731 5132 17740
rect 5080 17697 5089 17731
rect 5089 17697 5123 17731
rect 5123 17697 5132 17731
rect 5080 17688 5132 17697
rect 5264 17731 5316 17740
rect 5264 17697 5273 17731
rect 5273 17697 5307 17731
rect 5307 17697 5316 17731
rect 5264 17688 5316 17697
rect 5448 17688 5500 17740
rect 5632 17731 5684 17740
rect 5632 17697 5641 17731
rect 5641 17697 5675 17731
rect 5675 17697 5684 17731
rect 5632 17688 5684 17697
rect 5908 17688 5960 17740
rect 6552 17756 6604 17808
rect 6276 17688 6328 17740
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 6460 17729 6512 17740
rect 6460 17695 6469 17729
rect 6469 17695 6503 17729
rect 6503 17695 6512 17729
rect 6460 17688 6512 17695
rect 7380 17756 7432 17808
rect 7748 17824 7800 17876
rect 6552 17620 6604 17672
rect 7196 17731 7248 17740
rect 7196 17697 7205 17731
rect 7205 17697 7239 17731
rect 7239 17697 7248 17731
rect 7196 17688 7248 17697
rect 6828 17663 6880 17672
rect 6828 17629 6837 17663
rect 6837 17629 6871 17663
rect 6871 17629 6880 17663
rect 6828 17620 6880 17629
rect 1584 17484 1636 17536
rect 2044 17484 2096 17536
rect 2504 17484 2556 17536
rect 3424 17484 3476 17536
rect 3700 17484 3752 17536
rect 4804 17484 4856 17536
rect 6276 17595 6328 17604
rect 6276 17561 6285 17595
rect 6285 17561 6319 17595
rect 6319 17561 6328 17595
rect 6276 17552 6328 17561
rect 6828 17484 6880 17536
rect 7288 17552 7340 17604
rect 7656 17731 7708 17740
rect 7656 17697 7665 17731
rect 7665 17697 7699 17731
rect 7699 17697 7708 17731
rect 7656 17688 7708 17697
rect 8024 17688 8076 17740
rect 8668 17824 8720 17876
rect 8392 17799 8444 17808
rect 8392 17765 8401 17799
rect 8401 17765 8435 17799
rect 8435 17765 8444 17799
rect 8392 17756 8444 17765
rect 8576 17756 8628 17808
rect 9680 17824 9732 17876
rect 8484 17731 8536 17740
rect 8484 17697 8493 17731
rect 8493 17697 8527 17731
rect 8527 17697 8536 17731
rect 8484 17688 8536 17697
rect 8668 17731 8720 17740
rect 8668 17697 8677 17731
rect 8677 17697 8711 17731
rect 8711 17697 8720 17731
rect 8668 17688 8720 17697
rect 9404 17731 9456 17740
rect 9404 17697 9413 17731
rect 9413 17697 9447 17731
rect 9447 17697 9456 17731
rect 9404 17688 9456 17697
rect 9864 17688 9916 17740
rect 9128 17620 9180 17672
rect 9680 17620 9732 17672
rect 8300 17552 8352 17604
rect 9036 17552 9088 17604
rect 9404 17552 9456 17604
rect 9496 17552 9548 17604
rect 7564 17484 7616 17536
rect 8392 17484 8444 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 10062 17382 10114 17434
rect 10126 17382 10178 17434
rect 10190 17382 10242 17434
rect 10254 17382 10306 17434
rect 10318 17382 10370 17434
rect 2136 17280 2188 17332
rect 112 17212 164 17264
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 1952 17076 2004 17128
rect 2228 17119 2280 17128
rect 2228 17085 2237 17119
rect 2237 17085 2271 17119
rect 2271 17085 2280 17119
rect 2228 17076 2280 17085
rect 3056 17212 3108 17264
rect 3148 17212 3200 17264
rect 3424 17144 3476 17196
rect 4068 17280 4120 17332
rect 6828 17280 6880 17332
rect 7656 17280 7708 17332
rect 5080 17212 5132 17264
rect 5816 17212 5868 17264
rect 3976 17144 4028 17196
rect 664 17008 716 17060
rect 2596 16940 2648 16992
rect 2964 17119 3016 17128
rect 2964 17085 2973 17119
rect 2973 17085 3007 17119
rect 3007 17085 3016 17119
rect 2964 17076 3016 17085
rect 3700 17008 3752 17060
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 4068 17119 4120 17128
rect 4068 17085 4077 17119
rect 4077 17085 4111 17119
rect 4111 17085 4120 17119
rect 4068 17076 4120 17085
rect 4344 17076 4396 17128
rect 4620 17119 4672 17128
rect 4620 17085 4629 17119
rect 4629 17085 4663 17119
rect 4663 17085 4672 17119
rect 4620 17076 4672 17085
rect 3884 16940 3936 16992
rect 4528 17008 4580 17060
rect 4804 17119 4856 17128
rect 4804 17085 4813 17119
rect 4813 17085 4847 17119
rect 4847 17085 4856 17119
rect 4804 17076 4856 17085
rect 5080 17051 5132 17060
rect 5080 17017 5089 17051
rect 5089 17017 5123 17051
rect 5123 17017 5132 17051
rect 5080 17008 5132 17017
rect 5172 16940 5224 16992
rect 5448 16940 5500 16992
rect 5724 17144 5776 17196
rect 6000 17144 6052 17196
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 7196 17144 7248 17196
rect 8024 17144 8076 17196
rect 8208 17144 8260 17196
rect 6092 17119 6144 17128
rect 6092 17085 6101 17119
rect 6101 17085 6135 17119
rect 6135 17085 6144 17119
rect 6092 17076 6144 17085
rect 7380 17119 7432 17128
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 6276 17008 6328 17060
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 10416 17280 10468 17332
rect 9036 17144 9088 17196
rect 6092 16940 6144 16992
rect 7748 16940 7800 16992
rect 8024 16940 8076 16992
rect 8484 17008 8536 17060
rect 9956 17076 10008 17128
rect 9496 17008 9548 17060
rect 9680 17051 9732 17060
rect 9680 17017 9714 17051
rect 9714 17017 9732 17051
rect 9680 17008 9732 17017
rect 8392 16940 8444 16992
rect 10232 17008 10284 17060
rect 9864 16940 9916 16992
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 10722 16838 10774 16890
rect 10786 16838 10838 16890
rect 10850 16838 10902 16890
rect 10914 16838 10966 16890
rect 10978 16838 11030 16890
rect 4988 16779 5040 16788
rect 4988 16745 4997 16779
rect 4997 16745 5031 16779
rect 5031 16745 5040 16779
rect 4988 16736 5040 16745
rect 5724 16736 5776 16788
rect 6460 16779 6512 16788
rect 6460 16745 6469 16779
rect 6469 16745 6503 16779
rect 6503 16745 6512 16779
rect 6460 16736 6512 16745
rect 6828 16736 6880 16788
rect 3056 16668 3108 16720
rect 4436 16668 4488 16720
rect 1584 16600 1636 16652
rect 2044 16643 2096 16652
rect 2044 16609 2053 16643
rect 2053 16609 2087 16643
rect 2087 16609 2096 16643
rect 2044 16600 2096 16609
rect 2964 16600 3016 16652
rect 388 16532 440 16584
rect 1952 16532 2004 16584
rect 2228 16575 2280 16584
rect 2228 16541 2237 16575
rect 2237 16541 2271 16575
rect 2271 16541 2280 16575
rect 2228 16532 2280 16541
rect 2780 16532 2832 16584
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 3424 16643 3476 16652
rect 3424 16609 3433 16643
rect 3433 16609 3467 16643
rect 3467 16609 3476 16643
rect 3424 16600 3476 16609
rect 5816 16600 5868 16652
rect 6000 16643 6052 16652
rect 6000 16609 6009 16643
rect 6009 16609 6043 16643
rect 6043 16609 6052 16643
rect 6000 16600 6052 16609
rect 6092 16643 6144 16652
rect 6092 16609 6101 16643
rect 6101 16609 6135 16643
rect 6135 16609 6144 16643
rect 6092 16600 6144 16609
rect 7012 16668 7064 16720
rect 7288 16779 7340 16788
rect 7288 16745 7297 16779
rect 7297 16745 7331 16779
rect 7331 16745 7340 16779
rect 7288 16736 7340 16745
rect 7840 16736 7892 16788
rect 8668 16736 8720 16788
rect 7472 16668 7524 16720
rect 7748 16711 7800 16720
rect 7748 16677 7757 16711
rect 7757 16677 7791 16711
rect 7791 16677 7800 16711
rect 7748 16668 7800 16677
rect 8300 16668 8352 16720
rect 9772 16736 9824 16788
rect 10508 16736 10560 16788
rect 6736 16600 6788 16652
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 7932 16600 7984 16652
rect 3516 16575 3568 16584
rect 3516 16541 3525 16575
rect 3525 16541 3559 16575
rect 3559 16541 3568 16575
rect 3516 16532 3568 16541
rect 3884 16575 3936 16584
rect 3884 16541 3893 16575
rect 3893 16541 3927 16575
rect 3927 16541 3936 16575
rect 3884 16532 3936 16541
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 6552 16532 6604 16584
rect 8944 16643 8996 16652
rect 8944 16609 8953 16643
rect 8953 16609 8987 16643
rect 8987 16609 8996 16643
rect 8944 16600 8996 16609
rect 9128 16600 9180 16652
rect 4988 16464 5040 16516
rect 6276 16464 6328 16516
rect 10232 16668 10284 16720
rect 11060 16668 11112 16720
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 11336 16600 11388 16652
rect 9956 16464 10008 16516
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 10324 16464 10376 16516
rect 11060 16464 11112 16516
rect 2780 16439 2832 16448
rect 2780 16405 2789 16439
rect 2789 16405 2823 16439
rect 2823 16405 2832 16439
rect 2780 16396 2832 16405
rect 2964 16439 3016 16448
rect 2964 16405 2973 16439
rect 2973 16405 3007 16439
rect 3007 16405 3016 16439
rect 2964 16396 3016 16405
rect 3516 16396 3568 16448
rect 4252 16396 4304 16448
rect 4804 16396 4856 16448
rect 9404 16439 9456 16448
rect 9404 16405 9413 16439
rect 9413 16405 9447 16439
rect 9447 16405 9456 16439
rect 9404 16396 9456 16405
rect 9496 16396 9548 16448
rect 10140 16396 10192 16448
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 10062 16294 10114 16346
rect 10126 16294 10178 16346
rect 10190 16294 10242 16346
rect 10254 16294 10306 16346
rect 10318 16294 10370 16346
rect 940 16192 992 16244
rect 2412 16235 2464 16244
rect 2412 16201 2421 16235
rect 2421 16201 2455 16235
rect 2455 16201 2464 16235
rect 2412 16192 2464 16201
rect 2780 16192 2832 16244
rect 6368 16192 6420 16244
rect 6828 16192 6880 16244
rect 7564 16192 7616 16244
rect 8668 16192 8720 16244
rect 8852 16192 8904 16244
rect 9956 16192 10008 16244
rect 1676 15988 1728 16040
rect 1952 15988 2004 16040
rect 2504 16056 2556 16108
rect 3056 16124 3108 16176
rect 3424 16056 3476 16108
rect 2504 15920 2556 15972
rect 3148 15988 3200 16040
rect 3516 15988 3568 16040
rect 4252 16099 4304 16108
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 5448 16124 5500 16176
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 4896 16031 4948 16040
rect 4896 15997 4905 16031
rect 4905 15997 4939 16031
rect 4939 15997 4948 16031
rect 4896 15988 4948 15997
rect 8576 16031 8628 16040
rect 8576 15997 8585 16031
rect 8585 15997 8619 16031
rect 8619 15997 8628 16031
rect 8576 15988 8628 15997
rect 9312 16056 9364 16108
rect 9404 16056 9456 16108
rect 1400 15852 1452 15904
rect 2320 15852 2372 15904
rect 6276 15920 6328 15972
rect 8852 16031 8904 16040
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 9772 15920 9824 15972
rect 9312 15852 9364 15904
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 10722 15750 10774 15802
rect 10786 15750 10838 15802
rect 10850 15750 10902 15802
rect 10914 15750 10966 15802
rect 10978 15750 11030 15802
rect 2504 15648 2556 15700
rect 4068 15648 4120 15700
rect 6184 15691 6236 15700
rect 6184 15657 6193 15691
rect 6193 15657 6227 15691
rect 6227 15657 6236 15691
rect 6184 15648 6236 15657
rect 1952 15580 2004 15632
rect 2136 15555 2188 15564
rect 2136 15521 2145 15555
rect 2145 15521 2179 15555
rect 2179 15521 2188 15555
rect 2136 15512 2188 15521
rect 2688 15555 2740 15564
rect 2688 15521 2697 15555
rect 2697 15521 2731 15555
rect 2731 15521 2740 15555
rect 2688 15512 2740 15521
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 4160 15580 4212 15632
rect 4988 15580 5040 15632
rect 6828 15648 6880 15700
rect 7104 15648 7156 15700
rect 7656 15648 7708 15700
rect 8392 15648 8444 15700
rect 8576 15691 8628 15700
rect 8576 15657 8585 15691
rect 8585 15657 8619 15691
rect 8619 15657 8628 15691
rect 8576 15648 8628 15657
rect 9312 15691 9364 15700
rect 9312 15657 9321 15691
rect 9321 15657 9355 15691
rect 9355 15657 9364 15691
rect 9312 15648 9364 15657
rect 9496 15648 9548 15700
rect 7472 15580 7524 15632
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 2596 15444 2648 15496
rect 2872 15444 2924 15496
rect 1768 15376 1820 15428
rect 3700 15555 3752 15564
rect 3700 15521 3709 15555
rect 3709 15521 3743 15555
rect 3743 15521 3752 15555
rect 3700 15512 3752 15521
rect 4068 15444 4120 15496
rect 4804 15555 4856 15564
rect 4804 15521 4813 15555
rect 4813 15521 4847 15555
rect 4847 15521 4856 15555
rect 4804 15512 4856 15521
rect 6276 15512 6328 15564
rect 6552 15555 6604 15564
rect 6552 15521 6561 15555
rect 6561 15521 6595 15555
rect 6595 15521 6604 15555
rect 6552 15512 6604 15521
rect 6736 15555 6788 15564
rect 6736 15521 6745 15555
rect 6745 15521 6779 15555
rect 6779 15521 6788 15555
rect 6736 15512 6788 15521
rect 5816 15444 5868 15496
rect 7196 15512 7248 15564
rect 7288 15512 7340 15564
rect 7840 15555 7892 15564
rect 7840 15521 7849 15555
rect 7849 15521 7883 15555
rect 7883 15521 7892 15555
rect 7840 15512 7892 15521
rect 8208 15512 8260 15564
rect 8392 15555 8444 15564
rect 8392 15521 8401 15555
rect 8401 15521 8435 15555
rect 8435 15521 8444 15555
rect 8392 15512 8444 15521
rect 8668 15555 8720 15564
rect 8668 15521 8677 15555
rect 8677 15521 8711 15555
rect 8711 15521 8720 15555
rect 8668 15512 8720 15521
rect 9772 15580 9824 15632
rect 10692 15580 10744 15632
rect 9312 15512 9364 15564
rect 9496 15555 9548 15564
rect 9496 15521 9505 15555
rect 9505 15521 9539 15555
rect 9539 15521 9548 15555
rect 9496 15512 9548 15521
rect 9956 15555 10008 15564
rect 9956 15521 9965 15555
rect 9965 15521 9999 15555
rect 9999 15521 10008 15555
rect 9956 15512 10008 15521
rect 4344 15376 4396 15428
rect 4620 15419 4672 15428
rect 4620 15385 4629 15419
rect 4629 15385 4663 15419
rect 4663 15385 4672 15419
rect 4620 15376 4672 15385
rect 4804 15376 4856 15428
rect 2044 15308 2096 15360
rect 2964 15308 3016 15360
rect 3332 15308 3384 15360
rect 8852 15376 8904 15428
rect 8944 15419 8996 15428
rect 8944 15385 8953 15419
rect 8953 15385 8987 15419
rect 8987 15385 8996 15419
rect 8944 15376 8996 15385
rect 9220 15376 9272 15428
rect 8208 15308 8260 15360
rect 8576 15308 8628 15360
rect 9588 15444 9640 15496
rect 9404 15308 9456 15360
rect 10600 15308 10652 15360
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 10062 15206 10114 15258
rect 10126 15206 10178 15258
rect 10190 15206 10242 15258
rect 10254 15206 10306 15258
rect 10318 15206 10370 15258
rect 2228 15147 2280 15156
rect 2228 15113 2237 15147
rect 2237 15113 2271 15147
rect 2271 15113 2280 15147
rect 2228 15104 2280 15113
rect 2320 15104 2372 15156
rect 4160 15104 4212 15156
rect 4620 15104 4672 15156
rect 1492 15036 1544 15088
rect 2136 14968 2188 15020
rect 1584 14900 1636 14952
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 2412 14900 2464 14952
rect 1952 14832 2004 14884
rect 2688 15036 2740 15088
rect 2688 14943 2740 14952
rect 2688 14909 2697 14943
rect 2697 14909 2731 14943
rect 2731 14909 2740 14943
rect 2688 14900 2740 14909
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 2872 14900 2924 14909
rect 204 14764 256 14816
rect 1492 14764 1544 14816
rect 1676 14764 1728 14816
rect 2688 14764 2740 14816
rect 2872 14764 2924 14816
rect 3148 15036 3200 15088
rect 6092 15104 6144 15156
rect 7012 15104 7064 15156
rect 3700 14968 3752 15020
rect 5540 15036 5592 15088
rect 8116 15104 8168 15156
rect 8760 15104 8812 15156
rect 8944 15104 8996 15156
rect 9404 15104 9456 15156
rect 9956 15104 10008 15156
rect 3976 14900 4028 14952
rect 5356 14968 5408 15020
rect 6184 14968 6236 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 7748 14968 7800 15020
rect 4712 14900 4764 14952
rect 4896 14943 4948 14952
rect 4896 14909 4905 14943
rect 4905 14909 4939 14943
rect 4939 14909 4948 14943
rect 4896 14900 4948 14909
rect 5080 14943 5132 14952
rect 5080 14909 5089 14943
rect 5089 14909 5123 14943
rect 5123 14909 5132 14943
rect 5080 14900 5132 14909
rect 5816 14943 5868 14952
rect 5816 14909 5825 14943
rect 5825 14909 5859 14943
rect 5859 14909 5868 14943
rect 5816 14900 5868 14909
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 6276 14943 6328 14952
rect 3332 14875 3384 14884
rect 3332 14841 3341 14875
rect 3341 14841 3375 14875
rect 3375 14841 3384 14875
rect 3332 14832 3384 14841
rect 3424 14832 3476 14884
rect 3884 14832 3936 14884
rect 4344 14832 4396 14884
rect 6276 14909 6285 14943
rect 6285 14909 6319 14943
rect 6319 14909 6328 14943
rect 6276 14900 6328 14909
rect 6460 14900 6512 14952
rect 7104 14900 7156 14952
rect 7380 14943 7432 14952
rect 7380 14909 7389 14943
rect 7389 14909 7423 14943
rect 7423 14909 7432 14943
rect 7380 14900 7432 14909
rect 8576 15036 8628 15088
rect 9588 15036 9640 15088
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 8668 14968 8720 15020
rect 8944 14968 8996 15020
rect 9404 14968 9456 15020
rect 10232 14968 10284 15020
rect 6092 14875 6144 14884
rect 6092 14841 6101 14875
rect 6101 14841 6135 14875
rect 6135 14841 6144 14875
rect 6092 14832 6144 14841
rect 6920 14832 6972 14884
rect 4160 14764 4212 14816
rect 5356 14807 5408 14816
rect 5356 14773 5383 14807
rect 5383 14773 5408 14807
rect 5356 14764 5408 14773
rect 7288 14832 7340 14884
rect 8760 14832 8812 14884
rect 10324 14943 10376 14952
rect 10324 14909 10333 14943
rect 10333 14909 10367 14943
rect 10367 14909 10376 14943
rect 10324 14900 10376 14909
rect 10692 14900 10744 14952
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 8944 14764 8996 14816
rect 10324 14764 10376 14816
rect 10416 14764 10468 14816
rect 10600 14764 10652 14816
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 10722 14662 10774 14714
rect 10786 14662 10838 14714
rect 10850 14662 10902 14714
rect 10914 14662 10966 14714
rect 10978 14662 11030 14714
rect 1768 14560 1820 14612
rect 1952 14560 2004 14612
rect 2136 14560 2188 14612
rect 2596 14560 2648 14612
rect 2688 14560 2740 14612
rect 3240 14560 3292 14612
rect 3516 14560 3568 14612
rect 4344 14560 4396 14612
rect 5356 14560 5408 14612
rect 5448 14560 5500 14612
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2504 14467 2556 14476
rect 2504 14433 2513 14467
rect 2513 14433 2547 14467
rect 2547 14433 2556 14467
rect 2504 14424 2556 14433
rect 2596 14467 2648 14476
rect 2596 14433 2605 14467
rect 2605 14433 2639 14467
rect 2639 14433 2648 14467
rect 2596 14424 2648 14433
rect 3148 14424 3200 14476
rect 3240 14424 3292 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 2412 14356 2464 14408
rect 3516 14467 3568 14476
rect 3516 14433 3525 14467
rect 3525 14433 3559 14467
rect 3559 14433 3568 14467
rect 3516 14424 3568 14433
rect 3976 14492 4028 14544
rect 4160 14467 4212 14476
rect 4160 14433 4169 14467
rect 4169 14433 4203 14467
rect 4203 14433 4212 14467
rect 4160 14424 4212 14433
rect 4712 14467 4764 14476
rect 4712 14433 4721 14467
rect 4721 14433 4755 14467
rect 4755 14433 4764 14467
rect 4712 14424 4764 14433
rect 5080 14492 5132 14544
rect 7380 14560 7432 14612
rect 6644 14492 6696 14544
rect 3884 14356 3936 14408
rect 2596 14220 2648 14272
rect 4160 14288 4212 14340
rect 5356 14356 5408 14408
rect 4896 14220 4948 14272
rect 5080 14263 5132 14272
rect 5080 14229 5089 14263
rect 5089 14229 5123 14263
rect 5123 14229 5132 14263
rect 5080 14220 5132 14229
rect 5356 14220 5408 14272
rect 5816 14424 5868 14476
rect 7196 14492 7248 14544
rect 7472 14492 7524 14544
rect 7748 14603 7800 14612
rect 7748 14569 7757 14603
rect 7757 14569 7791 14603
rect 7791 14569 7800 14603
rect 7748 14560 7800 14569
rect 7840 14560 7892 14612
rect 8668 14603 8720 14612
rect 8668 14569 8670 14603
rect 8670 14569 8704 14603
rect 8704 14569 8720 14603
rect 8668 14560 8720 14569
rect 7656 14492 7708 14544
rect 9772 14560 9824 14612
rect 10232 14603 10284 14612
rect 10232 14569 10241 14603
rect 10241 14569 10275 14603
rect 10275 14569 10284 14603
rect 10232 14560 10284 14569
rect 10416 14603 10468 14612
rect 10416 14569 10425 14603
rect 10425 14569 10459 14603
rect 10459 14569 10468 14603
rect 10416 14560 10468 14569
rect 7380 14424 7432 14476
rect 8944 14492 8996 14544
rect 8392 14467 8444 14476
rect 8392 14433 8401 14467
rect 8401 14433 8435 14467
rect 8435 14433 8444 14467
rect 8392 14424 8444 14433
rect 6276 14356 6328 14408
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 6000 14288 6052 14340
rect 7288 14356 7340 14408
rect 7380 14288 7432 14340
rect 8116 14288 8168 14340
rect 8760 14467 8812 14476
rect 8760 14433 8769 14467
rect 8769 14433 8803 14467
rect 8803 14433 8812 14467
rect 8760 14424 8812 14433
rect 10600 14492 10652 14544
rect 8852 14356 8904 14408
rect 9772 14424 9824 14476
rect 9404 14356 9456 14408
rect 10324 14467 10376 14476
rect 10324 14433 10333 14467
rect 10333 14433 10367 14467
rect 10367 14433 10376 14467
rect 10324 14424 10376 14433
rect 11060 14424 11112 14476
rect 10600 14356 10652 14408
rect 10324 14288 10376 14340
rect 11152 14288 11204 14340
rect 5816 14220 5868 14272
rect 7196 14220 7248 14272
rect 8576 14220 8628 14272
rect 9496 14220 9548 14272
rect 9772 14220 9824 14272
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 10062 14118 10114 14170
rect 10126 14118 10178 14170
rect 10190 14118 10242 14170
rect 10254 14118 10306 14170
rect 10318 14118 10370 14170
rect 1400 14016 1452 14068
rect 3424 14016 3476 14068
rect 4712 14016 4764 14068
rect 6276 14016 6328 14068
rect 8484 14016 8536 14068
rect 8852 14016 8904 14068
rect 1400 13880 1452 13932
rect 1676 13880 1728 13932
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 2596 13880 2648 13932
rect 3240 13948 3292 14000
rect 3700 13948 3752 14000
rect 4344 13948 4396 14000
rect 4896 13948 4948 14000
rect 5356 13948 5408 14000
rect 5448 13948 5500 14000
rect 7012 13948 7064 14000
rect 8760 13948 8812 14000
rect 8944 13991 8996 14000
rect 8944 13957 8953 13991
rect 8953 13957 8987 13991
rect 8987 13957 8996 13991
rect 8944 13948 8996 13957
rect 1124 13855 1176 13864
rect 1124 13821 1133 13855
rect 1133 13821 1167 13855
rect 1167 13821 1176 13855
rect 1124 13812 1176 13821
rect 1952 13812 2004 13864
rect 2320 13812 2372 13864
rect 3424 13812 3476 13864
rect 7380 13880 7432 13932
rect 8116 13880 8168 13932
rect 11336 14016 11388 14068
rect 9588 13991 9640 14000
rect 9588 13957 9597 13991
rect 9597 13957 9631 13991
rect 9631 13957 9640 13991
rect 9588 13948 9640 13957
rect 2228 13744 2280 13796
rect 3148 13744 3200 13796
rect 3332 13744 3384 13796
rect 3884 13812 3936 13864
rect 4160 13812 4212 13864
rect 5632 13812 5684 13864
rect 6184 13855 6236 13864
rect 6184 13821 6193 13855
rect 6193 13821 6227 13855
rect 6227 13821 6236 13855
rect 6184 13812 6236 13821
rect 7196 13812 7248 13864
rect 8484 13812 8536 13864
rect 4712 13744 4764 13796
rect 4988 13744 5040 13796
rect 6092 13744 6144 13796
rect 7104 13744 7156 13796
rect 9220 13744 9272 13796
rect 9496 13744 9548 13796
rect 10600 13744 10652 13796
rect 1768 13676 1820 13728
rect 4068 13719 4120 13728
rect 4068 13685 4077 13719
rect 4077 13685 4111 13719
rect 4111 13685 4120 13719
rect 4068 13676 4120 13685
rect 6460 13676 6512 13728
rect 8760 13676 8812 13728
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 10722 13574 10774 13626
rect 10786 13574 10838 13626
rect 10850 13574 10902 13626
rect 10914 13574 10966 13626
rect 10978 13574 11030 13626
rect 1492 13472 1544 13524
rect 1952 13515 2004 13524
rect 1952 13481 1961 13515
rect 1961 13481 1995 13515
rect 1995 13481 2004 13515
rect 1952 13472 2004 13481
rect 2688 13472 2740 13524
rect 2320 13404 2372 13456
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 2044 13379 2096 13388
rect 2044 13345 2053 13379
rect 2053 13345 2087 13379
rect 2087 13345 2096 13379
rect 2044 13336 2096 13345
rect 2872 13336 2924 13388
rect 3240 13379 3292 13388
rect 3240 13345 3249 13379
rect 3249 13345 3283 13379
rect 3283 13345 3292 13379
rect 3240 13336 3292 13345
rect 4068 13472 4120 13524
rect 3700 13404 3752 13456
rect 3332 13268 3384 13320
rect 3792 13379 3844 13388
rect 3792 13345 3801 13379
rect 3801 13345 3835 13379
rect 3835 13345 3844 13379
rect 3792 13336 3844 13345
rect 4160 13404 4212 13456
rect 4528 13472 4580 13524
rect 4896 13472 4948 13524
rect 7932 13472 7984 13524
rect 4620 13379 4672 13388
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 4896 13379 4948 13388
rect 4896 13345 4905 13379
rect 4905 13345 4939 13379
rect 4939 13345 4948 13379
rect 4896 13336 4948 13345
rect 4160 13268 4212 13320
rect 4344 13311 4396 13320
rect 4344 13277 4353 13311
rect 4353 13277 4387 13311
rect 4387 13277 4396 13311
rect 7012 13404 7064 13456
rect 4344 13268 4396 13277
rect 2780 13175 2832 13184
rect 2780 13141 2789 13175
rect 2789 13141 2823 13175
rect 2823 13141 2832 13175
rect 2780 13132 2832 13141
rect 2964 13175 3016 13184
rect 2964 13141 2973 13175
rect 2973 13141 3007 13175
rect 3007 13141 3016 13175
rect 2964 13132 3016 13141
rect 3332 13132 3384 13184
rect 3884 13200 3936 13252
rect 6368 13336 6420 13388
rect 6552 13336 6604 13388
rect 6920 13336 6972 13388
rect 7932 13379 7984 13388
rect 7932 13345 7941 13379
rect 7941 13345 7975 13379
rect 7975 13345 7984 13379
rect 7932 13336 7984 13345
rect 8116 13379 8168 13388
rect 8116 13345 8125 13379
rect 8125 13345 8159 13379
rect 8159 13345 8168 13379
rect 8116 13336 8168 13345
rect 9220 13472 9272 13524
rect 9588 13404 9640 13456
rect 8484 13379 8536 13388
rect 8484 13345 8493 13379
rect 8493 13345 8527 13379
rect 8527 13345 8536 13379
rect 8484 13336 8536 13345
rect 9864 13336 9916 13388
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 7012 13268 7064 13320
rect 9220 13268 9272 13320
rect 9588 13268 9640 13320
rect 7288 13200 7340 13252
rect 4896 13132 4948 13184
rect 4988 13175 5040 13184
rect 4988 13141 4997 13175
rect 4997 13141 5031 13175
rect 5031 13141 5040 13175
rect 4988 13132 5040 13141
rect 7656 13175 7708 13184
rect 7656 13141 7665 13175
rect 7665 13141 7699 13175
rect 7699 13141 7708 13175
rect 7656 13132 7708 13141
rect 8024 13132 8076 13184
rect 9496 13132 9548 13184
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 10062 13030 10114 13082
rect 10126 13030 10178 13082
rect 10190 13030 10242 13082
rect 10254 13030 10306 13082
rect 10318 13030 10370 13082
rect 2596 12928 2648 12980
rect 3148 12928 3200 12980
rect 3516 12928 3568 12980
rect 9128 12971 9180 12980
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 9956 12928 10008 12980
rect 20 12724 72 12776
rect 4620 12860 4672 12912
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 1308 12724 1360 12776
rect 2228 12724 2280 12776
rect 2780 12792 2832 12844
rect 2688 12699 2740 12708
rect 2688 12665 2697 12699
rect 2697 12665 2731 12699
rect 2731 12665 2740 12699
rect 2688 12656 2740 12665
rect 2412 12588 2464 12640
rect 3148 12724 3200 12776
rect 4160 12792 4212 12844
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 5356 12860 5408 12912
rect 8668 12860 8720 12912
rect 9312 12860 9364 12912
rect 4528 12767 4580 12776
rect 4528 12733 4537 12767
rect 4537 12733 4571 12767
rect 4571 12733 4580 12767
rect 4528 12724 4580 12733
rect 5448 12724 5500 12776
rect 6000 12767 6052 12776
rect 6000 12733 6009 12767
rect 6009 12733 6043 12767
rect 6043 12733 6052 12767
rect 6000 12724 6052 12733
rect 6092 12767 6144 12776
rect 6092 12733 6101 12767
rect 6101 12733 6135 12767
rect 6135 12733 6144 12767
rect 6092 12724 6144 12733
rect 6184 12724 6236 12776
rect 2872 12656 2924 12708
rect 3700 12656 3752 12708
rect 4160 12656 4212 12708
rect 5080 12699 5132 12708
rect 5080 12665 5089 12699
rect 5089 12665 5123 12699
rect 5123 12665 5132 12699
rect 5080 12656 5132 12665
rect 5724 12656 5776 12708
rect 7012 12724 7064 12776
rect 7196 12699 7248 12708
rect 7196 12665 7205 12699
rect 7205 12665 7239 12699
rect 7239 12665 7248 12699
rect 7196 12656 7248 12665
rect 8024 12792 8076 12844
rect 7656 12724 7708 12776
rect 7748 12767 7800 12776
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 7840 12767 7892 12776
rect 7840 12733 7849 12767
rect 7849 12733 7883 12767
rect 7883 12733 7892 12767
rect 7840 12724 7892 12733
rect 7932 12767 7984 12776
rect 7932 12733 7941 12767
rect 7941 12733 7975 12767
rect 7975 12733 7984 12767
rect 7932 12724 7984 12733
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 9680 12792 9732 12844
rect 10140 12767 10192 12776
rect 10140 12733 10149 12767
rect 10149 12733 10183 12767
rect 10183 12733 10192 12767
rect 10140 12724 10192 12733
rect 10416 12767 10468 12776
rect 10416 12733 10425 12767
rect 10425 12733 10459 12767
rect 10459 12733 10468 12767
rect 10416 12724 10468 12733
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 9680 12656 9732 12708
rect 10324 12656 10376 12708
rect 3424 12588 3476 12640
rect 3792 12588 3844 12640
rect 7104 12588 7156 12640
rect 7472 12588 7524 12640
rect 7656 12588 7708 12640
rect 7840 12588 7892 12640
rect 8484 12588 8536 12640
rect 9496 12588 9548 12640
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 10722 12486 10774 12538
rect 10786 12486 10838 12538
rect 10850 12486 10902 12538
rect 10914 12486 10966 12538
rect 10978 12486 11030 12538
rect 1584 12384 1636 12436
rect 2228 12359 2280 12368
rect 2228 12325 2237 12359
rect 2237 12325 2271 12359
rect 2271 12325 2280 12359
rect 2228 12316 2280 12325
rect 1676 12248 1728 12300
rect 1768 12248 1820 12300
rect 2688 12427 2740 12436
rect 2688 12393 2697 12427
rect 2697 12393 2731 12427
rect 2731 12393 2740 12427
rect 2688 12384 2740 12393
rect 3056 12384 3108 12436
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 4988 12384 5040 12436
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 2504 12316 2556 12368
rect 2688 12248 2740 12300
rect 2780 12248 2832 12300
rect 3792 12291 3844 12300
rect 3792 12257 3801 12291
rect 3801 12257 3835 12291
rect 3835 12257 3844 12291
rect 3792 12248 3844 12257
rect 4068 12248 4120 12300
rect 4896 12316 4948 12368
rect 5540 12316 5592 12368
rect 6736 12384 6788 12436
rect 7196 12316 7248 12368
rect 2964 12180 3016 12232
rect 3332 12223 3384 12232
rect 3332 12189 3341 12223
rect 3341 12189 3375 12223
rect 3375 12189 3384 12223
rect 3332 12180 3384 12189
rect 4896 12180 4948 12232
rect 1952 12112 2004 12164
rect 2688 12112 2740 12164
rect 4804 12155 4856 12164
rect 4804 12121 4813 12155
rect 4813 12121 4847 12155
rect 4847 12121 4856 12155
rect 4804 12112 4856 12121
rect 4988 12112 5040 12164
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 5356 12248 5408 12300
rect 6368 12291 6420 12300
rect 6368 12257 6377 12291
rect 6377 12257 6411 12291
rect 6411 12257 6420 12291
rect 6368 12248 6420 12257
rect 7104 12248 7156 12300
rect 7380 12248 7432 12300
rect 8484 12384 8536 12436
rect 9312 12384 9364 12436
rect 10140 12384 10192 12436
rect 7932 12316 7984 12368
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 8116 12248 8168 12300
rect 10600 12359 10652 12368
rect 10600 12325 10609 12359
rect 10609 12325 10643 12359
rect 10643 12325 10652 12359
rect 10600 12316 10652 12325
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 6460 12180 6512 12232
rect 7012 12223 7064 12232
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9128 12291 9180 12300
rect 9128 12257 9137 12291
rect 9137 12257 9171 12291
rect 9171 12257 9180 12291
rect 9128 12248 9180 12257
rect 9312 12291 9364 12300
rect 9312 12257 9321 12291
rect 9321 12257 9355 12291
rect 9355 12257 9364 12291
rect 9312 12248 9364 12257
rect 9772 12291 9824 12300
rect 9772 12257 9781 12291
rect 9781 12257 9815 12291
rect 9815 12257 9824 12291
rect 9772 12248 9824 12257
rect 10416 12291 10468 12300
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 9220 12180 9272 12232
rect 10508 12180 10560 12232
rect 5264 12112 5316 12164
rect 6644 12112 6696 12164
rect 10600 12112 10652 12164
rect 1492 12044 1544 12096
rect 2044 12087 2096 12096
rect 2044 12053 2053 12087
rect 2053 12053 2087 12087
rect 2087 12053 2096 12087
rect 2044 12044 2096 12053
rect 2320 12044 2372 12096
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 4712 12044 4764 12096
rect 6184 12044 6236 12096
rect 6736 12044 6788 12096
rect 8116 12044 8168 12096
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 10062 11942 10114 11994
rect 10126 11942 10178 11994
rect 10190 11942 10242 11994
rect 10254 11942 10306 11994
rect 10318 11942 10370 11994
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 3240 11883 3292 11892
rect 3240 11849 3249 11883
rect 3249 11849 3283 11883
rect 3283 11849 3292 11883
rect 3240 11840 3292 11849
rect 3332 11840 3384 11892
rect 5908 11840 5960 11892
rect 6736 11883 6788 11892
rect 6736 11849 6745 11883
rect 6745 11849 6779 11883
rect 6779 11849 6788 11883
rect 6736 11840 6788 11849
rect 7012 11840 7064 11892
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 1400 11704 1452 11756
rect 1584 11679 1636 11688
rect 1584 11645 1593 11679
rect 1593 11645 1627 11679
rect 1627 11645 1636 11679
rect 1584 11636 1636 11645
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 2320 11704 2372 11756
rect 2504 11636 2556 11688
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 3516 11636 3568 11688
rect 5632 11636 5684 11688
rect 6184 11679 6236 11688
rect 6184 11645 6193 11679
rect 6193 11645 6227 11679
rect 6227 11645 6236 11679
rect 6184 11636 6236 11645
rect 6920 11679 6972 11688
rect 6920 11645 6929 11679
rect 6929 11645 6963 11679
rect 6963 11645 6972 11679
rect 6920 11636 6972 11645
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 8024 11704 8076 11756
rect 4804 11568 4856 11620
rect 8484 11704 8536 11756
rect 9128 11840 9180 11892
rect 10508 11840 10560 11892
rect 8852 11704 8904 11756
rect 9772 11704 9824 11756
rect 10140 11704 10192 11756
rect 10048 11679 10100 11688
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10048 11636 10100 11645
rect 10600 11679 10652 11688
rect 10600 11645 10609 11679
rect 10609 11645 10643 11679
rect 10643 11645 10652 11679
rect 10600 11636 10652 11645
rect 11060 11636 11112 11688
rect 1400 11543 1452 11552
rect 1400 11509 1409 11543
rect 1409 11509 1443 11543
rect 1443 11509 1452 11543
rect 1400 11500 1452 11509
rect 1584 11500 1636 11552
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 6184 11500 6236 11552
rect 7380 11500 7432 11552
rect 8024 11500 8076 11552
rect 8668 11500 8720 11552
rect 9588 11568 9640 11620
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 10722 11398 10774 11450
rect 10786 11398 10838 11450
rect 10850 11398 10902 11450
rect 10914 11398 10966 11450
rect 10978 11398 11030 11450
rect 1768 11339 1820 11348
rect 1768 11305 1777 11339
rect 1777 11305 1811 11339
rect 1811 11305 1820 11339
rect 1768 11296 1820 11305
rect 2044 11296 2096 11348
rect 4068 11296 4120 11348
rect 4252 11296 4304 11348
rect 4712 11339 4764 11348
rect 4712 11305 4721 11339
rect 4721 11305 4755 11339
rect 4755 11305 4764 11339
rect 4712 11296 4764 11305
rect 4896 11339 4948 11348
rect 4896 11305 4905 11339
rect 4905 11305 4939 11339
rect 4939 11305 4948 11339
rect 4896 11296 4948 11305
rect 1952 11228 2004 11280
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 2320 11160 2372 11212
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 1860 11024 1912 11076
rect 3424 11160 3476 11212
rect 3976 11160 4028 11212
rect 4252 11203 4304 11212
rect 4252 11169 4261 11203
rect 4261 11169 4295 11203
rect 4295 11169 4304 11203
rect 4252 11160 4304 11169
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 4712 11160 4764 11212
rect 5264 11160 5316 11212
rect 5816 11296 5868 11348
rect 6184 11339 6236 11348
rect 6184 11305 6193 11339
rect 6193 11305 6227 11339
rect 6227 11305 6236 11339
rect 6184 11296 6236 11305
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 8852 11271 8904 11280
rect 8852 11237 8861 11271
rect 8861 11237 8895 11271
rect 8895 11237 8904 11271
rect 8852 11228 8904 11237
rect 9496 11228 9548 11280
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 5908 11160 5960 11212
rect 6460 11160 6512 11212
rect 8576 11160 8628 11212
rect 8760 11160 8812 11212
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9128 11160 9180 11212
rect 9404 11203 9456 11212
rect 9404 11169 9413 11203
rect 9413 11169 9447 11203
rect 9447 11169 9456 11203
rect 9404 11160 9456 11169
rect 9588 11160 9640 11212
rect 3608 11024 3660 11076
rect 5632 11067 5684 11076
rect 5632 11033 5641 11067
rect 5641 11033 5675 11067
rect 5675 11033 5684 11067
rect 5632 11024 5684 11033
rect 6644 11135 6696 11144
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6644 11092 6696 11101
rect 7196 11092 7248 11144
rect 9772 11092 9824 11144
rect 10600 11092 10652 11144
rect 7840 11024 7892 11076
rect 7932 11024 7984 11076
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 10062 10854 10114 10906
rect 10126 10854 10178 10906
rect 10190 10854 10242 10906
rect 10254 10854 10306 10906
rect 10318 10854 10370 10906
rect 1952 10752 2004 10804
rect 2228 10795 2280 10804
rect 2228 10761 2237 10795
rect 2237 10761 2271 10795
rect 2271 10761 2280 10795
rect 2228 10752 2280 10761
rect 5448 10752 5500 10804
rect 6276 10752 6328 10804
rect 6644 10752 6696 10804
rect 7472 10752 7524 10804
rect 3240 10684 3292 10736
rect 4160 10684 4212 10736
rect 4344 10684 4396 10736
rect 1124 10591 1176 10600
rect 1124 10557 1133 10591
rect 1133 10557 1167 10591
rect 1167 10557 1176 10591
rect 1124 10548 1176 10557
rect 1308 10591 1360 10600
rect 1308 10557 1317 10591
rect 1317 10557 1351 10591
rect 1351 10557 1360 10591
rect 1308 10548 1360 10557
rect 2320 10591 2372 10600
rect 2320 10557 2329 10591
rect 2329 10557 2363 10591
rect 2363 10557 2372 10591
rect 2320 10548 2372 10557
rect 3976 10659 4028 10668
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 3792 10548 3844 10600
rect 5724 10684 5776 10736
rect 6460 10684 6512 10736
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 5632 10591 5684 10600
rect 5632 10557 5641 10591
rect 5641 10557 5675 10591
rect 5675 10557 5684 10591
rect 5632 10548 5684 10557
rect 7196 10684 7248 10736
rect 7932 10684 7984 10736
rect 4712 10480 4764 10532
rect 6276 10480 6328 10532
rect 3332 10412 3384 10464
rect 5448 10412 5500 10464
rect 6368 10412 6420 10464
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 8208 10616 8260 10668
rect 7012 10523 7064 10532
rect 7012 10489 7021 10523
rect 7021 10489 7055 10523
rect 7055 10489 7064 10523
rect 7932 10591 7984 10600
rect 7932 10557 7941 10591
rect 7941 10557 7975 10591
rect 7975 10557 7984 10591
rect 7932 10548 7984 10557
rect 8852 10548 8904 10600
rect 9312 10548 9364 10600
rect 9772 10591 9824 10600
rect 9772 10557 9781 10591
rect 9781 10557 9815 10591
rect 9815 10557 9824 10591
rect 9772 10548 9824 10557
rect 7012 10480 7064 10489
rect 8944 10455 8996 10464
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 10600 10412 10652 10464
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 10722 10310 10774 10362
rect 10786 10310 10838 10362
rect 10850 10310 10902 10362
rect 10914 10310 10966 10362
rect 10978 10310 11030 10362
rect 1308 10208 1360 10260
rect 1768 10208 1820 10260
rect 2320 10208 2372 10260
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 2688 10072 2740 10124
rect 2872 10072 2924 10124
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 2780 10004 2832 10056
rect 3792 10115 3844 10124
rect 3792 10081 3801 10115
rect 3801 10081 3835 10115
rect 3835 10081 3844 10115
rect 3792 10072 3844 10081
rect 3884 10115 3936 10124
rect 3884 10081 3893 10115
rect 3893 10081 3927 10115
rect 3927 10081 3936 10115
rect 3884 10072 3936 10081
rect 6000 10140 6052 10192
rect 4160 10004 4212 10056
rect 4896 10115 4948 10124
rect 4896 10081 4905 10115
rect 4905 10081 4939 10115
rect 4939 10081 4948 10115
rect 4896 10072 4948 10081
rect 5448 10072 5500 10124
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 3976 9936 4028 9988
rect 4712 9936 4764 9988
rect 1676 9911 1728 9920
rect 1676 9877 1685 9911
rect 1685 9877 1719 9911
rect 1719 9877 1728 9911
rect 1676 9868 1728 9877
rect 2596 9868 2648 9920
rect 5908 9936 5960 9988
rect 6184 10115 6236 10124
rect 6184 10081 6193 10115
rect 6193 10081 6227 10115
rect 6227 10081 6236 10115
rect 6184 10072 6236 10081
rect 6276 10072 6328 10124
rect 7012 10251 7064 10260
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 7288 10208 7340 10260
rect 9404 10208 9456 10260
rect 10416 10251 10468 10260
rect 10416 10217 10425 10251
rect 10425 10217 10459 10251
rect 10459 10217 10468 10251
rect 10416 10208 10468 10217
rect 9496 10140 9548 10192
rect 6736 10072 6788 10124
rect 7196 10072 7248 10124
rect 8852 10115 8904 10124
rect 8852 10081 8861 10115
rect 8861 10081 8895 10115
rect 8895 10081 8904 10115
rect 8852 10072 8904 10081
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 6368 9936 6420 9988
rect 8668 9936 8720 9988
rect 9680 10004 9732 10056
rect 9772 10004 9824 10056
rect 9956 9979 10008 9988
rect 9956 9945 9965 9979
rect 9965 9945 9999 9979
rect 9999 9945 10008 9979
rect 10600 10140 10652 10192
rect 9956 9936 10008 9945
rect 6184 9868 6236 9920
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 10062 9766 10114 9818
rect 10126 9766 10178 9818
rect 10190 9766 10242 9818
rect 10254 9766 10306 9818
rect 10318 9766 10370 9818
rect 4896 9664 4948 9716
rect 6276 9664 6328 9716
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 6736 9707 6788 9716
rect 6736 9673 6745 9707
rect 6745 9673 6779 9707
rect 6779 9673 6788 9707
rect 6736 9664 6788 9673
rect 8852 9664 8904 9716
rect 1860 9596 1912 9648
rect 3516 9596 3568 9648
rect 4252 9596 4304 9648
rect 5080 9596 5132 9648
rect 5356 9596 5408 9648
rect 6000 9639 6052 9648
rect 6000 9605 6009 9639
rect 6009 9605 6043 9639
rect 6043 9605 6052 9639
rect 6000 9596 6052 9605
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 1308 9460 1360 9512
rect 2596 9460 2648 9512
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 2320 9392 2372 9444
rect 3884 9392 3936 9444
rect 4712 9460 4764 9512
rect 4988 9460 5040 9512
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5724 9571 5776 9580
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 7288 9528 7340 9580
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 9772 9664 9824 9716
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 9496 9596 9548 9648
rect 5080 9460 5132 9469
rect 5448 9460 5500 9512
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 7196 9460 7248 9512
rect 8484 9460 8536 9512
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 9496 9503 9548 9512
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 9956 9460 10008 9512
rect 10600 9460 10652 9512
rect 6000 9392 6052 9444
rect 6736 9392 6788 9444
rect 10508 9392 10560 9444
rect 7196 9324 7248 9376
rect 7840 9324 7892 9376
rect 8944 9324 8996 9376
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 10722 9222 10774 9274
rect 10786 9222 10838 9274
rect 10850 9222 10902 9274
rect 10914 9222 10966 9274
rect 10978 9222 11030 9274
rect 1308 9163 1360 9172
rect 1308 9129 1317 9163
rect 1317 9129 1351 9163
rect 1351 9129 1360 9163
rect 1308 9120 1360 9129
rect 2872 9120 2924 9172
rect 3976 9120 4028 9172
rect 4160 9120 4212 9172
rect 4712 9163 4764 9172
rect 4712 9129 4721 9163
rect 4721 9129 4755 9163
rect 4755 9129 4764 9163
rect 4712 9120 4764 9129
rect 5080 9120 5132 9172
rect 7656 9120 7708 9172
rect 9496 9120 9548 9172
rect 1952 9027 2004 9036
rect 1952 8993 1961 9027
rect 1961 8993 1995 9027
rect 1995 8993 2004 9027
rect 1952 8984 2004 8993
rect 2688 9052 2740 9104
rect 2320 8984 2372 9036
rect 940 8916 992 8968
rect 1400 8916 1452 8968
rect 3240 9027 3292 9036
rect 3240 8993 3249 9027
rect 3249 8993 3283 9027
rect 3283 8993 3292 9027
rect 3240 8984 3292 8993
rect 3332 8916 3384 8968
rect 3516 8984 3568 9036
rect 3884 9027 3936 9036
rect 3884 8993 3893 9027
rect 3893 8993 3927 9027
rect 3927 8993 3936 9027
rect 3884 8984 3936 8993
rect 4160 8984 4212 9036
rect 8300 9052 8352 9104
rect 5080 8984 5132 9036
rect 6092 8984 6144 9036
rect 8668 8984 8720 9036
rect 9220 9095 9272 9104
rect 9220 9061 9229 9095
rect 9229 9061 9263 9095
rect 9263 9061 9272 9095
rect 9220 9052 9272 9061
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 8024 8959 8076 8968
rect 8024 8925 8033 8959
rect 8033 8925 8067 8959
rect 8067 8925 8076 8959
rect 8024 8916 8076 8925
rect 2596 8848 2648 8900
rect 6092 8848 6144 8900
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 8484 8916 8536 8968
rect 9496 8916 9548 8968
rect 10600 8916 10652 8968
rect 8576 8848 8628 8900
rect 7932 8780 7984 8832
rect 8300 8780 8352 8832
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 10062 8678 10114 8730
rect 10126 8678 10178 8730
rect 10190 8678 10242 8730
rect 10254 8678 10306 8730
rect 10318 8678 10370 8730
rect 4160 8619 4212 8628
rect 4160 8585 4169 8619
rect 4169 8585 4203 8619
rect 4203 8585 4212 8619
rect 4160 8576 4212 8585
rect 7748 8576 7800 8628
rect 8576 8576 8628 8628
rect 9588 8619 9640 8628
rect 9588 8585 9597 8619
rect 9597 8585 9631 8619
rect 9631 8585 9640 8619
rect 9588 8576 9640 8585
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 2136 8508 2188 8560
rect 8024 8508 8076 8560
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 3516 8372 3568 8424
rect 7932 8372 7984 8424
rect 3240 8236 3292 8288
rect 3516 8236 3568 8288
rect 4160 8304 4212 8356
rect 7840 8347 7892 8356
rect 7840 8313 7849 8347
rect 7849 8313 7883 8347
rect 7883 8313 7892 8347
rect 7840 8304 7892 8313
rect 9404 8508 9456 8560
rect 10416 8508 10468 8560
rect 8300 8440 8352 8492
rect 8852 8440 8904 8492
rect 8208 8304 8260 8356
rect 8576 8347 8628 8356
rect 8576 8313 8585 8347
rect 8585 8313 8619 8347
rect 8619 8313 8628 8347
rect 8576 8304 8628 8313
rect 8300 8236 8352 8288
rect 8944 8415 8996 8424
rect 8944 8381 8953 8415
rect 8953 8381 8987 8415
rect 8987 8381 8996 8415
rect 8944 8372 8996 8381
rect 9404 8372 9456 8424
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 10048 8415 10100 8424
rect 10048 8381 10057 8415
rect 10057 8381 10091 8415
rect 10091 8381 10100 8415
rect 10048 8372 10100 8381
rect 10140 8347 10192 8356
rect 10140 8313 10149 8347
rect 10149 8313 10183 8347
rect 10183 8313 10192 8347
rect 10140 8304 10192 8313
rect 9128 8236 9180 8288
rect 9404 8236 9456 8288
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 10722 8134 10774 8186
rect 10786 8134 10838 8186
rect 10850 8134 10902 8186
rect 10914 8134 10966 8186
rect 10978 8134 11030 8186
rect 2136 8032 2188 8084
rect 2504 8032 2556 8084
rect 6552 8032 6604 8084
rect 8392 8032 8444 8084
rect 1400 7896 1452 7948
rect 1952 7939 2004 7948
rect 1952 7905 1961 7939
rect 1961 7905 1995 7939
rect 1995 7905 2004 7939
rect 1952 7896 2004 7905
rect 3148 7896 3200 7948
rect 6460 7939 6512 7948
rect 6460 7905 6469 7939
rect 6469 7905 6503 7939
rect 6503 7905 6512 7939
rect 6460 7896 6512 7905
rect 6552 7896 6604 7948
rect 7380 7896 7432 7948
rect 2504 7828 2556 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 7656 7939 7708 7948
rect 7656 7905 7665 7939
rect 7665 7905 7699 7939
rect 7699 7905 7708 7939
rect 7656 7896 7708 7905
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 7932 7964 7984 8016
rect 9128 7964 9180 8016
rect 10140 8032 10192 8084
rect 6736 7828 6788 7837
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 7564 7828 7616 7880
rect 7656 7760 7708 7812
rect 8392 7937 8444 7948
rect 8392 7903 8401 7937
rect 8401 7903 8435 7937
rect 8435 7903 8444 7937
rect 8392 7896 8444 7903
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 8392 7692 8444 7744
rect 8944 7939 8996 7948
rect 8944 7905 8953 7939
rect 8953 7905 8987 7939
rect 8987 7905 8996 7939
rect 8944 7896 8996 7905
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 10416 7939 10468 7948
rect 10416 7905 10425 7939
rect 10425 7905 10459 7939
rect 10459 7905 10468 7939
rect 10416 7896 10468 7905
rect 9864 7828 9916 7880
rect 9956 7828 10008 7880
rect 9404 7760 9456 7812
rect 10048 7803 10100 7812
rect 10048 7769 10057 7803
rect 10057 7769 10091 7803
rect 10091 7769 10100 7803
rect 10048 7760 10100 7769
rect 9772 7692 9824 7744
rect 10508 7692 10560 7744
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 10062 7590 10114 7642
rect 10126 7590 10178 7642
rect 10190 7590 10242 7642
rect 10254 7590 10306 7642
rect 10318 7590 10370 7642
rect 1584 7488 1636 7540
rect 1400 7420 1452 7472
rect 1584 7352 1636 7404
rect 2136 7488 2188 7540
rect 3148 7488 3200 7540
rect 4068 7488 4120 7540
rect 6736 7531 6788 7540
rect 6736 7497 6745 7531
rect 6745 7497 6779 7531
rect 6779 7497 6788 7531
rect 6736 7488 6788 7497
rect 2412 7463 2464 7472
rect 2412 7429 2421 7463
rect 2421 7429 2455 7463
rect 2455 7429 2464 7463
rect 2412 7420 2464 7429
rect 5540 7420 5592 7472
rect 7380 7488 7432 7540
rect 7564 7531 7616 7540
rect 7564 7497 7573 7531
rect 7573 7497 7607 7531
rect 7607 7497 7616 7531
rect 7564 7488 7616 7497
rect 7656 7531 7708 7540
rect 7656 7497 7665 7531
rect 7665 7497 7699 7531
rect 7699 7497 7708 7531
rect 7656 7488 7708 7497
rect 8944 7488 8996 7540
rect 9680 7488 9732 7540
rect 2780 7352 2832 7404
rect 2412 7284 2464 7336
rect 2872 7284 2924 7336
rect 3516 7284 3568 7336
rect 3884 7284 3936 7336
rect 4252 7284 4304 7336
rect 5080 7284 5132 7336
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 5908 7327 5960 7336
rect 5908 7293 5917 7327
rect 5917 7293 5951 7327
rect 5951 7293 5960 7327
rect 5908 7284 5960 7293
rect 2228 7216 2280 7268
rect 5816 7216 5868 7268
rect 6184 7327 6236 7336
rect 6184 7293 6193 7327
rect 6193 7293 6227 7327
rect 6227 7293 6236 7327
rect 6184 7284 6236 7293
rect 6368 7327 6420 7336
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 6552 7284 6604 7336
rect 7564 7352 7616 7404
rect 6460 7216 6512 7268
rect 6736 7216 6788 7268
rect 1584 7148 1636 7200
rect 1860 7148 1912 7200
rect 3516 7148 3568 7200
rect 4988 7148 5040 7200
rect 6276 7191 6328 7200
rect 6276 7157 6285 7191
rect 6285 7157 6319 7191
rect 6319 7157 6328 7191
rect 6276 7148 6328 7157
rect 6552 7148 6604 7200
rect 7012 7148 7064 7200
rect 7196 7284 7248 7336
rect 8760 7352 8812 7404
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 8484 7284 8536 7336
rect 9128 7284 9180 7336
rect 9864 7284 9916 7336
rect 9956 7284 10008 7336
rect 10508 7327 10560 7336
rect 10508 7293 10517 7327
rect 10517 7293 10551 7327
rect 10551 7293 10560 7327
rect 10508 7284 10560 7293
rect 8760 7216 8812 7268
rect 9864 7148 9916 7200
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 10722 7046 10774 7098
rect 10786 7046 10838 7098
rect 10850 7046 10902 7098
rect 10914 7046 10966 7098
rect 10978 7046 11030 7098
rect 2228 6987 2280 6996
rect 2228 6953 2237 6987
rect 2237 6953 2271 6987
rect 2271 6953 2280 6987
rect 2228 6944 2280 6953
rect 1952 6876 2004 6928
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 1492 6740 1544 6792
rect 2228 6851 2280 6860
rect 2228 6817 2237 6851
rect 2237 6817 2271 6851
rect 2271 6817 2280 6851
rect 2228 6808 2280 6817
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 2688 6851 2740 6860
rect 2688 6817 2697 6851
rect 2697 6817 2731 6851
rect 2731 6817 2740 6851
rect 2688 6808 2740 6817
rect 2872 6808 2924 6860
rect 3884 6944 3936 6996
rect 5908 6944 5960 6996
rect 8208 6944 8260 6996
rect 9128 6944 9180 6996
rect 9588 6944 9640 6996
rect 3240 6851 3292 6860
rect 3240 6817 3249 6851
rect 3249 6817 3283 6851
rect 3283 6817 3292 6851
rect 3240 6808 3292 6817
rect 4068 6808 4120 6860
rect 4712 6808 4764 6860
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 1400 6672 1452 6724
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 6184 6808 6236 6860
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 6920 6808 6972 6860
rect 7472 6876 7524 6928
rect 5172 6672 5224 6724
rect 6828 6740 6880 6792
rect 8024 6851 8076 6860
rect 8024 6817 8033 6851
rect 8033 6817 8067 6851
rect 8067 6817 8076 6851
rect 8024 6808 8076 6817
rect 8208 6808 8260 6860
rect 9220 6808 9272 6860
rect 9496 6808 9548 6860
rect 1492 6604 1544 6656
rect 3424 6604 3476 6656
rect 3884 6604 3936 6656
rect 4620 6604 4672 6656
rect 5540 6604 5592 6656
rect 6828 6604 6880 6656
rect 8852 6740 8904 6792
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 10062 6502 10114 6554
rect 10126 6502 10178 6554
rect 10190 6502 10242 6554
rect 10254 6502 10306 6554
rect 10318 6502 10370 6554
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 3516 6400 3568 6452
rect 1400 6196 1452 6248
rect 2044 6196 2096 6248
rect 2136 6239 2188 6248
rect 2136 6205 2145 6239
rect 2145 6205 2179 6239
rect 2179 6205 2188 6239
rect 2136 6196 2188 6205
rect 1952 6128 2004 6180
rect 3240 6239 3292 6248
rect 3240 6205 3249 6239
rect 3249 6205 3283 6239
rect 3283 6205 3292 6239
rect 3240 6196 3292 6205
rect 3424 6239 3476 6248
rect 3424 6205 3433 6239
rect 3433 6205 3467 6239
rect 3467 6205 3476 6239
rect 3424 6196 3476 6205
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 5264 6400 5316 6452
rect 5724 6400 5776 6452
rect 6368 6443 6420 6452
rect 6368 6409 6377 6443
rect 6377 6409 6411 6443
rect 6411 6409 6420 6443
rect 6368 6400 6420 6409
rect 7104 6443 7156 6452
rect 7104 6409 7113 6443
rect 7113 6409 7147 6443
rect 7147 6409 7156 6443
rect 7104 6400 7156 6409
rect 3792 6375 3844 6384
rect 3792 6341 3801 6375
rect 3801 6341 3835 6375
rect 3835 6341 3844 6375
rect 3792 6332 3844 6341
rect 4252 6264 4304 6316
rect 7288 6332 7340 6384
rect 4988 6239 5040 6248
rect 4988 6205 4997 6239
rect 4997 6205 5031 6239
rect 5031 6205 5040 6239
rect 4988 6196 5040 6205
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 5540 6196 5592 6205
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 6460 6239 6512 6248
rect 6460 6205 6469 6239
rect 6469 6205 6503 6239
rect 6503 6205 6512 6239
rect 6460 6196 6512 6205
rect 7380 6264 7432 6316
rect 7472 6264 7524 6316
rect 5080 6128 5132 6180
rect 5908 6128 5960 6180
rect 6092 6128 6144 6180
rect 6552 6128 6604 6180
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 6920 6196 6972 6205
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 8116 6196 8168 6248
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 10416 6196 10468 6248
rect 7104 6128 7156 6180
rect 2412 6060 2464 6112
rect 2964 6060 3016 6112
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 10722 5958 10774 6010
rect 10786 5958 10838 6010
rect 10850 5958 10902 6010
rect 10914 5958 10966 6010
rect 10978 5958 11030 6010
rect 2412 5856 2464 5908
rect 3056 5856 3108 5908
rect 7196 5856 7248 5908
rect 8116 5899 8168 5908
rect 8116 5865 8125 5899
rect 8125 5865 8159 5899
rect 8159 5865 8168 5899
rect 8116 5856 8168 5865
rect 9128 5856 9180 5908
rect 10416 5899 10468 5908
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 5080 5788 5132 5840
rect 1860 5720 1912 5772
rect 2412 5720 2464 5772
rect 1492 5652 1544 5704
rect 1952 5652 2004 5704
rect 2136 5584 2188 5636
rect 5816 5720 5868 5772
rect 5540 5652 5592 5704
rect 6460 5652 6512 5704
rect 5356 5584 5408 5636
rect 5908 5584 5960 5636
rect 5724 5516 5776 5568
rect 6828 5788 6880 5840
rect 7288 5720 7340 5772
rect 7840 5763 7892 5772
rect 7840 5729 7849 5763
rect 7849 5729 7883 5763
rect 7883 5729 7892 5763
rect 7840 5720 7892 5729
rect 8852 5788 8904 5840
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 8944 5720 8996 5772
rect 9588 5720 9640 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 8024 5584 8076 5636
rect 8576 5516 8628 5568
rect 9404 5516 9456 5568
rect 10416 5652 10468 5704
rect 10692 5720 10744 5772
rect 10692 5559 10744 5568
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 10062 5414 10114 5466
rect 10126 5414 10178 5466
rect 10190 5414 10242 5466
rect 10254 5414 10306 5466
rect 10318 5414 10370 5466
rect 2136 5355 2188 5364
rect 2136 5321 2145 5355
rect 2145 5321 2179 5355
rect 2179 5321 2188 5355
rect 2136 5312 2188 5321
rect 6920 5355 6972 5364
rect 6920 5321 6929 5355
rect 6929 5321 6963 5355
rect 6963 5321 6972 5355
rect 6920 5312 6972 5321
rect 7104 5312 7156 5364
rect 8484 5312 8536 5364
rect 9404 5355 9456 5364
rect 9404 5321 9413 5355
rect 9413 5321 9447 5355
rect 9447 5321 9456 5355
rect 9404 5312 9456 5321
rect 4068 5244 4120 5296
rect 5816 5287 5868 5296
rect 5816 5253 5825 5287
rect 5825 5253 5859 5287
rect 5859 5253 5868 5287
rect 5816 5244 5868 5253
rect 9588 5287 9640 5296
rect 9588 5253 9597 5287
rect 9597 5253 9631 5287
rect 9631 5253 9640 5287
rect 9588 5244 9640 5253
rect 1676 5176 1728 5228
rect 1492 5108 1544 5160
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 1400 5040 1452 5092
rect 1768 5083 1820 5092
rect 1768 5049 1777 5083
rect 1777 5049 1811 5083
rect 1811 5049 1820 5083
rect 1768 5040 1820 5049
rect 2044 5040 2096 5092
rect 3148 5108 3200 5160
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 5448 5151 5500 5160
rect 5448 5117 5457 5151
rect 5457 5117 5491 5151
rect 5491 5117 5500 5151
rect 5448 5108 5500 5117
rect 6000 5108 6052 5160
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 7288 5151 7340 5160
rect 7288 5117 7297 5151
rect 7297 5117 7331 5151
rect 7331 5117 7340 5151
rect 7288 5108 7340 5117
rect 9864 5219 9916 5228
rect 9864 5185 9873 5219
rect 9873 5185 9907 5219
rect 9907 5185 9916 5219
rect 9864 5176 9916 5185
rect 10692 5219 10744 5228
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 5356 4972 5408 5024
rect 6736 4972 6788 5024
rect 7196 4972 7248 5024
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 8668 4972 8720 5024
rect 9404 5108 9456 5160
rect 9772 5108 9824 5160
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 9496 4972 9548 5024
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 10722 4870 10774 4922
rect 10786 4870 10838 4922
rect 10850 4870 10902 4922
rect 10914 4870 10966 4922
rect 10978 4870 11030 4922
rect 1400 4768 1452 4820
rect 2228 4743 2280 4752
rect 2228 4709 2237 4743
rect 2237 4709 2271 4743
rect 2271 4709 2280 4743
rect 2228 4700 2280 4709
rect 1952 4675 2004 4684
rect 1952 4641 1961 4675
rect 1961 4641 1995 4675
rect 1995 4641 2004 4675
rect 1952 4632 2004 4641
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 3516 4768 3568 4820
rect 5448 4768 5500 4820
rect 7840 4811 7892 4820
rect 7840 4777 7849 4811
rect 7849 4777 7883 4811
rect 7883 4777 7892 4811
rect 7840 4768 7892 4777
rect 1860 4539 1912 4548
rect 1860 4505 1869 4539
rect 1869 4505 1903 4539
rect 1903 4505 1912 4539
rect 1860 4496 1912 4505
rect 1584 4428 1636 4480
rect 2964 4496 3016 4548
rect 4528 4700 4580 4752
rect 4896 4700 4948 4752
rect 8944 4811 8996 4820
rect 8944 4777 8953 4811
rect 8953 4777 8987 4811
rect 8987 4777 8996 4811
rect 8944 4768 8996 4777
rect 9680 4768 9732 4820
rect 4252 4632 4304 4684
rect 4712 4632 4764 4684
rect 6000 4632 6052 4684
rect 5448 4564 5500 4616
rect 7288 4675 7340 4684
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 8024 4675 8076 4684
rect 8024 4641 8033 4675
rect 8033 4641 8067 4675
rect 8067 4641 8076 4675
rect 8024 4632 8076 4641
rect 7840 4496 7892 4548
rect 8668 4743 8720 4752
rect 8668 4709 8677 4743
rect 8677 4709 8711 4743
rect 8711 4709 8720 4743
rect 8668 4700 8720 4709
rect 9404 4700 9456 4752
rect 9772 4743 9824 4752
rect 9772 4709 9781 4743
rect 9781 4709 9815 4743
rect 9815 4709 9824 4743
rect 9772 4700 9824 4709
rect 9956 4811 10008 4820
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 10416 4768 10468 4820
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 9220 4564 9272 4616
rect 9496 4564 9548 4616
rect 10600 4564 10652 4616
rect 6092 4428 6144 4480
rect 7564 4428 7616 4480
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 8484 4428 8536 4437
rect 8576 4428 8628 4480
rect 9772 4428 9824 4480
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 10062 4326 10114 4378
rect 10126 4326 10178 4378
rect 10190 4326 10242 4378
rect 10254 4326 10306 4378
rect 10318 4326 10370 4378
rect 1400 4267 1452 4276
rect 1400 4233 1409 4267
rect 1409 4233 1443 4267
rect 1443 4233 1452 4267
rect 1400 4224 1452 4233
rect 1952 4224 2004 4276
rect 3332 4224 3384 4276
rect 4528 4224 4580 4276
rect 5724 4224 5776 4276
rect 7196 4224 7248 4276
rect 2320 4156 2372 4208
rect 2504 4156 2556 4208
rect 1768 4088 1820 4140
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 2964 4156 3016 4208
rect 1952 4020 2004 4072
rect 1676 3952 1728 4004
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 4252 4156 4304 4208
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 4712 4020 4764 4029
rect 2044 3884 2096 3936
rect 2596 3884 2648 3936
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 5540 4131 5592 4140
rect 5540 4097 5549 4131
rect 5549 4097 5583 4131
rect 5583 4097 5592 4131
rect 8024 4156 8076 4208
rect 5540 4088 5592 4097
rect 4988 4063 5040 4072
rect 4988 4029 4997 4063
rect 4997 4029 5031 4063
rect 5031 4029 5040 4063
rect 4988 4020 5040 4029
rect 5080 4063 5132 4072
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 5356 4063 5408 4072
rect 5356 4029 5365 4063
rect 5365 4029 5399 4063
rect 5399 4029 5408 4063
rect 5356 4020 5408 4029
rect 5264 3952 5316 4004
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 5724 4020 5776 4029
rect 6000 4020 6052 4072
rect 4712 3884 4764 3893
rect 5448 3884 5500 3936
rect 6092 3927 6144 3936
rect 6092 3893 6101 3927
rect 6101 3893 6135 3927
rect 6135 3893 6144 3927
rect 6092 3884 6144 3893
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 7932 4020 7984 4072
rect 8484 4156 8536 4208
rect 9312 4224 9364 4276
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9772 4020 9824 4072
rect 8852 3884 8904 3936
rect 9680 3884 9732 3936
rect 10600 3884 10652 3936
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 10722 3782 10774 3834
rect 10786 3782 10838 3834
rect 10850 3782 10902 3834
rect 10914 3782 10966 3834
rect 10978 3782 11030 3834
rect 3516 3680 3568 3732
rect 2596 3655 2648 3664
rect 2596 3621 2605 3655
rect 2605 3621 2639 3655
rect 2639 3621 2648 3655
rect 2596 3612 2648 3621
rect 4252 3544 4304 3596
rect 6092 3680 6144 3732
rect 6184 3680 6236 3732
rect 8300 3680 8352 3732
rect 4712 3612 4764 3664
rect 5356 3612 5408 3664
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 2320 3476 2372 3528
rect 2412 3476 2464 3528
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 5540 3476 5592 3528
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 7564 3544 7616 3596
rect 8116 3612 8168 3664
rect 9128 3680 9180 3732
rect 6736 3476 6788 3528
rect 7288 3476 7340 3528
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 8852 3587 8904 3596
rect 8852 3553 8861 3587
rect 8861 3553 8895 3587
rect 8895 3553 8904 3587
rect 8852 3544 8904 3553
rect 9588 3544 9640 3596
rect 7748 3408 7800 3460
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 2504 3340 2556 3392
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 5724 3340 5776 3392
rect 5908 3383 5960 3392
rect 5908 3349 5917 3383
rect 5917 3349 5951 3383
rect 5951 3349 5960 3383
rect 5908 3340 5960 3349
rect 7288 3340 7340 3392
rect 7932 3340 7984 3392
rect 8024 3340 8076 3392
rect 8760 3340 8812 3392
rect 8852 3340 8904 3392
rect 9128 3340 9180 3392
rect 10508 3340 10560 3392
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 10062 3238 10114 3290
rect 10126 3238 10178 3290
rect 10190 3238 10242 3290
rect 10254 3238 10306 3290
rect 10318 3238 10370 3290
rect 3608 3136 3660 3188
rect 6184 3136 6236 3188
rect 7196 3179 7248 3188
rect 7196 3145 7205 3179
rect 7205 3145 7239 3179
rect 7239 3145 7248 3179
rect 7196 3136 7248 3145
rect 8300 3136 8352 3188
rect 8944 3136 8996 3188
rect 9680 3136 9732 3188
rect 10600 3136 10652 3188
rect 2228 3068 2280 3120
rect 1032 3043 1084 3052
rect 1032 3009 1041 3043
rect 1041 3009 1075 3043
rect 1075 3009 1084 3043
rect 1032 3000 1084 3009
rect 2504 2932 2556 2984
rect 5264 3068 5316 3120
rect 4436 3000 4488 3052
rect 4988 3000 5040 3052
rect 5356 3000 5408 3052
rect 2872 2932 2924 2984
rect 3056 2932 3108 2984
rect 5080 2932 5132 2984
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 7932 2932 7984 2984
rect 10508 2975 10560 2984
rect 10508 2941 10517 2975
rect 10517 2941 10551 2975
rect 10551 2941 10560 2975
rect 10508 2932 10560 2941
rect 2964 2864 3016 2916
rect 4620 2864 4672 2916
rect 4896 2864 4948 2916
rect 6644 2864 6696 2916
rect 7288 2864 7340 2916
rect 7748 2864 7800 2916
rect 7840 2907 7892 2916
rect 7840 2873 7849 2907
rect 7849 2873 7883 2907
rect 7883 2873 7892 2907
rect 7840 2864 7892 2873
rect 8760 2907 8812 2916
rect 8760 2873 8769 2907
rect 8769 2873 8803 2907
rect 8803 2873 8812 2907
rect 8760 2864 8812 2873
rect 1584 2796 1636 2848
rect 1676 2796 1728 2848
rect 2136 2796 2188 2848
rect 2872 2839 2924 2848
rect 2872 2805 2881 2839
rect 2881 2805 2915 2839
rect 2915 2805 2924 2839
rect 2872 2796 2924 2805
rect 3148 2796 3200 2848
rect 7012 2839 7064 2848
rect 7012 2805 7021 2839
rect 7021 2805 7055 2839
rect 7055 2805 7064 2839
rect 7012 2796 7064 2805
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 10722 2694 10774 2746
rect 10786 2694 10838 2746
rect 10850 2694 10902 2746
rect 10914 2694 10966 2746
rect 10978 2694 11030 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 2872 2592 2924 2644
rect 7840 2592 7892 2644
rect 8024 2635 8076 2644
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 8300 2592 8352 2644
rect 8944 2592 8996 2644
rect 2320 2524 2372 2576
rect 1400 2456 1452 2508
rect 2136 2456 2188 2508
rect 2504 2456 2556 2508
rect 2596 2456 2648 2508
rect 3240 2456 3292 2508
rect 3516 2524 3568 2576
rect 5172 2456 5224 2508
rect 9036 2524 9088 2576
rect 7104 2456 7156 2508
rect 9496 2524 9548 2576
rect 1492 2388 1544 2440
rect 2044 2388 2096 2440
rect 3332 2388 3384 2440
rect 1584 2320 1636 2372
rect 2780 2320 2832 2372
rect 3608 2320 3660 2372
rect 3424 2252 3476 2304
rect 4068 2252 4120 2304
rect 4160 2295 4212 2304
rect 4160 2261 4169 2295
rect 4169 2261 4203 2295
rect 4203 2261 4212 2295
rect 4160 2252 4212 2261
rect 6920 2252 6972 2304
rect 8300 2252 8352 2304
rect 8760 2252 8812 2304
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 10062 2150 10114 2202
rect 10126 2150 10178 2202
rect 10190 2150 10242 2202
rect 10254 2150 10306 2202
rect 10318 2150 10370 2202
rect 1584 2091 1636 2100
rect 1584 2057 1593 2091
rect 1593 2057 1627 2091
rect 1627 2057 1636 2091
rect 1584 2048 1636 2057
rect 3516 2048 3568 2100
rect 1492 1912 1544 1964
rect 1400 1887 1452 1896
rect 1400 1853 1409 1887
rect 1409 1853 1443 1887
rect 1443 1853 1452 1887
rect 1400 1844 1452 1853
rect 2964 1844 3016 1896
rect 3608 1980 3660 2032
rect 3332 1912 3384 1964
rect 5172 2091 5224 2100
rect 5172 2057 5181 2091
rect 5181 2057 5215 2091
rect 5215 2057 5224 2091
rect 5172 2048 5224 2057
rect 6920 2091 6972 2100
rect 6920 2057 6929 2091
rect 6929 2057 6963 2091
rect 6963 2057 6972 2091
rect 6920 2048 6972 2057
rect 7104 2091 7156 2100
rect 7104 2057 7113 2091
rect 7113 2057 7147 2091
rect 7147 2057 7156 2091
rect 7104 2048 7156 2057
rect 7012 1980 7064 2032
rect 8116 2048 8168 2100
rect 8760 2091 8812 2100
rect 8760 2057 8769 2091
rect 8769 2057 8803 2091
rect 8803 2057 8812 2091
rect 8760 2048 8812 2057
rect 9864 2048 9916 2100
rect 9496 1980 9548 2032
rect 7564 1955 7616 1964
rect 7564 1921 7573 1955
rect 7573 1921 7607 1955
rect 7607 1921 7616 1955
rect 7564 1912 7616 1921
rect 7748 1955 7800 1964
rect 7748 1921 7757 1955
rect 7757 1921 7791 1955
rect 7791 1921 7800 1955
rect 7748 1912 7800 1921
rect 3148 1776 3200 1828
rect 3608 1844 3660 1896
rect 3516 1819 3568 1828
rect 3516 1785 3525 1819
rect 3525 1785 3559 1819
rect 3559 1785 3568 1819
rect 3516 1776 3568 1785
rect 4068 1819 4120 1828
rect 4068 1785 4102 1819
rect 4102 1785 4120 1819
rect 4068 1776 4120 1785
rect 7196 1844 7248 1896
rect 7932 1887 7984 1896
rect 7932 1853 7941 1887
rect 7941 1853 7975 1887
rect 7975 1853 7984 1887
rect 7932 1844 7984 1853
rect 9128 1844 9180 1896
rect 4252 1776 4304 1828
rect 2596 1708 2648 1760
rect 3240 1708 3292 1760
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 10722 1606 10774 1658
rect 10786 1606 10838 1658
rect 10850 1606 10902 1658
rect 10914 1606 10966 1658
rect 10978 1606 11030 1658
rect 2320 1504 2372 1556
rect 2964 1504 3016 1556
rect 3056 1436 3108 1488
rect 2044 1368 2096 1420
rect 2320 1411 2372 1420
rect 2320 1377 2329 1411
rect 2329 1377 2363 1411
rect 2363 1377 2372 1411
rect 2320 1368 2372 1377
rect 3332 1436 3384 1488
rect 3516 1436 3568 1488
rect 3240 1368 3292 1420
rect 4160 1436 4212 1488
rect 1952 1300 2004 1352
rect 4252 1343 4304 1352
rect 4252 1309 4261 1343
rect 4261 1309 4295 1343
rect 4295 1309 4304 1343
rect 4252 1300 4304 1309
rect 4804 1300 4856 1352
rect 3516 1164 3568 1216
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 10062 1062 10114 1114
rect 10126 1062 10178 1114
rect 10190 1062 10242 1114
rect 10254 1062 10306 1114
rect 10318 1062 10370 1114
rect 3240 1003 3292 1012
rect 3240 969 3249 1003
rect 3249 969 3283 1003
rect 3283 969 3292 1003
rect 3240 960 3292 969
rect 3424 1003 3476 1012
rect 3424 969 3433 1003
rect 3433 969 3467 1003
rect 3467 969 3476 1003
rect 3424 960 3476 969
rect 2780 756 2832 808
rect 3056 688 3108 740
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
rect 10722 518 10774 570
rect 10786 518 10838 570
rect 10850 518 10902 570
rect 10914 518 10966 570
rect 10978 518 11030 570
<< metal2 >>
rect 570 43602 626 43900
rect 492 43574 626 43602
rect 386 41712 442 41721
rect 308 41670 386 41698
rect 204 41200 256 41206
rect 204 41142 256 41148
rect 112 37800 164 37806
rect 112 37742 164 37748
rect 20 32224 72 32230
rect 20 32166 72 32172
rect 32 30394 60 32166
rect 20 30388 72 30394
rect 20 30330 72 30336
rect 20 29504 72 29510
rect 20 29446 72 29452
rect 32 27538 60 29446
rect 124 28694 152 37742
rect 216 35193 244 41142
rect 308 38049 336 41670
rect 386 41647 442 41656
rect 388 40928 440 40934
rect 388 40870 440 40876
rect 400 38282 428 40870
rect 388 38276 440 38282
rect 388 38218 440 38224
rect 294 38040 350 38049
rect 294 37975 350 37984
rect 202 35184 258 35193
rect 202 35119 258 35128
rect 492 34542 520 43574
rect 570 43500 626 43574
rect 1122 43616 1178 43900
rect 1674 43602 1730 43900
rect 3330 43602 3386 43900
rect 1122 43500 1178 43560
rect 1504 43574 1730 43602
rect 1216 42152 1268 42158
rect 1216 42094 1268 42100
rect 1400 42152 1452 42158
rect 1400 42094 1452 42100
rect 572 42016 624 42022
rect 572 41958 624 41964
rect 584 40361 612 41958
rect 1124 41676 1176 41682
rect 1124 41618 1176 41624
rect 756 41608 808 41614
rect 1136 41585 1164 41618
rect 756 41550 808 41556
rect 1122 41576 1178 41585
rect 662 41440 718 41449
rect 662 41375 718 41384
rect 676 40934 704 41375
rect 664 40928 716 40934
rect 664 40870 716 40876
rect 664 40724 716 40730
rect 664 40666 716 40672
rect 570 40352 626 40361
rect 570 40287 626 40296
rect 572 39500 624 39506
rect 572 39442 624 39448
rect 584 35222 612 39442
rect 676 39098 704 40666
rect 664 39092 716 39098
rect 664 39034 716 39040
rect 768 38554 796 41550
rect 1122 41511 1178 41520
rect 1032 41472 1084 41478
rect 1032 41414 1084 41420
rect 1122 41440 1178 41449
rect 846 40624 902 40633
rect 846 40559 902 40568
rect 756 38548 808 38554
rect 756 38490 808 38496
rect 860 38010 888 40559
rect 940 40384 992 40390
rect 940 40326 992 40332
rect 952 39545 980 40326
rect 1044 40089 1072 41414
rect 1122 41375 1178 41384
rect 1030 40080 1086 40089
rect 1030 40015 1086 40024
rect 938 39536 994 39545
rect 938 39471 994 39480
rect 1136 39420 1164 41375
rect 952 39392 1164 39420
rect 848 38004 900 38010
rect 848 37946 900 37952
rect 754 36816 810 36825
rect 754 36751 810 36760
rect 662 36272 718 36281
rect 662 36207 718 36216
rect 572 35216 624 35222
rect 572 35158 624 35164
rect 204 34536 256 34542
rect 204 34478 256 34484
rect 480 34536 532 34542
rect 480 34478 532 34484
rect 112 28688 164 28694
rect 112 28630 164 28636
rect 112 28552 164 28558
rect 112 28494 164 28500
rect 124 28014 152 28494
rect 112 28008 164 28014
rect 112 27950 164 27956
rect 20 27532 72 27538
rect 20 27474 72 27480
rect 110 27024 166 27033
rect 110 26959 166 26968
rect 18 26072 74 26081
rect 18 26007 74 26016
rect 32 12782 60 26007
rect 124 24410 152 26959
rect 112 24404 164 24410
rect 112 24346 164 24352
rect 216 22710 244 34478
rect 388 32020 440 32026
rect 388 31962 440 31968
rect 294 31784 350 31793
rect 294 31719 350 31728
rect 400 31754 428 31962
rect 400 31726 612 31754
rect 308 29050 336 31719
rect 478 31512 534 31521
rect 478 31447 534 31456
rect 388 30388 440 30394
rect 388 30330 440 30336
rect 400 29170 428 30330
rect 492 29209 520 31447
rect 478 29200 534 29209
rect 388 29164 440 29170
rect 478 29135 534 29144
rect 388 29106 440 29112
rect 308 29022 520 29050
rect 386 28928 442 28937
rect 308 28886 386 28914
rect 204 22704 256 22710
rect 204 22646 256 22652
rect 110 22264 166 22273
rect 110 22199 166 22208
rect 124 17270 152 22199
rect 204 19440 256 19446
rect 308 19417 336 28886
rect 386 28863 442 28872
rect 388 28824 440 28830
rect 388 28766 440 28772
rect 400 25673 428 28766
rect 386 25664 442 25673
rect 386 25599 442 25608
rect 388 24608 440 24614
rect 388 24550 440 24556
rect 400 23497 428 24550
rect 386 23488 442 23497
rect 386 23423 442 23432
rect 388 23316 440 23322
rect 388 23258 440 23264
rect 204 19382 256 19388
rect 294 19408 350 19417
rect 112 17264 164 17270
rect 112 17206 164 17212
rect 216 14822 244 19382
rect 294 19343 350 19352
rect 400 17678 428 23258
rect 492 23186 520 29022
rect 480 23180 532 23186
rect 480 23122 532 23128
rect 584 19446 612 31726
rect 676 29073 704 36207
rect 662 29064 718 29073
rect 662 28999 718 29008
rect 662 28656 718 28665
rect 662 28591 718 28600
rect 676 24682 704 28591
rect 664 24676 716 24682
rect 664 24618 716 24624
rect 664 24404 716 24410
rect 664 24346 716 24352
rect 572 19440 624 19446
rect 572 19382 624 19388
rect 572 19304 624 19310
rect 572 19246 624 19252
rect 584 18902 612 19246
rect 572 18896 624 18902
rect 572 18838 624 18844
rect 676 18057 704 24346
rect 768 22642 796 36751
rect 952 34490 980 39392
rect 1124 39296 1176 39302
rect 1122 39264 1124 39273
rect 1176 39264 1178 39273
rect 1122 39199 1178 39208
rect 1032 38888 1084 38894
rect 1030 38856 1032 38865
rect 1084 38856 1086 38865
rect 1030 38791 1086 38800
rect 1124 38820 1176 38826
rect 1124 38762 1176 38768
rect 1136 38214 1164 38762
rect 1124 38208 1176 38214
rect 1124 38150 1176 38156
rect 1136 37942 1164 38150
rect 1124 37936 1176 37942
rect 1124 37878 1176 37884
rect 1136 37754 1164 37878
rect 1044 37726 1164 37754
rect 1044 37466 1072 37726
rect 1124 37664 1176 37670
rect 1124 37606 1176 37612
rect 1032 37460 1084 37466
rect 1032 37402 1084 37408
rect 1044 36718 1072 37402
rect 1136 37330 1164 37606
rect 1124 37324 1176 37330
rect 1124 37266 1176 37272
rect 1136 36922 1164 37266
rect 1124 36916 1176 36922
rect 1124 36858 1176 36864
rect 1032 36712 1084 36718
rect 1032 36654 1084 36660
rect 1044 36258 1072 36654
rect 1044 36242 1164 36258
rect 1044 36236 1176 36242
rect 1044 36230 1124 36236
rect 1124 36178 1176 36184
rect 1032 36032 1084 36038
rect 1032 35974 1084 35980
rect 1044 34592 1072 35974
rect 1122 35184 1178 35193
rect 1122 35119 1124 35128
rect 1176 35119 1178 35128
rect 1124 35090 1176 35096
rect 1124 34944 1176 34950
rect 1122 34912 1124 34921
rect 1176 34912 1178 34921
rect 1122 34847 1178 34856
rect 1044 34564 1164 34592
rect 952 34462 1072 34490
rect 940 34400 992 34406
rect 938 34368 940 34377
rect 992 34368 994 34377
rect 938 34303 994 34312
rect 1044 34134 1072 34462
rect 1032 34128 1084 34134
rect 1032 34070 1084 34076
rect 1136 33538 1164 34564
rect 1044 33510 1164 33538
rect 848 33312 900 33318
rect 848 33254 900 33260
rect 860 33114 888 33254
rect 848 33108 900 33114
rect 848 33050 900 33056
rect 860 31482 888 33050
rect 1044 32858 1072 33510
rect 1124 33448 1176 33454
rect 1124 33390 1176 33396
rect 1136 32978 1164 33390
rect 1124 32972 1176 32978
rect 1124 32914 1176 32920
rect 1044 32830 1164 32858
rect 1032 31884 1084 31890
rect 1032 31826 1084 31832
rect 940 31680 992 31686
rect 940 31622 992 31628
rect 848 31476 900 31482
rect 848 31418 900 31424
rect 860 30258 888 31418
rect 848 30252 900 30258
rect 848 30194 900 30200
rect 848 29028 900 29034
rect 848 28970 900 28976
rect 860 28626 888 28970
rect 848 28620 900 28626
rect 848 28562 900 28568
rect 860 28150 888 28562
rect 952 28490 980 31622
rect 1044 30938 1072 31826
rect 1136 31521 1164 32830
rect 1122 31512 1178 31521
rect 1122 31447 1178 31456
rect 1122 31376 1178 31385
rect 1122 31311 1178 31320
rect 1032 30932 1084 30938
rect 1032 30874 1084 30880
rect 1032 30728 1084 30734
rect 1032 30670 1084 30676
rect 1044 29617 1072 30670
rect 1030 29608 1086 29617
rect 1030 29543 1086 29552
rect 1030 29472 1086 29481
rect 1030 29407 1086 29416
rect 1044 29102 1072 29407
rect 1136 29306 1164 31311
rect 1228 30172 1256 42094
rect 1412 41750 1440 42094
rect 1400 41744 1452 41750
rect 1400 41686 1452 41692
rect 1308 40588 1360 40594
rect 1308 40530 1360 40536
rect 1320 40497 1348 40530
rect 1412 40526 1440 41686
rect 1504 41206 1532 43574
rect 1674 43500 1730 43574
rect 3068 43574 3386 43602
rect 1768 42900 1820 42906
rect 1768 42842 1820 42848
rect 2136 42900 2188 42906
rect 2136 42842 2188 42848
rect 1584 42560 1636 42566
rect 1584 42502 1636 42508
rect 1596 42158 1624 42502
rect 1584 42152 1636 42158
rect 1584 42094 1636 42100
rect 1584 41472 1636 41478
rect 1584 41414 1636 41420
rect 1780 41414 1808 42842
rect 2044 42696 2096 42702
rect 2044 42638 2096 42644
rect 1492 41200 1544 41206
rect 1492 41142 1544 41148
rect 1596 41070 1624 41414
rect 1780 41386 1900 41414
rect 1676 41200 1728 41206
rect 1780 41154 1808 41386
rect 1728 41148 1808 41154
rect 1676 41142 1808 41148
rect 1688 41126 1808 41142
rect 1584 41064 1636 41070
rect 1584 41006 1636 41012
rect 1492 40996 1544 41002
rect 1492 40938 1544 40944
rect 1768 40996 1820 41002
rect 1768 40938 1820 40944
rect 1504 40882 1532 40938
rect 1504 40854 1624 40882
rect 1492 40588 1544 40594
rect 1492 40530 1544 40536
rect 1400 40520 1452 40526
rect 1306 40488 1362 40497
rect 1400 40462 1452 40468
rect 1306 40423 1362 40432
rect 1308 40384 1360 40390
rect 1308 40326 1360 40332
rect 1320 39817 1348 40326
rect 1306 39808 1362 39817
rect 1306 39743 1362 39752
rect 1306 39536 1362 39545
rect 1412 39522 1440 40462
rect 1504 39681 1532 40530
rect 1596 39982 1624 40854
rect 1676 40588 1728 40594
rect 1676 40530 1728 40536
rect 1584 39976 1636 39982
rect 1584 39918 1636 39924
rect 1490 39672 1546 39681
rect 1596 39642 1624 39918
rect 1688 39642 1716 40530
rect 1490 39607 1546 39616
rect 1584 39636 1636 39642
rect 1584 39578 1636 39584
rect 1676 39636 1728 39642
rect 1676 39578 1728 39584
rect 1412 39494 1532 39522
rect 1306 39471 1362 39480
rect 1320 38962 1348 39471
rect 1504 39438 1532 39494
rect 1584 39500 1636 39506
rect 1584 39442 1636 39448
rect 1492 39432 1544 39438
rect 1492 39374 1544 39380
rect 1400 39024 1452 39030
rect 1400 38966 1452 38972
rect 1308 38956 1360 38962
rect 1308 38898 1360 38904
rect 1412 38654 1440 38966
rect 1504 38962 1532 39374
rect 1492 38956 1544 38962
rect 1492 38898 1544 38904
rect 1320 38626 1440 38654
rect 1320 38418 1348 38626
rect 1308 38412 1360 38418
rect 1308 38354 1360 38360
rect 1320 36650 1348 38354
rect 1504 38350 1532 38898
rect 1492 38344 1544 38350
rect 1492 38286 1544 38292
rect 1504 37330 1532 38286
rect 1596 37806 1624 39442
rect 1676 39364 1728 39370
rect 1676 39306 1728 39312
rect 1688 38758 1716 39306
rect 1676 38752 1728 38758
rect 1676 38694 1728 38700
rect 1688 38282 1716 38694
rect 1780 38554 1808 40938
rect 1872 40497 1900 41386
rect 2056 40934 2084 42638
rect 2148 42634 2176 42842
rect 3068 42770 3096 43574
rect 3330 43500 3386 43574
rect 3882 43500 3938 43900
rect 4434 43602 4490 43900
rect 4172 43574 4490 43602
rect 3896 42770 3924 43500
rect 2320 42764 2372 42770
rect 2320 42706 2372 42712
rect 3056 42764 3108 42770
rect 3056 42706 3108 42712
rect 3884 42764 3936 42770
rect 3884 42706 3936 42712
rect 2136 42628 2188 42634
rect 2136 42570 2188 42576
rect 2228 41744 2280 41750
rect 2228 41686 2280 41692
rect 2134 41168 2190 41177
rect 2134 41103 2190 41112
rect 2044 40928 2096 40934
rect 2044 40870 2096 40876
rect 1858 40488 1914 40497
rect 1858 40423 1914 40432
rect 1860 40384 1912 40390
rect 1860 40326 1912 40332
rect 1872 39982 1900 40326
rect 2056 40118 2084 40870
rect 2044 40112 2096 40118
rect 1964 40060 2044 40066
rect 1964 40054 2096 40060
rect 1964 40038 2084 40054
rect 1964 39982 1992 40038
rect 1860 39976 1912 39982
rect 1860 39918 1912 39924
rect 1952 39976 2004 39982
rect 1952 39918 2004 39924
rect 2044 39976 2096 39982
rect 2044 39918 2096 39924
rect 2056 39574 2084 39918
rect 1952 39568 2004 39574
rect 1952 39510 2004 39516
rect 2044 39568 2096 39574
rect 2044 39510 2096 39516
rect 1860 39296 1912 39302
rect 1860 39238 1912 39244
rect 1872 39098 1900 39238
rect 1860 39092 1912 39098
rect 1860 39034 1912 39040
rect 1872 38593 1900 39034
rect 1858 38584 1914 38593
rect 1768 38548 1820 38554
rect 1858 38519 1914 38528
rect 1768 38490 1820 38496
rect 1676 38276 1728 38282
rect 1676 38218 1728 38224
rect 1688 37890 1716 38218
rect 1780 37992 1808 38490
rect 1964 38418 1992 39510
rect 1952 38412 2004 38418
rect 1952 38354 2004 38360
rect 2148 38010 2176 41103
rect 2240 41070 2268 41686
rect 2228 41064 2280 41070
rect 2228 41006 2280 41012
rect 2226 40488 2282 40497
rect 2226 40423 2282 40432
rect 2136 38004 2188 38010
rect 1780 37964 1900 37992
rect 1688 37862 1808 37890
rect 1584 37800 1636 37806
rect 1584 37742 1636 37748
rect 1676 37664 1728 37670
rect 1676 37606 1728 37612
rect 1584 37392 1636 37398
rect 1584 37334 1636 37340
rect 1492 37324 1544 37330
rect 1492 37266 1544 37272
rect 1400 36780 1452 36786
rect 1504 36768 1532 37266
rect 1452 36740 1532 36768
rect 1400 36722 1452 36728
rect 1308 36644 1360 36650
rect 1308 36586 1360 36592
rect 1412 36310 1440 36722
rect 1400 36304 1452 36310
rect 1400 36246 1452 36252
rect 1412 35680 1440 36246
rect 1492 35692 1544 35698
rect 1412 35652 1492 35680
rect 1492 35634 1544 35640
rect 1596 35630 1624 37334
rect 1688 37330 1716 37606
rect 1676 37324 1728 37330
rect 1676 37266 1728 37272
rect 1780 37126 1808 37862
rect 1872 37738 1900 37964
rect 2136 37946 2188 37952
rect 1952 37800 2004 37806
rect 1952 37742 2004 37748
rect 1860 37732 1912 37738
rect 1860 37674 1912 37680
rect 1768 37120 1820 37126
rect 1768 37062 1820 37068
rect 1780 36718 1808 37062
rect 1768 36712 1820 36718
rect 1768 36654 1820 36660
rect 1780 36310 1808 36654
rect 1768 36304 1820 36310
rect 1768 36246 1820 36252
rect 1308 35624 1360 35630
rect 1308 35566 1360 35572
rect 1584 35624 1636 35630
rect 1584 35566 1636 35572
rect 1320 34746 1348 35566
rect 1768 35488 1820 35494
rect 1768 35430 1820 35436
rect 1780 35154 1808 35430
rect 1858 35184 1914 35193
rect 1584 35148 1636 35154
rect 1584 35090 1636 35096
rect 1768 35148 1820 35154
rect 1858 35119 1914 35128
rect 1768 35090 1820 35096
rect 1308 34740 1360 34746
rect 1308 34682 1360 34688
rect 1308 33992 1360 33998
rect 1308 33934 1360 33940
rect 1320 32552 1348 33934
rect 1596 33862 1624 35090
rect 1780 34524 1808 35090
rect 1872 35086 1900 35119
rect 1860 35080 1912 35086
rect 1860 35022 1912 35028
rect 1872 34626 1900 35022
rect 1964 34785 1992 37742
rect 2136 37732 2188 37738
rect 2136 37674 2188 37680
rect 1950 34776 2006 34785
rect 1950 34711 2006 34720
rect 1872 34598 2084 34626
rect 1780 34496 1900 34524
rect 1584 33856 1636 33862
rect 1584 33798 1636 33804
rect 1400 33448 1452 33454
rect 1400 33390 1452 33396
rect 1412 32910 1440 33390
rect 1492 32972 1544 32978
rect 1492 32914 1544 32920
rect 1584 32972 1636 32978
rect 1584 32914 1636 32920
rect 1400 32904 1452 32910
rect 1400 32846 1452 32852
rect 1320 32524 1440 32552
rect 1308 32292 1360 32298
rect 1308 32234 1360 32240
rect 1320 31278 1348 32234
rect 1412 31958 1440 32524
rect 1400 31952 1452 31958
rect 1400 31894 1452 31900
rect 1308 31272 1360 31278
rect 1504 31260 1532 32914
rect 1596 32230 1624 32914
rect 1768 32836 1820 32842
rect 1768 32778 1820 32784
rect 1584 32224 1636 32230
rect 1584 32166 1636 32172
rect 1780 31657 1808 32778
rect 1872 32450 1900 34496
rect 1952 34060 2004 34066
rect 1952 34002 2004 34008
rect 1964 33658 1992 34002
rect 1952 33652 2004 33658
rect 1952 33594 2004 33600
rect 1952 33516 2004 33522
rect 1952 33458 2004 33464
rect 1964 32570 1992 33458
rect 2056 33318 2084 34598
rect 2044 33312 2096 33318
rect 2044 33254 2096 33260
rect 2056 33153 2084 33254
rect 2042 33144 2098 33153
rect 2148 33130 2176 37674
rect 2240 37244 2268 40423
rect 2332 39982 2360 42706
rect 2504 42560 2556 42566
rect 2504 42502 2556 42508
rect 2320 39976 2372 39982
rect 2320 39918 2372 39924
rect 2516 39794 2544 42502
rect 3662 42460 3970 42469
rect 3662 42458 3668 42460
rect 3724 42458 3748 42460
rect 3804 42458 3828 42460
rect 3884 42458 3908 42460
rect 3964 42458 3970 42460
rect 3724 42406 3726 42458
rect 3906 42406 3908 42458
rect 3662 42404 3668 42406
rect 3724 42404 3748 42406
rect 3804 42404 3828 42406
rect 3884 42404 3908 42406
rect 3964 42404 3970 42406
rect 3662 42395 3970 42404
rect 2964 42220 3016 42226
rect 2964 42162 3016 42168
rect 2872 42152 2924 42158
rect 2872 42094 2924 42100
rect 2780 42016 2832 42022
rect 2780 41958 2832 41964
rect 2688 41200 2740 41206
rect 2688 41142 2740 41148
rect 2596 40452 2648 40458
rect 2596 40394 2648 40400
rect 2608 40186 2636 40394
rect 2596 40180 2648 40186
rect 2596 40122 2648 40128
rect 2700 39914 2728 41142
rect 2792 41070 2820 41958
rect 2780 41064 2832 41070
rect 2780 41006 2832 41012
rect 2792 40338 2820 41006
rect 2884 40458 2912 42094
rect 2872 40452 2924 40458
rect 2872 40394 2924 40400
rect 2792 40310 2912 40338
rect 2884 40050 2912 40310
rect 2976 40225 3004 42162
rect 3700 42152 3752 42158
rect 3700 42094 3752 42100
rect 3056 42016 3108 42022
rect 3056 41958 3108 41964
rect 3068 40905 3096 41958
rect 3712 41818 3740 42094
rect 4172 42090 4200 43574
rect 4434 43500 4490 43574
rect 4986 43500 5042 43900
rect 5538 43602 5594 43900
rect 5816 43648 5868 43654
rect 5538 43596 5816 43602
rect 5538 43590 5868 43596
rect 6090 43602 6146 43900
rect 5538 43574 5856 43590
rect 6090 43574 6224 43602
rect 5538 43500 5594 43574
rect 6090 43500 6146 43574
rect 4322 43004 4630 43013
rect 4322 43002 4328 43004
rect 4384 43002 4408 43004
rect 4464 43002 4488 43004
rect 4544 43002 4568 43004
rect 4624 43002 4630 43004
rect 4384 42950 4386 43002
rect 4566 42950 4568 43002
rect 4322 42948 4328 42950
rect 4384 42948 4408 42950
rect 4464 42948 4488 42950
rect 4544 42948 4568 42950
rect 4624 42948 4630 42950
rect 4322 42939 4630 42948
rect 4252 42696 4304 42702
rect 4252 42638 4304 42644
rect 4712 42696 4764 42702
rect 4712 42638 4764 42644
rect 4160 42084 4212 42090
rect 4160 42026 4212 42032
rect 3700 41812 3752 41818
rect 3700 41754 3752 41760
rect 3332 41744 3384 41750
rect 3332 41686 3384 41692
rect 3240 41676 3292 41682
rect 3240 41618 3292 41624
rect 3054 40896 3110 40905
rect 3054 40831 3110 40840
rect 3252 40730 3280 41618
rect 3240 40724 3292 40730
rect 3240 40666 3292 40672
rect 3240 40588 3292 40594
rect 3240 40530 3292 40536
rect 3056 40384 3108 40390
rect 3056 40326 3108 40332
rect 2962 40216 3018 40225
rect 3068 40186 3096 40326
rect 2962 40151 3018 40160
rect 3056 40180 3108 40186
rect 3056 40122 3108 40128
rect 3252 40118 3280 40530
rect 3240 40112 3292 40118
rect 3240 40054 3292 40060
rect 2872 40044 2924 40050
rect 2872 39986 2924 39992
rect 2688 39908 2740 39914
rect 2688 39850 2740 39856
rect 2964 39908 3016 39914
rect 2964 39850 3016 39856
rect 3056 39908 3108 39914
rect 3056 39850 3108 39856
rect 2516 39766 2820 39794
rect 2594 39672 2650 39681
rect 2594 39607 2650 39616
rect 2412 39500 2464 39506
rect 2412 39442 2464 39448
rect 2318 38584 2374 38593
rect 2424 38554 2452 39442
rect 2318 38519 2374 38528
rect 2412 38548 2464 38554
rect 2332 38486 2360 38519
rect 2412 38490 2464 38496
rect 2320 38480 2372 38486
rect 2320 38422 2372 38428
rect 2424 37942 2452 38490
rect 2504 38208 2556 38214
rect 2504 38150 2556 38156
rect 2516 38010 2544 38150
rect 2504 38004 2556 38010
rect 2504 37946 2556 37952
rect 2412 37936 2464 37942
rect 2412 37878 2464 37884
rect 2320 37800 2372 37806
rect 2320 37742 2372 37748
rect 2332 37369 2360 37742
rect 2504 37732 2556 37738
rect 2504 37674 2556 37680
rect 2318 37360 2374 37369
rect 2318 37295 2374 37304
rect 2240 37216 2452 37244
rect 2228 36168 2280 36174
rect 2228 36110 2280 36116
rect 2240 35086 2268 36110
rect 2228 35080 2280 35086
rect 2228 35022 2280 35028
rect 2320 35080 2372 35086
rect 2320 35022 2372 35028
rect 2240 33522 2268 35022
rect 2332 34746 2360 35022
rect 2320 34740 2372 34746
rect 2320 34682 2372 34688
rect 2320 33584 2372 33590
rect 2320 33526 2372 33532
rect 2228 33516 2280 33522
rect 2228 33458 2280 33464
rect 2148 33102 2268 33130
rect 2042 33079 2098 33088
rect 2044 32972 2096 32978
rect 2044 32914 2096 32920
rect 2136 32972 2188 32978
rect 2136 32914 2188 32920
rect 2056 32881 2084 32914
rect 2042 32872 2098 32881
rect 2042 32807 2098 32816
rect 2044 32768 2096 32774
rect 2044 32710 2096 32716
rect 1952 32564 2004 32570
rect 1952 32506 2004 32512
rect 1872 32422 1992 32450
rect 1964 31890 1992 32422
rect 1952 31884 2004 31890
rect 1952 31826 2004 31832
rect 1766 31648 1822 31657
rect 1766 31583 1822 31592
rect 2056 31464 2084 32710
rect 2148 31822 2176 32914
rect 2240 32042 2268 33102
rect 2332 32366 2360 33526
rect 2424 32774 2452 37216
rect 2516 35154 2544 37674
rect 2504 35148 2556 35154
rect 2504 35090 2556 35096
rect 2608 35034 2636 39607
rect 2792 39001 2820 39766
rect 2778 38992 2834 39001
rect 2778 38927 2834 38936
rect 2688 37256 2740 37262
rect 2688 37198 2740 37204
rect 2700 36378 2728 37198
rect 2688 36372 2740 36378
rect 2688 36314 2740 36320
rect 2516 35006 2636 35034
rect 2516 34134 2544 35006
rect 2596 34944 2648 34950
rect 2700 34921 2728 36314
rect 2792 36088 2820 38927
rect 2870 38448 2926 38457
rect 2870 38383 2926 38392
rect 2884 37330 2912 38383
rect 2976 38282 3004 39850
rect 3068 39030 3096 39850
rect 3148 39568 3200 39574
rect 3148 39510 3200 39516
rect 3056 39024 3108 39030
rect 3056 38966 3108 38972
rect 2964 38276 3016 38282
rect 2964 38218 3016 38224
rect 2962 38040 3018 38049
rect 2962 37975 2964 37984
rect 3016 37975 3018 37984
rect 3056 38004 3108 38010
rect 2964 37946 3016 37952
rect 3056 37946 3108 37952
rect 3068 37670 3096 37946
rect 3056 37664 3108 37670
rect 3056 37606 3108 37612
rect 2872 37324 2924 37330
rect 2872 37266 2924 37272
rect 2872 36644 2924 36650
rect 2872 36586 2924 36592
rect 2884 36417 2912 36586
rect 2870 36408 2926 36417
rect 2870 36343 2926 36352
rect 2884 36242 2912 36343
rect 2872 36236 2924 36242
rect 2872 36178 2924 36184
rect 2792 36060 2912 36088
rect 2778 36000 2834 36009
rect 2778 35935 2834 35944
rect 2792 35290 2820 35935
rect 2780 35284 2832 35290
rect 2780 35226 2832 35232
rect 2884 35154 2912 36060
rect 3068 35850 3096 37606
rect 3160 36242 3188 39510
rect 3252 38486 3280 40054
rect 3344 39982 3372 41686
rect 3712 41682 3740 41754
rect 3700 41676 3752 41682
rect 3700 41618 3752 41624
rect 3712 41562 3740 41618
rect 3528 41534 3740 41562
rect 3424 41472 3476 41478
rect 3424 41414 3476 41420
rect 3436 40050 3464 41414
rect 3528 41138 3556 41534
rect 3662 41372 3970 41381
rect 3662 41370 3668 41372
rect 3724 41370 3748 41372
rect 3804 41370 3828 41372
rect 3884 41370 3908 41372
rect 3964 41370 3970 41372
rect 3724 41318 3726 41370
rect 3906 41318 3908 41370
rect 3662 41316 3668 41318
rect 3724 41316 3748 41318
rect 3804 41316 3828 41318
rect 3884 41316 3908 41318
rect 3964 41316 3970 41318
rect 3662 41307 3970 41316
rect 3516 41132 3568 41138
rect 3516 41074 3568 41080
rect 4068 40996 4120 41002
rect 4068 40938 4120 40944
rect 3516 40520 3568 40526
rect 3516 40462 3568 40468
rect 3424 40044 3476 40050
rect 3424 39986 3476 39992
rect 3332 39976 3384 39982
rect 3528 39930 3556 40462
rect 3662 40284 3970 40293
rect 3662 40282 3668 40284
rect 3724 40282 3748 40284
rect 3804 40282 3828 40284
rect 3884 40282 3908 40284
rect 3964 40282 3970 40284
rect 3724 40230 3726 40282
rect 3906 40230 3908 40282
rect 3662 40228 3668 40230
rect 3724 40228 3748 40230
rect 3804 40228 3828 40230
rect 3884 40228 3908 40230
rect 3964 40228 3970 40230
rect 3662 40219 3970 40228
rect 4080 40186 4108 40938
rect 3700 40180 3752 40186
rect 3700 40122 3752 40128
rect 4068 40180 4120 40186
rect 4068 40122 4120 40128
rect 3332 39918 3384 39924
rect 3436 39902 3556 39930
rect 3606 39944 3662 39953
rect 3332 39296 3384 39302
rect 3332 39238 3384 39244
rect 3240 38480 3292 38486
rect 3240 38422 3292 38428
rect 3252 37856 3280 38422
rect 3344 38010 3372 39238
rect 3332 38004 3384 38010
rect 3332 37946 3384 37952
rect 3332 37868 3384 37874
rect 3252 37828 3332 37856
rect 3332 37810 3384 37816
rect 3238 37768 3294 37777
rect 3238 37703 3294 37712
rect 3252 36258 3280 37703
rect 3332 37460 3384 37466
rect 3332 37402 3384 37408
rect 3344 36786 3372 37402
rect 3436 37398 3464 39902
rect 3606 39879 3662 39888
rect 3620 39574 3648 39879
rect 3608 39568 3660 39574
rect 3608 39510 3660 39516
rect 3712 39386 3740 40122
rect 4160 39636 4212 39642
rect 4160 39578 4212 39584
rect 3528 39358 3740 39386
rect 4068 39432 4120 39438
rect 4068 39374 4120 39380
rect 3528 38570 3556 39358
rect 3662 39196 3970 39205
rect 3662 39194 3668 39196
rect 3724 39194 3748 39196
rect 3804 39194 3828 39196
rect 3884 39194 3908 39196
rect 3964 39194 3970 39196
rect 3724 39142 3726 39194
rect 3906 39142 3908 39194
rect 3662 39140 3668 39142
rect 3724 39140 3748 39142
rect 3804 39140 3828 39142
rect 3884 39140 3908 39142
rect 3964 39140 3970 39142
rect 3662 39131 3970 39140
rect 3700 39092 3752 39098
rect 3700 39034 3752 39040
rect 3528 38542 3648 38570
rect 3516 38412 3568 38418
rect 3516 38354 3568 38360
rect 3528 38214 3556 38354
rect 3620 38321 3648 38542
rect 3712 38486 3740 39034
rect 4080 38978 4108 39374
rect 3804 38950 4108 38978
rect 3804 38554 3832 38950
rect 3884 38888 3936 38894
rect 3936 38836 4108 38842
rect 3884 38830 4108 38836
rect 3896 38814 4108 38830
rect 4172 38826 4200 39578
rect 3792 38548 3844 38554
rect 3792 38490 3844 38496
rect 4080 38486 4108 38814
rect 4160 38820 4212 38826
rect 4160 38762 4212 38768
rect 3700 38480 3752 38486
rect 4068 38480 4120 38486
rect 3700 38422 3752 38428
rect 3790 38448 3846 38457
rect 4068 38422 4120 38428
rect 3790 38383 3792 38392
rect 3844 38383 3846 38392
rect 3792 38354 3844 38360
rect 3606 38312 3662 38321
rect 3606 38247 3662 38256
rect 3516 38208 3568 38214
rect 3516 38150 3568 38156
rect 3424 37392 3476 37398
rect 3424 37334 3476 37340
rect 3424 37256 3476 37262
rect 3424 37198 3476 37204
rect 3332 36780 3384 36786
rect 3332 36722 3384 36728
rect 3436 36310 3464 37198
rect 3528 36650 3556 38150
rect 3662 38108 3970 38117
rect 3662 38106 3668 38108
rect 3724 38106 3748 38108
rect 3804 38106 3828 38108
rect 3884 38106 3908 38108
rect 3964 38106 3970 38108
rect 3724 38054 3726 38106
rect 3906 38054 3908 38106
rect 3662 38052 3668 38054
rect 3724 38052 3748 38054
rect 3804 38052 3828 38054
rect 3884 38052 3908 38054
rect 3964 38052 3970 38054
rect 3662 38043 3970 38052
rect 3884 38004 3936 38010
rect 3884 37946 3936 37952
rect 3606 37904 3662 37913
rect 3606 37839 3662 37848
rect 3620 37806 3648 37839
rect 3608 37800 3660 37806
rect 3608 37742 3660 37748
rect 3896 37330 3924 37946
rect 3976 37936 4028 37942
rect 3976 37878 4028 37884
rect 3988 37330 4016 37878
rect 3884 37324 3936 37330
rect 3884 37266 3936 37272
rect 3976 37324 4028 37330
rect 3976 37266 4028 37272
rect 3662 37020 3970 37029
rect 3662 37018 3668 37020
rect 3724 37018 3748 37020
rect 3804 37018 3828 37020
rect 3884 37018 3908 37020
rect 3964 37018 3970 37020
rect 3724 36966 3726 37018
rect 3906 36966 3908 37018
rect 3662 36964 3668 36966
rect 3724 36964 3748 36966
rect 3804 36964 3828 36966
rect 3884 36964 3908 36966
rect 3964 36964 3970 36966
rect 3662 36955 3970 36964
rect 3790 36816 3846 36825
rect 3790 36751 3846 36760
rect 3516 36644 3568 36650
rect 3516 36586 3568 36592
rect 3804 36378 3832 36751
rect 4080 36718 4108 38422
rect 4160 38208 4212 38214
rect 4160 38150 4212 38156
rect 4172 37330 4200 38150
rect 4264 37806 4292 42638
rect 4344 42628 4396 42634
rect 4344 42570 4396 42576
rect 4356 42129 4384 42570
rect 4342 42120 4398 42129
rect 4342 42055 4398 42064
rect 4356 42022 4384 42055
rect 4344 42016 4396 42022
rect 4344 41958 4396 41964
rect 4322 41916 4630 41925
rect 4322 41914 4328 41916
rect 4384 41914 4408 41916
rect 4464 41914 4488 41916
rect 4544 41914 4568 41916
rect 4624 41914 4630 41916
rect 4384 41862 4386 41914
rect 4566 41862 4568 41914
rect 4322 41860 4328 41862
rect 4384 41860 4408 41862
rect 4464 41860 4488 41862
rect 4544 41860 4568 41862
rect 4624 41860 4630 41862
rect 4322 41851 4630 41860
rect 4724 41274 4752 42638
rect 4804 42628 4856 42634
rect 4804 42570 4856 42576
rect 4816 41478 4844 42570
rect 4896 42560 4948 42566
rect 4896 42502 4948 42508
rect 4908 42090 4936 42502
rect 4896 42084 4948 42090
rect 4896 42026 4948 42032
rect 4804 41472 4856 41478
rect 4804 41414 4856 41420
rect 4712 41268 4764 41274
rect 4712 41210 4764 41216
rect 4322 40828 4630 40837
rect 4322 40826 4328 40828
rect 4384 40826 4408 40828
rect 4464 40826 4488 40828
rect 4544 40826 4568 40828
rect 4624 40826 4630 40828
rect 4384 40774 4386 40826
rect 4566 40774 4568 40826
rect 4322 40772 4328 40774
rect 4384 40772 4408 40774
rect 4464 40772 4488 40774
rect 4544 40772 4568 40774
rect 4624 40772 4630 40774
rect 4322 40763 4630 40772
rect 4816 40526 4844 41414
rect 4896 41200 4948 41206
rect 4896 41142 4948 41148
rect 4908 40934 4936 41142
rect 5000 41070 5028 43500
rect 5632 42832 5684 42838
rect 5632 42774 5684 42780
rect 5356 42560 5408 42566
rect 5356 42502 5408 42508
rect 5080 42016 5132 42022
rect 5080 41958 5132 41964
rect 4988 41064 5040 41070
rect 4988 41006 5040 41012
rect 4896 40928 4948 40934
rect 4896 40870 4948 40876
rect 4988 40928 5040 40934
rect 4988 40870 5040 40876
rect 5000 40594 5028 40870
rect 5092 40730 5120 41958
rect 5368 41750 5396 42502
rect 5356 41744 5408 41750
rect 5356 41686 5408 41692
rect 5172 41676 5224 41682
rect 5172 41618 5224 41624
rect 5184 40934 5212 41618
rect 5172 40928 5224 40934
rect 5172 40870 5224 40876
rect 5264 40928 5316 40934
rect 5264 40870 5316 40876
rect 5356 40928 5408 40934
rect 5356 40870 5408 40876
rect 5080 40724 5132 40730
rect 5080 40666 5132 40672
rect 4988 40588 5040 40594
rect 4988 40530 5040 40536
rect 5080 40588 5132 40594
rect 5080 40530 5132 40536
rect 4528 40520 4580 40526
rect 4528 40462 4580 40468
rect 4804 40520 4856 40526
rect 4804 40462 4856 40468
rect 4896 40520 4948 40526
rect 5092 40474 5120 40530
rect 4896 40462 4948 40468
rect 4540 39846 4568 40462
rect 4620 40384 4672 40390
rect 4620 40326 4672 40332
rect 4632 40050 4660 40326
rect 4620 40044 4672 40050
rect 4620 39986 4672 39992
rect 4528 39840 4580 39846
rect 4528 39782 4580 39788
rect 4712 39840 4764 39846
rect 4712 39782 4764 39788
rect 4322 39740 4630 39749
rect 4322 39738 4328 39740
rect 4384 39738 4408 39740
rect 4464 39738 4488 39740
rect 4544 39738 4568 39740
rect 4624 39738 4630 39740
rect 4384 39686 4386 39738
rect 4566 39686 4568 39738
rect 4322 39684 4328 39686
rect 4384 39684 4408 39686
rect 4464 39684 4488 39686
rect 4544 39684 4568 39686
rect 4624 39684 4630 39686
rect 4322 39675 4630 39684
rect 4724 39642 4752 39782
rect 4712 39636 4764 39642
rect 4712 39578 4764 39584
rect 4322 38652 4630 38661
rect 4322 38650 4328 38652
rect 4384 38650 4408 38652
rect 4464 38650 4488 38652
rect 4544 38650 4568 38652
rect 4624 38650 4630 38652
rect 4384 38598 4386 38650
rect 4566 38598 4568 38650
rect 4322 38596 4328 38598
rect 4384 38596 4408 38598
rect 4464 38596 4488 38598
rect 4544 38596 4568 38598
rect 4624 38596 4630 38598
rect 4322 38587 4630 38596
rect 4724 38418 4752 39578
rect 4816 39438 4844 40462
rect 4908 40186 4936 40462
rect 5000 40446 5120 40474
rect 4896 40180 4948 40186
rect 4896 40122 4948 40128
rect 4908 39545 4936 40122
rect 4894 39536 4950 39545
rect 4894 39471 4950 39480
rect 4804 39432 4856 39438
rect 4804 39374 4856 39380
rect 4896 39432 4948 39438
rect 4896 39374 4948 39380
rect 4712 38412 4764 38418
rect 4712 38354 4764 38360
rect 4436 38276 4488 38282
rect 4436 38218 4488 38224
rect 4448 38185 4476 38218
rect 4434 38176 4490 38185
rect 4434 38111 4490 38120
rect 4724 37806 4752 38354
rect 4816 37874 4844 39374
rect 4804 37868 4856 37874
rect 4804 37810 4856 37816
rect 4252 37800 4304 37806
rect 4252 37742 4304 37748
rect 4712 37800 4764 37806
rect 4712 37742 4764 37748
rect 4252 37664 4304 37670
rect 4252 37606 4304 37612
rect 4712 37664 4764 37670
rect 4712 37606 4764 37612
rect 4160 37324 4212 37330
rect 4160 37266 4212 37272
rect 4264 36718 4292 37606
rect 4322 37564 4630 37573
rect 4322 37562 4328 37564
rect 4384 37562 4408 37564
rect 4464 37562 4488 37564
rect 4544 37562 4568 37564
rect 4624 37562 4630 37564
rect 4384 37510 4386 37562
rect 4566 37510 4568 37562
rect 4322 37508 4328 37510
rect 4384 37508 4408 37510
rect 4464 37508 4488 37510
rect 4544 37508 4568 37510
rect 4624 37508 4630 37510
rect 4322 37499 4630 37508
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 4068 36712 4120 36718
rect 4068 36654 4120 36660
rect 4252 36712 4304 36718
rect 4252 36654 4304 36660
rect 4632 36666 4660 37062
rect 4724 36922 4752 37606
rect 4816 37262 4844 37810
rect 4804 37256 4856 37262
rect 4804 37198 4856 37204
rect 4908 37074 4936 39374
rect 5000 38865 5028 40446
rect 5276 40089 5304 40870
rect 5262 40080 5318 40089
rect 5262 40015 5318 40024
rect 5172 39976 5224 39982
rect 5368 39964 5396 40870
rect 5644 40458 5672 42774
rect 6196 42770 6224 43574
rect 6642 43500 6698 43900
rect 7194 43500 7250 43900
rect 7746 43616 7802 43900
rect 7746 43500 7802 43560
rect 8298 43500 8354 43900
rect 8850 43500 8906 43900
rect 10508 43648 10560 43654
rect 10508 43590 10560 43596
rect 6656 42838 6684 43500
rect 6644 42832 6696 42838
rect 6644 42774 6696 42780
rect 7208 42770 7236 43500
rect 6184 42764 6236 42770
rect 6184 42706 6236 42712
rect 7196 42764 7248 42770
rect 7196 42706 7248 42712
rect 7012 42696 7064 42702
rect 7012 42638 7064 42644
rect 7748 42696 7800 42702
rect 7748 42638 7800 42644
rect 5816 42628 5868 42634
rect 5816 42570 5868 42576
rect 6184 42628 6236 42634
rect 6184 42570 6236 42576
rect 5828 42265 5856 42570
rect 5814 42256 5870 42265
rect 5814 42191 5870 42200
rect 6092 42220 6144 42226
rect 6092 42162 6144 42168
rect 6000 42152 6052 42158
rect 6000 42094 6052 42100
rect 5724 42084 5776 42090
rect 5724 42026 5776 42032
rect 5736 41682 5764 42026
rect 6012 41682 6040 42094
rect 5724 41676 5776 41682
rect 5724 41618 5776 41624
rect 6000 41676 6052 41682
rect 6000 41618 6052 41624
rect 5632 40452 5684 40458
rect 5632 40394 5684 40400
rect 5172 39918 5224 39924
rect 5276 39936 5396 39964
rect 5448 39976 5500 39982
rect 5080 39908 5132 39914
rect 5080 39850 5132 39856
rect 5092 39506 5120 39850
rect 5080 39500 5132 39506
rect 5080 39442 5132 39448
rect 5092 39098 5120 39442
rect 5080 39092 5132 39098
rect 5080 39034 5132 39040
rect 4986 38856 5042 38865
rect 4986 38791 5042 38800
rect 4816 37046 4936 37074
rect 4712 36916 4764 36922
rect 4712 36858 4764 36864
rect 3884 36576 3936 36582
rect 3884 36518 3936 36524
rect 3792 36372 3844 36378
rect 3792 36314 3844 36320
rect 3896 36310 3924 36518
rect 3424 36304 3476 36310
rect 3148 36236 3200 36242
rect 3252 36230 3372 36258
rect 3424 36246 3476 36252
rect 3884 36304 3936 36310
rect 3884 36246 3936 36252
rect 4080 36242 4108 36654
rect 4632 36638 4752 36666
rect 4322 36476 4630 36485
rect 4322 36474 4328 36476
rect 4384 36474 4408 36476
rect 4464 36474 4488 36476
rect 4544 36474 4568 36476
rect 4624 36474 4630 36476
rect 4384 36422 4386 36474
rect 4566 36422 4568 36474
rect 4322 36420 4328 36422
rect 4384 36420 4408 36422
rect 4464 36420 4488 36422
rect 4544 36420 4568 36422
rect 4624 36420 4630 36422
rect 4322 36411 4630 36420
rect 3148 36178 3200 36184
rect 3160 36038 3188 36178
rect 3148 36032 3200 36038
rect 3148 35974 3200 35980
rect 3068 35822 3280 35850
rect 3056 35556 3108 35562
rect 3056 35498 3108 35504
rect 3068 35154 3096 35498
rect 3148 35488 3200 35494
rect 3148 35430 3200 35436
rect 3160 35154 3188 35430
rect 2872 35148 2924 35154
rect 2872 35090 2924 35096
rect 3056 35148 3108 35154
rect 3056 35090 3108 35096
rect 3148 35148 3200 35154
rect 3148 35090 3200 35096
rect 2596 34886 2648 34892
rect 2686 34912 2742 34921
rect 2608 34542 2636 34886
rect 2686 34847 2742 34856
rect 2688 34740 2740 34746
rect 2688 34682 2740 34688
rect 2700 34649 2728 34682
rect 2884 34678 2912 35090
rect 2962 35048 3018 35057
rect 2962 34983 3018 34992
rect 2872 34672 2924 34678
rect 2686 34640 2742 34649
rect 2872 34614 2924 34620
rect 2976 34610 3004 34983
rect 2686 34575 2742 34584
rect 2964 34604 3016 34610
rect 2964 34546 3016 34552
rect 2596 34536 2648 34542
rect 2596 34478 2648 34484
rect 2780 34400 2832 34406
rect 2976 34354 3004 34546
rect 3056 34536 3108 34542
rect 3056 34478 3108 34484
rect 2780 34342 2832 34348
rect 2504 34128 2556 34134
rect 2504 34070 2556 34076
rect 2504 33856 2556 33862
rect 2504 33798 2556 33804
rect 2516 33318 2544 33798
rect 2504 33312 2556 33318
rect 2792 33289 2820 34342
rect 2884 34326 3004 34354
rect 2504 33254 2556 33260
rect 2778 33280 2834 33289
rect 2516 33017 2544 33254
rect 2778 33215 2834 33224
rect 2502 33008 2558 33017
rect 2502 32943 2558 32952
rect 2688 32972 2740 32978
rect 2688 32914 2740 32920
rect 2700 32774 2728 32914
rect 2412 32768 2464 32774
rect 2412 32710 2464 32716
rect 2504 32768 2556 32774
rect 2504 32710 2556 32716
rect 2688 32768 2740 32774
rect 2688 32710 2740 32716
rect 2412 32496 2464 32502
rect 2412 32438 2464 32444
rect 2320 32360 2372 32366
rect 2424 32337 2452 32438
rect 2320 32302 2372 32308
rect 2410 32328 2466 32337
rect 2516 32298 2544 32710
rect 2700 32366 2728 32710
rect 2884 32586 2912 34326
rect 2964 33856 3016 33862
rect 3068 33844 3096 34478
rect 3148 34468 3200 34474
rect 3148 34410 3200 34416
rect 3160 33998 3188 34410
rect 3148 33992 3200 33998
rect 3148 33934 3200 33940
rect 3016 33816 3096 33844
rect 2964 33798 3016 33804
rect 3056 33448 3108 33454
rect 3056 33390 3108 33396
rect 2964 33312 3016 33318
rect 2964 33254 3016 33260
rect 2976 32842 3004 33254
rect 3068 32978 3096 33390
rect 3056 32972 3108 32978
rect 3056 32914 3108 32920
rect 2964 32836 3016 32842
rect 2964 32778 3016 32784
rect 2792 32558 2912 32586
rect 2688 32360 2740 32366
rect 2688 32302 2740 32308
rect 2410 32263 2466 32272
rect 2504 32292 2556 32298
rect 2424 32178 2452 32263
rect 2504 32234 2556 32240
rect 2688 32224 2740 32230
rect 2424 32150 2636 32178
rect 2688 32166 2740 32172
rect 2240 32014 2452 32042
rect 2318 31920 2374 31929
rect 2228 31884 2280 31890
rect 2318 31855 2374 31864
rect 2228 31826 2280 31832
rect 2136 31816 2188 31822
rect 2136 31758 2188 31764
rect 1872 31436 2084 31464
rect 1584 31272 1636 31278
rect 1504 31232 1584 31260
rect 1308 31214 1360 31220
rect 1584 31214 1636 31220
rect 1400 31136 1452 31142
rect 1400 31078 1452 31084
rect 1308 30864 1360 30870
rect 1308 30806 1360 30812
rect 1320 30326 1348 30806
rect 1412 30598 1440 31078
rect 1492 30796 1544 30802
rect 1492 30738 1544 30744
rect 1400 30592 1452 30598
rect 1400 30534 1452 30540
rect 1504 30394 1532 30738
rect 1596 30666 1624 31214
rect 1768 31136 1820 31142
rect 1766 31104 1768 31113
rect 1820 31104 1822 31113
rect 1766 31039 1822 31048
rect 1584 30660 1636 30666
rect 1584 30602 1636 30608
rect 1676 30592 1728 30598
rect 1676 30534 1728 30540
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 1492 30388 1544 30394
rect 1492 30330 1544 30336
rect 1308 30320 1360 30326
rect 1308 30262 1360 30268
rect 1228 30144 1440 30172
rect 1216 29640 1268 29646
rect 1214 29608 1216 29617
rect 1268 29608 1270 29617
rect 1214 29543 1270 29552
rect 1412 29322 1440 30144
rect 1124 29300 1176 29306
rect 1124 29242 1176 29248
rect 1320 29294 1440 29322
rect 1320 29186 1348 29294
rect 1504 29238 1532 30330
rect 1584 30116 1636 30122
rect 1584 30058 1636 30064
rect 1596 29560 1624 30058
rect 1688 29714 1716 30534
rect 1780 29714 1808 30534
rect 1872 29714 1900 31436
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 1964 30938 1992 31282
rect 2240 31278 2268 31826
rect 2332 31328 2360 31855
rect 2424 31686 2452 32014
rect 2412 31680 2464 31686
rect 2412 31622 2464 31628
rect 2332 31300 2452 31328
rect 2228 31272 2280 31278
rect 2228 31214 2280 31220
rect 2044 31136 2096 31142
rect 2044 31078 2096 31084
rect 1952 30932 2004 30938
rect 1952 30874 2004 30880
rect 2056 30802 2084 31078
rect 1952 30796 2004 30802
rect 1952 30738 2004 30744
rect 2044 30796 2096 30802
rect 2096 30756 2176 30784
rect 2044 30738 2096 30744
rect 1676 29708 1728 29714
rect 1676 29650 1728 29656
rect 1768 29708 1820 29714
rect 1768 29650 1820 29656
rect 1860 29708 1912 29714
rect 1860 29650 1912 29656
rect 1676 29572 1728 29578
rect 1596 29532 1676 29560
rect 1676 29514 1728 29520
rect 1228 29158 1348 29186
rect 1400 29232 1452 29238
rect 1400 29174 1452 29180
rect 1492 29232 1544 29238
rect 1492 29174 1544 29180
rect 1032 29096 1084 29102
rect 1032 29038 1084 29044
rect 1124 29096 1176 29102
rect 1124 29038 1176 29044
rect 1032 28960 1084 28966
rect 1032 28902 1084 28908
rect 940 28484 992 28490
rect 940 28426 992 28432
rect 848 28144 900 28150
rect 952 28121 980 28426
rect 848 28086 900 28092
rect 938 28112 994 28121
rect 938 28047 994 28056
rect 938 27976 994 27985
rect 938 27911 994 27920
rect 848 27872 900 27878
rect 846 27840 848 27849
rect 900 27840 902 27849
rect 846 27775 902 27784
rect 952 27402 980 27911
rect 940 27396 992 27402
rect 940 27338 992 27344
rect 848 27328 900 27334
rect 1044 27282 1072 28902
rect 1136 28121 1164 29038
rect 1228 29034 1256 29158
rect 1216 29028 1268 29034
rect 1216 28970 1268 28976
rect 1122 28112 1178 28121
rect 1122 28047 1178 28056
rect 1124 28008 1176 28014
rect 1124 27950 1176 27956
rect 1136 27334 1164 27950
rect 1228 27577 1256 28970
rect 1308 28960 1360 28966
rect 1308 28902 1360 28908
rect 1320 28801 1348 28902
rect 1306 28792 1362 28801
rect 1306 28727 1362 28736
rect 1308 28688 1360 28694
rect 1308 28630 1360 28636
rect 1320 28529 1348 28630
rect 1306 28520 1362 28529
rect 1306 28455 1362 28464
rect 1308 28416 1360 28422
rect 1308 28358 1360 28364
rect 1214 27568 1270 27577
rect 1214 27503 1270 27512
rect 848 27270 900 27276
rect 860 26994 888 27270
rect 952 27254 1072 27282
rect 1124 27328 1176 27334
rect 1124 27270 1176 27276
rect 1216 27328 1268 27334
rect 1216 27270 1268 27276
rect 848 26988 900 26994
rect 848 26930 900 26936
rect 848 26444 900 26450
rect 848 26386 900 26392
rect 860 25770 888 26386
rect 848 25764 900 25770
rect 848 25706 900 25712
rect 860 25226 888 25706
rect 952 25480 980 27254
rect 1122 27160 1178 27169
rect 1228 27130 1256 27270
rect 1122 27095 1178 27104
rect 1216 27124 1268 27130
rect 1030 26888 1086 26897
rect 1030 26823 1086 26832
rect 1044 26790 1072 26823
rect 1032 26784 1084 26790
rect 1032 26726 1084 26732
rect 1044 26450 1072 26726
rect 1136 26586 1164 27095
rect 1216 27066 1268 27072
rect 1320 26926 1348 28358
rect 1412 28014 1440 29174
rect 1504 28082 1532 29174
rect 1584 28484 1636 28490
rect 1584 28426 1636 28432
rect 1492 28076 1544 28082
rect 1492 28018 1544 28024
rect 1400 28008 1452 28014
rect 1400 27950 1452 27956
rect 1398 27840 1454 27849
rect 1398 27775 1454 27784
rect 1412 27674 1440 27775
rect 1400 27668 1452 27674
rect 1400 27610 1452 27616
rect 1398 27568 1454 27577
rect 1398 27503 1454 27512
rect 1308 26920 1360 26926
rect 1308 26862 1360 26868
rect 1216 26784 1268 26790
rect 1216 26726 1268 26732
rect 1124 26580 1176 26586
rect 1124 26522 1176 26528
rect 1032 26444 1084 26450
rect 1032 26386 1084 26392
rect 1044 25809 1072 26386
rect 1124 26240 1176 26246
rect 1124 26182 1176 26188
rect 1030 25800 1086 25809
rect 1030 25735 1086 25744
rect 952 25452 1072 25480
rect 940 25356 992 25362
rect 940 25298 992 25304
rect 848 25220 900 25226
rect 848 25162 900 25168
rect 848 24132 900 24138
rect 848 24074 900 24080
rect 860 23322 888 24074
rect 952 23905 980 25298
rect 1044 24410 1072 25452
rect 1136 25294 1164 26182
rect 1228 25378 1256 26726
rect 1412 26450 1440 27503
rect 1400 26444 1452 26450
rect 1320 26404 1400 26432
rect 1320 25838 1348 26404
rect 1400 26386 1452 26392
rect 1504 26330 1532 28018
rect 1596 27946 1624 28426
rect 1584 27940 1636 27946
rect 1584 27882 1636 27888
rect 1584 27464 1636 27470
rect 1582 27432 1584 27441
rect 1688 27452 1716 29514
rect 1780 29170 1808 29650
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1780 28558 1808 29106
rect 1768 28552 1820 28558
rect 1768 28494 1820 28500
rect 1872 28218 1900 29650
rect 1964 29306 1992 30738
rect 2042 30560 2098 30569
rect 2042 30495 2098 30504
rect 2056 30190 2084 30495
rect 2044 30184 2096 30190
rect 2044 30126 2096 30132
rect 1952 29300 2004 29306
rect 1952 29242 2004 29248
rect 1950 28792 2006 28801
rect 1950 28727 1952 28736
rect 2004 28727 2006 28736
rect 1952 28698 2004 28704
rect 1952 28620 2004 28626
rect 1952 28562 2004 28568
rect 1860 28212 1912 28218
rect 1780 28172 1860 28200
rect 1780 27606 1808 28172
rect 1860 28154 1912 28160
rect 1860 28008 1912 28014
rect 1860 27950 1912 27956
rect 1768 27600 1820 27606
rect 1768 27542 1820 27548
rect 1872 27538 1900 27950
rect 1964 27674 1992 28562
rect 2056 27690 2084 30126
rect 2148 29730 2176 30756
rect 2240 30734 2268 31214
rect 2320 31204 2372 31210
rect 2320 31146 2372 31152
rect 2332 30977 2360 31146
rect 2318 30968 2374 30977
rect 2318 30903 2374 30912
rect 2228 30728 2280 30734
rect 2228 30670 2280 30676
rect 2226 30288 2282 30297
rect 2226 30223 2282 30232
rect 2240 30190 2268 30223
rect 2228 30184 2280 30190
rect 2332 30161 2360 30903
rect 2228 30126 2280 30132
rect 2318 30152 2374 30161
rect 2318 30087 2374 30096
rect 2228 30048 2280 30054
rect 2228 29990 2280 29996
rect 2240 29850 2268 29990
rect 2228 29844 2280 29850
rect 2228 29786 2280 29792
rect 2148 29714 2268 29730
rect 2148 29708 2280 29714
rect 2148 29702 2228 29708
rect 2228 29650 2280 29656
rect 2136 29640 2188 29646
rect 2136 29582 2188 29588
rect 2148 29345 2176 29582
rect 2134 29336 2190 29345
rect 2134 29271 2190 29280
rect 2136 29232 2188 29238
rect 2136 29174 2188 29180
rect 2148 28626 2176 29174
rect 2240 28966 2268 29650
rect 2332 29646 2360 30087
rect 2320 29640 2372 29646
rect 2320 29582 2372 29588
rect 2320 29504 2372 29510
rect 2320 29446 2372 29452
rect 2228 28960 2280 28966
rect 2228 28902 2280 28908
rect 2240 28762 2268 28902
rect 2228 28756 2280 28762
rect 2228 28698 2280 28704
rect 2136 28620 2188 28626
rect 2136 28562 2188 28568
rect 2136 28484 2188 28490
rect 2136 28426 2188 28432
rect 2148 27985 2176 28426
rect 2228 28416 2280 28422
rect 2228 28358 2280 28364
rect 2240 28082 2268 28358
rect 2228 28076 2280 28082
rect 2228 28018 2280 28024
rect 2134 27976 2190 27985
rect 2134 27911 2190 27920
rect 2136 27872 2188 27878
rect 2188 27832 2268 27860
rect 2136 27814 2188 27820
rect 2134 27704 2190 27713
rect 1952 27668 2004 27674
rect 2056 27662 2134 27690
rect 2134 27639 2190 27648
rect 1952 27610 2004 27616
rect 1950 27568 2006 27577
rect 1860 27532 1912 27538
rect 1950 27503 2006 27512
rect 2044 27532 2096 27538
rect 1860 27474 1912 27480
rect 1768 27464 1820 27470
rect 1636 27432 1638 27441
rect 1688 27424 1768 27452
rect 1768 27406 1820 27412
rect 1582 27367 1638 27376
rect 1676 27328 1728 27334
rect 1582 27296 1638 27305
rect 1676 27270 1728 27276
rect 1582 27231 1638 27240
rect 1596 26625 1624 27231
rect 1582 26616 1638 26625
rect 1688 26586 1716 27270
rect 1780 26874 1808 27406
rect 1872 26994 1900 27474
rect 1860 26988 1912 26994
rect 1860 26930 1912 26936
rect 1780 26858 1900 26874
rect 1768 26852 1900 26858
rect 1820 26846 1900 26852
rect 1768 26794 1820 26800
rect 1582 26551 1638 26560
rect 1676 26580 1728 26586
rect 1676 26522 1728 26528
rect 1674 26480 1730 26489
rect 1730 26424 1808 26432
rect 1674 26415 1676 26424
rect 1728 26404 1808 26424
rect 1676 26386 1728 26392
rect 1400 26308 1452 26314
rect 1504 26302 1624 26330
rect 1400 26250 1452 26256
rect 1412 26042 1440 26250
rect 1492 26240 1544 26246
rect 1492 26182 1544 26188
rect 1400 26036 1452 26042
rect 1400 25978 1452 25984
rect 1398 25936 1454 25945
rect 1504 25906 1532 26182
rect 1596 25974 1624 26302
rect 1674 26208 1730 26217
rect 1674 26143 1730 26152
rect 1584 25968 1636 25974
rect 1584 25910 1636 25916
rect 1398 25871 1400 25880
rect 1452 25871 1454 25880
rect 1492 25900 1544 25906
rect 1400 25842 1452 25848
rect 1492 25842 1544 25848
rect 1308 25832 1360 25838
rect 1308 25774 1360 25780
rect 1228 25350 1348 25378
rect 1504 25362 1532 25842
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1596 25430 1624 25638
rect 1584 25424 1636 25430
rect 1584 25366 1636 25372
rect 1124 25288 1176 25294
rect 1124 25230 1176 25236
rect 1216 25288 1268 25294
rect 1216 25230 1268 25236
rect 1032 24404 1084 24410
rect 1032 24346 1084 24352
rect 1030 24304 1086 24313
rect 1030 24239 1086 24248
rect 938 23896 994 23905
rect 938 23831 994 23840
rect 848 23316 900 23322
rect 848 23258 900 23264
rect 846 23216 902 23225
rect 846 23151 902 23160
rect 860 22778 888 23151
rect 940 22976 992 22982
rect 938 22944 940 22953
rect 992 22944 994 22953
rect 938 22879 994 22888
rect 848 22772 900 22778
rect 848 22714 900 22720
rect 756 22636 808 22642
rect 756 22578 808 22584
rect 940 22568 992 22574
rect 940 22510 992 22516
rect 952 22409 980 22510
rect 938 22400 994 22409
rect 938 22335 994 22344
rect 756 22024 808 22030
rect 756 21966 808 21972
rect 662 18048 718 18057
rect 662 17983 718 17992
rect 388 17672 440 17678
rect 388 17614 440 17620
rect 294 17504 350 17513
rect 294 17439 350 17448
rect 308 16674 336 17439
rect 570 17096 626 17105
rect 570 17031 626 17040
rect 664 17060 716 17066
rect 386 16688 442 16697
rect 308 16646 386 16674
rect 386 16623 442 16632
rect 388 16584 440 16590
rect 388 16526 440 16532
rect 204 14816 256 14822
rect 204 14758 256 14764
rect 20 12776 72 12782
rect 20 12718 72 12724
rect 400 5273 428 16526
rect 584 12073 612 17031
rect 664 17002 716 17008
rect 570 12064 626 12073
rect 570 11999 626 12008
rect 676 5545 704 17002
rect 768 12345 796 21966
rect 848 19236 900 19242
rect 848 19178 900 19184
rect 860 18630 888 19178
rect 952 18970 980 22335
rect 1044 21690 1072 24239
rect 1228 23644 1256 25230
rect 1320 24954 1348 25350
rect 1492 25356 1544 25362
rect 1492 25298 1544 25304
rect 1400 25152 1452 25158
rect 1400 25094 1452 25100
rect 1308 24948 1360 24954
rect 1308 24890 1360 24896
rect 1412 24818 1440 25094
rect 1504 24818 1532 25298
rect 1584 25220 1636 25226
rect 1584 25162 1636 25168
rect 1400 24812 1452 24818
rect 1320 24772 1400 24800
rect 1320 24274 1348 24772
rect 1400 24754 1452 24760
rect 1492 24812 1544 24818
rect 1492 24754 1544 24760
rect 1398 24712 1454 24721
rect 1398 24647 1454 24656
rect 1492 24676 1544 24682
rect 1412 24342 1440 24647
rect 1492 24618 1544 24624
rect 1400 24336 1452 24342
rect 1400 24278 1452 24284
rect 1308 24268 1360 24274
rect 1308 24210 1360 24216
rect 1306 24032 1362 24041
rect 1306 23967 1362 23976
rect 1136 23616 1256 23644
rect 1032 21684 1084 21690
rect 1032 21626 1084 21632
rect 1136 20641 1164 23616
rect 1320 23322 1348 23967
rect 1400 23588 1452 23594
rect 1400 23530 1452 23536
rect 1412 23497 1440 23530
rect 1398 23488 1454 23497
rect 1398 23423 1454 23432
rect 1308 23316 1360 23322
rect 1308 23258 1360 23264
rect 1400 23316 1452 23322
rect 1400 23258 1452 23264
rect 1216 23180 1268 23186
rect 1216 23122 1268 23128
rect 1228 23089 1256 23122
rect 1214 23080 1270 23089
rect 1214 23015 1270 23024
rect 1308 22704 1360 22710
rect 1308 22646 1360 22652
rect 1320 22545 1348 22646
rect 1306 22536 1362 22545
rect 1216 22500 1268 22506
rect 1306 22471 1362 22480
rect 1216 22442 1268 22448
rect 1122 20632 1178 20641
rect 1122 20567 1178 20576
rect 1228 20330 1256 22442
rect 1412 21593 1440 23258
rect 1398 21584 1454 21593
rect 1398 21519 1454 21528
rect 1308 21480 1360 21486
rect 1308 21422 1360 21428
rect 1320 21146 1348 21422
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1308 21140 1360 21146
rect 1308 21082 1360 21088
rect 1412 21010 1440 21286
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1216 20324 1268 20330
rect 1136 20284 1216 20312
rect 1032 19712 1084 19718
rect 1032 19654 1084 19660
rect 940 18964 992 18970
rect 940 18906 992 18912
rect 848 18624 900 18630
rect 848 18566 900 18572
rect 860 17814 888 18566
rect 848 17808 900 17814
rect 848 17750 900 17756
rect 848 17672 900 17678
rect 848 17614 900 17620
rect 860 15881 888 17614
rect 938 17232 994 17241
rect 938 17167 994 17176
rect 952 16250 980 17167
rect 940 16244 992 16250
rect 940 16186 992 16192
rect 938 16144 994 16153
rect 938 16079 994 16088
rect 846 15872 902 15881
rect 846 15807 902 15816
rect 754 12336 810 12345
rect 754 12271 810 12280
rect 952 8974 980 16079
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 662 5536 718 5545
rect 662 5471 718 5480
rect 386 5264 442 5273
rect 386 5199 442 5208
rect 386 4992 442 5001
rect 386 4927 442 4936
rect 400 4457 428 4927
rect 386 4448 442 4457
rect 386 4383 442 4392
rect 1044 3058 1072 19654
rect 1136 19446 1164 20284
rect 1216 20266 1268 20272
rect 1216 19848 1268 19854
rect 1216 19790 1268 19796
rect 1124 19440 1176 19446
rect 1124 19382 1176 19388
rect 1124 19304 1176 19310
rect 1124 19246 1176 19252
rect 1136 18290 1164 19246
rect 1124 18284 1176 18290
rect 1124 18226 1176 18232
rect 1124 17536 1176 17542
rect 1124 17478 1176 17484
rect 1136 16969 1164 17478
rect 1122 16960 1178 16969
rect 1122 16895 1178 16904
rect 1122 16824 1178 16833
rect 1122 16759 1178 16768
rect 1136 13870 1164 16759
rect 1124 13864 1176 13870
rect 1124 13806 1176 13812
rect 1136 10606 1164 13806
rect 1228 12617 1256 19790
rect 1320 19310 1348 20703
rect 1398 20496 1454 20505
rect 1398 20431 1400 20440
rect 1452 20431 1454 20440
rect 1400 20402 1452 20408
rect 1504 19378 1532 24618
rect 1596 23322 1624 25162
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1688 23202 1716 26143
rect 1780 25702 1808 26404
rect 1768 25696 1820 25702
rect 1768 25638 1820 25644
rect 1780 24449 1808 25638
rect 1766 24440 1822 24449
rect 1766 24375 1822 24384
rect 1768 24268 1820 24274
rect 1768 24210 1820 24216
rect 1780 23730 1808 24210
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1596 23174 1716 23202
rect 1596 21570 1624 23174
rect 1872 23118 1900 26846
rect 1964 26450 1992 27503
rect 2044 27474 2096 27480
rect 2056 26586 2084 27474
rect 2044 26580 2096 26586
rect 2044 26522 2096 26528
rect 1952 26444 2004 26450
rect 1952 26386 2004 26392
rect 2044 26444 2096 26450
rect 2044 26386 2096 26392
rect 1952 26240 2004 26246
rect 1952 26182 2004 26188
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 1768 22976 1820 22982
rect 1768 22918 1820 22924
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 1688 22681 1716 22714
rect 1674 22672 1730 22681
rect 1674 22607 1730 22616
rect 1780 22574 1808 22918
rect 1676 22568 1728 22574
rect 1676 22510 1728 22516
rect 1768 22568 1820 22574
rect 1768 22510 1820 22516
rect 1688 21690 1716 22510
rect 1780 22098 1808 22510
rect 1872 22234 1900 22918
rect 1860 22228 1912 22234
rect 1860 22170 1912 22176
rect 1768 22092 1820 22098
rect 1768 22034 1820 22040
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 1676 21684 1728 21690
rect 1676 21626 1728 21632
rect 1596 21542 1808 21570
rect 1584 21480 1636 21486
rect 1584 21422 1636 21428
rect 1596 20806 1624 21422
rect 1676 21004 1728 21010
rect 1676 20946 1728 20952
rect 1584 20800 1636 20806
rect 1584 20742 1636 20748
rect 1596 20466 1624 20742
rect 1688 20534 1716 20946
rect 1676 20528 1728 20534
rect 1676 20470 1728 20476
rect 1584 20460 1636 20466
rect 1584 20402 1636 20408
rect 1596 19922 1624 20402
rect 1688 19990 1716 20470
rect 1780 20346 1808 21542
rect 1872 21146 1900 22034
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 1780 20318 1900 20346
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1676 19984 1728 19990
rect 1676 19926 1728 19932
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1308 19304 1360 19310
rect 1308 19246 1360 19252
rect 1398 19272 1454 19281
rect 1320 17746 1348 19246
rect 1398 19207 1454 19216
rect 1412 18834 1440 19207
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1400 18148 1452 18154
rect 1400 18090 1452 18096
rect 1308 17740 1360 17746
rect 1308 17682 1360 17688
rect 1412 15910 1440 18090
rect 1504 17241 1532 18906
rect 1780 18834 1808 20198
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1584 18692 1636 18698
rect 1584 18634 1636 18640
rect 1596 18222 1624 18634
rect 1584 18216 1636 18222
rect 1584 18158 1636 18164
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1688 17882 1716 18158
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1596 16658 1624 17478
rect 1780 17202 1808 18770
rect 1872 17921 1900 20318
rect 1964 20058 1992 26182
rect 2056 24585 2084 26386
rect 2148 26314 2176 27639
rect 2240 26450 2268 27832
rect 2228 26444 2280 26450
rect 2228 26386 2280 26392
rect 2136 26308 2188 26314
rect 2136 26250 2188 26256
rect 2228 26308 2280 26314
rect 2228 26250 2280 26256
rect 2148 25294 2176 26250
rect 2240 25945 2268 26250
rect 2332 26246 2360 29446
rect 2424 28506 2452 31300
rect 2608 31142 2636 32150
rect 2700 31890 2728 32166
rect 2688 31884 2740 31890
rect 2688 31826 2740 31832
rect 2792 31793 2820 32558
rect 2872 32360 2924 32366
rect 2872 32302 2924 32308
rect 2778 31784 2834 31793
rect 2778 31719 2834 31728
rect 2884 31482 2912 32302
rect 3068 31754 3096 32914
rect 3160 32348 3188 33934
rect 3252 32502 3280 35822
rect 3344 35306 3372 36230
rect 3516 36236 3568 36242
rect 3516 36178 3568 36184
rect 4068 36236 4120 36242
rect 4120 36196 4200 36224
rect 4068 36178 4120 36184
rect 3344 35278 3464 35306
rect 3436 35222 3464 35278
rect 3332 35216 3384 35222
rect 3332 35158 3384 35164
rect 3424 35216 3476 35222
rect 3424 35158 3476 35164
rect 3240 32496 3292 32502
rect 3240 32438 3292 32444
rect 3240 32360 3292 32366
rect 3160 32320 3240 32348
rect 3240 32302 3292 32308
rect 3252 31958 3280 32302
rect 3240 31952 3292 31958
rect 3146 31920 3202 31929
rect 3344 31929 3372 35158
rect 3424 35080 3476 35086
rect 3424 35022 3476 35028
rect 3436 34542 3464 35022
rect 3424 34536 3476 34542
rect 3424 34478 3476 34484
rect 3528 34474 3556 36178
rect 3662 35932 3970 35941
rect 3662 35930 3668 35932
rect 3724 35930 3748 35932
rect 3804 35930 3828 35932
rect 3884 35930 3908 35932
rect 3964 35930 3970 35932
rect 3724 35878 3726 35930
rect 3906 35878 3908 35930
rect 3662 35876 3668 35878
rect 3724 35876 3748 35878
rect 3804 35876 3828 35878
rect 3884 35876 3908 35878
rect 3964 35876 3970 35878
rect 3662 35867 3970 35876
rect 4066 35864 4122 35873
rect 3884 35828 3936 35834
rect 3884 35770 3936 35776
rect 3976 35828 4028 35834
rect 4066 35799 4122 35808
rect 3976 35770 4028 35776
rect 3896 34932 3924 35770
rect 3988 35630 4016 35770
rect 4080 35766 4108 35799
rect 4068 35760 4120 35766
rect 4068 35702 4120 35708
rect 4172 35630 4200 36196
rect 4252 35692 4304 35698
rect 4252 35634 4304 35640
rect 3976 35624 4028 35630
rect 3976 35566 4028 35572
rect 4160 35624 4212 35630
rect 4160 35566 4212 35572
rect 3974 35184 4030 35193
rect 3974 35119 3976 35128
rect 4028 35119 4030 35128
rect 3976 35090 4028 35096
rect 3896 34904 4108 34932
rect 3662 34844 3970 34853
rect 3662 34842 3668 34844
rect 3724 34842 3748 34844
rect 3804 34842 3828 34844
rect 3884 34842 3908 34844
rect 3964 34842 3970 34844
rect 3724 34790 3726 34842
rect 3906 34790 3908 34842
rect 3662 34788 3668 34790
rect 3724 34788 3748 34790
rect 3804 34788 3828 34790
rect 3884 34788 3908 34790
rect 3964 34788 3970 34790
rect 3662 34779 3970 34788
rect 4080 34785 4108 34904
rect 4066 34776 4122 34785
rect 3608 34740 3660 34746
rect 4066 34711 4122 34720
rect 3608 34682 3660 34688
rect 3516 34468 3568 34474
rect 3516 34410 3568 34416
rect 3620 34354 3648 34682
rect 3974 34640 4030 34649
rect 3974 34575 3976 34584
rect 4028 34575 4030 34584
rect 3976 34546 4028 34552
rect 3792 34536 3844 34542
rect 3790 34504 3792 34513
rect 4068 34536 4120 34542
rect 3844 34504 3846 34513
rect 4068 34478 4120 34484
rect 3790 34439 3846 34448
rect 3528 34326 3648 34354
rect 3424 34060 3476 34066
rect 3424 34002 3476 34008
rect 3436 33658 3464 34002
rect 3424 33652 3476 33658
rect 3424 33594 3476 33600
rect 3528 33538 3556 34326
rect 3662 33756 3970 33765
rect 3662 33754 3668 33756
rect 3724 33754 3748 33756
rect 3804 33754 3828 33756
rect 3884 33754 3908 33756
rect 3964 33754 3970 33756
rect 3724 33702 3726 33754
rect 3906 33702 3908 33754
rect 3662 33700 3668 33702
rect 3724 33700 3748 33702
rect 3804 33700 3828 33702
rect 3884 33700 3908 33702
rect 3964 33700 3970 33702
rect 3662 33691 3970 33700
rect 3436 33510 3556 33538
rect 3240 31894 3292 31900
rect 3330 31920 3386 31929
rect 3146 31855 3202 31864
rect 2976 31726 3096 31754
rect 2872 31476 2924 31482
rect 2872 31418 2924 31424
rect 2780 31408 2832 31414
rect 2976 31362 3004 31726
rect 3160 31482 3188 31855
rect 3148 31476 3200 31482
rect 3148 31418 3200 31424
rect 2832 31356 3004 31362
rect 2780 31350 3004 31356
rect 2792 31334 3004 31350
rect 2872 31204 2924 31210
rect 2872 31146 2924 31152
rect 2596 31136 2648 31142
rect 2596 31078 2648 31084
rect 2596 30796 2648 30802
rect 2596 30738 2648 30744
rect 2688 30796 2740 30802
rect 2688 30738 2740 30744
rect 2608 30374 2636 30738
rect 2516 30346 2636 30374
rect 2516 28801 2544 30346
rect 2596 29844 2648 29850
rect 2700 29832 2728 30738
rect 2780 30660 2832 30666
rect 2780 30602 2832 30608
rect 2648 29804 2728 29832
rect 2792 29832 2820 30602
rect 2884 30394 2912 31146
rect 2976 30938 3004 31334
rect 3056 31340 3108 31346
rect 3056 31282 3108 31288
rect 2964 30932 3016 30938
rect 2964 30874 3016 30880
rect 2964 30592 3016 30598
rect 2962 30560 2964 30569
rect 3016 30560 3018 30569
rect 2962 30495 3018 30504
rect 2872 30388 2924 30394
rect 2872 30330 2924 30336
rect 2964 30184 3016 30190
rect 3068 30172 3096 31282
rect 3016 30144 3096 30172
rect 2964 30126 3016 30132
rect 3160 30122 3188 31418
rect 3252 31278 3280 31894
rect 3330 31855 3386 31864
rect 3330 31784 3386 31793
rect 3330 31719 3386 31728
rect 3240 31272 3292 31278
rect 3240 31214 3292 31220
rect 3240 31136 3292 31142
rect 3240 31078 3292 31084
rect 3252 30394 3280 31078
rect 3344 30938 3372 31719
rect 3436 30977 3464 33510
rect 3976 33312 4028 33318
rect 3974 33280 3976 33289
rect 4080 33300 4108 34478
rect 4028 33280 4108 33300
rect 4030 33272 4108 33280
rect 3974 33215 4030 33224
rect 3698 33008 3754 33017
rect 3516 32972 3568 32978
rect 3698 32943 3700 32952
rect 3516 32914 3568 32920
rect 3752 32943 3754 32952
rect 3700 32914 3752 32920
rect 3528 32570 3556 32914
rect 4068 32768 4120 32774
rect 4068 32710 4120 32716
rect 3662 32668 3970 32677
rect 3662 32666 3668 32668
rect 3724 32666 3748 32668
rect 3804 32666 3828 32668
rect 3884 32666 3908 32668
rect 3964 32666 3970 32668
rect 3724 32614 3726 32666
rect 3906 32614 3908 32666
rect 3662 32612 3668 32614
rect 3724 32612 3748 32614
rect 3804 32612 3828 32614
rect 3884 32612 3908 32614
rect 3964 32612 3970 32614
rect 3662 32603 3970 32612
rect 3516 32564 3568 32570
rect 3516 32506 3568 32512
rect 3528 32450 3556 32506
rect 3700 32496 3752 32502
rect 3528 32422 3648 32450
rect 3700 32438 3752 32444
rect 3516 32224 3568 32230
rect 3516 32166 3568 32172
rect 3528 31113 3556 32166
rect 3620 31793 3648 32422
rect 3606 31784 3662 31793
rect 3606 31719 3662 31728
rect 3712 31686 3740 32438
rect 3884 32360 3936 32366
rect 3804 32320 3884 32348
rect 3804 32026 3832 32320
rect 3884 32302 3936 32308
rect 3792 32020 3844 32026
rect 3792 31962 3844 31968
rect 3700 31680 3752 31686
rect 3700 31622 3752 31628
rect 3662 31580 3970 31589
rect 3662 31578 3668 31580
rect 3724 31578 3748 31580
rect 3804 31578 3828 31580
rect 3884 31578 3908 31580
rect 3964 31578 3970 31580
rect 3724 31526 3726 31578
rect 3906 31526 3908 31578
rect 3662 31524 3668 31526
rect 3724 31524 3748 31526
rect 3804 31524 3828 31526
rect 3884 31524 3908 31526
rect 3964 31524 3970 31526
rect 3662 31515 3970 31524
rect 4080 31464 4108 32710
rect 3988 31436 4108 31464
rect 3514 31104 3570 31113
rect 3514 31039 3570 31048
rect 3422 30968 3478 30977
rect 3332 30932 3384 30938
rect 3422 30903 3478 30912
rect 3332 30874 3384 30880
rect 3424 30864 3476 30870
rect 3516 30864 3568 30870
rect 3424 30806 3476 30812
rect 3514 30832 3516 30841
rect 3568 30832 3570 30841
rect 3330 30696 3386 30705
rect 3330 30631 3386 30640
rect 3240 30388 3292 30394
rect 3240 30330 3292 30336
rect 3148 30116 3200 30122
rect 3148 30058 3200 30064
rect 3252 30036 3280 30330
rect 3344 30190 3372 30631
rect 3436 30190 3464 30806
rect 3514 30767 3570 30776
rect 3516 30728 3568 30734
rect 3516 30670 3568 30676
rect 3332 30184 3384 30190
rect 3332 30126 3384 30132
rect 3424 30184 3476 30190
rect 3424 30126 3476 30132
rect 3252 30008 3464 30036
rect 2872 29844 2924 29850
rect 2792 29804 2872 29832
rect 2596 29786 2648 29792
rect 2872 29786 2924 29792
rect 2502 28792 2558 28801
rect 2502 28727 2558 28736
rect 2424 28478 2544 28506
rect 2412 28416 2464 28422
rect 2412 28358 2464 28364
rect 2424 27538 2452 28358
rect 2412 27532 2464 27538
rect 2412 27474 2464 27480
rect 2410 27024 2466 27033
rect 2410 26959 2412 26968
rect 2464 26959 2466 26968
rect 2412 26930 2464 26936
rect 2516 26874 2544 28478
rect 2608 28257 2636 29786
rect 3436 29782 3464 30008
rect 3424 29776 3476 29782
rect 2870 29744 2926 29753
rect 2792 29688 2870 29696
rect 2792 29668 2872 29688
rect 2688 29504 2740 29510
rect 2688 29446 2740 29452
rect 2700 28529 2728 29446
rect 2792 28665 2820 29668
rect 2924 29679 2926 29688
rect 3146 29744 3202 29753
rect 3424 29718 3476 29724
rect 3146 29679 3202 29688
rect 3332 29708 3384 29714
rect 2872 29650 2924 29656
rect 3160 29646 3188 29679
rect 3332 29650 3384 29656
rect 3148 29640 3200 29646
rect 3148 29582 3200 29588
rect 2964 29504 3016 29510
rect 2964 29446 3016 29452
rect 2870 29200 2926 29209
rect 2870 29135 2926 29144
rect 2884 29080 2912 29135
rect 2872 29074 2924 29080
rect 2872 29016 2924 29022
rect 2872 28960 2924 28966
rect 2870 28928 2872 28937
rect 2924 28928 2926 28937
rect 2870 28863 2926 28872
rect 2976 28762 3004 29446
rect 3056 29232 3108 29238
rect 3056 29174 3108 29180
rect 2964 28756 3016 28762
rect 2964 28698 3016 28704
rect 2778 28656 2834 28665
rect 2778 28591 2834 28600
rect 2872 28620 2924 28626
rect 3068 28608 3096 29174
rect 3160 29170 3188 29582
rect 3148 29164 3200 29170
rect 3148 29106 3200 29112
rect 3344 29034 3372 29650
rect 3240 29028 3292 29034
rect 3240 28970 3292 28976
rect 3332 29028 3384 29034
rect 3332 28970 3384 28976
rect 3252 28744 3280 28970
rect 3332 28756 3384 28762
rect 3252 28716 3332 28744
rect 3332 28698 3384 28704
rect 3344 28626 3372 28698
rect 3332 28620 3384 28626
rect 3068 28580 3188 28608
rect 2872 28562 2924 28568
rect 2686 28520 2742 28529
rect 2686 28455 2742 28464
rect 2780 28484 2832 28490
rect 2780 28426 2832 28432
rect 2594 28248 2650 28257
rect 2594 28183 2650 28192
rect 2608 28082 2636 28183
rect 2792 28132 2820 28426
rect 2884 28257 2912 28562
rect 2964 28416 3016 28422
rect 2964 28358 3016 28364
rect 2870 28248 2926 28257
rect 2870 28183 2926 28192
rect 2976 28200 3004 28358
rect 3160 28218 3188 28580
rect 3332 28562 3384 28568
rect 3240 28552 3292 28558
rect 3240 28494 3292 28500
rect 3056 28212 3108 28218
rect 2976 28172 3056 28200
rect 3056 28154 3108 28160
rect 3148 28212 3200 28218
rect 3148 28154 3200 28160
rect 2792 28104 3004 28132
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 2594 27976 2650 27985
rect 2594 27911 2650 27920
rect 2688 27940 2740 27946
rect 2608 27334 2636 27911
rect 2688 27882 2740 27888
rect 2700 27713 2728 27882
rect 2780 27872 2832 27878
rect 2780 27814 2832 27820
rect 2870 27840 2926 27849
rect 2686 27704 2742 27713
rect 2686 27639 2742 27648
rect 2792 27606 2820 27814
rect 2870 27775 2926 27784
rect 2780 27600 2832 27606
rect 2780 27542 2832 27548
rect 2688 27532 2740 27538
rect 2688 27474 2740 27480
rect 2596 27328 2648 27334
rect 2700 27305 2728 27474
rect 2780 27328 2832 27334
rect 2596 27270 2648 27276
rect 2686 27296 2742 27305
rect 2780 27270 2832 27276
rect 2686 27231 2742 27240
rect 2792 27130 2820 27270
rect 2688 27124 2740 27130
rect 2688 27066 2740 27072
rect 2780 27124 2832 27130
rect 2780 27066 2832 27072
rect 2594 27024 2650 27033
rect 2594 26959 2596 26968
rect 2648 26959 2650 26968
rect 2596 26930 2648 26936
rect 2412 26852 2464 26858
rect 2516 26846 2636 26874
rect 2412 26794 2464 26800
rect 2424 26382 2452 26794
rect 2504 26784 2556 26790
rect 2504 26726 2556 26732
rect 2516 26450 2544 26726
rect 2504 26444 2556 26450
rect 2504 26386 2556 26392
rect 2412 26376 2464 26382
rect 2412 26318 2464 26324
rect 2502 26344 2558 26353
rect 2502 26279 2558 26288
rect 2320 26240 2372 26246
rect 2320 26182 2372 26188
rect 2410 26208 2466 26217
rect 2410 26143 2466 26152
rect 2318 26072 2374 26081
rect 2318 26007 2320 26016
rect 2372 26007 2374 26016
rect 2320 25978 2372 25984
rect 2226 25936 2282 25945
rect 2226 25871 2282 25880
rect 2228 25832 2280 25838
rect 2228 25774 2280 25780
rect 2320 25832 2372 25838
rect 2320 25774 2372 25780
rect 2240 25362 2268 25774
rect 2228 25356 2280 25362
rect 2228 25298 2280 25304
rect 2136 25288 2188 25294
rect 2136 25230 2188 25236
rect 2042 24576 2098 24585
rect 2042 24511 2098 24520
rect 2042 24440 2098 24449
rect 2042 24375 2098 24384
rect 2056 23186 2084 24375
rect 2148 23186 2176 25230
rect 2240 24750 2268 25298
rect 2332 24993 2360 25774
rect 2424 25430 2452 26143
rect 2516 25974 2544 26279
rect 2608 25974 2636 26846
rect 2700 26489 2728 27066
rect 2780 26580 2832 26586
rect 2780 26522 2832 26528
rect 2686 26480 2742 26489
rect 2686 26415 2742 26424
rect 2688 26240 2740 26246
rect 2688 26182 2740 26188
rect 2504 25968 2556 25974
rect 2504 25910 2556 25916
rect 2596 25968 2648 25974
rect 2596 25910 2648 25916
rect 2504 25832 2556 25838
rect 2504 25774 2556 25780
rect 2596 25832 2648 25838
rect 2596 25774 2648 25780
rect 2516 25498 2544 25774
rect 2608 25537 2636 25774
rect 2594 25528 2650 25537
rect 2504 25492 2556 25498
rect 2594 25463 2650 25472
rect 2504 25434 2556 25440
rect 2412 25424 2464 25430
rect 2412 25366 2464 25372
rect 2410 25120 2466 25129
rect 2410 25055 2466 25064
rect 2318 24984 2374 24993
rect 2318 24919 2374 24928
rect 2424 24857 2452 25055
rect 2410 24848 2466 24857
rect 2332 24806 2410 24834
rect 2228 24744 2280 24750
rect 2228 24686 2280 24692
rect 2240 24206 2268 24686
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2240 23662 2268 24142
rect 2228 23656 2280 23662
rect 2228 23598 2280 23604
rect 2332 23594 2360 24806
rect 2410 24783 2466 24792
rect 2504 24812 2556 24818
rect 2556 24772 2636 24800
rect 2504 24754 2556 24760
rect 2412 24744 2464 24750
rect 2412 24686 2464 24692
rect 2424 23866 2452 24686
rect 2608 24614 2636 24772
rect 2504 24608 2556 24614
rect 2504 24550 2556 24556
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 2516 24274 2544 24550
rect 2594 24304 2650 24313
rect 2504 24268 2556 24274
rect 2594 24239 2596 24248
rect 2504 24210 2556 24216
rect 2648 24239 2650 24248
rect 2596 24210 2648 24216
rect 2412 23860 2464 23866
rect 2412 23802 2464 23808
rect 2516 23798 2544 24210
rect 2596 24064 2648 24070
rect 2596 24006 2648 24012
rect 2504 23792 2556 23798
rect 2504 23734 2556 23740
rect 2502 23624 2558 23633
rect 2320 23588 2372 23594
rect 2502 23559 2558 23568
rect 2320 23530 2372 23536
rect 2226 23216 2282 23225
rect 2044 23180 2096 23186
rect 2044 23122 2096 23128
rect 2136 23180 2188 23186
rect 2226 23151 2228 23160
rect 2136 23122 2188 23128
rect 2280 23151 2282 23160
rect 2320 23180 2372 23186
rect 2228 23122 2280 23128
rect 2320 23122 2372 23128
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 2056 21672 2084 23122
rect 2148 21842 2176 23122
rect 2228 23044 2280 23050
rect 2228 22986 2280 22992
rect 2240 22409 2268 22986
rect 2226 22400 2282 22409
rect 2226 22335 2282 22344
rect 2332 22234 2360 23122
rect 2424 22778 2452 23122
rect 2412 22772 2464 22778
rect 2412 22714 2464 22720
rect 2320 22228 2372 22234
rect 2320 22170 2372 22176
rect 2320 22024 2372 22030
rect 2320 21966 2372 21972
rect 2148 21814 2268 21842
rect 2056 21644 2176 21672
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2056 21010 2084 21490
rect 2148 21146 2176 21644
rect 2240 21622 2268 21814
rect 2228 21616 2280 21622
rect 2228 21558 2280 21564
rect 2332 21468 2360 21966
rect 2424 21554 2452 22714
rect 2516 22438 2544 23559
rect 2608 23322 2636 24006
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 2596 22704 2648 22710
rect 2596 22646 2648 22652
rect 2504 22432 2556 22438
rect 2502 22400 2504 22409
rect 2556 22400 2558 22409
rect 2502 22335 2558 22344
rect 2502 22264 2558 22273
rect 2502 22199 2558 22208
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 2240 21440 2360 21468
rect 2240 21350 2268 21440
rect 2516 21418 2544 22199
rect 2608 21729 2636 22646
rect 2700 22522 2728 26182
rect 2792 25430 2820 26522
rect 2780 25424 2832 25430
rect 2778 25392 2780 25401
rect 2832 25392 2834 25401
rect 2778 25327 2834 25336
rect 2780 25288 2832 25294
rect 2780 25230 2832 25236
rect 2792 24886 2820 25230
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 2780 24676 2832 24682
rect 2780 24618 2832 24624
rect 2792 23769 2820 24618
rect 2778 23760 2834 23769
rect 2778 23695 2834 23704
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2792 22642 2820 23462
rect 2884 22982 2912 27775
rect 2976 25945 3004 28104
rect 3148 28076 3200 28082
rect 3148 28018 3200 28024
rect 3056 27396 3108 27402
rect 3056 27338 3108 27344
rect 3068 27169 3096 27338
rect 3054 27160 3110 27169
rect 3054 27095 3110 27104
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 3068 26217 3096 26318
rect 3054 26208 3110 26217
rect 3054 26143 3110 26152
rect 3056 25968 3108 25974
rect 2962 25936 3018 25945
rect 3056 25910 3108 25916
rect 2962 25871 3018 25880
rect 2964 25832 3016 25838
rect 2964 25774 3016 25780
rect 2976 25498 3004 25774
rect 3068 25702 3096 25910
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 2964 25492 3016 25498
rect 2964 25434 3016 25440
rect 2964 25356 3016 25362
rect 2964 25298 3016 25304
rect 3056 25356 3108 25362
rect 3056 25298 3108 25304
rect 2976 24206 3004 25298
rect 2964 24200 3016 24206
rect 3068 24177 3096 25298
rect 2964 24142 3016 24148
rect 3054 24168 3110 24177
rect 3054 24103 3056 24112
rect 3108 24103 3110 24112
rect 3056 24074 3108 24080
rect 3068 23746 3096 24074
rect 2976 23718 3096 23746
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2700 22494 2820 22522
rect 2688 22432 2740 22438
rect 2688 22374 2740 22380
rect 2700 22098 2728 22374
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2594 21720 2650 21729
rect 2594 21655 2650 21664
rect 2596 21616 2648 21622
rect 2596 21558 2648 21564
rect 2504 21412 2556 21418
rect 2504 21354 2556 21360
rect 2228 21344 2280 21350
rect 2228 21286 2280 21292
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2136 21140 2188 21146
rect 2136 21082 2188 21088
rect 2044 21004 2096 21010
rect 2044 20946 2096 20952
rect 2134 20632 2190 20641
rect 2134 20567 2190 20576
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 2056 19514 2084 20334
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 2148 18970 2176 20567
rect 2240 20398 2268 21286
rect 2332 21010 2360 21286
rect 2504 21140 2556 21146
rect 2504 21082 2556 21088
rect 2516 21010 2544 21082
rect 2320 21004 2372 21010
rect 2320 20946 2372 20952
rect 2504 21004 2556 21010
rect 2504 20946 2556 20952
rect 2608 20992 2636 21558
rect 2700 21418 2728 22034
rect 2688 21412 2740 21418
rect 2688 21354 2740 21360
rect 2688 21004 2740 21010
rect 2608 20964 2688 20992
rect 2516 20398 2544 20946
rect 2608 20602 2636 20964
rect 2688 20946 2740 20952
rect 2792 20890 2820 22494
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 2884 21894 2912 22374
rect 2976 22234 3004 23718
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 3068 23497 3096 23598
rect 3054 23488 3110 23497
rect 3054 23423 3110 23432
rect 3068 22710 3096 23423
rect 3056 22704 3108 22710
rect 3056 22646 3108 22652
rect 3054 22400 3110 22409
rect 3054 22335 3110 22344
rect 2964 22228 3016 22234
rect 2964 22170 3016 22176
rect 2964 22092 3016 22098
rect 2964 22034 3016 22040
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2884 21486 2912 21830
rect 2872 21480 2924 21486
rect 2872 21422 2924 21428
rect 2700 20862 2820 20890
rect 2596 20596 2648 20602
rect 2596 20538 2648 20544
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 2240 19854 2268 20334
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2240 19310 2268 19790
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 2056 18426 2084 18770
rect 2148 18766 2176 18906
rect 2240 18766 2268 19246
rect 2332 18834 2360 19858
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1858 17912 1914 17921
rect 1858 17847 1914 17856
rect 1860 17604 1912 17610
rect 1860 17546 1912 17552
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1780 16130 1808 17138
rect 1688 16102 1808 16130
rect 1688 16046 1716 16102
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1768 15428 1820 15434
rect 1768 15370 1820 15376
rect 1492 15088 1544 15094
rect 1492 15030 1544 15036
rect 1504 14822 1532 15030
rect 1780 14958 1808 15370
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 14074 1440 14350
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1308 12776 1360 12782
rect 1308 12718 1360 12724
rect 1214 12608 1270 12617
rect 1214 12543 1270 12552
rect 1320 10606 1348 12718
rect 1412 11762 1440 13874
rect 1504 13530 1532 14418
rect 1492 13524 1544 13530
rect 1492 13466 1544 13472
rect 1596 12442 1624 14894
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1766 14784 1822 14793
rect 1688 13938 1716 14758
rect 1766 14719 1822 14728
rect 1780 14618 1808 14719
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1674 13832 1730 13841
rect 1674 13767 1730 13776
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1688 12306 1716 13767
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1780 13394 1808 13670
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1872 12481 1900 17546
rect 1964 17134 1992 18022
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 2056 16658 2084 17478
rect 2148 17338 2176 17682
rect 2240 17678 2268 18702
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2332 18290 2360 18566
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2424 18136 2452 19722
rect 2516 19310 2544 19926
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2608 19378 2636 19858
rect 2700 19718 2728 20862
rect 2780 20392 2832 20398
rect 2778 20360 2780 20369
rect 2832 20360 2834 20369
rect 2778 20295 2834 20304
rect 2884 19990 2912 21422
rect 2976 21026 3004 22034
rect 3068 22001 3096 22335
rect 3054 21992 3110 22001
rect 3054 21927 3110 21936
rect 3054 21720 3110 21729
rect 3160 21690 3188 28018
rect 3252 27470 3280 28494
rect 3240 27464 3292 27470
rect 3240 27406 3292 27412
rect 3252 27334 3280 27406
rect 3240 27328 3292 27334
rect 3240 27270 3292 27276
rect 3238 27160 3294 27169
rect 3238 27095 3294 27104
rect 3252 25974 3280 27095
rect 3344 27033 3372 28562
rect 3528 28506 3556 30670
rect 3988 30666 4016 31436
rect 4068 31272 4120 31278
rect 4068 31214 4120 31220
rect 4080 30818 4108 31214
rect 4172 30938 4200 35566
rect 4264 35290 4292 35634
rect 4322 35388 4630 35397
rect 4322 35386 4328 35388
rect 4384 35386 4408 35388
rect 4464 35386 4488 35388
rect 4544 35386 4568 35388
rect 4624 35386 4630 35388
rect 4384 35334 4386 35386
rect 4566 35334 4568 35386
rect 4322 35332 4328 35334
rect 4384 35332 4408 35334
rect 4464 35332 4488 35334
rect 4544 35332 4568 35334
rect 4624 35332 4630 35334
rect 4322 35323 4630 35332
rect 4252 35284 4304 35290
rect 4252 35226 4304 35232
rect 4344 35080 4396 35086
rect 4344 35022 4396 35028
rect 4618 35048 4674 35057
rect 4356 34746 4384 35022
rect 4618 34983 4674 34992
rect 4344 34740 4396 34746
rect 4344 34682 4396 34688
rect 4632 34678 4660 34983
rect 4620 34672 4672 34678
rect 4620 34614 4672 34620
rect 4252 34604 4304 34610
rect 4252 34546 4304 34552
rect 4264 33454 4292 34546
rect 4620 34536 4672 34542
rect 4724 34524 4752 36638
rect 4816 35494 4844 37046
rect 4896 36032 4948 36038
rect 4896 35974 4948 35980
rect 4804 35488 4856 35494
rect 4804 35430 4856 35436
rect 4672 34496 4752 34524
rect 4804 34536 4856 34542
rect 4620 34478 4672 34484
rect 4908 34524 4936 35974
rect 5000 35494 5028 38791
rect 5184 38729 5212 39918
rect 5276 39438 5304 39936
rect 5448 39918 5500 39924
rect 5356 39840 5408 39846
rect 5356 39782 5408 39788
rect 5264 39432 5316 39438
rect 5264 39374 5316 39380
rect 5170 38720 5226 38729
rect 5170 38655 5226 38664
rect 5368 38554 5396 39782
rect 5460 39574 5488 39918
rect 5540 39840 5592 39846
rect 5540 39782 5592 39788
rect 5448 39568 5500 39574
rect 5448 39510 5500 39516
rect 5356 38548 5408 38554
rect 5356 38490 5408 38496
rect 5552 37806 5580 39782
rect 5632 39432 5684 39438
rect 5632 39374 5684 39380
rect 5736 39386 5764 41618
rect 5908 41472 5960 41478
rect 5908 41414 5960 41420
rect 5920 41070 5948 41414
rect 6104 41138 6132 42162
rect 6196 41414 6224 42570
rect 6552 42356 6604 42362
rect 6552 42298 6604 42304
rect 6460 42016 6512 42022
rect 6460 41958 6512 41964
rect 6472 41546 6500 41958
rect 6460 41540 6512 41546
rect 6460 41482 6512 41488
rect 6472 41414 6500 41482
rect 6196 41386 6316 41414
rect 6092 41132 6144 41138
rect 6092 41074 6144 41080
rect 5908 41064 5960 41070
rect 5908 41006 5960 41012
rect 6104 40730 6132 41074
rect 6092 40724 6144 40730
rect 6092 40666 6144 40672
rect 6184 40656 6236 40662
rect 6184 40598 6236 40604
rect 5816 40520 5868 40526
rect 5816 40462 5868 40468
rect 5828 39506 5856 40462
rect 6196 40089 6224 40598
rect 6182 40080 6238 40089
rect 6182 40015 6238 40024
rect 6288 39953 6316 41386
rect 6380 41386 6500 41414
rect 6274 39944 6330 39953
rect 6274 39879 6330 39888
rect 5998 39808 6054 39817
rect 5998 39743 6054 39752
rect 5816 39500 5868 39506
rect 5816 39442 5868 39448
rect 5644 39030 5672 39374
rect 5736 39358 5856 39386
rect 5724 39296 5776 39302
rect 5724 39238 5776 39244
rect 5736 39098 5764 39238
rect 5724 39092 5776 39098
rect 5724 39034 5776 39040
rect 5632 39024 5684 39030
rect 5632 38966 5684 38972
rect 5722 38584 5778 38593
rect 5722 38519 5778 38528
rect 5632 38412 5684 38418
rect 5632 38354 5684 38360
rect 5644 38010 5672 38354
rect 5632 38004 5684 38010
rect 5632 37946 5684 37952
rect 5448 37800 5500 37806
rect 5448 37742 5500 37748
rect 5540 37800 5592 37806
rect 5540 37742 5592 37748
rect 5460 37330 5488 37742
rect 5172 37324 5224 37330
rect 5172 37266 5224 37272
rect 5264 37324 5316 37330
rect 5264 37266 5316 37272
rect 5356 37324 5408 37330
rect 5356 37266 5408 37272
rect 5448 37324 5500 37330
rect 5448 37266 5500 37272
rect 5632 37324 5684 37330
rect 5632 37266 5684 37272
rect 5080 37256 5132 37262
rect 5080 37198 5132 37204
rect 4988 35488 5040 35494
rect 4988 35430 5040 35436
rect 5092 35086 5120 37198
rect 5184 36378 5212 37266
rect 5172 36372 5224 36378
rect 5172 36314 5224 36320
rect 5184 35630 5212 36314
rect 5172 35624 5224 35630
rect 5172 35566 5224 35572
rect 5172 35488 5224 35494
rect 5172 35430 5224 35436
rect 4988 35080 5040 35086
rect 4988 35022 5040 35028
rect 5080 35080 5132 35086
rect 5080 35022 5132 35028
rect 5000 34746 5028 35022
rect 5184 35018 5212 35430
rect 5276 35306 5304 37266
rect 5368 36718 5396 37266
rect 5460 36825 5488 37266
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5446 36816 5502 36825
rect 5446 36751 5502 36760
rect 5356 36712 5408 36718
rect 5356 36654 5408 36660
rect 5368 36038 5396 36654
rect 5552 36242 5580 37130
rect 5540 36236 5592 36242
rect 5540 36178 5592 36184
rect 5356 36032 5408 36038
rect 5356 35974 5408 35980
rect 5448 35828 5500 35834
rect 5448 35770 5500 35776
rect 5276 35278 5396 35306
rect 5264 35148 5316 35154
rect 5264 35090 5316 35096
rect 5172 35012 5224 35018
rect 5172 34954 5224 34960
rect 5078 34912 5134 34921
rect 5078 34847 5134 34856
rect 4988 34740 5040 34746
rect 4988 34682 5040 34688
rect 4856 34496 4936 34524
rect 4804 34478 4856 34484
rect 4896 34400 4948 34406
rect 4896 34342 4948 34348
rect 4322 34300 4630 34309
rect 4322 34298 4328 34300
rect 4384 34298 4408 34300
rect 4464 34298 4488 34300
rect 4544 34298 4568 34300
rect 4624 34298 4630 34300
rect 4384 34246 4386 34298
rect 4566 34246 4568 34298
rect 4322 34244 4328 34246
rect 4384 34244 4408 34246
rect 4464 34244 4488 34246
rect 4544 34244 4568 34246
rect 4624 34244 4630 34246
rect 4322 34235 4630 34244
rect 4908 34066 4936 34342
rect 4896 34060 4948 34066
rect 4896 34002 4948 34008
rect 4528 33924 4580 33930
rect 4528 33866 4580 33872
rect 4252 33448 4304 33454
rect 4252 33390 4304 33396
rect 4540 33318 4568 33866
rect 5092 33454 5120 34847
rect 5170 34776 5226 34785
rect 5276 34746 5304 35090
rect 5368 34950 5396 35278
rect 5460 35154 5488 35770
rect 5644 35222 5672 37266
rect 5632 35216 5684 35222
rect 5632 35158 5684 35164
rect 5448 35148 5500 35154
rect 5448 35090 5500 35096
rect 5356 34944 5408 34950
rect 5356 34886 5408 34892
rect 5170 34711 5172 34720
rect 5224 34711 5226 34720
rect 5264 34740 5316 34746
rect 5172 34682 5224 34688
rect 5264 34682 5316 34688
rect 5368 34542 5396 34886
rect 5356 34536 5408 34542
rect 5170 34504 5226 34513
rect 5356 34478 5408 34484
rect 5170 34439 5226 34448
rect 5264 34468 5316 34474
rect 5184 34066 5212 34439
rect 5264 34410 5316 34416
rect 5276 34066 5304 34410
rect 5460 34406 5488 35090
rect 5736 34490 5764 38519
rect 5828 37466 5856 39358
rect 5908 39092 5960 39098
rect 5908 39034 5960 39040
rect 5920 38894 5948 39034
rect 5908 38888 5960 38894
rect 5908 38830 5960 38836
rect 5908 38752 5960 38758
rect 5908 38694 5960 38700
rect 5920 38554 5948 38694
rect 5908 38548 5960 38554
rect 5908 38490 5960 38496
rect 5816 37460 5868 37466
rect 5816 37402 5868 37408
rect 5814 36816 5870 36825
rect 5814 36751 5870 36760
rect 5908 36780 5960 36786
rect 5828 36718 5856 36751
rect 5908 36722 5960 36728
rect 5816 36712 5868 36718
rect 5816 36654 5868 36660
rect 5814 36272 5870 36281
rect 5814 36207 5870 36216
rect 5828 35601 5856 36207
rect 5814 35592 5870 35601
rect 5814 35527 5870 35536
rect 5816 35488 5868 35494
rect 5816 35430 5868 35436
rect 5828 35290 5856 35430
rect 5816 35284 5868 35290
rect 5816 35226 5868 35232
rect 5920 34785 5948 36722
rect 6012 36122 6040 39743
rect 6092 39500 6144 39506
rect 6092 39442 6144 39448
rect 6104 37806 6132 39442
rect 6276 38344 6328 38350
rect 6276 38286 6328 38292
rect 6288 37874 6316 38286
rect 6276 37868 6328 37874
rect 6276 37810 6328 37816
rect 6092 37800 6144 37806
rect 6092 37742 6144 37748
rect 6104 37398 6132 37742
rect 6184 37732 6236 37738
rect 6184 37674 6236 37680
rect 6276 37732 6328 37738
rect 6276 37674 6328 37680
rect 6196 37466 6224 37674
rect 6184 37460 6236 37466
rect 6184 37402 6236 37408
rect 6092 37392 6144 37398
rect 6092 37334 6144 37340
rect 6288 37330 6316 37674
rect 6276 37324 6328 37330
rect 6276 37266 6328 37272
rect 6092 36780 6144 36786
rect 6092 36722 6144 36728
rect 6104 36242 6132 36722
rect 6184 36712 6236 36718
rect 6184 36654 6236 36660
rect 6196 36378 6224 36654
rect 6184 36372 6236 36378
rect 6184 36314 6236 36320
rect 6288 36310 6316 37266
rect 6276 36304 6328 36310
rect 6276 36246 6328 36252
rect 6092 36236 6144 36242
rect 6092 36178 6144 36184
rect 6276 36168 6328 36174
rect 6012 36094 6132 36122
rect 6276 36110 6328 36116
rect 6000 35488 6052 35494
rect 6000 35430 6052 35436
rect 6012 35154 6040 35430
rect 6000 35148 6052 35154
rect 6000 35090 6052 35096
rect 6000 35012 6052 35018
rect 6000 34954 6052 34960
rect 5906 34776 5962 34785
rect 5906 34711 5962 34720
rect 5552 34462 5764 34490
rect 5448 34400 5500 34406
rect 5354 34368 5410 34377
rect 5448 34342 5500 34348
rect 5354 34303 5410 34312
rect 5368 34202 5396 34303
rect 5356 34196 5408 34202
rect 5356 34138 5408 34144
rect 5172 34060 5224 34066
rect 5172 34002 5224 34008
rect 5264 34060 5316 34066
rect 5264 34002 5316 34008
rect 5552 33658 5580 34462
rect 5632 34400 5684 34406
rect 5632 34342 5684 34348
rect 5644 34066 5672 34342
rect 5632 34060 5684 34066
rect 5632 34002 5684 34008
rect 5816 34060 5868 34066
rect 5816 34002 5868 34008
rect 5724 33924 5776 33930
rect 5724 33866 5776 33872
rect 5540 33652 5592 33658
rect 5540 33594 5592 33600
rect 5538 33552 5594 33561
rect 5538 33487 5594 33496
rect 5552 33454 5580 33487
rect 5736 33454 5764 33866
rect 5828 33522 5856 34002
rect 6012 33946 6040 34954
rect 6104 33998 6132 36094
rect 6184 35624 6236 35630
rect 6184 35566 6236 35572
rect 6196 35086 6224 35566
rect 6184 35080 6236 35086
rect 6184 35022 6236 35028
rect 6196 34678 6224 35022
rect 6184 34672 6236 34678
rect 6184 34614 6236 34620
rect 6288 34626 6316 36110
rect 6380 35222 6408 41386
rect 6564 41018 6592 42298
rect 6644 41744 6696 41750
rect 6642 41712 6644 41721
rect 6696 41712 6698 41721
rect 6642 41647 6698 41656
rect 6736 41200 6788 41206
rect 6736 41142 6788 41148
rect 6472 40990 6592 41018
rect 6472 40066 6500 40990
rect 6552 40928 6604 40934
rect 6552 40870 6604 40876
rect 6644 40928 6696 40934
rect 6644 40870 6696 40876
rect 6564 40730 6592 40870
rect 6552 40724 6604 40730
rect 6552 40666 6604 40672
rect 6656 40089 6684 40870
rect 6748 40594 6776 41142
rect 6736 40588 6788 40594
rect 6736 40530 6788 40536
rect 6642 40080 6698 40089
rect 6472 40038 6592 40066
rect 6460 39908 6512 39914
rect 6460 39850 6512 39856
rect 6472 39506 6500 39850
rect 6564 39642 6592 40038
rect 6642 40015 6698 40024
rect 6644 39908 6696 39914
rect 6644 39850 6696 39856
rect 6656 39642 6684 39850
rect 6552 39636 6604 39642
rect 6552 39578 6604 39584
rect 6644 39636 6696 39642
rect 6644 39578 6696 39584
rect 6460 39500 6512 39506
rect 6460 39442 6512 39448
rect 6472 37126 6500 39442
rect 6748 39030 6776 40530
rect 7024 39846 7052 42638
rect 7656 42628 7708 42634
rect 7656 42570 7708 42576
rect 7668 42226 7696 42570
rect 7656 42220 7708 42226
rect 7656 42162 7708 42168
rect 7380 42152 7432 42158
rect 7380 42094 7432 42100
rect 7392 41682 7420 42094
rect 7564 42084 7616 42090
rect 7564 42026 7616 42032
rect 7380 41676 7432 41682
rect 7380 41618 7432 41624
rect 7576 41449 7604 42026
rect 7668 41750 7696 42162
rect 7760 42090 7788 42638
rect 8116 42220 8168 42226
rect 8116 42162 8168 42168
rect 7748 42084 7800 42090
rect 7748 42026 7800 42032
rect 7656 41744 7708 41750
rect 7656 41686 7708 41692
rect 7760 41585 7788 42026
rect 8128 41818 8156 42162
rect 8208 42016 8260 42022
rect 8208 41958 8260 41964
rect 8116 41812 8168 41818
rect 8116 41754 8168 41760
rect 7840 41676 7892 41682
rect 7840 41618 7892 41624
rect 7746 41576 7802 41585
rect 7746 41511 7802 41520
rect 7656 41472 7708 41478
rect 7562 41440 7618 41449
rect 7656 41414 7708 41420
rect 7562 41375 7618 41384
rect 7470 41304 7526 41313
rect 7668 41290 7696 41414
rect 7470 41239 7526 41248
rect 7576 41262 7696 41290
rect 7012 39840 7064 39846
rect 7012 39782 7064 39788
rect 7104 39840 7156 39846
rect 7104 39782 7156 39788
rect 7116 39642 7144 39782
rect 7104 39636 7156 39642
rect 7104 39578 7156 39584
rect 7380 39636 7432 39642
rect 7380 39578 7432 39584
rect 7104 39500 7156 39506
rect 7104 39442 7156 39448
rect 6826 39400 6882 39409
rect 6826 39335 6882 39344
rect 6920 39364 6972 39370
rect 6840 39098 6868 39335
rect 6920 39306 6972 39312
rect 6828 39092 6880 39098
rect 6828 39034 6880 39040
rect 6644 39024 6696 39030
rect 6644 38966 6696 38972
rect 6736 39024 6788 39030
rect 6736 38966 6788 38972
rect 6656 37330 6684 38966
rect 6736 38888 6788 38894
rect 6736 38830 6788 38836
rect 6748 38214 6776 38830
rect 6828 38820 6880 38826
rect 6828 38762 6880 38768
rect 6736 38208 6788 38214
rect 6736 38150 6788 38156
rect 6748 37806 6776 38150
rect 6840 37806 6868 38762
rect 6932 38350 6960 39306
rect 7116 38758 7144 39442
rect 7196 39432 7248 39438
rect 7196 39374 7248 39380
rect 7288 39432 7340 39438
rect 7288 39374 7340 39380
rect 7208 38962 7236 39374
rect 7300 39098 7328 39374
rect 7288 39092 7340 39098
rect 7288 39034 7340 39040
rect 7286 38992 7342 39001
rect 7196 38956 7248 38962
rect 7286 38927 7342 38936
rect 7196 38898 7248 38904
rect 7300 38894 7328 38927
rect 7288 38888 7340 38894
rect 7288 38830 7340 38836
rect 7104 38752 7156 38758
rect 7104 38694 7156 38700
rect 7012 38412 7064 38418
rect 7012 38354 7064 38360
rect 6920 38344 6972 38350
rect 6918 38312 6920 38321
rect 6972 38312 6974 38321
rect 6918 38247 6974 38256
rect 6736 37800 6788 37806
rect 6736 37742 6788 37748
rect 6828 37800 6880 37806
rect 6880 37760 6960 37788
rect 6828 37742 6880 37748
rect 6736 37664 6788 37670
rect 6736 37606 6788 37612
rect 6826 37632 6882 37641
rect 6748 37369 6776 37606
rect 6826 37567 6882 37576
rect 6734 37360 6790 37369
rect 6644 37324 6696 37330
rect 6734 37295 6790 37304
rect 6644 37266 6696 37272
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 6460 37120 6512 37126
rect 6460 37062 6512 37068
rect 6564 36718 6592 37198
rect 6552 36712 6604 36718
rect 6552 36654 6604 36660
rect 6564 36378 6592 36654
rect 6644 36644 6696 36650
rect 6644 36586 6696 36592
rect 6552 36372 6604 36378
rect 6552 36314 6604 36320
rect 6460 36168 6512 36174
rect 6460 36110 6512 36116
rect 6472 35290 6500 36110
rect 6656 35766 6684 36586
rect 6644 35760 6696 35766
rect 6644 35702 6696 35708
rect 6734 35728 6790 35737
rect 6734 35663 6790 35672
rect 6552 35556 6604 35562
rect 6552 35498 6604 35504
rect 6460 35284 6512 35290
rect 6460 35226 6512 35232
rect 6368 35216 6420 35222
rect 6368 35158 6420 35164
rect 6564 35086 6592 35498
rect 6644 35148 6696 35154
rect 6644 35090 6696 35096
rect 6552 35080 6604 35086
rect 6552 35022 6604 35028
rect 6656 34649 6684 35090
rect 6642 34640 6698 34649
rect 6288 34598 6408 34626
rect 6276 34536 6328 34542
rect 6276 34478 6328 34484
rect 6288 34202 6316 34478
rect 6276 34196 6328 34202
rect 6276 34138 6328 34144
rect 5920 33918 6040 33946
rect 6092 33992 6144 33998
rect 6380 33969 6408 34598
rect 6642 34575 6698 34584
rect 6656 34542 6684 34575
rect 6644 34536 6696 34542
rect 6644 34478 6696 34484
rect 6552 34400 6604 34406
rect 6552 34342 6604 34348
rect 6092 33934 6144 33940
rect 6366 33960 6422 33969
rect 5816 33516 5868 33522
rect 5816 33458 5868 33464
rect 5080 33448 5132 33454
rect 5080 33390 5132 33396
rect 5540 33448 5592 33454
rect 5540 33390 5592 33396
rect 5724 33448 5776 33454
rect 5724 33390 5776 33396
rect 4528 33312 4580 33318
rect 4528 33254 4580 33260
rect 5172 33312 5224 33318
rect 5172 33254 5224 33260
rect 4322 33212 4630 33221
rect 4322 33210 4328 33212
rect 4384 33210 4408 33212
rect 4464 33210 4488 33212
rect 4544 33210 4568 33212
rect 4624 33210 4630 33212
rect 4384 33158 4386 33210
rect 4566 33158 4568 33210
rect 4322 33156 4328 33158
rect 4384 33156 4408 33158
rect 4464 33156 4488 33158
rect 4544 33156 4568 33158
rect 4624 33156 4630 33158
rect 4322 33147 4630 33156
rect 4344 33108 4396 33114
rect 4344 33050 4396 33056
rect 4356 32978 4384 33050
rect 4434 33008 4490 33017
rect 4252 32972 4304 32978
rect 4252 32914 4304 32920
rect 4344 32972 4396 32978
rect 4434 32943 4490 32952
rect 4896 32972 4948 32978
rect 4344 32914 4396 32920
rect 4264 31414 4292 32914
rect 4448 32230 4476 32943
rect 4896 32914 4948 32920
rect 4908 32881 4936 32914
rect 4894 32872 4950 32881
rect 4620 32836 4672 32842
rect 4672 32796 4752 32824
rect 4894 32807 4950 32816
rect 4620 32778 4672 32784
rect 4436 32224 4488 32230
rect 4436 32166 4488 32172
rect 4322 32124 4630 32133
rect 4322 32122 4328 32124
rect 4384 32122 4408 32124
rect 4464 32122 4488 32124
rect 4544 32122 4568 32124
rect 4624 32122 4630 32124
rect 4384 32070 4386 32122
rect 4566 32070 4568 32122
rect 4322 32068 4328 32070
rect 4384 32068 4408 32070
rect 4464 32068 4488 32070
rect 4544 32068 4568 32070
rect 4624 32068 4630 32070
rect 4322 32059 4630 32068
rect 4724 32026 4752 32796
rect 4804 32292 4856 32298
rect 4804 32234 4856 32240
rect 4712 32020 4764 32026
rect 4632 31980 4712 32008
rect 4434 31920 4490 31929
rect 4434 31855 4436 31864
rect 4488 31855 4490 31864
rect 4436 31826 4488 31832
rect 4252 31408 4304 31414
rect 4252 31350 4304 31356
rect 4264 31142 4292 31350
rect 4632 31142 4660 31980
rect 4712 31962 4764 31968
rect 4710 31784 4766 31793
rect 4710 31719 4766 31728
rect 4252 31136 4304 31142
rect 4252 31078 4304 31084
rect 4620 31136 4672 31142
rect 4620 31078 4672 31084
rect 4160 30932 4212 30938
rect 4160 30874 4212 30880
rect 4264 30870 4292 31078
rect 4322 31036 4630 31045
rect 4322 31034 4328 31036
rect 4384 31034 4408 31036
rect 4464 31034 4488 31036
rect 4544 31034 4568 31036
rect 4624 31034 4630 31036
rect 4384 30982 4386 31034
rect 4566 30982 4568 31034
rect 4322 30980 4328 30982
rect 4384 30980 4408 30982
rect 4464 30980 4488 30982
rect 4544 30980 4568 30982
rect 4624 30980 4630 30982
rect 4322 30971 4630 30980
rect 4436 30932 4488 30938
rect 4436 30874 4488 30880
rect 4252 30864 4304 30870
rect 4080 30790 4200 30818
rect 4252 30806 4304 30812
rect 3976 30660 4028 30666
rect 3976 30602 4028 30608
rect 3662 30492 3970 30501
rect 3662 30490 3668 30492
rect 3724 30490 3748 30492
rect 3804 30490 3828 30492
rect 3884 30490 3908 30492
rect 3964 30490 3970 30492
rect 3724 30438 3726 30490
rect 3906 30438 3908 30490
rect 3662 30436 3668 30438
rect 3724 30436 3748 30438
rect 3804 30436 3828 30438
rect 3884 30436 3908 30438
rect 3964 30436 3970 30438
rect 3662 30427 3970 30436
rect 3884 30184 3936 30190
rect 3884 30126 3936 30132
rect 3896 29753 3924 30126
rect 4068 29776 4120 29782
rect 3882 29744 3938 29753
rect 4068 29718 4120 29724
rect 3882 29679 3938 29688
rect 3662 29404 3970 29413
rect 3662 29402 3668 29404
rect 3724 29402 3748 29404
rect 3804 29402 3828 29404
rect 3884 29402 3908 29404
rect 3964 29402 3970 29404
rect 3724 29350 3726 29402
rect 3906 29350 3908 29402
rect 3662 29348 3668 29350
rect 3724 29348 3748 29350
rect 3804 29348 3828 29350
rect 3884 29348 3908 29350
rect 3964 29348 3970 29350
rect 3662 29339 3970 29348
rect 3606 29200 3662 29209
rect 3606 29135 3662 29144
rect 3974 29200 4030 29209
rect 3974 29135 4030 29144
rect 3620 28937 3648 29135
rect 3884 28960 3936 28966
rect 3606 28928 3662 28937
rect 3884 28902 3936 28908
rect 3606 28863 3662 28872
rect 3608 28620 3660 28626
rect 3608 28562 3660 28568
rect 3620 28529 3648 28562
rect 3427 28478 3556 28506
rect 3606 28520 3662 28529
rect 3427 28132 3455 28478
rect 3606 28455 3662 28464
rect 3896 28422 3924 28902
rect 3988 28529 4016 29135
rect 4080 29102 4108 29718
rect 4068 29096 4120 29102
rect 4068 29038 4120 29044
rect 4080 28762 4108 29038
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 3974 28520 4030 28529
rect 3974 28455 4030 28464
rect 3608 28416 3660 28422
rect 3528 28376 3608 28404
rect 3528 28200 3556 28376
rect 3608 28358 3660 28364
rect 3884 28416 3936 28422
rect 3884 28358 3936 28364
rect 3662 28316 3970 28325
rect 3662 28314 3668 28316
rect 3724 28314 3748 28316
rect 3804 28314 3828 28316
rect 3884 28314 3908 28316
rect 3964 28314 3970 28316
rect 3724 28262 3726 28314
rect 3906 28262 3908 28314
rect 3662 28260 3668 28262
rect 3724 28260 3748 28262
rect 3804 28260 3828 28262
rect 3884 28260 3908 28262
rect 3964 28260 3970 28262
rect 3662 28251 3970 28260
rect 3608 28212 3660 28218
rect 3528 28172 3608 28200
rect 3608 28154 3660 28160
rect 3884 28212 3936 28218
rect 3884 28154 3936 28160
rect 3427 28104 3556 28132
rect 3528 28014 3556 28104
rect 3700 28076 3752 28082
rect 3700 28018 3752 28024
rect 3792 28076 3844 28082
rect 3792 28018 3844 28024
rect 3516 28008 3568 28014
rect 3516 27950 3568 27956
rect 3712 27713 3740 28018
rect 3698 27704 3754 27713
rect 3698 27639 3754 27648
rect 3804 27606 3832 28018
rect 3896 27849 3924 28154
rect 4068 28144 4120 28150
rect 4068 28086 4120 28092
rect 3882 27840 3938 27849
rect 3882 27775 3938 27784
rect 4080 27674 4108 28086
rect 4068 27668 4120 27674
rect 4068 27610 4120 27616
rect 3792 27600 3844 27606
rect 3792 27542 3844 27548
rect 3976 27532 4028 27538
rect 4172 27520 4200 30790
rect 4344 30660 4396 30666
rect 4344 30602 4396 30608
rect 4252 30592 4304 30598
rect 4252 30534 4304 30540
rect 4264 30326 4292 30534
rect 4356 30394 4384 30602
rect 4344 30388 4396 30394
rect 4344 30330 4396 30336
rect 4252 30320 4304 30326
rect 4252 30262 4304 30268
rect 4448 30190 4476 30874
rect 4436 30184 4488 30190
rect 4436 30126 4488 30132
rect 4724 30122 4752 31719
rect 4816 30598 4844 32234
rect 4908 31793 4936 32807
rect 4988 32768 5040 32774
rect 4988 32710 5040 32716
rect 5080 32768 5132 32774
rect 5080 32710 5132 32716
rect 4894 31784 4950 31793
rect 4894 31719 4950 31728
rect 4896 31408 4948 31414
rect 4896 31350 4948 31356
rect 4908 30734 4936 31350
rect 5000 31278 5028 32710
rect 4988 31272 5040 31278
rect 4988 31214 5040 31220
rect 4986 30968 5042 30977
rect 4986 30903 5042 30912
rect 5000 30734 5028 30903
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 4988 30728 5040 30734
rect 4988 30670 5040 30676
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 4802 30424 4858 30433
rect 4802 30359 4858 30368
rect 4816 30258 4844 30359
rect 4804 30252 4856 30258
rect 4804 30194 4856 30200
rect 4896 30184 4948 30190
rect 5000 30172 5028 30670
rect 5092 30394 5120 32710
rect 5184 31929 5212 33254
rect 5816 33040 5868 33046
rect 5816 32982 5868 32988
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 5552 32881 5580 32914
rect 5632 32904 5684 32910
rect 5538 32872 5594 32881
rect 5632 32846 5684 32852
rect 5724 32904 5776 32910
rect 5724 32846 5776 32852
rect 5538 32807 5594 32816
rect 5552 32502 5580 32807
rect 5540 32496 5592 32502
rect 5446 32464 5502 32473
rect 5540 32438 5592 32444
rect 5446 32399 5502 32408
rect 5460 32366 5488 32399
rect 5264 32360 5316 32366
rect 5264 32302 5316 32308
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 5170 31920 5226 31929
rect 5170 31855 5226 31864
rect 5276 31872 5304 32302
rect 5356 32224 5408 32230
rect 5540 32224 5592 32230
rect 5408 32184 5488 32212
rect 5356 32166 5408 32172
rect 5276 31844 5396 31872
rect 5264 31748 5316 31754
rect 5264 31690 5316 31696
rect 5172 31680 5224 31686
rect 5172 31622 5224 31628
rect 5080 30388 5132 30394
rect 5080 30330 5132 30336
rect 5080 30252 5132 30258
rect 5080 30194 5132 30200
rect 4948 30144 5028 30172
rect 4896 30126 4948 30132
rect 4712 30116 4764 30122
rect 4712 30058 4764 30064
rect 4804 30116 4856 30122
rect 4804 30058 4856 30064
rect 4252 30048 4304 30054
rect 4252 29990 4304 29996
rect 4264 28626 4292 29990
rect 4322 29948 4630 29957
rect 4322 29946 4328 29948
rect 4384 29946 4408 29948
rect 4464 29946 4488 29948
rect 4544 29946 4568 29948
rect 4624 29946 4630 29948
rect 4384 29894 4386 29946
rect 4566 29894 4568 29946
rect 4322 29892 4328 29894
rect 4384 29892 4408 29894
rect 4464 29892 4488 29894
rect 4544 29892 4568 29894
rect 4624 29892 4630 29894
rect 4322 29883 4630 29892
rect 4816 29850 4844 30058
rect 4804 29844 4856 29850
rect 4804 29786 4856 29792
rect 4344 29776 4396 29782
rect 4344 29718 4396 29724
rect 4710 29744 4766 29753
rect 4356 28966 4384 29718
rect 4710 29679 4766 29688
rect 4724 29646 4752 29679
rect 4712 29640 4764 29646
rect 4712 29582 4764 29588
rect 4620 29232 4672 29238
rect 4618 29200 4620 29209
rect 4672 29200 4674 29209
rect 4618 29135 4674 29144
rect 4344 28960 4396 28966
rect 4344 28902 4396 28908
rect 4322 28860 4630 28869
rect 4322 28858 4328 28860
rect 4384 28858 4408 28860
rect 4464 28858 4488 28860
rect 4544 28858 4568 28860
rect 4624 28858 4630 28860
rect 4384 28806 4386 28858
rect 4566 28806 4568 28858
rect 4322 28804 4328 28806
rect 4384 28804 4408 28806
rect 4464 28804 4488 28806
rect 4544 28804 4568 28806
rect 4624 28804 4630 28806
rect 4322 28795 4630 28804
rect 4252 28620 4304 28626
rect 4252 28562 4304 28568
rect 4620 28620 4672 28626
rect 4620 28562 4672 28568
rect 4436 28552 4488 28558
rect 4436 28494 4488 28500
rect 4252 28484 4304 28490
rect 4252 28426 4304 28432
rect 4264 27606 4292 28426
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 4356 28014 4384 28358
rect 4448 28218 4476 28494
rect 4528 28416 4580 28422
rect 4528 28358 4580 28364
rect 4436 28212 4488 28218
rect 4436 28154 4488 28160
rect 4344 28008 4396 28014
rect 4344 27950 4396 27956
rect 4540 27878 4568 28358
rect 4632 27985 4660 28562
rect 4724 28472 4752 29582
rect 4816 28966 4844 29786
rect 4908 29714 4936 30126
rect 4896 29708 4948 29714
rect 4896 29650 4948 29656
rect 5092 29594 5120 30194
rect 5184 30122 5212 31622
rect 5276 31521 5304 31690
rect 5262 31512 5318 31521
rect 5262 31447 5318 31456
rect 5264 31340 5316 31346
rect 5264 31282 5316 31288
rect 5276 30394 5304 31282
rect 5368 31210 5396 31844
rect 5356 31204 5408 31210
rect 5460 31192 5488 32184
rect 5540 32166 5592 32172
rect 5552 32026 5580 32166
rect 5540 32020 5592 32026
rect 5540 31962 5592 31968
rect 5540 31748 5592 31754
rect 5540 31690 5592 31696
rect 5552 31346 5580 31690
rect 5644 31482 5672 32846
rect 5736 31958 5764 32846
rect 5828 32434 5856 32982
rect 5920 32978 5948 33918
rect 6366 33895 6422 33904
rect 6000 33856 6052 33862
rect 6000 33798 6052 33804
rect 6012 33386 6040 33798
rect 6564 33454 6592 34342
rect 6276 33448 6328 33454
rect 6276 33390 6328 33396
rect 6368 33448 6420 33454
rect 6552 33448 6604 33454
rect 6420 33408 6500 33436
rect 6368 33390 6420 33396
rect 6000 33380 6052 33386
rect 6000 33322 6052 33328
rect 5908 32972 5960 32978
rect 5960 32932 6224 32960
rect 5908 32914 5960 32920
rect 6000 32836 6052 32842
rect 6000 32778 6052 32784
rect 5908 32768 5960 32774
rect 5906 32736 5908 32745
rect 5960 32736 5962 32745
rect 5906 32671 5962 32680
rect 5908 32564 5960 32570
rect 5908 32506 5960 32512
rect 5816 32428 5868 32434
rect 5816 32370 5868 32376
rect 5920 32337 5948 32506
rect 5906 32328 5962 32337
rect 5816 32292 5868 32298
rect 5906 32263 5962 32272
rect 5816 32234 5868 32240
rect 5828 31958 5856 32234
rect 5906 32056 5962 32065
rect 5906 31991 5962 32000
rect 5724 31952 5776 31958
rect 5724 31894 5776 31900
rect 5816 31952 5868 31958
rect 5816 31894 5868 31900
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 5540 31204 5592 31210
rect 5460 31164 5540 31192
rect 5356 31146 5408 31152
rect 5540 31146 5592 31152
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5356 30796 5408 30802
rect 5356 30738 5408 30744
rect 5540 30796 5592 30802
rect 5540 30738 5592 30744
rect 5264 30388 5316 30394
rect 5264 30330 5316 30336
rect 5368 30258 5396 30738
rect 5552 30326 5580 30738
rect 5644 30666 5672 31078
rect 5736 30938 5764 31894
rect 5816 31816 5868 31822
rect 5816 31758 5868 31764
rect 5828 31192 5856 31758
rect 5920 31521 5948 31991
rect 6012 31804 6040 32778
rect 6196 32722 6224 32932
rect 6288 32745 6316 33390
rect 6368 33312 6420 33318
rect 6368 33254 6420 33260
rect 6380 32910 6408 33254
rect 6368 32904 6420 32910
rect 6368 32846 6420 32852
rect 6472 32756 6500 33408
rect 6552 33390 6604 33396
rect 6564 32842 6592 33390
rect 6748 33153 6776 35663
rect 6840 35154 6868 37567
rect 6932 37466 6960 37760
rect 6920 37460 6972 37466
rect 6920 37402 6972 37408
rect 6920 37256 6972 37262
rect 6920 37198 6972 37204
rect 6932 36582 6960 37198
rect 7024 37194 7052 38354
rect 7116 38282 7144 38694
rect 7300 38418 7328 38830
rect 7392 38486 7420 39578
rect 7484 39506 7512 41239
rect 7576 39506 7604 41262
rect 7852 40730 7880 41618
rect 8022 41576 8078 41585
rect 8022 41511 8078 41520
rect 7932 40996 7984 41002
rect 7932 40938 7984 40944
rect 7944 40730 7972 40938
rect 7840 40724 7892 40730
rect 7840 40666 7892 40672
rect 7932 40724 7984 40730
rect 7932 40666 7984 40672
rect 8036 40390 8064 41511
rect 8024 40384 8076 40390
rect 8024 40326 8076 40332
rect 8220 40186 8248 41958
rect 8312 41177 8340 43500
rect 10520 42838 10548 43590
rect 10722 43004 11030 43013
rect 10722 43002 10728 43004
rect 10784 43002 10808 43004
rect 10864 43002 10888 43004
rect 10944 43002 10968 43004
rect 11024 43002 11030 43004
rect 10784 42950 10786 43002
rect 10966 42950 10968 43002
rect 10722 42948 10728 42950
rect 10784 42948 10808 42950
rect 10864 42948 10888 42950
rect 10944 42948 10968 42950
rect 11024 42948 11030 42950
rect 10722 42939 11030 42948
rect 10324 42832 10376 42838
rect 10508 42832 10560 42838
rect 10376 42792 10456 42820
rect 10324 42774 10376 42780
rect 8392 42764 8444 42770
rect 8392 42706 8444 42712
rect 8484 42764 8536 42770
rect 8484 42706 8536 42712
rect 8668 42764 8720 42770
rect 8668 42706 8720 42712
rect 8852 42764 8904 42770
rect 8852 42706 8904 42712
rect 9220 42764 9272 42770
rect 9220 42706 9272 42712
rect 8404 42362 8432 42706
rect 8392 42356 8444 42362
rect 8392 42298 8444 42304
rect 8392 42152 8444 42158
rect 8392 42094 8444 42100
rect 8404 41818 8432 42094
rect 8392 41812 8444 41818
rect 8392 41754 8444 41760
rect 8392 41676 8444 41682
rect 8392 41618 8444 41624
rect 8404 41313 8432 41618
rect 8390 41304 8446 41313
rect 8496 41274 8524 42706
rect 8680 42362 8708 42706
rect 8668 42356 8720 42362
rect 8668 42298 8720 42304
rect 8668 42084 8720 42090
rect 8668 42026 8720 42032
rect 8576 41472 8628 41478
rect 8576 41414 8628 41420
rect 8390 41239 8446 41248
rect 8484 41268 8536 41274
rect 8484 41210 8536 41216
rect 8588 41206 8616 41414
rect 8576 41200 8628 41206
rect 8298 41168 8354 41177
rect 8576 41142 8628 41148
rect 8298 41103 8354 41112
rect 8300 41064 8352 41070
rect 8300 41006 8352 41012
rect 8392 41064 8444 41070
rect 8392 41006 8444 41012
rect 8576 41064 8628 41070
rect 8576 41006 8628 41012
rect 8312 40769 8340 41006
rect 8298 40760 8354 40769
rect 8298 40695 8354 40704
rect 8404 40662 8432 41006
rect 8484 40724 8536 40730
rect 8484 40666 8536 40672
rect 8392 40656 8444 40662
rect 8392 40598 8444 40604
rect 8496 40594 8524 40666
rect 8300 40588 8352 40594
rect 8300 40530 8352 40536
rect 8484 40588 8536 40594
rect 8484 40530 8536 40536
rect 8312 40186 8340 40530
rect 8392 40520 8444 40526
rect 8392 40462 8444 40468
rect 8208 40180 8260 40186
rect 8208 40122 8260 40128
rect 8300 40180 8352 40186
rect 8300 40122 8352 40128
rect 8024 40112 8076 40118
rect 8024 40054 8076 40060
rect 7840 39976 7892 39982
rect 7840 39918 7892 39924
rect 7472 39500 7524 39506
rect 7472 39442 7524 39448
rect 7564 39500 7616 39506
rect 7748 39500 7800 39506
rect 7564 39442 7616 39448
rect 7668 39460 7748 39488
rect 7576 39001 7604 39442
rect 7668 39137 7696 39460
rect 7748 39442 7800 39448
rect 7654 39128 7710 39137
rect 7654 39063 7710 39072
rect 7562 38992 7618 39001
rect 7562 38927 7618 38936
rect 7472 38888 7524 38894
rect 7472 38830 7524 38836
rect 7564 38888 7616 38894
rect 7564 38830 7616 38836
rect 7484 38554 7512 38830
rect 7472 38548 7524 38554
rect 7472 38490 7524 38496
rect 7380 38480 7432 38486
rect 7380 38422 7432 38428
rect 7470 38448 7526 38457
rect 7288 38412 7340 38418
rect 7470 38383 7526 38392
rect 7288 38354 7340 38360
rect 7378 38312 7434 38321
rect 7104 38276 7156 38282
rect 7378 38247 7434 38256
rect 7104 38218 7156 38224
rect 7288 38208 7340 38214
rect 7288 38150 7340 38156
rect 7104 37868 7156 37874
rect 7156 37828 7236 37856
rect 7104 37810 7156 37816
rect 7208 37398 7236 37828
rect 7196 37392 7248 37398
rect 7196 37334 7248 37340
rect 7012 37188 7064 37194
rect 7012 37130 7064 37136
rect 7208 36718 7236 37334
rect 7196 36712 7248 36718
rect 7196 36654 7248 36660
rect 7104 36644 7156 36650
rect 7104 36586 7156 36592
rect 6920 36576 6972 36582
rect 6920 36518 6972 36524
rect 6932 36038 6960 36518
rect 7116 36038 7144 36586
rect 7194 36544 7250 36553
rect 7194 36479 7250 36488
rect 6920 36032 6972 36038
rect 6920 35974 6972 35980
rect 7104 36032 7156 36038
rect 7104 35974 7156 35980
rect 6920 35284 6972 35290
rect 6920 35226 6972 35232
rect 6828 35148 6880 35154
rect 6828 35090 6880 35096
rect 6932 34542 6960 35226
rect 7208 35222 7236 36479
rect 7300 35834 7328 38150
rect 7392 37330 7420 38247
rect 7484 38214 7512 38383
rect 7472 38208 7524 38214
rect 7472 38150 7524 38156
rect 7576 38010 7604 38830
rect 7668 38457 7696 39063
rect 7748 38888 7800 38894
rect 7748 38830 7800 38836
rect 7760 38554 7788 38830
rect 7852 38593 7880 39918
rect 7932 38888 7984 38894
rect 7932 38830 7984 38836
rect 7838 38584 7894 38593
rect 7748 38548 7800 38554
rect 7838 38519 7894 38528
rect 7748 38490 7800 38496
rect 7654 38448 7710 38457
rect 7838 38448 7894 38457
rect 7654 38383 7710 38392
rect 7748 38412 7800 38418
rect 7838 38383 7894 38392
rect 7748 38354 7800 38360
rect 7656 38208 7708 38214
rect 7760 38185 7788 38354
rect 7656 38150 7708 38156
rect 7746 38176 7802 38185
rect 7564 38004 7616 38010
rect 7564 37946 7616 37952
rect 7668 37330 7696 38150
rect 7746 38111 7802 38120
rect 7748 37936 7800 37942
rect 7748 37878 7800 37884
rect 7760 37777 7788 37878
rect 7746 37768 7802 37777
rect 7746 37703 7802 37712
rect 7852 37618 7880 38383
rect 7944 38010 7972 38830
rect 8036 38418 8064 40054
rect 8404 39982 8432 40462
rect 8588 40390 8616 41006
rect 8680 40730 8708 42026
rect 8758 41576 8814 41585
rect 8758 41511 8760 41520
rect 8812 41511 8814 41520
rect 8760 41482 8812 41488
rect 8864 41414 8892 42706
rect 9036 42560 9088 42566
rect 9036 42502 9088 42508
rect 9048 41750 9076 42502
rect 9128 42356 9180 42362
rect 9128 42298 9180 42304
rect 9036 41744 9088 41750
rect 9036 41686 9088 41692
rect 8772 41386 8892 41414
rect 8772 41313 8800 41386
rect 8758 41304 8814 41313
rect 9048 41274 9076 41686
rect 8758 41239 8814 41248
rect 8852 41268 8904 41274
rect 8852 41210 8904 41216
rect 9036 41268 9088 41274
rect 9036 41210 9088 41216
rect 8864 41070 8892 41210
rect 8760 41064 8812 41070
rect 8760 41006 8812 41012
rect 8852 41064 8904 41070
rect 8852 41006 8904 41012
rect 8668 40724 8720 40730
rect 8668 40666 8720 40672
rect 8666 40624 8722 40633
rect 8666 40559 8668 40568
rect 8720 40559 8722 40568
rect 8668 40530 8720 40536
rect 8576 40384 8628 40390
rect 8576 40326 8628 40332
rect 8576 40044 8628 40050
rect 8680 40032 8708 40530
rect 8772 40225 8800 41006
rect 8758 40216 8814 40225
rect 8864 40186 8892 41006
rect 9140 40746 9168 42298
rect 9232 41682 9260 42706
rect 9772 42628 9824 42634
rect 9772 42570 9824 42576
rect 9680 42220 9732 42226
rect 9680 42162 9732 42168
rect 9496 41744 9548 41750
rect 9496 41686 9548 41692
rect 9220 41676 9272 41682
rect 9220 41618 9272 41624
rect 9232 41070 9260 41618
rect 9220 41064 9272 41070
rect 9220 41006 9272 41012
rect 9404 41064 9456 41070
rect 9508 41052 9536 41686
rect 9692 41426 9720 42162
rect 9784 42022 9812 42570
rect 10062 42460 10370 42469
rect 10062 42458 10068 42460
rect 10124 42458 10148 42460
rect 10204 42458 10228 42460
rect 10284 42458 10308 42460
rect 10364 42458 10370 42460
rect 10124 42406 10126 42458
rect 10306 42406 10308 42458
rect 10062 42404 10068 42406
rect 10124 42404 10148 42406
rect 10204 42404 10228 42406
rect 10284 42404 10308 42406
rect 10364 42404 10370 42406
rect 10062 42395 10370 42404
rect 9772 42016 9824 42022
rect 9772 41958 9824 41964
rect 9956 42016 10008 42022
rect 9956 41958 10008 41964
rect 9784 41818 9812 41958
rect 9772 41812 9824 41818
rect 9772 41754 9824 41760
rect 9772 41676 9824 41682
rect 9772 41618 9824 41624
rect 9456 41024 9536 41052
rect 9404 41006 9456 41012
rect 8944 40724 8996 40730
rect 9140 40718 9260 40746
rect 8944 40666 8996 40672
rect 8956 40594 8984 40666
rect 9128 40656 9180 40662
rect 9128 40598 9180 40604
rect 8944 40588 8996 40594
rect 8944 40530 8996 40536
rect 9036 40384 9088 40390
rect 9140 40372 9168 40598
rect 9088 40344 9168 40372
rect 9036 40326 9088 40332
rect 8758 40151 8814 40160
rect 8852 40180 8904 40186
rect 8852 40122 8904 40128
rect 8628 40004 8708 40032
rect 8758 40080 8814 40089
rect 8758 40015 8814 40024
rect 8576 39986 8628 39992
rect 8392 39976 8444 39982
rect 8114 39944 8170 39953
rect 8392 39918 8444 39924
rect 8772 39914 8800 40015
rect 8114 39879 8170 39888
rect 8668 39908 8720 39914
rect 8128 39846 8156 39879
rect 8668 39850 8720 39856
rect 8760 39908 8812 39914
rect 8760 39850 8812 39856
rect 8116 39840 8168 39846
rect 8116 39782 8168 39788
rect 8484 39840 8536 39846
rect 8484 39782 8536 39788
rect 8576 39840 8628 39846
rect 8576 39782 8628 39788
rect 8208 39500 8260 39506
rect 8128 39460 8208 39488
rect 8024 38412 8076 38418
rect 8024 38354 8076 38360
rect 7932 38004 7984 38010
rect 7932 37946 7984 37952
rect 7760 37590 7880 37618
rect 7380 37324 7432 37330
rect 7380 37266 7432 37272
rect 7656 37324 7708 37330
rect 7656 37266 7708 37272
rect 7470 37224 7526 37233
rect 7380 37188 7432 37194
rect 7470 37159 7526 37168
rect 7380 37130 7432 37136
rect 7392 36854 7420 37130
rect 7380 36848 7432 36854
rect 7380 36790 7432 36796
rect 7484 36122 7512 37159
rect 7760 36666 7788 37590
rect 7840 37460 7892 37466
rect 7840 37402 7892 37408
rect 7668 36638 7788 36666
rect 7564 36576 7616 36582
rect 7564 36518 7616 36524
rect 7392 36094 7512 36122
rect 7392 35873 7420 36094
rect 7472 36032 7524 36038
rect 7472 35974 7524 35980
rect 7378 35864 7434 35873
rect 7288 35828 7340 35834
rect 7378 35799 7434 35808
rect 7288 35770 7340 35776
rect 7484 35272 7512 35974
rect 7300 35244 7512 35272
rect 7196 35216 7248 35222
rect 7196 35158 7248 35164
rect 7300 34542 7328 35244
rect 7380 35148 7432 35154
rect 7380 35090 7432 35096
rect 7472 35148 7524 35154
rect 7472 35090 7524 35096
rect 7392 34542 7420 35090
rect 6920 34536 6972 34542
rect 6920 34478 6972 34484
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 7380 34536 7432 34542
rect 7380 34478 7432 34484
rect 7104 34060 7156 34066
rect 7104 34002 7156 34008
rect 6828 33856 6880 33862
rect 6828 33798 6880 33804
rect 6920 33856 6972 33862
rect 6920 33798 6972 33804
rect 6734 33144 6790 33153
rect 6840 33114 6868 33798
rect 6932 33658 6960 33798
rect 6920 33652 6972 33658
rect 6920 33594 6972 33600
rect 7116 33454 7144 34002
rect 7194 33960 7250 33969
rect 7194 33895 7250 33904
rect 7104 33448 7156 33454
rect 7104 33390 7156 33396
rect 7104 33312 7156 33318
rect 7104 33254 7156 33260
rect 6734 33079 6736 33088
rect 6788 33079 6790 33088
rect 6828 33108 6880 33114
rect 6736 33050 6788 33056
rect 6828 33050 6880 33056
rect 6828 32972 6880 32978
rect 6828 32914 6880 32920
rect 7012 32972 7064 32978
rect 7012 32914 7064 32920
rect 6736 32904 6788 32910
rect 6656 32864 6736 32892
rect 6552 32836 6604 32842
rect 6552 32778 6604 32784
rect 6104 32694 6224 32722
rect 6274 32736 6330 32745
rect 6104 32570 6132 32694
rect 6274 32671 6330 32680
rect 6380 32728 6500 32756
rect 6182 32600 6238 32609
rect 6092 32564 6144 32570
rect 6182 32535 6238 32544
rect 6092 32506 6144 32512
rect 6104 32065 6132 32506
rect 6196 32434 6224 32535
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 6276 32360 6328 32366
rect 6276 32302 6328 32308
rect 6184 32292 6236 32298
rect 6184 32234 6236 32240
rect 6090 32056 6146 32065
rect 6090 31991 6146 32000
rect 6092 31952 6144 31958
rect 6090 31920 6092 31929
rect 6144 31920 6146 31929
rect 6090 31855 6146 31864
rect 6092 31816 6144 31822
rect 6012 31776 6092 31804
rect 6092 31758 6144 31764
rect 5906 31512 5962 31521
rect 5962 31456 6040 31464
rect 5906 31447 5908 31456
rect 5960 31436 6040 31456
rect 5908 31418 5960 31424
rect 5908 31204 5960 31210
rect 5828 31164 5908 31192
rect 5908 31146 5960 31152
rect 5814 30968 5870 30977
rect 5724 30932 5776 30938
rect 5814 30903 5870 30912
rect 5724 30874 5776 30880
rect 5632 30660 5684 30666
rect 5632 30602 5684 30608
rect 5540 30320 5592 30326
rect 5540 30262 5592 30268
rect 5356 30252 5408 30258
rect 5356 30194 5408 30200
rect 5644 30138 5672 30602
rect 5736 30274 5764 30874
rect 5828 30802 5856 30903
rect 5816 30796 5868 30802
rect 5816 30738 5868 30744
rect 5920 30705 5948 31146
rect 5906 30696 5962 30705
rect 5906 30631 5962 30640
rect 5906 30560 5962 30569
rect 5906 30495 5962 30504
rect 5814 30424 5870 30433
rect 5814 30359 5816 30368
rect 5868 30359 5870 30368
rect 5816 30330 5868 30336
rect 5736 30246 5856 30274
rect 5172 30116 5224 30122
rect 5172 30058 5224 30064
rect 5460 30110 5672 30138
rect 5724 30184 5776 30190
rect 5724 30126 5776 30132
rect 5460 29850 5488 30110
rect 5540 30048 5592 30054
rect 5540 29990 5592 29996
rect 5448 29844 5500 29850
rect 5448 29786 5500 29792
rect 5356 29708 5408 29714
rect 5356 29650 5408 29656
rect 5092 29566 5212 29594
rect 4988 29504 5040 29510
rect 4988 29446 5040 29452
rect 5080 29504 5132 29510
rect 5080 29446 5132 29452
rect 4804 28960 4856 28966
rect 4804 28902 4856 28908
rect 4896 28960 4948 28966
rect 5000 28937 5028 29446
rect 5092 29238 5120 29446
rect 5080 29232 5132 29238
rect 5080 29174 5132 29180
rect 5080 28960 5132 28966
rect 4896 28902 4948 28908
rect 4986 28928 5042 28937
rect 4816 28540 4844 28902
rect 4908 28694 4936 28902
rect 5080 28902 5132 28908
rect 4986 28863 5042 28872
rect 4986 28792 5042 28801
rect 4986 28727 5042 28736
rect 4896 28688 4948 28694
rect 4896 28630 4948 28636
rect 5000 28558 5028 28727
rect 4988 28552 5040 28558
rect 4816 28512 4936 28540
rect 4724 28444 4844 28472
rect 4816 28121 4844 28444
rect 4802 28112 4858 28121
rect 4802 28047 4804 28056
rect 4856 28047 4858 28056
rect 4804 28018 4856 28024
rect 4908 28014 4936 28512
rect 4988 28494 5040 28500
rect 4986 28112 5042 28121
rect 4986 28047 5042 28056
rect 4712 28008 4764 28014
rect 4618 27976 4674 27985
rect 4712 27950 4764 27956
rect 4896 28008 4948 28014
rect 4896 27950 4948 27956
rect 4618 27911 4674 27920
rect 4528 27872 4580 27878
rect 4528 27814 4580 27820
rect 4322 27772 4630 27781
rect 4322 27770 4328 27772
rect 4384 27770 4408 27772
rect 4464 27770 4488 27772
rect 4544 27770 4568 27772
rect 4624 27770 4630 27772
rect 4384 27718 4386 27770
rect 4566 27718 4568 27770
rect 4322 27716 4328 27718
rect 4384 27716 4408 27718
rect 4464 27716 4488 27718
rect 4544 27716 4568 27718
rect 4624 27716 4630 27718
rect 4322 27707 4630 27716
rect 4252 27600 4304 27606
rect 4620 27600 4672 27606
rect 4252 27542 4304 27548
rect 4526 27568 4582 27577
rect 4028 27492 4200 27520
rect 4620 27542 4672 27548
rect 4526 27503 4582 27512
rect 3976 27474 4028 27480
rect 3516 27464 3568 27470
rect 3514 27432 3516 27441
rect 3568 27432 3570 27441
rect 3514 27367 3570 27376
rect 3662 27228 3970 27237
rect 3662 27226 3668 27228
rect 3724 27226 3748 27228
rect 3804 27226 3828 27228
rect 3884 27226 3908 27228
rect 3964 27226 3970 27228
rect 3724 27174 3726 27226
rect 3906 27174 3908 27226
rect 3662 27172 3668 27174
rect 3724 27172 3748 27174
rect 3804 27172 3828 27174
rect 3884 27172 3908 27174
rect 3964 27172 3970 27174
rect 3662 27163 3970 27172
rect 3424 27124 3476 27130
rect 3424 27066 3476 27072
rect 3330 27024 3386 27033
rect 3330 26959 3386 26968
rect 3330 26480 3386 26489
rect 3330 26415 3386 26424
rect 3240 25968 3292 25974
rect 3240 25910 3292 25916
rect 3240 25696 3292 25702
rect 3240 25638 3292 25644
rect 3054 21655 3110 21664
rect 3148 21684 3200 21690
rect 3068 21350 3096 21655
rect 3148 21626 3200 21632
rect 3148 21480 3200 21486
rect 3146 21448 3148 21457
rect 3200 21448 3202 21457
rect 3146 21383 3202 21392
rect 3056 21344 3108 21350
rect 3252 21332 3280 25638
rect 3344 24750 3372 26415
rect 3436 25906 3464 27066
rect 4080 27062 4108 27492
rect 4160 27328 4212 27334
rect 4160 27270 4212 27276
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3528 26042 3556 26930
rect 3608 26920 3660 26926
rect 3608 26862 3660 26868
rect 4068 26920 4120 26926
rect 4068 26862 4120 26868
rect 3620 26246 3648 26862
rect 3700 26852 3752 26858
rect 3700 26794 3752 26800
rect 3712 26586 3740 26794
rect 4080 26761 4108 26862
rect 4066 26752 4122 26761
rect 4066 26687 4122 26696
rect 3790 26616 3846 26625
rect 3700 26580 3752 26586
rect 4080 26586 4108 26687
rect 4172 26625 4200 27270
rect 4342 27160 4398 27169
rect 4252 27124 4304 27130
rect 4342 27095 4398 27104
rect 4252 27066 4304 27072
rect 4158 26616 4214 26625
rect 3790 26551 3846 26560
rect 4068 26580 4120 26586
rect 3700 26522 3752 26528
rect 3804 26314 3832 26551
rect 4158 26551 4214 26560
rect 4068 26522 4120 26528
rect 3974 26480 4030 26489
rect 3974 26415 4030 26424
rect 3792 26308 3844 26314
rect 3988 26296 4016 26415
rect 3988 26268 4200 26296
rect 3792 26250 3844 26256
rect 3608 26240 3660 26246
rect 3608 26182 3660 26188
rect 3662 26140 3970 26149
rect 3662 26138 3668 26140
rect 3724 26138 3748 26140
rect 3804 26138 3828 26140
rect 3884 26138 3908 26140
rect 3964 26138 3970 26140
rect 3724 26086 3726 26138
rect 3906 26086 3908 26138
rect 3662 26084 3668 26086
rect 3724 26084 3748 26086
rect 3804 26084 3828 26086
rect 3884 26084 3908 26086
rect 3964 26084 3970 26086
rect 3662 26075 3970 26084
rect 3516 26036 3568 26042
rect 3516 25978 3568 25984
rect 3884 25968 3936 25974
rect 3514 25936 3570 25945
rect 3424 25900 3476 25906
rect 3698 25936 3754 25945
rect 3620 25906 3698 25922
rect 3514 25871 3570 25880
rect 3608 25900 3698 25906
rect 3424 25842 3476 25848
rect 3424 25356 3476 25362
rect 3424 25298 3476 25304
rect 3436 24954 3464 25298
rect 3424 24948 3476 24954
rect 3424 24890 3476 24896
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 3424 24744 3476 24750
rect 3528 24732 3556 25871
rect 3660 25894 3698 25900
rect 3884 25910 3936 25916
rect 3974 25936 4030 25945
rect 3698 25871 3754 25880
rect 3608 25842 3660 25848
rect 3896 25838 3924 25910
rect 3974 25871 4030 25880
rect 3792 25832 3844 25838
rect 3606 25800 3662 25809
rect 3792 25774 3844 25780
rect 3884 25832 3936 25838
rect 3884 25774 3936 25780
rect 3606 25735 3662 25744
rect 3620 25294 3648 25735
rect 3698 25664 3754 25673
rect 3698 25599 3754 25608
rect 3712 25430 3740 25599
rect 3700 25424 3752 25430
rect 3804 25401 3832 25774
rect 3884 25696 3936 25702
rect 3884 25638 3936 25644
rect 3700 25366 3752 25372
rect 3790 25392 3846 25401
rect 3790 25327 3846 25336
rect 3608 25288 3660 25294
rect 3700 25288 3752 25294
rect 3608 25230 3660 25236
rect 3698 25256 3700 25265
rect 3896 25265 3924 25638
rect 3988 25362 4016 25871
rect 4172 25820 4200 26268
rect 4264 26160 4292 27066
rect 4356 26926 4384 27095
rect 4540 26994 4568 27503
rect 4632 27418 4660 27542
rect 4724 27538 4752 27950
rect 4804 27940 4856 27946
rect 4804 27882 4856 27888
rect 4712 27532 4764 27538
rect 4712 27474 4764 27480
rect 4632 27390 4752 27418
rect 4618 27296 4674 27305
rect 4618 27231 4674 27240
rect 4528 26988 4580 26994
rect 4528 26930 4580 26936
rect 4344 26920 4396 26926
rect 4342 26888 4344 26897
rect 4396 26888 4398 26897
rect 4342 26823 4398 26832
rect 4632 26790 4660 27231
rect 4724 27130 4752 27390
rect 4712 27124 4764 27130
rect 4712 27066 4764 27072
rect 4712 26852 4764 26858
rect 4712 26794 4764 26800
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4322 26684 4630 26693
rect 4322 26682 4328 26684
rect 4384 26682 4408 26684
rect 4464 26682 4488 26684
rect 4544 26682 4568 26684
rect 4624 26682 4630 26684
rect 4384 26630 4386 26682
rect 4566 26630 4568 26682
rect 4322 26628 4328 26630
rect 4384 26628 4408 26630
rect 4464 26628 4488 26630
rect 4544 26628 4568 26630
rect 4624 26628 4630 26630
rect 4322 26619 4630 26628
rect 4724 26586 4752 26794
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 4712 26580 4764 26586
rect 4712 26522 4764 26528
rect 4528 26512 4580 26518
rect 4434 26480 4490 26489
rect 4528 26454 4580 26460
rect 4434 26415 4490 26424
rect 4264 26132 4384 26160
rect 4252 26036 4304 26042
rect 4252 25978 4304 25984
rect 4080 25792 4200 25820
rect 3976 25356 4028 25362
rect 3976 25298 4028 25304
rect 3752 25256 3754 25265
rect 3698 25191 3754 25200
rect 3882 25256 3938 25265
rect 3882 25191 3938 25200
rect 3662 25052 3970 25061
rect 3662 25050 3668 25052
rect 3724 25050 3748 25052
rect 3804 25050 3828 25052
rect 3884 25050 3908 25052
rect 3964 25050 3970 25052
rect 3724 24998 3726 25050
rect 3906 24998 3908 25050
rect 3662 24996 3668 24998
rect 3724 24996 3748 24998
rect 3804 24996 3828 24998
rect 3884 24996 3908 24998
rect 3964 24996 3970 24998
rect 3662 24987 3970 24996
rect 3976 24948 4028 24954
rect 3976 24890 4028 24896
rect 3700 24744 3752 24750
rect 3528 24704 3700 24732
rect 3424 24686 3476 24692
rect 3344 24342 3372 24686
rect 3332 24336 3384 24342
rect 3332 24278 3384 24284
rect 3344 24206 3372 24278
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 3344 23254 3372 24142
rect 3332 23248 3384 23254
rect 3332 23190 3384 23196
rect 3344 22438 3372 23190
rect 3436 23186 3464 24686
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3424 23180 3476 23186
rect 3424 23122 3476 23128
rect 3436 22574 3464 23122
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3332 22432 3384 22438
rect 3332 22374 3384 22380
rect 3436 22386 3464 22510
rect 3528 22506 3556 24210
rect 3620 24070 3648 24704
rect 3700 24686 3752 24692
rect 3884 24676 3936 24682
rect 3884 24618 3936 24624
rect 3896 24410 3924 24618
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3698 24304 3754 24313
rect 3698 24239 3754 24248
rect 3882 24304 3938 24313
rect 3882 24239 3938 24248
rect 3712 24206 3740 24239
rect 3700 24200 3752 24206
rect 3700 24142 3752 24148
rect 3896 24138 3924 24239
rect 3988 24138 4016 24890
rect 4080 24750 4108 25792
rect 4264 25752 4292 25978
rect 4172 25724 4292 25752
rect 4172 25673 4200 25724
rect 4356 25684 4384 26132
rect 4448 25770 4476 26415
rect 4540 26217 4568 26454
rect 4526 26208 4582 26217
rect 4526 26143 4582 26152
rect 4632 26081 4660 26522
rect 4724 26450 4752 26522
rect 4712 26444 4764 26450
rect 4712 26386 4764 26392
rect 4618 26072 4674 26081
rect 4618 26007 4674 26016
rect 4816 25888 4844 27882
rect 4908 26858 4936 27950
rect 5000 27606 5028 28047
rect 5092 27878 5120 28902
rect 5080 27872 5132 27878
rect 5080 27814 5132 27820
rect 4988 27600 5040 27606
rect 4988 27542 5040 27548
rect 5080 27532 5132 27538
rect 5080 27474 5132 27480
rect 4988 27328 5040 27334
rect 4988 27270 5040 27276
rect 4896 26852 4948 26858
rect 4896 26794 4948 26800
rect 4894 26752 4950 26761
rect 4894 26687 4950 26696
rect 4804 25860 4844 25888
rect 4712 25832 4764 25838
rect 4804 25786 4832 25860
rect 4764 25780 4832 25786
rect 4712 25774 4832 25780
rect 4436 25764 4488 25770
rect 4724 25758 4832 25774
rect 4908 25770 4936 26687
rect 5000 26160 5028 27270
rect 5092 26858 5120 27474
rect 5080 26852 5132 26858
rect 5080 26794 5132 26800
rect 5080 26444 5132 26450
rect 5080 26386 5132 26392
rect 5092 26353 5120 26386
rect 5078 26344 5134 26353
rect 5078 26279 5134 26288
rect 5000 26132 5120 26160
rect 4986 26072 5042 26081
rect 4986 26007 5042 26016
rect 5000 25974 5028 26007
rect 4988 25968 5040 25974
rect 4988 25910 5040 25916
rect 4988 25832 5040 25838
rect 5092 25820 5120 26132
rect 5040 25792 5120 25820
rect 4988 25774 5040 25780
rect 4896 25764 4948 25770
rect 4436 25706 4488 25712
rect 4896 25706 4948 25712
rect 4158 25664 4214 25673
rect 4158 25599 4214 25608
rect 4264 25656 4384 25684
rect 4804 25696 4856 25702
rect 4264 25480 4292 25656
rect 4804 25638 4856 25644
rect 4322 25596 4630 25605
rect 4322 25594 4328 25596
rect 4384 25594 4408 25596
rect 4464 25594 4488 25596
rect 4544 25594 4568 25596
rect 4624 25594 4630 25596
rect 4384 25542 4386 25594
rect 4566 25542 4568 25594
rect 4322 25540 4328 25542
rect 4384 25540 4408 25542
rect 4464 25540 4488 25542
rect 4544 25540 4568 25542
rect 4624 25540 4630 25542
rect 4322 25531 4630 25540
rect 4710 25528 4766 25537
rect 4620 25492 4672 25498
rect 4264 25452 4384 25480
rect 4160 25220 4212 25226
rect 4160 25162 4212 25168
rect 4172 24954 4200 25162
rect 4356 25140 4384 25452
rect 4540 25452 4620 25480
rect 4540 25344 4568 25452
rect 4816 25498 4844 25638
rect 5000 25537 5028 25774
rect 4986 25528 5042 25537
rect 4710 25463 4766 25472
rect 4804 25492 4856 25498
rect 4620 25434 4672 25440
rect 4524 25316 4568 25344
rect 4524 25208 4552 25316
rect 4620 25288 4672 25294
rect 4620 25230 4672 25236
rect 4524 25180 4568 25208
rect 4436 25152 4488 25158
rect 4356 25112 4436 25140
rect 4436 25094 4488 25100
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 4068 24744 4120 24750
rect 4068 24686 4120 24692
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4080 24342 4108 24686
rect 4068 24336 4120 24342
rect 4068 24278 4120 24284
rect 4068 24200 4120 24206
rect 4068 24142 4120 24148
rect 3884 24132 3936 24138
rect 3884 24074 3936 24080
rect 3976 24132 4028 24138
rect 3976 24074 4028 24080
rect 3608 24064 3660 24070
rect 3608 24006 3660 24012
rect 3662 23964 3970 23973
rect 3662 23962 3668 23964
rect 3724 23962 3748 23964
rect 3804 23962 3828 23964
rect 3884 23962 3908 23964
rect 3964 23962 3970 23964
rect 3724 23910 3726 23962
rect 3906 23910 3908 23962
rect 3662 23908 3668 23910
rect 3724 23908 3748 23910
rect 3804 23908 3828 23910
rect 3884 23908 3908 23910
rect 3964 23908 3970 23910
rect 3662 23899 3970 23908
rect 4080 23662 4108 24142
rect 3608 23656 3660 23662
rect 3606 23624 3608 23633
rect 4068 23656 4120 23662
rect 3660 23624 3662 23633
rect 4068 23598 4120 23604
rect 3606 23559 3662 23568
rect 3792 23520 3844 23526
rect 3792 23462 3844 23468
rect 3804 23186 3832 23462
rect 4080 23254 4108 23598
rect 4068 23248 4120 23254
rect 4068 23190 4120 23196
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3662 22876 3970 22885
rect 3662 22874 3668 22876
rect 3724 22874 3748 22876
rect 3804 22874 3828 22876
rect 3884 22874 3908 22876
rect 3964 22874 3970 22876
rect 3724 22822 3726 22874
rect 3906 22822 3908 22874
rect 3662 22820 3668 22822
rect 3724 22820 3748 22822
rect 3804 22820 3828 22822
rect 3884 22820 3908 22822
rect 3964 22820 3970 22822
rect 3662 22811 3970 22820
rect 4172 22692 4200 24686
rect 4540 24596 4568 25180
rect 4632 24818 4660 25230
rect 4724 24886 4752 25463
rect 4986 25463 5042 25472
rect 4804 25434 4856 25440
rect 5000 25378 5028 25463
rect 4816 25350 5028 25378
rect 4816 24954 4844 25350
rect 4896 25288 4948 25294
rect 4894 25256 4896 25265
rect 4948 25256 4950 25265
rect 4894 25191 4950 25200
rect 4988 25152 5040 25158
rect 4986 25120 4988 25129
rect 5040 25120 5042 25129
rect 4986 25055 5042 25064
rect 4894 24984 4950 24993
rect 4804 24948 4856 24954
rect 4894 24919 4950 24928
rect 4804 24890 4856 24896
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 4264 24568 4568 24596
rect 4264 22817 4292 24568
rect 4322 24508 4630 24517
rect 4322 24506 4328 24508
rect 4384 24506 4408 24508
rect 4464 24506 4488 24508
rect 4544 24506 4568 24508
rect 4624 24506 4630 24508
rect 4384 24454 4386 24506
rect 4566 24454 4568 24506
rect 4322 24452 4328 24454
rect 4384 24452 4408 24454
rect 4464 24452 4488 24454
rect 4544 24452 4568 24454
rect 4624 24452 4630 24454
rect 4322 24443 4630 24452
rect 4528 24404 4580 24410
rect 4528 24346 4580 24352
rect 4540 24070 4568 24346
rect 4724 24342 4752 24822
rect 4816 24750 4844 24890
rect 4804 24744 4856 24750
rect 4804 24686 4856 24692
rect 4712 24336 4764 24342
rect 4712 24278 4764 24284
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 4712 24132 4764 24138
rect 4712 24074 4764 24080
rect 4436 24064 4488 24070
rect 4436 24006 4488 24012
rect 4528 24064 4580 24070
rect 4528 24006 4580 24012
rect 4448 23594 4476 24006
rect 4436 23588 4488 23594
rect 4436 23530 4488 23536
rect 4322 23420 4630 23429
rect 4322 23418 4328 23420
rect 4384 23418 4408 23420
rect 4464 23418 4488 23420
rect 4544 23418 4568 23420
rect 4624 23418 4630 23420
rect 4384 23366 4386 23418
rect 4566 23366 4568 23418
rect 4322 23364 4328 23366
rect 4384 23364 4408 23366
rect 4464 23364 4488 23366
rect 4544 23364 4568 23366
rect 4624 23364 4630 23366
rect 4322 23355 4630 23364
rect 4434 23216 4490 23225
rect 4724 23186 4752 24074
rect 4816 24041 4844 24210
rect 4802 24032 4858 24041
rect 4802 23967 4858 23976
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4434 23151 4490 23160
rect 4620 23180 4672 23186
rect 4250 22808 4306 22817
rect 4448 22778 4476 23151
rect 4620 23122 4672 23128
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4528 23112 4580 23118
rect 4528 23054 4580 23060
rect 4250 22743 4306 22752
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 3790 22672 3846 22681
rect 3700 22636 3752 22642
rect 4172 22664 4384 22692
rect 3790 22607 3846 22616
rect 3700 22578 3752 22584
rect 3516 22500 3568 22506
rect 3516 22442 3568 22448
rect 3712 22386 3740 22578
rect 3436 22358 3740 22386
rect 3332 22228 3384 22234
rect 3332 22170 3384 22176
rect 3700 22228 3752 22234
rect 3700 22170 3752 22176
rect 3344 22098 3372 22170
rect 3712 22098 3740 22170
rect 3804 22098 3832 22607
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 4068 22432 4120 22438
rect 3882 22400 3938 22409
rect 4068 22374 4120 22380
rect 3882 22335 3938 22344
rect 3896 22098 3924 22335
rect 4080 22098 4108 22374
rect 4172 22166 4200 22510
rect 4252 22500 4304 22506
rect 4252 22442 4304 22448
rect 4160 22160 4212 22166
rect 4158 22128 4160 22137
rect 4212 22128 4214 22137
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 3792 22092 3844 22098
rect 3792 22034 3844 22040
rect 3884 22092 3936 22098
rect 3884 22034 3936 22040
rect 4068 22092 4120 22098
rect 4264 22098 4292 22442
rect 4356 22438 4384 22664
rect 4540 22642 4568 23054
rect 4528 22636 4580 22642
rect 4528 22578 4580 22584
rect 4632 22506 4660 23122
rect 4620 22500 4672 22506
rect 4620 22442 4672 22448
rect 4724 22438 4752 23122
rect 4816 23118 4844 23462
rect 4804 23112 4856 23118
rect 4804 23054 4856 23060
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4322 22332 4630 22341
rect 4322 22330 4328 22332
rect 4384 22330 4408 22332
rect 4464 22330 4488 22332
rect 4544 22330 4568 22332
rect 4624 22330 4630 22332
rect 4384 22278 4386 22330
rect 4566 22278 4568 22330
rect 4322 22276 4328 22278
rect 4384 22276 4408 22278
rect 4464 22276 4488 22278
rect 4544 22276 4568 22278
rect 4624 22276 4630 22278
rect 4322 22267 4630 22276
rect 4710 22264 4766 22273
rect 4436 22228 4488 22234
rect 4710 22199 4712 22208
rect 4436 22170 4488 22176
rect 4764 22199 4766 22208
rect 4712 22170 4764 22176
rect 4448 22137 4476 22170
rect 4434 22128 4490 22137
rect 4158 22063 4214 22072
rect 4252 22092 4304 22098
rect 4068 22034 4120 22040
rect 4816 22094 4844 23054
rect 4434 22063 4490 22072
rect 4540 22066 4844 22094
rect 4252 22034 4304 22040
rect 3804 21978 3832 22034
rect 4344 22024 4396 22030
rect 3424 21956 3476 21962
rect 3804 21950 4200 21978
rect 4344 21966 4396 21972
rect 3424 21898 3476 21904
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3344 21486 3372 21830
rect 3436 21690 3464 21898
rect 3662 21788 3970 21797
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3792 21616 3844 21622
rect 3792 21558 3844 21564
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 4066 21584 4122 21593
rect 3332 21480 3384 21486
rect 3608 21480 3660 21486
rect 3384 21440 3556 21468
rect 3332 21422 3384 21428
rect 3056 21286 3108 21292
rect 3160 21321 3280 21332
rect 3160 21312 3294 21321
rect 3160 21304 3238 21312
rect 2976 20998 3096 21026
rect 3160 21010 3188 21304
rect 3238 21247 3294 21256
rect 3330 21176 3386 21185
rect 3330 21111 3386 21120
rect 3344 21078 3372 21111
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 3332 21072 3384 21078
rect 3332 21014 3384 21020
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 2872 19984 2924 19990
rect 2778 19952 2834 19961
rect 2872 19926 2924 19932
rect 2778 19887 2780 19896
rect 2832 19887 2834 19896
rect 2780 19858 2832 19864
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2688 19440 2740 19446
rect 2688 19382 2740 19388
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2516 18834 2544 19246
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 2608 18766 2636 19314
rect 2700 18834 2728 19382
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2332 18108 2452 18136
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2240 17134 2268 17614
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2240 16590 2268 17070
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 1964 16046 1992 16526
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 2332 15910 2360 18108
rect 2410 18048 2466 18057
rect 2608 18034 2636 18702
rect 2410 17983 2466 17992
rect 2516 18006 2636 18034
rect 2424 16250 2452 17983
rect 2516 17678 2544 18006
rect 2792 17864 2820 19450
rect 2976 19360 3004 20878
rect 3068 19514 3096 20998
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3146 20904 3202 20913
rect 3146 20839 3148 20848
rect 3200 20839 3202 20848
rect 3148 20810 3200 20816
rect 3252 20058 3280 21014
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3332 20868 3384 20874
rect 3332 20810 3384 20816
rect 3344 20777 3372 20810
rect 3330 20768 3386 20777
rect 3330 20703 3386 20712
rect 3330 20632 3386 20641
rect 3330 20567 3386 20576
rect 3344 20330 3372 20567
rect 3436 20534 3464 20946
rect 3528 20602 3556 21440
rect 3608 21422 3660 21428
rect 3620 21010 3648 21422
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3712 21010 3740 21286
rect 3804 21078 3832 21558
rect 3988 21486 4016 21558
rect 4066 21519 4122 21528
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 4080 21418 4108 21519
rect 3884 21412 3936 21418
rect 3884 21354 3936 21360
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 3792 21072 3844 21078
rect 3792 21014 3844 21020
rect 3896 21010 3924 21354
rect 4066 21312 4122 21321
rect 4066 21247 4122 21256
rect 4080 21010 4108 21247
rect 3608 21004 3660 21010
rect 3608 20946 3660 20952
rect 3700 21004 3752 21010
rect 3700 20946 3752 20952
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 4066 20496 4122 20505
rect 3332 20324 3384 20330
rect 3332 20266 3384 20272
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 2884 19332 3004 19360
rect 2884 18902 2912 19332
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 2872 18896 2924 18902
rect 2872 18838 2924 18844
rect 2884 18714 2912 18838
rect 3068 18834 3096 19110
rect 3160 18873 3188 19858
rect 3240 19848 3292 19854
rect 3238 19816 3240 19825
rect 3292 19816 3294 19825
rect 3238 19751 3294 19760
rect 3238 19408 3294 19417
rect 3344 19378 3372 19994
rect 3436 19394 3464 20470
rect 4066 20431 4122 20440
rect 4080 20398 4108 20431
rect 3700 20392 3752 20398
rect 3700 20334 3752 20340
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 3516 20256 3568 20262
rect 3516 20198 3568 20204
rect 3528 19514 3556 20198
rect 3712 20058 3740 20334
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 3700 20052 3752 20058
rect 3700 19994 3752 20000
rect 3988 19990 4016 20266
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 4172 19922 4200 21950
rect 4252 21888 4304 21894
rect 4356 21865 4384 21966
rect 4252 21830 4304 21836
rect 4342 21856 4398 21865
rect 4264 20942 4292 21830
rect 4342 21791 4398 21800
rect 4342 21720 4398 21729
rect 4342 21655 4344 21664
rect 4396 21655 4398 21664
rect 4344 21626 4396 21632
rect 4436 21616 4488 21622
rect 4342 21584 4398 21593
rect 4540 21604 4568 22066
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4488 21576 4568 21604
rect 4436 21558 4488 21564
rect 4342 21519 4398 21528
rect 4356 21486 4384 21519
rect 4344 21480 4396 21486
rect 4344 21422 4396 21428
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 4724 21146 4752 21966
rect 4908 21842 4936 24919
rect 4988 24880 5040 24886
rect 4988 24822 5040 24828
rect 5000 24614 5028 24822
rect 4988 24608 5040 24614
rect 4988 24550 5040 24556
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 5092 24449 5120 24550
rect 5078 24440 5134 24449
rect 5078 24375 5134 24384
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 5000 23254 5028 24142
rect 5080 24064 5132 24070
rect 5080 24006 5132 24012
rect 5092 23866 5120 24006
rect 5080 23860 5132 23866
rect 5080 23802 5132 23808
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4988 23248 5040 23254
rect 4988 23190 5040 23196
rect 5092 23186 5120 23598
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 5080 22976 5132 22982
rect 5080 22918 5132 22924
rect 5092 22817 5120 22918
rect 5078 22808 5134 22817
rect 5078 22743 5134 22752
rect 5184 22624 5212 29566
rect 5262 29336 5318 29345
rect 5262 29271 5318 29280
rect 5276 27402 5304 29271
rect 5368 27538 5396 29650
rect 5460 29034 5488 29786
rect 5552 29102 5580 29990
rect 5630 29880 5686 29889
rect 5630 29815 5632 29824
rect 5684 29815 5686 29824
rect 5632 29786 5684 29792
rect 5632 29708 5684 29714
rect 5632 29650 5684 29656
rect 5644 29170 5672 29650
rect 5736 29617 5764 30126
rect 5722 29608 5778 29617
rect 5722 29543 5778 29552
rect 5724 29504 5776 29510
rect 5724 29446 5776 29452
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 5540 29096 5592 29102
rect 5540 29038 5592 29044
rect 5448 29028 5500 29034
rect 5448 28970 5500 28976
rect 5552 28994 5580 29038
rect 5552 28966 5672 28994
rect 5446 28656 5502 28665
rect 5446 28591 5448 28600
rect 5500 28591 5502 28600
rect 5448 28562 5500 28568
rect 5538 28520 5594 28529
rect 5538 28455 5594 28464
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5460 27606 5488 28358
rect 5448 27600 5500 27606
rect 5448 27542 5500 27548
rect 5356 27532 5408 27538
rect 5356 27474 5408 27480
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5264 27396 5316 27402
rect 5264 27338 5316 27344
rect 5356 27396 5408 27402
rect 5356 27338 5408 27344
rect 5368 26586 5396 27338
rect 5264 26580 5316 26586
rect 5264 26522 5316 26528
rect 5356 26580 5408 26586
rect 5356 26522 5408 26528
rect 5276 25945 5304 26522
rect 5356 26444 5408 26450
rect 5356 26386 5408 26392
rect 5368 26081 5396 26386
rect 5354 26072 5410 26081
rect 5354 26007 5410 26016
rect 5262 25936 5318 25945
rect 5262 25871 5318 25880
rect 5276 24954 5304 25871
rect 5368 25362 5396 26007
rect 5356 25356 5408 25362
rect 5356 25298 5408 25304
rect 5356 25220 5408 25226
rect 5356 25162 5408 25168
rect 5368 25129 5396 25162
rect 5354 25120 5410 25129
rect 5354 25055 5410 25064
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 5356 24676 5408 24682
rect 5460 24664 5488 27406
rect 5552 26926 5580 28455
rect 5644 27946 5672 28966
rect 5632 27940 5684 27946
rect 5632 27882 5684 27888
rect 5644 27713 5672 27882
rect 5630 27704 5686 27713
rect 5736 27674 5764 29446
rect 5828 29102 5856 30246
rect 5920 30190 5948 30495
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5920 29345 5948 30126
rect 5906 29336 5962 29345
rect 5906 29271 5962 29280
rect 5816 29096 5868 29102
rect 5816 29038 5868 29044
rect 5816 28960 5868 28966
rect 5814 28928 5816 28937
rect 5868 28928 5870 28937
rect 5814 28863 5870 28872
rect 5816 28688 5868 28694
rect 5816 28630 5868 28636
rect 5630 27639 5686 27648
rect 5724 27668 5776 27674
rect 5540 26920 5592 26926
rect 5540 26862 5592 26868
rect 5644 26790 5672 27639
rect 5724 27610 5776 27616
rect 5724 27532 5776 27538
rect 5724 27474 5776 27480
rect 5632 26784 5684 26790
rect 5632 26726 5684 26732
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5552 26382 5580 26522
rect 5632 26512 5684 26518
rect 5632 26454 5684 26460
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5540 26240 5592 26246
rect 5540 26182 5592 26188
rect 5552 25498 5580 26182
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5538 25256 5594 25265
rect 5538 25191 5594 25200
rect 5552 24886 5580 25191
rect 5540 24880 5592 24886
rect 5540 24822 5592 24828
rect 5408 24636 5488 24664
rect 5356 24618 5408 24624
rect 5262 24576 5318 24585
rect 5262 24511 5318 24520
rect 5446 24576 5502 24585
rect 5446 24511 5502 24520
rect 5276 24426 5304 24511
rect 5460 24426 5488 24511
rect 5276 24398 5488 24426
rect 5264 24336 5316 24342
rect 5264 24278 5316 24284
rect 5356 24336 5408 24342
rect 5552 24324 5580 24822
rect 5644 24750 5672 26454
rect 5736 26081 5764 27474
rect 5828 27334 5856 28630
rect 5920 27878 5948 29271
rect 6012 27946 6040 31436
rect 6104 31278 6132 31758
rect 6196 31754 6224 32234
rect 6184 31748 6236 31754
rect 6184 31690 6236 31696
rect 6196 31385 6224 31690
rect 6182 31376 6238 31385
rect 6182 31311 6238 31320
rect 6288 31278 6316 32302
rect 6380 31822 6408 32728
rect 6460 32496 6512 32502
rect 6460 32438 6512 32444
rect 6368 31816 6420 31822
rect 6368 31758 6420 31764
rect 6380 31414 6408 31758
rect 6368 31408 6420 31414
rect 6368 31350 6420 31356
rect 6472 31346 6500 32438
rect 6552 32360 6604 32366
rect 6552 32302 6604 32308
rect 6564 31482 6592 32302
rect 6552 31476 6604 31482
rect 6552 31418 6604 31424
rect 6460 31340 6512 31346
rect 6460 31282 6512 31288
rect 6656 31278 6684 32864
rect 6736 32846 6788 32852
rect 6736 32768 6788 32774
rect 6736 32710 6788 32716
rect 6748 31958 6776 32710
rect 6840 32026 6868 32914
rect 6920 32768 6972 32774
rect 6920 32710 6972 32716
rect 6932 32570 6960 32710
rect 6920 32564 6972 32570
rect 6920 32506 6972 32512
rect 6932 32201 6960 32506
rect 7024 32298 7052 32914
rect 7116 32774 7144 33254
rect 7104 32768 7156 32774
rect 7104 32710 7156 32716
rect 7116 32570 7144 32710
rect 7104 32564 7156 32570
rect 7104 32506 7156 32512
rect 7208 32450 7236 33895
rect 7300 32774 7328 34478
rect 7380 34060 7432 34066
rect 7380 34002 7432 34008
rect 7392 33697 7420 34002
rect 7378 33688 7434 33697
rect 7378 33623 7434 33632
rect 7380 33380 7432 33386
rect 7380 33322 7432 33328
rect 7392 33289 7420 33322
rect 7378 33280 7434 33289
rect 7378 33215 7434 33224
rect 7484 33153 7512 35090
rect 7470 33144 7526 33153
rect 7576 33130 7604 36518
rect 7668 33862 7696 36638
rect 7748 36576 7800 36582
rect 7748 36518 7800 36524
rect 7760 36242 7788 36518
rect 7748 36236 7800 36242
rect 7748 36178 7800 36184
rect 7852 35834 7880 37402
rect 8036 37346 8064 38354
rect 8128 38321 8156 39460
rect 8208 39442 8260 39448
rect 8496 39438 8524 39782
rect 8484 39432 8536 39438
rect 8312 39392 8484 39420
rect 8312 39250 8340 39392
rect 8484 39374 8536 39380
rect 8220 39222 8340 39250
rect 8220 39030 8248 39222
rect 8390 39128 8446 39137
rect 8300 39092 8352 39098
rect 8390 39063 8392 39072
rect 8300 39034 8352 39040
rect 8444 39063 8446 39072
rect 8392 39034 8444 39040
rect 8208 39024 8260 39030
rect 8312 39001 8340 39034
rect 8208 38966 8260 38972
rect 8298 38992 8354 39001
rect 8298 38927 8354 38936
rect 8392 38956 8444 38962
rect 8392 38898 8444 38904
rect 8208 38888 8260 38894
rect 8208 38830 8260 38836
rect 8300 38888 8352 38894
rect 8404 38842 8432 38898
rect 8352 38836 8432 38842
rect 8300 38830 8432 38836
rect 8114 38312 8170 38321
rect 8114 38247 8170 38256
rect 8116 38208 8168 38214
rect 8116 38150 8168 38156
rect 8128 37942 8156 38150
rect 8116 37936 8168 37942
rect 8116 37878 8168 37884
rect 8220 37466 8248 38830
rect 8312 38814 8432 38830
rect 8300 38752 8352 38758
rect 8484 38752 8536 38758
rect 8352 38712 8432 38740
rect 8300 38694 8352 38700
rect 8300 38480 8352 38486
rect 8404 38457 8432 38712
rect 8484 38694 8536 38700
rect 8300 38422 8352 38428
rect 8390 38448 8446 38457
rect 8312 38298 8340 38422
rect 8390 38383 8392 38392
rect 8444 38383 8446 38392
rect 8392 38354 8444 38360
rect 8496 38321 8524 38694
rect 8588 38593 8616 39782
rect 8680 39681 8708 39850
rect 8772 39817 8800 39850
rect 8944 39840 8996 39846
rect 8758 39808 8814 39817
rect 8758 39743 8814 39752
rect 8864 39800 8944 39828
rect 8666 39672 8722 39681
rect 8864 39658 8892 39800
rect 8944 39782 8996 39788
rect 8666 39607 8722 39616
rect 8772 39630 8892 39658
rect 8944 39636 8996 39642
rect 8668 39296 8720 39302
rect 8668 39238 8720 39244
rect 8680 38758 8708 39238
rect 8668 38752 8720 38758
rect 8668 38694 8720 38700
rect 8574 38584 8630 38593
rect 8574 38519 8630 38528
rect 8772 38321 8800 39630
rect 8944 39578 8996 39584
rect 8956 39506 8984 39578
rect 8944 39500 8996 39506
rect 8944 39442 8996 39448
rect 9036 39500 9088 39506
rect 9036 39442 9088 39448
rect 8852 39296 8904 39302
rect 8852 39238 8904 39244
rect 8864 38894 8892 39238
rect 8956 39030 8984 39442
rect 8944 39024 8996 39030
rect 8944 38966 8996 38972
rect 8852 38888 8904 38894
rect 8852 38830 8904 38836
rect 8944 38888 8996 38894
rect 8944 38830 8996 38836
rect 8956 38554 8984 38830
rect 8944 38548 8996 38554
rect 8944 38490 8996 38496
rect 8944 38412 8996 38418
rect 8944 38354 8996 38360
rect 8482 38312 8538 38321
rect 8312 38270 8432 38298
rect 8404 37913 8432 38270
rect 8482 38247 8538 38256
rect 8758 38312 8814 38321
rect 8758 38247 8814 38256
rect 8482 38176 8538 38185
rect 8956 38162 8984 38354
rect 8482 38111 8538 38120
rect 8936 38134 8984 38162
rect 8496 37992 8524 38111
rect 8936 37992 8964 38134
rect 8496 37964 8616 37992
rect 8390 37904 8446 37913
rect 8588 37874 8616 37964
rect 8772 37964 8964 37992
rect 8390 37839 8446 37848
rect 8576 37868 8628 37874
rect 8404 37806 8432 37839
rect 8576 37810 8628 37816
rect 8392 37800 8444 37806
rect 8772 37754 8800 37964
rect 9048 37924 9076 39442
rect 9140 38457 9168 40344
rect 9232 38554 9260 40718
rect 9404 40724 9456 40730
rect 9404 40666 9456 40672
rect 9416 40186 9444 40666
rect 9508 40633 9536 41024
rect 9600 41398 9720 41426
rect 9494 40624 9550 40633
rect 9494 40559 9550 40568
rect 9404 40180 9456 40186
rect 9404 40122 9456 40128
rect 9404 39432 9456 39438
rect 9508 39420 9536 40559
rect 9600 40390 9628 41398
rect 9784 41290 9812 41618
rect 9864 41472 9916 41478
rect 9864 41414 9916 41420
rect 9692 41274 9812 41290
rect 9680 41268 9812 41274
rect 9732 41262 9812 41268
rect 9680 41210 9732 41216
rect 9680 40520 9732 40526
rect 9680 40462 9732 40468
rect 9588 40384 9640 40390
rect 9588 40326 9640 40332
rect 9600 39642 9628 40326
rect 9588 39636 9640 39642
rect 9588 39578 9640 39584
rect 9456 39392 9536 39420
rect 9692 39386 9720 40462
rect 9876 39914 9904 41414
rect 9968 40168 9996 41958
rect 10062 41372 10370 41381
rect 10062 41370 10068 41372
rect 10124 41370 10148 41372
rect 10204 41370 10228 41372
rect 10284 41370 10308 41372
rect 10364 41370 10370 41372
rect 10124 41318 10126 41370
rect 10306 41318 10308 41370
rect 10062 41316 10068 41318
rect 10124 41316 10148 41318
rect 10204 41316 10228 41318
rect 10284 41316 10308 41318
rect 10364 41316 10370 41318
rect 10062 41307 10370 41316
rect 10140 40996 10192 41002
rect 10140 40938 10192 40944
rect 10152 40730 10180 40938
rect 10324 40928 10376 40934
rect 10324 40870 10376 40876
rect 10140 40724 10192 40730
rect 10140 40666 10192 40672
rect 10336 40594 10364 40870
rect 10140 40588 10192 40594
rect 10140 40530 10192 40536
rect 10324 40588 10376 40594
rect 10324 40530 10376 40536
rect 10152 40390 10180 40530
rect 10428 40458 10456 42792
rect 10508 42774 10560 42780
rect 10600 42764 10652 42770
rect 10600 42706 10652 42712
rect 10508 42288 10560 42294
rect 10508 42230 10560 42236
rect 10416 40452 10468 40458
rect 10416 40394 10468 40400
rect 10140 40384 10192 40390
rect 10140 40326 10192 40332
rect 10062 40284 10370 40293
rect 10062 40282 10068 40284
rect 10124 40282 10148 40284
rect 10204 40282 10228 40284
rect 10284 40282 10308 40284
rect 10364 40282 10370 40284
rect 10124 40230 10126 40282
rect 10306 40230 10308 40282
rect 10062 40228 10068 40230
rect 10124 40228 10148 40230
rect 10204 40228 10228 40230
rect 10284 40228 10308 40230
rect 10364 40228 10370 40230
rect 10062 40219 10370 40228
rect 9968 40140 10180 40168
rect 10048 40044 10100 40050
rect 10048 39986 10100 39992
rect 9864 39908 9916 39914
rect 9864 39850 9916 39856
rect 9956 39840 10008 39846
rect 9956 39782 10008 39788
rect 9772 39636 9824 39642
rect 9772 39578 9824 39584
rect 9404 39374 9456 39380
rect 9312 38752 9364 38758
rect 9312 38694 9364 38700
rect 9220 38548 9272 38554
rect 9220 38490 9272 38496
rect 9126 38448 9182 38457
rect 9324 38434 9352 38694
rect 9126 38383 9182 38392
rect 9232 38406 9352 38434
rect 9128 38276 9180 38282
rect 9128 38218 9180 38224
rect 9140 38010 9168 38218
rect 9232 38214 9260 38406
rect 9312 38344 9364 38350
rect 9312 38286 9364 38292
rect 9220 38208 9272 38214
rect 9220 38150 9272 38156
rect 9128 38004 9180 38010
rect 9324 37992 9352 38286
rect 9416 38185 9444 39374
rect 9600 39358 9720 39386
rect 9600 39098 9628 39358
rect 9680 39296 9732 39302
rect 9680 39238 9732 39244
rect 9588 39092 9640 39098
rect 9588 39034 9640 39040
rect 9588 38956 9640 38962
rect 9508 38916 9588 38944
rect 9402 38176 9458 38185
rect 9402 38111 9458 38120
rect 9180 37964 9260 37992
rect 9324 37964 9444 37992
rect 9128 37946 9180 37952
rect 8392 37742 8444 37748
rect 8208 37460 8260 37466
rect 8404 37448 8432 37742
rect 8588 37726 8800 37754
rect 8864 37896 9076 37924
rect 8208 37402 8260 37408
rect 8312 37420 8432 37448
rect 8482 37496 8538 37505
rect 8482 37431 8538 37440
rect 8036 37318 8248 37346
rect 8024 37256 8076 37262
rect 8024 37198 8076 37204
rect 7932 36848 7984 36854
rect 7930 36816 7932 36825
rect 7984 36816 7986 36825
rect 7930 36751 7986 36760
rect 7932 36712 7984 36718
rect 7932 36654 7984 36660
rect 7944 36378 7972 36654
rect 7932 36372 7984 36378
rect 7932 36314 7984 36320
rect 7840 35828 7892 35834
rect 7840 35770 7892 35776
rect 7852 35306 7880 35770
rect 7852 35278 7972 35306
rect 8036 35290 8064 37198
rect 8116 37188 8168 37194
rect 8116 37130 8168 37136
rect 8128 36242 8156 37130
rect 8220 36582 8248 37318
rect 8312 37126 8340 37420
rect 8392 37324 8444 37330
rect 8392 37266 8444 37272
rect 8300 37120 8352 37126
rect 8300 37062 8352 37068
rect 8312 36582 8340 37062
rect 8404 36718 8432 37266
rect 8392 36712 8444 36718
rect 8390 36680 8392 36689
rect 8444 36680 8446 36689
rect 8390 36615 8446 36624
rect 8208 36576 8260 36582
rect 8208 36518 8260 36524
rect 8300 36576 8352 36582
rect 8300 36518 8352 36524
rect 8116 36236 8168 36242
rect 8116 36178 8168 36184
rect 8220 35494 8248 36518
rect 8312 35698 8340 36518
rect 8404 36378 8432 36615
rect 8392 36372 8444 36378
rect 8392 36314 8444 36320
rect 8496 36242 8524 37431
rect 8588 37233 8616 37726
rect 8668 37664 8720 37670
rect 8668 37606 8720 37612
rect 8760 37664 8812 37670
rect 8760 37606 8812 37612
rect 8680 37505 8708 37606
rect 8666 37496 8722 37505
rect 8772 37466 8800 37606
rect 8666 37431 8722 37440
rect 8760 37460 8812 37466
rect 8574 37224 8630 37233
rect 8574 37159 8630 37168
rect 8680 36650 8708 37431
rect 8760 37402 8812 37408
rect 8864 37330 8892 37896
rect 9128 37800 9180 37806
rect 9048 37760 9128 37788
rect 8852 37324 8904 37330
rect 8852 37266 8904 37272
rect 8760 36712 8812 36718
rect 8760 36654 8812 36660
rect 8668 36644 8720 36650
rect 8668 36586 8720 36592
rect 8680 36242 8708 36586
rect 8484 36236 8536 36242
rect 8484 36178 8536 36184
rect 8668 36236 8720 36242
rect 8668 36178 8720 36184
rect 8390 36136 8446 36145
rect 8390 36071 8446 36080
rect 8404 36038 8432 36071
rect 8392 36032 8444 36038
rect 8496 36009 8524 36178
rect 8668 36032 8720 36038
rect 8392 35974 8444 35980
rect 8482 36000 8538 36009
rect 8300 35692 8352 35698
rect 8300 35634 8352 35640
rect 8208 35488 8260 35494
rect 8208 35430 8260 35436
rect 8404 35306 8432 35974
rect 8668 35974 8720 35980
rect 8482 35935 8538 35944
rect 8574 35728 8630 35737
rect 8574 35663 8630 35672
rect 8588 35630 8616 35663
rect 8576 35624 8628 35630
rect 8576 35566 8628 35572
rect 7748 35080 7800 35086
rect 7748 35022 7800 35028
rect 7656 33856 7708 33862
rect 7656 33798 7708 33804
rect 7656 33652 7708 33658
rect 7656 33594 7708 33600
rect 7668 33318 7696 33594
rect 7656 33312 7708 33318
rect 7656 33254 7708 33260
rect 7576 33102 7696 33130
rect 7470 33079 7526 33088
rect 7564 33040 7616 33046
rect 7564 32982 7616 32988
rect 7472 32972 7524 32978
rect 7472 32914 7524 32920
rect 7380 32836 7432 32842
rect 7380 32778 7432 32784
rect 7288 32768 7340 32774
rect 7288 32710 7340 32716
rect 7208 32422 7328 32450
rect 7392 32434 7420 32778
rect 7196 32360 7248 32366
rect 7196 32302 7248 32308
rect 7012 32292 7064 32298
rect 7012 32234 7064 32240
rect 6918 32192 6974 32201
rect 6918 32127 6974 32136
rect 6828 32020 6880 32026
rect 6828 31962 6880 31968
rect 6736 31952 6788 31958
rect 7024 31929 7052 32234
rect 7102 32056 7158 32065
rect 7102 31991 7158 32000
rect 6736 31894 6788 31900
rect 7010 31920 7066 31929
rect 6828 31884 6880 31890
rect 6880 31844 6960 31872
rect 7010 31855 7066 31864
rect 6828 31826 6880 31832
rect 6736 31816 6788 31822
rect 6734 31784 6736 31793
rect 6788 31784 6790 31793
rect 6790 31742 6868 31770
rect 6734 31719 6790 31728
rect 6736 31680 6788 31686
rect 6734 31648 6736 31657
rect 6788 31648 6790 31657
rect 6734 31583 6790 31592
rect 6840 31464 6868 31742
rect 6932 31686 6960 31844
rect 7116 31822 7144 31991
rect 7104 31816 7156 31822
rect 7010 31784 7066 31793
rect 7104 31758 7156 31764
rect 7208 31754 7236 32302
rect 7300 32042 7328 32422
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 7484 32366 7512 32914
rect 7472 32360 7524 32366
rect 7472 32302 7524 32308
rect 7300 32014 7512 32042
rect 7576 32026 7604 32982
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 7010 31719 7066 31728
rect 7196 31748 7248 31754
rect 6920 31680 6972 31686
rect 6920 31622 6972 31628
rect 6840 31436 6960 31464
rect 6736 31408 6788 31414
rect 6788 31368 6868 31396
rect 6736 31350 6788 31356
rect 6092 31272 6144 31278
rect 6092 31214 6144 31220
rect 6184 31272 6236 31278
rect 6184 31214 6236 31220
rect 6276 31272 6328 31278
rect 6276 31214 6328 31220
rect 6644 31272 6696 31278
rect 6644 31214 6696 31220
rect 6196 30598 6224 31214
rect 6288 30734 6316 31214
rect 6460 31204 6512 31210
rect 6460 31146 6512 31152
rect 6472 30938 6500 31146
rect 6656 30938 6684 31214
rect 6460 30932 6512 30938
rect 6380 30892 6460 30920
rect 6276 30728 6328 30734
rect 6276 30670 6328 30676
rect 6184 30592 6236 30598
rect 6184 30534 6236 30540
rect 6092 30388 6144 30394
rect 6196 30376 6224 30534
rect 6144 30348 6224 30376
rect 6092 30330 6144 30336
rect 6092 30184 6144 30190
rect 6092 30126 6144 30132
rect 6184 30184 6236 30190
rect 6184 30126 6236 30132
rect 6104 29850 6132 30126
rect 6092 29844 6144 29850
rect 6092 29786 6144 29792
rect 6092 29504 6144 29510
rect 6092 29446 6144 29452
rect 6000 27940 6052 27946
rect 6000 27882 6052 27888
rect 5908 27872 5960 27878
rect 6012 27849 6040 27882
rect 5908 27814 5960 27820
rect 5998 27840 6054 27849
rect 5920 27418 5948 27814
rect 5998 27775 6054 27784
rect 6012 27606 6040 27775
rect 6000 27600 6052 27606
rect 6000 27542 6052 27548
rect 5920 27390 6040 27418
rect 5816 27328 5868 27334
rect 5814 27296 5816 27305
rect 5868 27296 5870 27305
rect 5814 27231 5870 27240
rect 6012 26858 6040 27390
rect 6000 26852 6052 26858
rect 6000 26794 6052 26800
rect 5814 26752 5870 26761
rect 5814 26687 5870 26696
rect 5722 26072 5778 26081
rect 5722 26007 5778 26016
rect 5724 25968 5776 25974
rect 5722 25936 5724 25945
rect 5776 25936 5778 25945
rect 5722 25871 5778 25880
rect 5724 25832 5776 25838
rect 5724 25774 5776 25780
rect 5736 25702 5764 25774
rect 5724 25696 5776 25702
rect 5724 25638 5776 25644
rect 5736 24993 5764 25638
rect 5722 24984 5778 24993
rect 5722 24919 5778 24928
rect 5722 24848 5778 24857
rect 5722 24783 5724 24792
rect 5776 24783 5778 24792
rect 5724 24754 5776 24760
rect 5632 24744 5684 24750
rect 5630 24712 5632 24721
rect 5684 24712 5686 24721
rect 5630 24647 5686 24656
rect 5724 24676 5776 24682
rect 5724 24618 5776 24624
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5408 24296 5580 24324
rect 5356 24278 5408 24284
rect 5276 24188 5304 24278
rect 5356 24200 5408 24206
rect 5276 24160 5356 24188
rect 5356 24142 5408 24148
rect 5262 23896 5318 23905
rect 5460 23866 5488 24296
rect 5644 24256 5672 24550
rect 5736 24449 5764 24618
rect 5722 24440 5778 24449
rect 5722 24375 5778 24384
rect 5552 24228 5672 24256
rect 5828 24246 5856 26687
rect 6000 26580 6052 26586
rect 6000 26522 6052 26528
rect 5906 26480 5962 26489
rect 5906 26415 5962 26424
rect 5920 25906 5948 26415
rect 5908 25900 5960 25906
rect 5908 25842 5960 25848
rect 5906 25800 5962 25809
rect 5906 25735 5962 25744
rect 5920 25265 5948 25735
rect 5906 25256 5962 25265
rect 5906 25191 5962 25200
rect 5908 25152 5960 25158
rect 5908 25094 5960 25100
rect 5920 24857 5948 25094
rect 5906 24848 5962 24857
rect 5906 24783 5962 24792
rect 6012 24614 6040 26522
rect 6104 26450 6132 29446
rect 6196 29102 6224 30126
rect 6184 29096 6236 29102
rect 6184 29038 6236 29044
rect 6184 28960 6236 28966
rect 6184 28902 6236 28908
rect 6196 28257 6224 28902
rect 6288 28762 6316 30670
rect 6380 29714 6408 30892
rect 6460 30874 6512 30880
rect 6644 30932 6696 30938
rect 6644 30874 6696 30880
rect 6736 30932 6788 30938
rect 6736 30874 6788 30880
rect 6552 30592 6604 30598
rect 6550 30560 6552 30569
rect 6604 30560 6606 30569
rect 6550 30495 6606 30504
rect 6460 30388 6512 30394
rect 6460 30330 6512 30336
rect 6472 29714 6500 30330
rect 6552 30320 6604 30326
rect 6552 30262 6604 30268
rect 6564 30190 6592 30262
rect 6552 30184 6604 30190
rect 6552 30126 6604 30132
rect 6564 29714 6592 30126
rect 6748 29889 6776 30874
rect 6734 29880 6790 29889
rect 6734 29815 6790 29824
rect 6368 29708 6420 29714
rect 6368 29650 6420 29656
rect 6460 29708 6512 29714
rect 6460 29650 6512 29656
rect 6552 29708 6604 29714
rect 6552 29650 6604 29656
rect 6736 29708 6788 29714
rect 6736 29650 6788 29656
rect 6368 29504 6420 29510
rect 6368 29446 6420 29452
rect 6380 28937 6408 29446
rect 6472 29306 6500 29650
rect 6644 29572 6696 29578
rect 6644 29514 6696 29520
rect 6550 29336 6606 29345
rect 6460 29300 6512 29306
rect 6550 29271 6606 29280
rect 6460 29242 6512 29248
rect 6458 29200 6514 29209
rect 6458 29135 6514 29144
rect 6472 29034 6500 29135
rect 6460 29028 6512 29034
rect 6460 28970 6512 28976
rect 6366 28928 6422 28937
rect 6366 28863 6422 28872
rect 6276 28756 6328 28762
rect 6276 28698 6328 28704
rect 6182 28248 6238 28257
rect 6182 28183 6238 28192
rect 6184 28144 6236 28150
rect 6182 28112 6184 28121
rect 6236 28112 6238 28121
rect 6182 28047 6238 28056
rect 6184 28008 6236 28014
rect 6288 27996 6316 28698
rect 6380 28626 6408 28863
rect 6564 28626 6592 29271
rect 6656 28994 6684 29514
rect 6748 29102 6776 29650
rect 6840 29510 6868 31368
rect 6932 30326 6960 31436
rect 6920 30320 6972 30326
rect 6920 30262 6972 30268
rect 6920 30184 6972 30190
rect 6920 30126 6972 30132
rect 6828 29504 6880 29510
rect 6828 29446 6880 29452
rect 6932 29306 6960 30126
rect 6828 29300 6880 29306
rect 6828 29242 6880 29248
rect 6920 29300 6972 29306
rect 6920 29242 6972 29248
rect 6840 29186 6868 29242
rect 6840 29158 6960 29186
rect 6736 29096 6788 29102
rect 6736 29038 6788 29044
rect 6826 29064 6882 29073
rect 6826 28999 6882 29008
rect 6656 28966 6776 28994
rect 6368 28620 6420 28626
rect 6368 28562 6420 28568
rect 6460 28620 6512 28626
rect 6460 28562 6512 28568
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 6236 27968 6316 27996
rect 6184 27950 6236 27956
rect 6288 27538 6316 27968
rect 6276 27532 6328 27538
rect 6276 27474 6328 27480
rect 6184 27328 6236 27334
rect 6184 27270 6236 27276
rect 6274 27296 6330 27305
rect 6092 26444 6144 26450
rect 6196 26432 6224 27270
rect 6274 27231 6330 27240
rect 6288 26858 6316 27231
rect 6380 26994 6408 28562
rect 6472 27985 6500 28562
rect 6564 28014 6592 28562
rect 6748 28506 6776 28966
rect 6656 28478 6776 28506
rect 6552 28008 6604 28014
rect 6458 27976 6514 27985
rect 6552 27950 6604 27956
rect 6458 27911 6514 27920
rect 6656 27656 6684 28478
rect 6736 28008 6788 28014
rect 6736 27950 6788 27956
rect 6748 27713 6776 27950
rect 6564 27628 6684 27656
rect 6734 27704 6790 27713
rect 6734 27639 6790 27648
rect 6458 27024 6514 27033
rect 6368 26988 6420 26994
rect 6458 26959 6514 26968
rect 6368 26930 6420 26936
rect 6472 26926 6500 26959
rect 6460 26920 6512 26926
rect 6460 26862 6512 26868
rect 6276 26852 6328 26858
rect 6276 26794 6328 26800
rect 6368 26784 6420 26790
rect 6368 26726 6420 26732
rect 6380 26518 6408 26726
rect 6472 26625 6500 26862
rect 6458 26616 6514 26625
rect 6458 26551 6514 26560
rect 6368 26512 6420 26518
rect 6368 26454 6420 26460
rect 6276 26444 6328 26450
rect 6196 26404 6276 26432
rect 6092 26386 6144 26392
rect 6276 26386 6328 26392
rect 6276 26308 6328 26314
rect 6276 26250 6328 26256
rect 6460 26308 6512 26314
rect 6460 26250 6512 26256
rect 6184 25968 6236 25974
rect 6090 25936 6146 25945
rect 6184 25910 6236 25916
rect 6090 25871 6146 25880
rect 6104 25838 6132 25871
rect 6092 25832 6144 25838
rect 6092 25774 6144 25780
rect 6196 25430 6224 25910
rect 6184 25424 6236 25430
rect 6184 25366 6236 25372
rect 6288 25362 6316 26250
rect 6368 26240 6420 26246
rect 6368 26182 6420 26188
rect 6276 25356 6328 25362
rect 6276 25298 6328 25304
rect 6184 25220 6236 25226
rect 6184 25162 6236 25168
rect 6196 24868 6224 25162
rect 6276 24880 6328 24886
rect 6090 24848 6146 24857
rect 6196 24840 6276 24868
rect 6276 24822 6328 24828
rect 6090 24783 6146 24792
rect 6000 24608 6052 24614
rect 6000 24550 6052 24556
rect 5552 24120 5580 24228
rect 5828 24218 6040 24246
rect 5908 24132 5960 24138
rect 5552 24092 5672 24120
rect 5262 23831 5318 23840
rect 5448 23860 5500 23866
rect 5276 23662 5304 23831
rect 5448 23802 5500 23808
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 5368 23066 5396 23734
rect 5460 23662 5488 23802
rect 5448 23656 5500 23662
rect 5644 23633 5672 24092
rect 5908 24074 5960 24080
rect 5920 23644 5948 24074
rect 5448 23598 5500 23604
rect 5630 23624 5686 23633
rect 5460 23526 5488 23598
rect 5828 23616 5948 23644
rect 5630 23559 5686 23568
rect 5724 23588 5776 23594
rect 5724 23530 5776 23536
rect 5448 23520 5500 23526
rect 5448 23462 5500 23468
rect 5632 23520 5684 23526
rect 5736 23497 5764 23530
rect 5632 23462 5684 23468
rect 5722 23488 5778 23497
rect 5092 22596 5212 22624
rect 5276 23038 5396 23066
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 4816 21814 4936 21842
rect 4816 21486 4844 21814
rect 5000 21672 5028 22374
rect 4908 21644 5028 21672
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4802 21176 4858 21185
rect 4712 21140 4764 21146
rect 4802 21111 4858 21120
rect 4712 21082 4764 21088
rect 4724 21049 4752 21082
rect 4816 21078 4844 21111
rect 4804 21072 4856 21078
rect 4710 21040 4766 21049
rect 4804 21014 4856 21020
rect 4710 20975 4766 20984
rect 4252 20936 4304 20942
rect 4816 20913 4844 21014
rect 4908 21010 4936 21644
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 5000 21049 5028 21490
rect 4986 21040 5042 21049
rect 4896 21004 4948 21010
rect 4986 20975 5042 20984
rect 4896 20946 4948 20952
rect 4252 20878 4304 20884
rect 4802 20904 4858 20913
rect 4802 20839 4858 20848
rect 4712 20800 4764 20806
rect 4250 20768 4306 20777
rect 4712 20742 4764 20748
rect 4250 20703 4306 20712
rect 4264 20534 4292 20703
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 4080 19689 4108 19790
rect 4264 19786 4292 20334
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 4528 20052 4580 20058
rect 4580 20012 4660 20040
rect 4528 19994 4580 20000
rect 4526 19952 4582 19961
rect 4436 19916 4488 19922
rect 4526 19887 4582 19896
rect 4436 19858 4488 19864
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 4066 19680 4122 19689
rect 3662 19612 3970 19621
rect 4066 19615 4122 19624
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3700 19440 3752 19446
rect 3238 19343 3240 19352
rect 3292 19343 3294 19352
rect 3332 19372 3384 19378
rect 3240 19314 3292 19320
rect 3436 19366 3648 19394
rect 3700 19382 3752 19388
rect 3332 19314 3384 19320
rect 3146 18864 3202 18873
rect 3056 18828 3108 18834
rect 3146 18799 3202 18808
rect 3056 18770 3108 18776
rect 2884 18686 3004 18714
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2884 18222 2912 18566
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2976 18154 3004 18686
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2700 17836 2820 17864
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2700 17610 2728 17836
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2516 16114 2544 17478
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2686 16960 2742 16969
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2504 15972 2556 15978
rect 2504 15914 2556 15920
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2516 15706 2544 15914
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 1952 15632 2004 15638
rect 1952 15574 2004 15580
rect 1964 14890 1992 15574
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 2044 15360 2096 15366
rect 2044 15302 2096 15308
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 1964 14618 1992 14826
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2056 13938 2084 15302
rect 2148 15026 2176 15506
rect 2608 15502 2636 16934
rect 2686 16895 2742 16904
rect 2700 15570 2728 16895
rect 2792 16590 2820 17682
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 2884 17105 2912 17546
rect 2976 17134 3004 18090
rect 3068 17610 3096 18566
rect 3252 18306 3280 19314
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3160 18278 3280 18306
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 3160 17354 3188 18278
rect 3344 18222 3372 19110
rect 3436 18698 3464 19246
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3528 18834 3556 19110
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 3424 18692 3476 18698
rect 3424 18634 3476 18640
rect 3436 18358 3464 18634
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3422 18184 3478 18193
rect 3068 17326 3188 17354
rect 3068 17270 3096 17326
rect 3056 17264 3108 17270
rect 3148 17264 3200 17270
rect 3056 17206 3108 17212
rect 3146 17232 3148 17241
rect 3200 17232 3202 17241
rect 2964 17128 3016 17134
rect 2870 17096 2926 17105
rect 2964 17070 3016 17076
rect 2870 17031 2926 17040
rect 2884 16590 2912 17031
rect 2976 16658 3004 17070
rect 3068 16726 3096 17206
rect 3146 17167 3202 17176
rect 3056 16720 3108 16726
rect 3108 16680 3188 16708
rect 3056 16662 3108 16668
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2792 16250 2820 16390
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2778 15600 2834 15609
rect 2688 15564 2740 15570
rect 2976 15570 3004 16390
rect 3056 16176 3108 16182
rect 3056 16118 3108 16124
rect 2778 15535 2834 15544
rect 2964 15564 3016 15570
rect 2688 15506 2740 15512
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2226 15192 2282 15201
rect 2226 15127 2228 15136
rect 2280 15127 2282 15136
rect 2320 15156 2372 15162
rect 2228 15098 2280 15104
rect 2320 15098 2372 15104
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13530 1992 13806
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 1858 12472 1914 12481
rect 1858 12407 1914 12416
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1582 12064 1638 12073
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1400 11552 1452 11558
rect 1504 11529 1532 12038
rect 1582 11999 1638 12008
rect 1596 11694 1624 11999
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1584 11552 1636 11558
rect 1400 11494 1452 11500
rect 1490 11520 1546 11529
rect 1412 11257 1440 11494
rect 1584 11494 1636 11500
rect 1490 11455 1546 11464
rect 1398 11248 1454 11257
rect 1398 11183 1454 11192
rect 1596 10985 1624 11494
rect 1780 11354 1808 12242
rect 1964 12170 1992 13466
rect 2056 13394 2084 13874
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2056 12850 2084 13330
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 2044 12096 2096 12102
rect 1950 12064 2006 12073
rect 2044 12038 2096 12044
rect 1950 11999 2006 12008
rect 1964 11694 1992 11999
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 2056 11354 2084 12038
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1872 11082 1900 11154
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1124 10600 1176 10606
rect 1124 10542 1176 10548
rect 1308 10600 1360 10606
rect 1308 10542 1360 10548
rect 1320 10266 1348 10542
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1308 9512 1360 9518
rect 1308 9454 1360 9460
rect 1320 9178 1348 9454
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 7954 1440 8910
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1400 7472 1452 7478
rect 1400 7414 1452 7420
rect 1412 6730 1440 7414
rect 1504 6798 1532 9998
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9586 1716 9862
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 7546 1624 8434
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1596 7206 1624 7346
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1400 6724 1452 6730
rect 1400 6666 1452 6672
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5778 1440 6190
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5098 1440 5714
rect 1504 5710 1532 6598
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1504 5166 1532 5646
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1400 5092 1452 5098
rect 1400 5034 1452 5040
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1412 4282 1440 4762
rect 1596 4486 1624 7142
rect 1688 6866 1716 8366
rect 1780 8242 1808 10202
rect 1872 9654 1900 11018
rect 1964 10810 1992 11222
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1950 9072 2006 9081
rect 2006 9016 2084 9024
rect 1950 9007 1952 9016
rect 2004 8996 2084 9016
rect 1952 8978 2004 8984
rect 1780 8214 1900 8242
rect 1872 7290 1900 8214
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1780 7262 1900 7290
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1780 6202 1808 7262
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1872 6866 1900 7142
rect 1964 6934 1992 7890
rect 1952 6928 2004 6934
rect 1952 6870 2004 6876
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 2056 6254 2084 8996
rect 2148 8566 2176 14554
rect 2332 13870 2360 15098
rect 2424 15076 2452 15438
rect 2688 15088 2740 15094
rect 2424 15048 2688 15076
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2424 14414 2452 14894
rect 2608 14618 2636 15048
rect 2688 15030 2740 15036
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2700 14822 2728 14894
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2686 14648 2742 14657
rect 2596 14612 2648 14618
rect 2686 14583 2688 14592
rect 2596 14554 2648 14560
rect 2740 14583 2742 14592
rect 2688 14554 2740 14560
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2228 13796 2280 13802
rect 2228 13738 2280 13744
rect 2240 12782 2268 13738
rect 2320 13456 2372 13462
rect 2320 13398 2372 13404
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2228 12368 2280 12374
rect 2226 12336 2228 12345
rect 2280 12336 2282 12345
rect 2226 12271 2282 12280
rect 2332 12102 2360 13398
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11762 2360 12038
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 10810 2268 11086
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2332 10606 2360 11154
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2332 10266 2360 10542
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2332 9450 2360 9998
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2148 7546 2176 8026
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2228 7268 2280 7274
rect 2228 7210 2280 7216
rect 2240 7002 2268 7210
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 1688 6174 1808 6202
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 1952 6180 2004 6186
rect 1688 5234 1716 6174
rect 1952 6122 2004 6128
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1688 4010 1716 5170
rect 1768 5092 1820 5098
rect 1768 5034 1820 5040
rect 1780 4146 1808 5034
rect 1872 4554 1900 5714
rect 1964 5710 1992 6122
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 2148 5642 2176 6190
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 2148 5370 2176 5578
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2240 5250 2268 6802
rect 2148 5222 2268 5250
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 1964 4282 1992 4626
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1032 3052 1084 3058
rect 1032 2994 1084 3000
rect 1504 2910 1716 2938
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1412 1902 1440 2450
rect 1504 2446 1532 2910
rect 1688 2854 1716 2910
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1596 2650 1624 2790
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1504 1970 1532 2382
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 1596 2106 1624 2314
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1492 1964 1544 1970
rect 1492 1906 1544 1912
rect 1400 1896 1452 1902
rect 1400 1838 1452 1844
rect 1964 1358 1992 4014
rect 2056 3942 2084 5034
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2148 2854 2176 5222
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2240 4758 2268 4966
rect 2228 4752 2280 4758
rect 2228 4694 2280 4700
rect 2332 4690 2360 8978
rect 2424 7478 2452 12582
rect 2516 12374 2544 14418
rect 2608 14278 2636 14418
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2608 12986 2636 13874
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2608 12889 2636 12922
rect 2594 12880 2650 12889
rect 2594 12815 2650 12824
rect 2700 12714 2728 13466
rect 2792 13274 2820 15535
rect 2964 15506 3016 15512
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2884 14958 2912 15438
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2884 13433 2912 14758
rect 2870 13424 2926 13433
rect 2870 13359 2872 13368
rect 2924 13359 2926 13368
rect 2872 13330 2924 13336
rect 2976 13297 3004 15302
rect 2962 13288 3018 13297
rect 2792 13246 2912 13274
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2792 12850 2820 13126
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2688 12708 2740 12714
rect 2608 12668 2688 12696
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2608 11898 2636 12668
rect 2688 12650 2740 12656
rect 2686 12472 2742 12481
rect 2686 12407 2688 12416
rect 2740 12407 2742 12416
rect 2688 12378 2740 12384
rect 2686 12336 2742 12345
rect 2792 12306 2820 12786
rect 2884 12714 2912 13246
rect 2962 13223 3018 13232
rect 3068 13240 3096 16118
rect 3160 16046 3188 16680
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3160 14482 3188 15030
rect 3252 14618 3280 18158
rect 3422 18119 3478 18128
rect 3436 18068 3464 18119
rect 3344 18040 3464 18068
rect 3344 15366 3372 18040
rect 3528 17746 3556 18770
rect 3620 18630 3648 19366
rect 3712 19310 3740 19382
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3896 18737 3924 18770
rect 3882 18728 3938 18737
rect 3882 18663 3938 18672
rect 3988 18630 4016 19246
rect 4080 18970 4108 19450
rect 4264 19334 4292 19722
rect 4448 19514 4476 19858
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4540 19446 4568 19887
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 4172 19306 4292 19334
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4172 18850 4200 19306
rect 4342 19272 4398 19281
rect 4080 18822 4200 18850
rect 4264 19230 4342 19258
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 3976 18352 4028 18358
rect 3896 18312 3976 18340
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3436 17377 3464 17478
rect 3422 17368 3478 17377
rect 3422 17303 3478 17312
rect 3528 17218 3556 17546
rect 3712 17542 3740 18022
rect 3804 17649 3832 18090
rect 3896 17746 3924 18312
rect 3976 18294 4028 18300
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3988 17785 4016 18158
rect 4080 17882 4108 18822
rect 4264 18766 4292 19230
rect 4342 19207 4398 19216
rect 4526 19272 4582 19281
rect 4526 19207 4528 19216
rect 4580 19207 4582 19216
rect 4528 19178 4580 19184
rect 4632 19156 4660 20012
rect 4724 19378 4752 20742
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4816 20058 4844 20334
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4908 19786 4936 20946
rect 4988 20392 5040 20398
rect 5092 20369 5120 22596
rect 5276 22556 5304 23038
rect 5354 22944 5410 22953
rect 5354 22879 5410 22888
rect 5184 22528 5304 22556
rect 5184 22234 5212 22528
rect 5264 22432 5316 22438
rect 5264 22374 5316 22380
rect 5276 22273 5304 22374
rect 5262 22264 5318 22273
rect 5172 22228 5224 22234
rect 5262 22199 5318 22208
rect 5172 22170 5224 22176
rect 5276 22098 5304 22199
rect 5264 22092 5316 22098
rect 5264 22034 5316 22040
rect 5276 22001 5304 22034
rect 5262 21992 5318 22001
rect 5262 21927 5318 21936
rect 5170 21720 5226 21729
rect 5170 21655 5172 21664
rect 5224 21655 5226 21664
rect 5172 21626 5224 21632
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 5184 20777 5212 21490
rect 5368 21400 5396 22879
rect 5448 22704 5500 22710
rect 5446 22672 5448 22681
rect 5500 22672 5502 22681
rect 5446 22607 5502 22616
rect 5448 22500 5500 22506
rect 5448 22442 5500 22448
rect 5460 22166 5488 22442
rect 5448 22160 5500 22166
rect 5448 22102 5500 22108
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5460 21729 5488 21966
rect 5446 21720 5502 21729
rect 5446 21655 5502 21664
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5276 21372 5396 21400
rect 5170 20768 5226 20777
rect 5170 20703 5226 20712
rect 5172 20392 5224 20398
rect 4988 20334 5040 20340
rect 5078 20360 5134 20369
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4632 19128 4752 19156
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 4724 19009 4752 19128
rect 4710 19000 4766 19009
rect 4344 18964 4396 18970
rect 4710 18935 4766 18944
rect 4344 18906 4396 18912
rect 4356 18834 4384 18906
rect 4344 18828 4396 18834
rect 4724 18816 4752 18935
rect 4396 18788 4476 18816
rect 4344 18770 4396 18776
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4160 18624 4212 18630
rect 4158 18592 4160 18601
rect 4212 18592 4214 18601
rect 4158 18527 4214 18536
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 3974 17776 4030 17785
rect 3884 17740 3936 17746
rect 3974 17711 4030 17720
rect 3884 17682 3936 17688
rect 4068 17672 4120 17678
rect 3790 17640 3846 17649
rect 4068 17614 4120 17620
rect 3790 17575 3846 17584
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 4080 17338 4108 17614
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 3436 17202 3556 17218
rect 3424 17196 3556 17202
rect 3476 17190 3556 17196
rect 3424 17138 3476 17144
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3436 16114 3464 16594
rect 3528 16590 3556 17190
rect 3698 17232 3754 17241
rect 3698 17167 3754 17176
rect 3976 17196 4028 17202
rect 3712 17066 3740 17167
rect 3976 17138 4028 17144
rect 3884 17128 3936 17134
rect 3804 17088 3884 17116
rect 3700 17060 3752 17066
rect 3700 17002 3752 17008
rect 3804 16969 3832 17088
rect 3988 17105 4016 17138
rect 4068 17128 4120 17134
rect 3884 17070 3936 17076
rect 3974 17096 4030 17105
rect 4068 17070 4120 17076
rect 3974 17031 4030 17040
rect 3884 16992 3936 16998
rect 3790 16960 3846 16969
rect 3884 16934 3936 16940
rect 3790 16895 3846 16904
rect 3896 16590 3924 16934
rect 3516 16584 3568 16590
rect 3884 16584 3936 16590
rect 3516 16526 3568 16532
rect 3882 16552 3884 16561
rect 3936 16552 3938 16561
rect 3882 16487 3938 16496
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3528 16046 3556 16390
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 3698 16144 3754 16153
rect 3698 16079 3754 16088
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3712 15570 3740 16079
rect 4080 15706 4108 17070
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4172 15638 4200 18226
rect 4264 17746 4292 18702
rect 4342 18456 4398 18465
rect 4342 18391 4398 18400
rect 4356 18290 4384 18391
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4448 18086 4476 18788
rect 4540 18788 4844 18816
rect 4540 18290 4568 18788
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4528 18284 4580 18290
rect 4528 18226 4580 18232
rect 4632 18154 4660 18634
rect 4724 18465 4752 18634
rect 4710 18456 4766 18465
rect 4710 18391 4766 18400
rect 4620 18148 4672 18154
rect 4620 18090 4672 18096
rect 4436 18080 4488 18086
rect 4816 18057 4844 18788
rect 4436 18022 4488 18028
rect 4802 18048 4858 18057
rect 4322 17980 4630 17989
rect 4802 17983 4858 17992
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 4802 17912 4858 17921
rect 4344 17876 4396 17882
rect 4802 17847 4858 17856
rect 4344 17818 4396 17824
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4264 17241 4292 17682
rect 4250 17232 4306 17241
rect 4250 17167 4306 17176
rect 4356 17134 4384 17818
rect 4528 17808 4580 17814
rect 4528 17750 4580 17756
rect 4710 17776 4766 17785
rect 4436 17604 4488 17610
rect 4436 17546 4488 17552
rect 4448 17513 4476 17546
rect 4434 17504 4490 17513
rect 4434 17439 4490 17448
rect 4540 17320 4568 17750
rect 4620 17740 4672 17746
rect 4816 17746 4844 17847
rect 4710 17711 4766 17720
rect 4804 17740 4856 17746
rect 4620 17682 4672 17688
rect 4448 17292 4568 17320
rect 4344 17128 4396 17134
rect 4264 17088 4344 17116
rect 4264 16538 4292 17088
rect 4448 17105 4476 17292
rect 4526 17232 4582 17241
rect 4526 17167 4582 17176
rect 4344 17070 4396 17076
rect 4434 17096 4490 17105
rect 4540 17066 4568 17167
rect 4632 17134 4660 17682
rect 4724 17678 4752 17711
rect 4804 17682 4856 17688
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4434 17031 4490 17040
rect 4528 17060 4580 17066
rect 4528 17002 4580 17008
rect 4724 16969 4752 17614
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4816 17377 4844 17478
rect 4802 17368 4858 17377
rect 4802 17303 4858 17312
rect 4816 17134 4844 17303
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4710 16960 4766 16969
rect 4322 16892 4630 16901
rect 4710 16895 4766 16904
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 4264 16510 4384 16538
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4264 16114 4292 16390
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4356 15892 4384 16510
rect 4448 16114 4476 16662
rect 4710 16552 4766 16561
rect 4710 16487 4766 16496
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4724 16046 4752 16487
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4264 15864 4384 15892
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3712 15450 3740 15506
rect 3528 15422 3740 15450
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3332 14884 3384 14890
rect 3332 14826 3384 14832
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3252 14006 3280 14418
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 3146 13832 3202 13841
rect 3344 13802 3372 14826
rect 3436 14074 3464 14826
rect 3528 14618 3556 15422
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3436 13870 3464 14010
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3146 13767 3148 13776
rect 3200 13767 3202 13776
rect 3332 13796 3384 13802
rect 3148 13738 3200 13744
rect 3332 13738 3384 13744
rect 3238 13696 3294 13705
rect 3238 13631 3294 13640
rect 3252 13394 3280 13631
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3332 13320 3384 13326
rect 3238 13288 3294 13297
rect 3068 13212 3188 13240
rect 3384 13280 3464 13308
rect 3332 13262 3384 13268
rect 3238 13223 3294 13232
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 3054 13152 3110 13161
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2686 12271 2688 12280
rect 2740 12271 2742 12280
rect 2780 12300 2832 12306
rect 2688 12242 2740 12248
rect 2780 12242 2832 12248
rect 2976 12238 3004 13126
rect 3054 13087 3110 13096
rect 3068 12442 3096 13087
rect 3160 12986 3188 13212
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3160 12288 3188 12718
rect 3068 12260 3188 12288
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2516 8090 2544 11630
rect 2700 10248 2728 12106
rect 2962 12064 3018 12073
rect 2962 11999 3018 12008
rect 2778 11792 2834 11801
rect 2778 11727 2834 11736
rect 2792 11694 2820 11727
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2700 10220 2820 10248
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2608 9518 2636 9862
rect 2700 9518 2728 10066
rect 2792 10062 2820 10220
rect 2870 10160 2926 10169
rect 2870 10095 2872 10104
rect 2924 10095 2926 10104
rect 2872 10066 2924 10072
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2608 8906 2636 9454
rect 2700 9110 2728 9454
rect 2884 9178 2912 9454
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2424 6458 2452 7278
rect 2516 6866 2544 7822
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2688 6860 2740 6866
rect 2792 6848 2820 7346
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2884 6866 2912 7278
rect 2740 6820 2820 6848
rect 2872 6860 2924 6866
rect 2688 6802 2740 6808
rect 2872 6802 2924 6808
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5914 2452 6054
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2424 5778 2452 5850
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2332 4214 2360 4626
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2424 3534 2452 4082
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 3126 2268 3334
rect 2228 3120 2280 3126
rect 2228 3062 2280 3068
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 2136 2508 2188 2514
rect 2240 2496 2268 3062
rect 2332 2582 2360 3470
rect 2516 3398 2544 4150
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2608 3670 2636 3878
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 2990 2544 3334
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 2188 2468 2268 2496
rect 2136 2450 2188 2456
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2056 1426 2084 2382
rect 2332 1562 2360 2518
rect 2516 2514 2544 2926
rect 2608 2514 2636 3606
rect 2884 2990 2912 6802
rect 2976 6118 3004 11999
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 3068 5914 3096 12260
rect 3252 12186 3280 13223
rect 3332 13184 3384 13190
rect 3330 13152 3332 13161
rect 3384 13152 3386 13161
rect 3330 13087 3386 13096
rect 3436 12646 3464 13280
rect 3528 12986 3556 14418
rect 3712 14385 3740 14962
rect 3976 14952 4028 14958
rect 3974 14920 3976 14929
rect 4028 14920 4030 14929
rect 3884 14884 3936 14890
rect 3974 14855 4030 14864
rect 3884 14826 3936 14832
rect 3896 14793 3924 14826
rect 3882 14784 3938 14793
rect 3882 14719 3938 14728
rect 3896 14414 3924 14719
rect 3988 14550 4016 14855
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3884 14408 3936 14414
rect 3698 14376 3754 14385
rect 3884 14350 3936 14356
rect 3698 14311 3754 14320
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3790 13968 3846 13977
rect 3712 13462 3740 13942
rect 3790 13903 3846 13912
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3804 13394 3832 13903
rect 3884 13864 3936 13870
rect 4080 13818 4108 15438
rect 4264 15314 4292 15864
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 4816 15570 4844 16390
rect 4908 16046 4936 19722
rect 5000 19553 5028 20334
rect 5172 20334 5224 20340
rect 5078 20295 5134 20304
rect 4986 19544 5042 19553
rect 4986 19479 5042 19488
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 5000 18193 5028 19246
rect 5092 19174 5120 20295
rect 5184 20058 5212 20334
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 5276 18970 5304 21372
rect 5354 21312 5410 21321
rect 5354 21247 5410 21256
rect 5368 20942 5396 21247
rect 5460 21010 5488 21490
rect 5552 21185 5580 23054
rect 5644 22080 5672 23462
rect 5722 23423 5778 23432
rect 5828 23372 5856 23616
rect 5908 23520 5960 23526
rect 5908 23462 5960 23468
rect 5736 23344 5856 23372
rect 5736 22642 5764 23344
rect 5920 23186 5948 23462
rect 5816 23180 5868 23186
rect 5816 23122 5868 23128
rect 5908 23180 5960 23186
rect 5908 23122 5960 23128
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5828 22234 5856 23122
rect 5906 22944 5962 22953
rect 5906 22879 5962 22888
rect 5920 22778 5948 22879
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 5908 22636 5960 22642
rect 5908 22578 5960 22584
rect 5816 22228 5868 22234
rect 5816 22170 5868 22176
rect 5724 22092 5776 22098
rect 5644 22052 5724 22080
rect 5724 22034 5776 22040
rect 5920 22030 5948 22578
rect 5908 22024 5960 22030
rect 6012 22001 6040 24218
rect 6104 24206 6132 24783
rect 6276 24676 6328 24682
rect 6276 24618 6328 24624
rect 6184 24268 6236 24274
rect 6288 24256 6316 24618
rect 6380 24342 6408 26182
rect 6472 25129 6500 26250
rect 6564 25838 6592 27628
rect 6748 27606 6776 27639
rect 6736 27600 6788 27606
rect 6736 27542 6788 27548
rect 6736 26920 6788 26926
rect 6736 26862 6788 26868
rect 6748 26790 6776 26862
rect 6644 26784 6696 26790
rect 6644 26726 6696 26732
rect 6736 26784 6788 26790
rect 6736 26726 6788 26732
rect 6656 26450 6684 26726
rect 6734 26616 6790 26625
rect 6734 26551 6790 26560
rect 6644 26444 6696 26450
rect 6644 26386 6696 26392
rect 6748 26382 6776 26551
rect 6736 26376 6788 26382
rect 6736 26318 6788 26324
rect 6642 26208 6698 26217
rect 6642 26143 6698 26152
rect 6656 26042 6684 26143
rect 6644 26036 6696 26042
rect 6644 25978 6696 25984
rect 6736 26036 6788 26042
rect 6736 25978 6788 25984
rect 6748 25906 6776 25978
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6552 25832 6604 25838
rect 6552 25774 6604 25780
rect 6644 25832 6696 25838
rect 6644 25774 6696 25780
rect 6552 25696 6604 25702
rect 6656 25673 6684 25774
rect 6736 25696 6788 25702
rect 6552 25638 6604 25644
rect 6642 25664 6698 25673
rect 6564 25294 6592 25638
rect 6736 25638 6788 25644
rect 6642 25599 6698 25608
rect 6748 25537 6776 25638
rect 6734 25528 6790 25537
rect 6734 25463 6790 25472
rect 6736 25424 6788 25430
rect 6736 25366 6788 25372
rect 6644 25356 6696 25362
rect 6644 25298 6696 25304
rect 6552 25288 6604 25294
rect 6552 25230 6604 25236
rect 6458 25120 6514 25129
rect 6458 25055 6514 25064
rect 6472 24954 6500 25055
rect 6460 24948 6512 24954
rect 6460 24890 6512 24896
rect 6552 24608 6604 24614
rect 6458 24576 6514 24585
rect 6656 24596 6684 25298
rect 6604 24568 6684 24596
rect 6552 24550 6604 24556
rect 6458 24511 6514 24520
rect 6368 24336 6420 24342
rect 6368 24278 6420 24284
rect 6236 24228 6316 24256
rect 6184 24210 6236 24216
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6196 23905 6224 24210
rect 6380 24206 6408 24278
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6182 23896 6238 23905
rect 6182 23831 6238 23840
rect 6276 23588 6328 23594
rect 6196 23548 6276 23576
rect 6090 23352 6146 23361
rect 6090 23287 6146 23296
rect 6104 23186 6132 23287
rect 6196 23186 6224 23548
rect 6276 23530 6328 23536
rect 6274 23352 6330 23361
rect 6274 23287 6276 23296
rect 6328 23287 6330 23296
rect 6276 23258 6328 23264
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6184 23180 6236 23186
rect 6184 23122 6236 23128
rect 5908 21966 5960 21972
rect 5998 21992 6054 22001
rect 5998 21927 6054 21936
rect 5908 21616 5960 21622
rect 5908 21558 5960 21564
rect 5998 21584 6054 21593
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 5538 21176 5594 21185
rect 5538 21111 5594 21120
rect 5540 21072 5592 21078
rect 5540 21014 5592 21020
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5460 20874 5488 20946
rect 5448 20868 5500 20874
rect 5448 20810 5500 20816
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5460 19174 5488 19790
rect 5552 19378 5580 21014
rect 5644 20097 5672 21422
rect 5736 21010 5764 21422
rect 5816 21412 5868 21418
rect 5816 21354 5868 21360
rect 5724 21004 5776 21010
rect 5724 20946 5776 20952
rect 5724 20528 5776 20534
rect 5724 20470 5776 20476
rect 5736 20262 5764 20470
rect 5828 20398 5856 21354
rect 5920 21321 5948 21558
rect 5998 21519 6054 21528
rect 6012 21486 6040 21519
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 5906 21312 5962 21321
rect 5906 21247 5962 21256
rect 6104 21049 6132 23122
rect 6196 22778 6224 23122
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 6184 22772 6236 22778
rect 6184 22714 6236 22720
rect 6182 22672 6238 22681
rect 6182 22607 6238 22616
rect 6196 22574 6224 22607
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6196 22234 6224 22510
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6288 22166 6316 22986
rect 6276 22160 6328 22166
rect 6276 22102 6328 22108
rect 6274 21992 6330 22001
rect 6274 21927 6276 21936
rect 6328 21927 6330 21936
rect 6276 21898 6328 21904
rect 6184 21480 6236 21486
rect 6184 21422 6236 21428
rect 6276 21480 6328 21486
rect 6276 21422 6328 21428
rect 6090 21040 6146 21049
rect 6000 21004 6052 21010
rect 6090 20975 6146 20984
rect 6000 20946 6052 20952
rect 6012 20913 6040 20946
rect 5998 20904 6054 20913
rect 5998 20839 6054 20848
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 5816 20392 5868 20398
rect 5868 20352 5948 20380
rect 5816 20334 5868 20340
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5630 20088 5686 20097
rect 5630 20023 5632 20032
rect 5684 20023 5686 20032
rect 5632 19994 5684 20000
rect 5722 19816 5778 19825
rect 5722 19751 5778 19760
rect 5630 19680 5686 19689
rect 5630 19615 5686 19624
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5552 19281 5580 19314
rect 5644 19310 5672 19615
rect 5632 19304 5684 19310
rect 5538 19272 5594 19281
rect 5632 19246 5684 19252
rect 5538 19207 5594 19216
rect 5448 19168 5500 19174
rect 5644 19145 5672 19246
rect 5448 19110 5500 19116
rect 5630 19136 5686 19145
rect 5630 19071 5686 19080
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5078 18864 5134 18873
rect 5078 18799 5080 18808
rect 5132 18799 5134 18808
rect 5080 18770 5132 18776
rect 5080 18692 5132 18698
rect 5080 18634 5132 18640
rect 5092 18601 5120 18634
rect 5078 18592 5134 18601
rect 5078 18527 5134 18536
rect 5170 18456 5226 18465
rect 5170 18391 5172 18400
rect 5224 18391 5226 18400
rect 5172 18362 5224 18368
rect 5078 18320 5134 18329
rect 5078 18255 5134 18264
rect 5092 18222 5120 18255
rect 5080 18216 5132 18222
rect 4986 18184 5042 18193
rect 5172 18216 5224 18222
rect 5080 18158 5132 18164
rect 5170 18184 5172 18193
rect 5224 18184 5226 18193
rect 4986 18119 5042 18128
rect 5170 18119 5226 18128
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5170 18048 5226 18057
rect 5092 17882 5120 18022
rect 5170 17983 5226 17992
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5092 17270 5120 17682
rect 5080 17264 5132 17270
rect 5080 17206 5132 17212
rect 5184 17082 5212 17983
rect 5276 17785 5304 18906
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5262 17776 5318 17785
rect 5262 17711 5264 17720
rect 5316 17711 5318 17720
rect 5264 17682 5316 17688
rect 5262 17504 5318 17513
rect 5262 17439 5318 17448
rect 5092 17066 5212 17082
rect 5080 17060 5212 17066
rect 5132 17054 5212 17060
rect 5080 17002 5132 17008
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5000 16522 5028 16730
rect 4988 16516 5040 16522
rect 4988 16458 5040 16464
rect 5092 16402 5120 17002
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16590 5212 16934
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5092 16374 5212 16402
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4344 15428 4396 15434
rect 4344 15370 4396 15376
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4172 15286 4292 15314
rect 4172 15162 4200 15286
rect 4250 15192 4306 15201
rect 4160 15156 4212 15162
rect 4250 15127 4306 15136
rect 4160 15098 4212 15104
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14482 4200 14758
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4158 14376 4214 14385
rect 4158 14311 4160 14320
rect 4212 14311 4214 14320
rect 4160 14282 4212 14288
rect 3884 13806 3936 13812
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3896 13258 3924 13806
rect 3988 13790 4108 13818
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 3988 13410 4016 13790
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13530 4108 13670
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4172 13462 4200 13806
rect 4160 13456 4212 13462
rect 3988 13382 4108 13410
rect 4160 13398 4212 13404
rect 3884 13252 3936 13258
rect 3884 13194 3936 13200
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3160 12158 3280 12186
rect 3332 12232 3384 12238
rect 3712 12209 3740 12650
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3804 12306 3832 12582
rect 4080 12442 4108 13382
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4172 12850 4200 13262
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3332 12174 3384 12180
rect 3698 12200 3754 12209
rect 3160 7954 3188 12158
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3252 11898 3280 12038
rect 3344 11898 3372 12174
rect 3698 12135 3754 12144
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 3252 9042 3280 10678
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3252 8294 3280 8978
rect 3344 8974 3372 10406
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3160 7546 3188 7890
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3160 6361 3188 6734
rect 3146 6352 3202 6361
rect 3146 6287 3202 6296
rect 3252 6254 3280 6802
rect 3436 6746 3464 11154
rect 3528 9654 3556 11630
rect 3608 11552 3660 11558
rect 4080 11506 4108 12242
rect 3608 11494 3660 11500
rect 3620 11082 3648 11494
rect 3988 11478 4108 11506
rect 3988 11218 4016 11478
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3804 10130 3832 10542
rect 3882 10160 3938 10169
rect 3792 10124 3844 10130
rect 3882 10095 3884 10104
rect 3792 10066 3844 10072
rect 3936 10095 3938 10104
rect 3884 10066 3936 10072
rect 3988 9994 4016 10610
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3896 9042 3924 9386
rect 3988 9178 4016 9454
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3528 8430 3556 8978
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3528 7342 3556 8230
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 4080 7546 4108 11290
rect 4172 10742 4200 12650
rect 4264 11354 4292 15127
rect 4356 14890 4384 15370
rect 4632 15162 4660 15370
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4356 14006 4384 14554
rect 4724 14482 4752 14894
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4724 14074 4752 14418
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4342 13424 4398 13433
rect 4342 13359 4398 13368
rect 4356 13326 4384 13359
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4540 12782 4568 13466
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12918 4660 13330
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4724 12850 4752 13738
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 4724 12209 4752 12786
rect 4710 12200 4766 12209
rect 4816 12170 4844 15370
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4908 14278 4936 14894
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4908 13530 4936 13942
rect 5000 13802 5028 15574
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5092 14550 5120 14894
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 5080 14272 5132 14278
rect 5078 14240 5080 14249
rect 5132 14240 5134 14249
rect 5078 14175 5134 14184
rect 5184 13977 5212 16374
rect 5170 13968 5226 13977
rect 5170 13903 5226 13912
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4894 13424 4950 13433
rect 4894 13359 4896 13368
rect 4948 13359 4950 13368
rect 4896 13330 4948 13336
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4908 12374 4936 13126
rect 5000 12442 5028 13126
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 5092 12481 5120 12650
rect 5078 12472 5134 12481
rect 4988 12436 5040 12442
rect 5078 12407 5134 12416
rect 4988 12378 5040 12384
rect 4896 12368 4948 12374
rect 4948 12316 5212 12322
rect 4896 12310 5212 12316
rect 4908 12306 5212 12310
rect 4908 12300 5224 12306
rect 4908 12294 5172 12300
rect 5172 12242 5224 12248
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4710 12135 4766 12144
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 4724 11354 4752 12038
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4712 11212 4764 11218
rect 4816 11200 4844 11562
rect 4908 11354 4936 12174
rect 5276 12170 5304 17439
rect 5368 15026 5396 18362
rect 5460 17746 5488 18906
rect 5736 18902 5764 19751
rect 5828 19514 5856 20198
rect 5920 19922 5948 20352
rect 5908 19916 5960 19922
rect 5908 19858 5960 19864
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5920 19417 5948 19858
rect 6012 19514 6040 20538
rect 6104 20330 6132 20975
rect 6196 20584 6224 21422
rect 6288 21321 6316 21422
rect 6274 21312 6330 21321
rect 6274 21247 6330 21256
rect 6380 21078 6408 24006
rect 6368 21072 6420 21078
rect 6368 21014 6420 21020
rect 6196 20556 6316 20584
rect 6092 20324 6144 20330
rect 6092 20266 6144 20272
rect 6090 20088 6146 20097
rect 6090 20023 6146 20032
rect 6104 19990 6132 20023
rect 6092 19984 6144 19990
rect 6092 19926 6144 19932
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 5906 19408 5962 19417
rect 5828 19366 5906 19394
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5736 18737 5764 18838
rect 5722 18728 5778 18737
rect 5722 18663 5778 18672
rect 5538 18592 5594 18601
rect 5538 18527 5594 18536
rect 5552 18426 5580 18527
rect 5722 18456 5778 18465
rect 5540 18420 5592 18426
rect 5722 18391 5724 18400
rect 5540 18362 5592 18368
rect 5776 18391 5778 18400
rect 5724 18362 5776 18368
rect 5722 18320 5778 18329
rect 5828 18290 5856 19366
rect 5906 19343 5962 19352
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6012 18902 6040 19246
rect 6090 19000 6146 19009
rect 6090 18935 6146 18944
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 6104 18834 6132 18935
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 5920 18340 5948 18702
rect 6104 18630 6132 18770
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 6012 18358 6040 18566
rect 6090 18456 6146 18465
rect 6090 18391 6146 18400
rect 6000 18352 6052 18358
rect 5920 18312 5949 18340
rect 5722 18255 5724 18264
rect 5776 18255 5778 18264
rect 5816 18284 5868 18290
rect 5724 18226 5776 18232
rect 5816 18226 5868 18232
rect 5538 18184 5594 18193
rect 5538 18119 5594 18128
rect 5722 18184 5778 18193
rect 5921 18170 5949 18312
rect 6000 18294 6052 18300
rect 5722 18119 5778 18128
rect 5828 18142 5949 18170
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5460 16998 5488 17682
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 16833 5488 16934
rect 5446 16824 5502 16833
rect 5446 16759 5502 16768
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 14618 5396 14758
rect 5460 14618 5488 16118
rect 5552 15094 5580 18119
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5356 14408 5408 14414
rect 5552 14396 5580 15030
rect 5408 14368 5580 14396
rect 5356 14350 5408 14356
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 14006 5396 14214
rect 5356 14000 5408 14006
rect 5356 13942 5408 13948
rect 5448 14000 5500 14006
rect 5448 13942 5500 13948
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5368 12442 5396 12854
rect 5460 12782 5488 13942
rect 5644 13870 5672 17682
rect 5736 17649 5764 18119
rect 5828 18068 5856 18142
rect 5828 18040 5949 18068
rect 5921 17954 5949 18040
rect 5920 17926 5949 17954
rect 5920 17882 5948 17926
rect 5908 17876 5960 17882
rect 5908 17818 5960 17824
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 5722 17640 5778 17649
rect 5722 17575 5778 17584
rect 5736 17202 5764 17575
rect 5816 17264 5868 17270
rect 5816 17206 5868 17212
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5722 17096 5778 17105
rect 5722 17031 5778 17040
rect 5736 16794 5764 17031
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5828 16658 5856 17206
rect 5920 16697 5948 17682
rect 6012 17202 6040 18294
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6104 17134 6132 18391
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 6092 16992 6144 16998
rect 6012 16952 6092 16980
rect 5906 16688 5962 16697
rect 5816 16652 5868 16658
rect 6012 16658 6040 16952
rect 6092 16934 6144 16940
rect 5906 16623 5962 16632
rect 6000 16652 6052 16658
rect 5816 16594 5868 16600
rect 6000 16594 6052 16600
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5828 14958 5856 15438
rect 6104 15162 6132 16594
rect 6196 15706 6224 19790
rect 6288 19242 6316 20556
rect 6276 19236 6328 19242
rect 6276 19178 6328 19184
rect 6288 18970 6316 19178
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6380 18834 6408 21014
rect 6472 19310 6500 24511
rect 6564 24449 6592 24550
rect 6550 24440 6606 24449
rect 6550 24375 6606 24384
rect 6644 24404 6696 24410
rect 6644 24346 6696 24352
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 6564 23798 6592 24210
rect 6656 23798 6684 24346
rect 6748 24138 6776 25366
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6840 24018 6868 28999
rect 6932 28937 6960 29158
rect 7024 28994 7052 31719
rect 7196 31690 7248 31696
rect 7104 30728 7156 30734
rect 7104 30670 7156 30676
rect 7116 29850 7144 30670
rect 7208 30394 7236 31690
rect 7392 31482 7420 31826
rect 7484 31754 7512 32014
rect 7564 32020 7616 32026
rect 7564 31962 7616 31968
rect 7562 31920 7618 31929
rect 7668 31906 7696 33102
rect 7760 32065 7788 35022
rect 7840 34536 7892 34542
rect 7838 34504 7840 34513
rect 7892 34504 7894 34513
rect 7838 34439 7894 34448
rect 7838 34096 7894 34105
rect 7838 34031 7840 34040
rect 7892 34031 7894 34040
rect 7840 34002 7892 34008
rect 7852 33454 7880 34002
rect 7944 33538 7972 35278
rect 8024 35284 8076 35290
rect 8024 35226 8076 35232
rect 8220 35278 8432 35306
rect 8680 35290 8708 35974
rect 8772 35834 8800 36654
rect 8760 35828 8812 35834
rect 8760 35770 8812 35776
rect 8668 35284 8720 35290
rect 8220 35154 8248 35278
rect 8668 35226 8720 35232
rect 8298 35184 8354 35193
rect 8208 35148 8260 35154
rect 8864 35154 8892 37266
rect 8942 37224 8998 37233
rect 8942 37159 8944 37168
rect 8996 37159 8998 37168
rect 8944 37130 8996 37136
rect 8942 36408 8998 36417
rect 8942 36343 8998 36352
rect 8956 36310 8984 36343
rect 8944 36304 8996 36310
rect 8944 36246 8996 36252
rect 9048 36038 9076 37760
rect 9128 37742 9180 37748
rect 9128 37460 9180 37466
rect 9128 37402 9180 37408
rect 9140 36922 9168 37402
rect 9232 37398 9260 37964
rect 9416 37890 9444 37964
rect 9324 37862 9444 37890
rect 9324 37670 9352 37862
rect 9404 37800 9456 37806
rect 9508 37788 9536 38916
rect 9588 38898 9640 38904
rect 9692 38826 9720 39238
rect 9784 39098 9812 39578
rect 9968 39506 9996 39782
rect 9956 39500 10008 39506
rect 9956 39442 10008 39448
rect 10060 39302 10088 39986
rect 10152 39409 10180 40140
rect 10428 39914 10456 40394
rect 10520 40390 10548 42230
rect 10612 42226 10640 42706
rect 10600 42220 10652 42226
rect 10600 42162 10652 42168
rect 10722 41916 11030 41925
rect 10722 41914 10728 41916
rect 10784 41914 10808 41916
rect 10864 41914 10888 41916
rect 10944 41914 10968 41916
rect 11024 41914 11030 41916
rect 10784 41862 10786 41914
rect 10966 41862 10968 41914
rect 10722 41860 10728 41862
rect 10784 41860 10808 41862
rect 10864 41860 10888 41862
rect 10944 41860 10968 41862
rect 11024 41860 11030 41862
rect 10722 41851 11030 41860
rect 10692 41812 10744 41818
rect 10692 41754 10744 41760
rect 10600 41676 10652 41682
rect 10600 41618 10652 41624
rect 10508 40384 10560 40390
rect 10508 40326 10560 40332
rect 10416 39908 10468 39914
rect 10416 39850 10468 39856
rect 10232 39840 10284 39846
rect 10232 39782 10284 39788
rect 10244 39545 10272 39782
rect 10230 39536 10286 39545
rect 10230 39471 10286 39480
rect 10138 39400 10194 39409
rect 10138 39335 10194 39344
rect 10048 39296 10100 39302
rect 10048 39238 10100 39244
rect 10062 39196 10370 39205
rect 10062 39194 10068 39196
rect 10124 39194 10148 39196
rect 10204 39194 10228 39196
rect 10284 39194 10308 39196
rect 10364 39194 10370 39196
rect 10124 39142 10126 39194
rect 10306 39142 10308 39194
rect 10062 39140 10068 39142
rect 10124 39140 10148 39142
rect 10204 39140 10228 39142
rect 10284 39140 10308 39142
rect 10364 39140 10370 39142
rect 10062 39131 10370 39140
rect 9772 39092 9824 39098
rect 9772 39034 9824 39040
rect 9956 39024 10008 39030
rect 9862 38992 9918 39001
rect 9956 38966 10008 38972
rect 9862 38927 9918 38936
rect 9876 38894 9904 38927
rect 9864 38888 9916 38894
rect 9770 38856 9826 38865
rect 9680 38820 9732 38826
rect 9864 38830 9916 38836
rect 9770 38791 9826 38800
rect 9680 38762 9732 38768
rect 9680 38480 9732 38486
rect 9680 38422 9732 38428
rect 9588 38004 9640 38010
rect 9588 37946 9640 37952
rect 9600 37913 9628 37946
rect 9586 37904 9642 37913
rect 9586 37839 9642 37848
rect 9456 37760 9536 37788
rect 9404 37742 9456 37748
rect 9312 37664 9364 37670
rect 9404 37664 9456 37670
rect 9312 37606 9364 37612
rect 9402 37632 9404 37641
rect 9456 37632 9458 37641
rect 9402 37567 9458 37576
rect 9310 37496 9366 37505
rect 9310 37431 9366 37440
rect 9220 37392 9272 37398
rect 9220 37334 9272 37340
rect 9128 36916 9180 36922
rect 9128 36858 9180 36864
rect 9324 36718 9352 37431
rect 9402 37224 9458 37233
rect 9402 37159 9458 37168
rect 9128 36712 9180 36718
rect 9128 36654 9180 36660
rect 9312 36712 9364 36718
rect 9312 36654 9364 36660
rect 9140 36378 9168 36654
rect 9220 36576 9272 36582
rect 9218 36544 9220 36553
rect 9272 36544 9274 36553
rect 9218 36479 9274 36488
rect 9128 36372 9180 36378
rect 9128 36314 9180 36320
rect 9128 36236 9180 36242
rect 9128 36178 9180 36184
rect 9036 36032 9088 36038
rect 9036 35974 9088 35980
rect 9036 35692 9088 35698
rect 9036 35634 9088 35640
rect 8944 35624 8996 35630
rect 8944 35566 8996 35572
rect 8956 35154 8984 35566
rect 9048 35290 9076 35634
rect 9140 35306 9168 36178
rect 9220 35828 9272 35834
rect 9220 35770 9272 35776
rect 9232 35698 9260 35770
rect 9220 35692 9272 35698
rect 9220 35634 9272 35640
rect 9036 35284 9088 35290
rect 9140 35278 9260 35306
rect 9036 35226 9088 35232
rect 8298 35119 8300 35128
rect 8208 35090 8260 35096
rect 8352 35119 8354 35128
rect 8852 35148 8904 35154
rect 8300 35090 8352 35096
rect 8852 35090 8904 35096
rect 8944 35148 8996 35154
rect 8944 35090 8996 35096
rect 8760 35080 8812 35086
rect 8864 35057 8892 35090
rect 8760 35022 8812 35028
rect 8850 35048 8906 35057
rect 8208 35012 8260 35018
rect 8208 34954 8260 34960
rect 8024 34944 8076 34950
rect 8024 34886 8076 34892
rect 8036 34542 8064 34886
rect 8024 34536 8076 34542
rect 8024 34478 8076 34484
rect 8116 34536 8168 34542
rect 8116 34478 8168 34484
rect 7944 33510 8064 33538
rect 7840 33448 7892 33454
rect 7840 33390 7892 33396
rect 7932 33448 7984 33454
rect 7932 33390 7984 33396
rect 7840 33312 7892 33318
rect 7944 33289 7972 33390
rect 7840 33254 7892 33260
rect 7930 33280 7986 33289
rect 7852 32774 7880 33254
rect 7930 33215 7986 33224
rect 8036 33046 8064 33510
rect 8024 33040 8076 33046
rect 8024 32982 8076 32988
rect 7932 32904 7984 32910
rect 7932 32846 7984 32852
rect 8024 32904 8076 32910
rect 8024 32846 8076 32852
rect 7840 32768 7892 32774
rect 7840 32710 7892 32716
rect 7944 32609 7972 32846
rect 8036 32745 8064 32846
rect 8022 32736 8078 32745
rect 8022 32671 8078 32680
rect 7930 32600 7986 32609
rect 7840 32564 7892 32570
rect 7930 32535 7986 32544
rect 7840 32506 7892 32512
rect 7746 32056 7802 32065
rect 7852 32026 7880 32506
rect 8036 32502 8064 32671
rect 8024 32496 8076 32502
rect 8024 32438 8076 32444
rect 7932 32224 7984 32230
rect 7984 32184 8064 32212
rect 7932 32166 7984 32172
rect 7746 31991 7802 32000
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 7668 31878 7972 31906
rect 7562 31855 7564 31864
rect 7616 31855 7618 31864
rect 7564 31826 7616 31832
rect 7484 31726 7788 31754
rect 7564 31680 7616 31686
rect 7564 31622 7616 31628
rect 7470 31512 7526 31521
rect 7380 31476 7432 31482
rect 7576 31482 7604 31622
rect 7470 31447 7526 31456
rect 7564 31476 7616 31482
rect 7380 31418 7432 31424
rect 7380 31136 7432 31142
rect 7380 31078 7432 31084
rect 7392 30938 7420 31078
rect 7380 30932 7432 30938
rect 7380 30874 7432 30880
rect 7288 30864 7340 30870
rect 7288 30806 7340 30812
rect 7196 30388 7248 30394
rect 7196 30330 7248 30336
rect 7194 30288 7250 30297
rect 7194 30223 7196 30232
rect 7248 30223 7250 30232
rect 7196 30194 7248 30200
rect 7104 29844 7156 29850
rect 7104 29786 7156 29792
rect 7102 29608 7158 29617
rect 7102 29543 7158 29552
rect 7116 29510 7144 29543
rect 7104 29504 7156 29510
rect 7104 29446 7156 29452
rect 7196 29504 7248 29510
rect 7300 29481 7328 30806
rect 7484 30682 7512 31447
rect 7564 31418 7616 31424
rect 7656 31340 7708 31346
rect 7656 31282 7708 31288
rect 7562 30832 7618 30841
rect 7562 30767 7564 30776
rect 7616 30767 7618 30776
rect 7564 30738 7616 30744
rect 7392 30654 7512 30682
rect 7564 30660 7616 30666
rect 7196 29446 7248 29452
rect 7286 29472 7342 29481
rect 7102 29336 7158 29345
rect 7102 29271 7104 29280
rect 7156 29271 7158 29280
rect 7104 29242 7156 29248
rect 7208 29186 7236 29446
rect 7286 29407 7342 29416
rect 7116 29158 7236 29186
rect 7288 29232 7340 29238
rect 7288 29174 7340 29180
rect 7116 29102 7144 29158
rect 7104 29096 7156 29102
rect 7196 29096 7248 29102
rect 7104 29038 7156 29044
rect 7194 29064 7196 29073
rect 7248 29064 7250 29073
rect 7194 28999 7250 29008
rect 7024 28966 7144 28994
rect 6918 28928 6974 28937
rect 6918 28863 6974 28872
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 6932 28529 6960 28698
rect 7012 28620 7064 28626
rect 7012 28562 7064 28568
rect 6918 28520 6974 28529
rect 6918 28455 6974 28464
rect 7024 28082 7052 28562
rect 7116 28393 7144 28966
rect 7196 28688 7248 28694
rect 7196 28630 7248 28636
rect 7102 28384 7158 28393
rect 7102 28319 7158 28328
rect 7012 28076 7064 28082
rect 7012 28018 7064 28024
rect 6918 27976 6974 27985
rect 6918 27911 6920 27920
rect 6972 27911 6974 27920
rect 7104 27940 7156 27946
rect 6920 27882 6972 27888
rect 7104 27882 7156 27888
rect 6932 27470 6960 27882
rect 6920 27464 6972 27470
rect 6920 27406 6972 27412
rect 6920 27124 6972 27130
rect 6920 27066 6972 27072
rect 6932 26926 6960 27066
rect 7116 26926 7144 27882
rect 7208 27849 7236 28630
rect 7194 27840 7250 27849
rect 7194 27775 7250 27784
rect 7300 27577 7328 29174
rect 7392 28529 7420 30654
rect 7564 30602 7616 30608
rect 7472 30592 7524 30598
rect 7472 30534 7524 30540
rect 7484 30433 7512 30534
rect 7470 30424 7526 30433
rect 7470 30359 7526 30368
rect 7472 30048 7524 30054
rect 7472 29990 7524 29996
rect 7484 29714 7512 29990
rect 7472 29708 7524 29714
rect 7472 29650 7524 29656
rect 7472 29572 7524 29578
rect 7472 29514 7524 29520
rect 7378 28520 7434 28529
rect 7378 28455 7434 28464
rect 7380 28416 7432 28422
rect 7380 28358 7432 28364
rect 7392 27713 7420 28358
rect 7484 27878 7512 29514
rect 7472 27872 7524 27878
rect 7472 27814 7524 27820
rect 7378 27704 7434 27713
rect 7378 27639 7434 27648
rect 7380 27600 7432 27606
rect 7286 27568 7342 27577
rect 7196 27532 7248 27538
rect 7484 27554 7512 27814
rect 7432 27548 7512 27554
rect 7380 27542 7512 27548
rect 7392 27526 7512 27542
rect 7286 27503 7342 27512
rect 7196 27474 7248 27480
rect 7208 27130 7236 27474
rect 7300 27130 7328 27503
rect 7196 27124 7248 27130
rect 7196 27066 7248 27072
rect 7288 27124 7340 27130
rect 7288 27066 7340 27072
rect 7472 27124 7524 27130
rect 7472 27066 7524 27072
rect 7208 27033 7236 27066
rect 7380 27056 7432 27062
rect 7194 27024 7250 27033
rect 7380 26998 7432 27004
rect 7194 26959 7250 26968
rect 6920 26920 6972 26926
rect 7104 26920 7156 26926
rect 6920 26862 6972 26868
rect 7010 26888 7066 26897
rect 7104 26862 7156 26868
rect 7196 26920 7248 26926
rect 7196 26862 7248 26868
rect 7010 26823 7066 26832
rect 6918 26752 6974 26761
rect 6918 26687 6974 26696
rect 6932 25498 6960 26687
rect 7024 26518 7052 26823
rect 7012 26512 7064 26518
rect 7012 26454 7064 26460
rect 7012 26036 7064 26042
rect 7012 25978 7064 25984
rect 7024 25537 7052 25978
rect 7010 25528 7066 25537
rect 6920 25492 6972 25498
rect 7010 25463 7066 25472
rect 6920 25434 6972 25440
rect 6918 25392 6974 25401
rect 6918 25327 6974 25336
rect 7012 25356 7064 25362
rect 6932 24562 6960 25327
rect 7012 25298 7064 25304
rect 7024 24954 7052 25298
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 6932 24534 7052 24562
rect 6918 24440 6974 24449
rect 7024 24410 7052 24534
rect 6918 24375 6920 24384
rect 6972 24375 6974 24384
rect 7012 24404 7064 24410
rect 6920 24346 6972 24352
rect 7012 24346 7064 24352
rect 6932 24041 6960 24346
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 6748 23990 6868 24018
rect 6918 24032 6974 24041
rect 6552 23792 6604 23798
rect 6552 23734 6604 23740
rect 6644 23792 6696 23798
rect 6644 23734 6696 23740
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6644 23656 6696 23662
rect 6644 23598 6696 23604
rect 6564 23526 6592 23598
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6564 22982 6592 23462
rect 6552 22976 6604 22982
rect 6552 22918 6604 22924
rect 6656 22778 6684 23598
rect 6748 22794 6776 23990
rect 6918 23967 6974 23976
rect 6920 23588 6972 23594
rect 6920 23530 6972 23536
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 6840 22953 6868 23122
rect 6932 23118 6960 23530
rect 7024 23322 7052 24210
rect 7116 23848 7144 26862
rect 7208 26790 7236 26862
rect 7196 26784 7248 26790
rect 7196 26726 7248 26732
rect 7288 26784 7340 26790
rect 7288 26726 7340 26732
rect 7194 26480 7250 26489
rect 7194 26415 7196 26424
rect 7248 26415 7250 26424
rect 7196 26386 7248 26392
rect 7196 26240 7248 26246
rect 7196 26182 7248 26188
rect 7208 25838 7236 26182
rect 7300 25906 7328 26726
rect 7288 25900 7340 25906
rect 7392 25888 7420 26998
rect 7484 26246 7512 27066
rect 7576 26450 7604 30602
rect 7668 29714 7696 31282
rect 7760 30870 7788 31726
rect 7840 31408 7892 31414
rect 7840 31350 7892 31356
rect 7748 30864 7800 30870
rect 7748 30806 7800 30812
rect 7760 30161 7788 30806
rect 7746 30152 7802 30161
rect 7746 30087 7802 30096
rect 7748 30048 7800 30054
rect 7748 29990 7800 29996
rect 7656 29708 7708 29714
rect 7656 29650 7708 29656
rect 7760 29646 7788 29990
rect 7852 29714 7880 31350
rect 7944 30190 7972 31878
rect 7932 30184 7984 30190
rect 7932 30126 7984 30132
rect 7840 29708 7892 29714
rect 7840 29650 7892 29656
rect 7748 29640 7800 29646
rect 7748 29582 7800 29588
rect 7838 29608 7894 29617
rect 7838 29543 7894 29552
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 7654 28656 7710 28665
rect 7654 28591 7656 28600
rect 7708 28591 7710 28600
rect 7656 28562 7708 28568
rect 7656 28416 7708 28422
rect 7656 28358 7708 28364
rect 7668 27538 7696 28358
rect 7656 27532 7708 27538
rect 7656 27474 7708 27480
rect 7656 27328 7708 27334
rect 7656 27270 7708 27276
rect 7668 26858 7696 27270
rect 7760 26994 7788 28970
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7656 26852 7708 26858
rect 7656 26794 7708 26800
rect 7748 26852 7800 26858
rect 7748 26794 7800 26800
rect 7564 26444 7616 26450
rect 7564 26386 7616 26392
rect 7472 26240 7524 26246
rect 7470 26208 7472 26217
rect 7524 26208 7604 26228
rect 7526 26200 7604 26208
rect 7470 26143 7526 26152
rect 7576 25974 7604 26200
rect 7564 25968 7616 25974
rect 7564 25910 7616 25916
rect 7392 25860 7512 25888
rect 7288 25842 7340 25848
rect 7196 25832 7248 25838
rect 7196 25774 7248 25780
rect 7208 25362 7236 25774
rect 7380 25764 7432 25770
rect 7380 25706 7432 25712
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 7300 25498 7328 25638
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 7392 25378 7420 25706
rect 7196 25356 7248 25362
rect 7196 25298 7248 25304
rect 7300 25350 7420 25378
rect 7208 24750 7236 25298
rect 7300 24834 7328 25350
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7392 25129 7420 25230
rect 7378 25120 7434 25129
rect 7378 25055 7434 25064
rect 7484 24993 7512 25860
rect 7564 25832 7616 25838
rect 7564 25774 7616 25780
rect 7576 25362 7604 25774
rect 7668 25498 7696 26794
rect 7760 26586 7788 26794
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7852 26024 7880 29543
rect 7944 26217 7972 30126
rect 8036 29170 8064 32184
rect 8128 31657 8156 34478
rect 8220 33998 8248 34954
rect 8392 34672 8444 34678
rect 8392 34614 8444 34620
rect 8574 34640 8630 34649
rect 8404 34542 8432 34614
rect 8574 34575 8630 34584
rect 8588 34542 8616 34575
rect 8392 34536 8444 34542
rect 8576 34536 8628 34542
rect 8392 34478 8444 34484
rect 8482 34504 8538 34513
rect 8576 34478 8628 34484
rect 8668 34536 8720 34542
rect 8668 34478 8720 34484
rect 8482 34439 8538 34448
rect 8392 34400 8444 34406
rect 8392 34342 8444 34348
rect 8208 33992 8260 33998
rect 8206 33960 8208 33969
rect 8260 33960 8262 33969
rect 8206 33895 8262 33904
rect 8208 33856 8260 33862
rect 8208 33798 8260 33804
rect 8220 33674 8248 33798
rect 8220 33658 8340 33674
rect 8220 33652 8352 33658
rect 8220 33646 8300 33652
rect 8300 33594 8352 33600
rect 8206 33552 8262 33561
rect 8206 33487 8262 33496
rect 8220 32570 8248 33487
rect 8300 33450 8352 33456
rect 8404 33454 8432 34342
rect 8496 34066 8524 34439
rect 8680 34134 8708 34478
rect 8772 34474 8800 35022
rect 8850 34983 8906 34992
rect 8956 34746 8984 35090
rect 8944 34740 8996 34746
rect 8944 34682 8996 34688
rect 8760 34468 8812 34474
rect 8760 34410 8812 34416
rect 8956 34202 8984 34682
rect 8852 34196 8904 34202
rect 8852 34138 8904 34144
rect 8944 34196 8996 34202
rect 8944 34138 8996 34144
rect 8668 34128 8720 34134
rect 8574 34096 8630 34105
rect 8484 34060 8536 34066
rect 8864 34105 8892 34138
rect 8668 34070 8720 34076
rect 8850 34096 8906 34105
rect 8574 34031 8630 34040
rect 8760 34060 8812 34066
rect 8484 34002 8536 34008
rect 8588 33946 8616 34031
rect 9048 34066 9076 35226
rect 9128 35216 9180 35222
rect 9128 35158 9180 35164
rect 8850 34031 8906 34040
rect 8944 34060 8996 34066
rect 8760 34002 8812 34008
rect 8944 34002 8996 34008
rect 9036 34060 9088 34066
rect 9036 34002 9088 34008
rect 8772 33969 8800 34002
rect 8852 33992 8904 33998
rect 8496 33918 8616 33946
rect 8758 33960 8814 33969
rect 8300 33392 8352 33398
rect 8392 33448 8444 33454
rect 8312 33046 8340 33392
rect 8392 33390 8444 33396
rect 8390 33280 8446 33289
rect 8496 33266 8524 33918
rect 8852 33934 8904 33940
rect 8758 33895 8814 33904
rect 8760 33856 8812 33862
rect 8760 33798 8812 33804
rect 8668 33652 8720 33658
rect 8668 33594 8720 33600
rect 8574 33552 8630 33561
rect 8574 33487 8630 33496
rect 8588 33386 8616 33487
rect 8576 33380 8628 33386
rect 8576 33322 8628 33328
rect 8446 33238 8524 33266
rect 8390 33215 8446 33224
rect 8300 33040 8352 33046
rect 8300 32982 8352 32988
rect 8404 32978 8432 33215
rect 8680 32978 8708 33594
rect 8772 33289 8800 33798
rect 8758 33280 8814 33289
rect 8758 33215 8814 33224
rect 8758 33144 8814 33153
rect 8864 33114 8892 33934
rect 8758 33079 8814 33088
rect 8852 33108 8904 33114
rect 8772 32978 8800 33079
rect 8852 33050 8904 33056
rect 8392 32972 8444 32978
rect 8392 32914 8444 32920
rect 8668 32972 8720 32978
rect 8668 32914 8720 32920
rect 8760 32972 8812 32978
rect 8760 32914 8812 32920
rect 8300 32904 8352 32910
rect 8404 32881 8432 32914
rect 8300 32846 8352 32852
rect 8390 32872 8446 32881
rect 8208 32564 8260 32570
rect 8208 32506 8260 32512
rect 8312 32366 8340 32846
rect 8390 32807 8446 32816
rect 8576 32768 8628 32774
rect 8482 32736 8538 32745
rect 8576 32710 8628 32716
rect 8482 32671 8538 32680
rect 8300 32360 8352 32366
rect 8300 32302 8352 32308
rect 8208 32292 8260 32298
rect 8208 32234 8260 32240
rect 8392 32292 8444 32298
rect 8392 32234 8444 32240
rect 8220 31754 8248 32234
rect 8298 32056 8354 32065
rect 8298 31991 8300 32000
rect 8352 31991 8354 32000
rect 8300 31962 8352 31968
rect 8220 31726 8340 31754
rect 8208 31680 8260 31686
rect 8114 31648 8170 31657
rect 8208 31622 8260 31628
rect 8114 31583 8170 31592
rect 8128 31278 8156 31583
rect 8116 31272 8168 31278
rect 8116 31214 8168 31220
rect 8220 31142 8248 31622
rect 8312 31142 8340 31726
rect 8404 31482 8432 32234
rect 8392 31476 8444 31482
rect 8392 31418 8444 31424
rect 8404 31210 8432 31418
rect 8392 31204 8444 31210
rect 8392 31146 8444 31152
rect 8208 31136 8260 31142
rect 8208 31078 8260 31084
rect 8300 31136 8352 31142
rect 8300 31078 8352 31084
rect 8116 30796 8168 30802
rect 8116 30738 8168 30744
rect 8024 29164 8076 29170
rect 8024 29106 8076 29112
rect 8024 29028 8076 29034
rect 8024 28970 8076 28976
rect 8036 28937 8064 28970
rect 8022 28928 8078 28937
rect 8022 28863 8078 28872
rect 8036 27577 8064 28863
rect 8128 27946 8156 30738
rect 8220 30326 8248 31078
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 8312 30394 8340 30738
rect 8404 30598 8432 31146
rect 8392 30592 8444 30598
rect 8392 30534 8444 30540
rect 8496 30410 8524 32671
rect 8588 31414 8616 32710
rect 8680 32502 8708 32914
rect 8668 32496 8720 32502
rect 8668 32438 8720 32444
rect 8668 32360 8720 32366
rect 8668 32302 8720 32308
rect 8680 31804 8708 32302
rect 8864 32298 8892 33050
rect 8956 32609 8984 34002
rect 9036 33312 9088 33318
rect 9036 33254 9088 33260
rect 9048 33046 9076 33254
rect 9036 33040 9088 33046
rect 9036 32982 9088 32988
rect 8942 32600 8998 32609
rect 8942 32535 8998 32544
rect 9036 32496 9088 32502
rect 9036 32438 9088 32444
rect 8944 32360 8996 32366
rect 9048 32337 9076 32438
rect 8944 32302 8996 32308
rect 9034 32328 9090 32337
rect 8852 32292 8904 32298
rect 8852 32234 8904 32240
rect 8956 32178 8984 32302
rect 9140 32298 9168 35158
rect 9232 34728 9260 35278
rect 9324 35018 9352 36654
rect 9416 36242 9444 37159
rect 9508 36582 9536 37760
rect 9692 36854 9720 38422
rect 9784 38214 9812 38791
rect 9876 38554 9904 38830
rect 9864 38548 9916 38554
rect 9864 38490 9916 38496
rect 9968 38332 9996 38966
rect 10140 38888 10192 38894
rect 10138 38856 10140 38865
rect 10192 38856 10194 38865
rect 10138 38791 10194 38800
rect 10232 38752 10284 38758
rect 10232 38694 10284 38700
rect 10416 38752 10468 38758
rect 10416 38694 10468 38700
rect 10048 38344 10100 38350
rect 9968 38304 10048 38332
rect 10048 38286 10100 38292
rect 10244 38214 10272 38694
rect 10322 38584 10378 38593
rect 10322 38519 10378 38528
rect 10336 38214 10364 38519
rect 9772 38208 9824 38214
rect 9772 38150 9824 38156
rect 9956 38208 10008 38214
rect 9956 38150 10008 38156
rect 10232 38208 10284 38214
rect 10232 38150 10284 38156
rect 10324 38208 10376 38214
rect 10324 38150 10376 38156
rect 9784 37777 9812 38150
rect 9862 38040 9918 38049
rect 9862 37975 9918 37984
rect 9876 37874 9904 37975
rect 9864 37868 9916 37874
rect 9864 37810 9916 37816
rect 9968 37806 9996 38150
rect 10062 38108 10370 38117
rect 10062 38106 10068 38108
rect 10124 38106 10148 38108
rect 10204 38106 10228 38108
rect 10284 38106 10308 38108
rect 10364 38106 10370 38108
rect 10124 38054 10126 38106
rect 10306 38054 10308 38106
rect 10062 38052 10068 38054
rect 10124 38052 10148 38054
rect 10204 38052 10228 38054
rect 10284 38052 10308 38054
rect 10364 38052 10370 38054
rect 10062 38043 10370 38052
rect 9956 37800 10008 37806
rect 9770 37768 9826 37777
rect 9956 37742 10008 37748
rect 10428 37738 10456 38694
rect 10520 38418 10548 40326
rect 10612 39982 10640 41618
rect 10704 40934 10732 41754
rect 11060 41744 11112 41750
rect 11060 41686 11112 41692
rect 10692 40928 10744 40934
rect 10692 40870 10744 40876
rect 10722 40828 11030 40837
rect 10722 40826 10728 40828
rect 10784 40826 10808 40828
rect 10864 40826 10888 40828
rect 10944 40826 10968 40828
rect 11024 40826 11030 40828
rect 10784 40774 10786 40826
rect 10966 40774 10968 40826
rect 10722 40772 10728 40774
rect 10784 40772 10808 40774
rect 10864 40772 10888 40774
rect 10944 40772 10968 40774
rect 11024 40772 11030 40774
rect 10722 40763 11030 40772
rect 10692 40588 10744 40594
rect 10692 40530 10744 40536
rect 10704 40089 10732 40530
rect 10690 40080 10746 40089
rect 11072 40050 11100 41686
rect 11244 40112 11296 40118
rect 11244 40054 11296 40060
rect 10690 40015 10746 40024
rect 11060 40044 11112 40050
rect 11060 39986 11112 39992
rect 10600 39976 10652 39982
rect 10600 39918 10652 39924
rect 10690 39944 10746 39953
rect 10508 38412 10560 38418
rect 10508 38354 10560 38360
rect 10508 38276 10560 38282
rect 10508 38218 10560 38224
rect 10520 37942 10548 38218
rect 10508 37936 10560 37942
rect 10508 37878 10560 37884
rect 10508 37800 10560 37806
rect 10508 37742 10560 37748
rect 9770 37703 9826 37712
rect 9864 37732 9916 37738
rect 9864 37674 9916 37680
rect 10416 37732 10468 37738
rect 10416 37674 10468 37680
rect 9770 37360 9826 37369
rect 9770 37295 9826 37304
rect 9680 36848 9732 36854
rect 9680 36790 9732 36796
rect 9496 36576 9548 36582
rect 9496 36518 9548 36524
rect 9680 36576 9732 36582
rect 9680 36518 9732 36524
rect 9494 36408 9550 36417
rect 9494 36343 9550 36352
rect 9508 36242 9536 36343
rect 9404 36236 9456 36242
rect 9404 36178 9456 36184
rect 9496 36236 9548 36242
rect 9496 36178 9548 36184
rect 9312 35012 9364 35018
rect 9312 34954 9364 34960
rect 9312 34740 9364 34746
rect 9232 34700 9312 34728
rect 9232 34649 9260 34700
rect 9312 34682 9364 34688
rect 9218 34640 9274 34649
rect 9218 34575 9274 34584
rect 9218 34504 9274 34513
rect 9416 34474 9444 36178
rect 9692 36038 9720 36518
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 9680 35624 9732 35630
rect 9680 35566 9732 35572
rect 9784 35578 9812 37295
rect 9876 36922 9904 37674
rect 10520 37126 10548 37742
rect 10508 37120 10560 37126
rect 10508 37062 10560 37068
rect 10062 37020 10370 37029
rect 10062 37018 10068 37020
rect 10124 37018 10148 37020
rect 10204 37018 10228 37020
rect 10284 37018 10308 37020
rect 10364 37018 10370 37020
rect 10124 36966 10126 37018
rect 10306 36966 10308 37018
rect 10062 36964 10068 36966
rect 10124 36964 10148 36966
rect 10204 36964 10228 36966
rect 10284 36964 10308 36966
rect 10364 36964 10370 36966
rect 10062 36955 10370 36964
rect 9864 36916 9916 36922
rect 9864 36858 9916 36864
rect 10324 36916 10376 36922
rect 10324 36858 10376 36864
rect 9876 36689 9904 36858
rect 10140 36712 10192 36718
rect 9862 36680 9918 36689
rect 10140 36654 10192 36660
rect 9862 36615 9864 36624
rect 9916 36615 9918 36624
rect 9864 36586 9916 36592
rect 9956 36576 10008 36582
rect 9956 36518 10008 36524
rect 9968 36242 9996 36518
rect 9956 36236 10008 36242
rect 9956 36178 10008 36184
rect 10152 36122 10180 36654
rect 10336 36378 10364 36858
rect 10520 36650 10548 37062
rect 10612 36854 10640 39918
rect 10690 39879 10692 39888
rect 10744 39879 10746 39888
rect 10692 39850 10744 39856
rect 10722 39740 11030 39749
rect 10722 39738 10728 39740
rect 10784 39738 10808 39740
rect 10864 39738 10888 39740
rect 10944 39738 10968 39740
rect 11024 39738 11030 39740
rect 10784 39686 10786 39738
rect 10966 39686 10968 39738
rect 10722 39684 10728 39686
rect 10784 39684 10808 39686
rect 10864 39684 10888 39686
rect 10944 39684 10968 39686
rect 11024 39684 11030 39686
rect 10722 39675 11030 39684
rect 11072 39642 11100 39986
rect 11152 39908 11204 39914
rect 11152 39850 11204 39856
rect 11060 39636 11112 39642
rect 11060 39578 11112 39584
rect 10722 38652 11030 38661
rect 10722 38650 10728 38652
rect 10784 38650 10808 38652
rect 10864 38650 10888 38652
rect 10944 38650 10968 38652
rect 11024 38650 11030 38652
rect 10784 38598 10786 38650
rect 10966 38598 10968 38650
rect 10722 38596 10728 38598
rect 10784 38596 10808 38598
rect 10864 38596 10888 38598
rect 10944 38596 10968 38598
rect 11024 38596 11030 38598
rect 10722 38587 11030 38596
rect 11060 38208 11112 38214
rect 11060 38150 11112 38156
rect 10722 37564 11030 37573
rect 10722 37562 10728 37564
rect 10784 37562 10808 37564
rect 10864 37562 10888 37564
rect 10944 37562 10968 37564
rect 11024 37562 11030 37564
rect 10784 37510 10786 37562
rect 10966 37510 10968 37562
rect 10722 37508 10728 37510
rect 10784 37508 10808 37510
rect 10864 37508 10888 37510
rect 10944 37508 10968 37510
rect 11024 37508 11030 37510
rect 10722 37499 11030 37508
rect 11072 37330 11100 38150
rect 11060 37324 11112 37330
rect 11060 37266 11112 37272
rect 10600 36848 10652 36854
rect 10600 36790 10652 36796
rect 10692 36712 10744 36718
rect 10612 36660 10692 36666
rect 10612 36654 10744 36660
rect 10508 36644 10560 36650
rect 10508 36586 10560 36592
rect 10612 36638 10732 36654
rect 10324 36372 10376 36378
rect 10324 36314 10376 36320
rect 10612 36145 10640 36638
rect 10722 36476 11030 36485
rect 10722 36474 10728 36476
rect 10784 36474 10808 36476
rect 10864 36474 10888 36476
rect 10944 36474 10968 36476
rect 11024 36474 11030 36476
rect 10784 36422 10786 36474
rect 10966 36422 10968 36474
rect 10722 36420 10728 36422
rect 10784 36420 10808 36422
rect 10864 36420 10888 36422
rect 10944 36420 10968 36422
rect 11024 36420 11030 36422
rect 10722 36411 11030 36420
rect 9968 36094 10180 36122
rect 10598 36136 10654 36145
rect 9496 35488 9548 35494
rect 9496 35430 9548 35436
rect 9588 35488 9640 35494
rect 9588 35430 9640 35436
rect 9218 34439 9274 34448
rect 9404 34468 9456 34474
rect 9232 33590 9260 34439
rect 9404 34410 9456 34416
rect 9404 34196 9456 34202
rect 9404 34138 9456 34144
rect 9312 33924 9364 33930
rect 9312 33866 9364 33872
rect 9324 33658 9352 33866
rect 9312 33652 9364 33658
rect 9312 33594 9364 33600
rect 9220 33584 9272 33590
rect 9220 33526 9272 33532
rect 9312 33380 9364 33386
rect 9312 33322 9364 33328
rect 9220 33312 9272 33318
rect 9218 33280 9220 33289
rect 9272 33280 9274 33289
rect 9218 33215 9274 33224
rect 9034 32263 9090 32272
rect 9128 32292 9180 32298
rect 8864 32150 8984 32178
rect 8864 31822 8892 32150
rect 8942 32056 8998 32065
rect 9048 32042 9076 32263
rect 9128 32234 9180 32240
rect 9048 32014 9168 32042
rect 8942 31991 8998 32000
rect 8956 31958 8984 31991
rect 8944 31952 8996 31958
rect 8944 31894 8996 31900
rect 8852 31816 8904 31822
rect 8680 31793 8800 31804
rect 8680 31784 8814 31793
rect 8680 31776 8758 31784
rect 8852 31758 8904 31764
rect 8758 31719 8814 31728
rect 8668 31680 8720 31686
rect 8668 31622 8720 31628
rect 8576 31408 8628 31414
rect 8576 31350 8628 31356
rect 8576 31204 8628 31210
rect 8576 31146 8628 31152
rect 8300 30388 8352 30394
rect 8300 30330 8352 30336
rect 8404 30382 8524 30410
rect 8208 30320 8260 30326
rect 8208 30262 8260 30268
rect 8208 30184 8260 30190
rect 8208 30126 8260 30132
rect 8220 29850 8248 30126
rect 8300 30116 8352 30122
rect 8300 30058 8352 30064
rect 8208 29844 8260 29850
rect 8208 29786 8260 29792
rect 8206 29472 8262 29481
rect 8206 29407 8262 29416
rect 8220 29306 8248 29407
rect 8208 29300 8260 29306
rect 8208 29242 8260 29248
rect 8208 28620 8260 28626
rect 8208 28562 8260 28568
rect 8220 28393 8248 28562
rect 8312 28490 8340 30058
rect 8404 29238 8432 30382
rect 8484 30116 8536 30122
rect 8484 30058 8536 30064
rect 8392 29232 8444 29238
rect 8392 29174 8444 29180
rect 8392 29028 8444 29034
rect 8392 28970 8444 28976
rect 8404 28626 8432 28970
rect 8392 28620 8444 28626
rect 8392 28562 8444 28568
rect 8300 28484 8352 28490
rect 8300 28426 8352 28432
rect 8206 28384 8262 28393
rect 8206 28319 8262 28328
rect 8206 28248 8262 28257
rect 8206 28183 8262 28192
rect 8220 28150 8248 28183
rect 8208 28144 8260 28150
rect 8208 28086 8260 28092
rect 8208 28008 8260 28014
rect 8208 27950 8260 27956
rect 8116 27940 8168 27946
rect 8116 27882 8168 27888
rect 8022 27568 8078 27577
rect 8022 27503 8078 27512
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 8036 27062 8064 27406
rect 8128 27334 8156 27882
rect 8220 27713 8248 27950
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8206 27704 8262 27713
rect 8206 27639 8262 27648
rect 8312 27402 8340 27814
rect 8300 27396 8352 27402
rect 8300 27338 8352 27344
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 8114 27160 8170 27169
rect 8114 27095 8170 27104
rect 8024 27056 8076 27062
rect 8024 26998 8076 27004
rect 8024 26920 8076 26926
rect 8024 26862 8076 26868
rect 8036 26489 8064 26862
rect 8022 26480 8078 26489
rect 8128 26450 8156 27095
rect 8312 26926 8340 27338
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 8208 26852 8260 26858
rect 8208 26794 8260 26800
rect 8022 26415 8078 26424
rect 8116 26444 8168 26450
rect 7930 26208 7986 26217
rect 7930 26143 7986 26152
rect 7852 25996 7972 26024
rect 7838 25936 7894 25945
rect 7838 25871 7894 25880
rect 7852 25838 7880 25871
rect 7840 25832 7892 25838
rect 7760 25792 7840 25820
rect 7656 25492 7708 25498
rect 7656 25434 7708 25440
rect 7656 25390 7708 25396
rect 7564 25356 7616 25362
rect 7760 25362 7788 25792
rect 7840 25774 7892 25780
rect 7656 25332 7708 25338
rect 7748 25356 7800 25362
rect 7564 25298 7616 25304
rect 7668 25242 7696 25332
rect 7944 25344 7972 25996
rect 8036 25820 8064 26415
rect 8116 26386 8168 26392
rect 8128 25922 8156 26386
rect 8220 26042 8248 26794
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8312 26042 8340 26386
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 8128 25894 8248 25922
rect 8036 25792 8156 25820
rect 8024 25696 8076 25702
rect 8024 25638 8076 25644
rect 7748 25298 7800 25304
rect 7852 25316 7972 25344
rect 7576 25214 7696 25242
rect 7470 24984 7526 24993
rect 7470 24919 7526 24928
rect 7470 24848 7526 24857
rect 7300 24806 7420 24834
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7300 24392 7328 24686
rect 7392 24614 7420 24806
rect 7470 24783 7526 24792
rect 7484 24750 7512 24783
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 7208 24364 7328 24392
rect 7378 24440 7434 24449
rect 7378 24375 7434 24384
rect 7208 24274 7236 24364
rect 7288 24302 7340 24308
rect 7196 24268 7248 24274
rect 7392 24290 7420 24375
rect 7340 24262 7420 24290
rect 7470 24304 7526 24313
rect 7288 24244 7340 24250
rect 7470 24239 7472 24248
rect 7196 24210 7248 24216
rect 7524 24239 7526 24248
rect 7472 24210 7524 24216
rect 7288 24200 7340 24206
rect 7340 24160 7420 24188
rect 7288 24142 7340 24148
rect 7288 24064 7340 24070
rect 7392 24041 7420 24160
rect 7288 24006 7340 24012
rect 7378 24032 7434 24041
rect 7116 23820 7236 23848
rect 7104 23724 7156 23730
rect 7104 23666 7156 23672
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 6826 22944 6882 22953
rect 6826 22879 6882 22888
rect 6644 22772 6696 22778
rect 6748 22766 7052 22794
rect 7116 22778 7144 23666
rect 7208 23594 7236 23820
rect 7300 23662 7328 24006
rect 7378 23967 7434 23976
rect 7378 23896 7434 23905
rect 7378 23831 7434 23840
rect 7472 23860 7524 23866
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 7196 23588 7248 23594
rect 7196 23530 7248 23536
rect 6644 22714 6696 22720
rect 6734 22672 6790 22681
rect 6734 22607 6790 22616
rect 6552 22568 6604 22574
rect 6604 22516 6684 22522
rect 6552 22510 6684 22516
rect 6564 22494 6684 22510
rect 6748 22506 6776 22607
rect 6656 22438 6684 22494
rect 6736 22500 6788 22506
rect 6736 22442 6788 22448
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6734 22400 6790 22409
rect 6564 22001 6592 22374
rect 6734 22335 6790 22344
rect 6642 22264 6698 22273
rect 6642 22199 6644 22208
rect 6696 22199 6698 22208
rect 6644 22170 6696 22176
rect 6748 22098 6776 22335
rect 7024 22166 7052 22766
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7102 22672 7158 22681
rect 7102 22607 7158 22616
rect 7116 22438 7144 22607
rect 7208 22574 7236 23530
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7300 23089 7328 23122
rect 7286 23080 7342 23089
rect 7286 23015 7342 23024
rect 7288 22976 7340 22982
rect 7288 22918 7340 22924
rect 7196 22568 7248 22574
rect 7196 22510 7248 22516
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7102 22264 7158 22273
rect 7102 22199 7158 22208
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 7012 22160 7064 22166
rect 7012 22102 7064 22108
rect 6644 22092 6696 22098
rect 6644 22034 6696 22040
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6550 21992 6606 22001
rect 6550 21927 6606 21936
rect 6656 21706 6684 22034
rect 6932 21978 6960 22102
rect 6932 21950 7052 21978
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 6552 21684 6604 21690
rect 6656 21678 6776 21706
rect 6552 21626 6604 21632
rect 6564 20602 6592 21626
rect 6748 21554 6776 21678
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6826 21448 6882 21457
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6564 19990 6592 20402
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6368 18828 6420 18834
rect 6472 18816 6500 19246
rect 6552 18828 6604 18834
rect 6472 18788 6552 18816
rect 6368 18770 6420 18776
rect 6552 18770 6604 18776
rect 6380 18698 6408 18770
rect 6564 18698 6592 18770
rect 6368 18692 6420 18698
rect 6288 18652 6368 18680
rect 6288 17746 6316 18652
rect 6368 18634 6420 18640
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6564 18290 6592 18362
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6550 18184 6606 18193
rect 6368 18148 6420 18154
rect 6362 18096 6368 18136
rect 6550 18119 6552 18128
rect 6362 18090 6420 18096
rect 6604 18119 6606 18128
rect 6552 18090 6604 18096
rect 6362 18034 6390 18090
rect 6550 18048 6606 18057
rect 6362 18006 6408 18034
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6274 17640 6330 17649
rect 6274 17575 6276 17584
rect 6328 17575 6330 17584
rect 6276 17546 6328 17552
rect 6288 17377 6316 17546
rect 6274 17368 6330 17377
rect 6274 17303 6330 17312
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 6288 16522 6316 17002
rect 6380 16561 6408 18006
rect 6550 17983 6606 17992
rect 6564 17814 6592 17983
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6472 16794 6500 17682
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 6564 16674 6592 17614
rect 6656 17377 6684 21422
rect 6826 21383 6882 21392
rect 6736 21072 6788 21078
rect 6736 21014 6788 21020
rect 6748 20874 6776 21014
rect 6736 20868 6788 20874
rect 6736 20810 6788 20816
rect 6748 19904 6776 20810
rect 6840 20618 6868 21383
rect 6932 20942 6960 21830
rect 7024 21418 7052 21950
rect 7116 21622 7144 22199
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 7012 21140 7064 21146
rect 7116 21128 7144 21558
rect 7208 21486 7236 22374
rect 7300 21962 7328 22918
rect 7392 22794 7420 23831
rect 7576 23848 7604 25214
rect 7656 25152 7708 25158
rect 7760 25129 7788 25298
rect 7656 25094 7708 25100
rect 7746 25120 7802 25129
rect 7668 24750 7696 25094
rect 7746 25055 7802 25064
rect 7852 24868 7880 25316
rect 8036 25226 8064 25638
rect 7932 25220 7984 25226
rect 7932 25162 7984 25168
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 7760 24840 7880 24868
rect 7656 24744 7708 24750
rect 7656 24686 7708 24692
rect 7656 24608 7708 24614
rect 7656 24550 7708 24556
rect 7524 23820 7604 23848
rect 7472 23802 7524 23808
rect 7484 23254 7512 23802
rect 7668 23780 7696 24550
rect 7760 23905 7788 24840
rect 7944 24750 7972 25162
rect 8036 24857 8064 25162
rect 8022 24848 8078 24857
rect 8022 24783 8078 24792
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7932 24744 7984 24750
rect 8128 24698 8156 25792
rect 7932 24686 7984 24692
rect 7852 24206 7880 24686
rect 8036 24670 8156 24698
rect 8036 24562 8064 24670
rect 7944 24534 8064 24562
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7944 24120 7972 24534
rect 8128 24256 8156 24550
rect 7912 24092 7972 24120
rect 8036 24228 8156 24256
rect 7912 24018 7940 24092
rect 7852 23990 7940 24018
rect 7746 23896 7802 23905
rect 7852 23866 7880 23990
rect 7930 23896 7986 23905
rect 7746 23831 7802 23840
rect 7840 23860 7892 23866
rect 7930 23831 7986 23840
rect 7840 23802 7892 23808
rect 7576 23752 7696 23780
rect 7472 23248 7524 23254
rect 7472 23190 7524 23196
rect 7576 23118 7604 23752
rect 7748 23724 7800 23730
rect 7668 23684 7748 23712
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7392 22766 7512 22794
rect 7380 22704 7432 22710
rect 7380 22646 7432 22652
rect 7288 21956 7340 21962
rect 7288 21898 7340 21904
rect 7288 21616 7340 21622
rect 7288 21558 7340 21564
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7194 21312 7250 21321
rect 7194 21247 7250 21256
rect 7064 21100 7144 21128
rect 7012 21082 7064 21088
rect 7208 20942 7236 21247
rect 7300 21010 7328 21558
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 6920 20936 6972 20942
rect 7196 20936 7248 20942
rect 6972 20896 7052 20924
rect 6920 20878 6972 20884
rect 6840 20602 6960 20618
rect 6840 20596 6972 20602
rect 6840 20590 6920 20596
rect 6920 20538 6972 20544
rect 6826 20360 6882 20369
rect 6826 20295 6882 20304
rect 6840 20262 6868 20295
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 7024 19938 7052 20896
rect 7196 20878 7248 20884
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 7116 20466 7144 20742
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7286 20360 7342 20369
rect 7286 20295 7342 20304
rect 7300 20262 7328 20295
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 6828 19916 6880 19922
rect 6748 19876 6828 19904
rect 6828 19858 6880 19864
rect 6932 19910 7052 19938
rect 7104 19916 7156 19922
rect 6932 19854 6960 19910
rect 7104 19858 7156 19864
rect 7196 19916 7248 19922
rect 7196 19858 7248 19864
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6840 19310 6868 19722
rect 6932 19689 6960 19790
rect 6918 19680 6974 19689
rect 6918 19615 6974 19624
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6932 18970 6960 19246
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 6826 18864 6882 18873
rect 6826 18799 6882 18808
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 17882 6776 18566
rect 6840 18465 6868 18799
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6826 18456 6882 18465
rect 6826 18391 6882 18400
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6840 17762 6868 18294
rect 6932 18086 6960 18702
rect 7024 18170 7052 19790
rect 7116 19310 7144 19858
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7116 18630 7144 19246
rect 7208 18902 7236 19858
rect 7300 19718 7328 20198
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7300 19310 7328 19450
rect 7392 19446 7420 22646
rect 7484 22438 7512 22766
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7576 22001 7604 22918
rect 7668 22506 7696 23684
rect 7748 23666 7800 23672
rect 7838 23624 7894 23633
rect 7838 23559 7840 23568
rect 7892 23559 7894 23568
rect 7840 23530 7892 23536
rect 7944 23322 7972 23831
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 7656 22500 7708 22506
rect 7656 22442 7708 22448
rect 7562 21992 7618 22001
rect 7562 21927 7618 21936
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 7484 21010 7512 21626
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7576 20505 7604 21354
rect 7668 21350 7696 22442
rect 7760 22273 7788 23258
rect 7932 23180 7984 23186
rect 7932 23122 7984 23128
rect 7944 22710 7972 23122
rect 7932 22704 7984 22710
rect 7932 22646 7984 22652
rect 7840 22568 7892 22574
rect 7840 22510 7892 22516
rect 7932 22568 7984 22574
rect 7932 22510 7984 22516
rect 7746 22264 7802 22273
rect 7746 22199 7802 22208
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7760 21554 7788 22034
rect 7852 22030 7880 22510
rect 7944 22273 7972 22510
rect 7930 22264 7986 22273
rect 7930 22199 7932 22208
rect 7984 22199 7986 22208
rect 7932 22170 7984 22176
rect 8036 22114 8064 24228
rect 8116 24132 8168 24138
rect 8116 24074 8168 24080
rect 8128 23712 8156 24074
rect 8220 23866 8248 25894
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8128 23684 8248 23712
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 8128 22234 8156 23530
rect 8220 23361 8248 23684
rect 8206 23352 8262 23361
rect 8206 23287 8262 23296
rect 8208 23248 8260 23254
rect 8206 23216 8208 23225
rect 8260 23216 8262 23225
rect 8206 23151 8262 23160
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8220 22642 8248 23054
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 8036 22086 8156 22114
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7944 21622 7972 21830
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7668 20754 7696 21286
rect 7760 21146 7788 21490
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7852 21010 7880 21286
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 7838 20904 7894 20913
rect 7944 20890 7972 21422
rect 7894 20862 7972 20890
rect 8024 20936 8076 20942
rect 8024 20878 8076 20884
rect 7838 20839 7894 20848
rect 7668 20726 7788 20754
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7562 20496 7618 20505
rect 7562 20431 7618 20440
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7484 19854 7512 20198
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7380 19440 7432 19446
rect 7380 19382 7432 19388
rect 7288 19304 7340 19310
rect 7340 19264 7420 19292
rect 7288 19246 7340 19252
rect 7196 18896 7248 18902
rect 7196 18838 7248 18844
rect 7288 18896 7340 18902
rect 7288 18838 7340 18844
rect 7300 18698 7328 18838
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7104 18624 7156 18630
rect 7300 18601 7328 18634
rect 7104 18566 7156 18572
rect 7286 18592 7342 18601
rect 7286 18527 7342 18536
rect 7286 18456 7342 18465
rect 7286 18391 7342 18400
rect 7300 18222 7328 18391
rect 7288 18216 7340 18222
rect 7208 18176 7288 18204
rect 7024 18142 7144 18170
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6748 17734 6868 17762
rect 6642 17368 6698 17377
rect 6642 17303 6698 17312
rect 6472 16646 6592 16674
rect 6748 16658 6776 17734
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 17542 6868 17614
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6840 17338 6868 17478
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6826 17232 6882 17241
rect 6826 17167 6828 17176
rect 6880 17167 6882 17176
rect 6828 17138 6880 17144
rect 6826 16824 6882 16833
rect 6826 16759 6828 16768
rect 6880 16759 6882 16768
rect 6828 16730 6880 16736
rect 6826 16688 6882 16697
rect 6736 16652 6788 16658
rect 6366 16552 6422 16561
rect 6276 16516 6328 16522
rect 6366 16487 6422 16496
rect 6276 16458 6328 16464
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6288 15570 6316 15914
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6090 15056 6146 15065
rect 6090 14991 6146 15000
rect 6184 15020 6236 15026
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5828 14278 5856 14418
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5356 12436 5408 12442
rect 5644 12434 5672 13806
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5356 12378 5408 12384
rect 5460 12406 5672 12434
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4764 11172 4844 11200
rect 4712 11154 4764 11160
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9178 4200 9998
rect 4264 9654 4292 11154
rect 4356 10742 4384 11154
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 4724 9994 4752 10474
rect 4802 10160 4858 10169
rect 5000 10146 5028 12106
rect 5368 11370 5396 12242
rect 5184 11342 5396 11370
rect 4802 10095 4858 10104
rect 4896 10124 4948 10130
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 4724 9178 4752 9454
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4172 8634 4200 8978
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3344 6718 3464 6746
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3160 4826 3188 5102
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2976 4214 3004 4490
rect 3344 4282 3372 6718
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6254 3464 6598
rect 3528 6458 3556 7142
rect 3896 7002 3924 7278
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3896 6662 3924 6938
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3792 6384 3844 6390
rect 3790 6352 3792 6361
rect 3844 6352 3846 6361
rect 3790 6287 3846 6296
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 4080 5302 4108 6802
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3528 4826 3556 5170
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3528 3738 3556 4082
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2884 2650 2912 2790
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2608 1766 2636 2450
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2596 1760 2648 1766
rect 2596 1702 2648 1708
rect 2320 1556 2372 1562
rect 2320 1498 2372 1504
rect 2332 1426 2360 1498
rect 2044 1420 2096 1426
rect 2044 1362 2096 1368
rect 2320 1420 2372 1426
rect 2320 1362 2372 1368
rect 1952 1352 2004 1358
rect 1952 1294 2004 1300
rect 2792 814 2820 2314
rect 2976 1902 3004 2858
rect 2964 1896 3016 1902
rect 2964 1838 3016 1844
rect 3068 1578 3096 2926
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3160 1834 3188 2790
rect 3516 2576 3568 2582
rect 3516 2518 3568 2524
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3148 1828 3200 1834
rect 3148 1770 3200 1776
rect 3252 1766 3280 2450
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3344 1970 3372 2382
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 3240 1760 3292 1766
rect 3240 1702 3292 1708
rect 2976 1562 3096 1578
rect 2964 1556 3096 1562
rect 3016 1550 3096 1556
rect 2964 1498 3016 1504
rect 3344 1494 3372 1906
rect 3056 1488 3108 1494
rect 3056 1430 3108 1436
rect 3332 1488 3384 1494
rect 3332 1430 3384 1436
rect 2780 808 2832 814
rect 2780 750 2832 756
rect 3068 746 3096 1430
rect 3240 1420 3292 1426
rect 3240 1362 3292 1368
rect 3252 1018 3280 1362
rect 3436 1018 3464 2246
rect 3528 2106 3556 2518
rect 3620 2378 3648 3130
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 4172 2310 4200 8298
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4264 6322 4292 7278
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4632 6338 4660 6598
rect 4724 6458 4752 6802
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4252 6316 4304 6322
rect 4632 6310 4752 6338
rect 4252 6258 4304 6264
rect 4264 4690 4292 6258
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 4724 5522 4752 6310
rect 4816 5760 4844 10095
rect 5000 10118 5120 10146
rect 4896 10066 4948 10072
rect 4908 9722 4936 10066
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5000 9518 5028 9998
rect 5092 9654 5120 10118
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5092 9178 5120 9454
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5092 7342 5120 8978
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6866 5028 7142
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 5000 6254 5028 6802
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5092 6186 5120 7278
rect 5184 6730 5212 11342
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5276 10266 5304 11154
rect 5460 10810 5488 12406
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5460 10606 5488 10746
rect 5448 10600 5500 10606
rect 5368 10560 5448 10588
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5368 9738 5396 10560
rect 5448 10542 5500 10548
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5460 10130 5488 10406
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5368 9710 5488 9738
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5276 6458 5304 6802
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5092 5846 5120 6122
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 4816 5732 4936 5760
rect 4724 5494 4844 5522
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4540 4282 4568 4694
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4264 3602 4292 4150
rect 4540 4078 4568 4218
rect 4724 4078 4752 4626
rect 4816 4570 4844 5494
rect 4908 4758 4936 5732
rect 5368 5642 5396 9590
rect 5460 9518 5488 9710
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5552 7478 5580 12310
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5644 11082 5672 11630
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5736 10742 5764 12650
rect 5920 11898 5948 14894
rect 6104 14890 6132 14991
rect 6184 14962 6236 14968
rect 6092 14884 6144 14890
rect 6012 14844 6092 14872
rect 6012 14346 6040 14844
rect 6092 14826 6144 14832
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 6012 12782 6040 14282
rect 6196 13870 6224 14962
rect 6288 14958 6316 15506
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6288 14074 6316 14350
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6104 12782 6132 13738
rect 6196 12782 6224 13806
rect 6380 13546 6408 16186
rect 6472 14958 6500 16646
rect 6826 16623 6828 16632
rect 6736 16594 6788 16600
rect 6880 16623 6882 16632
rect 6828 16594 6880 16600
rect 6552 16584 6604 16590
rect 6550 16552 6552 16561
rect 6604 16552 6606 16561
rect 6550 16487 6606 16496
rect 6642 16416 6698 16425
rect 6642 16351 6698 16360
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6564 15337 6592 15506
rect 6550 15328 6606 15337
rect 6550 15263 6606 15272
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6472 13734 6500 14894
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6380 13518 6500 13546
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6380 12889 6408 13330
rect 6366 12880 6422 12889
rect 6366 12815 6422 12824
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5828 11218 5856 11290
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5632 10600 5684 10606
rect 5630 10568 5632 10577
rect 5684 10568 5686 10577
rect 5630 10503 5686 10512
rect 5736 9586 5764 10678
rect 5920 9994 5948 11154
rect 6012 10282 6040 12718
rect 6380 12306 6408 12815
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6472 12238 6500 13518
rect 6564 13394 6592 15263
rect 6656 14929 6684 16351
rect 6840 16250 6868 16594
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6642 14920 6698 14929
rect 6642 14855 6698 14864
rect 6656 14550 6684 14855
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6196 11694 6224 12038
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 11354 6224 11494
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6288 10538 6316 10746
rect 6472 10742 6500 11154
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6564 10588 6592 13330
rect 6656 12288 6684 14350
rect 6748 12442 6776 15506
rect 6840 13326 6868 15642
rect 6932 14890 6960 18022
rect 7024 16726 7052 18022
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7116 15706 7144 18142
rect 7208 17921 7236 18176
rect 7288 18158 7340 18164
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7194 17912 7250 17921
rect 7194 17847 7250 17856
rect 7196 17740 7248 17746
rect 7300 17728 7328 18022
rect 7392 17921 7420 19264
rect 7484 18329 7512 19654
rect 7576 18834 7604 20431
rect 7668 19417 7696 20538
rect 7760 20097 7788 20726
rect 7746 20088 7802 20097
rect 7746 20023 7802 20032
rect 7760 19854 7788 20023
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7654 19408 7710 19417
rect 7654 19343 7710 19352
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7760 18834 7788 19314
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7576 18358 7604 18770
rect 7564 18352 7616 18358
rect 7470 18320 7526 18329
rect 7656 18352 7708 18358
rect 7564 18294 7616 18300
rect 7654 18320 7656 18329
rect 7708 18320 7710 18329
rect 7470 18255 7526 18264
rect 7654 18255 7710 18264
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7656 18216 7708 18222
rect 7470 18184 7526 18193
rect 7656 18158 7708 18164
rect 7470 18119 7526 18128
rect 7378 17912 7434 17921
rect 7378 17847 7434 17856
rect 7380 17808 7432 17814
rect 7484 17796 7512 18119
rect 7562 17912 7618 17921
rect 7562 17847 7618 17856
rect 7668 17864 7696 18158
rect 7760 18057 7788 18226
rect 7746 18048 7802 18057
rect 7746 17983 7802 17992
rect 7748 17876 7800 17882
rect 7432 17768 7512 17796
rect 7380 17750 7432 17756
rect 7248 17700 7328 17728
rect 7576 17728 7604 17847
rect 7668 17836 7748 17864
rect 7748 17818 7800 17824
rect 7656 17740 7708 17746
rect 7576 17700 7656 17728
rect 7196 17682 7248 17688
rect 7656 17682 7708 17688
rect 7208 17202 7236 17682
rect 7470 17640 7526 17649
rect 7288 17604 7340 17610
rect 7470 17575 7526 17584
rect 7288 17546 7340 17552
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7300 16794 7328 17546
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7392 15722 7420 17070
rect 7484 16726 7512 17575
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7576 17377 7604 17478
rect 7562 17368 7618 17377
rect 7668 17338 7696 17682
rect 7562 17303 7618 17312
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7760 17134 7788 17818
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7576 16250 7604 17070
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7760 16726 7788 16934
rect 7852 16794 7880 20839
rect 8036 20330 8064 20878
rect 8024 20324 8076 20330
rect 8024 20266 8076 20272
rect 7932 19984 7984 19990
rect 7930 19952 7932 19961
rect 7984 19952 7986 19961
rect 7986 19910 8064 19938
rect 7930 19887 7986 19896
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7944 19514 7972 19654
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 8036 19394 8064 19910
rect 7944 19366 8064 19394
rect 7944 19174 7972 19366
rect 8128 19310 8156 22086
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8220 21593 8248 21966
rect 8206 21584 8262 21593
rect 8206 21519 8262 21528
rect 8312 20754 8340 25978
rect 8404 25906 8432 28562
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8496 25838 8524 30058
rect 8588 29850 8616 31146
rect 8680 30258 8708 31622
rect 8668 30252 8720 30258
rect 8668 30194 8720 30200
rect 8576 29844 8628 29850
rect 8576 29786 8628 29792
rect 8668 29708 8720 29714
rect 8668 29650 8720 29656
rect 8576 29572 8628 29578
rect 8576 29514 8628 29520
rect 8588 29238 8616 29514
rect 8576 29232 8628 29238
rect 8576 29174 8628 29180
rect 8576 29096 8628 29102
rect 8574 29064 8576 29073
rect 8628 29064 8630 29073
rect 8574 28999 8630 29008
rect 8576 28620 8628 28626
rect 8576 28562 8628 28568
rect 8588 27577 8616 28562
rect 8574 27568 8630 27577
rect 8574 27503 8630 27512
rect 8576 27464 8628 27470
rect 8576 27406 8628 27412
rect 8588 27033 8616 27406
rect 8574 27024 8630 27033
rect 8574 26959 8630 26968
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8588 26761 8616 26862
rect 8574 26752 8630 26761
rect 8574 26687 8630 26696
rect 8680 26518 8708 29650
rect 8772 29102 8800 31719
rect 8852 31136 8904 31142
rect 8852 31078 8904 31084
rect 8864 30569 8892 31078
rect 8956 30938 8984 31894
rect 9140 31890 9168 32014
rect 9232 32008 9260 33215
rect 9324 32473 9352 33322
rect 9416 33017 9444 34138
rect 9402 33008 9458 33017
rect 9402 32943 9458 32952
rect 9310 32464 9366 32473
rect 9310 32399 9366 32408
rect 9324 32366 9352 32399
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 9312 32020 9364 32026
rect 9232 31980 9312 32008
rect 9312 31962 9364 31968
rect 9036 31884 9088 31890
rect 9036 31826 9088 31832
rect 9128 31884 9180 31890
rect 9128 31826 9180 31832
rect 8944 30932 8996 30938
rect 8944 30874 8996 30880
rect 8944 30592 8996 30598
rect 8850 30560 8906 30569
rect 8944 30534 8996 30540
rect 8850 30495 8906 30504
rect 8852 30252 8904 30258
rect 8852 30194 8904 30200
rect 8760 29096 8812 29102
rect 8760 29038 8812 29044
rect 8760 28484 8812 28490
rect 8760 28426 8812 28432
rect 8772 27402 8800 28426
rect 8760 27396 8812 27402
rect 8760 27338 8812 27344
rect 8864 27010 8892 30194
rect 8956 29646 8984 30534
rect 8944 29640 8996 29646
rect 8944 29582 8996 29588
rect 8956 28626 8984 29582
rect 8944 28620 8996 28626
rect 8944 28562 8996 28568
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 8956 27674 8984 28018
rect 8944 27668 8996 27674
rect 8944 27610 8996 27616
rect 8942 27568 8998 27577
rect 8942 27503 8998 27512
rect 8956 27402 8984 27503
rect 8944 27396 8996 27402
rect 8944 27338 8996 27344
rect 8956 27305 8984 27338
rect 8942 27296 8998 27305
rect 8942 27231 8998 27240
rect 8772 26982 8892 27010
rect 8944 26988 8996 26994
rect 8668 26512 8720 26518
rect 8668 26454 8720 26460
rect 8576 26308 8628 26314
rect 8576 26250 8628 26256
rect 8484 25832 8536 25838
rect 8482 25800 8484 25809
rect 8536 25800 8538 25809
rect 8482 25735 8538 25744
rect 8588 25537 8616 26250
rect 8772 25673 8800 26982
rect 8944 26930 8996 26936
rect 8852 26920 8904 26926
rect 8852 26862 8904 26868
rect 8758 25664 8814 25673
rect 8758 25599 8814 25608
rect 8574 25528 8630 25537
rect 8484 25492 8536 25498
rect 8574 25463 8576 25472
rect 8484 25434 8536 25440
rect 8628 25463 8630 25472
rect 8576 25434 8628 25440
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 8404 24818 8432 25298
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8496 24682 8524 25434
rect 8574 25392 8630 25401
rect 8574 25327 8576 25336
rect 8628 25327 8630 25336
rect 8576 25298 8628 25304
rect 8588 24886 8616 25298
rect 8772 25294 8800 25599
rect 8864 25498 8892 26862
rect 8852 25492 8904 25498
rect 8852 25434 8904 25440
rect 8760 25288 8812 25294
rect 8760 25230 8812 25236
rect 8666 25120 8722 25129
rect 8666 25055 8722 25064
rect 8576 24880 8628 24886
rect 8576 24822 8628 24828
rect 8574 24712 8630 24721
rect 8392 24676 8444 24682
rect 8392 24618 8444 24624
rect 8484 24676 8536 24682
rect 8680 24682 8708 25055
rect 8852 24880 8904 24886
rect 8852 24822 8904 24828
rect 8574 24647 8630 24656
rect 8668 24676 8720 24682
rect 8484 24618 8536 24624
rect 8404 24070 8432 24618
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8390 23896 8446 23905
rect 8390 23831 8392 23840
rect 8444 23831 8446 23840
rect 8392 23802 8444 23808
rect 8390 23624 8446 23633
rect 8390 23559 8446 23568
rect 8404 22166 8432 23559
rect 8496 23186 8524 24618
rect 8588 24410 8616 24647
rect 8668 24618 8720 24624
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8574 24304 8630 24313
rect 8680 24290 8708 24618
rect 8864 24313 8892 24822
rect 8956 24342 8984 26930
rect 9048 26926 9076 31826
rect 9128 31748 9180 31754
rect 9128 31690 9180 31696
rect 9140 31657 9168 31690
rect 9126 31648 9182 31657
rect 9126 31583 9182 31592
rect 9324 31362 9352 31962
rect 9416 31482 9444 32943
rect 9508 32434 9536 35430
rect 9600 34202 9628 35430
rect 9588 34196 9640 34202
rect 9588 34138 9640 34144
rect 9588 33448 9640 33454
rect 9588 33390 9640 33396
rect 9600 32502 9628 33390
rect 9692 33114 9720 35566
rect 9784 35550 9904 35578
rect 9772 35488 9824 35494
rect 9772 35430 9824 35436
rect 9784 35222 9812 35430
rect 9772 35216 9824 35222
rect 9772 35158 9824 35164
rect 9772 34060 9824 34066
rect 9772 34002 9824 34008
rect 9784 33522 9812 34002
rect 9876 33697 9904 35550
rect 9968 35193 9996 36094
rect 10598 36071 10654 36080
rect 10062 35932 10370 35941
rect 10062 35930 10068 35932
rect 10124 35930 10148 35932
rect 10204 35930 10228 35932
rect 10284 35930 10308 35932
rect 10364 35930 10370 35932
rect 10124 35878 10126 35930
rect 10306 35878 10308 35930
rect 10062 35876 10068 35878
rect 10124 35876 10148 35878
rect 10204 35876 10228 35878
rect 10284 35876 10308 35878
rect 10364 35876 10370 35878
rect 10062 35867 10370 35876
rect 10416 35488 10468 35494
rect 10416 35430 10468 35436
rect 9954 35184 10010 35193
rect 9954 35119 10010 35128
rect 10428 34950 10456 35430
rect 10722 35388 11030 35397
rect 10722 35386 10728 35388
rect 10784 35386 10808 35388
rect 10864 35386 10888 35388
rect 10944 35386 10968 35388
rect 11024 35386 11030 35388
rect 10784 35334 10786 35386
rect 10966 35334 10968 35386
rect 10722 35332 10728 35334
rect 10784 35332 10808 35334
rect 10864 35332 10888 35334
rect 10944 35332 10968 35334
rect 11024 35332 11030 35334
rect 10722 35323 11030 35332
rect 10598 35048 10654 35057
rect 10598 34983 10654 34992
rect 10416 34944 10468 34950
rect 10416 34886 10468 34892
rect 10508 34944 10560 34950
rect 10508 34886 10560 34892
rect 10062 34844 10370 34853
rect 10062 34842 10068 34844
rect 10124 34842 10148 34844
rect 10204 34842 10228 34844
rect 10284 34842 10308 34844
rect 10364 34842 10370 34844
rect 10124 34790 10126 34842
rect 10306 34790 10308 34842
rect 10062 34788 10068 34790
rect 10124 34788 10148 34790
rect 10204 34788 10228 34790
rect 10284 34788 10308 34790
rect 10364 34788 10370 34790
rect 10062 34779 10370 34788
rect 9956 34672 10008 34678
rect 9956 34614 10008 34620
rect 9862 33688 9918 33697
rect 9862 33623 9918 33632
rect 9864 33584 9916 33590
rect 9864 33526 9916 33532
rect 9772 33516 9824 33522
rect 9772 33458 9824 33464
rect 9772 33312 9824 33318
rect 9772 33254 9824 33260
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 9680 32972 9732 32978
rect 9680 32914 9732 32920
rect 9588 32496 9640 32502
rect 9588 32438 9640 32444
rect 9496 32428 9548 32434
rect 9496 32370 9548 32376
rect 9588 32360 9640 32366
rect 9494 32328 9550 32337
rect 9588 32302 9640 32308
rect 9494 32263 9550 32272
rect 9508 31958 9536 32263
rect 9496 31952 9548 31958
rect 9496 31894 9548 31900
rect 9508 31822 9536 31894
rect 9496 31816 9548 31822
rect 9496 31758 9548 31764
rect 9404 31476 9456 31482
rect 9404 31418 9456 31424
rect 9324 31334 9536 31362
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 9128 30184 9180 30190
rect 9128 30126 9180 30132
rect 9140 29306 9168 30126
rect 9220 30116 9272 30122
rect 9220 30058 9272 30064
rect 9128 29300 9180 29306
rect 9128 29242 9180 29248
rect 9140 29073 9168 29242
rect 9126 29064 9182 29073
rect 9232 29034 9260 30058
rect 9312 29844 9364 29850
rect 9312 29786 9364 29792
rect 9126 28999 9182 29008
rect 9220 29028 9272 29034
rect 9220 28970 9272 28976
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 9140 28762 9168 28902
rect 9128 28756 9180 28762
rect 9128 28698 9180 28704
rect 9128 28620 9180 28626
rect 9232 28608 9260 28970
rect 9180 28580 9260 28608
rect 9128 28562 9180 28568
rect 9324 28558 9352 29786
rect 9416 29782 9444 30534
rect 9404 29776 9456 29782
rect 9404 29718 9456 29724
rect 9416 29510 9444 29718
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9508 28994 9536 31334
rect 9600 30394 9628 32302
rect 9692 31754 9720 32914
rect 9784 32298 9812 33254
rect 9772 32292 9824 32298
rect 9772 32234 9824 32240
rect 9692 31726 9812 31754
rect 9680 31680 9732 31686
rect 9680 31622 9732 31628
rect 9692 30870 9720 31622
rect 9680 30864 9732 30870
rect 9680 30806 9732 30812
rect 9784 30734 9812 31726
rect 9876 31278 9904 33526
rect 9968 33046 9996 34614
rect 10428 34610 10456 34886
rect 10416 34604 10468 34610
rect 10416 34546 10468 34552
rect 10140 34536 10192 34542
rect 10140 34478 10192 34484
rect 10324 34536 10376 34542
rect 10520 34490 10548 34886
rect 10612 34542 10640 34983
rect 11072 34762 11100 37266
rect 10980 34734 11100 34762
rect 10980 34542 11008 34734
rect 11060 34672 11112 34678
rect 11060 34614 11112 34620
rect 10324 34478 10376 34484
rect 10152 33930 10180 34478
rect 10232 34400 10284 34406
rect 10232 34342 10284 34348
rect 10140 33924 10192 33930
rect 10140 33866 10192 33872
rect 10244 33862 10272 34342
rect 10336 34066 10364 34478
rect 10428 34474 10548 34490
rect 10600 34536 10652 34542
rect 10968 34536 11020 34542
rect 10600 34478 10652 34484
rect 10966 34504 10968 34513
rect 11020 34504 11022 34513
rect 10416 34468 10548 34474
rect 10468 34462 10548 34468
rect 10416 34410 10468 34416
rect 10324 34060 10376 34066
rect 10324 34002 10376 34008
rect 10232 33856 10284 33862
rect 10232 33798 10284 33804
rect 10416 33856 10468 33862
rect 10416 33798 10468 33804
rect 10062 33756 10370 33765
rect 10062 33754 10068 33756
rect 10124 33754 10148 33756
rect 10204 33754 10228 33756
rect 10284 33754 10308 33756
rect 10364 33754 10370 33756
rect 10124 33702 10126 33754
rect 10306 33702 10308 33754
rect 10062 33700 10068 33702
rect 10124 33700 10148 33702
rect 10204 33700 10228 33702
rect 10284 33700 10308 33702
rect 10364 33700 10370 33702
rect 10062 33691 10370 33700
rect 10428 33590 10456 33798
rect 10416 33584 10468 33590
rect 10416 33526 10468 33532
rect 10140 33448 10192 33454
rect 10416 33448 10468 33454
rect 10140 33390 10192 33396
rect 10414 33416 10416 33425
rect 10468 33416 10470 33425
rect 9956 33040 10008 33046
rect 9956 32982 10008 32988
rect 10152 32756 10180 33390
rect 10414 33351 10470 33360
rect 10416 33312 10468 33318
rect 10416 33254 10468 33260
rect 9968 32728 10180 32756
rect 9968 31958 9996 32728
rect 10062 32668 10370 32677
rect 10062 32666 10068 32668
rect 10124 32666 10148 32668
rect 10204 32666 10228 32668
rect 10284 32666 10308 32668
rect 10364 32666 10370 32668
rect 10124 32614 10126 32666
rect 10306 32614 10308 32666
rect 10062 32612 10068 32614
rect 10124 32612 10148 32614
rect 10204 32612 10228 32614
rect 10284 32612 10308 32614
rect 10364 32612 10370 32614
rect 10062 32603 10370 32612
rect 10428 32026 10456 33254
rect 10520 32910 10548 34462
rect 10966 34439 11022 34448
rect 10600 34400 10652 34406
rect 10600 34342 10652 34348
rect 10612 34202 10640 34342
rect 10722 34300 11030 34309
rect 10722 34298 10728 34300
rect 10784 34298 10808 34300
rect 10864 34298 10888 34300
rect 10944 34298 10968 34300
rect 11024 34298 11030 34300
rect 10784 34246 10786 34298
rect 10966 34246 10968 34298
rect 10722 34244 10728 34246
rect 10784 34244 10808 34246
rect 10864 34244 10888 34246
rect 10944 34244 10968 34246
rect 11024 34244 11030 34246
rect 10722 34235 11030 34244
rect 10600 34196 10652 34202
rect 10600 34138 10652 34144
rect 10692 33924 10744 33930
rect 10692 33866 10744 33872
rect 10704 33658 10732 33866
rect 10692 33652 10744 33658
rect 10692 33594 10744 33600
rect 10722 33212 11030 33221
rect 10722 33210 10728 33212
rect 10784 33210 10808 33212
rect 10864 33210 10888 33212
rect 10944 33210 10968 33212
rect 11024 33210 11030 33212
rect 10784 33158 10786 33210
rect 10966 33158 10968 33210
rect 10722 33156 10728 33158
rect 10784 33156 10808 33158
rect 10864 33156 10888 33158
rect 10944 33156 10968 33158
rect 11024 33156 11030 33158
rect 10722 33147 11030 33156
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 10508 32904 10560 32910
rect 10508 32846 10560 32852
rect 10508 32564 10560 32570
rect 10508 32506 10560 32512
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10416 32020 10468 32026
rect 10416 31962 10468 31968
rect 9956 31952 10008 31958
rect 9956 31894 10008 31900
rect 10152 31822 10180 31962
rect 10520 31890 10548 32506
rect 10508 31884 10560 31890
rect 10508 31826 10560 31832
rect 9956 31816 10008 31822
rect 10048 31816 10100 31822
rect 9956 31758 10008 31764
rect 10046 31784 10048 31793
rect 10140 31816 10192 31822
rect 10100 31784 10102 31793
rect 9864 31272 9916 31278
rect 9864 31214 9916 31220
rect 9968 31142 9996 31758
rect 10140 31758 10192 31764
rect 10046 31719 10102 31728
rect 10062 31580 10370 31589
rect 10062 31578 10068 31580
rect 10124 31578 10148 31580
rect 10204 31578 10228 31580
rect 10284 31578 10308 31580
rect 10364 31578 10370 31580
rect 10124 31526 10126 31578
rect 10306 31526 10308 31578
rect 10062 31524 10068 31526
rect 10124 31524 10148 31526
rect 10204 31524 10228 31526
rect 10284 31524 10308 31526
rect 10364 31524 10370 31526
rect 10062 31515 10370 31524
rect 10508 31272 10560 31278
rect 10508 31214 10560 31220
rect 9956 31136 10008 31142
rect 9956 31078 10008 31084
rect 9772 30728 9824 30734
rect 9968 30705 9996 31078
rect 9772 30670 9824 30676
rect 9954 30696 10010 30705
rect 9954 30631 10010 30640
rect 10520 30598 10548 31214
rect 10612 31210 10640 33050
rect 10784 32836 10836 32842
rect 10784 32778 10836 32784
rect 10796 32434 10824 32778
rect 10888 32570 10916 33050
rect 10876 32564 10928 32570
rect 10876 32506 10928 32512
rect 10784 32428 10836 32434
rect 10784 32370 10836 32376
rect 10722 32124 11030 32133
rect 10722 32122 10728 32124
rect 10784 32122 10808 32124
rect 10864 32122 10888 32124
rect 10944 32122 10968 32124
rect 11024 32122 11030 32124
rect 10784 32070 10786 32122
rect 10966 32070 10968 32122
rect 10722 32068 10728 32070
rect 10784 32068 10808 32070
rect 10864 32068 10888 32070
rect 10944 32068 10968 32070
rect 11024 32068 11030 32070
rect 10722 32059 11030 32068
rect 10600 31204 10652 31210
rect 10600 31146 10652 31152
rect 10722 31036 11030 31045
rect 10722 31034 10728 31036
rect 10784 31034 10808 31036
rect 10864 31034 10888 31036
rect 10944 31034 10968 31036
rect 11024 31034 11030 31036
rect 10784 30982 10786 31034
rect 10966 30982 10968 31034
rect 10722 30980 10728 30982
rect 10784 30980 10808 30982
rect 10864 30980 10888 30982
rect 10944 30980 10968 30982
rect 11024 30980 11030 30982
rect 10722 30971 11030 30980
rect 10508 30592 10560 30598
rect 10508 30534 10560 30540
rect 10062 30492 10370 30501
rect 10062 30490 10068 30492
rect 10124 30490 10148 30492
rect 10204 30490 10228 30492
rect 10284 30490 10308 30492
rect 10364 30490 10370 30492
rect 10124 30438 10126 30490
rect 10306 30438 10308 30490
rect 10062 30436 10068 30438
rect 10124 30436 10148 30438
rect 10204 30436 10228 30438
rect 10284 30436 10308 30438
rect 10364 30436 10370 30438
rect 10062 30427 10370 30436
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9770 30288 9826 30297
rect 9770 30223 9826 30232
rect 9588 29504 9640 29510
rect 9588 29446 9640 29452
rect 9680 29504 9732 29510
rect 9680 29446 9732 29452
rect 9600 29306 9628 29446
rect 9588 29300 9640 29306
rect 9588 29242 9640 29248
rect 9508 28966 9628 28994
rect 9494 28792 9550 28801
rect 9494 28727 9550 28736
rect 9508 28694 9536 28727
rect 9404 28688 9456 28694
rect 9402 28656 9404 28665
rect 9496 28688 9548 28694
rect 9456 28656 9458 28665
rect 9496 28630 9548 28636
rect 9402 28591 9458 28600
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 9128 28008 9180 28014
rect 9126 27976 9128 27985
rect 9180 27976 9182 27985
rect 9324 27946 9352 28358
rect 9416 28082 9444 28494
rect 9496 28416 9548 28422
rect 9494 28384 9496 28393
rect 9548 28384 9550 28393
rect 9494 28319 9550 28328
rect 9508 28218 9536 28319
rect 9496 28212 9548 28218
rect 9496 28154 9548 28160
rect 9404 28076 9456 28082
rect 9404 28018 9456 28024
rect 9496 28076 9548 28082
rect 9496 28018 9548 28024
rect 9126 27911 9182 27920
rect 9312 27940 9364 27946
rect 9312 27882 9364 27888
rect 9220 27872 9272 27878
rect 9220 27814 9272 27820
rect 9128 27532 9180 27538
rect 9128 27474 9180 27480
rect 9140 27441 9168 27474
rect 9126 27432 9182 27441
rect 9126 27367 9182 27376
rect 9036 26920 9088 26926
rect 9128 26920 9180 26926
rect 9036 26862 9088 26868
rect 9126 26888 9128 26897
rect 9180 26888 9182 26897
rect 9048 26586 9076 26862
rect 9126 26823 9182 26832
rect 9128 26784 9180 26790
rect 9128 26726 9180 26732
rect 9036 26580 9088 26586
rect 9036 26522 9088 26528
rect 9036 26444 9088 26450
rect 9036 26386 9088 26392
rect 9048 25974 9076 26386
rect 9036 25968 9088 25974
rect 9036 25910 9088 25916
rect 9036 25696 9088 25702
rect 9036 25638 9088 25644
rect 9048 24342 9076 25638
rect 9140 25362 9168 26726
rect 9232 26314 9260 27814
rect 9324 26994 9352 27882
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 9324 26586 9352 26930
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 9312 26444 9364 26450
rect 9312 26386 9364 26392
rect 9324 26353 9352 26386
rect 9310 26344 9366 26353
rect 9220 26308 9272 26314
rect 9310 26279 9366 26288
rect 9220 26250 9272 26256
rect 9128 25356 9180 25362
rect 9128 25298 9180 25304
rect 9128 25220 9180 25226
rect 9128 25162 9180 25168
rect 9140 24993 9168 25162
rect 9126 24984 9182 24993
rect 9126 24919 9182 24928
rect 9232 24682 9260 26250
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9220 24676 9272 24682
rect 9220 24618 9272 24624
rect 9232 24449 9260 24618
rect 9324 24614 9352 26182
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9218 24440 9274 24449
rect 9218 24375 9274 24384
rect 8944 24336 8996 24342
rect 8630 24262 8708 24290
rect 8850 24304 8906 24313
rect 8760 24268 8812 24274
rect 8574 24239 8630 24248
rect 8588 23526 8616 24239
rect 8944 24278 8996 24284
rect 9036 24336 9088 24342
rect 9036 24278 9088 24284
rect 8850 24239 8906 24248
rect 8760 24210 8812 24216
rect 8666 24032 8722 24041
rect 8666 23967 8722 23976
rect 8680 23798 8708 23967
rect 8772 23798 8800 24210
rect 8864 24138 8892 24239
rect 8852 24132 8904 24138
rect 8852 24074 8904 24080
rect 8956 24041 8984 24278
rect 9128 24268 9180 24274
rect 9128 24210 9180 24216
rect 9036 24132 9088 24138
rect 9036 24074 9088 24080
rect 8942 24032 8998 24041
rect 8942 23967 8998 23976
rect 9048 23882 9076 24074
rect 8864 23854 9076 23882
rect 8668 23792 8720 23798
rect 8668 23734 8720 23740
rect 8760 23792 8812 23798
rect 8760 23734 8812 23740
rect 8666 23624 8722 23633
rect 8666 23559 8722 23568
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8484 23180 8536 23186
rect 8484 23122 8536 23128
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 8484 22976 8536 22982
rect 8484 22918 8536 22924
rect 8496 22642 8524 22918
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8588 22574 8616 23122
rect 8576 22568 8628 22574
rect 8574 22536 8576 22545
rect 8628 22536 8630 22545
rect 8574 22471 8630 22480
rect 8484 22432 8536 22438
rect 8484 22374 8536 22380
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 8390 21992 8446 22001
rect 8390 21927 8446 21936
rect 8404 21486 8432 21927
rect 8496 21486 8524 22374
rect 8680 22250 8708 23559
rect 8760 23180 8812 23186
rect 8760 23122 8812 23128
rect 8772 22778 8800 23122
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8588 22222 8708 22250
rect 8758 22264 8814 22273
rect 8588 22166 8616 22222
rect 8758 22199 8814 22208
rect 8576 22160 8628 22166
rect 8576 22102 8628 22108
rect 8772 22030 8800 22199
rect 8864 22166 8892 23854
rect 8944 23792 8996 23798
rect 9036 23792 9088 23798
rect 8944 23734 8996 23740
rect 9034 23760 9036 23769
rect 9088 23760 9090 23769
rect 8956 23662 8984 23734
rect 9034 23695 9090 23704
rect 8944 23656 8996 23662
rect 8944 23598 8996 23604
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 8956 22438 8984 23462
rect 9048 23322 9076 23598
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9034 23216 9090 23225
rect 9034 23151 9036 23160
rect 9088 23151 9090 23160
rect 9036 23122 9088 23128
rect 9140 22658 9168 24210
rect 9324 24206 9352 24550
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9220 24064 9272 24070
rect 9218 24032 9220 24041
rect 9272 24032 9274 24041
rect 9218 23967 9274 23976
rect 9218 23896 9274 23905
rect 9218 23831 9274 23840
rect 9232 23798 9260 23831
rect 9220 23792 9272 23798
rect 9220 23734 9272 23740
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9232 23322 9260 23598
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9048 22630 9168 22658
rect 9232 22642 9260 23258
rect 9324 23100 9352 24142
rect 9416 24041 9444 28018
rect 9508 27946 9536 28018
rect 9496 27940 9548 27946
rect 9496 27882 9548 27888
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9508 25498 9536 27270
rect 9600 26518 9628 28966
rect 9692 27606 9720 29446
rect 9784 28082 9812 30223
rect 10232 30048 10284 30054
rect 10232 29990 10284 29996
rect 10244 29782 10272 29990
rect 9956 29776 10008 29782
rect 9956 29718 10008 29724
rect 10232 29776 10284 29782
rect 10232 29718 10284 29724
rect 9968 29186 9996 29718
rect 10520 29578 10548 30534
rect 10722 29948 11030 29957
rect 10722 29946 10728 29948
rect 10784 29946 10808 29948
rect 10864 29946 10888 29948
rect 10944 29946 10968 29948
rect 11024 29946 11030 29948
rect 10784 29894 10786 29946
rect 10966 29894 10968 29946
rect 10722 29892 10728 29894
rect 10784 29892 10808 29894
rect 10864 29892 10888 29894
rect 10944 29892 10968 29894
rect 11024 29892 11030 29894
rect 10722 29883 11030 29892
rect 10692 29640 10744 29646
rect 10692 29582 10744 29588
rect 10508 29572 10560 29578
rect 10508 29514 10560 29520
rect 10416 29504 10468 29510
rect 10416 29446 10468 29452
rect 10062 29404 10370 29413
rect 10062 29402 10068 29404
rect 10124 29402 10148 29404
rect 10204 29402 10228 29404
rect 10284 29402 10308 29404
rect 10364 29402 10370 29404
rect 10124 29350 10126 29402
rect 10306 29350 10308 29402
rect 10062 29348 10068 29350
rect 10124 29348 10148 29350
rect 10204 29348 10228 29350
rect 10284 29348 10308 29350
rect 10364 29348 10370 29350
rect 10062 29339 10370 29348
rect 9968 29158 10088 29186
rect 9956 28620 10008 28626
rect 9876 28580 9956 28608
rect 9772 28076 9824 28082
rect 9772 28018 9824 28024
rect 9772 27940 9824 27946
rect 9772 27882 9824 27888
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9692 26926 9720 27542
rect 9680 26920 9732 26926
rect 9680 26862 9732 26868
rect 9588 26512 9640 26518
rect 9586 26480 9588 26489
rect 9640 26480 9642 26489
rect 9586 26415 9642 26424
rect 9692 26296 9720 26862
rect 9600 26268 9720 26296
rect 9600 26042 9628 26268
rect 9588 26036 9640 26042
rect 9588 25978 9640 25984
rect 9784 25922 9812 27882
rect 9600 25894 9812 25922
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9600 24682 9628 25894
rect 9678 25800 9734 25809
rect 9678 25735 9734 25744
rect 9692 24886 9720 25735
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9588 24676 9640 24682
rect 9588 24618 9640 24624
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9508 24274 9536 24550
rect 9496 24268 9548 24274
rect 9496 24210 9548 24216
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9600 24177 9628 24210
rect 9586 24168 9642 24177
rect 9586 24103 9642 24112
rect 9496 24064 9548 24070
rect 9402 24032 9458 24041
rect 9496 24006 9548 24012
rect 9402 23967 9458 23976
rect 9404 23588 9456 23594
rect 9404 23530 9456 23536
rect 9416 23225 9444 23530
rect 9402 23216 9458 23225
rect 9402 23151 9458 23160
rect 9324 23072 9444 23100
rect 9310 22944 9366 22953
rect 9310 22879 9366 22888
rect 9220 22636 9272 22642
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 8852 22160 8904 22166
rect 8850 22128 8852 22137
rect 8904 22128 8906 22137
rect 8850 22063 8906 22072
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8760 22024 8812 22030
rect 8956 22023 8984 22374
rect 9048 22080 9076 22630
rect 9220 22578 9272 22584
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 9140 22409 9168 22510
rect 9126 22400 9182 22409
rect 9126 22335 9182 22344
rect 9220 22092 9272 22098
rect 9048 22052 9168 22080
rect 8760 21966 8812 21972
rect 8864 21995 8984 22023
rect 8588 21690 8616 21966
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8484 21480 8536 21486
rect 8484 21422 8536 21428
rect 8576 21344 8628 21350
rect 8576 21286 8628 21292
rect 8588 21078 8616 21286
rect 8576 21072 8628 21078
rect 8576 21014 8628 21020
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8404 20777 8432 20810
rect 8220 20726 8340 20754
rect 8390 20768 8446 20777
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7944 18170 7972 19110
rect 8116 18760 8168 18766
rect 8022 18728 8078 18737
rect 8116 18702 8168 18708
rect 8022 18663 8078 18672
rect 8036 18290 8064 18663
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7944 18142 8064 18170
rect 7930 18048 7986 18057
rect 7930 17983 7986 17992
rect 7944 17134 7972 17983
rect 8036 17921 8064 18142
rect 8022 17912 8078 17921
rect 8022 17847 8078 17856
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8036 17202 8064 17682
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 8128 17048 8156 18702
rect 8220 17898 8248 20726
rect 8390 20703 8446 20712
rect 8482 20496 8538 20505
rect 8482 20431 8538 20440
rect 8496 20398 8524 20431
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8312 18465 8340 19858
rect 8392 19780 8444 19786
rect 8392 19722 8444 19728
rect 8404 18737 8432 19722
rect 8496 19242 8524 20334
rect 8588 19514 8616 20334
rect 8680 19990 8708 21490
rect 8760 21412 8812 21418
rect 8760 21354 8812 21360
rect 8668 19984 8720 19990
rect 8668 19926 8720 19932
rect 8666 19544 8722 19553
rect 8576 19508 8628 19514
rect 8666 19479 8668 19488
rect 8576 19450 8628 19456
rect 8720 19479 8722 19488
rect 8668 19450 8720 19456
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8390 18728 8446 18737
rect 8390 18663 8446 18672
rect 8298 18456 8354 18465
rect 8298 18391 8354 18400
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8220 17870 8340 17898
rect 8206 17640 8262 17649
rect 8312 17610 8340 17870
rect 8404 17814 8432 18158
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 8496 17746 8524 18090
rect 8588 17898 8616 19314
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8680 18290 8708 18770
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8588 17882 8708 17898
rect 8588 17876 8720 17882
rect 8588 17870 8668 17876
rect 8668 17818 8720 17824
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8496 17649 8524 17682
rect 8482 17640 8538 17649
rect 8206 17575 8262 17584
rect 8300 17604 8352 17610
rect 8220 17202 8248 17575
rect 8482 17575 8538 17584
rect 8300 17546 8352 17552
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8404 17082 8432 17478
rect 8312 17054 8432 17082
rect 8482 17096 8538 17105
rect 8128 17020 8248 17048
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 8114 16960 8170 16969
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 7944 16561 7972 16594
rect 7930 16552 7986 16561
rect 7930 16487 7986 16496
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7208 15694 7420 15722
rect 7656 15700 7708 15706
rect 7208 15570 7236 15694
rect 7656 15642 7708 15648
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 7024 14006 7052 15098
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7116 14396 7144 14894
rect 7300 14890 7328 15506
rect 7484 15026 7512 15574
rect 7562 15192 7618 15201
rect 7562 15127 7618 15136
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 14550 7236 14758
rect 7392 14618 7420 14894
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7484 14550 7512 14962
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7288 14408 7340 14414
rect 7116 14368 7288 14396
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 7116 13802 7144 14368
rect 7288 14350 7340 14356
rect 7392 14346 7420 14418
rect 7576 14362 7604 15127
rect 7668 14550 7696 15642
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7760 14618 7788 14962
rect 7852 14618 7880 15506
rect 7930 15464 7986 15473
rect 7930 15399 7986 15408
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7484 14334 7604 14362
rect 7196 14272 7248 14278
rect 7392 14249 7420 14282
rect 7196 14214 7248 14220
rect 7378 14240 7434 14249
rect 7208 13870 7236 14214
rect 7378 14175 7434 14184
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6656 12260 6868 12288
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6656 11150 6684 12106
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11898 6776 12038
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10810 6684 11086
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6840 10690 6868 12260
rect 6932 11694 6960 13330
rect 7024 13326 7052 13398
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7024 12782 7052 13262
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7116 12306 7144 12582
rect 7208 12374 7236 12650
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7024 11898 7052 12174
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7208 11150 7236 11630
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7196 10736 7248 10742
rect 6840 10662 7144 10690
rect 7196 10678 7248 10684
rect 6920 10600 6972 10606
rect 6564 10577 6920 10588
rect 6550 10568 6920 10577
rect 6276 10532 6328 10538
rect 6606 10560 6920 10568
rect 6920 10542 6972 10548
rect 6550 10503 6606 10512
rect 6276 10474 6328 10480
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6012 10254 6132 10282
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 6012 9654 6040 10134
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5736 7426 5764 9522
rect 6012 9450 6040 9590
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6104 9042 6132 10254
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6196 9926 6224 10066
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6288 9722 6316 10066
rect 6380 9994 6408 10406
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9722 6408 9930
rect 6748 9722 6776 10066
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 5552 7342 5580 7414
rect 5736 7398 6040 7426
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6254 5580 6598
rect 5736 6458 5764 7278
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5828 6254 5856 7210
rect 5920 7002 5948 7278
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5828 5930 5856 6190
rect 5920 6186 5948 6938
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5736 5902 5856 5930
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5552 5250 5580 5646
rect 5736 5574 5764 5902
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5828 5302 5856 5714
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 5368 5222 5580 5250
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5368 5166 5396 5222
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 5368 4706 5396 4966
rect 5460 4826 5488 5102
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5368 4678 5488 4706
rect 5460 4622 5488 4678
rect 5448 4616 5500 4622
rect 4816 4542 4936 4570
rect 5448 4558 5500 4564
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4712 4072 4764 4078
rect 4764 4020 4844 4026
rect 4712 4014 4844 4020
rect 4724 3998 4844 4014
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 4724 3670 4752 3878
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 3058 4476 3334
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4632 2922 4660 3538
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 3608 2032 3660 2038
rect 3608 1974 3660 1980
rect 3620 1902 3648 1974
rect 3608 1896 3660 1902
rect 3608 1838 3660 1844
rect 4080 1834 4108 2246
rect 3516 1828 3568 1834
rect 3516 1770 3568 1776
rect 4068 1828 4120 1834
rect 4068 1770 4120 1776
rect 3528 1494 3556 1770
rect 4172 1494 4200 2246
rect 4252 1828 4304 1834
rect 4252 1770 4304 1776
rect 3516 1488 3568 1494
rect 3516 1430 3568 1436
rect 4160 1488 4212 1494
rect 4160 1430 4212 1436
rect 3528 1222 3556 1430
rect 4264 1358 4292 1770
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 4816 1358 4844 3998
rect 4908 2922 4936 4542
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5000 3058 5028 4014
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5092 2990 5120 4014
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5276 3602 5304 3946
rect 5368 3670 5396 4014
rect 5460 3942 5488 4558
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5276 3126 5304 3538
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5368 3058 5396 3606
rect 5552 3534 5580 4082
rect 5736 4078 5764 4218
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5920 3398 5948 5578
rect 6012 5166 6040 7398
rect 6104 6746 6132 8842
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6564 7954 6592 8026
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6196 6866 6224 7278
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6866 6316 7142
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6104 6718 6224 6746
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6012 4690 6040 5102
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6012 4078 6040 4626
rect 6104 4486 6132 6122
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3738 6132 3878
rect 6196 3738 6224 6718
rect 6380 6458 6408 7278
rect 6472 7274 6500 7890
rect 6564 7342 6592 7890
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6472 5710 6500 6190
rect 6564 6186 6592 7142
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6564 5166 6592 6122
rect 6656 5234 6684 9454
rect 6748 9450 6776 9658
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6932 8294 6960 10542
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7024 10266 7052 10474
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6932 8266 7052 8294
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7546 6776 7822
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6748 5030 6776 7210
rect 6932 6866 6960 7686
rect 7024 7206 7052 8266
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6828 6792 6880 6798
rect 6918 6760 6974 6769
rect 6880 6740 6918 6746
rect 6828 6734 6918 6740
rect 6840 6718 6918 6734
rect 6918 6695 6974 6704
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 5846 6868 6598
rect 7116 6458 7144 10662
rect 7208 10606 7236 10678
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7300 10266 7328 13194
rect 7392 12306 7420 13874
rect 7484 12646 7512 14334
rect 7746 13696 7802 13705
rect 7746 13631 7802 13640
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7668 12782 7696 13126
rect 7760 12782 7788 13631
rect 7944 13530 7972 15399
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7944 13394 7972 13466
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 8036 13274 8064 16934
rect 8114 16895 8170 16904
rect 8128 15162 8156 16895
rect 8220 15570 8248 17020
rect 8312 16726 8340 17054
rect 8482 17031 8484 17040
rect 8536 17031 8538 17040
rect 8484 17002 8536 17008
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8300 16720 8352 16726
rect 8404 16697 8432 16934
rect 8300 16662 8352 16668
rect 8390 16688 8446 16697
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8220 15473 8248 15506
rect 8206 15464 8262 15473
rect 8206 15399 8262 15408
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8220 14958 8248 15302
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8128 13938 8156 14282
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8114 13560 8170 13569
rect 8114 13495 8170 13504
rect 8128 13394 8156 13495
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8036 13246 8248 13274
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7838 12880 7894 12889
rect 8036 12850 8064 13126
rect 7838 12815 7894 12824
rect 8024 12844 8076 12850
rect 7852 12782 7880 12815
rect 8024 12786 8076 12792
rect 7656 12776 7708 12782
rect 7576 12724 7656 12730
rect 7576 12718 7708 12724
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7576 12702 7696 12718
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7208 9518 7236 10066
rect 7300 9586 7328 10202
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 7342 7236 9318
rect 7392 8498 7420 11494
rect 7484 10810 7512 11630
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7392 7954 7420 8434
rect 7576 7970 7604 12702
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7668 9178 7696 12582
rect 7852 11082 7880 12582
rect 7944 12374 7972 12718
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 8036 12306 8064 12786
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8128 12306 8156 12718
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 11898 8156 12038
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8036 11558 8064 11698
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7852 10452 7880 11018
rect 7944 10742 7972 11018
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7944 10606 7972 10678
rect 8220 10674 8248 13246
rect 8312 12073 8340 16662
rect 8390 16623 8446 16632
rect 8588 16130 8616 17750
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8680 16794 8708 17682
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8496 16102 8616 16130
rect 8390 15736 8446 15745
rect 8390 15671 8392 15680
rect 8444 15671 8446 15680
rect 8392 15642 8444 15648
rect 8404 15570 8432 15642
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8390 15464 8446 15473
rect 8390 15399 8446 15408
rect 8404 14482 8432 15399
rect 8496 14521 8524 16102
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8588 15706 8616 15982
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8680 15570 8708 16186
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8588 15094 8616 15302
rect 8772 15162 8800 21354
rect 8864 20942 8892 21995
rect 9034 21992 9090 22001
rect 9034 21927 9090 21936
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 8956 21554 8984 21626
rect 9048 21593 9076 21927
rect 9034 21584 9090 21593
rect 8944 21548 8996 21554
rect 9034 21519 9090 21528
rect 8944 21490 8996 21496
rect 8944 21412 8996 21418
rect 8944 21354 8996 21360
rect 8852 20936 8904 20942
rect 8850 20904 8852 20913
rect 8904 20904 8906 20913
rect 8850 20839 8906 20848
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8864 19310 8892 19654
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8864 16250 8892 19110
rect 8956 16969 8984 21354
rect 9140 21078 9168 22052
rect 9220 22034 9272 22040
rect 9232 21690 9260 22034
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9218 21584 9274 21593
rect 9324 21554 9352 22879
rect 9416 22030 9444 23072
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9416 21729 9444 21966
rect 9402 21720 9458 21729
rect 9402 21655 9458 21664
rect 9218 21519 9274 21528
rect 9312 21548 9364 21554
rect 9232 21400 9260 21519
rect 9312 21490 9364 21496
rect 9232 21372 9352 21400
rect 9128 21072 9180 21078
rect 9128 21014 9180 21020
rect 9218 21040 9274 21049
rect 9218 20975 9274 20984
rect 9128 20936 9180 20942
rect 9034 20904 9090 20913
rect 9128 20878 9180 20884
rect 9034 20839 9090 20848
rect 9048 20210 9076 20839
rect 9140 20777 9168 20878
rect 9126 20768 9182 20777
rect 9126 20703 9182 20712
rect 9126 20224 9182 20233
rect 9048 20182 9126 20210
rect 9126 20159 9182 20168
rect 9140 19922 9168 20159
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9048 19174 9076 19858
rect 9126 19544 9182 19553
rect 9126 19479 9182 19488
rect 9140 19446 9168 19479
rect 9128 19440 9180 19446
rect 9128 19382 9180 19388
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 9140 18873 9168 19246
rect 9126 18864 9182 18873
rect 9126 18799 9182 18808
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 9048 18358 9076 18702
rect 9126 18592 9182 18601
rect 9232 18578 9260 20975
rect 9324 20482 9352 21372
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9416 20602 9444 20946
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9324 20454 9444 20482
rect 9508 20466 9536 24006
rect 9588 23656 9640 23662
rect 9586 23624 9588 23633
rect 9640 23624 9642 23633
rect 9586 23559 9642 23568
rect 9588 23520 9640 23526
rect 9586 23488 9588 23497
rect 9640 23488 9642 23497
rect 9586 23423 9642 23432
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 9600 22982 9628 23122
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9692 22710 9720 24686
rect 9784 24342 9812 25434
rect 9876 24410 9904 28580
rect 9956 28562 10008 28568
rect 10060 28506 10088 29158
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10152 28529 10180 28902
rect 10428 28626 10456 29446
rect 10704 28966 10732 29582
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10722 28860 11030 28869
rect 10722 28858 10728 28860
rect 10784 28858 10808 28860
rect 10864 28858 10888 28860
rect 10944 28858 10968 28860
rect 11024 28858 11030 28860
rect 10784 28806 10786 28858
rect 10966 28806 10968 28858
rect 10722 28804 10728 28806
rect 10784 28804 10808 28806
rect 10864 28804 10888 28806
rect 10944 28804 10968 28806
rect 11024 28804 11030 28806
rect 10722 28795 11030 28804
rect 10416 28620 10468 28626
rect 10416 28562 10468 28568
rect 9968 28478 10088 28506
rect 10138 28520 10194 28529
rect 9968 28200 9996 28478
rect 10138 28455 10194 28464
rect 10508 28484 10560 28490
rect 10508 28426 10560 28432
rect 10062 28316 10370 28325
rect 10062 28314 10068 28316
rect 10124 28314 10148 28316
rect 10204 28314 10228 28316
rect 10284 28314 10308 28316
rect 10364 28314 10370 28316
rect 10124 28262 10126 28314
rect 10306 28262 10308 28314
rect 10062 28260 10068 28262
rect 10124 28260 10148 28262
rect 10204 28260 10228 28262
rect 10284 28260 10308 28262
rect 10364 28260 10370 28262
rect 10062 28251 10370 28260
rect 10140 28212 10192 28218
rect 9968 28172 10088 28200
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 9968 26314 9996 28018
rect 10060 27946 10088 28172
rect 10140 28154 10192 28160
rect 10048 27940 10100 27946
rect 10048 27882 10100 27888
rect 10152 27441 10180 28154
rect 10416 28008 10468 28014
rect 10416 27950 10468 27956
rect 10138 27432 10194 27441
rect 10138 27367 10194 27376
rect 10062 27228 10370 27237
rect 10062 27226 10068 27228
rect 10124 27226 10148 27228
rect 10204 27226 10228 27228
rect 10284 27226 10308 27228
rect 10364 27226 10370 27228
rect 10124 27174 10126 27226
rect 10306 27174 10308 27226
rect 10062 27172 10068 27174
rect 10124 27172 10148 27174
rect 10204 27172 10228 27174
rect 10284 27172 10308 27174
rect 10364 27172 10370 27174
rect 10062 27163 10370 27172
rect 10140 27124 10192 27130
rect 10140 27066 10192 27072
rect 10046 27024 10102 27033
rect 10046 26959 10102 26968
rect 10060 26353 10088 26959
rect 10152 26450 10180 27066
rect 10140 26444 10192 26450
rect 10140 26386 10192 26392
rect 10046 26344 10102 26353
rect 9956 26308 10008 26314
rect 10046 26279 10102 26288
rect 9956 26250 10008 26256
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 9772 24336 9824 24342
rect 9772 24278 9824 24284
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9876 24070 9904 24142
rect 9864 24064 9916 24070
rect 9770 24032 9826 24041
rect 9864 24006 9916 24012
rect 9770 23967 9826 23976
rect 9784 23662 9812 23967
rect 9876 23780 9904 24006
rect 9968 23848 9996 26250
rect 10060 26246 10088 26279
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 10062 26140 10370 26149
rect 10062 26138 10068 26140
rect 10124 26138 10148 26140
rect 10204 26138 10228 26140
rect 10284 26138 10308 26140
rect 10364 26138 10370 26140
rect 10124 26086 10126 26138
rect 10306 26086 10308 26138
rect 10062 26084 10068 26086
rect 10124 26084 10148 26086
rect 10204 26084 10228 26086
rect 10284 26084 10308 26086
rect 10364 26084 10370 26086
rect 10062 26075 10370 26084
rect 10048 25968 10100 25974
rect 10048 25910 10100 25916
rect 10060 25226 10088 25910
rect 10048 25220 10100 25226
rect 10048 25162 10100 25168
rect 10062 25052 10370 25061
rect 10062 25050 10068 25052
rect 10124 25050 10148 25052
rect 10204 25050 10228 25052
rect 10284 25050 10308 25052
rect 10364 25050 10370 25052
rect 10124 24998 10126 25050
rect 10306 24998 10308 25050
rect 10062 24996 10068 24998
rect 10124 24996 10148 24998
rect 10204 24996 10228 24998
rect 10284 24996 10308 24998
rect 10364 24996 10370 24998
rect 10062 24987 10370 24996
rect 10232 24880 10284 24886
rect 10232 24822 10284 24828
rect 10048 24744 10100 24750
rect 10046 24712 10048 24721
rect 10100 24712 10102 24721
rect 10046 24647 10102 24656
rect 10140 24676 10192 24682
rect 10140 24618 10192 24624
rect 10152 24206 10180 24618
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10244 24070 10272 24822
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10336 24177 10364 24754
rect 10428 24274 10456 27950
rect 10520 26858 10548 28426
rect 11072 28150 11100 34614
rect 11060 28144 11112 28150
rect 11060 28086 11112 28092
rect 10600 28076 10652 28082
rect 10600 28018 10652 28024
rect 10508 26852 10560 26858
rect 10508 26794 10560 26800
rect 10508 26240 10560 26246
rect 10508 26182 10560 26188
rect 10520 25838 10548 26182
rect 10612 25838 10640 28018
rect 11058 27976 11114 27985
rect 11058 27911 11114 27920
rect 10722 27772 11030 27781
rect 10722 27770 10728 27772
rect 10784 27770 10808 27772
rect 10864 27770 10888 27772
rect 10944 27770 10968 27772
rect 11024 27770 11030 27772
rect 10784 27718 10786 27770
rect 10966 27718 10968 27770
rect 10722 27716 10728 27718
rect 10784 27716 10808 27718
rect 10864 27716 10888 27718
rect 10944 27716 10968 27718
rect 11024 27716 11030 27718
rect 10722 27707 11030 27716
rect 10690 27568 10746 27577
rect 10690 27503 10746 27512
rect 10704 27334 10732 27503
rect 10692 27328 10744 27334
rect 10692 27270 10744 27276
rect 10704 26897 10732 27270
rect 10690 26888 10746 26897
rect 10690 26823 10746 26832
rect 10722 26684 11030 26693
rect 10722 26682 10728 26684
rect 10784 26682 10808 26684
rect 10864 26682 10888 26684
rect 10944 26682 10968 26684
rect 11024 26682 11030 26684
rect 10784 26630 10786 26682
rect 10966 26630 10968 26682
rect 10722 26628 10728 26630
rect 10784 26628 10808 26630
rect 10864 26628 10888 26630
rect 10944 26628 10968 26630
rect 11024 26628 11030 26630
rect 10722 26619 11030 26628
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 10520 25362 10548 25774
rect 10508 25356 10560 25362
rect 10508 25298 10560 25304
rect 10520 24818 10548 25298
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10612 24750 10640 25774
rect 10722 25596 11030 25605
rect 10722 25594 10728 25596
rect 10784 25594 10808 25596
rect 10864 25594 10888 25596
rect 10944 25594 10968 25596
rect 11024 25594 11030 25596
rect 10784 25542 10786 25594
rect 10966 25542 10968 25594
rect 10722 25540 10728 25542
rect 10784 25540 10808 25542
rect 10864 25540 10888 25542
rect 10944 25540 10968 25542
rect 11024 25540 11030 25542
rect 10722 25531 11030 25540
rect 10690 25256 10746 25265
rect 11072 25242 11100 27911
rect 10690 25191 10746 25200
rect 10980 25214 11100 25242
rect 10600 24744 10652 24750
rect 10600 24686 10652 24692
rect 10508 24676 10560 24682
rect 10508 24618 10560 24624
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10322 24168 10378 24177
rect 10322 24103 10378 24112
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 10062 23964 10370 23973
rect 10062 23962 10068 23964
rect 10124 23962 10148 23964
rect 10204 23962 10228 23964
rect 10284 23962 10308 23964
rect 10364 23962 10370 23964
rect 10124 23910 10126 23962
rect 10306 23910 10308 23962
rect 10062 23908 10068 23910
rect 10124 23908 10148 23910
rect 10204 23908 10228 23910
rect 10284 23908 10308 23910
rect 10364 23908 10370 23910
rect 10062 23899 10370 23908
rect 10428 23866 10456 24210
rect 10140 23860 10192 23866
rect 9968 23820 10088 23848
rect 9876 23752 9996 23780
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9864 23520 9916 23526
rect 9864 23462 9916 23468
rect 9784 23118 9812 23462
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9680 22092 9732 22098
rect 9784 22080 9812 23054
rect 9732 22052 9812 22080
rect 9680 22034 9732 22040
rect 9692 22001 9720 22034
rect 9678 21992 9734 22001
rect 9678 21927 9734 21936
rect 9588 21888 9640 21894
rect 9586 21856 9588 21865
rect 9680 21888 9732 21894
rect 9640 21856 9642 21865
rect 9680 21830 9732 21836
rect 9586 21791 9642 21800
rect 9692 21593 9720 21830
rect 9678 21584 9734 21593
rect 9600 21542 9678 21570
rect 9600 21486 9628 21542
rect 9678 21519 9734 21528
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9770 21312 9826 21321
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9324 18766 9352 19246
rect 9416 19174 9444 20454
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 9508 19786 9536 20402
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9600 18902 9628 21286
rect 9770 21247 9826 21256
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9784 20754 9812 21247
rect 9876 21146 9904 23462
rect 9968 23089 9996 23752
rect 10060 23662 10088 23820
rect 10140 23802 10192 23808
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10152 23730 10180 23802
rect 10322 23760 10378 23769
rect 10140 23724 10192 23730
rect 10322 23695 10378 23704
rect 10140 23666 10192 23672
rect 10336 23662 10364 23695
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 10324 23656 10376 23662
rect 10376 23616 10456 23644
rect 10324 23598 10376 23604
rect 10322 23488 10378 23497
rect 10322 23423 10378 23432
rect 10336 23322 10364 23423
rect 10324 23316 10376 23322
rect 10324 23258 10376 23264
rect 10138 23216 10194 23225
rect 10138 23151 10140 23160
rect 10192 23151 10194 23160
rect 10140 23122 10192 23128
rect 9954 23080 10010 23089
rect 9954 23015 10010 23024
rect 9968 22080 9996 23015
rect 10062 22876 10370 22885
rect 10062 22874 10068 22876
rect 10124 22874 10148 22876
rect 10204 22874 10228 22876
rect 10284 22874 10308 22876
rect 10364 22874 10370 22876
rect 10124 22822 10126 22874
rect 10306 22822 10308 22874
rect 10062 22820 10068 22822
rect 10124 22820 10148 22822
rect 10204 22820 10228 22822
rect 10284 22820 10308 22822
rect 10364 22820 10370 22822
rect 10062 22811 10370 22820
rect 10428 22658 10456 23616
rect 10520 22982 10548 24618
rect 10704 24596 10732 25191
rect 10980 24682 11008 25214
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 10968 24676 11020 24682
rect 10968 24618 11020 24624
rect 10612 24568 10732 24596
rect 10612 24154 10640 24568
rect 10722 24508 11030 24517
rect 10722 24506 10728 24508
rect 10784 24506 10808 24508
rect 10864 24506 10888 24508
rect 10944 24506 10968 24508
rect 11024 24506 11030 24508
rect 10784 24454 10786 24506
rect 10966 24454 10968 24506
rect 10722 24452 10728 24454
rect 10784 24452 10808 24454
rect 10864 24452 10888 24454
rect 10944 24452 10968 24454
rect 11024 24452 11030 24454
rect 10722 24443 11030 24452
rect 10782 24304 10838 24313
rect 10782 24239 10838 24248
rect 10966 24304 11022 24313
rect 10966 24239 11022 24248
rect 10612 24126 10732 24154
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10336 22630 10456 22658
rect 10520 22642 10548 22918
rect 10508 22636 10560 22642
rect 10336 22166 10364 22630
rect 10508 22578 10560 22584
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10428 22234 10456 22510
rect 10416 22228 10468 22234
rect 10416 22170 10468 22176
rect 10324 22160 10376 22166
rect 10324 22102 10376 22108
rect 10048 22092 10100 22098
rect 9968 22052 10048 22080
rect 9968 21486 9996 22052
rect 10048 22034 10100 22040
rect 10416 22092 10468 22098
rect 10416 22034 10468 22040
rect 10062 21788 10370 21797
rect 10062 21786 10068 21788
rect 10124 21786 10148 21788
rect 10204 21786 10228 21788
rect 10284 21786 10308 21788
rect 10364 21786 10370 21788
rect 10124 21734 10126 21786
rect 10306 21734 10308 21786
rect 10062 21732 10068 21734
rect 10124 21732 10148 21734
rect 10204 21732 10228 21734
rect 10284 21732 10308 21734
rect 10364 21732 10370 21734
rect 10062 21723 10370 21732
rect 10428 21690 10456 22034
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9876 20874 9904 21082
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 9692 19514 9720 20742
rect 9784 20726 9904 20754
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9784 20262 9812 20334
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9784 19990 9812 20198
rect 9772 19984 9824 19990
rect 9772 19926 9824 19932
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9692 19292 9720 19450
rect 9772 19304 9824 19310
rect 9692 19264 9772 19292
rect 9772 19246 9824 19252
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9588 18896 9640 18902
rect 9588 18838 9640 18844
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9232 18550 9352 18578
rect 9126 18527 9182 18536
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9140 17678 9168 18527
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9048 17202 9076 17546
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 8942 16960 8998 16969
rect 8942 16895 8998 16904
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8864 15609 8892 15982
rect 8850 15600 8906 15609
rect 8850 15535 8906 15544
rect 8956 15434 8984 16594
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 8944 15428 8996 15434
rect 8944 15370 8996 15376
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8574 14920 8630 14929
rect 8574 14855 8630 14864
rect 8482 14512 8538 14521
rect 8392 14476 8444 14482
rect 8482 14447 8538 14456
rect 8392 14418 8444 14424
rect 8496 14074 8524 14447
rect 8588 14362 8616 14855
rect 8680 14618 8708 14962
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8772 14793 8800 14826
rect 8758 14784 8814 14793
rect 8758 14719 8814 14728
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8588 14334 8708 14362
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 13394 8524 13806
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8496 12646 8524 13330
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12442 8524 12582
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8496 12209 8524 12242
rect 8482 12200 8538 12209
rect 8482 12135 8538 12144
rect 8298 12064 8354 12073
rect 8298 11999 8354 12008
rect 8298 11792 8354 11801
rect 8298 11727 8354 11736
rect 8482 11792 8538 11801
rect 8482 11727 8484 11736
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7852 10424 7972 10452
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8634 7788 8910
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7852 8362 7880 9318
rect 7944 8838 7972 10424
rect 8312 9110 8340 11727
rect 8536 11727 8538 11736
rect 8484 11698 8536 11704
rect 8390 11656 8446 11665
rect 8390 11591 8446 11600
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 8036 8566 8064 8910
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7852 8242 7880 8298
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7484 7942 7604 7970
rect 7760 8214 7880 8242
rect 7760 7954 7788 8214
rect 7944 8022 7972 8366
rect 8220 8362 8248 8910
rect 8312 8838 8340 8910
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8312 8498 8340 8774
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7656 7948 7708 7954
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7300 6390 7328 7686
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6932 5710 6960 6190
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6932 5370 6960 5646
rect 7116 5370 7144 6122
rect 7208 5914 7236 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7300 5778 7328 6326
rect 7392 6322 7420 7482
rect 7484 6934 7512 7942
rect 7656 7890 7708 7896
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7576 7546 7604 7822
rect 7668 7818 7696 7890
rect 8312 7886 8340 8230
rect 8404 8090 8432 11591
rect 8588 11218 8616 14214
rect 8680 12918 8708 14334
rect 8772 14006 8800 14418
rect 8864 14414 8892 15370
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8956 15026 8984 15098
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8956 14550 8984 14758
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8668 12232 8720 12238
rect 8772 12220 8800 13670
rect 8864 12434 8892 14010
rect 8944 14000 8996 14006
rect 8942 13968 8944 13977
rect 8996 13968 8998 13977
rect 8942 13903 8998 13912
rect 8864 12406 8984 12434
rect 8720 12192 8800 12220
rect 8668 12174 8720 12180
rect 8680 11558 8708 12174
rect 8850 11792 8906 11801
rect 8850 11727 8852 11736
rect 8904 11727 8906 11736
rect 8852 11698 8904 11704
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8680 11098 8708 11494
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8588 11070 8708 11098
rect 8588 9518 8616 11070
rect 8668 9988 8720 9994
rect 8668 9930 8720 9936
rect 8680 9586 8708 9930
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8496 8974 8524 9454
rect 8680 9042 8708 9522
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7668 7546 7696 7754
rect 8404 7750 8432 7890
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7484 6322 7512 6870
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4282 7236 4966
rect 7300 4690 7328 5102
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5736 2990 5764 3334
rect 6196 3194 6224 3538
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 6656 2922 6684 3538
rect 6748 3534 6776 3878
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 7208 3194 7236 4218
rect 7300 3534 7328 4626
rect 7576 4486 7604 7346
rect 8496 7342 8524 8910
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8588 8634 8616 8842
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8588 8362 8616 8570
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8772 7410 8800 11154
rect 8864 10606 8892 11222
rect 8956 11218 8984 12406
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8864 9722 8892 10066
rect 8956 10062 8984 10406
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8220 6866 8248 6938
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 4826 7880 5714
rect 8036 5642 8064 6802
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8128 5914 8156 6190
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7852 4078 7880 4490
rect 7944 4078 7972 4966
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8036 4214 8064 4626
rect 8496 4486 8524 5306
rect 8588 4486 8616 5510
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8680 4758 8708 4966
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8496 4214 8524 4422
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5184 2106 5212 2450
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6932 2106 6960 2246
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 6920 2100 6972 2106
rect 6920 2042 6972 2048
rect 7024 2038 7052 2790
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7116 2106 7144 2450
rect 7104 2100 7156 2106
rect 7104 2042 7156 2048
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 7208 1902 7236 3130
rect 7300 2922 7328 3334
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7576 1970 7604 3538
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7760 2922 7788 3402
rect 8036 3398 8064 3975
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7944 2990 7972 3334
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7760 1970 7788 2858
rect 7852 2650 7880 2858
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 7748 1964 7800 1970
rect 7748 1906 7800 1912
rect 7944 1902 7972 2926
rect 8036 2650 8064 3334
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8128 2106 8156 3606
rect 8312 3602 8340 3674
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8312 3194 8340 3538
rect 8772 3482 8800 7210
rect 8864 6798 8892 8434
rect 8956 8430 8984 9318
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8956 7546 8984 7890
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8864 5846 8892 6734
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8956 4826 8984 5714
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8942 4040 8998 4049
rect 8942 3975 8998 3984
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8864 3602 8892 3878
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8772 3454 8892 3482
rect 8864 3398 8892 3454
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8772 2922 8800 3334
rect 8956 3194 8984 3975
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8956 2650 8984 3130
rect 9048 3058 9076 17138
rect 9126 16688 9182 16697
rect 9126 16623 9128 16632
rect 9180 16623 9182 16632
rect 9128 16594 9180 16600
rect 9232 16046 9260 18022
rect 9324 17105 9352 18550
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9416 17746 9444 18226
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9508 17610 9536 18634
rect 9600 18358 9628 18838
rect 9678 18728 9734 18737
rect 9678 18663 9680 18672
rect 9732 18663 9734 18672
rect 9680 18634 9732 18640
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9692 18222 9720 18634
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9784 17954 9812 19110
rect 9692 17926 9812 17954
rect 9692 17882 9720 17926
rect 9876 17898 9904 20726
rect 9680 17876 9732 17882
rect 9600 17836 9680 17864
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9310 17096 9366 17105
rect 9310 17031 9366 17040
rect 9416 16980 9444 17546
rect 9508 17066 9536 17546
rect 9496 17060 9548 17066
rect 9496 17002 9548 17008
rect 9324 16952 9444 16980
rect 9324 16114 9352 16952
rect 9402 16552 9458 16561
rect 9402 16487 9458 16496
rect 9416 16454 9444 16487
rect 9508 16454 9536 17002
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9232 15434 9260 15982
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 15706 9352 15846
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9416 15586 9444 16050
rect 9508 15706 9536 16390
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9324 15570 9444 15586
rect 9312 15564 9444 15570
rect 9364 15558 9444 15564
rect 9496 15564 9548 15570
rect 9312 15506 9364 15512
rect 9496 15506 9548 15512
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9218 15328 9274 15337
rect 9218 15263 9274 15272
rect 9232 13802 9260 15263
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9232 13530 9260 13738
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9232 13326 9260 13466
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9126 13016 9182 13025
rect 9126 12951 9128 12960
rect 9180 12951 9182 12960
rect 9128 12922 9180 12928
rect 9324 12918 9352 15506
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9416 15162 9444 15302
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9402 15056 9458 15065
rect 9402 14991 9404 15000
rect 9456 14991 9458 15000
rect 9404 14962 9456 14968
rect 9402 14512 9458 14521
rect 9402 14447 9458 14456
rect 9416 14414 9444 14447
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9508 14278 9536 15506
rect 9600 15502 9628 17836
rect 9680 17818 9732 17824
rect 9784 17870 9904 17898
rect 9680 17672 9732 17678
rect 9678 17640 9680 17649
rect 9732 17640 9734 17649
rect 9678 17575 9734 17584
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9692 16776 9720 17002
rect 9784 16969 9812 17870
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9876 16998 9904 17682
rect 9968 17134 9996 21422
rect 10140 21412 10192 21418
rect 10140 21354 10192 21360
rect 10152 21049 10180 21354
rect 10138 21040 10194 21049
rect 10138 20975 10194 20984
rect 10048 20936 10100 20942
rect 10046 20904 10048 20913
rect 10100 20904 10102 20913
rect 10046 20839 10102 20848
rect 10062 20700 10370 20709
rect 10062 20698 10068 20700
rect 10124 20698 10148 20700
rect 10204 20698 10228 20700
rect 10284 20698 10308 20700
rect 10364 20698 10370 20700
rect 10124 20646 10126 20698
rect 10306 20646 10308 20698
rect 10062 20644 10068 20646
rect 10124 20644 10148 20646
rect 10204 20644 10228 20646
rect 10284 20644 10308 20646
rect 10364 20644 10370 20646
rect 10062 20635 10370 20644
rect 10428 20618 10456 21626
rect 10520 21146 10548 22578
rect 10612 21962 10640 24006
rect 10704 23526 10732 24126
rect 10796 24041 10824 24239
rect 10782 24032 10838 24041
rect 10782 23967 10838 23976
rect 10980 23610 11008 24239
rect 11072 23730 11100 25094
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 10980 23582 11100 23610
rect 10692 23520 10744 23526
rect 10692 23462 10744 23468
rect 10722 23420 11030 23429
rect 10722 23418 10728 23420
rect 10784 23418 10808 23420
rect 10864 23418 10888 23420
rect 10944 23418 10968 23420
rect 11024 23418 11030 23420
rect 10784 23366 10786 23418
rect 10966 23366 10968 23418
rect 10722 23364 10728 23366
rect 10784 23364 10808 23366
rect 10864 23364 10888 23366
rect 10944 23364 10968 23366
rect 11024 23364 11030 23366
rect 10722 23355 11030 23364
rect 10692 23248 10744 23254
rect 10690 23216 10692 23225
rect 10744 23216 10746 23225
rect 10690 23151 10746 23160
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10796 22778 10824 22986
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 10722 22332 11030 22341
rect 10722 22330 10728 22332
rect 10784 22330 10808 22332
rect 10864 22330 10888 22332
rect 10944 22330 10968 22332
rect 11024 22330 11030 22332
rect 10784 22278 10786 22330
rect 10966 22278 10968 22330
rect 10722 22276 10728 22278
rect 10784 22276 10808 22278
rect 10864 22276 10888 22278
rect 10944 22276 10968 22278
rect 11024 22276 11030 22278
rect 10722 22267 11030 22276
rect 10692 22160 10744 22166
rect 10692 22102 10744 22108
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10598 21856 10654 21865
rect 10598 21791 10654 21800
rect 10508 21140 10560 21146
rect 10612 21128 10640 21791
rect 10704 21418 10732 22102
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10722 21244 11030 21253
rect 10722 21242 10728 21244
rect 10784 21242 10808 21244
rect 10864 21242 10888 21244
rect 10944 21242 10968 21244
rect 11024 21242 11030 21244
rect 10784 21190 10786 21242
rect 10966 21190 10968 21242
rect 10722 21188 10728 21190
rect 10784 21188 10808 21190
rect 10864 21188 10888 21190
rect 10944 21188 10968 21190
rect 11024 21188 11030 21190
rect 10722 21179 11030 21188
rect 10612 21100 10732 21128
rect 10508 21082 10560 21088
rect 10428 20590 10640 20618
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10062 19612 10370 19621
rect 10062 19610 10068 19612
rect 10124 19610 10148 19612
rect 10204 19610 10228 19612
rect 10284 19610 10308 19612
rect 10364 19610 10370 19612
rect 10124 19558 10126 19610
rect 10306 19558 10308 19610
rect 10062 19556 10068 19558
rect 10124 19556 10148 19558
rect 10204 19556 10228 19558
rect 10284 19556 10308 19558
rect 10364 19556 10370 19558
rect 10062 19547 10370 19556
rect 10428 19378 10456 19654
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10062 18524 10370 18533
rect 10062 18522 10068 18524
rect 10124 18522 10148 18524
rect 10204 18522 10228 18524
rect 10284 18522 10308 18524
rect 10364 18522 10370 18524
rect 10124 18470 10126 18522
rect 10306 18470 10308 18522
rect 10062 18468 10068 18470
rect 10124 18468 10148 18470
rect 10204 18468 10228 18470
rect 10284 18468 10308 18470
rect 10364 18468 10370 18470
rect 10062 18459 10370 18468
rect 10062 17436 10370 17445
rect 10062 17434 10068 17436
rect 10124 17434 10148 17436
rect 10204 17434 10228 17436
rect 10284 17434 10308 17436
rect 10364 17434 10370 17436
rect 10124 17382 10126 17434
rect 10306 17382 10308 17434
rect 10062 17380 10068 17382
rect 10124 17380 10148 17382
rect 10204 17380 10228 17382
rect 10284 17380 10308 17382
rect 10364 17380 10370 17382
rect 10062 17371 10370 17380
rect 10428 17338 10456 18906
rect 10520 18834 10548 20402
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10520 18290 10548 18770
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9864 16992 9916 16998
rect 9770 16960 9826 16969
rect 9864 16934 9916 16940
rect 9770 16895 9826 16904
rect 9772 16788 9824 16794
rect 9692 16748 9772 16776
rect 9772 16730 9824 16736
rect 9678 16688 9734 16697
rect 9678 16623 9734 16632
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9600 14793 9628 15030
rect 9586 14784 9642 14793
rect 9586 14719 9642 14728
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9600 14006 9628 14719
rect 9588 14000 9640 14006
rect 9494 13968 9550 13977
rect 9588 13942 9640 13948
rect 9494 13903 9550 13912
rect 9508 13802 9536 13903
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9600 13462 9628 13942
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9324 12442 9352 12718
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9140 11898 9168 12242
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9140 11218 9168 11834
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9232 9602 9260 12174
rect 9324 11200 9352 12242
rect 9416 11354 9444 12718
rect 9508 12646 9536 13126
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9508 11286 9536 12582
rect 9600 11626 9628 13262
rect 9692 12850 9720 16623
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9784 15745 9812 15914
rect 9770 15736 9826 15745
rect 9770 15671 9826 15680
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9784 14618 9812 15574
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9784 14278 9812 14418
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9876 13394 9904 16934
rect 9968 16658 9996 17070
rect 10232 17060 10284 17066
rect 10428 17048 10456 17274
rect 10232 17002 10284 17008
rect 10336 17020 10456 17048
rect 10244 16726 10272 17002
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9968 16250 9996 16458
rect 10152 16454 10180 16526
rect 10336 16522 10364 17020
rect 10612 16946 10640 20590
rect 10704 20369 10732 21100
rect 10690 20360 10746 20369
rect 10690 20295 10746 20304
rect 10722 20156 11030 20165
rect 10722 20154 10728 20156
rect 10784 20154 10808 20156
rect 10864 20154 10888 20156
rect 10944 20154 10968 20156
rect 11024 20154 11030 20156
rect 10784 20102 10786 20154
rect 10966 20102 10968 20154
rect 10722 20100 10728 20102
rect 10784 20100 10808 20102
rect 10864 20100 10888 20102
rect 10944 20100 10968 20102
rect 11024 20100 11030 20102
rect 10722 20091 11030 20100
rect 10722 19068 11030 19077
rect 10722 19066 10728 19068
rect 10784 19066 10808 19068
rect 10864 19066 10888 19068
rect 10944 19066 10968 19068
rect 11024 19066 11030 19068
rect 10784 19014 10786 19066
rect 10966 19014 10968 19066
rect 10722 19012 10728 19014
rect 10784 19012 10808 19014
rect 10864 19012 10888 19014
rect 10944 19012 10968 19014
rect 11024 19012 11030 19014
rect 10722 19003 11030 19012
rect 10722 17980 11030 17989
rect 10722 17978 10728 17980
rect 10784 17978 10808 17980
rect 10864 17978 10888 17980
rect 10944 17978 10968 17980
rect 11024 17978 11030 17980
rect 10784 17926 10786 17978
rect 10966 17926 10968 17978
rect 10722 17924 10728 17926
rect 10784 17924 10808 17926
rect 10864 17924 10888 17926
rect 10944 17924 10968 17926
rect 11024 17924 11030 17926
rect 10722 17915 11030 17924
rect 10428 16918 10640 16946
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10062 16348 10370 16357
rect 10062 16346 10068 16348
rect 10124 16346 10148 16348
rect 10204 16346 10228 16348
rect 10284 16346 10308 16348
rect 10364 16346 10370 16348
rect 10124 16294 10126 16346
rect 10306 16294 10308 16346
rect 10062 16292 10068 16294
rect 10124 16292 10148 16294
rect 10204 16292 10228 16294
rect 10284 16292 10308 16294
rect 10364 16292 10370 16294
rect 10062 16283 10370 16292
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 15162 9996 15506
rect 10062 15260 10370 15269
rect 10062 15258 10068 15260
rect 10124 15258 10148 15260
rect 10204 15258 10228 15260
rect 10284 15258 10308 15260
rect 10364 15258 10370 15260
rect 10124 15206 10126 15258
rect 10306 15206 10308 15258
rect 10062 15204 10068 15206
rect 10124 15204 10148 15206
rect 10204 15204 10228 15206
rect 10284 15204 10308 15206
rect 10364 15204 10370 15206
rect 10062 15195 10370 15204
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9954 15056 10010 15065
rect 9954 14991 10010 15000
rect 10232 15020 10284 15026
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9968 12986 9996 14991
rect 10232 14962 10284 14968
rect 10244 14618 10272 14962
rect 10324 14952 10376 14958
rect 10428 14940 10456 16918
rect 10722 16892 11030 16901
rect 10722 16890 10728 16892
rect 10784 16890 10808 16892
rect 10864 16890 10888 16892
rect 10944 16890 10968 16892
rect 11024 16890 11030 16892
rect 10784 16838 10786 16890
rect 10966 16838 10968 16890
rect 10722 16836 10728 16838
rect 10784 16836 10808 16838
rect 10864 16836 10888 16838
rect 10944 16836 10968 16838
rect 11024 16836 11030 16838
rect 10722 16827 11030 16836
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10376 14912 10456 14940
rect 10324 14894 10376 14900
rect 10336 14822 10364 14894
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10428 14618 10456 14758
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10336 14362 10364 14418
rect 10336 14346 10456 14362
rect 10324 14340 10456 14346
rect 10376 14334 10456 14340
rect 10324 14282 10376 14288
rect 10062 14172 10370 14181
rect 10062 14170 10068 14172
rect 10124 14170 10148 14172
rect 10204 14170 10228 14172
rect 10284 14170 10308 14172
rect 10364 14170 10370 14172
rect 10124 14118 10126 14170
rect 10306 14118 10308 14170
rect 10062 14116 10068 14118
rect 10124 14116 10148 14118
rect 10204 14116 10228 14118
rect 10284 14116 10308 14118
rect 10364 14116 10370 14118
rect 10062 14107 10370 14116
rect 10062 13084 10370 13093
rect 10062 13082 10068 13084
rect 10124 13082 10148 13084
rect 10204 13082 10228 13084
rect 10284 13082 10308 13084
rect 10364 13082 10370 13084
rect 10124 13030 10126 13082
rect 10306 13030 10308 13082
rect 10062 13028 10068 13030
rect 10124 13028 10148 13030
rect 10204 13028 10228 13030
rect 10284 13028 10308 13030
rect 10364 13028 10370 13030
rect 10062 13019 10370 13028
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 10428 12866 10456 14334
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 10336 12838 10456 12866
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9404 11212 9456 11218
rect 9324 11172 9404 11200
rect 9404 11154 9456 11160
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9140 9574 9260 9602
rect 9324 9586 9352 10542
rect 9416 10266 9444 11154
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9508 10198 9536 11222
rect 9600 11218 9628 11562
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 9508 9654 9536 10134
rect 9692 10062 9720 12650
rect 10152 12442 10180 12718
rect 10336 12714 10364 12838
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10428 12306 10456 12718
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 9784 11762 9812 12242
rect 10062 11996 10370 12005
rect 10062 11994 10068 11996
rect 10124 11994 10148 11996
rect 10204 11994 10228 11996
rect 10284 11994 10308 11996
rect 10364 11994 10370 11996
rect 10124 11942 10126 11994
rect 10306 11942 10308 11994
rect 10062 11940 10068 11942
rect 10124 11940 10148 11942
rect 10204 11940 10228 11942
rect 10284 11940 10308 11942
rect 10364 11940 10370 11942
rect 10062 11931 10370 11940
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9784 10606 9812 11086
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9784 9722 9812 9998
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9496 9648 9548 9654
rect 9416 9596 9496 9602
rect 9416 9590 9548 9596
rect 9312 9580 9364 9586
rect 9140 8378 9168 9574
rect 9312 9522 9364 9528
rect 9416 9574 9536 9590
rect 9218 9480 9274 9489
rect 9218 9415 9274 9424
rect 9232 9110 9260 9415
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 9416 8566 9444 9574
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9508 9178 9536 9454
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9416 8430 9444 8502
rect 9508 8430 9536 8910
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9600 8634 9628 8774
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9404 8424 9456 8430
rect 9140 8350 9352 8378
rect 9404 8366 9456 8372
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 8022 9168 8230
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 7002 9168 7278
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9232 6866 9260 7346
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9324 6202 9352 8350
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 7818 9444 8230
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9416 6848 9444 7754
rect 9692 7546 9720 7890
rect 9784 7750 9812 9658
rect 9876 7886 9904 11494
rect 10060 11354 10088 11630
rect 10152 11354 10180 11698
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10062 10908 10370 10917
rect 10062 10906 10068 10908
rect 10124 10906 10148 10908
rect 10204 10906 10228 10908
rect 10284 10906 10308 10908
rect 10364 10906 10370 10908
rect 10124 10854 10126 10906
rect 10306 10854 10308 10906
rect 10062 10852 10068 10854
rect 10124 10852 10148 10854
rect 10204 10852 10228 10854
rect 10284 10852 10308 10854
rect 10364 10852 10370 10854
rect 10062 10843 10370 10852
rect 10428 10266 10456 12242
rect 10520 12238 10548 16730
rect 11072 16726 11100 23582
rect 11164 18442 11192 39850
rect 11256 36786 11284 40054
rect 11244 36780 11296 36786
rect 11244 36722 11296 36728
rect 11244 33312 11296 33318
rect 11244 33254 11296 33260
rect 11256 29850 11284 33254
rect 11336 33040 11388 33046
rect 11336 32982 11388 32988
rect 11348 30054 11376 32982
rect 11336 30048 11388 30054
rect 11336 29990 11388 29996
rect 11244 29844 11296 29850
rect 11244 29786 11296 29792
rect 11242 29200 11298 29209
rect 11242 29135 11298 29144
rect 11256 27606 11284 29135
rect 11336 28552 11388 28558
rect 11336 28494 11388 28500
rect 11244 27600 11296 27606
rect 11244 27542 11296 27548
rect 11256 26625 11284 27542
rect 11348 26790 11376 28494
rect 11336 26784 11388 26790
rect 11336 26726 11388 26732
rect 11242 26616 11298 26625
rect 11242 26551 11298 26560
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 11256 24410 11284 26386
rect 11244 24404 11296 24410
rect 11244 24346 11296 24352
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11256 21350 11284 24142
rect 11348 23866 11376 26726
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11348 22574 11376 23462
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 11256 20210 11284 21082
rect 11348 20398 11376 22510
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 11256 20182 11376 20210
rect 11242 19272 11298 19281
rect 11242 19207 11298 19216
rect 11256 18902 11284 19207
rect 11244 18896 11296 18902
rect 11244 18838 11296 18844
rect 11164 18414 11284 18442
rect 11150 18320 11206 18329
rect 11150 18255 11206 18264
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10722 15804 11030 15813
rect 10722 15802 10728 15804
rect 10784 15802 10808 15804
rect 10864 15802 10888 15804
rect 10944 15802 10968 15804
rect 11024 15802 11030 15804
rect 10784 15750 10786 15802
rect 10966 15750 10968 15802
rect 10722 15748 10728 15750
rect 10784 15748 10808 15750
rect 10864 15748 10888 15750
rect 10944 15748 10968 15750
rect 11024 15748 11030 15750
rect 10722 15739 11030 15748
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10612 14822 10640 15302
rect 10704 14958 10732 15574
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14550 10640 14758
rect 10722 14716 11030 14725
rect 10722 14714 10728 14716
rect 10784 14714 10808 14716
rect 10864 14714 10888 14716
rect 10944 14714 10968 14716
rect 11024 14714 11030 14716
rect 10784 14662 10786 14714
rect 10966 14662 10968 14714
rect 10722 14660 10728 14662
rect 10784 14660 10808 14662
rect 10864 14660 10888 14662
rect 10944 14660 10968 14662
rect 11024 14660 11030 14662
rect 10722 14651 11030 14660
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 11072 14482 11100 16458
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10612 13802 10640 14350
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10722 13628 11030 13637
rect 10722 13626 10728 13628
rect 10784 13626 10808 13628
rect 10864 13626 10888 13628
rect 10944 13626 10968 13628
rect 11024 13626 11030 13628
rect 10784 13574 10786 13626
rect 10966 13574 10968 13626
rect 10722 13572 10728 13574
rect 10784 13572 10808 13574
rect 10864 13572 10888 13574
rect 10944 13572 10968 13574
rect 11024 13572 11030 13574
rect 10722 13563 11030 13572
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10612 12374 10640 12718
rect 10722 12540 11030 12549
rect 10722 12538 10728 12540
rect 10784 12538 10808 12540
rect 10864 12538 10888 12540
rect 10944 12538 10968 12540
rect 11024 12538 11030 12540
rect 10784 12486 10786 12538
rect 10966 12486 10968 12538
rect 10722 12484 10728 12486
rect 10784 12484 10808 12486
rect 10864 12484 10888 12486
rect 10944 12484 10968 12486
rect 11024 12484 11030 12486
rect 10722 12475 11030 12484
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11898 10548 12174
rect 10612 12170 10640 12310
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 11072 11694 11100 14418
rect 11164 14346 11192 18255
rect 11256 16561 11284 18414
rect 11348 16658 11376 20182
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11242 16552 11298 16561
rect 11242 16487 11298 16496
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11348 14074 11376 16594
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10612 11150 10640 11630
rect 10722 11452 11030 11461
rect 10722 11450 10728 11452
rect 10784 11450 10808 11452
rect 10864 11450 10888 11452
rect 10944 11450 10968 11452
rect 11024 11450 11030 11452
rect 10784 11398 10786 11450
rect 10966 11398 10968 11450
rect 10722 11396 10728 11398
rect 10784 11396 10808 11398
rect 10864 11396 10888 11398
rect 10944 11396 10968 11398
rect 11024 11396 11030 11398
rect 10722 11387 11030 11396
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10612 10198 10640 10406
rect 10722 10364 11030 10373
rect 10722 10362 10728 10364
rect 10784 10362 10808 10364
rect 10864 10362 10888 10364
rect 10944 10362 10968 10364
rect 11024 10362 11030 10364
rect 10784 10310 10786 10362
rect 10966 10310 10968 10362
rect 10722 10308 10728 10310
rect 10784 10308 10808 10310
rect 10864 10308 10888 10310
rect 10944 10308 10968 10310
rect 11024 10308 11030 10310
rect 10722 10299 11030 10308
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9968 9518 9996 9930
rect 10062 9820 10370 9829
rect 10062 9818 10068 9820
rect 10124 9818 10148 9820
rect 10204 9818 10228 9820
rect 10284 9818 10308 9820
rect 10364 9818 10370 9820
rect 10124 9766 10126 9818
rect 10306 9766 10308 9818
rect 10062 9764 10068 9766
rect 10124 9764 10148 9766
rect 10204 9764 10228 9766
rect 10284 9764 10308 9766
rect 10364 9764 10370 9766
rect 10062 9755 10370 9764
rect 10612 9518 10640 10134
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10062 8732 10370 8741
rect 10062 8730 10068 8732
rect 10124 8730 10148 8732
rect 10204 8730 10228 8732
rect 10284 8730 10308 8732
rect 10364 8730 10370 8732
rect 10124 8678 10126 8730
rect 10306 8678 10308 8730
rect 10062 8676 10068 8678
rect 10124 8676 10148 8678
rect 10204 8676 10228 8678
rect 10284 8676 10308 8678
rect 10364 8676 10370 8678
rect 10062 8667 10370 8676
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10520 8514 10548 9386
rect 10722 9276 11030 9285
rect 10722 9274 10728 9276
rect 10784 9274 10808 9276
rect 10864 9274 10888 9276
rect 10944 9274 10968 9276
rect 11024 9274 11030 9276
rect 10784 9222 10786 9274
rect 10966 9222 10968 9274
rect 10722 9220 10728 9222
rect 10784 9220 10808 9222
rect 10864 9220 10888 9222
rect 10944 9220 10968 9222
rect 11024 9220 11030 9222
rect 10722 9211 11030 9220
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8634 10640 8910
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9876 7342 9904 7822
rect 9968 7342 9996 7822
rect 10060 7818 10088 8366
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10152 8090 10180 8298
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10428 7954 10456 8502
rect 10520 8486 10640 8514
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10062 7644 10370 7653
rect 10062 7642 10068 7644
rect 10124 7642 10148 7644
rect 10204 7642 10228 7644
rect 10284 7642 10308 7644
rect 10364 7642 10370 7644
rect 10124 7590 10126 7642
rect 10306 7590 10308 7642
rect 10062 7588 10068 7590
rect 10124 7588 10148 7590
rect 10204 7588 10228 7590
rect 10284 7588 10308 7590
rect 10364 7588 10370 7590
rect 10062 7579 10370 7588
rect 10520 7342 10548 7686
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 9864 7200 9916 7206
rect 10612 7188 10640 8486
rect 10722 8188 11030 8197
rect 10722 8186 10728 8188
rect 10784 8186 10808 8188
rect 10864 8186 10888 8188
rect 10944 8186 10968 8188
rect 11024 8186 11030 8188
rect 10784 8134 10786 8186
rect 10966 8134 10968 8186
rect 10722 8132 10728 8134
rect 10784 8132 10808 8134
rect 10864 8132 10888 8134
rect 10944 8132 10968 8134
rect 11024 8132 11030 8134
rect 10722 8123 11030 8132
rect 9864 7142 9916 7148
rect 10520 7160 10640 7188
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9496 6860 9548 6866
rect 9416 6820 9496 6848
rect 9496 6802 9548 6808
rect 9140 5914 9168 6190
rect 9324 6174 9536 6202
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5370 9444 5510
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9508 5114 9536 6174
rect 9600 5930 9628 6938
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9600 5902 9720 5930
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9600 5302 9628 5714
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9416 4758 9444 5102
rect 9508 5086 9628 5114
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9232 4078 9260 4558
rect 9324 4282 9352 4626
rect 9508 4622 9536 4966
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9126 3768 9182 3777
rect 9126 3703 9128 3712
rect 9180 3703 9182 3712
rect 9128 3674 9180 3680
rect 9600 3602 9628 5086
rect 9692 4826 9720 5902
rect 9784 5166 9812 6598
rect 9876 5234 9904 7142
rect 10062 6556 10370 6565
rect 10062 6554 10068 6556
rect 10124 6554 10148 6556
rect 10204 6554 10228 6556
rect 10284 6554 10308 6556
rect 10364 6554 10370 6556
rect 10124 6502 10126 6554
rect 10306 6502 10308 6554
rect 10062 6500 10068 6502
rect 10124 6500 10148 6502
rect 10204 6500 10228 6502
rect 10284 6500 10308 6502
rect 10364 6500 10370 6502
rect 10062 6491 10370 6500
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5914 10456 6190
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10048 5772 10100 5778
rect 9968 5732 10048 5760
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9692 3942 9720 4762
rect 9784 4758 9812 5102
rect 9968 4826 9996 5732
rect 10048 5714 10100 5720
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10062 5468 10370 5477
rect 10062 5466 10068 5468
rect 10124 5466 10148 5468
rect 10204 5466 10228 5468
rect 10284 5466 10308 5468
rect 10364 5466 10370 5468
rect 10124 5414 10126 5466
rect 10306 5414 10308 5466
rect 10062 5412 10068 5414
rect 10124 5412 10148 5414
rect 10204 5412 10228 5414
rect 10284 5412 10308 5414
rect 10364 5412 10370 5414
rect 10062 5403 10370 5412
rect 10428 5166 10456 5646
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10428 4826 10456 5102
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9784 4078 9812 4422
rect 10062 4380 10370 4389
rect 10062 4378 10068 4380
rect 10124 4378 10148 4380
rect 10204 4378 10228 4380
rect 10284 4378 10308 4380
rect 10364 4378 10370 4380
rect 10124 4326 10126 4378
rect 10306 4326 10308 4378
rect 10062 4324 10068 4326
rect 10124 4324 10148 4326
rect 10204 4324 10228 4326
rect 10284 4324 10308 4326
rect 10364 4324 10370 4326
rect 10062 4315 10370 4324
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 8312 2310 8340 2586
rect 9048 2582 9076 2994
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8772 2106 8800 2246
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 8760 2100 8812 2106
rect 8760 2042 8812 2048
rect 9140 1902 9168 3334
rect 9600 3210 9628 3538
rect 9600 3194 9720 3210
rect 9600 3188 9732 3194
rect 9600 3182 9680 3188
rect 9680 3130 9732 3136
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9508 2038 9536 2518
rect 9876 2106 9904 4082
rect 10520 3398 10548 7160
rect 10722 7100 11030 7109
rect 10722 7098 10728 7100
rect 10784 7098 10808 7100
rect 10864 7098 10888 7100
rect 10944 7098 10968 7100
rect 11024 7098 11030 7100
rect 10784 7046 10786 7098
rect 10966 7046 10968 7098
rect 10722 7044 10728 7046
rect 10784 7044 10808 7046
rect 10864 7044 10888 7046
rect 10944 7044 10968 7046
rect 11024 7044 11030 7046
rect 10722 7035 11030 7044
rect 10722 6012 11030 6021
rect 10722 6010 10728 6012
rect 10784 6010 10808 6012
rect 10864 6010 10888 6012
rect 10944 6010 10968 6012
rect 11024 6010 11030 6012
rect 10784 5958 10786 6010
rect 10966 5958 10968 6010
rect 10722 5956 10728 5958
rect 10784 5956 10808 5958
rect 10864 5956 10888 5958
rect 10944 5956 10968 5958
rect 11024 5956 11030 5958
rect 10722 5947 11030 5956
rect 10692 5772 10744 5778
rect 10612 5732 10692 5760
rect 10612 4622 10640 5732
rect 10692 5714 10744 5720
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10704 5234 10732 5510
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10722 4924 11030 4933
rect 10722 4922 10728 4924
rect 10784 4922 10808 4924
rect 10864 4922 10888 4924
rect 10944 4922 10968 4924
rect 11024 4922 11030 4924
rect 10784 4870 10786 4922
rect 10966 4870 10968 4922
rect 10722 4868 10728 4870
rect 10784 4868 10808 4870
rect 10864 4868 10888 4870
rect 10944 4868 10968 4870
rect 11024 4868 11030 4870
rect 10722 4859 11030 4868
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10062 3292 10370 3301
rect 10062 3290 10068 3292
rect 10124 3290 10148 3292
rect 10204 3290 10228 3292
rect 10284 3290 10308 3292
rect 10364 3290 10370 3292
rect 10124 3238 10126 3290
rect 10306 3238 10308 3290
rect 10062 3236 10068 3238
rect 10124 3236 10148 3238
rect 10204 3236 10228 3238
rect 10284 3236 10308 3238
rect 10364 3236 10370 3238
rect 10062 3227 10370 3236
rect 10520 2990 10548 3334
rect 10612 3194 10640 3878
rect 10722 3836 11030 3845
rect 10722 3834 10728 3836
rect 10784 3834 10808 3836
rect 10864 3834 10888 3836
rect 10944 3834 10968 3836
rect 11024 3834 11030 3836
rect 10784 3782 10786 3834
rect 10966 3782 10968 3834
rect 10722 3780 10728 3782
rect 10784 3780 10808 3782
rect 10864 3780 10888 3782
rect 10944 3780 10968 3782
rect 11024 3780 11030 3782
rect 10722 3771 11030 3780
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10722 2748 11030 2757
rect 10722 2746 10728 2748
rect 10784 2746 10808 2748
rect 10864 2746 10888 2748
rect 10944 2746 10968 2748
rect 11024 2746 11030 2748
rect 10784 2694 10786 2746
rect 10966 2694 10968 2746
rect 10722 2692 10728 2694
rect 10784 2692 10808 2694
rect 10864 2692 10888 2694
rect 10944 2692 10968 2694
rect 11024 2692 11030 2694
rect 10722 2683 11030 2692
rect 10062 2204 10370 2213
rect 10062 2202 10068 2204
rect 10124 2202 10148 2204
rect 10204 2202 10228 2204
rect 10284 2202 10308 2204
rect 10364 2202 10370 2204
rect 10124 2150 10126 2202
rect 10306 2150 10308 2202
rect 10062 2148 10068 2150
rect 10124 2148 10148 2150
rect 10204 2148 10228 2150
rect 10284 2148 10308 2150
rect 10364 2148 10370 2150
rect 10062 2139 10370 2148
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 9496 2032 9548 2038
rect 9496 1974 9548 1980
rect 7196 1896 7248 1902
rect 7196 1838 7248 1844
rect 7932 1896 7984 1902
rect 7932 1838 7984 1844
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 10722 1660 11030 1669
rect 10722 1658 10728 1660
rect 10784 1658 10808 1660
rect 10864 1658 10888 1660
rect 10944 1658 10968 1660
rect 11024 1658 11030 1660
rect 10784 1606 10786 1658
rect 10966 1606 10968 1658
rect 10722 1604 10728 1606
rect 10784 1604 10808 1606
rect 10864 1604 10888 1606
rect 10944 1604 10968 1606
rect 11024 1604 11030 1606
rect 10722 1595 11030 1604
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 3516 1216 3568 1222
rect 3516 1158 3568 1164
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 10062 1116 10370 1125
rect 10062 1114 10068 1116
rect 10124 1114 10148 1116
rect 10204 1114 10228 1116
rect 10284 1114 10308 1116
rect 10364 1114 10370 1116
rect 10124 1062 10126 1114
rect 10306 1062 10308 1114
rect 10062 1060 10068 1062
rect 10124 1060 10148 1062
rect 10204 1060 10228 1062
rect 10284 1060 10308 1062
rect 10364 1060 10370 1062
rect 10062 1051 10370 1060
rect 3240 1012 3292 1018
rect 3240 954 3292 960
rect 3424 1012 3476 1018
rect 3424 954 3476 960
rect 3056 740 3108 746
rect 3056 682 3108 688
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 10722 572 11030 581
rect 10722 570 10728 572
rect 10784 570 10808 572
rect 10864 570 10888 572
rect 10944 570 10968 572
rect 11024 570 11030 572
rect 10784 518 10786 570
rect 10966 518 10968 570
rect 10722 516 10728 518
rect 10784 516 10808 518
rect 10864 516 10888 518
rect 10944 516 10968 518
rect 11024 516 11030 518
rect 10722 507 11030 516
<< via2 >>
rect 386 41656 442 41712
rect 294 37984 350 38040
rect 202 35128 258 35184
rect 1122 43560 1178 43616
rect 662 41384 718 41440
rect 570 40296 626 40352
rect 1122 41520 1178 41576
rect 846 40568 902 40624
rect 1122 41384 1178 41440
rect 1030 40024 1086 40080
rect 938 39480 994 39536
rect 754 36760 810 36816
rect 662 36216 718 36272
rect 110 26968 166 27024
rect 18 26016 74 26072
rect 294 31728 350 31784
rect 478 31456 534 31512
rect 478 29144 534 29200
rect 110 22208 166 22264
rect 386 28872 442 28928
rect 386 25608 442 25664
rect 386 23432 442 23488
rect 294 19352 350 19408
rect 662 29008 718 29064
rect 662 28600 718 28656
rect 1122 39244 1124 39264
rect 1124 39244 1176 39264
rect 1176 39244 1178 39264
rect 1122 39208 1178 39244
rect 1030 38836 1032 38856
rect 1032 38836 1084 38856
rect 1084 38836 1086 38856
rect 1030 38800 1086 38836
rect 1122 35148 1178 35184
rect 1122 35128 1124 35148
rect 1124 35128 1176 35148
rect 1176 35128 1178 35148
rect 1122 34892 1124 34912
rect 1124 34892 1176 34912
rect 1176 34892 1178 34912
rect 1122 34856 1178 34892
rect 938 34348 940 34368
rect 940 34348 992 34368
rect 992 34348 994 34368
rect 938 34312 994 34348
rect 1122 31456 1178 31512
rect 1122 31320 1178 31376
rect 1030 29552 1086 29608
rect 1030 29416 1086 29472
rect 1306 40432 1362 40488
rect 1306 39752 1362 39808
rect 1306 39480 1362 39536
rect 1490 39616 1546 39672
rect 2134 41112 2190 41168
rect 1858 40432 1914 40488
rect 1858 38528 1914 38584
rect 2226 40432 2282 40488
rect 1858 35128 1914 35184
rect 1950 34720 2006 34776
rect 2042 33088 2098 33144
rect 3668 42458 3724 42460
rect 3748 42458 3804 42460
rect 3828 42458 3884 42460
rect 3908 42458 3964 42460
rect 3668 42406 3714 42458
rect 3714 42406 3724 42458
rect 3748 42406 3778 42458
rect 3778 42406 3790 42458
rect 3790 42406 3804 42458
rect 3828 42406 3842 42458
rect 3842 42406 3854 42458
rect 3854 42406 3884 42458
rect 3908 42406 3918 42458
rect 3918 42406 3964 42458
rect 3668 42404 3724 42406
rect 3748 42404 3804 42406
rect 3828 42404 3884 42406
rect 3908 42404 3964 42406
rect 4328 43002 4384 43004
rect 4408 43002 4464 43004
rect 4488 43002 4544 43004
rect 4568 43002 4624 43004
rect 4328 42950 4374 43002
rect 4374 42950 4384 43002
rect 4408 42950 4438 43002
rect 4438 42950 4450 43002
rect 4450 42950 4464 43002
rect 4488 42950 4502 43002
rect 4502 42950 4514 43002
rect 4514 42950 4544 43002
rect 4568 42950 4578 43002
rect 4578 42950 4624 43002
rect 4328 42948 4384 42950
rect 4408 42948 4464 42950
rect 4488 42948 4544 42950
rect 4568 42948 4624 42950
rect 3054 40840 3110 40896
rect 2962 40160 3018 40216
rect 2594 39616 2650 39672
rect 2318 38528 2374 38584
rect 2318 37304 2374 37360
rect 2042 32816 2098 32872
rect 1766 31592 1822 31648
rect 2778 38936 2834 38992
rect 2870 38392 2926 38448
rect 2962 38004 3018 38040
rect 2962 37984 2964 38004
rect 2964 37984 3016 38004
rect 3016 37984 3018 38004
rect 2870 36352 2926 36408
rect 2778 35944 2834 36000
rect 3668 41370 3724 41372
rect 3748 41370 3804 41372
rect 3828 41370 3884 41372
rect 3908 41370 3964 41372
rect 3668 41318 3714 41370
rect 3714 41318 3724 41370
rect 3748 41318 3778 41370
rect 3778 41318 3790 41370
rect 3790 41318 3804 41370
rect 3828 41318 3842 41370
rect 3842 41318 3854 41370
rect 3854 41318 3884 41370
rect 3908 41318 3918 41370
rect 3918 41318 3964 41370
rect 3668 41316 3724 41318
rect 3748 41316 3804 41318
rect 3828 41316 3884 41318
rect 3908 41316 3964 41318
rect 3668 40282 3724 40284
rect 3748 40282 3804 40284
rect 3828 40282 3884 40284
rect 3908 40282 3964 40284
rect 3668 40230 3714 40282
rect 3714 40230 3724 40282
rect 3748 40230 3778 40282
rect 3778 40230 3790 40282
rect 3790 40230 3804 40282
rect 3828 40230 3842 40282
rect 3842 40230 3854 40282
rect 3854 40230 3884 40282
rect 3908 40230 3918 40282
rect 3918 40230 3964 40282
rect 3668 40228 3724 40230
rect 3748 40228 3804 40230
rect 3828 40228 3884 40230
rect 3908 40228 3964 40230
rect 3238 37712 3294 37768
rect 3606 39888 3662 39944
rect 3668 39194 3724 39196
rect 3748 39194 3804 39196
rect 3828 39194 3884 39196
rect 3908 39194 3964 39196
rect 3668 39142 3714 39194
rect 3714 39142 3724 39194
rect 3748 39142 3778 39194
rect 3778 39142 3790 39194
rect 3790 39142 3804 39194
rect 3828 39142 3842 39194
rect 3842 39142 3854 39194
rect 3854 39142 3884 39194
rect 3908 39142 3918 39194
rect 3918 39142 3964 39194
rect 3668 39140 3724 39142
rect 3748 39140 3804 39142
rect 3828 39140 3884 39142
rect 3908 39140 3964 39142
rect 3790 38412 3846 38448
rect 3790 38392 3792 38412
rect 3792 38392 3844 38412
rect 3844 38392 3846 38412
rect 3606 38256 3662 38312
rect 3668 38106 3724 38108
rect 3748 38106 3804 38108
rect 3828 38106 3884 38108
rect 3908 38106 3964 38108
rect 3668 38054 3714 38106
rect 3714 38054 3724 38106
rect 3748 38054 3778 38106
rect 3778 38054 3790 38106
rect 3790 38054 3804 38106
rect 3828 38054 3842 38106
rect 3842 38054 3854 38106
rect 3854 38054 3884 38106
rect 3908 38054 3918 38106
rect 3918 38054 3964 38106
rect 3668 38052 3724 38054
rect 3748 38052 3804 38054
rect 3828 38052 3884 38054
rect 3908 38052 3964 38054
rect 3606 37848 3662 37904
rect 3668 37018 3724 37020
rect 3748 37018 3804 37020
rect 3828 37018 3884 37020
rect 3908 37018 3964 37020
rect 3668 36966 3714 37018
rect 3714 36966 3724 37018
rect 3748 36966 3778 37018
rect 3778 36966 3790 37018
rect 3790 36966 3804 37018
rect 3828 36966 3842 37018
rect 3842 36966 3854 37018
rect 3854 36966 3884 37018
rect 3908 36966 3918 37018
rect 3918 36966 3964 37018
rect 3668 36964 3724 36966
rect 3748 36964 3804 36966
rect 3828 36964 3884 36966
rect 3908 36964 3964 36966
rect 3790 36760 3846 36816
rect 4342 42064 4398 42120
rect 4328 41914 4384 41916
rect 4408 41914 4464 41916
rect 4488 41914 4544 41916
rect 4568 41914 4624 41916
rect 4328 41862 4374 41914
rect 4374 41862 4384 41914
rect 4408 41862 4438 41914
rect 4438 41862 4450 41914
rect 4450 41862 4464 41914
rect 4488 41862 4502 41914
rect 4502 41862 4514 41914
rect 4514 41862 4544 41914
rect 4568 41862 4578 41914
rect 4578 41862 4624 41914
rect 4328 41860 4384 41862
rect 4408 41860 4464 41862
rect 4488 41860 4544 41862
rect 4568 41860 4624 41862
rect 4328 40826 4384 40828
rect 4408 40826 4464 40828
rect 4488 40826 4544 40828
rect 4568 40826 4624 40828
rect 4328 40774 4374 40826
rect 4374 40774 4384 40826
rect 4408 40774 4438 40826
rect 4438 40774 4450 40826
rect 4450 40774 4464 40826
rect 4488 40774 4502 40826
rect 4502 40774 4514 40826
rect 4514 40774 4544 40826
rect 4568 40774 4578 40826
rect 4578 40774 4624 40826
rect 4328 40772 4384 40774
rect 4408 40772 4464 40774
rect 4488 40772 4544 40774
rect 4568 40772 4624 40774
rect 4328 39738 4384 39740
rect 4408 39738 4464 39740
rect 4488 39738 4544 39740
rect 4568 39738 4624 39740
rect 4328 39686 4374 39738
rect 4374 39686 4384 39738
rect 4408 39686 4438 39738
rect 4438 39686 4450 39738
rect 4450 39686 4464 39738
rect 4488 39686 4502 39738
rect 4502 39686 4514 39738
rect 4514 39686 4544 39738
rect 4568 39686 4578 39738
rect 4578 39686 4624 39738
rect 4328 39684 4384 39686
rect 4408 39684 4464 39686
rect 4488 39684 4544 39686
rect 4568 39684 4624 39686
rect 4328 38650 4384 38652
rect 4408 38650 4464 38652
rect 4488 38650 4544 38652
rect 4568 38650 4624 38652
rect 4328 38598 4374 38650
rect 4374 38598 4384 38650
rect 4408 38598 4438 38650
rect 4438 38598 4450 38650
rect 4450 38598 4464 38650
rect 4488 38598 4502 38650
rect 4502 38598 4514 38650
rect 4514 38598 4544 38650
rect 4568 38598 4578 38650
rect 4578 38598 4624 38650
rect 4328 38596 4384 38598
rect 4408 38596 4464 38598
rect 4488 38596 4544 38598
rect 4568 38596 4624 38598
rect 4894 39480 4950 39536
rect 4434 38120 4490 38176
rect 4328 37562 4384 37564
rect 4408 37562 4464 37564
rect 4488 37562 4544 37564
rect 4568 37562 4624 37564
rect 4328 37510 4374 37562
rect 4374 37510 4384 37562
rect 4408 37510 4438 37562
rect 4438 37510 4450 37562
rect 4450 37510 4464 37562
rect 4488 37510 4502 37562
rect 4502 37510 4514 37562
rect 4514 37510 4544 37562
rect 4568 37510 4578 37562
rect 4578 37510 4624 37562
rect 4328 37508 4384 37510
rect 4408 37508 4464 37510
rect 4488 37508 4544 37510
rect 4568 37508 4624 37510
rect 5262 40024 5318 40080
rect 7746 43560 7802 43616
rect 5814 42200 5870 42256
rect 4986 38800 5042 38856
rect 4328 36474 4384 36476
rect 4408 36474 4464 36476
rect 4488 36474 4544 36476
rect 4568 36474 4624 36476
rect 4328 36422 4374 36474
rect 4374 36422 4384 36474
rect 4408 36422 4438 36474
rect 4438 36422 4450 36474
rect 4450 36422 4464 36474
rect 4488 36422 4502 36474
rect 4502 36422 4514 36474
rect 4514 36422 4544 36474
rect 4568 36422 4578 36474
rect 4578 36422 4624 36474
rect 4328 36420 4384 36422
rect 4408 36420 4464 36422
rect 4488 36420 4544 36422
rect 4568 36420 4624 36422
rect 2686 34856 2742 34912
rect 2962 34992 3018 35048
rect 2686 34584 2742 34640
rect 2778 33224 2834 33280
rect 2502 32952 2558 33008
rect 2410 32272 2466 32328
rect 2318 31864 2374 31920
rect 1766 31084 1768 31104
rect 1768 31084 1820 31104
rect 1820 31084 1822 31104
rect 1766 31048 1822 31084
rect 1214 29588 1216 29608
rect 1216 29588 1268 29608
rect 1268 29588 1270 29608
rect 1214 29552 1270 29588
rect 938 28056 994 28112
rect 938 27920 994 27976
rect 846 27820 848 27840
rect 848 27820 900 27840
rect 900 27820 902 27840
rect 846 27784 902 27820
rect 1122 28056 1178 28112
rect 1306 28736 1362 28792
rect 1306 28464 1362 28520
rect 1214 27512 1270 27568
rect 1122 27104 1178 27160
rect 1030 26832 1086 26888
rect 1398 27784 1454 27840
rect 1398 27512 1454 27568
rect 1030 25744 1086 25800
rect 2042 30504 2098 30560
rect 1950 28756 2006 28792
rect 1950 28736 1952 28756
rect 1952 28736 2004 28756
rect 2004 28736 2006 28756
rect 2318 30912 2374 30968
rect 2226 30232 2282 30288
rect 2318 30096 2374 30152
rect 2134 29280 2190 29336
rect 2134 27920 2190 27976
rect 2134 27648 2190 27704
rect 1950 27512 2006 27568
rect 1582 27412 1584 27432
rect 1584 27412 1636 27432
rect 1636 27412 1638 27432
rect 1582 27376 1638 27412
rect 1582 27240 1638 27296
rect 1582 26560 1638 26616
rect 1674 26444 1730 26480
rect 1674 26424 1676 26444
rect 1676 26424 1728 26444
rect 1728 26424 1730 26444
rect 1398 25900 1454 25936
rect 1674 26152 1730 26208
rect 1398 25880 1400 25900
rect 1400 25880 1452 25900
rect 1452 25880 1454 25900
rect 1030 24248 1086 24304
rect 938 23840 994 23896
rect 846 23160 902 23216
rect 938 22924 940 22944
rect 940 22924 992 22944
rect 992 22924 994 22944
rect 938 22888 994 22924
rect 938 22344 994 22400
rect 662 17992 718 18048
rect 294 17448 350 17504
rect 570 17040 626 17096
rect 386 16632 442 16688
rect 570 12008 626 12064
rect 1398 24656 1454 24712
rect 1306 23976 1362 24032
rect 1398 23432 1454 23488
rect 1214 23024 1270 23080
rect 1306 22480 1362 22536
rect 1122 20576 1178 20632
rect 1398 21528 1454 21584
rect 1306 20712 1362 20768
rect 938 17176 994 17232
rect 938 16088 994 16144
rect 846 15816 902 15872
rect 754 12280 810 12336
rect 662 5480 718 5536
rect 386 5208 442 5264
rect 386 4936 442 4992
rect 386 4392 442 4448
rect 1122 16904 1178 16960
rect 1122 16768 1178 16824
rect 1398 20460 1454 20496
rect 1398 20440 1400 20460
rect 1400 20440 1452 20460
rect 1452 20440 1454 20460
rect 1766 24384 1822 24440
rect 1674 22616 1730 22672
rect 1398 19216 1454 19272
rect 1490 17176 1546 17232
rect 2778 31728 2834 31784
rect 3146 31864 3202 31920
rect 3668 35930 3724 35932
rect 3748 35930 3804 35932
rect 3828 35930 3884 35932
rect 3908 35930 3964 35932
rect 3668 35878 3714 35930
rect 3714 35878 3724 35930
rect 3748 35878 3778 35930
rect 3778 35878 3790 35930
rect 3790 35878 3804 35930
rect 3828 35878 3842 35930
rect 3842 35878 3854 35930
rect 3854 35878 3884 35930
rect 3908 35878 3918 35930
rect 3918 35878 3964 35930
rect 3668 35876 3724 35878
rect 3748 35876 3804 35878
rect 3828 35876 3884 35878
rect 3908 35876 3964 35878
rect 4066 35808 4122 35864
rect 3974 35148 4030 35184
rect 3974 35128 3976 35148
rect 3976 35128 4028 35148
rect 4028 35128 4030 35148
rect 3668 34842 3724 34844
rect 3748 34842 3804 34844
rect 3828 34842 3884 34844
rect 3908 34842 3964 34844
rect 3668 34790 3714 34842
rect 3714 34790 3724 34842
rect 3748 34790 3778 34842
rect 3778 34790 3790 34842
rect 3790 34790 3804 34842
rect 3828 34790 3842 34842
rect 3842 34790 3854 34842
rect 3854 34790 3884 34842
rect 3908 34790 3918 34842
rect 3918 34790 3964 34842
rect 3668 34788 3724 34790
rect 3748 34788 3804 34790
rect 3828 34788 3884 34790
rect 3908 34788 3964 34790
rect 4066 34720 4122 34776
rect 3974 34604 4030 34640
rect 3974 34584 3976 34604
rect 3976 34584 4028 34604
rect 4028 34584 4030 34604
rect 3790 34484 3792 34504
rect 3792 34484 3844 34504
rect 3844 34484 3846 34504
rect 3790 34448 3846 34484
rect 3668 33754 3724 33756
rect 3748 33754 3804 33756
rect 3828 33754 3884 33756
rect 3908 33754 3964 33756
rect 3668 33702 3714 33754
rect 3714 33702 3724 33754
rect 3748 33702 3778 33754
rect 3778 33702 3790 33754
rect 3790 33702 3804 33754
rect 3828 33702 3842 33754
rect 3842 33702 3854 33754
rect 3854 33702 3884 33754
rect 3908 33702 3918 33754
rect 3918 33702 3964 33754
rect 3668 33700 3724 33702
rect 3748 33700 3804 33702
rect 3828 33700 3884 33702
rect 3908 33700 3964 33702
rect 2962 30540 2964 30560
rect 2964 30540 3016 30560
rect 3016 30540 3018 30560
rect 2962 30504 3018 30540
rect 3330 31864 3386 31920
rect 3330 31728 3386 31784
rect 3974 33260 3976 33280
rect 3976 33260 4028 33280
rect 4028 33260 4030 33280
rect 3974 33224 4030 33260
rect 3698 32972 3754 33008
rect 3698 32952 3700 32972
rect 3700 32952 3752 32972
rect 3752 32952 3754 32972
rect 3668 32666 3724 32668
rect 3748 32666 3804 32668
rect 3828 32666 3884 32668
rect 3908 32666 3964 32668
rect 3668 32614 3714 32666
rect 3714 32614 3724 32666
rect 3748 32614 3778 32666
rect 3778 32614 3790 32666
rect 3790 32614 3804 32666
rect 3828 32614 3842 32666
rect 3842 32614 3854 32666
rect 3854 32614 3884 32666
rect 3908 32614 3918 32666
rect 3918 32614 3964 32666
rect 3668 32612 3724 32614
rect 3748 32612 3804 32614
rect 3828 32612 3884 32614
rect 3908 32612 3964 32614
rect 3606 31728 3662 31784
rect 3668 31578 3724 31580
rect 3748 31578 3804 31580
rect 3828 31578 3884 31580
rect 3908 31578 3964 31580
rect 3668 31526 3714 31578
rect 3714 31526 3724 31578
rect 3748 31526 3778 31578
rect 3778 31526 3790 31578
rect 3790 31526 3804 31578
rect 3828 31526 3842 31578
rect 3842 31526 3854 31578
rect 3854 31526 3884 31578
rect 3908 31526 3918 31578
rect 3918 31526 3964 31578
rect 3668 31524 3724 31526
rect 3748 31524 3804 31526
rect 3828 31524 3884 31526
rect 3908 31524 3964 31526
rect 3514 31048 3570 31104
rect 3422 30912 3478 30968
rect 3514 30812 3516 30832
rect 3516 30812 3568 30832
rect 3568 30812 3570 30832
rect 3330 30640 3386 30696
rect 3514 30776 3570 30812
rect 2502 28736 2558 28792
rect 2410 26988 2466 27024
rect 2410 26968 2412 26988
rect 2412 26968 2464 26988
rect 2464 26968 2466 26988
rect 2870 29708 2926 29744
rect 2870 29688 2872 29708
rect 2872 29688 2924 29708
rect 2924 29688 2926 29708
rect 3146 29688 3202 29744
rect 2870 29144 2926 29200
rect 2870 28908 2872 28928
rect 2872 28908 2924 28928
rect 2924 28908 2926 28928
rect 2870 28872 2926 28908
rect 2778 28600 2834 28656
rect 2686 28464 2742 28520
rect 2594 28192 2650 28248
rect 2870 28192 2926 28248
rect 2594 27920 2650 27976
rect 2686 27648 2742 27704
rect 2870 27784 2926 27840
rect 2686 27240 2742 27296
rect 2594 26988 2650 27024
rect 2594 26968 2596 26988
rect 2596 26968 2648 26988
rect 2648 26968 2650 26988
rect 2502 26288 2558 26344
rect 2410 26152 2466 26208
rect 2318 26036 2374 26072
rect 2318 26016 2320 26036
rect 2320 26016 2372 26036
rect 2372 26016 2374 26036
rect 2226 25880 2282 25936
rect 2042 24520 2098 24576
rect 2042 24384 2098 24440
rect 2686 26424 2742 26480
rect 2594 25472 2650 25528
rect 2410 25064 2466 25120
rect 2318 24928 2374 24984
rect 2410 24792 2466 24848
rect 2594 24268 2650 24304
rect 2594 24248 2596 24268
rect 2596 24248 2648 24268
rect 2648 24248 2650 24268
rect 2502 23568 2558 23624
rect 2226 23180 2282 23216
rect 2226 23160 2228 23180
rect 2228 23160 2280 23180
rect 2280 23160 2282 23180
rect 2226 22344 2282 22400
rect 2502 22380 2504 22400
rect 2504 22380 2556 22400
rect 2556 22380 2558 22400
rect 2502 22344 2558 22380
rect 2502 22208 2558 22264
rect 2778 25372 2780 25392
rect 2780 25372 2832 25392
rect 2832 25372 2834 25392
rect 2778 25336 2834 25372
rect 2778 23704 2834 23760
rect 3054 27104 3110 27160
rect 3054 26152 3110 26208
rect 2962 25880 3018 25936
rect 3054 24132 3110 24168
rect 3054 24112 3056 24132
rect 3056 24112 3108 24132
rect 3108 24112 3110 24132
rect 2594 21664 2650 21720
rect 2134 20576 2190 20632
rect 3054 23432 3110 23488
rect 3054 22344 3110 22400
rect 1858 17856 1914 17912
rect 1214 12552 1270 12608
rect 1766 14728 1822 14784
rect 1674 13776 1730 13832
rect 2778 20340 2780 20360
rect 2780 20340 2832 20360
rect 2832 20340 2834 20360
rect 2778 20304 2834 20340
rect 3054 21936 3110 21992
rect 3054 21664 3110 21720
rect 3238 27104 3294 27160
rect 4328 35386 4384 35388
rect 4408 35386 4464 35388
rect 4488 35386 4544 35388
rect 4568 35386 4624 35388
rect 4328 35334 4374 35386
rect 4374 35334 4384 35386
rect 4408 35334 4438 35386
rect 4438 35334 4450 35386
rect 4450 35334 4464 35386
rect 4488 35334 4502 35386
rect 4502 35334 4514 35386
rect 4514 35334 4544 35386
rect 4568 35334 4578 35386
rect 4578 35334 4624 35386
rect 4328 35332 4384 35334
rect 4408 35332 4464 35334
rect 4488 35332 4544 35334
rect 4568 35332 4624 35334
rect 4618 34992 4674 35048
rect 5170 38664 5226 38720
rect 6182 40024 6238 40080
rect 6274 39888 6330 39944
rect 5998 39752 6054 39808
rect 5722 38528 5778 38584
rect 5446 36760 5502 36816
rect 5078 34856 5134 34912
rect 4328 34298 4384 34300
rect 4408 34298 4464 34300
rect 4488 34298 4544 34300
rect 4568 34298 4624 34300
rect 4328 34246 4374 34298
rect 4374 34246 4384 34298
rect 4408 34246 4438 34298
rect 4438 34246 4450 34298
rect 4450 34246 4464 34298
rect 4488 34246 4502 34298
rect 4502 34246 4514 34298
rect 4514 34246 4544 34298
rect 4568 34246 4578 34298
rect 4578 34246 4624 34298
rect 4328 34244 4384 34246
rect 4408 34244 4464 34246
rect 4488 34244 4544 34246
rect 4568 34244 4624 34246
rect 5170 34740 5226 34776
rect 5170 34720 5172 34740
rect 5172 34720 5224 34740
rect 5224 34720 5226 34740
rect 5170 34448 5226 34504
rect 5814 36760 5870 36816
rect 5814 36216 5870 36272
rect 5814 35536 5870 35592
rect 5906 34720 5962 34776
rect 5354 34312 5410 34368
rect 5538 33496 5594 33552
rect 6642 41692 6644 41712
rect 6644 41692 6696 41712
rect 6696 41692 6698 41712
rect 6642 41656 6698 41692
rect 6642 40024 6698 40080
rect 7746 41520 7802 41576
rect 7562 41384 7618 41440
rect 7470 41248 7526 41304
rect 6826 39344 6882 39400
rect 7286 38936 7342 38992
rect 6918 38292 6920 38312
rect 6920 38292 6972 38312
rect 6972 38292 6974 38312
rect 6918 38256 6974 38292
rect 6826 37576 6882 37632
rect 6734 37304 6790 37360
rect 6734 35672 6790 35728
rect 6642 34584 6698 34640
rect 4328 33210 4384 33212
rect 4408 33210 4464 33212
rect 4488 33210 4544 33212
rect 4568 33210 4624 33212
rect 4328 33158 4374 33210
rect 4374 33158 4384 33210
rect 4408 33158 4438 33210
rect 4438 33158 4450 33210
rect 4450 33158 4464 33210
rect 4488 33158 4502 33210
rect 4502 33158 4514 33210
rect 4514 33158 4544 33210
rect 4568 33158 4578 33210
rect 4578 33158 4624 33210
rect 4328 33156 4384 33158
rect 4408 33156 4464 33158
rect 4488 33156 4544 33158
rect 4568 33156 4624 33158
rect 4434 32952 4490 33008
rect 4894 32816 4950 32872
rect 4328 32122 4384 32124
rect 4408 32122 4464 32124
rect 4488 32122 4544 32124
rect 4568 32122 4624 32124
rect 4328 32070 4374 32122
rect 4374 32070 4384 32122
rect 4408 32070 4438 32122
rect 4438 32070 4450 32122
rect 4450 32070 4464 32122
rect 4488 32070 4502 32122
rect 4502 32070 4514 32122
rect 4514 32070 4544 32122
rect 4568 32070 4578 32122
rect 4578 32070 4624 32122
rect 4328 32068 4384 32070
rect 4408 32068 4464 32070
rect 4488 32068 4544 32070
rect 4568 32068 4624 32070
rect 4434 31884 4490 31920
rect 4434 31864 4436 31884
rect 4436 31864 4488 31884
rect 4488 31864 4490 31884
rect 4710 31728 4766 31784
rect 4328 31034 4384 31036
rect 4408 31034 4464 31036
rect 4488 31034 4544 31036
rect 4568 31034 4624 31036
rect 4328 30982 4374 31034
rect 4374 30982 4384 31034
rect 4408 30982 4438 31034
rect 4438 30982 4450 31034
rect 4450 30982 4464 31034
rect 4488 30982 4502 31034
rect 4502 30982 4514 31034
rect 4514 30982 4544 31034
rect 4568 30982 4578 31034
rect 4578 30982 4624 31034
rect 4328 30980 4384 30982
rect 4408 30980 4464 30982
rect 4488 30980 4544 30982
rect 4568 30980 4624 30982
rect 3668 30490 3724 30492
rect 3748 30490 3804 30492
rect 3828 30490 3884 30492
rect 3908 30490 3964 30492
rect 3668 30438 3714 30490
rect 3714 30438 3724 30490
rect 3748 30438 3778 30490
rect 3778 30438 3790 30490
rect 3790 30438 3804 30490
rect 3828 30438 3842 30490
rect 3842 30438 3854 30490
rect 3854 30438 3884 30490
rect 3908 30438 3918 30490
rect 3918 30438 3964 30490
rect 3668 30436 3724 30438
rect 3748 30436 3804 30438
rect 3828 30436 3884 30438
rect 3908 30436 3964 30438
rect 3882 29688 3938 29744
rect 3668 29402 3724 29404
rect 3748 29402 3804 29404
rect 3828 29402 3884 29404
rect 3908 29402 3964 29404
rect 3668 29350 3714 29402
rect 3714 29350 3724 29402
rect 3748 29350 3778 29402
rect 3778 29350 3790 29402
rect 3790 29350 3804 29402
rect 3828 29350 3842 29402
rect 3842 29350 3854 29402
rect 3854 29350 3884 29402
rect 3908 29350 3918 29402
rect 3918 29350 3964 29402
rect 3668 29348 3724 29350
rect 3748 29348 3804 29350
rect 3828 29348 3884 29350
rect 3908 29348 3964 29350
rect 3606 29144 3662 29200
rect 3974 29144 4030 29200
rect 3606 28872 3662 28928
rect 3606 28464 3662 28520
rect 3974 28464 4030 28520
rect 3668 28314 3724 28316
rect 3748 28314 3804 28316
rect 3828 28314 3884 28316
rect 3908 28314 3964 28316
rect 3668 28262 3714 28314
rect 3714 28262 3724 28314
rect 3748 28262 3778 28314
rect 3778 28262 3790 28314
rect 3790 28262 3804 28314
rect 3828 28262 3842 28314
rect 3842 28262 3854 28314
rect 3854 28262 3884 28314
rect 3908 28262 3918 28314
rect 3918 28262 3964 28314
rect 3668 28260 3724 28262
rect 3748 28260 3804 28262
rect 3828 28260 3884 28262
rect 3908 28260 3964 28262
rect 3698 27648 3754 27704
rect 3882 27784 3938 27840
rect 4894 31728 4950 31784
rect 4986 30912 5042 30968
rect 4802 30368 4858 30424
rect 5538 32816 5594 32872
rect 5446 32408 5502 32464
rect 5170 31864 5226 31920
rect 4328 29946 4384 29948
rect 4408 29946 4464 29948
rect 4488 29946 4544 29948
rect 4568 29946 4624 29948
rect 4328 29894 4374 29946
rect 4374 29894 4384 29946
rect 4408 29894 4438 29946
rect 4438 29894 4450 29946
rect 4450 29894 4464 29946
rect 4488 29894 4502 29946
rect 4502 29894 4514 29946
rect 4514 29894 4544 29946
rect 4568 29894 4578 29946
rect 4578 29894 4624 29946
rect 4328 29892 4384 29894
rect 4408 29892 4464 29894
rect 4488 29892 4544 29894
rect 4568 29892 4624 29894
rect 4710 29688 4766 29744
rect 4618 29180 4620 29200
rect 4620 29180 4672 29200
rect 4672 29180 4674 29200
rect 4618 29144 4674 29180
rect 4328 28858 4384 28860
rect 4408 28858 4464 28860
rect 4488 28858 4544 28860
rect 4568 28858 4624 28860
rect 4328 28806 4374 28858
rect 4374 28806 4384 28858
rect 4408 28806 4438 28858
rect 4438 28806 4450 28858
rect 4450 28806 4464 28858
rect 4488 28806 4502 28858
rect 4502 28806 4514 28858
rect 4514 28806 4544 28858
rect 4568 28806 4578 28858
rect 4578 28806 4624 28858
rect 4328 28804 4384 28806
rect 4408 28804 4464 28806
rect 4488 28804 4544 28806
rect 4568 28804 4624 28806
rect 5262 31456 5318 31512
rect 6366 33904 6422 33960
rect 5906 32716 5908 32736
rect 5908 32716 5960 32736
rect 5960 32716 5962 32736
rect 5906 32680 5962 32716
rect 5906 32272 5962 32328
rect 5906 32000 5962 32056
rect 8022 41520 8078 41576
rect 10728 43002 10784 43004
rect 10808 43002 10864 43004
rect 10888 43002 10944 43004
rect 10968 43002 11024 43004
rect 10728 42950 10774 43002
rect 10774 42950 10784 43002
rect 10808 42950 10838 43002
rect 10838 42950 10850 43002
rect 10850 42950 10864 43002
rect 10888 42950 10902 43002
rect 10902 42950 10914 43002
rect 10914 42950 10944 43002
rect 10968 42950 10978 43002
rect 10978 42950 11024 43002
rect 10728 42948 10784 42950
rect 10808 42948 10864 42950
rect 10888 42948 10944 42950
rect 10968 42948 11024 42950
rect 8390 41248 8446 41304
rect 8298 41112 8354 41168
rect 8298 40704 8354 40760
rect 7654 39072 7710 39128
rect 7562 38936 7618 38992
rect 7470 38392 7526 38448
rect 7378 38256 7434 38312
rect 7194 36488 7250 36544
rect 7838 38528 7894 38584
rect 7654 38392 7710 38448
rect 7838 38392 7894 38448
rect 7746 38120 7802 38176
rect 7746 37712 7802 37768
rect 8758 41540 8814 41576
rect 8758 41520 8760 41540
rect 8760 41520 8812 41540
rect 8812 41520 8814 41540
rect 8758 41248 8814 41304
rect 8666 40588 8722 40624
rect 8666 40568 8668 40588
rect 8668 40568 8720 40588
rect 8720 40568 8722 40588
rect 8758 40160 8814 40216
rect 10068 42458 10124 42460
rect 10148 42458 10204 42460
rect 10228 42458 10284 42460
rect 10308 42458 10364 42460
rect 10068 42406 10114 42458
rect 10114 42406 10124 42458
rect 10148 42406 10178 42458
rect 10178 42406 10190 42458
rect 10190 42406 10204 42458
rect 10228 42406 10242 42458
rect 10242 42406 10254 42458
rect 10254 42406 10284 42458
rect 10308 42406 10318 42458
rect 10318 42406 10364 42458
rect 10068 42404 10124 42406
rect 10148 42404 10204 42406
rect 10228 42404 10284 42406
rect 10308 42404 10364 42406
rect 8758 40024 8814 40080
rect 8114 39888 8170 39944
rect 7470 37168 7526 37224
rect 7378 35808 7434 35864
rect 6734 33108 6790 33144
rect 7194 33904 7250 33960
rect 6734 33088 6736 33108
rect 6736 33088 6788 33108
rect 6788 33088 6790 33108
rect 6274 32680 6330 32736
rect 6182 32544 6238 32600
rect 6090 32000 6146 32056
rect 6090 31900 6092 31920
rect 6092 31900 6144 31920
rect 6144 31900 6146 31920
rect 6090 31864 6146 31900
rect 5906 31476 5962 31512
rect 5906 31456 5908 31476
rect 5908 31456 5960 31476
rect 5960 31456 5962 31476
rect 5814 30912 5870 30968
rect 5906 30640 5962 30696
rect 5906 30504 5962 30560
rect 5814 30388 5870 30424
rect 5814 30368 5816 30388
rect 5816 30368 5868 30388
rect 5868 30368 5870 30388
rect 4986 28872 5042 28928
rect 4986 28736 5042 28792
rect 4802 28076 4858 28112
rect 4802 28056 4804 28076
rect 4804 28056 4856 28076
rect 4856 28056 4858 28076
rect 4986 28056 5042 28112
rect 4618 27920 4674 27976
rect 4328 27770 4384 27772
rect 4408 27770 4464 27772
rect 4488 27770 4544 27772
rect 4568 27770 4624 27772
rect 4328 27718 4374 27770
rect 4374 27718 4384 27770
rect 4408 27718 4438 27770
rect 4438 27718 4450 27770
rect 4450 27718 4464 27770
rect 4488 27718 4502 27770
rect 4502 27718 4514 27770
rect 4514 27718 4544 27770
rect 4568 27718 4578 27770
rect 4578 27718 4624 27770
rect 4328 27716 4384 27718
rect 4408 27716 4464 27718
rect 4488 27716 4544 27718
rect 4568 27716 4624 27718
rect 4526 27512 4582 27568
rect 3514 27412 3516 27432
rect 3516 27412 3568 27432
rect 3568 27412 3570 27432
rect 3514 27376 3570 27412
rect 3668 27226 3724 27228
rect 3748 27226 3804 27228
rect 3828 27226 3884 27228
rect 3908 27226 3964 27228
rect 3668 27174 3714 27226
rect 3714 27174 3724 27226
rect 3748 27174 3778 27226
rect 3778 27174 3790 27226
rect 3790 27174 3804 27226
rect 3828 27174 3842 27226
rect 3842 27174 3854 27226
rect 3854 27174 3884 27226
rect 3908 27174 3918 27226
rect 3918 27174 3964 27226
rect 3668 27172 3724 27174
rect 3748 27172 3804 27174
rect 3828 27172 3884 27174
rect 3908 27172 3964 27174
rect 3330 26968 3386 27024
rect 3330 26424 3386 26480
rect 3146 21428 3148 21448
rect 3148 21428 3200 21448
rect 3200 21428 3202 21448
rect 3146 21392 3202 21428
rect 4066 26696 4122 26752
rect 3790 26560 3846 26616
rect 4342 27104 4398 27160
rect 4158 26560 4214 26616
rect 3974 26424 4030 26480
rect 3668 26138 3724 26140
rect 3748 26138 3804 26140
rect 3828 26138 3884 26140
rect 3908 26138 3964 26140
rect 3668 26086 3714 26138
rect 3714 26086 3724 26138
rect 3748 26086 3778 26138
rect 3778 26086 3790 26138
rect 3790 26086 3804 26138
rect 3828 26086 3842 26138
rect 3842 26086 3854 26138
rect 3854 26086 3884 26138
rect 3908 26086 3918 26138
rect 3918 26086 3964 26138
rect 3668 26084 3724 26086
rect 3748 26084 3804 26086
rect 3828 26084 3884 26086
rect 3908 26084 3964 26086
rect 3514 25880 3570 25936
rect 3698 25880 3754 25936
rect 3974 25880 4030 25936
rect 3606 25744 3662 25800
rect 3698 25608 3754 25664
rect 3790 25336 3846 25392
rect 4618 27240 4674 27296
rect 4342 26868 4344 26888
rect 4344 26868 4396 26888
rect 4396 26868 4398 26888
rect 4342 26832 4398 26868
rect 4328 26682 4384 26684
rect 4408 26682 4464 26684
rect 4488 26682 4544 26684
rect 4568 26682 4624 26684
rect 4328 26630 4374 26682
rect 4374 26630 4384 26682
rect 4408 26630 4438 26682
rect 4438 26630 4450 26682
rect 4450 26630 4464 26682
rect 4488 26630 4502 26682
rect 4502 26630 4514 26682
rect 4514 26630 4544 26682
rect 4568 26630 4578 26682
rect 4578 26630 4624 26682
rect 4328 26628 4384 26630
rect 4408 26628 4464 26630
rect 4488 26628 4544 26630
rect 4568 26628 4624 26630
rect 4434 26424 4490 26480
rect 3698 25236 3700 25256
rect 3700 25236 3752 25256
rect 3752 25236 3754 25256
rect 3698 25200 3754 25236
rect 3882 25200 3938 25256
rect 3668 25050 3724 25052
rect 3748 25050 3804 25052
rect 3828 25050 3884 25052
rect 3908 25050 3964 25052
rect 3668 24998 3714 25050
rect 3714 24998 3724 25050
rect 3748 24998 3778 25050
rect 3778 24998 3790 25050
rect 3790 24998 3804 25050
rect 3828 24998 3842 25050
rect 3842 24998 3854 25050
rect 3854 24998 3884 25050
rect 3908 24998 3918 25050
rect 3918 24998 3964 25050
rect 3668 24996 3724 24998
rect 3748 24996 3804 24998
rect 3828 24996 3884 24998
rect 3908 24996 3964 24998
rect 3698 24248 3754 24304
rect 3882 24248 3938 24304
rect 4526 26152 4582 26208
rect 4618 26016 4674 26072
rect 4894 26696 4950 26752
rect 5078 26288 5134 26344
rect 4986 26016 5042 26072
rect 4158 25608 4214 25664
rect 4328 25594 4384 25596
rect 4408 25594 4464 25596
rect 4488 25594 4544 25596
rect 4568 25594 4624 25596
rect 4328 25542 4374 25594
rect 4374 25542 4384 25594
rect 4408 25542 4438 25594
rect 4438 25542 4450 25594
rect 4450 25542 4464 25594
rect 4488 25542 4502 25594
rect 4502 25542 4514 25594
rect 4514 25542 4544 25594
rect 4568 25542 4578 25594
rect 4578 25542 4624 25594
rect 4328 25540 4384 25542
rect 4408 25540 4464 25542
rect 4488 25540 4544 25542
rect 4568 25540 4624 25542
rect 4710 25472 4766 25528
rect 3668 23962 3724 23964
rect 3748 23962 3804 23964
rect 3828 23962 3884 23964
rect 3908 23962 3964 23964
rect 3668 23910 3714 23962
rect 3714 23910 3724 23962
rect 3748 23910 3778 23962
rect 3778 23910 3790 23962
rect 3790 23910 3804 23962
rect 3828 23910 3842 23962
rect 3842 23910 3854 23962
rect 3854 23910 3884 23962
rect 3908 23910 3918 23962
rect 3918 23910 3964 23962
rect 3668 23908 3724 23910
rect 3748 23908 3804 23910
rect 3828 23908 3884 23910
rect 3908 23908 3964 23910
rect 3606 23604 3608 23624
rect 3608 23604 3660 23624
rect 3660 23604 3662 23624
rect 3606 23568 3662 23604
rect 3668 22874 3724 22876
rect 3748 22874 3804 22876
rect 3828 22874 3884 22876
rect 3908 22874 3964 22876
rect 3668 22822 3714 22874
rect 3714 22822 3724 22874
rect 3748 22822 3778 22874
rect 3778 22822 3790 22874
rect 3790 22822 3804 22874
rect 3828 22822 3842 22874
rect 3842 22822 3854 22874
rect 3854 22822 3884 22874
rect 3908 22822 3918 22874
rect 3918 22822 3964 22874
rect 3668 22820 3724 22822
rect 3748 22820 3804 22822
rect 3828 22820 3884 22822
rect 3908 22820 3964 22822
rect 4986 25472 5042 25528
rect 4894 25236 4896 25256
rect 4896 25236 4948 25256
rect 4948 25236 4950 25256
rect 4894 25200 4950 25236
rect 4986 25100 4988 25120
rect 4988 25100 5040 25120
rect 5040 25100 5042 25120
rect 4986 25064 5042 25100
rect 4894 24928 4950 24984
rect 4328 24506 4384 24508
rect 4408 24506 4464 24508
rect 4488 24506 4544 24508
rect 4568 24506 4624 24508
rect 4328 24454 4374 24506
rect 4374 24454 4384 24506
rect 4408 24454 4438 24506
rect 4438 24454 4450 24506
rect 4450 24454 4464 24506
rect 4488 24454 4502 24506
rect 4502 24454 4514 24506
rect 4514 24454 4544 24506
rect 4568 24454 4578 24506
rect 4578 24454 4624 24506
rect 4328 24452 4384 24454
rect 4408 24452 4464 24454
rect 4488 24452 4544 24454
rect 4568 24452 4624 24454
rect 4328 23418 4384 23420
rect 4408 23418 4464 23420
rect 4488 23418 4544 23420
rect 4568 23418 4624 23420
rect 4328 23366 4374 23418
rect 4374 23366 4384 23418
rect 4408 23366 4438 23418
rect 4438 23366 4450 23418
rect 4450 23366 4464 23418
rect 4488 23366 4502 23418
rect 4502 23366 4514 23418
rect 4514 23366 4544 23418
rect 4568 23366 4578 23418
rect 4578 23366 4624 23418
rect 4328 23364 4384 23366
rect 4408 23364 4464 23366
rect 4488 23364 4544 23366
rect 4568 23364 4624 23366
rect 4434 23160 4490 23216
rect 4802 23976 4858 24032
rect 4250 22752 4306 22808
rect 3790 22616 3846 22672
rect 3882 22344 3938 22400
rect 4158 22108 4160 22128
rect 4160 22108 4212 22128
rect 4212 22108 4214 22128
rect 4158 22072 4214 22108
rect 4328 22330 4384 22332
rect 4408 22330 4464 22332
rect 4488 22330 4544 22332
rect 4568 22330 4624 22332
rect 4328 22278 4374 22330
rect 4374 22278 4384 22330
rect 4408 22278 4438 22330
rect 4438 22278 4450 22330
rect 4450 22278 4464 22330
rect 4488 22278 4502 22330
rect 4502 22278 4514 22330
rect 4514 22278 4544 22330
rect 4568 22278 4578 22330
rect 4578 22278 4624 22330
rect 4328 22276 4384 22278
rect 4408 22276 4464 22278
rect 4488 22276 4544 22278
rect 4568 22276 4624 22278
rect 4710 22228 4766 22264
rect 4710 22208 4712 22228
rect 4712 22208 4764 22228
rect 4764 22208 4766 22228
rect 4434 22072 4490 22128
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 3238 21256 3294 21312
rect 3330 21120 3386 21176
rect 2778 19916 2834 19952
rect 2778 19896 2780 19916
rect 2780 19896 2832 19916
rect 2832 19896 2834 19916
rect 2410 17992 2466 18048
rect 3146 20868 3202 20904
rect 3146 20848 3148 20868
rect 3148 20848 3200 20868
rect 3200 20848 3202 20868
rect 3330 20712 3386 20768
rect 3330 20576 3386 20632
rect 4066 21528 4122 21584
rect 4066 21256 4122 21312
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 3238 19796 3240 19816
rect 3240 19796 3292 19816
rect 3292 19796 3294 19816
rect 3238 19760 3294 19796
rect 3238 19372 3294 19408
rect 4066 20440 4122 20496
rect 4342 21800 4398 21856
rect 4342 21684 4398 21720
rect 4342 21664 4344 21684
rect 4344 21664 4396 21684
rect 4396 21664 4398 21684
rect 4342 21528 4398 21584
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 5078 24384 5134 24440
rect 5078 22752 5134 22808
rect 5262 29280 5318 29336
rect 5630 29844 5686 29880
rect 5630 29824 5632 29844
rect 5632 29824 5684 29844
rect 5684 29824 5686 29844
rect 5722 29552 5778 29608
rect 5446 28620 5502 28656
rect 5446 28600 5448 28620
rect 5448 28600 5500 28620
rect 5500 28600 5502 28620
rect 5538 28464 5594 28520
rect 5354 26016 5410 26072
rect 5262 25880 5318 25936
rect 5354 25064 5410 25120
rect 5630 27648 5686 27704
rect 5906 29280 5962 29336
rect 5814 28908 5816 28928
rect 5816 28908 5868 28928
rect 5868 28908 5870 28928
rect 5814 28872 5870 28908
rect 5538 25200 5594 25256
rect 5262 24520 5318 24576
rect 5446 24520 5502 24576
rect 6182 31320 6238 31376
rect 7378 33632 7434 33688
rect 7378 33224 7434 33280
rect 7470 33088 7526 33144
rect 8390 39092 8446 39128
rect 8390 39072 8392 39092
rect 8392 39072 8444 39092
rect 8444 39072 8446 39092
rect 8298 38936 8354 38992
rect 8114 38256 8170 38312
rect 8390 38412 8446 38448
rect 8390 38392 8392 38412
rect 8392 38392 8444 38412
rect 8444 38392 8446 38412
rect 8758 39752 8814 39808
rect 8666 39616 8722 39672
rect 8574 38528 8630 38584
rect 8482 38256 8538 38312
rect 8758 38256 8814 38312
rect 8482 38120 8538 38176
rect 8390 37848 8446 37904
rect 9494 40568 9550 40624
rect 10068 41370 10124 41372
rect 10148 41370 10204 41372
rect 10228 41370 10284 41372
rect 10308 41370 10364 41372
rect 10068 41318 10114 41370
rect 10114 41318 10124 41370
rect 10148 41318 10178 41370
rect 10178 41318 10190 41370
rect 10190 41318 10204 41370
rect 10228 41318 10242 41370
rect 10242 41318 10254 41370
rect 10254 41318 10284 41370
rect 10308 41318 10318 41370
rect 10318 41318 10364 41370
rect 10068 41316 10124 41318
rect 10148 41316 10204 41318
rect 10228 41316 10284 41318
rect 10308 41316 10364 41318
rect 10068 40282 10124 40284
rect 10148 40282 10204 40284
rect 10228 40282 10284 40284
rect 10308 40282 10364 40284
rect 10068 40230 10114 40282
rect 10114 40230 10124 40282
rect 10148 40230 10178 40282
rect 10178 40230 10190 40282
rect 10190 40230 10204 40282
rect 10228 40230 10242 40282
rect 10242 40230 10254 40282
rect 10254 40230 10284 40282
rect 10308 40230 10318 40282
rect 10318 40230 10364 40282
rect 10068 40228 10124 40230
rect 10148 40228 10204 40230
rect 10228 40228 10284 40230
rect 10308 40228 10364 40230
rect 9126 38392 9182 38448
rect 9402 38120 9458 38176
rect 8482 37440 8538 37496
rect 7930 36796 7932 36816
rect 7932 36796 7984 36816
rect 7984 36796 7986 36816
rect 7930 36760 7986 36796
rect 8390 36660 8392 36680
rect 8392 36660 8444 36680
rect 8444 36660 8446 36680
rect 8390 36624 8446 36660
rect 8666 37440 8722 37496
rect 8574 37168 8630 37224
rect 8390 36080 8446 36136
rect 8482 35944 8538 36000
rect 8574 35672 8630 35728
rect 6918 32136 6974 32192
rect 7102 32000 7158 32056
rect 7010 31864 7066 31920
rect 6734 31764 6736 31784
rect 6736 31764 6788 31784
rect 6788 31764 6790 31784
rect 6734 31728 6790 31764
rect 6734 31628 6736 31648
rect 6736 31628 6788 31648
rect 6788 31628 6790 31648
rect 6734 31592 6790 31628
rect 7010 31728 7066 31784
rect 5998 27784 6054 27840
rect 5814 27276 5816 27296
rect 5816 27276 5868 27296
rect 5868 27276 5870 27296
rect 5814 27240 5870 27276
rect 5814 26696 5870 26752
rect 5722 26016 5778 26072
rect 5722 25916 5724 25936
rect 5724 25916 5776 25936
rect 5776 25916 5778 25936
rect 5722 25880 5778 25916
rect 5722 24928 5778 24984
rect 5722 24812 5778 24848
rect 5722 24792 5724 24812
rect 5724 24792 5776 24812
rect 5776 24792 5778 24812
rect 5630 24692 5632 24712
rect 5632 24692 5684 24712
rect 5684 24692 5686 24712
rect 5630 24656 5686 24692
rect 5262 23840 5318 23896
rect 5722 24384 5778 24440
rect 5906 26424 5962 26480
rect 5906 25744 5962 25800
rect 5906 25200 5962 25256
rect 5906 24792 5962 24848
rect 6550 30540 6552 30560
rect 6552 30540 6604 30560
rect 6604 30540 6606 30560
rect 6550 30504 6606 30540
rect 6734 29824 6790 29880
rect 6550 29280 6606 29336
rect 6458 29144 6514 29200
rect 6366 28872 6422 28928
rect 6182 28192 6238 28248
rect 6182 28092 6184 28112
rect 6184 28092 6236 28112
rect 6236 28092 6238 28112
rect 6182 28056 6238 28092
rect 6826 29008 6882 29064
rect 6274 27240 6330 27296
rect 6458 27920 6514 27976
rect 6734 27648 6790 27704
rect 6458 26968 6514 27024
rect 6458 26560 6514 26616
rect 6090 25880 6146 25936
rect 6090 24792 6146 24848
rect 5630 23568 5686 23624
rect 4802 21120 4858 21176
rect 4710 20984 4766 21040
rect 4986 20984 5042 21040
rect 4802 20848 4858 20904
rect 4250 20712 4306 20768
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 4526 19896 4582 19952
rect 4066 19624 4122 19680
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 3238 19352 3240 19372
rect 3240 19352 3292 19372
rect 3292 19352 3294 19372
rect 3146 18808 3202 18864
rect 2686 16904 2742 16960
rect 3146 17212 3148 17232
rect 3148 17212 3200 17232
rect 3200 17212 3202 17232
rect 2870 17040 2926 17096
rect 3146 17176 3202 17212
rect 2778 15544 2834 15600
rect 2226 15156 2282 15192
rect 2226 15136 2228 15156
rect 2228 15136 2280 15156
rect 2280 15136 2282 15156
rect 1858 12416 1914 12472
rect 1582 12008 1638 12064
rect 1490 11464 1546 11520
rect 1398 11192 1454 11248
rect 1950 12008 2006 12064
rect 1582 10920 1638 10976
rect 1950 9036 2006 9072
rect 1950 9016 1952 9036
rect 1952 9016 2004 9036
rect 2004 9016 2006 9036
rect 2686 14612 2742 14648
rect 2686 14592 2688 14612
rect 2688 14592 2740 14612
rect 2740 14592 2742 14612
rect 2226 12316 2228 12336
rect 2228 12316 2280 12336
rect 2280 12316 2282 12336
rect 2226 12280 2282 12316
rect 2594 12824 2650 12880
rect 2870 13388 2926 13424
rect 2870 13368 2872 13388
rect 2872 13368 2924 13388
rect 2924 13368 2926 13388
rect 2686 12436 2742 12472
rect 2686 12416 2688 12436
rect 2688 12416 2740 12436
rect 2740 12416 2742 12436
rect 2686 12300 2742 12336
rect 2962 13232 3018 13288
rect 3422 18128 3478 18184
rect 3882 18672 3938 18728
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 3422 17312 3478 17368
rect 4342 19216 4398 19272
rect 4526 19236 4582 19272
rect 4526 19216 4528 19236
rect 4528 19216 4580 19236
rect 4580 19216 4582 19236
rect 5354 22888 5410 22944
rect 5262 22208 5318 22264
rect 5262 21936 5318 21992
rect 5170 21684 5226 21720
rect 5170 21664 5172 21684
rect 5172 21664 5224 21684
rect 5224 21664 5226 21684
rect 5446 22652 5448 22672
rect 5448 22652 5500 22672
rect 5500 22652 5502 22672
rect 5446 22616 5502 22652
rect 5446 21664 5502 21720
rect 5170 20712 5226 20768
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 4710 18944 4766 19000
rect 4158 18572 4160 18592
rect 4160 18572 4212 18592
rect 4212 18572 4214 18592
rect 4158 18536 4214 18572
rect 3974 17720 4030 17776
rect 3790 17584 3846 17640
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 3698 17176 3754 17232
rect 3974 17040 4030 17096
rect 3790 16904 3846 16960
rect 3882 16532 3884 16552
rect 3884 16532 3936 16552
rect 3936 16532 3938 16552
rect 3882 16496 3938 16532
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 3698 16088 3754 16144
rect 4342 18400 4398 18456
rect 4710 18400 4766 18456
rect 4802 17992 4858 18048
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 4802 17856 4858 17912
rect 4250 17176 4306 17232
rect 4434 17448 4490 17504
rect 4710 17720 4766 17776
rect 4526 17176 4582 17232
rect 4434 17040 4490 17096
rect 4802 17312 4858 17368
rect 4710 16904 4766 16960
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 4710 16496 4766 16552
rect 3146 13796 3202 13832
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 3146 13776 3148 13796
rect 3148 13776 3200 13796
rect 3200 13776 3202 13796
rect 3238 13640 3294 13696
rect 3238 13232 3294 13288
rect 2686 12280 2688 12300
rect 2688 12280 2740 12300
rect 2740 12280 2742 12300
rect 3054 13096 3110 13152
rect 2962 12008 3018 12064
rect 2778 11736 2834 11792
rect 2870 10124 2926 10160
rect 2870 10104 2872 10124
rect 2872 10104 2924 10124
rect 2924 10104 2926 10124
rect 3330 13132 3332 13152
rect 3332 13132 3384 13152
rect 3384 13132 3386 13152
rect 3330 13096 3386 13132
rect 3974 14900 3976 14920
rect 3976 14900 4028 14920
rect 4028 14900 4030 14920
rect 3974 14864 4030 14900
rect 3882 14728 3938 14784
rect 3698 14320 3754 14376
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 3790 13912 3846 13968
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 5078 20304 5134 20360
rect 4986 19488 5042 19544
rect 5354 21256 5410 21312
rect 5722 23432 5778 23488
rect 5906 22888 5962 22944
rect 6734 26560 6790 26616
rect 6642 26152 6698 26208
rect 6642 25608 6698 25664
rect 6734 25472 6790 25528
rect 6458 25064 6514 25120
rect 6458 24520 6514 24576
rect 6182 23840 6238 23896
rect 6090 23296 6146 23352
rect 6274 23316 6330 23352
rect 6274 23296 6276 23316
rect 6276 23296 6328 23316
rect 6328 23296 6330 23316
rect 5998 21936 6054 21992
rect 5538 21120 5594 21176
rect 5998 21528 6054 21584
rect 5906 21256 5962 21312
rect 6182 22616 6238 22672
rect 6274 21956 6330 21992
rect 6274 21936 6276 21956
rect 6276 21936 6328 21956
rect 6328 21936 6330 21956
rect 6090 20984 6146 21040
rect 5998 20848 6054 20904
rect 5630 20052 5686 20088
rect 5630 20032 5632 20052
rect 5632 20032 5684 20052
rect 5684 20032 5686 20052
rect 5722 19760 5778 19816
rect 5630 19624 5686 19680
rect 5538 19216 5594 19272
rect 5630 19080 5686 19136
rect 5078 18828 5134 18864
rect 5078 18808 5080 18828
rect 5080 18808 5132 18828
rect 5132 18808 5134 18828
rect 5078 18536 5134 18592
rect 5170 18420 5226 18456
rect 5170 18400 5172 18420
rect 5172 18400 5224 18420
rect 5224 18400 5226 18420
rect 5078 18264 5134 18320
rect 4986 18128 5042 18184
rect 5170 18164 5172 18184
rect 5172 18164 5224 18184
rect 5224 18164 5226 18184
rect 5170 18128 5226 18164
rect 5170 17992 5226 18048
rect 5262 17740 5318 17776
rect 5262 17720 5264 17740
rect 5264 17720 5316 17740
rect 5316 17720 5318 17740
rect 5262 17448 5318 17504
rect 4250 15136 4306 15192
rect 4158 14340 4214 14376
rect 4158 14320 4160 14340
rect 4160 14320 4212 14340
rect 4212 14320 4214 14340
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 3698 12144 3754 12200
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 3146 6296 3202 6352
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 3882 10124 3938 10160
rect 3882 10104 3884 10124
rect 3884 10104 3936 10124
rect 3936 10104 3938 10124
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 4342 13368 4398 13424
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 4710 12144 4766 12200
rect 5078 14220 5080 14240
rect 5080 14220 5132 14240
rect 5132 14220 5134 14240
rect 5078 14184 5134 14220
rect 5170 13912 5226 13968
rect 4894 13388 4950 13424
rect 4894 13368 4896 13388
rect 4896 13368 4948 13388
rect 4948 13368 4950 13388
rect 5078 12416 5134 12472
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 6274 21256 6330 21312
rect 6090 20032 6146 20088
rect 5722 18672 5778 18728
rect 5538 18536 5594 18592
rect 5722 18420 5778 18456
rect 5722 18400 5724 18420
rect 5724 18400 5776 18420
rect 5776 18400 5778 18420
rect 5722 18284 5778 18320
rect 5906 19352 5962 19408
rect 6090 18944 6146 19000
rect 6090 18400 6146 18456
rect 5722 18264 5724 18284
rect 5724 18264 5776 18284
rect 5776 18264 5778 18284
rect 5538 18128 5594 18184
rect 5722 18128 5778 18184
rect 5446 16768 5502 16824
rect 5722 17584 5778 17640
rect 5722 17040 5778 17096
rect 5906 16632 5962 16688
rect 6550 24384 6606 24440
rect 7562 31884 7618 31920
rect 7562 31864 7564 31884
rect 7564 31864 7616 31884
rect 7616 31864 7618 31884
rect 7838 34484 7840 34504
rect 7840 34484 7892 34504
rect 7892 34484 7894 34504
rect 7838 34448 7894 34484
rect 7838 34060 7894 34096
rect 7838 34040 7840 34060
rect 7840 34040 7892 34060
rect 7892 34040 7894 34060
rect 8298 35148 8354 35184
rect 8942 37188 8998 37224
rect 8942 37168 8944 37188
rect 8944 37168 8996 37188
rect 8996 37168 8998 37188
rect 8942 36352 8998 36408
rect 10728 41914 10784 41916
rect 10808 41914 10864 41916
rect 10888 41914 10944 41916
rect 10968 41914 11024 41916
rect 10728 41862 10774 41914
rect 10774 41862 10784 41914
rect 10808 41862 10838 41914
rect 10838 41862 10850 41914
rect 10850 41862 10864 41914
rect 10888 41862 10902 41914
rect 10902 41862 10914 41914
rect 10914 41862 10944 41914
rect 10968 41862 10978 41914
rect 10978 41862 11024 41914
rect 10728 41860 10784 41862
rect 10808 41860 10864 41862
rect 10888 41860 10944 41862
rect 10968 41860 11024 41862
rect 10230 39480 10286 39536
rect 10138 39344 10194 39400
rect 10068 39194 10124 39196
rect 10148 39194 10204 39196
rect 10228 39194 10284 39196
rect 10308 39194 10364 39196
rect 10068 39142 10114 39194
rect 10114 39142 10124 39194
rect 10148 39142 10178 39194
rect 10178 39142 10190 39194
rect 10190 39142 10204 39194
rect 10228 39142 10242 39194
rect 10242 39142 10254 39194
rect 10254 39142 10284 39194
rect 10308 39142 10318 39194
rect 10318 39142 10364 39194
rect 10068 39140 10124 39142
rect 10148 39140 10204 39142
rect 10228 39140 10284 39142
rect 10308 39140 10364 39142
rect 9862 38936 9918 38992
rect 9770 38800 9826 38856
rect 9586 37848 9642 37904
rect 9402 37612 9404 37632
rect 9404 37612 9456 37632
rect 9456 37612 9458 37632
rect 9402 37576 9458 37612
rect 9310 37440 9366 37496
rect 9402 37168 9458 37224
rect 9218 36524 9220 36544
rect 9220 36524 9272 36544
rect 9272 36524 9274 36544
rect 9218 36488 9274 36524
rect 8298 35128 8300 35148
rect 8300 35128 8352 35148
rect 8352 35128 8354 35148
rect 7930 33224 7986 33280
rect 8022 32680 8078 32736
rect 7930 32544 7986 32600
rect 7746 32000 7802 32056
rect 7470 31456 7526 31512
rect 7194 30252 7250 30288
rect 7194 30232 7196 30252
rect 7196 30232 7248 30252
rect 7248 30232 7250 30252
rect 7102 29552 7158 29608
rect 7562 30796 7618 30832
rect 7562 30776 7564 30796
rect 7564 30776 7616 30796
rect 7616 30776 7618 30796
rect 7102 29300 7158 29336
rect 7102 29280 7104 29300
rect 7104 29280 7156 29300
rect 7156 29280 7158 29300
rect 7286 29416 7342 29472
rect 7194 29044 7196 29064
rect 7196 29044 7248 29064
rect 7248 29044 7250 29064
rect 7194 29008 7250 29044
rect 6918 28872 6974 28928
rect 6918 28464 6974 28520
rect 7102 28328 7158 28384
rect 6918 27940 6974 27976
rect 6918 27920 6920 27940
rect 6920 27920 6972 27940
rect 6972 27920 6974 27940
rect 7194 27784 7250 27840
rect 7470 30368 7526 30424
rect 7378 28464 7434 28520
rect 7378 27648 7434 27704
rect 7286 27512 7342 27568
rect 7194 26968 7250 27024
rect 7010 26832 7066 26888
rect 6918 26696 6974 26752
rect 7010 25472 7066 25528
rect 6918 25336 6974 25392
rect 6918 24404 6974 24440
rect 6918 24384 6920 24404
rect 6920 24384 6972 24404
rect 6972 24384 6974 24404
rect 6918 23976 6974 24032
rect 7194 26444 7250 26480
rect 7194 26424 7196 26444
rect 7196 26424 7248 26444
rect 7248 26424 7250 26444
rect 7746 30096 7802 30152
rect 7838 29552 7894 29608
rect 7654 28620 7710 28656
rect 7654 28600 7656 28620
rect 7656 28600 7708 28620
rect 7708 28600 7710 28620
rect 7470 26188 7472 26208
rect 7472 26188 7524 26208
rect 7524 26188 7526 26208
rect 7470 26152 7526 26188
rect 7378 25064 7434 25120
rect 8574 34584 8630 34640
rect 8482 34448 8538 34504
rect 8206 33940 8208 33960
rect 8208 33940 8260 33960
rect 8260 33940 8262 33960
rect 8206 33904 8262 33940
rect 8206 33496 8262 33552
rect 8850 34992 8906 35048
rect 8574 34040 8630 34096
rect 8850 34040 8906 34096
rect 8390 33224 8446 33280
rect 8758 33904 8814 33960
rect 8574 33496 8630 33552
rect 8758 33224 8814 33280
rect 8758 33088 8814 33144
rect 8390 32816 8446 32872
rect 8482 32680 8538 32736
rect 8298 32020 8354 32056
rect 8298 32000 8300 32020
rect 8300 32000 8352 32020
rect 8352 32000 8354 32020
rect 8114 31592 8170 31648
rect 8022 28872 8078 28928
rect 8942 32544 8998 32600
rect 9034 32272 9090 32328
rect 10138 38836 10140 38856
rect 10140 38836 10192 38856
rect 10192 38836 10194 38856
rect 10138 38800 10194 38836
rect 10322 38528 10378 38584
rect 9862 37984 9918 38040
rect 10068 38106 10124 38108
rect 10148 38106 10204 38108
rect 10228 38106 10284 38108
rect 10308 38106 10364 38108
rect 10068 38054 10114 38106
rect 10114 38054 10124 38106
rect 10148 38054 10178 38106
rect 10178 38054 10190 38106
rect 10190 38054 10204 38106
rect 10228 38054 10242 38106
rect 10242 38054 10254 38106
rect 10254 38054 10284 38106
rect 10308 38054 10318 38106
rect 10318 38054 10364 38106
rect 10068 38052 10124 38054
rect 10148 38052 10204 38054
rect 10228 38052 10284 38054
rect 10308 38052 10364 38054
rect 9770 37712 9826 37768
rect 10728 40826 10784 40828
rect 10808 40826 10864 40828
rect 10888 40826 10944 40828
rect 10968 40826 11024 40828
rect 10728 40774 10774 40826
rect 10774 40774 10784 40826
rect 10808 40774 10838 40826
rect 10838 40774 10850 40826
rect 10850 40774 10864 40826
rect 10888 40774 10902 40826
rect 10902 40774 10914 40826
rect 10914 40774 10944 40826
rect 10968 40774 10978 40826
rect 10978 40774 11024 40826
rect 10728 40772 10784 40774
rect 10808 40772 10864 40774
rect 10888 40772 10944 40774
rect 10968 40772 11024 40774
rect 10690 40024 10746 40080
rect 9770 37304 9826 37360
rect 9494 36352 9550 36408
rect 9218 34584 9274 34640
rect 9218 34448 9274 34504
rect 10068 37018 10124 37020
rect 10148 37018 10204 37020
rect 10228 37018 10284 37020
rect 10308 37018 10364 37020
rect 10068 36966 10114 37018
rect 10114 36966 10124 37018
rect 10148 36966 10178 37018
rect 10178 36966 10190 37018
rect 10190 36966 10204 37018
rect 10228 36966 10242 37018
rect 10242 36966 10254 37018
rect 10254 36966 10284 37018
rect 10308 36966 10318 37018
rect 10318 36966 10364 37018
rect 10068 36964 10124 36966
rect 10148 36964 10204 36966
rect 10228 36964 10284 36966
rect 10308 36964 10364 36966
rect 9862 36644 9918 36680
rect 9862 36624 9864 36644
rect 9864 36624 9916 36644
rect 9916 36624 9918 36644
rect 10690 39908 10746 39944
rect 10690 39888 10692 39908
rect 10692 39888 10744 39908
rect 10744 39888 10746 39908
rect 10728 39738 10784 39740
rect 10808 39738 10864 39740
rect 10888 39738 10944 39740
rect 10968 39738 11024 39740
rect 10728 39686 10774 39738
rect 10774 39686 10784 39738
rect 10808 39686 10838 39738
rect 10838 39686 10850 39738
rect 10850 39686 10864 39738
rect 10888 39686 10902 39738
rect 10902 39686 10914 39738
rect 10914 39686 10944 39738
rect 10968 39686 10978 39738
rect 10978 39686 11024 39738
rect 10728 39684 10784 39686
rect 10808 39684 10864 39686
rect 10888 39684 10944 39686
rect 10968 39684 11024 39686
rect 10728 38650 10784 38652
rect 10808 38650 10864 38652
rect 10888 38650 10944 38652
rect 10968 38650 11024 38652
rect 10728 38598 10774 38650
rect 10774 38598 10784 38650
rect 10808 38598 10838 38650
rect 10838 38598 10850 38650
rect 10850 38598 10864 38650
rect 10888 38598 10902 38650
rect 10902 38598 10914 38650
rect 10914 38598 10944 38650
rect 10968 38598 10978 38650
rect 10978 38598 11024 38650
rect 10728 38596 10784 38598
rect 10808 38596 10864 38598
rect 10888 38596 10944 38598
rect 10968 38596 11024 38598
rect 10728 37562 10784 37564
rect 10808 37562 10864 37564
rect 10888 37562 10944 37564
rect 10968 37562 11024 37564
rect 10728 37510 10774 37562
rect 10774 37510 10784 37562
rect 10808 37510 10838 37562
rect 10838 37510 10850 37562
rect 10850 37510 10864 37562
rect 10888 37510 10902 37562
rect 10902 37510 10914 37562
rect 10914 37510 10944 37562
rect 10968 37510 10978 37562
rect 10978 37510 11024 37562
rect 10728 37508 10784 37510
rect 10808 37508 10864 37510
rect 10888 37508 10944 37510
rect 10968 37508 11024 37510
rect 10728 36474 10784 36476
rect 10808 36474 10864 36476
rect 10888 36474 10944 36476
rect 10968 36474 11024 36476
rect 10728 36422 10774 36474
rect 10774 36422 10784 36474
rect 10808 36422 10838 36474
rect 10838 36422 10850 36474
rect 10850 36422 10864 36474
rect 10888 36422 10902 36474
rect 10902 36422 10914 36474
rect 10914 36422 10944 36474
rect 10968 36422 10978 36474
rect 10978 36422 11024 36474
rect 10728 36420 10784 36422
rect 10808 36420 10864 36422
rect 10888 36420 10944 36422
rect 10968 36420 11024 36422
rect 9218 33260 9220 33280
rect 9220 33260 9272 33280
rect 9272 33260 9274 33280
rect 9218 33224 9274 33260
rect 8942 32000 8998 32056
rect 8758 31728 8814 31784
rect 8206 29416 8262 29472
rect 8206 28328 8262 28384
rect 8206 28192 8262 28248
rect 8022 27512 8078 27568
rect 8206 27648 8262 27704
rect 8114 27104 8170 27160
rect 8022 26424 8078 26480
rect 7930 26152 7986 26208
rect 7838 25880 7894 25936
rect 7470 24928 7526 24984
rect 7470 24792 7526 24848
rect 7378 24384 7434 24440
rect 7470 24268 7526 24304
rect 7470 24248 7472 24268
rect 7472 24248 7524 24268
rect 7524 24248 7526 24268
rect 6826 22888 6882 22944
rect 7378 23976 7434 24032
rect 7378 23840 7434 23896
rect 6734 22616 6790 22672
rect 6734 22344 6790 22400
rect 6642 22228 6698 22264
rect 6642 22208 6644 22228
rect 6644 22208 6696 22228
rect 6696 22208 6698 22228
rect 7102 22616 7158 22672
rect 7286 23024 7342 23080
rect 7102 22208 7158 22264
rect 6550 21936 6606 21992
rect 6550 18148 6606 18184
rect 6550 18128 6552 18148
rect 6552 18128 6604 18148
rect 6604 18128 6606 18148
rect 6274 17604 6330 17640
rect 6274 17584 6276 17604
rect 6276 17584 6328 17604
rect 6328 17584 6330 17604
rect 6274 17312 6330 17368
rect 6550 17992 6606 18048
rect 6826 21392 6882 21448
rect 7746 25064 7802 25120
rect 8022 24792 8078 24848
rect 7746 23840 7802 23896
rect 7930 23840 7986 23896
rect 7194 21256 7250 21312
rect 6826 20304 6882 20360
rect 7286 20304 7342 20360
rect 6918 19624 6974 19680
rect 6826 18808 6882 18864
rect 6826 18400 6882 18456
rect 7838 23588 7894 23624
rect 7838 23568 7840 23588
rect 7840 23568 7892 23588
rect 7892 23568 7894 23588
rect 7562 21936 7618 21992
rect 7746 22208 7802 22264
rect 7930 22228 7986 22264
rect 7930 22208 7932 22228
rect 7932 22208 7984 22228
rect 7984 22208 7986 22228
rect 8206 23296 8262 23352
rect 8206 23196 8208 23216
rect 8208 23196 8260 23216
rect 8260 23196 8262 23216
rect 8206 23160 8262 23196
rect 7838 20848 7894 20904
rect 7562 20440 7618 20496
rect 7286 18536 7342 18592
rect 7286 18400 7342 18456
rect 6642 17312 6698 17368
rect 6826 17196 6882 17232
rect 6826 17176 6828 17196
rect 6828 17176 6880 17196
rect 6880 17176 6882 17196
rect 6826 16788 6882 16824
rect 6826 16768 6828 16788
rect 6828 16768 6880 16788
rect 6880 16768 6882 16788
rect 6366 16496 6422 16552
rect 6090 15000 6146 15056
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 4802 10104 4858 10160
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 3790 6332 3792 6352
rect 3792 6332 3844 6352
rect 3844 6332 3846 6352
rect 3790 6296 3846 6332
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 6826 16652 6882 16688
rect 6826 16632 6828 16652
rect 6828 16632 6880 16652
rect 6880 16632 6882 16652
rect 6550 16532 6552 16552
rect 6552 16532 6604 16552
rect 6604 16532 6606 16552
rect 6550 16496 6606 16532
rect 6642 16360 6698 16416
rect 6550 15272 6606 15328
rect 6366 12824 6422 12880
rect 5630 10548 5632 10568
rect 5632 10548 5684 10568
rect 5684 10548 5686 10568
rect 5630 10512 5686 10548
rect 6642 14864 6698 14920
rect 7194 17856 7250 17912
rect 7746 20032 7802 20088
rect 7654 19352 7710 19408
rect 7470 18264 7526 18320
rect 7654 18300 7656 18320
rect 7656 18300 7708 18320
rect 7708 18300 7710 18320
rect 7654 18264 7710 18300
rect 7470 18128 7526 18184
rect 7378 17856 7434 17912
rect 7562 17856 7618 17912
rect 7746 17992 7802 18048
rect 7470 17584 7526 17640
rect 7562 17312 7618 17368
rect 7930 19932 7932 19952
rect 7932 19932 7984 19952
rect 7984 19932 7986 19952
rect 7930 19896 7986 19932
rect 8206 21528 8262 21584
rect 8574 29044 8576 29064
rect 8576 29044 8628 29064
rect 8628 29044 8630 29064
rect 8574 29008 8630 29044
rect 8574 27512 8630 27568
rect 8574 26968 8630 27024
rect 8574 26696 8630 26752
rect 9402 32952 9458 33008
rect 9310 32408 9366 32464
rect 8850 30504 8906 30560
rect 8942 27512 8998 27568
rect 8942 27240 8998 27296
rect 8482 25780 8484 25800
rect 8484 25780 8536 25800
rect 8536 25780 8538 25800
rect 8482 25744 8538 25780
rect 8758 25608 8814 25664
rect 8574 25492 8630 25528
rect 8574 25472 8576 25492
rect 8576 25472 8628 25492
rect 8628 25472 8630 25492
rect 8574 25356 8630 25392
rect 8574 25336 8576 25356
rect 8576 25336 8628 25356
rect 8628 25336 8630 25356
rect 8666 25064 8722 25120
rect 8574 24656 8630 24712
rect 8390 23860 8446 23896
rect 8390 23840 8392 23860
rect 8392 23840 8444 23860
rect 8444 23840 8446 23860
rect 8390 23568 8446 23624
rect 8574 24248 8630 24304
rect 9126 31592 9182 31648
rect 10598 36080 10654 36136
rect 10068 35930 10124 35932
rect 10148 35930 10204 35932
rect 10228 35930 10284 35932
rect 10308 35930 10364 35932
rect 10068 35878 10114 35930
rect 10114 35878 10124 35930
rect 10148 35878 10178 35930
rect 10178 35878 10190 35930
rect 10190 35878 10204 35930
rect 10228 35878 10242 35930
rect 10242 35878 10254 35930
rect 10254 35878 10284 35930
rect 10308 35878 10318 35930
rect 10318 35878 10364 35930
rect 10068 35876 10124 35878
rect 10148 35876 10204 35878
rect 10228 35876 10284 35878
rect 10308 35876 10364 35878
rect 9954 35128 10010 35184
rect 10728 35386 10784 35388
rect 10808 35386 10864 35388
rect 10888 35386 10944 35388
rect 10968 35386 11024 35388
rect 10728 35334 10774 35386
rect 10774 35334 10784 35386
rect 10808 35334 10838 35386
rect 10838 35334 10850 35386
rect 10850 35334 10864 35386
rect 10888 35334 10902 35386
rect 10902 35334 10914 35386
rect 10914 35334 10944 35386
rect 10968 35334 10978 35386
rect 10978 35334 11024 35386
rect 10728 35332 10784 35334
rect 10808 35332 10864 35334
rect 10888 35332 10944 35334
rect 10968 35332 11024 35334
rect 10598 34992 10654 35048
rect 10068 34842 10124 34844
rect 10148 34842 10204 34844
rect 10228 34842 10284 34844
rect 10308 34842 10364 34844
rect 10068 34790 10114 34842
rect 10114 34790 10124 34842
rect 10148 34790 10178 34842
rect 10178 34790 10190 34842
rect 10190 34790 10204 34842
rect 10228 34790 10242 34842
rect 10242 34790 10254 34842
rect 10254 34790 10284 34842
rect 10308 34790 10318 34842
rect 10318 34790 10364 34842
rect 10068 34788 10124 34790
rect 10148 34788 10204 34790
rect 10228 34788 10284 34790
rect 10308 34788 10364 34790
rect 9862 33632 9918 33688
rect 9494 32272 9550 32328
rect 9126 29008 9182 29064
rect 10966 34484 10968 34504
rect 10968 34484 11020 34504
rect 11020 34484 11022 34504
rect 10068 33754 10124 33756
rect 10148 33754 10204 33756
rect 10228 33754 10284 33756
rect 10308 33754 10364 33756
rect 10068 33702 10114 33754
rect 10114 33702 10124 33754
rect 10148 33702 10178 33754
rect 10178 33702 10190 33754
rect 10190 33702 10204 33754
rect 10228 33702 10242 33754
rect 10242 33702 10254 33754
rect 10254 33702 10284 33754
rect 10308 33702 10318 33754
rect 10318 33702 10364 33754
rect 10068 33700 10124 33702
rect 10148 33700 10204 33702
rect 10228 33700 10284 33702
rect 10308 33700 10364 33702
rect 10414 33396 10416 33416
rect 10416 33396 10468 33416
rect 10468 33396 10470 33416
rect 10414 33360 10470 33396
rect 10068 32666 10124 32668
rect 10148 32666 10204 32668
rect 10228 32666 10284 32668
rect 10308 32666 10364 32668
rect 10068 32614 10114 32666
rect 10114 32614 10124 32666
rect 10148 32614 10178 32666
rect 10178 32614 10190 32666
rect 10190 32614 10204 32666
rect 10228 32614 10242 32666
rect 10242 32614 10254 32666
rect 10254 32614 10284 32666
rect 10308 32614 10318 32666
rect 10318 32614 10364 32666
rect 10068 32612 10124 32614
rect 10148 32612 10204 32614
rect 10228 32612 10284 32614
rect 10308 32612 10364 32614
rect 10966 34448 11022 34484
rect 10728 34298 10784 34300
rect 10808 34298 10864 34300
rect 10888 34298 10944 34300
rect 10968 34298 11024 34300
rect 10728 34246 10774 34298
rect 10774 34246 10784 34298
rect 10808 34246 10838 34298
rect 10838 34246 10850 34298
rect 10850 34246 10864 34298
rect 10888 34246 10902 34298
rect 10902 34246 10914 34298
rect 10914 34246 10944 34298
rect 10968 34246 10978 34298
rect 10978 34246 11024 34298
rect 10728 34244 10784 34246
rect 10808 34244 10864 34246
rect 10888 34244 10944 34246
rect 10968 34244 11024 34246
rect 10728 33210 10784 33212
rect 10808 33210 10864 33212
rect 10888 33210 10944 33212
rect 10968 33210 11024 33212
rect 10728 33158 10774 33210
rect 10774 33158 10784 33210
rect 10808 33158 10838 33210
rect 10838 33158 10850 33210
rect 10850 33158 10864 33210
rect 10888 33158 10902 33210
rect 10902 33158 10914 33210
rect 10914 33158 10944 33210
rect 10968 33158 10978 33210
rect 10978 33158 11024 33210
rect 10728 33156 10784 33158
rect 10808 33156 10864 33158
rect 10888 33156 10944 33158
rect 10968 33156 11024 33158
rect 10046 31764 10048 31784
rect 10048 31764 10100 31784
rect 10100 31764 10102 31784
rect 10046 31728 10102 31764
rect 10068 31578 10124 31580
rect 10148 31578 10204 31580
rect 10228 31578 10284 31580
rect 10308 31578 10364 31580
rect 10068 31526 10114 31578
rect 10114 31526 10124 31578
rect 10148 31526 10178 31578
rect 10178 31526 10190 31578
rect 10190 31526 10204 31578
rect 10228 31526 10242 31578
rect 10242 31526 10254 31578
rect 10254 31526 10284 31578
rect 10308 31526 10318 31578
rect 10318 31526 10364 31578
rect 10068 31524 10124 31526
rect 10148 31524 10204 31526
rect 10228 31524 10284 31526
rect 10308 31524 10364 31526
rect 9954 30640 10010 30696
rect 10728 32122 10784 32124
rect 10808 32122 10864 32124
rect 10888 32122 10944 32124
rect 10968 32122 11024 32124
rect 10728 32070 10774 32122
rect 10774 32070 10784 32122
rect 10808 32070 10838 32122
rect 10838 32070 10850 32122
rect 10850 32070 10864 32122
rect 10888 32070 10902 32122
rect 10902 32070 10914 32122
rect 10914 32070 10944 32122
rect 10968 32070 10978 32122
rect 10978 32070 11024 32122
rect 10728 32068 10784 32070
rect 10808 32068 10864 32070
rect 10888 32068 10944 32070
rect 10968 32068 11024 32070
rect 10728 31034 10784 31036
rect 10808 31034 10864 31036
rect 10888 31034 10944 31036
rect 10968 31034 11024 31036
rect 10728 30982 10774 31034
rect 10774 30982 10784 31034
rect 10808 30982 10838 31034
rect 10838 30982 10850 31034
rect 10850 30982 10864 31034
rect 10888 30982 10902 31034
rect 10902 30982 10914 31034
rect 10914 30982 10944 31034
rect 10968 30982 10978 31034
rect 10978 30982 11024 31034
rect 10728 30980 10784 30982
rect 10808 30980 10864 30982
rect 10888 30980 10944 30982
rect 10968 30980 11024 30982
rect 10068 30490 10124 30492
rect 10148 30490 10204 30492
rect 10228 30490 10284 30492
rect 10308 30490 10364 30492
rect 10068 30438 10114 30490
rect 10114 30438 10124 30490
rect 10148 30438 10178 30490
rect 10178 30438 10190 30490
rect 10190 30438 10204 30490
rect 10228 30438 10242 30490
rect 10242 30438 10254 30490
rect 10254 30438 10284 30490
rect 10308 30438 10318 30490
rect 10318 30438 10364 30490
rect 10068 30436 10124 30438
rect 10148 30436 10204 30438
rect 10228 30436 10284 30438
rect 10308 30436 10364 30438
rect 9770 30232 9826 30288
rect 9494 28736 9550 28792
rect 9402 28636 9404 28656
rect 9404 28636 9456 28656
rect 9456 28636 9458 28656
rect 9402 28600 9458 28636
rect 9126 27956 9128 27976
rect 9128 27956 9180 27976
rect 9180 27956 9182 27976
rect 9126 27920 9182 27956
rect 9494 28364 9496 28384
rect 9496 28364 9548 28384
rect 9548 28364 9550 28384
rect 9494 28328 9550 28364
rect 9126 27376 9182 27432
rect 9126 26868 9128 26888
rect 9128 26868 9180 26888
rect 9180 26868 9182 26888
rect 9126 26832 9182 26868
rect 9310 26288 9366 26344
rect 9126 24928 9182 24984
rect 9218 24384 9274 24440
rect 8850 24248 8906 24304
rect 8666 23976 8722 24032
rect 8942 23976 8998 24032
rect 8666 23568 8722 23624
rect 8574 22516 8576 22536
rect 8576 22516 8628 22536
rect 8628 22516 8630 22536
rect 8574 22480 8630 22516
rect 8390 21936 8446 21992
rect 8758 22208 8814 22264
rect 9034 23740 9036 23760
rect 9036 23740 9088 23760
rect 9088 23740 9090 23760
rect 9034 23704 9090 23740
rect 9034 23180 9090 23216
rect 9034 23160 9036 23180
rect 9036 23160 9088 23180
rect 9088 23160 9090 23180
rect 9218 24012 9220 24032
rect 9220 24012 9272 24032
rect 9272 24012 9274 24032
rect 9218 23976 9274 24012
rect 9218 23840 9274 23896
rect 10728 29946 10784 29948
rect 10808 29946 10864 29948
rect 10888 29946 10944 29948
rect 10968 29946 11024 29948
rect 10728 29894 10774 29946
rect 10774 29894 10784 29946
rect 10808 29894 10838 29946
rect 10838 29894 10850 29946
rect 10850 29894 10864 29946
rect 10888 29894 10902 29946
rect 10902 29894 10914 29946
rect 10914 29894 10944 29946
rect 10968 29894 10978 29946
rect 10978 29894 11024 29946
rect 10728 29892 10784 29894
rect 10808 29892 10864 29894
rect 10888 29892 10944 29894
rect 10968 29892 11024 29894
rect 10068 29402 10124 29404
rect 10148 29402 10204 29404
rect 10228 29402 10284 29404
rect 10308 29402 10364 29404
rect 10068 29350 10114 29402
rect 10114 29350 10124 29402
rect 10148 29350 10178 29402
rect 10178 29350 10190 29402
rect 10190 29350 10204 29402
rect 10228 29350 10242 29402
rect 10242 29350 10254 29402
rect 10254 29350 10284 29402
rect 10308 29350 10318 29402
rect 10318 29350 10364 29402
rect 10068 29348 10124 29350
rect 10148 29348 10204 29350
rect 10228 29348 10284 29350
rect 10308 29348 10364 29350
rect 9586 26460 9588 26480
rect 9588 26460 9640 26480
rect 9640 26460 9642 26480
rect 9586 26424 9642 26460
rect 9678 25744 9734 25800
rect 9586 24112 9642 24168
rect 9402 23976 9458 24032
rect 9402 23160 9458 23216
rect 9310 22888 9366 22944
rect 8850 22108 8852 22128
rect 8852 22108 8904 22128
rect 8904 22108 8906 22128
rect 8850 22072 8906 22108
rect 9126 22344 9182 22400
rect 8022 18672 8078 18728
rect 7930 17992 7986 18048
rect 8022 17856 8078 17912
rect 8390 20712 8446 20768
rect 8482 20440 8538 20496
rect 8666 19508 8722 19544
rect 8666 19488 8668 19508
rect 8668 19488 8720 19508
rect 8720 19488 8722 19508
rect 8390 18672 8446 18728
rect 8298 18400 8354 18456
rect 8206 17584 8262 17640
rect 8482 17584 8538 17640
rect 8482 17060 8538 17096
rect 7930 16496 7986 16552
rect 7562 15136 7618 15192
rect 7930 15408 7986 15464
rect 7378 14184 7434 14240
rect 6550 10512 6606 10568
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 6918 6704 6974 6760
rect 7746 13640 7802 13696
rect 8114 16904 8170 16960
rect 8482 17040 8484 17060
rect 8484 17040 8536 17060
rect 8536 17040 8538 17060
rect 8206 15408 8262 15464
rect 8114 13504 8170 13560
rect 7838 12824 7894 12880
rect 8390 16632 8446 16688
rect 8390 15700 8446 15736
rect 8390 15680 8392 15700
rect 8392 15680 8444 15700
rect 8444 15680 8446 15700
rect 8390 15408 8446 15464
rect 9034 21936 9090 21992
rect 9034 21528 9090 21584
rect 8850 20884 8852 20904
rect 8852 20884 8904 20904
rect 8904 20884 8906 20904
rect 8850 20848 8906 20884
rect 9218 21528 9274 21584
rect 9402 21664 9458 21720
rect 9218 20984 9274 21040
rect 9034 20848 9090 20904
rect 9126 20712 9182 20768
rect 9126 20168 9182 20224
rect 9126 19488 9182 19544
rect 9126 18808 9182 18864
rect 9126 18536 9182 18592
rect 9586 23604 9588 23624
rect 9588 23604 9640 23624
rect 9640 23604 9642 23624
rect 9586 23568 9642 23604
rect 9586 23468 9588 23488
rect 9588 23468 9640 23488
rect 9640 23468 9642 23488
rect 9586 23432 9642 23468
rect 10728 28858 10784 28860
rect 10808 28858 10864 28860
rect 10888 28858 10944 28860
rect 10968 28858 11024 28860
rect 10728 28806 10774 28858
rect 10774 28806 10784 28858
rect 10808 28806 10838 28858
rect 10838 28806 10850 28858
rect 10850 28806 10864 28858
rect 10888 28806 10902 28858
rect 10902 28806 10914 28858
rect 10914 28806 10944 28858
rect 10968 28806 10978 28858
rect 10978 28806 11024 28858
rect 10728 28804 10784 28806
rect 10808 28804 10864 28806
rect 10888 28804 10944 28806
rect 10968 28804 11024 28806
rect 10138 28464 10194 28520
rect 10068 28314 10124 28316
rect 10148 28314 10204 28316
rect 10228 28314 10284 28316
rect 10308 28314 10364 28316
rect 10068 28262 10114 28314
rect 10114 28262 10124 28314
rect 10148 28262 10178 28314
rect 10178 28262 10190 28314
rect 10190 28262 10204 28314
rect 10228 28262 10242 28314
rect 10242 28262 10254 28314
rect 10254 28262 10284 28314
rect 10308 28262 10318 28314
rect 10318 28262 10364 28314
rect 10068 28260 10124 28262
rect 10148 28260 10204 28262
rect 10228 28260 10284 28262
rect 10308 28260 10364 28262
rect 10138 27376 10194 27432
rect 10068 27226 10124 27228
rect 10148 27226 10204 27228
rect 10228 27226 10284 27228
rect 10308 27226 10364 27228
rect 10068 27174 10114 27226
rect 10114 27174 10124 27226
rect 10148 27174 10178 27226
rect 10178 27174 10190 27226
rect 10190 27174 10204 27226
rect 10228 27174 10242 27226
rect 10242 27174 10254 27226
rect 10254 27174 10284 27226
rect 10308 27174 10318 27226
rect 10318 27174 10364 27226
rect 10068 27172 10124 27174
rect 10148 27172 10204 27174
rect 10228 27172 10284 27174
rect 10308 27172 10364 27174
rect 10046 26968 10102 27024
rect 10046 26288 10102 26344
rect 9770 23976 9826 24032
rect 10068 26138 10124 26140
rect 10148 26138 10204 26140
rect 10228 26138 10284 26140
rect 10308 26138 10364 26140
rect 10068 26086 10114 26138
rect 10114 26086 10124 26138
rect 10148 26086 10178 26138
rect 10178 26086 10190 26138
rect 10190 26086 10204 26138
rect 10228 26086 10242 26138
rect 10242 26086 10254 26138
rect 10254 26086 10284 26138
rect 10308 26086 10318 26138
rect 10318 26086 10364 26138
rect 10068 26084 10124 26086
rect 10148 26084 10204 26086
rect 10228 26084 10284 26086
rect 10308 26084 10364 26086
rect 10068 25050 10124 25052
rect 10148 25050 10204 25052
rect 10228 25050 10284 25052
rect 10308 25050 10364 25052
rect 10068 24998 10114 25050
rect 10114 24998 10124 25050
rect 10148 24998 10178 25050
rect 10178 24998 10190 25050
rect 10190 24998 10204 25050
rect 10228 24998 10242 25050
rect 10242 24998 10254 25050
rect 10254 24998 10284 25050
rect 10308 24998 10318 25050
rect 10318 24998 10364 25050
rect 10068 24996 10124 24998
rect 10148 24996 10204 24998
rect 10228 24996 10284 24998
rect 10308 24996 10364 24998
rect 10046 24692 10048 24712
rect 10048 24692 10100 24712
rect 10100 24692 10102 24712
rect 10046 24656 10102 24692
rect 11058 27920 11114 27976
rect 10728 27770 10784 27772
rect 10808 27770 10864 27772
rect 10888 27770 10944 27772
rect 10968 27770 11024 27772
rect 10728 27718 10774 27770
rect 10774 27718 10784 27770
rect 10808 27718 10838 27770
rect 10838 27718 10850 27770
rect 10850 27718 10864 27770
rect 10888 27718 10902 27770
rect 10902 27718 10914 27770
rect 10914 27718 10944 27770
rect 10968 27718 10978 27770
rect 10978 27718 11024 27770
rect 10728 27716 10784 27718
rect 10808 27716 10864 27718
rect 10888 27716 10944 27718
rect 10968 27716 11024 27718
rect 10690 27512 10746 27568
rect 10690 26832 10746 26888
rect 10728 26682 10784 26684
rect 10808 26682 10864 26684
rect 10888 26682 10944 26684
rect 10968 26682 11024 26684
rect 10728 26630 10774 26682
rect 10774 26630 10784 26682
rect 10808 26630 10838 26682
rect 10838 26630 10850 26682
rect 10850 26630 10864 26682
rect 10888 26630 10902 26682
rect 10902 26630 10914 26682
rect 10914 26630 10944 26682
rect 10968 26630 10978 26682
rect 10978 26630 11024 26682
rect 10728 26628 10784 26630
rect 10808 26628 10864 26630
rect 10888 26628 10944 26630
rect 10968 26628 11024 26630
rect 10728 25594 10784 25596
rect 10808 25594 10864 25596
rect 10888 25594 10944 25596
rect 10968 25594 11024 25596
rect 10728 25542 10774 25594
rect 10774 25542 10784 25594
rect 10808 25542 10838 25594
rect 10838 25542 10850 25594
rect 10850 25542 10864 25594
rect 10888 25542 10902 25594
rect 10902 25542 10914 25594
rect 10914 25542 10944 25594
rect 10968 25542 10978 25594
rect 10978 25542 11024 25594
rect 10728 25540 10784 25542
rect 10808 25540 10864 25542
rect 10888 25540 10944 25542
rect 10968 25540 11024 25542
rect 10690 25200 10746 25256
rect 10322 24112 10378 24168
rect 10068 23962 10124 23964
rect 10148 23962 10204 23964
rect 10228 23962 10284 23964
rect 10308 23962 10364 23964
rect 10068 23910 10114 23962
rect 10114 23910 10124 23962
rect 10148 23910 10178 23962
rect 10178 23910 10190 23962
rect 10190 23910 10204 23962
rect 10228 23910 10242 23962
rect 10242 23910 10254 23962
rect 10254 23910 10284 23962
rect 10308 23910 10318 23962
rect 10318 23910 10364 23962
rect 10068 23908 10124 23910
rect 10148 23908 10204 23910
rect 10228 23908 10284 23910
rect 10308 23908 10364 23910
rect 9678 21936 9734 21992
rect 9586 21836 9588 21856
rect 9588 21836 9640 21856
rect 9640 21836 9642 21856
rect 9586 21800 9642 21836
rect 9678 21528 9734 21584
rect 9770 21256 9826 21312
rect 10322 23704 10378 23760
rect 10322 23432 10378 23488
rect 10138 23180 10194 23216
rect 10138 23160 10140 23180
rect 10140 23160 10192 23180
rect 10192 23160 10194 23180
rect 9954 23024 10010 23080
rect 10068 22874 10124 22876
rect 10148 22874 10204 22876
rect 10228 22874 10284 22876
rect 10308 22874 10364 22876
rect 10068 22822 10114 22874
rect 10114 22822 10124 22874
rect 10148 22822 10178 22874
rect 10178 22822 10190 22874
rect 10190 22822 10204 22874
rect 10228 22822 10242 22874
rect 10242 22822 10254 22874
rect 10254 22822 10284 22874
rect 10308 22822 10318 22874
rect 10318 22822 10364 22874
rect 10068 22820 10124 22822
rect 10148 22820 10204 22822
rect 10228 22820 10284 22822
rect 10308 22820 10364 22822
rect 10728 24506 10784 24508
rect 10808 24506 10864 24508
rect 10888 24506 10944 24508
rect 10968 24506 11024 24508
rect 10728 24454 10774 24506
rect 10774 24454 10784 24506
rect 10808 24454 10838 24506
rect 10838 24454 10850 24506
rect 10850 24454 10864 24506
rect 10888 24454 10902 24506
rect 10902 24454 10914 24506
rect 10914 24454 10944 24506
rect 10968 24454 10978 24506
rect 10978 24454 11024 24506
rect 10728 24452 10784 24454
rect 10808 24452 10864 24454
rect 10888 24452 10944 24454
rect 10968 24452 11024 24454
rect 10782 24248 10838 24304
rect 10966 24248 11022 24304
rect 10068 21786 10124 21788
rect 10148 21786 10204 21788
rect 10228 21786 10284 21788
rect 10308 21786 10364 21788
rect 10068 21734 10114 21786
rect 10114 21734 10124 21786
rect 10148 21734 10178 21786
rect 10178 21734 10190 21786
rect 10190 21734 10204 21786
rect 10228 21734 10242 21786
rect 10242 21734 10254 21786
rect 10254 21734 10284 21786
rect 10308 21734 10318 21786
rect 10318 21734 10364 21786
rect 10068 21732 10124 21734
rect 10148 21732 10204 21734
rect 10228 21732 10284 21734
rect 10308 21732 10364 21734
rect 8942 16904 8998 16960
rect 8850 15544 8906 15600
rect 8574 14864 8630 14920
rect 8482 14456 8538 14512
rect 8758 14728 8814 14784
rect 8482 12144 8538 12200
rect 8298 12008 8354 12064
rect 8298 11736 8354 11792
rect 8482 11756 8538 11792
rect 8482 11736 8484 11756
rect 8484 11736 8536 11756
rect 8536 11736 8538 11756
rect 8390 11600 8446 11656
rect 8942 13948 8944 13968
rect 8944 13948 8996 13968
rect 8996 13948 8998 13968
rect 8942 13912 8998 13948
rect 8850 11756 8906 11792
rect 8850 11736 8852 11756
rect 8852 11736 8904 11756
rect 8904 11736 8906 11756
rect 8022 3984 8078 4040
rect 8942 3984 8998 4040
rect 9126 16652 9182 16688
rect 9126 16632 9128 16652
rect 9128 16632 9180 16652
rect 9180 16632 9182 16652
rect 9678 18692 9734 18728
rect 9678 18672 9680 18692
rect 9680 18672 9732 18692
rect 9732 18672 9734 18692
rect 9310 17040 9366 17096
rect 9402 16496 9458 16552
rect 9218 15272 9274 15328
rect 9126 12980 9182 13016
rect 9126 12960 9128 12980
rect 9128 12960 9180 12980
rect 9180 12960 9182 12980
rect 9402 15020 9458 15056
rect 9402 15000 9404 15020
rect 9404 15000 9456 15020
rect 9456 15000 9458 15020
rect 9402 14456 9458 14512
rect 9678 17620 9680 17640
rect 9680 17620 9732 17640
rect 9732 17620 9734 17640
rect 9678 17584 9734 17620
rect 10138 20984 10194 21040
rect 10046 20884 10048 20904
rect 10048 20884 10100 20904
rect 10100 20884 10102 20904
rect 10046 20848 10102 20884
rect 10068 20698 10124 20700
rect 10148 20698 10204 20700
rect 10228 20698 10284 20700
rect 10308 20698 10364 20700
rect 10068 20646 10114 20698
rect 10114 20646 10124 20698
rect 10148 20646 10178 20698
rect 10178 20646 10190 20698
rect 10190 20646 10204 20698
rect 10228 20646 10242 20698
rect 10242 20646 10254 20698
rect 10254 20646 10284 20698
rect 10308 20646 10318 20698
rect 10318 20646 10364 20698
rect 10068 20644 10124 20646
rect 10148 20644 10204 20646
rect 10228 20644 10284 20646
rect 10308 20644 10364 20646
rect 10782 23976 10838 24032
rect 10728 23418 10784 23420
rect 10808 23418 10864 23420
rect 10888 23418 10944 23420
rect 10968 23418 11024 23420
rect 10728 23366 10774 23418
rect 10774 23366 10784 23418
rect 10808 23366 10838 23418
rect 10838 23366 10850 23418
rect 10850 23366 10864 23418
rect 10888 23366 10902 23418
rect 10902 23366 10914 23418
rect 10914 23366 10944 23418
rect 10968 23366 10978 23418
rect 10978 23366 11024 23418
rect 10728 23364 10784 23366
rect 10808 23364 10864 23366
rect 10888 23364 10944 23366
rect 10968 23364 11024 23366
rect 10690 23196 10692 23216
rect 10692 23196 10744 23216
rect 10744 23196 10746 23216
rect 10690 23160 10746 23196
rect 10728 22330 10784 22332
rect 10808 22330 10864 22332
rect 10888 22330 10944 22332
rect 10968 22330 11024 22332
rect 10728 22278 10774 22330
rect 10774 22278 10784 22330
rect 10808 22278 10838 22330
rect 10838 22278 10850 22330
rect 10850 22278 10864 22330
rect 10888 22278 10902 22330
rect 10902 22278 10914 22330
rect 10914 22278 10944 22330
rect 10968 22278 10978 22330
rect 10978 22278 11024 22330
rect 10728 22276 10784 22278
rect 10808 22276 10864 22278
rect 10888 22276 10944 22278
rect 10968 22276 11024 22278
rect 10598 21800 10654 21856
rect 10728 21242 10784 21244
rect 10808 21242 10864 21244
rect 10888 21242 10944 21244
rect 10968 21242 11024 21244
rect 10728 21190 10774 21242
rect 10774 21190 10784 21242
rect 10808 21190 10838 21242
rect 10838 21190 10850 21242
rect 10850 21190 10864 21242
rect 10888 21190 10902 21242
rect 10902 21190 10914 21242
rect 10914 21190 10944 21242
rect 10968 21190 10978 21242
rect 10978 21190 11024 21242
rect 10728 21188 10784 21190
rect 10808 21188 10864 21190
rect 10888 21188 10944 21190
rect 10968 21188 11024 21190
rect 10068 19610 10124 19612
rect 10148 19610 10204 19612
rect 10228 19610 10284 19612
rect 10308 19610 10364 19612
rect 10068 19558 10114 19610
rect 10114 19558 10124 19610
rect 10148 19558 10178 19610
rect 10178 19558 10190 19610
rect 10190 19558 10204 19610
rect 10228 19558 10242 19610
rect 10242 19558 10254 19610
rect 10254 19558 10284 19610
rect 10308 19558 10318 19610
rect 10318 19558 10364 19610
rect 10068 19556 10124 19558
rect 10148 19556 10204 19558
rect 10228 19556 10284 19558
rect 10308 19556 10364 19558
rect 10068 18522 10124 18524
rect 10148 18522 10204 18524
rect 10228 18522 10284 18524
rect 10308 18522 10364 18524
rect 10068 18470 10114 18522
rect 10114 18470 10124 18522
rect 10148 18470 10178 18522
rect 10178 18470 10190 18522
rect 10190 18470 10204 18522
rect 10228 18470 10242 18522
rect 10242 18470 10254 18522
rect 10254 18470 10284 18522
rect 10308 18470 10318 18522
rect 10318 18470 10364 18522
rect 10068 18468 10124 18470
rect 10148 18468 10204 18470
rect 10228 18468 10284 18470
rect 10308 18468 10364 18470
rect 10068 17434 10124 17436
rect 10148 17434 10204 17436
rect 10228 17434 10284 17436
rect 10308 17434 10364 17436
rect 10068 17382 10114 17434
rect 10114 17382 10124 17434
rect 10148 17382 10178 17434
rect 10178 17382 10190 17434
rect 10190 17382 10204 17434
rect 10228 17382 10242 17434
rect 10242 17382 10254 17434
rect 10254 17382 10284 17434
rect 10308 17382 10318 17434
rect 10318 17382 10364 17434
rect 10068 17380 10124 17382
rect 10148 17380 10204 17382
rect 10228 17380 10284 17382
rect 10308 17380 10364 17382
rect 9770 16904 9826 16960
rect 9678 16632 9734 16688
rect 9586 14728 9642 14784
rect 9494 13912 9550 13968
rect 9770 15680 9826 15736
rect 10690 20304 10746 20360
rect 10728 20154 10784 20156
rect 10808 20154 10864 20156
rect 10888 20154 10944 20156
rect 10968 20154 11024 20156
rect 10728 20102 10774 20154
rect 10774 20102 10784 20154
rect 10808 20102 10838 20154
rect 10838 20102 10850 20154
rect 10850 20102 10864 20154
rect 10888 20102 10902 20154
rect 10902 20102 10914 20154
rect 10914 20102 10944 20154
rect 10968 20102 10978 20154
rect 10978 20102 11024 20154
rect 10728 20100 10784 20102
rect 10808 20100 10864 20102
rect 10888 20100 10944 20102
rect 10968 20100 11024 20102
rect 10728 19066 10784 19068
rect 10808 19066 10864 19068
rect 10888 19066 10944 19068
rect 10968 19066 11024 19068
rect 10728 19014 10774 19066
rect 10774 19014 10784 19066
rect 10808 19014 10838 19066
rect 10838 19014 10850 19066
rect 10850 19014 10864 19066
rect 10888 19014 10902 19066
rect 10902 19014 10914 19066
rect 10914 19014 10944 19066
rect 10968 19014 10978 19066
rect 10978 19014 11024 19066
rect 10728 19012 10784 19014
rect 10808 19012 10864 19014
rect 10888 19012 10944 19014
rect 10968 19012 11024 19014
rect 10728 17978 10784 17980
rect 10808 17978 10864 17980
rect 10888 17978 10944 17980
rect 10968 17978 11024 17980
rect 10728 17926 10774 17978
rect 10774 17926 10784 17978
rect 10808 17926 10838 17978
rect 10838 17926 10850 17978
rect 10850 17926 10864 17978
rect 10888 17926 10902 17978
rect 10902 17926 10914 17978
rect 10914 17926 10944 17978
rect 10968 17926 10978 17978
rect 10978 17926 11024 17978
rect 10728 17924 10784 17926
rect 10808 17924 10864 17926
rect 10888 17924 10944 17926
rect 10968 17924 11024 17926
rect 10068 16346 10124 16348
rect 10148 16346 10204 16348
rect 10228 16346 10284 16348
rect 10308 16346 10364 16348
rect 10068 16294 10114 16346
rect 10114 16294 10124 16346
rect 10148 16294 10178 16346
rect 10178 16294 10190 16346
rect 10190 16294 10204 16346
rect 10228 16294 10242 16346
rect 10242 16294 10254 16346
rect 10254 16294 10284 16346
rect 10308 16294 10318 16346
rect 10318 16294 10364 16346
rect 10068 16292 10124 16294
rect 10148 16292 10204 16294
rect 10228 16292 10284 16294
rect 10308 16292 10364 16294
rect 10068 15258 10124 15260
rect 10148 15258 10204 15260
rect 10228 15258 10284 15260
rect 10308 15258 10364 15260
rect 10068 15206 10114 15258
rect 10114 15206 10124 15258
rect 10148 15206 10178 15258
rect 10178 15206 10190 15258
rect 10190 15206 10204 15258
rect 10228 15206 10242 15258
rect 10242 15206 10254 15258
rect 10254 15206 10284 15258
rect 10308 15206 10318 15258
rect 10318 15206 10364 15258
rect 10068 15204 10124 15206
rect 10148 15204 10204 15206
rect 10228 15204 10284 15206
rect 10308 15204 10364 15206
rect 9954 15000 10010 15056
rect 10728 16890 10784 16892
rect 10808 16890 10864 16892
rect 10888 16890 10944 16892
rect 10968 16890 11024 16892
rect 10728 16838 10774 16890
rect 10774 16838 10784 16890
rect 10808 16838 10838 16890
rect 10838 16838 10850 16890
rect 10850 16838 10864 16890
rect 10888 16838 10902 16890
rect 10902 16838 10914 16890
rect 10914 16838 10944 16890
rect 10968 16838 10978 16890
rect 10978 16838 11024 16890
rect 10728 16836 10784 16838
rect 10808 16836 10864 16838
rect 10888 16836 10944 16838
rect 10968 16836 11024 16838
rect 10068 14170 10124 14172
rect 10148 14170 10204 14172
rect 10228 14170 10284 14172
rect 10308 14170 10364 14172
rect 10068 14118 10114 14170
rect 10114 14118 10124 14170
rect 10148 14118 10178 14170
rect 10178 14118 10190 14170
rect 10190 14118 10204 14170
rect 10228 14118 10242 14170
rect 10242 14118 10254 14170
rect 10254 14118 10284 14170
rect 10308 14118 10318 14170
rect 10318 14118 10364 14170
rect 10068 14116 10124 14118
rect 10148 14116 10204 14118
rect 10228 14116 10284 14118
rect 10308 14116 10364 14118
rect 10068 13082 10124 13084
rect 10148 13082 10204 13084
rect 10228 13082 10284 13084
rect 10308 13082 10364 13084
rect 10068 13030 10114 13082
rect 10114 13030 10124 13082
rect 10148 13030 10178 13082
rect 10178 13030 10190 13082
rect 10190 13030 10204 13082
rect 10228 13030 10242 13082
rect 10242 13030 10254 13082
rect 10254 13030 10284 13082
rect 10308 13030 10318 13082
rect 10318 13030 10364 13082
rect 10068 13028 10124 13030
rect 10148 13028 10204 13030
rect 10228 13028 10284 13030
rect 10308 13028 10364 13030
rect 10068 11994 10124 11996
rect 10148 11994 10204 11996
rect 10228 11994 10284 11996
rect 10308 11994 10364 11996
rect 10068 11942 10114 11994
rect 10114 11942 10124 11994
rect 10148 11942 10178 11994
rect 10178 11942 10190 11994
rect 10190 11942 10204 11994
rect 10228 11942 10242 11994
rect 10242 11942 10254 11994
rect 10254 11942 10284 11994
rect 10308 11942 10318 11994
rect 10318 11942 10364 11994
rect 10068 11940 10124 11942
rect 10148 11940 10204 11942
rect 10228 11940 10284 11942
rect 10308 11940 10364 11942
rect 9218 9424 9274 9480
rect 10068 10906 10124 10908
rect 10148 10906 10204 10908
rect 10228 10906 10284 10908
rect 10308 10906 10364 10908
rect 10068 10854 10114 10906
rect 10114 10854 10124 10906
rect 10148 10854 10178 10906
rect 10178 10854 10190 10906
rect 10190 10854 10204 10906
rect 10228 10854 10242 10906
rect 10242 10854 10254 10906
rect 10254 10854 10284 10906
rect 10308 10854 10318 10906
rect 10318 10854 10364 10906
rect 10068 10852 10124 10854
rect 10148 10852 10204 10854
rect 10228 10852 10284 10854
rect 10308 10852 10364 10854
rect 11242 29144 11298 29200
rect 11242 26560 11298 26616
rect 11242 19216 11298 19272
rect 11150 18264 11206 18320
rect 10728 15802 10784 15804
rect 10808 15802 10864 15804
rect 10888 15802 10944 15804
rect 10968 15802 11024 15804
rect 10728 15750 10774 15802
rect 10774 15750 10784 15802
rect 10808 15750 10838 15802
rect 10838 15750 10850 15802
rect 10850 15750 10864 15802
rect 10888 15750 10902 15802
rect 10902 15750 10914 15802
rect 10914 15750 10944 15802
rect 10968 15750 10978 15802
rect 10978 15750 11024 15802
rect 10728 15748 10784 15750
rect 10808 15748 10864 15750
rect 10888 15748 10944 15750
rect 10968 15748 11024 15750
rect 10728 14714 10784 14716
rect 10808 14714 10864 14716
rect 10888 14714 10944 14716
rect 10968 14714 11024 14716
rect 10728 14662 10774 14714
rect 10774 14662 10784 14714
rect 10808 14662 10838 14714
rect 10838 14662 10850 14714
rect 10850 14662 10864 14714
rect 10888 14662 10902 14714
rect 10902 14662 10914 14714
rect 10914 14662 10944 14714
rect 10968 14662 10978 14714
rect 10978 14662 11024 14714
rect 10728 14660 10784 14662
rect 10808 14660 10864 14662
rect 10888 14660 10944 14662
rect 10968 14660 11024 14662
rect 10728 13626 10784 13628
rect 10808 13626 10864 13628
rect 10888 13626 10944 13628
rect 10968 13626 11024 13628
rect 10728 13574 10774 13626
rect 10774 13574 10784 13626
rect 10808 13574 10838 13626
rect 10838 13574 10850 13626
rect 10850 13574 10864 13626
rect 10888 13574 10902 13626
rect 10902 13574 10914 13626
rect 10914 13574 10944 13626
rect 10968 13574 10978 13626
rect 10978 13574 11024 13626
rect 10728 13572 10784 13574
rect 10808 13572 10864 13574
rect 10888 13572 10944 13574
rect 10968 13572 11024 13574
rect 10728 12538 10784 12540
rect 10808 12538 10864 12540
rect 10888 12538 10944 12540
rect 10968 12538 11024 12540
rect 10728 12486 10774 12538
rect 10774 12486 10784 12538
rect 10808 12486 10838 12538
rect 10838 12486 10850 12538
rect 10850 12486 10864 12538
rect 10888 12486 10902 12538
rect 10902 12486 10914 12538
rect 10914 12486 10944 12538
rect 10968 12486 10978 12538
rect 10978 12486 11024 12538
rect 10728 12484 10784 12486
rect 10808 12484 10864 12486
rect 10888 12484 10944 12486
rect 10968 12484 11024 12486
rect 11242 16496 11298 16552
rect 10728 11450 10784 11452
rect 10808 11450 10864 11452
rect 10888 11450 10944 11452
rect 10968 11450 11024 11452
rect 10728 11398 10774 11450
rect 10774 11398 10784 11450
rect 10808 11398 10838 11450
rect 10838 11398 10850 11450
rect 10850 11398 10864 11450
rect 10888 11398 10902 11450
rect 10902 11398 10914 11450
rect 10914 11398 10944 11450
rect 10968 11398 10978 11450
rect 10978 11398 11024 11450
rect 10728 11396 10784 11398
rect 10808 11396 10864 11398
rect 10888 11396 10944 11398
rect 10968 11396 11024 11398
rect 10728 10362 10784 10364
rect 10808 10362 10864 10364
rect 10888 10362 10944 10364
rect 10968 10362 11024 10364
rect 10728 10310 10774 10362
rect 10774 10310 10784 10362
rect 10808 10310 10838 10362
rect 10838 10310 10850 10362
rect 10850 10310 10864 10362
rect 10888 10310 10902 10362
rect 10902 10310 10914 10362
rect 10914 10310 10944 10362
rect 10968 10310 10978 10362
rect 10978 10310 11024 10362
rect 10728 10308 10784 10310
rect 10808 10308 10864 10310
rect 10888 10308 10944 10310
rect 10968 10308 11024 10310
rect 10068 9818 10124 9820
rect 10148 9818 10204 9820
rect 10228 9818 10284 9820
rect 10308 9818 10364 9820
rect 10068 9766 10114 9818
rect 10114 9766 10124 9818
rect 10148 9766 10178 9818
rect 10178 9766 10190 9818
rect 10190 9766 10204 9818
rect 10228 9766 10242 9818
rect 10242 9766 10254 9818
rect 10254 9766 10284 9818
rect 10308 9766 10318 9818
rect 10318 9766 10364 9818
rect 10068 9764 10124 9766
rect 10148 9764 10204 9766
rect 10228 9764 10284 9766
rect 10308 9764 10364 9766
rect 10068 8730 10124 8732
rect 10148 8730 10204 8732
rect 10228 8730 10284 8732
rect 10308 8730 10364 8732
rect 10068 8678 10114 8730
rect 10114 8678 10124 8730
rect 10148 8678 10178 8730
rect 10178 8678 10190 8730
rect 10190 8678 10204 8730
rect 10228 8678 10242 8730
rect 10242 8678 10254 8730
rect 10254 8678 10284 8730
rect 10308 8678 10318 8730
rect 10318 8678 10364 8730
rect 10068 8676 10124 8678
rect 10148 8676 10204 8678
rect 10228 8676 10284 8678
rect 10308 8676 10364 8678
rect 10728 9274 10784 9276
rect 10808 9274 10864 9276
rect 10888 9274 10944 9276
rect 10968 9274 11024 9276
rect 10728 9222 10774 9274
rect 10774 9222 10784 9274
rect 10808 9222 10838 9274
rect 10838 9222 10850 9274
rect 10850 9222 10864 9274
rect 10888 9222 10902 9274
rect 10902 9222 10914 9274
rect 10914 9222 10944 9274
rect 10968 9222 10978 9274
rect 10978 9222 11024 9274
rect 10728 9220 10784 9222
rect 10808 9220 10864 9222
rect 10888 9220 10944 9222
rect 10968 9220 11024 9222
rect 10068 7642 10124 7644
rect 10148 7642 10204 7644
rect 10228 7642 10284 7644
rect 10308 7642 10364 7644
rect 10068 7590 10114 7642
rect 10114 7590 10124 7642
rect 10148 7590 10178 7642
rect 10178 7590 10190 7642
rect 10190 7590 10204 7642
rect 10228 7590 10242 7642
rect 10242 7590 10254 7642
rect 10254 7590 10284 7642
rect 10308 7590 10318 7642
rect 10318 7590 10364 7642
rect 10068 7588 10124 7590
rect 10148 7588 10204 7590
rect 10228 7588 10284 7590
rect 10308 7588 10364 7590
rect 10728 8186 10784 8188
rect 10808 8186 10864 8188
rect 10888 8186 10944 8188
rect 10968 8186 11024 8188
rect 10728 8134 10774 8186
rect 10774 8134 10784 8186
rect 10808 8134 10838 8186
rect 10838 8134 10850 8186
rect 10850 8134 10864 8186
rect 10888 8134 10902 8186
rect 10902 8134 10914 8186
rect 10914 8134 10944 8186
rect 10968 8134 10978 8186
rect 10978 8134 11024 8186
rect 10728 8132 10784 8134
rect 10808 8132 10864 8134
rect 10888 8132 10944 8134
rect 10968 8132 11024 8134
rect 9126 3732 9182 3768
rect 9126 3712 9128 3732
rect 9128 3712 9180 3732
rect 9180 3712 9182 3732
rect 10068 6554 10124 6556
rect 10148 6554 10204 6556
rect 10228 6554 10284 6556
rect 10308 6554 10364 6556
rect 10068 6502 10114 6554
rect 10114 6502 10124 6554
rect 10148 6502 10178 6554
rect 10178 6502 10190 6554
rect 10190 6502 10204 6554
rect 10228 6502 10242 6554
rect 10242 6502 10254 6554
rect 10254 6502 10284 6554
rect 10308 6502 10318 6554
rect 10318 6502 10364 6554
rect 10068 6500 10124 6502
rect 10148 6500 10204 6502
rect 10228 6500 10284 6502
rect 10308 6500 10364 6502
rect 10068 5466 10124 5468
rect 10148 5466 10204 5468
rect 10228 5466 10284 5468
rect 10308 5466 10364 5468
rect 10068 5414 10114 5466
rect 10114 5414 10124 5466
rect 10148 5414 10178 5466
rect 10178 5414 10190 5466
rect 10190 5414 10204 5466
rect 10228 5414 10242 5466
rect 10242 5414 10254 5466
rect 10254 5414 10284 5466
rect 10308 5414 10318 5466
rect 10318 5414 10364 5466
rect 10068 5412 10124 5414
rect 10148 5412 10204 5414
rect 10228 5412 10284 5414
rect 10308 5412 10364 5414
rect 10068 4378 10124 4380
rect 10148 4378 10204 4380
rect 10228 4378 10284 4380
rect 10308 4378 10364 4380
rect 10068 4326 10114 4378
rect 10114 4326 10124 4378
rect 10148 4326 10178 4378
rect 10178 4326 10190 4378
rect 10190 4326 10204 4378
rect 10228 4326 10242 4378
rect 10242 4326 10254 4378
rect 10254 4326 10284 4378
rect 10308 4326 10318 4378
rect 10318 4326 10364 4378
rect 10068 4324 10124 4326
rect 10148 4324 10204 4326
rect 10228 4324 10284 4326
rect 10308 4324 10364 4326
rect 10728 7098 10784 7100
rect 10808 7098 10864 7100
rect 10888 7098 10944 7100
rect 10968 7098 11024 7100
rect 10728 7046 10774 7098
rect 10774 7046 10784 7098
rect 10808 7046 10838 7098
rect 10838 7046 10850 7098
rect 10850 7046 10864 7098
rect 10888 7046 10902 7098
rect 10902 7046 10914 7098
rect 10914 7046 10944 7098
rect 10968 7046 10978 7098
rect 10978 7046 11024 7098
rect 10728 7044 10784 7046
rect 10808 7044 10864 7046
rect 10888 7044 10944 7046
rect 10968 7044 11024 7046
rect 10728 6010 10784 6012
rect 10808 6010 10864 6012
rect 10888 6010 10944 6012
rect 10968 6010 11024 6012
rect 10728 5958 10774 6010
rect 10774 5958 10784 6010
rect 10808 5958 10838 6010
rect 10838 5958 10850 6010
rect 10850 5958 10864 6010
rect 10888 5958 10902 6010
rect 10902 5958 10914 6010
rect 10914 5958 10944 6010
rect 10968 5958 10978 6010
rect 10978 5958 11024 6010
rect 10728 5956 10784 5958
rect 10808 5956 10864 5958
rect 10888 5956 10944 5958
rect 10968 5956 11024 5958
rect 10728 4922 10784 4924
rect 10808 4922 10864 4924
rect 10888 4922 10944 4924
rect 10968 4922 11024 4924
rect 10728 4870 10774 4922
rect 10774 4870 10784 4922
rect 10808 4870 10838 4922
rect 10838 4870 10850 4922
rect 10850 4870 10864 4922
rect 10888 4870 10902 4922
rect 10902 4870 10914 4922
rect 10914 4870 10944 4922
rect 10968 4870 10978 4922
rect 10978 4870 11024 4922
rect 10728 4868 10784 4870
rect 10808 4868 10864 4870
rect 10888 4868 10944 4870
rect 10968 4868 11024 4870
rect 10068 3290 10124 3292
rect 10148 3290 10204 3292
rect 10228 3290 10284 3292
rect 10308 3290 10364 3292
rect 10068 3238 10114 3290
rect 10114 3238 10124 3290
rect 10148 3238 10178 3290
rect 10178 3238 10190 3290
rect 10190 3238 10204 3290
rect 10228 3238 10242 3290
rect 10242 3238 10254 3290
rect 10254 3238 10284 3290
rect 10308 3238 10318 3290
rect 10318 3238 10364 3290
rect 10068 3236 10124 3238
rect 10148 3236 10204 3238
rect 10228 3236 10284 3238
rect 10308 3236 10364 3238
rect 10728 3834 10784 3836
rect 10808 3834 10864 3836
rect 10888 3834 10944 3836
rect 10968 3834 11024 3836
rect 10728 3782 10774 3834
rect 10774 3782 10784 3834
rect 10808 3782 10838 3834
rect 10838 3782 10850 3834
rect 10850 3782 10864 3834
rect 10888 3782 10902 3834
rect 10902 3782 10914 3834
rect 10914 3782 10944 3834
rect 10968 3782 10978 3834
rect 10978 3782 11024 3834
rect 10728 3780 10784 3782
rect 10808 3780 10864 3782
rect 10888 3780 10944 3782
rect 10968 3780 11024 3782
rect 10728 2746 10784 2748
rect 10808 2746 10864 2748
rect 10888 2746 10944 2748
rect 10968 2746 11024 2748
rect 10728 2694 10774 2746
rect 10774 2694 10784 2746
rect 10808 2694 10838 2746
rect 10838 2694 10850 2746
rect 10850 2694 10864 2746
rect 10888 2694 10902 2746
rect 10902 2694 10914 2746
rect 10914 2694 10944 2746
rect 10968 2694 10978 2746
rect 10978 2694 11024 2746
rect 10728 2692 10784 2694
rect 10808 2692 10864 2694
rect 10888 2692 10944 2694
rect 10968 2692 11024 2694
rect 10068 2202 10124 2204
rect 10148 2202 10204 2204
rect 10228 2202 10284 2204
rect 10308 2202 10364 2204
rect 10068 2150 10114 2202
rect 10114 2150 10124 2202
rect 10148 2150 10178 2202
rect 10178 2150 10190 2202
rect 10190 2150 10204 2202
rect 10228 2150 10242 2202
rect 10242 2150 10254 2202
rect 10254 2150 10284 2202
rect 10308 2150 10318 2202
rect 10318 2150 10364 2202
rect 10068 2148 10124 2150
rect 10148 2148 10204 2150
rect 10228 2148 10284 2150
rect 10308 2148 10364 2150
rect 10728 1658 10784 1660
rect 10808 1658 10864 1660
rect 10888 1658 10944 1660
rect 10968 1658 11024 1660
rect 10728 1606 10774 1658
rect 10774 1606 10784 1658
rect 10808 1606 10838 1658
rect 10838 1606 10850 1658
rect 10850 1606 10864 1658
rect 10888 1606 10902 1658
rect 10902 1606 10914 1658
rect 10914 1606 10944 1658
rect 10968 1606 10978 1658
rect 10978 1606 11024 1658
rect 10728 1604 10784 1606
rect 10808 1604 10864 1606
rect 10888 1604 10944 1606
rect 10968 1604 11024 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 10068 1114 10124 1116
rect 10148 1114 10204 1116
rect 10228 1114 10284 1116
rect 10308 1114 10364 1116
rect 10068 1062 10114 1114
rect 10114 1062 10124 1114
rect 10148 1062 10178 1114
rect 10178 1062 10190 1114
rect 10190 1062 10204 1114
rect 10228 1062 10242 1114
rect 10242 1062 10254 1114
rect 10254 1062 10284 1114
rect 10308 1062 10318 1114
rect 10318 1062 10364 1114
rect 10068 1060 10124 1062
rect 10148 1060 10204 1062
rect 10228 1060 10284 1062
rect 10308 1060 10364 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
rect 10728 570 10784 572
rect 10808 570 10864 572
rect 10888 570 10944 572
rect 10968 570 11024 572
rect 10728 518 10774 570
rect 10774 518 10784 570
rect 10808 518 10838 570
rect 10838 518 10850 570
rect 10850 518 10864 570
rect 10888 518 10902 570
rect 10902 518 10914 570
rect 10914 518 10944 570
rect 10968 518 10978 570
rect 10978 518 11024 570
rect 10728 516 10784 518
rect 10808 516 10864 518
rect 10888 516 10944 518
rect 10968 516 11024 518
<< metal3 >>
rect 974 43556 980 43620
rect 1044 43618 1050 43620
rect 1117 43618 1183 43621
rect 1044 43616 1183 43618
rect 1044 43560 1122 43616
rect 1178 43560 1183 43616
rect 1044 43558 1183 43560
rect 1044 43556 1050 43558
rect 1117 43555 1183 43558
rect 7741 43620 7807 43621
rect 7741 43616 7788 43620
rect 7852 43618 7858 43620
rect 7741 43560 7746 43616
rect 7741 43556 7788 43560
rect 7852 43558 7898 43618
rect 7852 43556 7858 43558
rect 7741 43555 7807 43556
rect 4318 43008 4634 43009
rect 4318 42944 4324 43008
rect 4388 42944 4404 43008
rect 4468 42944 4484 43008
rect 4548 42944 4564 43008
rect 4628 42944 4634 43008
rect 4318 42943 4634 42944
rect 10718 43008 11034 43009
rect 10718 42944 10724 43008
rect 10788 42944 10804 43008
rect 10868 42944 10884 43008
rect 10948 42944 10964 43008
rect 11028 42944 11034 43008
rect 10718 42943 11034 42944
rect 3658 42464 3974 42465
rect 3658 42400 3664 42464
rect 3728 42400 3744 42464
rect 3808 42400 3824 42464
rect 3888 42400 3904 42464
rect 3968 42400 3974 42464
rect 3658 42399 3974 42400
rect 10058 42464 10374 42465
rect 10058 42400 10064 42464
rect 10128 42400 10144 42464
rect 10208 42400 10224 42464
rect 10288 42400 10304 42464
rect 10368 42400 10374 42464
rect 10058 42399 10374 42400
rect 5574 42196 5580 42260
rect 5644 42258 5650 42260
rect 5809 42258 5875 42261
rect 5644 42256 5875 42258
rect 5644 42200 5814 42256
rect 5870 42200 5875 42256
rect 5644 42198 5875 42200
rect 5644 42196 5650 42198
rect 5809 42195 5875 42198
rect 4337 42122 4403 42125
rect 5206 42122 5212 42124
rect 4337 42120 5212 42122
rect 4337 42064 4342 42120
rect 4398 42064 5212 42120
rect 4337 42062 5212 42064
rect 4337 42059 4403 42062
rect 5206 42060 5212 42062
rect 5276 42060 5282 42124
rect 4318 41920 4634 41921
rect 4318 41856 4324 41920
rect 4388 41856 4404 41920
rect 4468 41856 4484 41920
rect 4548 41856 4564 41920
rect 4628 41856 4634 41920
rect 4318 41855 4634 41856
rect 10718 41920 11034 41921
rect 10718 41856 10724 41920
rect 10788 41856 10804 41920
rect 10868 41856 10884 41920
rect 10948 41856 10964 41920
rect 11028 41856 11034 41920
rect 10718 41855 11034 41856
rect 0 41717 400 41744
rect 0 41712 447 41717
rect 6637 41716 6703 41717
rect 6637 41714 6684 41716
rect 0 41656 386 41712
rect 442 41656 447 41712
rect 0 41651 447 41656
rect 6592 41712 6684 41714
rect 6592 41656 6642 41712
rect 6592 41654 6684 41656
rect 6637 41652 6684 41654
rect 6748 41652 6754 41716
rect 6637 41651 6703 41652
rect 0 41624 400 41651
rect 1117 41580 1183 41581
rect 1117 41576 1164 41580
rect 1228 41578 1234 41580
rect 7741 41578 7807 41581
rect 1117 41520 1122 41576
rect 1117 41516 1164 41520
rect 1228 41518 1274 41578
rect 3374 41576 7807 41578
rect 3374 41520 7746 41576
rect 7802 41520 7807 41576
rect 3374 41518 7807 41520
rect 1228 41516 1234 41518
rect 1117 41515 1183 41516
rect 0 41442 400 41472
rect 657 41442 723 41445
rect 0 41440 723 41442
rect 0 41384 662 41440
rect 718 41384 723 41440
rect 0 41382 723 41384
rect 0 41352 400 41382
rect 657 41379 723 41382
rect 1117 41442 1183 41445
rect 3374 41442 3434 41518
rect 7741 41515 7807 41518
rect 8017 41578 8083 41581
rect 8753 41578 8819 41581
rect 8017 41576 8819 41578
rect 8017 41520 8022 41576
rect 8078 41520 8758 41576
rect 8814 41520 8819 41576
rect 8017 41518 8819 41520
rect 8017 41515 8083 41518
rect 8753 41515 8819 41518
rect 1117 41440 3434 41442
rect 1117 41384 1122 41440
rect 1178 41384 3434 41440
rect 1117 41382 3434 41384
rect 7557 41442 7623 41445
rect 7966 41442 7972 41444
rect 7557 41440 7972 41442
rect 7557 41384 7562 41440
rect 7618 41384 7972 41440
rect 7557 41382 7972 41384
rect 1117 41379 1183 41382
rect 7557 41379 7623 41382
rect 7966 41380 7972 41382
rect 8036 41380 8042 41444
rect 3658 41376 3974 41377
rect 3658 41312 3664 41376
rect 3728 41312 3744 41376
rect 3808 41312 3824 41376
rect 3888 41312 3904 41376
rect 3968 41312 3974 41376
rect 3658 41311 3974 41312
rect 10058 41376 10374 41377
rect 10058 41312 10064 41376
rect 10128 41312 10144 41376
rect 10208 41312 10224 41376
rect 10288 41312 10304 41376
rect 10368 41312 10374 41376
rect 10058 41311 10374 41312
rect 7465 41306 7531 41309
rect 8385 41306 8451 41309
rect 8753 41306 8819 41309
rect 7465 41304 8451 41306
rect 7465 41248 7470 41304
rect 7526 41248 8390 41304
rect 8446 41248 8451 41304
rect 7465 41246 8451 41248
rect 7465 41243 7531 41246
rect 8385 41243 8451 41246
rect 8526 41304 8819 41306
rect 8526 41248 8758 41304
rect 8814 41248 8819 41304
rect 8526 41246 8819 41248
rect 0 41170 400 41200
rect 2129 41170 2195 41173
rect 0 41168 2195 41170
rect 0 41112 2134 41168
rect 2190 41112 2195 41168
rect 0 41110 2195 41112
rect 0 41080 400 41110
rect 2129 41107 2195 41110
rect 2630 41108 2636 41172
rect 2700 41170 2706 41172
rect 8293 41170 8359 41173
rect 2700 41168 8359 41170
rect 2700 41112 8298 41168
rect 8354 41112 8359 41168
rect 2700 41110 8359 41112
rect 2700 41108 2706 41110
rect 8293 41107 8359 41110
rect 3366 40972 3372 41036
rect 3436 41034 3442 41036
rect 8526 41034 8586 41246
rect 8753 41243 8819 41246
rect 3436 40974 8586 41034
rect 3436 40972 3442 40974
rect 0 40898 400 40928
rect 3049 40898 3115 40901
rect 0 40896 3115 40898
rect 0 40840 3054 40896
rect 3110 40840 3115 40896
rect 0 40838 3115 40840
rect 0 40808 400 40838
rect 3049 40835 3115 40838
rect 4318 40832 4634 40833
rect 4318 40768 4324 40832
rect 4388 40768 4404 40832
rect 4468 40768 4484 40832
rect 4548 40768 4564 40832
rect 4628 40768 4634 40832
rect 4318 40767 4634 40768
rect 10718 40832 11034 40833
rect 10718 40768 10724 40832
rect 10788 40768 10804 40832
rect 10868 40768 10884 40832
rect 10948 40768 10964 40832
rect 11028 40768 11034 40832
rect 10718 40767 11034 40768
rect 8293 40760 8359 40765
rect 8293 40704 8298 40760
rect 8354 40704 8359 40760
rect 8293 40699 8359 40704
rect 0 40626 400 40656
rect 841 40626 907 40629
rect 0 40624 907 40626
rect 0 40568 846 40624
rect 902 40568 907 40624
rect 0 40566 907 40568
rect 8296 40626 8356 40699
rect 8661 40626 8727 40629
rect 9489 40626 9555 40629
rect 8296 40624 9555 40626
rect 8296 40568 8666 40624
rect 8722 40568 9494 40624
rect 9550 40568 9555 40624
rect 8296 40566 9555 40568
rect 0 40536 400 40566
rect 841 40563 907 40566
rect 8661 40563 8727 40566
rect 9489 40563 9555 40566
rect 1301 40490 1367 40493
rect 1853 40490 1919 40493
rect 2221 40490 2287 40493
rect 1301 40488 1410 40490
rect 1301 40432 1306 40488
rect 1362 40432 1410 40488
rect 1301 40427 1410 40432
rect 1853 40488 2287 40490
rect 1853 40432 1858 40488
rect 1914 40432 2226 40488
rect 2282 40432 2287 40488
rect 1853 40430 2287 40432
rect 1853 40427 1919 40430
rect 2221 40427 2287 40430
rect 0 40354 400 40384
rect 565 40354 631 40357
rect 0 40352 631 40354
rect 0 40296 570 40352
rect 626 40296 631 40352
rect 0 40294 631 40296
rect 0 40264 400 40294
rect 565 40291 631 40294
rect 0 40082 400 40112
rect 1025 40082 1091 40085
rect 0 40080 1091 40082
rect 0 40024 1030 40080
rect 1086 40024 1091 40080
rect 0 40022 1091 40024
rect 0 39992 400 40022
rect 1025 40019 1091 40022
rect 1350 39946 1410 40427
rect 3658 40288 3974 40289
rect 3658 40224 3664 40288
rect 3728 40224 3744 40288
rect 3808 40224 3824 40288
rect 3888 40224 3904 40288
rect 3968 40224 3974 40288
rect 3658 40223 3974 40224
rect 10058 40288 10374 40289
rect 10058 40224 10064 40288
rect 10128 40224 10144 40288
rect 10208 40224 10224 40288
rect 10288 40224 10304 40288
rect 10368 40224 10374 40288
rect 10058 40223 10374 40224
rect 1894 40156 1900 40220
rect 1964 40218 1970 40220
rect 2957 40218 3023 40221
rect 1964 40216 3023 40218
rect 1964 40160 2962 40216
rect 3018 40160 3023 40216
rect 1964 40158 3023 40160
rect 1964 40156 1970 40158
rect 2957 40155 3023 40158
rect 4838 40156 4844 40220
rect 4908 40218 4914 40220
rect 8753 40218 8819 40221
rect 4908 40216 8819 40218
rect 4908 40160 8758 40216
rect 8814 40160 8819 40216
rect 4908 40158 8819 40160
rect 4908 40156 4914 40158
rect 8753 40155 8819 40158
rect 4102 40020 4108 40084
rect 4172 40082 4178 40084
rect 5257 40082 5323 40085
rect 4172 40080 5323 40082
rect 4172 40024 5262 40080
rect 5318 40024 5323 40080
rect 4172 40022 5323 40024
rect 4172 40020 4178 40022
rect 5257 40019 5323 40022
rect 5942 40020 5948 40084
rect 6012 40082 6018 40084
rect 6177 40082 6243 40085
rect 6012 40080 6243 40082
rect 6012 40024 6182 40080
rect 6238 40024 6243 40080
rect 6012 40022 6243 40024
rect 6012 40020 6018 40022
rect 6177 40019 6243 40022
rect 6494 40020 6500 40084
rect 6564 40082 6570 40084
rect 6637 40082 6703 40085
rect 6564 40080 6703 40082
rect 6564 40024 6642 40080
rect 6698 40024 6703 40080
rect 6564 40022 6703 40024
rect 6564 40020 6570 40022
rect 6637 40019 6703 40022
rect 8753 40082 8819 40085
rect 10685 40082 10751 40085
rect 8753 40080 10751 40082
rect 8753 40024 8758 40080
rect 8814 40024 10690 40080
rect 10746 40024 10751 40080
rect 8753 40022 10751 40024
rect 8753 40019 8819 40022
rect 10685 40019 10751 40022
rect 2078 39946 2084 39948
rect 1350 39886 2084 39946
rect 2078 39884 2084 39886
rect 2148 39884 2154 39948
rect 3601 39946 3667 39949
rect 6269 39946 6335 39949
rect 3601 39944 6335 39946
rect 3601 39888 3606 39944
rect 3662 39888 6274 39944
rect 6330 39888 6335 39944
rect 3601 39886 6335 39888
rect 3601 39883 3667 39886
rect 6269 39883 6335 39886
rect 8109 39946 8175 39949
rect 10685 39946 10751 39949
rect 8109 39944 10751 39946
rect 8109 39888 8114 39944
rect 8170 39888 10690 39944
rect 10746 39888 10751 39944
rect 8109 39886 10751 39888
rect 8109 39883 8175 39886
rect 10685 39883 10751 39886
rect 0 39810 400 39840
rect 1301 39810 1367 39813
rect 0 39808 1367 39810
rect 0 39752 1306 39808
rect 1362 39752 1367 39808
rect 0 39750 1367 39752
rect 0 39720 400 39750
rect 1301 39747 1367 39750
rect 5993 39810 6059 39813
rect 8753 39810 8819 39813
rect 5993 39808 8819 39810
rect 5993 39752 5998 39808
rect 6054 39752 8758 39808
rect 8814 39752 8819 39808
rect 5993 39750 8819 39752
rect 5993 39747 6059 39750
rect 8753 39747 8819 39750
rect 4318 39744 4634 39745
rect 4318 39680 4324 39744
rect 4388 39680 4404 39744
rect 4468 39680 4484 39744
rect 4548 39680 4564 39744
rect 4628 39680 4634 39744
rect 4318 39679 4634 39680
rect 10718 39744 11034 39745
rect 10718 39680 10724 39744
rect 10788 39680 10804 39744
rect 10868 39680 10884 39744
rect 10948 39680 10964 39744
rect 11028 39680 11034 39744
rect 10718 39679 11034 39680
rect 1485 39674 1551 39677
rect 2589 39674 2655 39677
rect 1485 39672 2655 39674
rect 1485 39616 1490 39672
rect 1546 39616 2594 39672
rect 2650 39616 2655 39672
rect 1485 39614 2655 39616
rect 1485 39611 1551 39614
rect 2589 39611 2655 39614
rect 8661 39674 8727 39677
rect 9438 39674 9444 39676
rect 8661 39672 9444 39674
rect 8661 39616 8666 39672
rect 8722 39616 9444 39672
rect 8661 39614 9444 39616
rect 8661 39611 8727 39614
rect 9438 39612 9444 39614
rect 9508 39612 9514 39676
rect 0 39538 400 39568
rect 933 39538 999 39541
rect 0 39536 999 39538
rect 0 39480 938 39536
rect 994 39480 999 39536
rect 0 39478 999 39480
rect 0 39448 400 39478
rect 933 39475 999 39478
rect 1301 39538 1367 39541
rect 4889 39538 4955 39541
rect 1301 39536 4955 39538
rect 1301 39480 1306 39536
rect 1362 39480 4894 39536
rect 4950 39480 4955 39536
rect 1301 39478 4955 39480
rect 1301 39475 1367 39478
rect 4889 39475 4955 39478
rect 8334 39476 8340 39540
rect 8404 39538 8410 39540
rect 10225 39538 10291 39541
rect 8404 39536 10291 39538
rect 8404 39480 10230 39536
rect 10286 39480 10291 39536
rect 8404 39478 10291 39480
rect 8404 39476 8410 39478
rect 10225 39475 10291 39478
rect 2078 39340 2084 39404
rect 2148 39402 2154 39404
rect 6821 39402 6887 39405
rect 2148 39400 6887 39402
rect 2148 39344 6826 39400
rect 6882 39344 6887 39400
rect 2148 39342 6887 39344
rect 2148 39340 2154 39342
rect 6821 39339 6887 39342
rect 7598 39340 7604 39404
rect 7668 39402 7674 39404
rect 10133 39402 10199 39405
rect 7668 39400 10199 39402
rect 7668 39344 10138 39400
rect 10194 39344 10199 39400
rect 7668 39342 10199 39344
rect 7668 39340 7674 39342
rect 10133 39339 10199 39342
rect 0 39266 400 39296
rect 1117 39266 1183 39269
rect 0 39264 1183 39266
rect 0 39208 1122 39264
rect 1178 39208 1183 39264
rect 0 39206 1183 39208
rect 0 39176 400 39206
rect 1117 39203 1183 39206
rect 3658 39200 3974 39201
rect 3658 39136 3664 39200
rect 3728 39136 3744 39200
rect 3808 39136 3824 39200
rect 3888 39136 3904 39200
rect 3968 39136 3974 39200
rect 3658 39135 3974 39136
rect 10058 39200 10374 39201
rect 10058 39136 10064 39200
rect 10128 39136 10144 39200
rect 10208 39136 10224 39200
rect 10288 39136 10304 39200
rect 10368 39136 10374 39200
rect 10058 39135 10374 39136
rect 7649 39130 7715 39133
rect 8385 39130 8451 39133
rect 7649 39128 8451 39130
rect 7649 39072 7654 39128
rect 7710 39072 8390 39128
rect 8446 39072 8451 39128
rect 7649 39070 8451 39072
rect 7649 39067 7715 39070
rect 8385 39067 8451 39070
rect 2773 38994 2839 38997
rect 7281 38994 7347 38997
rect 7557 38994 7623 38997
rect 2773 38992 7623 38994
rect 2773 38936 2778 38992
rect 2834 38936 7286 38992
rect 7342 38936 7562 38992
rect 7618 38936 7623 38992
rect 2773 38934 7623 38936
rect 2773 38931 2839 38934
rect 7281 38931 7347 38934
rect 7557 38931 7623 38934
rect 8293 38994 8359 38997
rect 9857 38994 9923 38997
rect 8293 38992 9923 38994
rect 8293 38936 8298 38992
rect 8354 38936 9862 38992
rect 9918 38936 9923 38992
rect 8293 38934 9923 38936
rect 8293 38931 8359 38934
rect 9857 38931 9923 38934
rect 1025 38858 1091 38861
rect 4981 38858 5047 38861
rect 1025 38856 5047 38858
rect 1025 38800 1030 38856
rect 1086 38800 4986 38856
rect 5042 38800 5047 38856
rect 1025 38798 5047 38800
rect 1025 38795 1091 38798
rect 4981 38795 5047 38798
rect 9765 38858 9831 38861
rect 10133 38858 10199 38861
rect 9765 38856 10199 38858
rect 9765 38800 9770 38856
rect 9826 38800 10138 38856
rect 10194 38800 10199 38856
rect 9765 38798 10199 38800
rect 9765 38795 9831 38798
rect 10133 38795 10199 38798
rect 5022 38660 5028 38724
rect 5092 38722 5098 38724
rect 5165 38722 5231 38725
rect 5092 38720 5231 38722
rect 5092 38664 5170 38720
rect 5226 38664 5231 38720
rect 5092 38662 5231 38664
rect 5092 38660 5098 38662
rect 5165 38659 5231 38662
rect 4318 38656 4634 38657
rect 4318 38592 4324 38656
rect 4388 38592 4404 38656
rect 4468 38592 4484 38656
rect 4548 38592 4564 38656
rect 4628 38592 4634 38656
rect 4318 38591 4634 38592
rect 10718 38656 11034 38657
rect 10718 38592 10724 38656
rect 10788 38592 10804 38656
rect 10868 38592 10884 38656
rect 10948 38592 10964 38656
rect 11028 38592 11034 38656
rect 10718 38591 11034 38592
rect 1853 38586 1919 38589
rect 2313 38586 2379 38589
rect 1853 38584 2379 38586
rect 1853 38528 1858 38584
rect 1914 38528 2318 38584
rect 2374 38528 2379 38584
rect 1853 38526 2379 38528
rect 1853 38523 1919 38526
rect 2313 38523 2379 38526
rect 5717 38586 5783 38589
rect 7833 38586 7899 38589
rect 8569 38586 8635 38589
rect 10317 38586 10383 38589
rect 5717 38584 7899 38586
rect 5717 38528 5722 38584
rect 5778 38528 7838 38584
rect 7894 38528 7899 38584
rect 5717 38526 7899 38528
rect 5717 38523 5783 38526
rect 7833 38523 7899 38526
rect 7974 38584 8635 38586
rect 7974 38528 8574 38584
rect 8630 38528 8635 38584
rect 7974 38526 8635 38528
rect 2865 38450 2931 38453
rect 3785 38450 3851 38453
rect 5574 38450 5580 38452
rect 2865 38448 5580 38450
rect 2865 38392 2870 38448
rect 2926 38392 3790 38448
rect 3846 38392 5580 38448
rect 2865 38390 5580 38392
rect 2865 38387 2931 38390
rect 3785 38387 3851 38390
rect 5574 38388 5580 38390
rect 5644 38388 5650 38452
rect 7465 38450 7531 38453
rect 7649 38450 7715 38453
rect 7465 38448 7715 38450
rect 7465 38392 7470 38448
rect 7526 38392 7654 38448
rect 7710 38392 7715 38448
rect 7465 38390 7715 38392
rect 7465 38387 7531 38390
rect 7649 38387 7715 38390
rect 7833 38450 7899 38453
rect 7974 38450 8034 38526
rect 8569 38523 8635 38526
rect 8710 38584 10383 38586
rect 8710 38528 10322 38584
rect 10378 38528 10383 38584
rect 8710 38526 10383 38528
rect 7833 38448 8034 38450
rect 7833 38392 7838 38448
rect 7894 38392 8034 38448
rect 7833 38390 8034 38392
rect 8385 38450 8451 38453
rect 8710 38450 8770 38526
rect 10317 38523 10383 38526
rect 9121 38452 9187 38453
rect 9070 38450 9076 38452
rect 8385 38448 8770 38450
rect 8385 38392 8390 38448
rect 8446 38392 8770 38448
rect 8385 38390 8770 38392
rect 9030 38390 9076 38450
rect 9140 38448 9187 38452
rect 9182 38392 9187 38448
rect 7833 38387 7899 38390
rect 8385 38387 8451 38390
rect 9070 38388 9076 38390
rect 9140 38388 9187 38392
rect 9121 38387 9187 38388
rect 3601 38314 3667 38317
rect 3374 38312 3667 38314
rect 3374 38256 3606 38312
rect 3662 38256 3667 38312
rect 3374 38254 3667 38256
rect 289 38042 355 38045
rect 2957 38042 3023 38045
rect 3374 38042 3434 38254
rect 3601 38251 3667 38254
rect 6913 38314 6979 38317
rect 7373 38314 7439 38317
rect 8109 38314 8175 38317
rect 8477 38316 8543 38317
rect 8753 38316 8819 38317
rect 8477 38314 8524 38316
rect 6913 38312 8175 38314
rect 6913 38256 6918 38312
rect 6974 38256 7378 38312
rect 7434 38256 8114 38312
rect 8170 38256 8175 38312
rect 6913 38254 8175 38256
rect 8432 38312 8524 38314
rect 8432 38256 8482 38312
rect 8432 38254 8524 38256
rect 6913 38251 6979 38254
rect 7373 38251 7439 38254
rect 8109 38251 8175 38254
rect 8477 38252 8524 38254
rect 8588 38252 8594 38316
rect 8702 38252 8708 38316
rect 8772 38314 8819 38316
rect 8772 38312 8864 38314
rect 8814 38256 8864 38312
rect 8772 38254 8864 38256
rect 8772 38252 8819 38254
rect 8477 38251 8543 38252
rect 8753 38251 8819 38252
rect 4429 38178 4495 38181
rect 7741 38178 7807 38181
rect 8150 38178 8156 38180
rect 4429 38176 8156 38178
rect 4429 38120 4434 38176
rect 4490 38120 7746 38176
rect 7802 38120 8156 38176
rect 4429 38118 8156 38120
rect 4429 38115 4495 38118
rect 7741 38115 7807 38118
rect 8150 38116 8156 38118
rect 8220 38178 8226 38180
rect 8477 38178 8543 38181
rect 8220 38176 8543 38178
rect 8220 38120 8482 38176
rect 8538 38120 8543 38176
rect 8220 38118 8543 38120
rect 8220 38116 8226 38118
rect 8477 38115 8543 38118
rect 9254 38116 9260 38180
rect 9324 38178 9330 38180
rect 9397 38178 9463 38181
rect 9324 38176 9463 38178
rect 9324 38120 9402 38176
rect 9458 38120 9463 38176
rect 9324 38118 9463 38120
rect 9324 38116 9330 38118
rect 9397 38115 9463 38118
rect 3658 38112 3974 38113
rect 3658 38048 3664 38112
rect 3728 38048 3744 38112
rect 3808 38048 3824 38112
rect 3888 38048 3904 38112
rect 3968 38048 3974 38112
rect 3658 38047 3974 38048
rect 10058 38112 10374 38113
rect 10058 38048 10064 38112
rect 10128 38048 10144 38112
rect 10208 38048 10224 38112
rect 10288 38048 10304 38112
rect 10368 38048 10374 38112
rect 10058 38047 10374 38048
rect 289 38040 3023 38042
rect 289 37984 294 38040
rect 350 37984 2962 38040
rect 3018 37984 3023 38040
rect 289 37982 3023 37984
rect 289 37979 355 37982
rect 2957 37979 3023 37982
rect 3190 37982 3434 38042
rect 3190 37773 3250 37982
rect 8886 37980 8892 38044
rect 8956 38042 8962 38044
rect 9857 38042 9923 38045
rect 8956 38040 9923 38042
rect 8956 37984 9862 38040
rect 9918 37984 9923 38040
rect 8956 37982 9923 37984
rect 8956 37980 8962 37982
rect 9857 37979 9923 37982
rect 3366 37844 3372 37908
rect 3436 37906 3442 37908
rect 3601 37906 3667 37909
rect 3436 37904 3667 37906
rect 3436 37848 3606 37904
rect 3662 37848 3667 37904
rect 3436 37846 3667 37848
rect 3436 37844 3442 37846
rect 3601 37843 3667 37846
rect 8385 37906 8451 37909
rect 9581 37906 9647 37909
rect 8385 37904 9647 37906
rect 8385 37848 8390 37904
rect 8446 37848 9586 37904
rect 9642 37848 9647 37904
rect 8385 37846 9647 37848
rect 8385 37843 8451 37846
rect 9581 37843 9647 37846
rect 3190 37768 3299 37773
rect 3190 37712 3238 37768
rect 3294 37712 3299 37768
rect 3190 37710 3299 37712
rect 3233 37707 3299 37710
rect 7741 37770 7807 37773
rect 9765 37770 9831 37773
rect 7741 37768 9831 37770
rect 7741 37712 7746 37768
rect 7802 37712 9770 37768
rect 9826 37712 9831 37768
rect 7741 37710 9831 37712
rect 7741 37707 7807 37710
rect 9765 37707 9831 37710
rect 6821 37634 6887 37637
rect 9397 37634 9463 37637
rect 6821 37632 9463 37634
rect 6821 37576 6826 37632
rect 6882 37576 9402 37632
rect 9458 37576 9463 37632
rect 6821 37574 9463 37576
rect 6821 37571 6887 37574
rect 9397 37571 9463 37574
rect 4318 37568 4634 37569
rect 4318 37504 4324 37568
rect 4388 37504 4404 37568
rect 4468 37504 4484 37568
rect 4548 37504 4564 37568
rect 4628 37504 4634 37568
rect 4318 37503 4634 37504
rect 10718 37568 11034 37569
rect 10718 37504 10724 37568
rect 10788 37504 10804 37568
rect 10868 37504 10884 37568
rect 10948 37504 10964 37568
rect 11028 37504 11034 37568
rect 10718 37503 11034 37504
rect 8477 37500 8543 37501
rect 8477 37498 8524 37500
rect 8432 37496 8524 37498
rect 8432 37440 8482 37496
rect 8432 37438 8524 37440
rect 8477 37436 8524 37438
rect 8588 37436 8594 37500
rect 8661 37498 8727 37501
rect 8886 37498 8892 37500
rect 8661 37496 8892 37498
rect 8661 37440 8666 37496
rect 8722 37440 8892 37496
rect 8661 37438 8892 37440
rect 8477 37435 8543 37436
rect 8661 37435 8727 37438
rect 8886 37436 8892 37438
rect 8956 37436 8962 37500
rect 9305 37498 9371 37501
rect 9438 37498 9444 37500
rect 9305 37496 9444 37498
rect 9305 37440 9310 37496
rect 9366 37440 9444 37496
rect 9305 37438 9444 37440
rect 9305 37435 9371 37438
rect 9438 37436 9444 37438
rect 9508 37436 9514 37500
rect 1342 37300 1348 37364
rect 1412 37362 1418 37364
rect 2313 37362 2379 37365
rect 1412 37360 2379 37362
rect 1412 37304 2318 37360
rect 2374 37304 2379 37360
rect 1412 37302 2379 37304
rect 1412 37300 1418 37302
rect 2313 37299 2379 37302
rect 6729 37362 6795 37365
rect 9765 37362 9831 37365
rect 6729 37360 9831 37362
rect 6729 37304 6734 37360
rect 6790 37304 9770 37360
rect 9826 37304 9831 37360
rect 6729 37302 9831 37304
rect 6729 37299 6795 37302
rect 9765 37299 9831 37302
rect 7465 37226 7531 37229
rect 8569 37226 8635 37229
rect 7465 37224 8635 37226
rect 7465 37168 7470 37224
rect 7526 37168 8574 37224
rect 8630 37168 8635 37224
rect 7465 37166 8635 37168
rect 7465 37163 7531 37166
rect 8569 37163 8635 37166
rect 8937 37226 9003 37229
rect 9254 37226 9260 37228
rect 8937 37224 9260 37226
rect 8937 37168 8942 37224
rect 8998 37168 9260 37224
rect 8937 37166 9260 37168
rect 8937 37163 9003 37166
rect 9254 37164 9260 37166
rect 9324 37226 9330 37228
rect 9397 37226 9463 37229
rect 9324 37224 9463 37226
rect 9324 37168 9402 37224
rect 9458 37168 9463 37224
rect 9324 37166 9463 37168
rect 9324 37164 9330 37166
rect 9397 37163 9463 37166
rect 0 37092 400 37120
rect 0 37028 382 37092
rect 446 37028 452 37092
rect 5574 37028 5580 37092
rect 5644 37090 5650 37092
rect 8518 37090 8524 37092
rect 5644 37030 8524 37090
rect 5644 37028 5650 37030
rect 8518 37028 8524 37030
rect 8588 37028 8594 37092
rect 0 37000 400 37028
rect 3658 37024 3974 37025
rect 3658 36960 3664 37024
rect 3728 36960 3744 37024
rect 3808 36960 3824 37024
rect 3888 36960 3904 37024
rect 3968 36960 3974 37024
rect 3658 36959 3974 36960
rect 10058 37024 10374 37025
rect 10058 36960 10064 37024
rect 10128 36960 10144 37024
rect 10208 36960 10224 37024
rect 10288 36960 10304 37024
rect 10368 36960 10374 37024
rect 10058 36959 10374 36960
rect 0 36818 400 36848
rect 749 36818 815 36821
rect 0 36816 815 36818
rect 0 36760 754 36816
rect 810 36760 815 36816
rect 0 36758 815 36760
rect 0 36728 400 36758
rect 749 36755 815 36758
rect 3785 36818 3851 36821
rect 5441 36820 5507 36821
rect 5390 36818 5396 36820
rect 3785 36816 5396 36818
rect 5460 36818 5507 36820
rect 5809 36818 5875 36821
rect 5460 36816 5875 36818
rect 3785 36760 3790 36816
rect 3846 36760 5396 36816
rect 5502 36760 5814 36816
rect 5870 36760 5875 36816
rect 3785 36758 5396 36760
rect 3785 36755 3851 36758
rect 5390 36756 5396 36758
rect 5460 36758 5875 36760
rect 5460 36756 5507 36758
rect 5441 36755 5507 36756
rect 5809 36755 5875 36758
rect 6126 36756 6132 36820
rect 6196 36818 6202 36820
rect 7925 36818 7991 36821
rect 8334 36818 8340 36820
rect 6196 36816 8340 36818
rect 6196 36760 7930 36816
rect 7986 36760 8340 36816
rect 6196 36758 8340 36760
rect 6196 36756 6202 36758
rect 7925 36755 7991 36758
rect 8334 36756 8340 36758
rect 8404 36756 8410 36820
rect 8385 36682 8451 36685
rect 9857 36682 9923 36685
rect 8385 36680 9923 36682
rect 8385 36624 8390 36680
rect 8446 36624 9862 36680
rect 9918 36624 9923 36680
rect 8385 36622 9923 36624
rect 8385 36619 8451 36622
rect 9857 36619 9923 36622
rect 0 36546 400 36576
rect 7189 36546 7255 36549
rect 9213 36546 9279 36549
rect 0 36486 2790 36546
rect 0 36456 400 36486
rect 0 36274 400 36304
rect 657 36274 723 36277
rect 0 36272 723 36274
rect 0 36216 662 36272
rect 718 36216 723 36272
rect 0 36214 723 36216
rect 2730 36274 2790 36486
rect 7189 36544 9279 36546
rect 7189 36488 7194 36544
rect 7250 36488 9218 36544
rect 9274 36488 9279 36544
rect 7189 36486 9279 36488
rect 7189 36483 7255 36486
rect 9213 36483 9279 36486
rect 4318 36480 4634 36481
rect 4318 36416 4324 36480
rect 4388 36416 4404 36480
rect 4468 36416 4484 36480
rect 4548 36416 4564 36480
rect 4628 36416 4634 36480
rect 4318 36415 4634 36416
rect 10718 36480 11034 36481
rect 10718 36416 10724 36480
rect 10788 36416 10804 36480
rect 10868 36416 10884 36480
rect 10948 36416 10964 36480
rect 11028 36416 11034 36480
rect 10718 36415 11034 36416
rect 2865 36410 2931 36413
rect 3182 36410 3188 36412
rect 2865 36408 3188 36410
rect 2865 36352 2870 36408
rect 2926 36352 3188 36408
rect 2865 36350 3188 36352
rect 2865 36347 2931 36350
rect 3182 36348 3188 36350
rect 3252 36348 3258 36412
rect 8937 36410 9003 36413
rect 9070 36410 9076 36412
rect 8937 36408 9076 36410
rect 8937 36352 8942 36408
rect 8998 36352 9076 36408
rect 8937 36350 9076 36352
rect 8937 36347 9003 36350
rect 9070 36348 9076 36350
rect 9140 36410 9146 36412
rect 9489 36410 9555 36413
rect 9140 36408 9555 36410
rect 9140 36352 9494 36408
rect 9550 36352 9555 36408
rect 9140 36350 9555 36352
rect 9140 36348 9146 36350
rect 9489 36347 9555 36350
rect 5809 36274 5875 36277
rect 2730 36272 5875 36274
rect 2730 36216 5814 36272
rect 5870 36216 5875 36272
rect 2730 36214 5875 36216
rect 0 36184 400 36214
rect 657 36211 723 36214
rect 5809 36211 5875 36214
rect 4838 36138 4844 36140
rect 2822 36078 4844 36138
rect 2822 36005 2882 36078
rect 4838 36076 4844 36078
rect 4908 36076 4914 36140
rect 8385 36138 8451 36141
rect 10593 36138 10659 36141
rect 8385 36136 10659 36138
rect 8385 36080 8390 36136
rect 8446 36080 10598 36136
rect 10654 36080 10659 36136
rect 8385 36078 10659 36080
rect 8385 36075 8451 36078
rect 10593 36075 10659 36078
rect 2773 36000 2882 36005
rect 2773 35944 2778 36000
rect 2834 35944 2882 36000
rect 2773 35942 2882 35944
rect 8477 36002 8543 36005
rect 9070 36002 9076 36004
rect 8477 36000 9076 36002
rect 8477 35944 8482 36000
rect 8538 35944 9076 36000
rect 8477 35942 9076 35944
rect 2773 35939 2839 35942
rect 8477 35939 8543 35942
rect 9070 35940 9076 35942
rect 9140 35940 9146 36004
rect 3658 35936 3974 35937
rect 3658 35872 3664 35936
rect 3728 35872 3744 35936
rect 3808 35872 3824 35936
rect 3888 35872 3904 35936
rect 3968 35872 3974 35936
rect 3658 35871 3974 35872
rect 10058 35936 10374 35937
rect 10058 35872 10064 35936
rect 10128 35872 10144 35936
rect 10208 35872 10224 35936
rect 10288 35872 10304 35936
rect 10368 35872 10374 35936
rect 10058 35871 10374 35872
rect 4061 35866 4127 35869
rect 7373 35866 7439 35869
rect 4061 35864 7439 35866
rect 4061 35808 4066 35864
rect 4122 35808 7378 35864
rect 7434 35808 7439 35864
rect 4061 35806 7439 35808
rect 4061 35803 4127 35806
rect 7373 35803 7439 35806
rect 6729 35730 6795 35733
rect 8150 35730 8156 35732
rect 6729 35728 8156 35730
rect 6729 35672 6734 35728
rect 6790 35672 8156 35728
rect 6729 35670 8156 35672
rect 6729 35667 6795 35670
rect 8150 35668 8156 35670
rect 8220 35730 8226 35732
rect 8569 35730 8635 35733
rect 8220 35728 8635 35730
rect 8220 35672 8574 35728
rect 8630 35672 8635 35728
rect 8220 35670 8635 35672
rect 8220 35668 8226 35670
rect 8569 35667 8635 35670
rect 5809 35594 5875 35597
rect 7046 35594 7052 35596
rect 5809 35592 7052 35594
rect 5809 35536 5814 35592
rect 5870 35536 7052 35592
rect 5809 35534 7052 35536
rect 5809 35531 5875 35534
rect 7046 35532 7052 35534
rect 7116 35532 7122 35596
rect 4318 35392 4634 35393
rect 4318 35328 4324 35392
rect 4388 35328 4404 35392
rect 4468 35328 4484 35392
rect 4548 35328 4564 35392
rect 4628 35328 4634 35392
rect 4318 35327 4634 35328
rect 10718 35392 11034 35393
rect 10718 35328 10724 35392
rect 10788 35328 10804 35392
rect 10868 35328 10884 35392
rect 10948 35328 10964 35392
rect 11028 35328 11034 35392
rect 10718 35327 11034 35328
rect 197 35186 263 35189
rect 422 35186 428 35188
rect 197 35184 428 35186
rect 197 35128 202 35184
rect 258 35128 428 35184
rect 197 35126 428 35128
rect 197 35123 263 35126
rect 422 35124 428 35126
rect 492 35186 498 35188
rect 1117 35186 1183 35189
rect 1853 35188 1919 35189
rect 1853 35186 1900 35188
rect 492 35184 1183 35186
rect 492 35128 1122 35184
rect 1178 35128 1183 35184
rect 492 35126 1183 35128
rect 1808 35184 1900 35186
rect 1808 35128 1858 35184
rect 1808 35126 1900 35128
rect 492 35124 498 35126
rect 1117 35123 1183 35126
rect 1853 35124 1900 35126
rect 1964 35124 1970 35188
rect 3969 35186 4035 35189
rect 8293 35186 8359 35189
rect 9254 35186 9260 35188
rect 3969 35184 9260 35186
rect 3969 35128 3974 35184
rect 4030 35128 8298 35184
rect 8354 35128 9260 35184
rect 3969 35126 9260 35128
rect 1853 35123 1919 35124
rect 3969 35123 4035 35126
rect 8293 35123 8359 35126
rect 9254 35124 9260 35126
rect 9324 35186 9330 35188
rect 9949 35186 10015 35189
rect 9324 35184 10015 35186
rect 9324 35128 9954 35184
rect 10010 35128 10015 35184
rect 9324 35126 10015 35128
rect 9324 35124 9330 35126
rect 9949 35123 10015 35126
rect 974 34988 980 35052
rect 1044 35050 1050 35052
rect 2957 35050 3023 35053
rect 1044 35048 3023 35050
rect 1044 34992 2962 35048
rect 3018 34992 3023 35048
rect 1044 34990 3023 34992
rect 1044 34988 1050 34990
rect 2957 34987 3023 34990
rect 4613 35050 4679 35053
rect 5390 35050 5396 35052
rect 4613 35048 5396 35050
rect 4613 34992 4618 35048
rect 4674 34992 5396 35048
rect 4613 34990 5396 34992
rect 4613 34987 4679 34990
rect 5390 34988 5396 34990
rect 5460 34988 5466 35052
rect 8845 35050 8911 35053
rect 10593 35050 10659 35053
rect 8845 35048 10659 35050
rect 8845 34992 8850 35048
rect 8906 34992 10598 35048
rect 10654 34992 10659 35048
rect 8845 34990 10659 34992
rect 8845 34987 8911 34990
rect 10593 34987 10659 34990
rect 0 34914 400 34944
rect 1117 34914 1183 34917
rect 0 34912 1183 34914
rect 0 34856 1122 34912
rect 1178 34856 1183 34912
rect 0 34854 1183 34856
rect 0 34824 400 34854
rect 1117 34851 1183 34854
rect 2446 34852 2452 34916
rect 2516 34914 2522 34916
rect 2681 34914 2747 34917
rect 2516 34912 2747 34914
rect 2516 34856 2686 34912
rect 2742 34856 2747 34912
rect 2516 34854 2747 34856
rect 2516 34852 2522 34854
rect 2681 34851 2747 34854
rect 5073 34914 5139 34917
rect 7782 34914 7788 34916
rect 5073 34912 7788 34914
rect 5073 34856 5078 34912
rect 5134 34856 7788 34912
rect 5073 34854 7788 34856
rect 5073 34851 5139 34854
rect 7782 34852 7788 34854
rect 7852 34852 7858 34916
rect 3658 34848 3974 34849
rect 3658 34784 3664 34848
rect 3728 34784 3744 34848
rect 3808 34784 3824 34848
rect 3888 34784 3904 34848
rect 3968 34784 3974 34848
rect 3658 34783 3974 34784
rect 10058 34848 10374 34849
rect 10058 34784 10064 34848
rect 10128 34784 10144 34848
rect 10208 34784 10224 34848
rect 10288 34784 10304 34848
rect 10368 34784 10374 34848
rect 10058 34783 10374 34784
rect 1945 34780 2011 34781
rect 1894 34778 1900 34780
rect 1854 34718 1900 34778
rect 1964 34776 2011 34780
rect 2006 34720 2011 34776
rect 1894 34716 1900 34718
rect 1964 34716 2011 34720
rect 1945 34715 2011 34716
rect 4061 34778 4127 34781
rect 5165 34778 5231 34781
rect 5901 34778 5967 34781
rect 4061 34776 5967 34778
rect 4061 34720 4066 34776
rect 4122 34720 5170 34776
rect 5226 34720 5906 34776
rect 5962 34720 5967 34776
rect 4061 34718 5967 34720
rect 4061 34715 4127 34718
rect 5165 34715 5231 34718
rect 5901 34715 5967 34718
rect 0 34642 400 34672
rect 2681 34642 2747 34645
rect 0 34640 2747 34642
rect 0 34584 2686 34640
rect 2742 34584 2747 34640
rect 0 34582 2747 34584
rect 0 34552 400 34582
rect 2681 34579 2747 34582
rect 3969 34642 4035 34645
rect 4102 34642 4108 34644
rect 3969 34640 4108 34642
rect 3969 34584 3974 34640
rect 4030 34584 4108 34640
rect 3969 34582 4108 34584
rect 3969 34579 4035 34582
rect 4102 34580 4108 34582
rect 4172 34580 4178 34644
rect 6637 34642 6703 34645
rect 8569 34642 8635 34645
rect 9213 34642 9279 34645
rect 6637 34640 9279 34642
rect 6637 34584 6642 34640
rect 6698 34584 8574 34640
rect 8630 34584 9218 34640
rect 9274 34584 9279 34640
rect 6637 34582 9279 34584
rect 6637 34579 6703 34582
rect 8569 34579 8635 34582
rect 9213 34579 9279 34582
rect 3785 34506 3851 34509
rect 5165 34508 5231 34509
rect 4838 34506 4844 34508
rect 3785 34504 4844 34506
rect 3785 34448 3790 34504
rect 3846 34448 4844 34504
rect 3785 34446 4844 34448
rect 3785 34443 3851 34446
rect 4838 34444 4844 34446
rect 4908 34444 4914 34508
rect 5165 34504 5212 34508
rect 5276 34506 5282 34508
rect 7833 34506 7899 34509
rect 8150 34506 8156 34508
rect 5165 34448 5170 34504
rect 5165 34444 5212 34448
rect 5276 34446 5322 34506
rect 7833 34504 8156 34506
rect 7833 34448 7838 34504
rect 7894 34448 8156 34504
rect 7833 34446 8156 34448
rect 5276 34444 5282 34446
rect 5165 34443 5231 34444
rect 7833 34443 7899 34446
rect 8150 34444 8156 34446
rect 8220 34444 8226 34508
rect 8477 34506 8543 34509
rect 9213 34506 9279 34509
rect 10961 34506 11027 34509
rect 8477 34504 11027 34506
rect 8477 34448 8482 34504
rect 8538 34448 9218 34504
rect 9274 34448 10966 34504
rect 11022 34448 11027 34504
rect 8477 34446 11027 34448
rect 8477 34443 8543 34446
rect 9213 34443 9279 34446
rect 10961 34443 11027 34446
rect 0 34370 400 34400
rect 933 34370 999 34373
rect 0 34368 999 34370
rect 0 34312 938 34368
rect 994 34312 999 34368
rect 0 34310 999 34312
rect 0 34280 400 34310
rect 933 34307 999 34310
rect 5349 34370 5415 34373
rect 8702 34370 8708 34372
rect 5349 34368 8708 34370
rect 5349 34312 5354 34368
rect 5410 34312 8708 34368
rect 5349 34310 8708 34312
rect 5349 34307 5415 34310
rect 8702 34308 8708 34310
rect 8772 34308 8778 34372
rect 4318 34304 4634 34305
rect 4318 34240 4324 34304
rect 4388 34240 4404 34304
rect 4468 34240 4484 34304
rect 4548 34240 4564 34304
rect 4628 34240 4634 34304
rect 4318 34239 4634 34240
rect 10718 34304 11034 34305
rect 10718 34240 10724 34304
rect 10788 34240 10804 34304
rect 10868 34240 10884 34304
rect 10948 34240 10964 34304
rect 11028 34240 11034 34304
rect 10718 34239 11034 34240
rect 3366 34036 3372 34100
rect 3436 34098 3442 34100
rect 5390 34098 5396 34100
rect 3436 34038 5396 34098
rect 3436 34036 3442 34038
rect 5390 34036 5396 34038
rect 5460 34036 5466 34100
rect 7833 34098 7899 34101
rect 7966 34098 7972 34100
rect 7833 34096 7972 34098
rect 7833 34040 7838 34096
rect 7894 34040 7972 34096
rect 7833 34038 7972 34040
rect 7833 34035 7899 34038
rect 7966 34036 7972 34038
rect 8036 34036 8042 34100
rect 8569 34098 8635 34101
rect 8845 34098 8911 34101
rect 8569 34096 8911 34098
rect 8569 34040 8574 34096
rect 8630 34040 8850 34096
rect 8906 34040 8911 34096
rect 8569 34038 8911 34040
rect 8569 34035 8635 34038
rect 8845 34035 8911 34038
rect 6361 33962 6427 33965
rect 7189 33962 7255 33965
rect 6361 33960 7255 33962
rect 6361 33904 6366 33960
rect 6422 33904 7194 33960
rect 7250 33904 7255 33960
rect 6361 33902 7255 33904
rect 6361 33899 6427 33902
rect 7189 33899 7255 33902
rect 8201 33960 8267 33965
rect 8201 33904 8206 33960
rect 8262 33904 8267 33960
rect 8201 33899 8267 33904
rect 8753 33962 8819 33965
rect 10542 33962 10548 33964
rect 8753 33960 10548 33962
rect 8753 33904 8758 33960
rect 8814 33904 10548 33960
rect 8753 33902 10548 33904
rect 8753 33899 8819 33902
rect 10542 33900 10548 33902
rect 10612 33900 10618 33964
rect 8204 33826 8264 33899
rect 8204 33766 8632 33826
rect 3658 33760 3974 33761
rect 3658 33696 3664 33760
rect 3728 33696 3744 33760
rect 3808 33696 3824 33760
rect 3888 33696 3904 33760
rect 3968 33696 3974 33760
rect 3658 33695 3974 33696
rect 7373 33690 7439 33693
rect 7373 33688 8264 33690
rect 7373 33632 7378 33688
rect 7434 33632 8264 33688
rect 7373 33630 8264 33632
rect 7373 33627 7439 33630
rect 8204 33557 8264 33630
rect 8572 33557 8632 33766
rect 10058 33760 10374 33761
rect 10058 33696 10064 33760
rect 10128 33696 10144 33760
rect 10208 33696 10224 33760
rect 10288 33696 10304 33760
rect 10368 33696 10374 33760
rect 10058 33695 10374 33696
rect 9438 33628 9444 33692
rect 9508 33690 9514 33692
rect 9857 33690 9923 33693
rect 9508 33688 9923 33690
rect 9508 33632 9862 33688
rect 9918 33632 9923 33688
rect 9508 33630 9923 33632
rect 9508 33628 9514 33630
rect 9857 33627 9923 33630
rect 5533 33554 5599 33557
rect 7598 33554 7604 33556
rect 5533 33552 7604 33554
rect 5533 33496 5538 33552
rect 5594 33496 7604 33552
rect 5533 33494 7604 33496
rect 5533 33491 5599 33494
rect 7598 33492 7604 33494
rect 7668 33492 7674 33556
rect 8201 33552 8267 33557
rect 8201 33496 8206 33552
rect 8262 33496 8267 33552
rect 8201 33491 8267 33496
rect 8569 33552 8635 33557
rect 8569 33496 8574 33552
rect 8630 33496 8635 33552
rect 8569 33491 8635 33496
rect 8150 33356 8156 33420
rect 8220 33418 8226 33420
rect 10409 33418 10475 33421
rect 8220 33416 10475 33418
rect 8220 33360 10414 33416
rect 10470 33360 10475 33416
rect 8220 33358 10475 33360
rect 8220 33356 8226 33358
rect 10409 33355 10475 33358
rect 1526 33220 1532 33284
rect 1596 33282 1602 33284
rect 2773 33282 2839 33285
rect 1596 33280 2839 33282
rect 1596 33224 2778 33280
rect 2834 33224 2839 33280
rect 1596 33222 2839 33224
rect 1596 33220 1602 33222
rect 2773 33219 2839 33222
rect 3366 33220 3372 33284
rect 3436 33282 3442 33284
rect 3969 33282 4035 33285
rect 3436 33280 4035 33282
rect 3436 33224 3974 33280
rect 4030 33224 4035 33280
rect 3436 33222 4035 33224
rect 3436 33220 3442 33222
rect 3969 33219 4035 33222
rect 7373 33282 7439 33285
rect 7925 33282 7991 33285
rect 8385 33282 8451 33285
rect 7373 33280 7850 33282
rect 7373 33224 7378 33280
rect 7434 33224 7850 33280
rect 7373 33222 7850 33224
rect 7373 33219 7439 33222
rect 4318 33216 4634 33217
rect 4318 33152 4324 33216
rect 4388 33152 4404 33216
rect 4468 33152 4484 33216
rect 4548 33152 4564 33216
rect 4628 33152 4634 33216
rect 4318 33151 4634 33152
rect 2037 33146 2103 33149
rect 2262 33146 2268 33148
rect 2037 33144 2268 33146
rect 2037 33088 2042 33144
rect 2098 33088 2268 33144
rect 2037 33086 2268 33088
rect 2037 33083 2103 33086
rect 2262 33084 2268 33086
rect 2332 33084 2338 33148
rect 6729 33146 6795 33149
rect 7465 33148 7531 33149
rect 6862 33146 6868 33148
rect 6729 33144 6868 33146
rect 6729 33088 6734 33144
rect 6790 33088 6868 33144
rect 6729 33086 6868 33088
rect 6729 33083 6795 33086
rect 6862 33084 6868 33086
rect 6932 33084 6938 33148
rect 7414 33084 7420 33148
rect 7484 33146 7531 33148
rect 7790 33146 7850 33222
rect 7925 33280 8451 33282
rect 7925 33224 7930 33280
rect 7986 33224 8390 33280
rect 8446 33224 8451 33280
rect 7925 33222 8451 33224
rect 7925 33219 7991 33222
rect 8385 33219 8451 33222
rect 8753 33282 8819 33285
rect 9213 33282 9279 33285
rect 8753 33280 9279 33282
rect 8753 33224 8758 33280
rect 8814 33224 9218 33280
rect 9274 33224 9279 33280
rect 8753 33222 9279 33224
rect 8753 33219 8819 33222
rect 9213 33219 9279 33222
rect 10718 33216 11034 33217
rect 10718 33152 10724 33216
rect 10788 33152 10804 33216
rect 10868 33152 10884 33216
rect 10948 33152 10964 33216
rect 11028 33152 11034 33216
rect 10718 33151 11034 33152
rect 8753 33146 8819 33149
rect 7484 33144 7576 33146
rect 7526 33088 7576 33144
rect 7484 33086 7576 33088
rect 7790 33144 8819 33146
rect 7790 33088 8758 33144
rect 8814 33088 8819 33144
rect 7790 33086 8819 33088
rect 7484 33084 7531 33086
rect 7465 33083 7531 33084
rect 8753 33083 8819 33086
rect 974 32948 980 33012
rect 1044 33010 1050 33012
rect 2497 33010 2563 33013
rect 1044 33008 2563 33010
rect 1044 32952 2502 33008
rect 2558 32952 2563 33008
rect 1044 32950 2563 32952
rect 1044 32948 1050 32950
rect 2497 32947 2563 32950
rect 3693 33010 3759 33013
rect 4429 33010 4495 33013
rect 9397 33010 9463 33013
rect 3693 33008 9463 33010
rect 3693 32952 3698 33008
rect 3754 32952 4434 33008
rect 4490 32952 9402 33008
rect 9458 32952 9463 33008
rect 3693 32950 9463 32952
rect 3693 32947 3759 32950
rect 4429 32947 4495 32950
rect 9397 32947 9463 32950
rect 2037 32874 2103 32877
rect 4889 32874 4955 32877
rect 2037 32872 4955 32874
rect 2037 32816 2042 32872
rect 2098 32816 4894 32872
rect 4950 32816 4955 32872
rect 2037 32814 4955 32816
rect 2037 32811 2103 32814
rect 4889 32811 4955 32814
rect 5533 32874 5599 32877
rect 8385 32874 8451 32877
rect 5533 32872 8451 32874
rect 5533 32816 5538 32872
rect 5594 32816 8390 32872
rect 8446 32816 8451 32872
rect 5533 32814 8451 32816
rect 5533 32811 5599 32814
rect 8385 32811 8451 32814
rect 5758 32676 5764 32740
rect 5828 32738 5834 32740
rect 5901 32738 5967 32741
rect 5828 32736 5967 32738
rect 5828 32680 5906 32736
rect 5962 32680 5967 32736
rect 5828 32678 5967 32680
rect 5828 32676 5834 32678
rect 5901 32675 5967 32678
rect 6269 32738 6335 32741
rect 8017 32738 8083 32741
rect 6269 32736 8083 32738
rect 6269 32680 6274 32736
rect 6330 32680 8022 32736
rect 8078 32680 8083 32736
rect 6269 32678 8083 32680
rect 6269 32675 6335 32678
rect 8017 32675 8083 32678
rect 8477 32738 8543 32741
rect 9070 32738 9076 32740
rect 8477 32736 9076 32738
rect 8477 32680 8482 32736
rect 8538 32680 9076 32736
rect 8477 32678 9076 32680
rect 8477 32675 8543 32678
rect 9070 32676 9076 32678
rect 9140 32676 9146 32740
rect 3658 32672 3974 32673
rect 3658 32608 3664 32672
rect 3728 32608 3744 32672
rect 3808 32608 3824 32672
rect 3888 32608 3904 32672
rect 3968 32608 3974 32672
rect 3658 32607 3974 32608
rect 10058 32672 10374 32673
rect 10058 32608 10064 32672
rect 10128 32608 10144 32672
rect 10208 32608 10224 32672
rect 10288 32608 10304 32672
rect 10368 32608 10374 32672
rect 10058 32607 10374 32608
rect 6177 32604 6243 32605
rect 6126 32540 6132 32604
rect 6196 32602 6243 32604
rect 7925 32604 7991 32605
rect 6196 32600 6288 32602
rect 6238 32544 6288 32600
rect 6196 32542 6288 32544
rect 7925 32600 7972 32604
rect 8036 32602 8042 32604
rect 8937 32602 9003 32605
rect 9070 32602 9076 32604
rect 7925 32544 7930 32600
rect 6196 32540 6243 32542
rect 6177 32539 6243 32540
rect 7925 32540 7972 32544
rect 8036 32542 8082 32602
rect 8937 32600 9076 32602
rect 8937 32544 8942 32600
rect 8998 32544 9076 32600
rect 8937 32542 9076 32544
rect 8036 32540 8042 32542
rect 7925 32539 7991 32540
rect 8937 32539 9003 32542
rect 9070 32540 9076 32542
rect 9140 32540 9146 32604
rect 5441 32466 5507 32469
rect 5574 32466 5580 32468
rect 5441 32464 5580 32466
rect 5441 32408 5446 32464
rect 5502 32408 5580 32464
rect 5441 32406 5580 32408
rect 5441 32403 5507 32406
rect 5574 32404 5580 32406
rect 5644 32404 5650 32468
rect 9305 32466 9371 32469
rect 5766 32464 9506 32466
rect 5766 32408 9310 32464
rect 9366 32408 9506 32464
rect 5766 32406 9506 32408
rect 2405 32330 2471 32333
rect 5766 32330 5826 32406
rect 9305 32403 9371 32406
rect 9446 32333 9506 32406
rect 2405 32328 2790 32330
rect 2405 32272 2410 32328
rect 2466 32272 2790 32328
rect 2405 32270 2790 32272
rect 2405 32267 2471 32270
rect 2730 32194 2790 32270
rect 4110 32270 5826 32330
rect 5901 32330 5967 32333
rect 9029 32330 9095 32333
rect 5901 32328 9095 32330
rect 5901 32272 5906 32328
rect 5962 32272 9034 32328
rect 9090 32272 9095 32328
rect 5901 32270 9095 32272
rect 9446 32328 9555 32333
rect 9446 32272 9494 32328
rect 9550 32272 9555 32328
rect 9446 32270 9555 32272
rect 4110 32194 4170 32270
rect 5901 32267 5967 32270
rect 9029 32267 9095 32270
rect 9489 32267 9555 32270
rect 2730 32134 4170 32194
rect 2313 31924 2379 31925
rect 2262 31860 2268 31924
rect 2332 31922 2379 31924
rect 3141 31922 3207 31925
rect 3325 31922 3391 31925
rect 2332 31920 2424 31922
rect 2374 31864 2424 31920
rect 2332 31862 2424 31864
rect 3141 31920 3391 31922
rect 3141 31864 3146 31920
rect 3202 31864 3330 31920
rect 3386 31864 3391 31920
rect 3141 31862 3391 31864
rect 2332 31860 2379 31862
rect 2313 31859 2379 31860
rect 3141 31859 3207 31862
rect 3325 31859 3391 31862
rect 289 31786 355 31789
rect 2773 31786 2839 31789
rect 289 31784 2839 31786
rect 289 31728 294 31784
rect 350 31728 2778 31784
rect 2834 31728 2839 31784
rect 289 31726 2839 31728
rect 289 31723 355 31726
rect 2773 31723 2839 31726
rect 3325 31786 3391 31789
rect 3601 31786 3667 31789
rect 3325 31784 3667 31786
rect 3325 31728 3330 31784
rect 3386 31728 3606 31784
rect 3662 31728 3667 31784
rect 3325 31726 3667 31728
rect 4110 31786 4170 32134
rect 6913 32194 6979 32197
rect 6913 32192 7620 32194
rect 6913 32136 6918 32192
rect 6974 32136 7620 32192
rect 6913 32134 7620 32136
rect 6913 32131 6979 32134
rect 4318 32128 4634 32129
rect 4318 32064 4324 32128
rect 4388 32064 4404 32128
rect 4468 32064 4484 32128
rect 4548 32064 4564 32128
rect 4628 32064 4634 32128
rect 4318 32063 4634 32064
rect 5901 32058 5967 32061
rect 6085 32058 6151 32061
rect 5901 32056 6151 32058
rect 5901 32000 5906 32056
rect 5962 32000 6090 32056
rect 6146 32000 6151 32056
rect 5901 31998 6151 32000
rect 5901 31995 5967 31998
rect 6085 31995 6151 31998
rect 6862 31996 6868 32060
rect 6932 32058 6938 32060
rect 7097 32058 7163 32061
rect 6932 32056 7163 32058
rect 6932 32000 7102 32056
rect 7158 32000 7163 32056
rect 6932 31998 7163 32000
rect 6932 31996 6938 31998
rect 7097 31995 7163 31998
rect 7560 31925 7620 32134
rect 10718 32128 11034 32129
rect 10718 32064 10724 32128
rect 10788 32064 10804 32128
rect 10868 32064 10884 32128
rect 10948 32064 10964 32128
rect 11028 32064 11034 32128
rect 10718 32063 11034 32064
rect 7741 32060 7807 32061
rect 7741 32056 7788 32060
rect 7852 32058 7858 32060
rect 7741 32000 7746 32056
rect 7741 31996 7788 32000
rect 7852 31998 7898 32058
rect 7852 31996 7858 31998
rect 7966 31996 7972 32060
rect 8036 32058 8042 32060
rect 8293 32058 8359 32061
rect 8036 32056 8359 32058
rect 8036 32000 8298 32056
rect 8354 32000 8359 32056
rect 8036 31998 8359 32000
rect 8036 31996 8042 31998
rect 7741 31995 7807 31996
rect 8293 31995 8359 31998
rect 8937 32058 9003 32061
rect 9070 32058 9076 32060
rect 8937 32056 9076 32058
rect 8937 32000 8942 32056
rect 8998 32000 9076 32056
rect 8937 31998 9076 32000
rect 8937 31995 9003 31998
rect 9070 31996 9076 31998
rect 9140 31996 9146 32060
rect 4429 31922 4495 31925
rect 5165 31922 5231 31925
rect 4429 31920 5231 31922
rect 4429 31864 4434 31920
rect 4490 31864 5170 31920
rect 5226 31864 5231 31920
rect 4429 31862 5231 31864
rect 4429 31859 4495 31862
rect 5165 31859 5231 31862
rect 6085 31922 6151 31925
rect 7005 31922 7071 31925
rect 6085 31920 7071 31922
rect 6085 31864 6090 31920
rect 6146 31864 7010 31920
rect 7066 31864 7071 31920
rect 6085 31862 7071 31864
rect 6085 31859 6151 31862
rect 7005 31859 7071 31862
rect 7557 31920 7623 31925
rect 7557 31864 7562 31920
rect 7618 31864 7623 31920
rect 7557 31859 7623 31864
rect 4705 31786 4771 31789
rect 4110 31784 4771 31786
rect 4110 31728 4710 31784
rect 4766 31728 4771 31784
rect 4110 31726 4771 31728
rect 3325 31723 3391 31726
rect 3601 31723 3667 31726
rect 4705 31723 4771 31726
rect 4889 31786 4955 31789
rect 5206 31786 5212 31788
rect 4889 31784 5212 31786
rect 4889 31728 4894 31784
rect 4950 31728 5212 31784
rect 4889 31726 5212 31728
rect 4889 31723 4955 31726
rect 5206 31724 5212 31726
rect 5276 31724 5282 31788
rect 6729 31786 6795 31789
rect 7005 31786 7071 31789
rect 7414 31786 7420 31788
rect 6729 31784 6930 31786
rect 6729 31728 6734 31784
rect 6790 31728 6930 31784
rect 6729 31726 6930 31728
rect 6729 31723 6795 31726
rect 1761 31652 1827 31653
rect 1710 31588 1716 31652
rect 1780 31650 1827 31652
rect 1780 31648 1872 31650
rect 1822 31592 1872 31648
rect 1780 31590 1872 31592
rect 1780 31588 1827 31590
rect 5758 31588 5764 31652
rect 5828 31650 5834 31652
rect 6729 31650 6795 31653
rect 5828 31648 6795 31650
rect 5828 31592 6734 31648
rect 6790 31592 6795 31648
rect 5828 31590 6795 31592
rect 6870 31650 6930 31726
rect 7005 31784 7420 31786
rect 7005 31728 7010 31784
rect 7066 31728 7420 31784
rect 7005 31726 7420 31728
rect 7005 31723 7071 31726
rect 7414 31724 7420 31726
rect 7484 31724 7490 31788
rect 8753 31786 8819 31789
rect 10041 31786 10107 31789
rect 8753 31784 10107 31786
rect 8753 31728 8758 31784
rect 8814 31728 10046 31784
rect 10102 31728 10107 31784
rect 8753 31726 10107 31728
rect 8753 31723 8819 31726
rect 10041 31723 10107 31726
rect 8109 31650 8175 31653
rect 9121 31652 9187 31653
rect 6870 31648 8175 31650
rect 6870 31592 8114 31648
rect 8170 31592 8175 31648
rect 6870 31590 8175 31592
rect 5828 31588 5834 31590
rect 1761 31587 1827 31588
rect 6729 31587 6795 31590
rect 8109 31587 8175 31590
rect 9070 31588 9076 31652
rect 9140 31650 9187 31652
rect 9140 31648 9232 31650
rect 9182 31592 9232 31648
rect 9140 31590 9232 31592
rect 9140 31588 9187 31590
rect 9121 31587 9187 31588
rect 3658 31584 3974 31585
rect 3658 31520 3664 31584
rect 3728 31520 3744 31584
rect 3808 31520 3824 31584
rect 3888 31520 3904 31584
rect 3968 31520 3974 31584
rect 3658 31519 3974 31520
rect 10058 31584 10374 31585
rect 10058 31520 10064 31584
rect 10128 31520 10144 31584
rect 10208 31520 10224 31584
rect 10288 31520 10304 31584
rect 10368 31520 10374 31584
rect 10058 31519 10374 31520
rect 473 31514 539 31517
rect 1117 31514 1183 31517
rect 473 31512 1183 31514
rect 473 31456 478 31512
rect 534 31456 1122 31512
rect 1178 31456 1183 31512
rect 473 31454 1183 31456
rect 473 31451 539 31454
rect 1117 31451 1183 31454
rect 5257 31514 5323 31517
rect 5901 31514 5967 31517
rect 5257 31512 5967 31514
rect 5257 31456 5262 31512
rect 5318 31456 5906 31512
rect 5962 31456 5967 31512
rect 5257 31454 5967 31456
rect 5257 31451 5323 31454
rect 5901 31451 5967 31454
rect 7465 31514 7531 31517
rect 7782 31514 7788 31516
rect 7465 31512 7788 31514
rect 7465 31456 7470 31512
rect 7526 31456 7788 31512
rect 7465 31454 7788 31456
rect 7465 31451 7531 31454
rect 7782 31452 7788 31454
rect 7852 31452 7858 31516
rect 1117 31378 1183 31381
rect 1526 31378 1532 31380
rect 1117 31376 1532 31378
rect 1117 31320 1122 31376
rect 1178 31320 1532 31376
rect 1117 31318 1532 31320
rect 1117 31315 1183 31318
rect 1526 31316 1532 31318
rect 1596 31316 1602 31380
rect 6177 31376 6243 31381
rect 6177 31320 6182 31376
rect 6238 31320 6243 31376
rect 6177 31315 6243 31320
rect 1761 31108 1827 31109
rect 1710 31044 1716 31108
rect 1780 31106 1827 31108
rect 3509 31106 3575 31109
rect 1780 31104 1872 31106
rect 1822 31048 1872 31104
rect 1780 31046 1872 31048
rect 3509 31104 3618 31106
rect 3509 31048 3514 31104
rect 3570 31048 3618 31104
rect 1780 31044 1827 31046
rect 1761 31043 1827 31044
rect 3509 31043 3618 31048
rect 2313 30970 2379 30973
rect 3417 30970 3483 30973
rect 2313 30968 3483 30970
rect 2313 30912 2318 30968
rect 2374 30912 3422 30968
rect 3478 30912 3483 30968
rect 2313 30910 3483 30912
rect 2313 30907 2379 30910
rect 3417 30907 3483 30910
rect 3558 30837 3618 31043
rect 4318 31040 4634 31041
rect 4318 30976 4324 31040
rect 4388 30976 4404 31040
rect 4468 30976 4484 31040
rect 4548 30976 4564 31040
rect 4628 30976 4634 31040
rect 4318 30975 4634 30976
rect 4981 30970 5047 30973
rect 5574 30970 5580 30972
rect 4981 30968 5580 30970
rect 4981 30912 4986 30968
rect 5042 30912 5580 30968
rect 4981 30910 5580 30912
rect 4981 30907 5047 30910
rect 5574 30908 5580 30910
rect 5644 30908 5650 30972
rect 5809 30970 5875 30973
rect 6180 30970 6240 31315
rect 10718 31040 11034 31041
rect 10718 30976 10724 31040
rect 10788 30976 10804 31040
rect 10868 30976 10884 31040
rect 10948 30976 10964 31040
rect 11028 30976 11034 31040
rect 10718 30975 11034 30976
rect 5809 30968 6240 30970
rect 5809 30912 5814 30968
rect 5870 30912 6240 30968
rect 5809 30910 6240 30912
rect 5809 30907 5875 30910
rect 3509 30834 3618 30837
rect 5574 30834 5580 30836
rect 3509 30832 5580 30834
rect 3509 30776 3514 30832
rect 3570 30776 5580 30832
rect 3509 30774 5580 30776
rect 3509 30771 3575 30774
rect 5574 30772 5580 30774
rect 5644 30772 5650 30836
rect 6494 30772 6500 30836
rect 6564 30834 6570 30836
rect 7414 30834 7420 30836
rect 6564 30774 7420 30834
rect 6564 30772 6570 30774
rect 7414 30772 7420 30774
rect 7484 30834 7490 30836
rect 7557 30834 7623 30837
rect 7484 30832 7623 30834
rect 7484 30776 7562 30832
rect 7618 30776 7623 30832
rect 7484 30774 7623 30776
rect 7484 30772 7490 30774
rect 7557 30771 7623 30774
rect 3325 30698 3391 30701
rect 5901 30698 5967 30701
rect 3325 30696 5967 30698
rect 3325 30640 3330 30696
rect 3386 30640 5906 30696
rect 5962 30640 5967 30696
rect 3325 30638 5967 30640
rect 3325 30635 3391 30638
rect 5901 30635 5967 30638
rect 9622 30636 9628 30700
rect 9692 30698 9698 30700
rect 9949 30698 10015 30701
rect 9692 30696 10015 30698
rect 9692 30640 9954 30696
rect 10010 30640 10015 30696
rect 9692 30638 10015 30640
rect 9692 30636 9698 30638
rect 9949 30635 10015 30638
rect 2037 30562 2103 30565
rect 2957 30562 3023 30565
rect 2037 30560 3023 30562
rect 2037 30504 2042 30560
rect 2098 30504 2962 30560
rect 3018 30504 3023 30560
rect 2037 30502 3023 30504
rect 2037 30499 2103 30502
rect 2957 30499 3023 30502
rect 5758 30500 5764 30564
rect 5828 30562 5834 30564
rect 5901 30562 5967 30565
rect 6545 30564 6611 30565
rect 6494 30562 6500 30564
rect 5828 30560 5967 30562
rect 5828 30504 5906 30560
rect 5962 30504 5967 30560
rect 5828 30502 5967 30504
rect 6454 30502 6500 30562
rect 6564 30560 6611 30564
rect 6606 30504 6611 30560
rect 5828 30500 5834 30502
rect 5901 30499 5967 30502
rect 6494 30500 6500 30502
rect 6564 30500 6611 30504
rect 6545 30499 6611 30500
rect 8845 30562 8911 30565
rect 9806 30562 9812 30564
rect 8845 30560 9812 30562
rect 8845 30504 8850 30560
rect 8906 30504 9812 30560
rect 8845 30502 9812 30504
rect 8845 30499 8911 30502
rect 9806 30500 9812 30502
rect 9876 30500 9882 30564
rect 3658 30496 3974 30497
rect 3658 30432 3664 30496
rect 3728 30432 3744 30496
rect 3808 30432 3824 30496
rect 3888 30432 3904 30496
rect 3968 30432 3974 30496
rect 3658 30431 3974 30432
rect 10058 30496 10374 30497
rect 10058 30432 10064 30496
rect 10128 30432 10144 30496
rect 10208 30432 10224 30496
rect 10288 30432 10304 30496
rect 10368 30432 10374 30496
rect 10058 30431 10374 30432
rect 606 30364 612 30428
rect 676 30426 682 30428
rect 1342 30426 1348 30428
rect 676 30366 1348 30426
rect 676 30364 682 30366
rect 1342 30364 1348 30366
rect 1412 30364 1418 30428
rect 4102 30364 4108 30428
rect 4172 30426 4178 30428
rect 4797 30426 4863 30429
rect 4172 30424 4863 30426
rect 4172 30368 4802 30424
rect 4858 30368 4863 30424
rect 4172 30366 4863 30368
rect 4172 30364 4178 30366
rect 4797 30363 4863 30366
rect 5809 30426 5875 30429
rect 6678 30426 6684 30428
rect 5809 30424 6684 30426
rect 5809 30368 5814 30424
rect 5870 30368 6684 30424
rect 5809 30366 6684 30368
rect 5809 30363 5875 30366
rect 6678 30364 6684 30366
rect 6748 30426 6754 30428
rect 7465 30426 7531 30429
rect 6748 30424 7531 30426
rect 6748 30368 7470 30424
rect 7526 30368 7531 30424
rect 6748 30366 7531 30368
rect 6748 30364 6754 30366
rect 7465 30363 7531 30366
rect 2078 30228 2084 30292
rect 2148 30290 2154 30292
rect 2221 30290 2287 30293
rect 7189 30292 7255 30293
rect 2148 30288 2287 30290
rect 2148 30232 2226 30288
rect 2282 30232 2287 30288
rect 2148 30230 2287 30232
rect 2148 30228 2154 30230
rect 2221 30227 2287 30230
rect 2630 30228 2636 30292
rect 2700 30290 2706 30292
rect 5942 30290 5948 30292
rect 2700 30230 5948 30290
rect 2700 30228 2706 30230
rect 5942 30228 5948 30230
rect 6012 30228 6018 30292
rect 7189 30290 7236 30292
rect 7144 30288 7236 30290
rect 7144 30232 7194 30288
rect 7144 30230 7236 30232
rect 7189 30228 7236 30230
rect 7300 30228 7306 30292
rect 9254 30228 9260 30292
rect 9324 30290 9330 30292
rect 9765 30290 9831 30293
rect 9324 30288 9831 30290
rect 9324 30232 9770 30288
rect 9826 30232 9831 30288
rect 9324 30230 9831 30232
rect 9324 30228 9330 30230
rect 7189 30227 7255 30228
rect 9765 30227 9831 30230
rect 2313 30154 2379 30157
rect 2313 30152 5458 30154
rect 2313 30096 2318 30152
rect 2374 30096 5458 30152
rect 2313 30094 5458 30096
rect 2313 30091 2379 30094
rect 5398 30018 5458 30094
rect 5758 30092 5764 30156
rect 5828 30154 5834 30156
rect 7192 30154 7252 30227
rect 5828 30094 7252 30154
rect 7741 30154 7807 30157
rect 7741 30152 7850 30154
rect 7741 30096 7746 30152
rect 7802 30096 7850 30152
rect 5828 30092 5834 30094
rect 7741 30091 7850 30096
rect 7046 30018 7052 30020
rect 5398 29958 7052 30018
rect 7046 29956 7052 29958
rect 7116 29956 7122 30020
rect 4318 29952 4634 29953
rect 4318 29888 4324 29952
rect 4388 29888 4404 29952
rect 4468 29888 4484 29952
rect 4548 29888 4564 29952
rect 4628 29888 4634 29952
rect 4318 29887 4634 29888
rect 5625 29882 5691 29885
rect 6729 29882 6795 29885
rect 5582 29880 5691 29882
rect 5582 29824 5630 29880
rect 5686 29824 5691 29880
rect 5582 29819 5691 29824
rect 6686 29880 6795 29882
rect 6686 29824 6734 29880
rect 6790 29824 6795 29880
rect 6686 29819 6795 29824
rect 2078 29746 2084 29748
rect 1028 29686 2084 29746
rect 1028 29613 1088 29686
rect 2078 29684 2084 29686
rect 2148 29684 2154 29748
rect 2446 29684 2452 29748
rect 2516 29746 2522 29748
rect 2865 29746 2931 29749
rect 3141 29748 3207 29749
rect 3141 29746 3188 29748
rect 2516 29744 2931 29746
rect 2516 29688 2870 29744
rect 2926 29688 2931 29744
rect 2516 29686 2931 29688
rect 3096 29744 3188 29746
rect 3252 29746 3258 29748
rect 3877 29746 3943 29749
rect 4705 29746 4771 29749
rect 3252 29744 4771 29746
rect 3096 29688 3146 29744
rect 3252 29688 3882 29744
rect 3938 29688 4710 29744
rect 4766 29688 4771 29744
rect 3096 29686 3188 29688
rect 2516 29684 2522 29686
rect 2865 29683 2931 29686
rect 3141 29684 3188 29686
rect 3252 29686 4771 29688
rect 3252 29684 3258 29686
rect 3141 29683 3207 29684
rect 3877 29683 3943 29686
rect 4705 29683 4771 29686
rect 238 29548 244 29612
rect 308 29610 314 29612
rect 1025 29610 1091 29613
rect 308 29608 1091 29610
rect 308 29552 1030 29608
rect 1086 29552 1091 29608
rect 308 29550 1091 29552
rect 308 29548 314 29550
rect 1025 29547 1091 29550
rect 1209 29610 1275 29613
rect 1342 29610 1348 29612
rect 1209 29608 1348 29610
rect 1209 29552 1214 29608
rect 1270 29552 1348 29608
rect 1209 29550 1348 29552
rect 1209 29547 1275 29550
rect 1342 29548 1348 29550
rect 1412 29548 1418 29612
rect 5582 29610 5642 29819
rect 6686 29746 6746 29819
rect 5720 29686 6746 29746
rect 5720 29613 5780 29686
rect 7790 29613 7850 30091
rect 10718 29952 11034 29953
rect 10718 29888 10724 29952
rect 10788 29888 10804 29952
rect 10868 29888 10884 29952
rect 10948 29888 10964 29952
rect 11028 29888 11034 29952
rect 10718 29887 11034 29888
rect 2730 29550 5642 29610
rect 5717 29608 5783 29613
rect 5717 29552 5722 29608
rect 5778 29552 5783 29608
rect 1025 29474 1091 29477
rect 2730 29474 2790 29550
rect 5717 29547 5783 29552
rect 5942 29548 5948 29612
rect 6012 29610 6018 29612
rect 7097 29610 7163 29613
rect 6012 29608 7163 29610
rect 6012 29552 7102 29608
rect 7158 29552 7163 29608
rect 6012 29550 7163 29552
rect 7790 29608 7899 29613
rect 7790 29552 7838 29608
rect 7894 29552 7899 29608
rect 7790 29550 7899 29552
rect 6012 29548 6018 29550
rect 7097 29547 7163 29550
rect 7833 29547 7899 29550
rect 1025 29472 2790 29474
rect 1025 29416 1030 29472
rect 1086 29416 2790 29472
rect 1025 29414 2790 29416
rect 1025 29411 1091 29414
rect 4102 29412 4108 29476
rect 4172 29474 4178 29476
rect 5720 29474 5780 29547
rect 4172 29414 5780 29474
rect 4172 29412 4178 29414
rect 6310 29412 6316 29476
rect 6380 29474 6386 29476
rect 7281 29474 7347 29477
rect 8201 29474 8267 29477
rect 6380 29472 7347 29474
rect 6380 29416 7286 29472
rect 7342 29416 7347 29472
rect 6380 29414 7347 29416
rect 6380 29412 6386 29414
rect 7281 29411 7347 29414
rect 7468 29472 8267 29474
rect 7468 29416 8206 29472
rect 8262 29416 8267 29472
rect 7468 29414 8267 29416
rect 3658 29408 3974 29409
rect 3658 29344 3664 29408
rect 3728 29344 3744 29408
rect 3808 29344 3824 29408
rect 3888 29344 3904 29408
rect 3968 29344 3974 29408
rect 3658 29343 3974 29344
rect 974 29276 980 29340
rect 1044 29338 1050 29340
rect 2129 29338 2195 29341
rect 1044 29336 2195 29338
rect 1044 29280 2134 29336
rect 2190 29280 2195 29336
rect 1044 29278 2195 29280
rect 1044 29276 1050 29278
rect 2129 29275 2195 29278
rect 4838 29276 4844 29340
rect 4908 29338 4914 29340
rect 5257 29338 5323 29341
rect 4908 29336 5323 29338
rect 4908 29280 5262 29336
rect 5318 29280 5323 29336
rect 4908 29278 5323 29280
rect 4908 29276 4914 29278
rect 5257 29275 5323 29278
rect 5901 29338 5967 29341
rect 6545 29338 6611 29341
rect 5901 29336 6611 29338
rect 5901 29280 5906 29336
rect 5962 29280 6550 29336
rect 6606 29280 6611 29336
rect 5901 29278 6611 29280
rect 5901 29275 5967 29278
rect 6545 29275 6611 29278
rect 7097 29338 7163 29341
rect 7468 29338 7528 29414
rect 8201 29411 8267 29414
rect 10058 29408 10374 29409
rect 10058 29344 10064 29408
rect 10128 29344 10144 29408
rect 10208 29344 10224 29408
rect 10288 29344 10304 29408
rect 10368 29344 10374 29408
rect 10058 29343 10374 29344
rect 7097 29336 7528 29338
rect 7097 29280 7102 29336
rect 7158 29280 7528 29336
rect 7097 29278 7528 29280
rect 7606 29278 9690 29338
rect 7097 29275 7163 29278
rect 473 29202 539 29205
rect 2446 29202 2452 29204
rect 473 29200 2452 29202
rect 473 29144 478 29200
rect 534 29144 2452 29200
rect 473 29142 2452 29144
rect 473 29139 539 29142
rect 2446 29140 2452 29142
rect 2516 29140 2522 29204
rect 2865 29202 2931 29205
rect 3366 29202 3372 29204
rect 2865 29200 3372 29202
rect 2865 29144 2870 29200
rect 2926 29144 3372 29200
rect 2865 29142 3372 29144
rect 2865 29139 2931 29142
rect 3366 29140 3372 29142
rect 3436 29202 3442 29204
rect 3601 29202 3667 29205
rect 3436 29200 3667 29202
rect 3436 29144 3606 29200
rect 3662 29144 3667 29200
rect 3436 29142 3667 29144
rect 3436 29140 3442 29142
rect 3601 29139 3667 29142
rect 3969 29202 4035 29205
rect 4613 29202 4679 29205
rect 3969 29200 4679 29202
rect 3969 29144 3974 29200
rect 4030 29144 4618 29200
rect 4674 29144 4679 29200
rect 3969 29142 4679 29144
rect 3969 29139 4035 29142
rect 4613 29139 4679 29142
rect 4838 29140 4844 29204
rect 4908 29202 4914 29204
rect 5206 29202 5212 29204
rect 4908 29142 5212 29202
rect 4908 29140 4914 29142
rect 5206 29140 5212 29142
rect 5276 29140 5282 29204
rect 6453 29202 6519 29205
rect 7606 29202 7666 29278
rect 9438 29202 9444 29204
rect 6453 29200 7666 29202
rect 6453 29144 6458 29200
rect 6514 29144 7666 29200
rect 6453 29142 7666 29144
rect 7790 29142 9444 29202
rect 6453 29139 6519 29142
rect 657 29066 723 29069
rect 1526 29066 1532 29068
rect 657 29064 1532 29066
rect 657 29008 662 29064
rect 718 29008 1532 29064
rect 657 29006 1532 29008
rect 657 29003 723 29006
rect 1526 29004 1532 29006
rect 1596 29004 1602 29068
rect 2814 29004 2820 29068
rect 2884 29066 2890 29068
rect 6821 29066 6887 29069
rect 2884 29064 6887 29066
rect 2884 29008 6826 29064
rect 6882 29008 6887 29064
rect 2884 29006 6887 29008
rect 2884 29004 2890 29006
rect 6821 29003 6887 29006
rect 7189 29066 7255 29069
rect 7790 29068 7850 29142
rect 9438 29140 9444 29142
rect 9508 29140 9514 29204
rect 9630 29202 9690 29278
rect 11237 29202 11303 29205
rect 9630 29200 11303 29202
rect 9630 29144 11242 29200
rect 11298 29144 11303 29200
rect 9630 29142 11303 29144
rect 11237 29139 11303 29142
rect 7782 29066 7788 29068
rect 7189 29064 7788 29066
rect 7189 29008 7194 29064
rect 7250 29008 7788 29064
rect 7189 29006 7788 29008
rect 7189 29003 7255 29006
rect 7782 29004 7788 29006
rect 7852 29004 7858 29068
rect 8569 29066 8635 29069
rect 8702 29066 8708 29068
rect 8569 29064 8708 29066
rect 8569 29008 8574 29064
rect 8630 29008 8708 29064
rect 8569 29006 8708 29008
rect 8569 29003 8635 29006
rect 8702 29004 8708 29006
rect 8772 29004 8778 29068
rect 9121 29066 9187 29069
rect 9078 29064 9187 29066
rect 9078 29008 9126 29064
rect 9182 29008 9187 29064
rect 9078 29003 9187 29008
rect 0 28933 400 28960
rect 0 28928 447 28933
rect 2865 28930 2931 28933
rect 0 28872 386 28928
rect 442 28872 447 28928
rect 0 28867 447 28872
rect 1534 28928 2931 28930
rect 1534 28872 2870 28928
rect 2926 28872 2931 28928
rect 1534 28870 2931 28872
rect 0 28840 400 28867
rect 790 28732 796 28796
rect 860 28794 866 28796
rect 1301 28794 1367 28797
rect 860 28792 1367 28794
rect 860 28736 1306 28792
rect 1362 28736 1367 28792
rect 860 28734 1367 28736
rect 860 28732 866 28734
rect 1301 28731 1367 28734
rect 0 28658 400 28688
rect 657 28658 723 28661
rect 0 28656 723 28658
rect 0 28600 662 28656
rect 718 28600 723 28656
rect 0 28598 723 28600
rect 0 28568 400 28598
rect 657 28595 723 28598
rect 1301 28520 1367 28525
rect 1301 28464 1306 28520
rect 1362 28464 1367 28520
rect 1301 28459 1367 28464
rect 0 28386 400 28416
rect 1304 28386 1364 28459
rect 0 28326 1364 28386
rect 0 28296 400 28326
rect 0 28114 400 28144
rect 933 28114 999 28117
rect 0 28112 999 28114
rect 0 28056 938 28112
rect 994 28056 999 28112
rect 0 28054 999 28056
rect 0 28024 400 28054
rect 933 28051 999 28054
rect 1117 28114 1183 28117
rect 1117 28112 1456 28114
rect 1117 28056 1122 28112
rect 1178 28056 1456 28112
rect 1117 28054 1456 28056
rect 1117 28051 1183 28054
rect 933 27978 999 27981
rect 1158 27978 1164 27980
rect 933 27976 1164 27978
rect 933 27920 938 27976
rect 994 27920 1164 27976
rect 933 27918 1164 27920
rect 933 27915 999 27918
rect 1158 27916 1164 27918
rect 1228 27916 1234 27980
rect 1396 27845 1456 28054
rect 238 27780 244 27844
rect 308 27842 314 27844
rect 841 27842 907 27845
rect 1158 27842 1164 27844
rect 308 27840 1164 27842
rect 308 27784 846 27840
rect 902 27784 1164 27840
rect 308 27782 1164 27784
rect 308 27780 314 27782
rect 841 27779 907 27782
rect 1158 27780 1164 27782
rect 1228 27780 1234 27844
rect 1393 27840 1459 27845
rect 1393 27784 1398 27840
rect 1454 27784 1459 27840
rect 1393 27779 1459 27784
rect 238 27508 244 27572
rect 308 27570 314 27572
rect 1209 27570 1275 27573
rect 308 27568 1275 27570
rect 308 27512 1214 27568
rect 1270 27512 1275 27568
rect 308 27510 1275 27512
rect 308 27508 314 27510
rect 1209 27507 1275 27510
rect 1393 27570 1459 27573
rect 1534 27570 1594 28870
rect 2865 28867 2931 28870
rect 3366 28868 3372 28932
rect 3436 28930 3442 28932
rect 3601 28930 3667 28933
rect 3436 28928 3667 28930
rect 3436 28872 3606 28928
rect 3662 28872 3667 28928
rect 3436 28870 3667 28872
rect 3436 28868 3442 28870
rect 3601 28867 3667 28870
rect 4981 28932 5047 28933
rect 4981 28928 5028 28932
rect 5092 28930 5098 28932
rect 5809 28930 5875 28933
rect 6361 28930 6427 28933
rect 4981 28872 4986 28928
rect 4981 28868 5028 28872
rect 5092 28870 5138 28930
rect 5809 28928 6427 28930
rect 5809 28872 5814 28928
rect 5870 28872 6366 28928
rect 6422 28872 6427 28928
rect 5809 28870 6427 28872
rect 5092 28868 5098 28870
rect 4981 28867 5047 28868
rect 5809 28867 5875 28870
rect 6361 28867 6427 28870
rect 6913 28930 6979 28933
rect 8017 28930 8083 28933
rect 6913 28928 8083 28930
rect 6913 28872 6918 28928
rect 6974 28872 8022 28928
rect 8078 28872 8083 28928
rect 6913 28870 8083 28872
rect 6913 28867 6979 28870
rect 8017 28867 8083 28870
rect 4318 28864 4634 28865
rect 4318 28800 4324 28864
rect 4388 28800 4404 28864
rect 4468 28800 4484 28864
rect 4548 28800 4564 28864
rect 4628 28800 4634 28864
rect 4318 28799 4634 28800
rect 1945 28794 2011 28797
rect 2262 28794 2268 28796
rect 1945 28792 2268 28794
rect 1945 28736 1950 28792
rect 2006 28736 2268 28792
rect 1945 28734 2268 28736
rect 1945 28731 2011 28734
rect 2262 28732 2268 28734
rect 2332 28794 2338 28796
rect 2497 28794 2563 28797
rect 2332 28792 2563 28794
rect 2332 28736 2502 28792
rect 2558 28736 2563 28792
rect 2332 28734 2563 28736
rect 2332 28732 2338 28734
rect 2497 28731 2563 28734
rect 2814 28732 2820 28796
rect 2884 28794 2890 28796
rect 4102 28794 4108 28796
rect 2884 28734 4108 28794
rect 2884 28732 2890 28734
rect 4102 28732 4108 28734
rect 4172 28732 4178 28796
rect 4981 28794 5047 28797
rect 6126 28794 6132 28796
rect 4981 28792 6132 28794
rect 4981 28736 4986 28792
rect 5042 28736 6132 28792
rect 4981 28734 6132 28736
rect 4981 28731 5047 28734
rect 6126 28732 6132 28734
rect 6196 28794 6202 28796
rect 9078 28794 9138 29003
rect 10718 28864 11034 28865
rect 10718 28800 10724 28864
rect 10788 28800 10804 28864
rect 10868 28800 10884 28864
rect 10948 28800 10964 28864
rect 11028 28800 11034 28864
rect 10718 28799 11034 28800
rect 9489 28794 9555 28797
rect 6196 28792 9555 28794
rect 6196 28736 9494 28792
rect 9550 28736 9555 28792
rect 6196 28734 9555 28736
rect 6196 28732 6202 28734
rect 9489 28731 9555 28734
rect 2773 28658 2839 28661
rect 5441 28658 5507 28661
rect 6310 28658 6316 28660
rect 2773 28656 6316 28658
rect 2773 28600 2778 28656
rect 2834 28600 5446 28656
rect 5502 28600 6316 28656
rect 2773 28598 6316 28600
rect 2773 28595 2839 28598
rect 5441 28595 5507 28598
rect 6310 28596 6316 28598
rect 6380 28658 6386 28660
rect 7649 28658 7715 28661
rect 6380 28656 7715 28658
rect 6380 28600 7654 28656
rect 7710 28600 7715 28656
rect 6380 28598 7715 28600
rect 6380 28596 6386 28598
rect 7649 28595 7715 28598
rect 9397 28656 9463 28661
rect 9397 28600 9402 28656
rect 9458 28600 9463 28656
rect 9397 28595 9463 28600
rect 2681 28522 2747 28525
rect 2998 28522 3004 28524
rect 2681 28520 3004 28522
rect 2681 28464 2686 28520
rect 2742 28464 3004 28520
rect 2681 28462 3004 28464
rect 2681 28459 2747 28462
rect 2998 28460 3004 28462
rect 3068 28460 3074 28524
rect 3366 28460 3372 28524
rect 3436 28522 3442 28524
rect 3601 28522 3667 28525
rect 3436 28520 3667 28522
rect 3436 28464 3606 28520
rect 3662 28464 3667 28520
rect 3436 28462 3667 28464
rect 3436 28460 3442 28462
rect 3601 28459 3667 28462
rect 3969 28522 4035 28525
rect 4102 28522 4108 28524
rect 3969 28520 4108 28522
rect 3969 28464 3974 28520
rect 4030 28464 4108 28520
rect 3969 28462 4108 28464
rect 3969 28459 4035 28462
rect 4102 28460 4108 28462
rect 4172 28460 4178 28524
rect 5533 28522 5599 28525
rect 6913 28522 6979 28525
rect 7373 28524 7439 28525
rect 7373 28522 7420 28524
rect 5533 28520 6979 28522
rect 5533 28464 5538 28520
rect 5594 28464 6918 28520
rect 6974 28464 6979 28520
rect 5533 28462 6979 28464
rect 7332 28520 7420 28522
rect 7484 28522 7490 28524
rect 9400 28522 9460 28595
rect 10133 28522 10199 28525
rect 7332 28464 7378 28520
rect 7332 28462 7420 28464
rect 5533 28459 5599 28462
rect 6913 28459 6979 28462
rect 7373 28460 7420 28462
rect 7484 28462 9460 28522
rect 9630 28520 10199 28522
rect 9630 28464 10138 28520
rect 10194 28464 10199 28520
rect 9630 28462 10199 28464
rect 7484 28460 7490 28462
rect 7373 28459 7439 28460
rect 2078 28324 2084 28388
rect 2148 28386 2154 28388
rect 6494 28386 6500 28388
rect 2148 28326 3434 28386
rect 2148 28324 2154 28326
rect 2078 28188 2084 28252
rect 2148 28250 2154 28252
rect 2589 28250 2655 28253
rect 2865 28250 2931 28253
rect 2148 28248 2655 28250
rect 2148 28192 2594 28248
rect 2650 28192 2655 28248
rect 2148 28190 2655 28192
rect 2148 28188 2154 28190
rect 2589 28187 2655 28190
rect 2822 28248 2931 28250
rect 2822 28192 2870 28248
rect 2926 28192 2931 28248
rect 2822 28187 2931 28192
rect 2998 28188 3004 28252
rect 3068 28250 3074 28252
rect 3068 28190 3296 28250
rect 3068 28188 3074 28190
rect 2129 27978 2195 27981
rect 2589 27978 2655 27981
rect 2129 27976 2655 27978
rect 2129 27920 2134 27976
rect 2190 27920 2594 27976
rect 2650 27920 2655 27976
rect 2129 27918 2655 27920
rect 2129 27915 2195 27918
rect 2589 27915 2655 27918
rect 2822 27845 2882 28187
rect 2822 27840 2931 27845
rect 2822 27784 2870 27840
rect 2926 27784 2931 27840
rect 2822 27782 2931 27784
rect 3236 27842 3296 28190
rect 3374 28114 3434 28326
rect 4110 28326 6500 28386
rect 3658 28320 3974 28321
rect 3658 28256 3664 28320
rect 3728 28256 3744 28320
rect 3808 28256 3824 28320
rect 3888 28256 3904 28320
rect 3968 28256 3974 28320
rect 3658 28255 3974 28256
rect 4110 28114 4170 28326
rect 6494 28324 6500 28326
rect 6564 28324 6570 28388
rect 7097 28386 7163 28389
rect 8201 28386 8267 28389
rect 7097 28384 8267 28386
rect 7097 28328 7102 28384
rect 7158 28328 8206 28384
rect 8262 28328 8267 28384
rect 7097 28326 8267 28328
rect 7097 28323 7163 28326
rect 8201 28323 8267 28326
rect 9489 28386 9555 28389
rect 9630 28386 9690 28462
rect 10133 28459 10199 28462
rect 9489 28384 9690 28386
rect 9489 28328 9494 28384
rect 9550 28328 9690 28384
rect 9489 28326 9690 28328
rect 9489 28323 9555 28326
rect 10058 28320 10374 28321
rect 10058 28256 10064 28320
rect 10128 28256 10144 28320
rect 10208 28256 10224 28320
rect 10288 28256 10304 28320
rect 10368 28256 10374 28320
rect 10058 28255 10374 28256
rect 6177 28250 6243 28253
rect 8201 28250 8267 28253
rect 6177 28248 8267 28250
rect 6177 28192 6182 28248
rect 6238 28192 8206 28248
rect 8262 28192 8267 28248
rect 6177 28190 8267 28192
rect 6177 28187 6243 28190
rect 8201 28187 8267 28190
rect 3374 28054 4170 28114
rect 4797 28114 4863 28117
rect 4981 28114 5047 28117
rect 6177 28116 6243 28117
rect 6126 28114 6132 28116
rect 4797 28112 5047 28114
rect 4797 28056 4802 28112
rect 4858 28056 4986 28112
rect 5042 28056 5047 28112
rect 4797 28054 5047 28056
rect 6086 28054 6132 28114
rect 6196 28112 6243 28116
rect 6238 28056 6243 28112
rect 4797 28051 4863 28054
rect 4981 28051 5047 28054
rect 6126 28052 6132 28054
rect 6196 28052 6243 28056
rect 6177 28051 6243 28052
rect 4613 27978 4679 27981
rect 4156 27976 4679 27978
rect 4156 27920 4618 27976
rect 4674 27920 4679 27976
rect 4156 27918 4679 27920
rect 4984 27978 5044 28051
rect 6453 27978 6519 27981
rect 6913 27978 6979 27981
rect 4984 27976 6979 27978
rect 4984 27920 6458 27976
rect 6514 27920 6918 27976
rect 6974 27920 6979 27976
rect 4984 27918 6979 27920
rect 3877 27842 3943 27845
rect 3236 27840 3943 27842
rect 3236 27784 3882 27840
rect 3938 27784 3943 27840
rect 3236 27782 3943 27784
rect 2865 27779 2931 27782
rect 3877 27779 3943 27782
rect 2129 27706 2195 27709
rect 2681 27706 2747 27709
rect 2129 27704 2747 27706
rect 2129 27648 2134 27704
rect 2190 27648 2686 27704
rect 2742 27648 2747 27704
rect 2129 27646 2747 27648
rect 2129 27643 2195 27646
rect 2681 27643 2747 27646
rect 3182 27644 3188 27708
rect 3252 27706 3258 27708
rect 3693 27706 3759 27709
rect 3252 27704 3759 27706
rect 3252 27648 3698 27704
rect 3754 27648 3759 27704
rect 3252 27646 3759 27648
rect 3252 27644 3258 27646
rect 3693 27643 3759 27646
rect 1393 27568 1594 27570
rect 1393 27512 1398 27568
rect 1454 27512 1594 27568
rect 1393 27510 1594 27512
rect 1945 27570 2011 27573
rect 4156 27570 4216 27918
rect 4613 27915 4679 27918
rect 6453 27915 6519 27918
rect 6913 27915 6979 27918
rect 8518 27916 8524 27980
rect 8588 27978 8594 27980
rect 9121 27978 9187 27981
rect 8588 27976 9187 27978
rect 8588 27920 9126 27976
rect 9182 27920 9187 27976
rect 8588 27918 9187 27920
rect 8588 27916 8594 27918
rect 9121 27915 9187 27918
rect 10542 27916 10548 27980
rect 10612 27978 10618 27980
rect 11053 27978 11119 27981
rect 10612 27976 11119 27978
rect 10612 27920 11058 27976
rect 11114 27920 11119 27976
rect 10612 27918 11119 27920
rect 10612 27916 10618 27918
rect 11053 27915 11119 27918
rect 5993 27842 6059 27845
rect 7189 27842 7255 27845
rect 5993 27840 7255 27842
rect 5993 27784 5998 27840
rect 6054 27784 7194 27840
rect 7250 27784 7255 27840
rect 5993 27782 7255 27784
rect 5993 27779 6059 27782
rect 7189 27779 7255 27782
rect 4318 27776 4634 27777
rect 4318 27712 4324 27776
rect 4388 27712 4404 27776
rect 4468 27712 4484 27776
rect 4548 27712 4564 27776
rect 4628 27712 4634 27776
rect 4318 27711 4634 27712
rect 10718 27776 11034 27777
rect 10718 27712 10724 27776
rect 10788 27712 10804 27776
rect 10868 27712 10884 27776
rect 10948 27712 10964 27776
rect 11028 27712 11034 27776
rect 10718 27711 11034 27712
rect 5625 27706 5691 27709
rect 6729 27706 6795 27709
rect 5625 27704 6795 27706
rect 5625 27648 5630 27704
rect 5686 27648 6734 27704
rect 6790 27648 6795 27704
rect 5625 27646 6795 27648
rect 5625 27643 5691 27646
rect 6729 27643 6795 27646
rect 7373 27706 7439 27709
rect 7598 27706 7604 27708
rect 7373 27704 7604 27706
rect 7373 27648 7378 27704
rect 7434 27648 7604 27704
rect 7373 27646 7604 27648
rect 7373 27643 7439 27646
rect 7598 27644 7604 27646
rect 7668 27644 7674 27708
rect 8201 27706 8267 27709
rect 8201 27704 9690 27706
rect 8201 27648 8206 27704
rect 8262 27648 9690 27704
rect 8201 27646 9690 27648
rect 8201 27643 8267 27646
rect 1945 27568 4216 27570
rect 1945 27512 1950 27568
rect 2006 27512 4216 27568
rect 1945 27510 4216 27512
rect 1393 27507 1459 27510
rect 1945 27507 2011 27510
rect 606 27372 612 27436
rect 676 27434 682 27436
rect 1577 27434 1643 27437
rect 3509 27434 3575 27437
rect 676 27432 1643 27434
rect 676 27376 1582 27432
rect 1638 27376 1643 27432
rect 676 27374 1643 27376
rect 676 27372 682 27374
rect 1577 27371 1643 27374
rect 1764 27432 3575 27434
rect 1764 27376 3514 27432
rect 3570 27376 3575 27432
rect 1764 27374 3575 27376
rect 4156 27434 4216 27510
rect 4521 27570 4587 27573
rect 7281 27570 7347 27573
rect 4521 27568 7347 27570
rect 4521 27512 4526 27568
rect 4582 27512 7286 27568
rect 7342 27512 7347 27568
rect 4521 27510 7347 27512
rect 4521 27507 4587 27510
rect 7281 27507 7347 27510
rect 8017 27570 8083 27573
rect 8569 27570 8635 27573
rect 8937 27570 9003 27573
rect 8017 27568 8448 27570
rect 8017 27512 8022 27568
rect 8078 27512 8448 27568
rect 8017 27510 8448 27512
rect 8017 27507 8083 27510
rect 5206 27434 5212 27436
rect 4156 27374 5212 27434
rect 1577 27298 1643 27301
rect 1764 27298 1824 27374
rect 3509 27371 3575 27374
rect 5206 27372 5212 27374
rect 5276 27434 5282 27436
rect 8388 27434 8448 27510
rect 8569 27568 9003 27570
rect 8569 27512 8574 27568
rect 8630 27512 8942 27568
rect 8998 27512 9003 27568
rect 8569 27510 9003 27512
rect 9630 27570 9690 27646
rect 10685 27570 10751 27573
rect 9630 27568 10751 27570
rect 9630 27512 10690 27568
rect 10746 27512 10751 27568
rect 9630 27510 10751 27512
rect 8569 27507 8635 27510
rect 8937 27507 9003 27510
rect 10685 27507 10751 27510
rect 9121 27434 9187 27437
rect 5276 27374 7068 27434
rect 5276 27372 5282 27374
rect 1577 27296 1824 27298
rect 1577 27240 1582 27296
rect 1638 27240 1824 27296
rect 1577 27238 1824 27240
rect 2681 27298 2747 27301
rect 4613 27298 4679 27301
rect 5206 27298 5212 27300
rect 2681 27296 3296 27298
rect 2681 27240 2686 27296
rect 2742 27240 3296 27296
rect 2681 27238 3296 27240
rect 1577 27235 1643 27238
rect 2681 27235 2747 27238
rect 3236 27165 3296 27238
rect 4613 27296 5212 27298
rect 4613 27240 4618 27296
rect 4674 27240 5212 27296
rect 4613 27238 5212 27240
rect 4613 27235 4679 27238
rect 5206 27236 5212 27238
rect 5276 27236 5282 27300
rect 5809 27298 5875 27301
rect 5942 27298 5948 27300
rect 5809 27296 5948 27298
rect 5809 27240 5814 27296
rect 5870 27240 5948 27296
rect 5809 27238 5948 27240
rect 5809 27235 5875 27238
rect 5942 27236 5948 27238
rect 6012 27298 6018 27300
rect 6269 27298 6335 27301
rect 6012 27296 6335 27298
rect 6012 27240 6274 27296
rect 6330 27240 6335 27296
rect 6012 27238 6335 27240
rect 6012 27236 6018 27238
rect 6269 27235 6335 27238
rect 3658 27232 3974 27233
rect 3658 27168 3664 27232
rect 3728 27168 3744 27232
rect 3808 27168 3824 27232
rect 3888 27168 3904 27232
rect 3968 27168 3974 27232
rect 3658 27167 3974 27168
rect 1117 27162 1183 27165
rect 3049 27162 3115 27165
rect 1117 27160 3115 27162
rect 1117 27104 1122 27160
rect 1178 27104 3054 27160
rect 3110 27104 3115 27160
rect 1117 27102 3115 27104
rect 1117 27099 1183 27102
rect 3049 27099 3115 27102
rect 3233 27160 3299 27165
rect 3233 27104 3238 27160
rect 3294 27104 3299 27160
rect 3233 27099 3299 27104
rect 4337 27162 4403 27165
rect 5758 27162 5764 27164
rect 4337 27160 5764 27162
rect 4337 27104 4342 27160
rect 4398 27104 5764 27160
rect 4337 27102 5764 27104
rect 4337 27099 4403 27102
rect 5758 27100 5764 27102
rect 5828 27100 5834 27164
rect 105 27026 171 27029
rect 1894 27026 1900 27028
rect 105 27024 1900 27026
rect 105 26968 110 27024
rect 166 26968 1900 27024
rect 105 26966 1900 26968
rect 105 26963 171 26966
rect 1894 26964 1900 26966
rect 1964 27026 1970 27028
rect 2405 27026 2471 27029
rect 1964 27024 2471 27026
rect 1964 26968 2410 27024
rect 2466 26968 2471 27024
rect 1964 26966 2471 26968
rect 1964 26964 1970 26966
rect 2405 26963 2471 26966
rect 2589 27026 2655 27029
rect 3325 27026 3391 27029
rect 2589 27024 6010 27026
rect 2589 26968 2594 27024
rect 2650 26968 3330 27024
rect 3386 26968 6010 27024
rect 2589 26966 6010 26968
rect 2589 26963 2655 26966
rect 3325 26963 3391 26966
rect 1025 26890 1091 26893
rect 3366 26890 3372 26892
rect 1025 26888 3372 26890
rect 1025 26832 1030 26888
rect 1086 26832 3372 26888
rect 1025 26830 3372 26832
rect 1025 26827 1091 26830
rect 3366 26828 3372 26830
rect 3436 26828 3442 26892
rect 4337 26890 4403 26893
rect 4337 26888 4952 26890
rect 4337 26832 4342 26888
rect 4398 26832 4952 26888
rect 4337 26830 4952 26832
rect 4337 26827 4403 26830
rect 4892 26757 4952 26830
rect 3366 26692 3372 26756
rect 3436 26754 3442 26756
rect 4061 26754 4127 26757
rect 3436 26752 4127 26754
rect 3436 26696 4066 26752
rect 4122 26696 4127 26752
rect 3436 26694 4127 26696
rect 3436 26692 3442 26694
rect 4061 26691 4127 26694
rect 4889 26752 4955 26757
rect 4889 26696 4894 26752
rect 4950 26696 4955 26752
rect 4889 26691 4955 26696
rect 5574 26692 5580 26756
rect 5644 26754 5650 26756
rect 5809 26754 5875 26757
rect 5644 26752 5875 26754
rect 5644 26696 5814 26752
rect 5870 26696 5875 26752
rect 5644 26694 5875 26696
rect 5950 26754 6010 26966
rect 6310 26964 6316 27028
rect 6380 27026 6386 27028
rect 6453 27026 6519 27029
rect 6380 27024 6519 27026
rect 6380 26968 6458 27024
rect 6514 26968 6519 27024
rect 6380 26966 6519 26968
rect 6380 26964 6386 26966
rect 6453 26963 6519 26966
rect 7008 26893 7068 27374
rect 8388 27432 9187 27434
rect 8388 27376 9126 27432
rect 9182 27376 9187 27432
rect 8388 27374 9187 27376
rect 8109 27162 8175 27165
rect 8388 27162 8448 27374
rect 9121 27371 9187 27374
rect 10133 27434 10199 27437
rect 10542 27434 10548 27436
rect 10133 27432 10548 27434
rect 10133 27376 10138 27432
rect 10194 27376 10548 27432
rect 10133 27374 10548 27376
rect 10133 27371 10199 27374
rect 10542 27372 10548 27374
rect 10612 27372 10618 27436
rect 8937 27298 9003 27301
rect 9438 27298 9444 27300
rect 8937 27296 9444 27298
rect 8937 27240 8942 27296
rect 8998 27240 9444 27296
rect 8937 27238 9444 27240
rect 8937 27235 9003 27238
rect 9438 27236 9444 27238
rect 9508 27236 9514 27300
rect 10058 27232 10374 27233
rect 10058 27168 10064 27232
rect 10128 27168 10144 27232
rect 10208 27168 10224 27232
rect 10288 27168 10304 27232
rect 10368 27168 10374 27232
rect 10058 27167 10374 27168
rect 8109 27160 8448 27162
rect 8109 27104 8114 27160
rect 8170 27104 8448 27160
rect 8109 27102 8448 27104
rect 8109 27099 8175 27102
rect 7189 27026 7255 27029
rect 8569 27026 8635 27029
rect 10041 27026 10107 27029
rect 7189 27024 10107 27026
rect 7189 26968 7194 27024
rect 7250 26968 8574 27024
rect 8630 26968 10046 27024
rect 10102 26968 10107 27024
rect 7189 26966 10107 26968
rect 7189 26963 7255 26966
rect 8569 26963 8635 26966
rect 10041 26963 10107 26966
rect 7005 26888 7071 26893
rect 7005 26832 7010 26888
rect 7066 26832 7071 26888
rect 7005 26827 7071 26832
rect 9121 26890 9187 26893
rect 9254 26890 9260 26892
rect 9121 26888 9260 26890
rect 9121 26832 9126 26888
rect 9182 26832 9260 26888
rect 9121 26830 9260 26832
rect 9121 26827 9187 26830
rect 9254 26828 9260 26830
rect 9324 26828 9330 26892
rect 10685 26890 10751 26893
rect 11278 26890 11284 26892
rect 10685 26888 11284 26890
rect 10685 26832 10690 26888
rect 10746 26832 11284 26888
rect 10685 26830 11284 26832
rect 10685 26827 10751 26830
rect 11278 26828 11284 26830
rect 11348 26828 11354 26892
rect 6913 26754 6979 26757
rect 8569 26754 8635 26757
rect 5950 26752 8635 26754
rect 5950 26696 6918 26752
rect 6974 26696 8574 26752
rect 8630 26696 8635 26752
rect 5950 26694 8635 26696
rect 5644 26692 5650 26694
rect 5809 26691 5875 26694
rect 6913 26691 6979 26694
rect 8569 26691 8635 26694
rect 4318 26688 4634 26689
rect 4318 26624 4324 26688
rect 4388 26624 4404 26688
rect 4468 26624 4484 26688
rect 4548 26624 4564 26688
rect 4628 26624 4634 26688
rect 4318 26623 4634 26624
rect 10718 26688 11034 26689
rect 10718 26624 10724 26688
rect 10788 26624 10804 26688
rect 10868 26624 10884 26688
rect 10948 26624 10964 26688
rect 11028 26624 11034 26688
rect 10718 26623 11034 26624
rect 1577 26618 1643 26621
rect 3785 26618 3851 26621
rect 1577 26616 2330 26618
rect 1577 26560 1582 26616
rect 1638 26560 2330 26616
rect 1577 26558 2330 26560
rect 1577 26555 1643 26558
rect 1669 26482 1735 26485
rect 2078 26482 2084 26484
rect 1669 26480 2084 26482
rect 1669 26424 1674 26480
rect 1730 26424 2084 26480
rect 1669 26422 2084 26424
rect 1669 26419 1735 26422
rect 2078 26420 2084 26422
rect 2148 26420 2154 26484
rect 1342 26148 1348 26212
rect 1412 26210 1418 26212
rect 1669 26210 1735 26213
rect 1412 26208 1735 26210
rect 1412 26152 1674 26208
rect 1730 26152 1735 26208
rect 1412 26150 1735 26152
rect 1412 26148 1418 26150
rect 1669 26147 1735 26150
rect 2270 26077 2330 26558
rect 2500 26616 3851 26618
rect 2500 26560 3790 26616
rect 3846 26560 3851 26616
rect 2500 26558 3851 26560
rect 2500 26349 2560 26558
rect 3785 26555 3851 26558
rect 4153 26616 4219 26621
rect 4153 26560 4158 26616
rect 4214 26560 4219 26616
rect 4153 26555 4219 26560
rect 5574 26556 5580 26620
rect 5644 26618 5650 26620
rect 6453 26618 6519 26621
rect 5644 26616 6519 26618
rect 5644 26560 6458 26616
rect 6514 26560 6519 26616
rect 5644 26558 6519 26560
rect 5644 26556 5650 26558
rect 6453 26555 6519 26558
rect 6729 26618 6795 26621
rect 10542 26618 10548 26620
rect 6729 26616 10548 26618
rect 6729 26560 6734 26616
rect 6790 26560 10548 26616
rect 6729 26558 10548 26560
rect 6729 26555 6795 26558
rect 10542 26556 10548 26558
rect 10612 26556 10618 26620
rect 11094 26556 11100 26620
rect 11164 26618 11170 26620
rect 11237 26618 11303 26621
rect 11164 26616 11303 26618
rect 11164 26560 11242 26616
rect 11298 26560 11303 26616
rect 11164 26558 11303 26560
rect 11164 26556 11170 26558
rect 11237 26555 11303 26558
rect 2681 26482 2747 26485
rect 3325 26482 3391 26485
rect 2681 26480 3391 26482
rect 2681 26424 2686 26480
rect 2742 26424 3330 26480
rect 3386 26424 3391 26480
rect 2681 26422 3391 26424
rect 2681 26419 2747 26422
rect 3325 26419 3391 26422
rect 3969 26482 4035 26485
rect 4156 26482 4216 26555
rect 3969 26480 4216 26482
rect 3969 26424 3974 26480
rect 4030 26424 4216 26480
rect 3969 26422 4216 26424
rect 4429 26482 4495 26485
rect 5901 26482 5967 26485
rect 4429 26480 5967 26482
rect 4429 26424 4434 26480
rect 4490 26424 5906 26480
rect 5962 26424 5967 26480
rect 4429 26422 5967 26424
rect 3969 26419 4035 26422
rect 4429 26419 4495 26422
rect 5901 26419 5967 26422
rect 7046 26420 7052 26484
rect 7116 26482 7122 26484
rect 7189 26482 7255 26485
rect 7116 26480 7255 26482
rect 7116 26424 7194 26480
rect 7250 26424 7255 26480
rect 7116 26422 7255 26424
rect 7116 26420 7122 26422
rect 7189 26419 7255 26422
rect 8017 26482 8083 26485
rect 9581 26482 9647 26485
rect 8017 26480 9647 26482
rect 8017 26424 8022 26480
rect 8078 26424 9586 26480
rect 9642 26424 9647 26480
rect 8017 26422 9647 26424
rect 8017 26419 8083 26422
rect 9581 26419 9647 26422
rect 2497 26344 2563 26349
rect 4838 26346 4844 26348
rect 2497 26288 2502 26344
rect 2558 26288 2563 26344
rect 2497 26283 2563 26288
rect 3328 26286 4844 26346
rect 2405 26210 2471 26213
rect 3049 26210 3115 26213
rect 3182 26210 3188 26212
rect 2405 26208 3188 26210
rect 2405 26152 2410 26208
rect 2466 26152 3054 26208
rect 3110 26152 3188 26208
rect 2405 26150 3188 26152
rect 2405 26147 2471 26150
rect 3049 26147 3115 26150
rect 3182 26148 3188 26150
rect 3252 26148 3258 26212
rect 13 26074 79 26077
rect 1710 26074 1716 26076
rect 13 26072 1716 26074
rect 13 26016 18 26072
rect 74 26016 1716 26072
rect 13 26014 1716 26016
rect 13 26011 79 26014
rect 1710 26012 1716 26014
rect 1780 26012 1786 26076
rect 2270 26072 2379 26077
rect 2270 26016 2318 26072
rect 2374 26016 2379 26072
rect 2270 26014 2379 26016
rect 2313 26011 2379 26014
rect 3182 26012 3188 26076
rect 3252 26074 3258 26076
rect 3328 26074 3388 26286
rect 4838 26284 4844 26286
rect 4908 26284 4914 26348
rect 5073 26346 5139 26349
rect 6310 26346 6316 26348
rect 5073 26344 6316 26346
rect 5073 26288 5078 26344
rect 5134 26288 6316 26344
rect 5073 26286 6316 26288
rect 5073 26283 5139 26286
rect 6310 26284 6316 26286
rect 6380 26284 6386 26348
rect 8150 26346 8156 26348
rect 6456 26286 8156 26346
rect 4521 26210 4587 26213
rect 4700 26210 4706 26212
rect 4521 26208 4706 26210
rect 4521 26152 4526 26208
rect 4582 26152 4706 26208
rect 4521 26150 4706 26152
rect 4521 26147 4587 26150
rect 4700 26148 4706 26150
rect 4770 26148 4776 26212
rect 5758 26148 5764 26212
rect 5828 26210 5834 26212
rect 6456 26210 6516 26286
rect 8150 26284 8156 26286
rect 8220 26284 8226 26348
rect 8886 26284 8892 26348
rect 8956 26346 8962 26348
rect 9305 26346 9371 26349
rect 10041 26346 10107 26349
rect 8956 26344 9371 26346
rect 8956 26288 9310 26344
rect 9366 26288 9371 26344
rect 8956 26286 9371 26288
rect 8956 26284 8962 26286
rect 9305 26283 9371 26286
rect 9676 26344 10107 26346
rect 9676 26288 10046 26344
rect 10102 26288 10107 26344
rect 9676 26286 10107 26288
rect 5828 26150 6516 26210
rect 6637 26210 6703 26213
rect 7465 26210 7531 26213
rect 6637 26208 7531 26210
rect 6637 26152 6642 26208
rect 6698 26152 7470 26208
rect 7526 26152 7531 26208
rect 6637 26150 7531 26152
rect 5828 26148 5834 26150
rect 6637 26147 6703 26150
rect 7465 26147 7531 26150
rect 7925 26210 7991 26213
rect 8150 26210 8156 26212
rect 7925 26208 8156 26210
rect 7925 26152 7930 26208
rect 7986 26152 8156 26208
rect 7925 26150 8156 26152
rect 7925 26147 7991 26150
rect 8150 26148 8156 26150
rect 8220 26148 8226 26212
rect 3658 26144 3974 26145
rect 3658 26080 3664 26144
rect 3728 26080 3744 26144
rect 3808 26080 3824 26144
rect 3888 26080 3904 26144
rect 3968 26080 3974 26144
rect 3658 26079 3974 26080
rect 3252 26014 3388 26074
rect 4613 26074 4679 26077
rect 4981 26074 5047 26077
rect 4613 26072 5047 26074
rect 4613 26016 4618 26072
rect 4674 26016 4986 26072
rect 5042 26016 5047 26072
rect 4613 26014 5047 26016
rect 3252 26012 3258 26014
rect 4613 26011 4679 26014
rect 4981 26011 5047 26014
rect 5349 26074 5415 26077
rect 5717 26074 5783 26077
rect 8334 26074 8340 26076
rect 5349 26072 5642 26074
rect 5349 26016 5354 26072
rect 5410 26016 5642 26072
rect 5349 26014 5642 26016
rect 5349 26011 5415 26014
rect 1393 25938 1459 25941
rect 1526 25938 1532 25940
rect 1393 25936 1532 25938
rect 1393 25880 1398 25936
rect 1454 25880 1532 25936
rect 1393 25878 1532 25880
rect 1393 25875 1459 25878
rect 1526 25876 1532 25878
rect 1596 25876 1602 25940
rect 1710 25876 1716 25940
rect 1780 25938 1786 25940
rect 2221 25938 2287 25941
rect 1780 25936 2287 25938
rect 1780 25880 2226 25936
rect 2282 25880 2287 25936
rect 1780 25878 2287 25880
rect 1780 25876 1786 25878
rect 2221 25875 2287 25878
rect 2957 25938 3023 25941
rect 3509 25938 3575 25941
rect 2957 25936 3575 25938
rect 2957 25880 2962 25936
rect 3018 25880 3514 25936
rect 3570 25880 3575 25936
rect 2957 25878 3575 25880
rect 2957 25875 3023 25878
rect 3509 25875 3575 25878
rect 3693 25938 3759 25941
rect 3969 25938 4035 25941
rect 5257 25938 5323 25941
rect 3693 25936 3802 25938
rect 3693 25880 3698 25936
rect 3754 25880 3802 25936
rect 3693 25875 3802 25880
rect 3969 25936 5323 25938
rect 3969 25880 3974 25936
rect 4030 25880 5262 25936
rect 5318 25880 5323 25936
rect 3969 25878 5323 25880
rect 5582 25938 5642 26014
rect 5717 26072 8340 26074
rect 5717 26016 5722 26072
rect 5778 26016 8340 26072
rect 5717 26014 8340 26016
rect 5717 26011 5783 26014
rect 8334 26012 8340 26014
rect 8404 26012 8410 26076
rect 5717 25938 5783 25941
rect 5582 25936 5783 25938
rect 5582 25880 5722 25936
rect 5778 25880 5783 25936
rect 5582 25878 5783 25880
rect 3969 25875 4035 25878
rect 5257 25875 5323 25878
rect 5717 25875 5783 25878
rect 6085 25938 6151 25941
rect 6494 25938 6500 25940
rect 6085 25936 6500 25938
rect 6085 25880 6090 25936
rect 6146 25880 6500 25936
rect 6085 25878 6500 25880
rect 6085 25875 6151 25878
rect 6494 25876 6500 25878
rect 6564 25876 6570 25940
rect 7833 25938 7899 25941
rect 7966 25938 7972 25940
rect 7833 25936 7972 25938
rect 7833 25880 7838 25936
rect 7894 25880 7972 25936
rect 7833 25878 7972 25880
rect 7833 25875 7899 25878
rect 7966 25876 7972 25878
rect 8036 25876 8042 25940
rect 1025 25802 1091 25805
rect 1342 25802 1348 25804
rect 1025 25800 1348 25802
rect 1025 25744 1030 25800
rect 1086 25744 1348 25800
rect 1025 25742 1348 25744
rect 1025 25739 1091 25742
rect 1342 25740 1348 25742
rect 1412 25740 1418 25804
rect 1894 25740 1900 25804
rect 1964 25802 1970 25804
rect 2998 25802 3004 25804
rect 1964 25742 3004 25802
rect 1964 25740 1970 25742
rect 2998 25740 3004 25742
rect 3068 25740 3074 25804
rect 3182 25740 3188 25804
rect 3252 25802 3258 25804
rect 3601 25802 3667 25805
rect 3252 25800 3667 25802
rect 3252 25744 3606 25800
rect 3662 25744 3667 25800
rect 3252 25742 3667 25744
rect 3742 25802 3802 25875
rect 9676 25805 9736 26286
rect 10041 26283 10107 26286
rect 10058 26144 10374 26145
rect 10058 26080 10064 26144
rect 10128 26080 10144 26144
rect 10208 26080 10224 26144
rect 10288 26080 10304 26144
rect 10368 26080 10374 26144
rect 10058 26079 10374 26080
rect 5901 25802 5967 25805
rect 3742 25800 5967 25802
rect 3742 25744 5906 25800
rect 5962 25744 5967 25800
rect 3742 25742 5967 25744
rect 3252 25740 3258 25742
rect 3601 25739 3667 25742
rect 5901 25739 5967 25742
rect 6310 25740 6316 25804
rect 6380 25802 6386 25804
rect 8477 25802 8543 25805
rect 6380 25800 8543 25802
rect 6380 25744 8482 25800
rect 8538 25744 8543 25800
rect 6380 25742 8543 25744
rect 6380 25740 6386 25742
rect 8477 25739 8543 25742
rect 9673 25800 9739 25805
rect 9673 25744 9678 25800
rect 9734 25744 9739 25800
rect 9673 25739 9739 25744
rect 381 25666 447 25669
rect 3182 25666 3188 25668
rect 381 25664 3188 25666
rect 381 25608 386 25664
rect 442 25608 3188 25664
rect 381 25606 3188 25608
rect 381 25603 447 25606
rect 3182 25604 3188 25606
rect 3252 25604 3258 25668
rect 3693 25666 3759 25669
rect 4153 25666 4219 25669
rect 5758 25666 5764 25668
rect 3693 25664 4219 25666
rect 3693 25608 3698 25664
rect 3754 25608 4158 25664
rect 4214 25608 4219 25664
rect 3693 25606 4219 25608
rect 3693 25603 3759 25606
rect 4153 25603 4219 25606
rect 4708 25606 5764 25666
rect 4318 25600 4634 25601
rect 4318 25536 4324 25600
rect 4388 25536 4404 25600
rect 4468 25536 4484 25600
rect 4548 25536 4564 25600
rect 4628 25536 4634 25600
rect 4318 25535 4634 25536
rect 4708 25533 4768 25606
rect 5758 25604 5764 25606
rect 5828 25604 5834 25668
rect 6637 25666 6703 25669
rect 8753 25666 8819 25669
rect 6637 25664 8819 25666
rect 6637 25608 6642 25664
rect 6698 25608 8758 25664
rect 8814 25608 8819 25664
rect 6637 25606 8819 25608
rect 6637 25603 6703 25606
rect 8753 25603 8819 25606
rect 10718 25600 11034 25601
rect 10718 25536 10724 25600
rect 10788 25536 10804 25600
rect 10868 25536 10884 25600
rect 10948 25536 10964 25600
rect 11028 25536 11034 25600
rect 10718 25535 11034 25536
rect 2589 25530 2655 25533
rect 2589 25528 4170 25530
rect 2589 25472 2594 25528
rect 2650 25472 4170 25528
rect 2589 25470 4170 25472
rect 2589 25467 2655 25470
rect 2078 25332 2084 25396
rect 2148 25394 2154 25396
rect 2773 25394 2839 25397
rect 2148 25392 2839 25394
rect 2148 25336 2778 25392
rect 2834 25336 2839 25392
rect 2148 25334 2839 25336
rect 2148 25332 2154 25334
rect 2773 25331 2839 25334
rect 2998 25332 3004 25396
rect 3068 25394 3074 25396
rect 3785 25394 3851 25397
rect 3068 25392 3851 25394
rect 3068 25336 3790 25392
rect 3846 25336 3851 25392
rect 3068 25334 3851 25336
rect 4110 25394 4170 25470
rect 4705 25528 4771 25533
rect 4705 25472 4710 25528
rect 4766 25472 4771 25528
rect 4705 25467 4771 25472
rect 4981 25530 5047 25533
rect 6729 25530 6795 25533
rect 4981 25528 6795 25530
rect 4981 25472 4986 25528
rect 5042 25472 6734 25528
rect 6790 25472 6795 25528
rect 4981 25470 6795 25472
rect 4981 25467 5047 25470
rect 6729 25467 6795 25470
rect 7005 25530 7071 25533
rect 8569 25530 8635 25533
rect 7005 25528 8635 25530
rect 7005 25472 7010 25528
rect 7066 25472 8574 25528
rect 8630 25472 8635 25528
rect 7005 25470 8635 25472
rect 7005 25467 7071 25470
rect 8569 25467 8635 25470
rect 6913 25394 6979 25397
rect 8569 25394 8635 25397
rect 9254 25394 9260 25396
rect 4110 25392 6979 25394
rect 4110 25336 6918 25392
rect 6974 25336 6979 25392
rect 4110 25334 6979 25336
rect 3068 25332 3074 25334
rect 3785 25331 3851 25334
rect 6913 25331 6979 25334
rect 7054 25392 9260 25394
rect 7054 25336 8574 25392
rect 8630 25336 9260 25392
rect 7054 25334 9260 25336
rect 3366 25196 3372 25260
rect 3436 25258 3442 25260
rect 3693 25258 3759 25261
rect 3436 25256 3759 25258
rect 3436 25200 3698 25256
rect 3754 25200 3759 25256
rect 3436 25198 3759 25200
rect 3436 25196 3442 25198
rect 3693 25195 3759 25198
rect 3877 25258 3943 25261
rect 4889 25258 4955 25261
rect 5206 25258 5212 25260
rect 3877 25256 4768 25258
rect 3877 25200 3882 25256
rect 3938 25200 4768 25256
rect 3877 25198 4768 25200
rect 3877 25195 3943 25198
rect 2262 25060 2268 25124
rect 2332 25122 2338 25124
rect 2405 25122 2471 25125
rect 2332 25120 2471 25122
rect 2332 25064 2410 25120
rect 2466 25064 2471 25120
rect 2332 25062 2471 25064
rect 4708 25122 4768 25198
rect 4889 25256 5212 25258
rect 4889 25200 4894 25256
rect 4950 25200 5212 25256
rect 4889 25198 5212 25200
rect 4889 25195 4955 25198
rect 5206 25196 5212 25198
rect 5276 25258 5282 25260
rect 5533 25258 5599 25261
rect 5276 25256 5599 25258
rect 5276 25200 5538 25256
rect 5594 25200 5599 25256
rect 5276 25198 5599 25200
rect 5276 25196 5282 25198
rect 5533 25195 5599 25198
rect 5901 25258 5967 25261
rect 7054 25258 7114 25334
rect 8569 25331 8635 25334
rect 9254 25332 9260 25334
rect 9324 25332 9330 25396
rect 5901 25256 7114 25258
rect 5901 25200 5906 25256
rect 5962 25200 7114 25256
rect 5901 25198 7114 25200
rect 5901 25195 5967 25198
rect 8518 25196 8524 25260
rect 8588 25258 8594 25260
rect 10685 25258 10751 25261
rect 8588 25256 10751 25258
rect 8588 25200 10690 25256
rect 10746 25200 10751 25256
rect 8588 25198 10751 25200
rect 8588 25196 8594 25198
rect 10685 25195 10751 25198
rect 4981 25122 5047 25125
rect 5349 25122 5415 25125
rect 6453 25124 6519 25125
rect 6453 25122 6500 25124
rect 4708 25120 5047 25122
rect 4708 25064 4986 25120
rect 5042 25064 5047 25120
rect 4708 25062 5047 25064
rect 2332 25060 2338 25062
rect 2405 25059 2471 25062
rect 4981 25059 5047 25062
rect 5168 25120 5415 25122
rect 5168 25064 5354 25120
rect 5410 25064 5415 25120
rect 5168 25062 5415 25064
rect 6372 25120 6500 25122
rect 6564 25122 6570 25124
rect 7373 25122 7439 25125
rect 6564 25120 7439 25122
rect 6372 25064 6458 25120
rect 6564 25064 7378 25120
rect 7434 25064 7439 25120
rect 6372 25062 6500 25064
rect 3658 25056 3974 25057
rect 3658 24992 3664 25056
rect 3728 24992 3744 25056
rect 3808 24992 3824 25056
rect 3888 24992 3904 25056
rect 3968 24992 3974 25056
rect 3658 24991 3974 24992
rect 2313 24988 2379 24989
rect 2262 24986 2268 24988
rect 2222 24926 2268 24986
rect 2332 24984 2379 24988
rect 2374 24928 2379 24984
rect 2262 24924 2268 24926
rect 2332 24924 2379 24928
rect 2313 24923 2379 24924
rect 4889 24986 4955 24989
rect 5168 24986 5228 25062
rect 5349 25059 5415 25062
rect 6453 25060 6500 25062
rect 6564 25062 7439 25064
rect 6564 25060 6570 25062
rect 6453 25059 6519 25060
rect 7373 25059 7439 25062
rect 7741 25122 7807 25125
rect 8518 25122 8524 25124
rect 7741 25120 8524 25122
rect 7741 25064 7746 25120
rect 7802 25064 8524 25120
rect 7741 25062 8524 25064
rect 7741 25059 7807 25062
rect 8518 25060 8524 25062
rect 8588 25060 8594 25124
rect 8661 25122 8727 25125
rect 8886 25122 8892 25124
rect 8661 25120 8892 25122
rect 8661 25064 8666 25120
rect 8722 25064 8892 25120
rect 8661 25062 8892 25064
rect 8661 25059 8727 25062
rect 8886 25060 8892 25062
rect 8956 25060 8962 25124
rect 10058 25056 10374 25057
rect 10058 24992 10064 25056
rect 10128 24992 10144 25056
rect 10208 24992 10224 25056
rect 10288 24992 10304 25056
rect 10368 24992 10374 25056
rect 10058 24991 10374 24992
rect 5717 24986 5783 24989
rect 4889 24984 5228 24986
rect 4889 24928 4894 24984
rect 4950 24928 5228 24984
rect 4889 24926 5228 24928
rect 5352 24984 5783 24986
rect 5352 24928 5722 24984
rect 5778 24928 5783 24984
rect 5352 24926 5783 24928
rect 4889 24923 4955 24926
rect 5352 24870 5412 24926
rect 5717 24923 5783 24926
rect 7465 24986 7531 24989
rect 7966 24986 7972 24988
rect 7465 24984 7972 24986
rect 7465 24928 7470 24984
rect 7526 24928 7972 24984
rect 7465 24926 7972 24928
rect 7465 24923 7531 24926
rect 7966 24924 7972 24926
rect 8036 24924 8042 24988
rect 8886 24924 8892 24988
rect 8956 24986 8962 24988
rect 9121 24986 9187 24989
rect 8956 24984 9187 24986
rect 8956 24928 9126 24984
rect 9182 24928 9187 24984
rect 8956 24926 9187 24928
rect 8956 24924 8962 24926
rect 9121 24923 9187 24926
rect 2405 24850 2471 24853
rect 5260 24850 5412 24870
rect 2405 24848 5412 24850
rect 2405 24792 2410 24848
rect 2466 24810 5412 24848
rect 5717 24850 5783 24853
rect 5901 24850 5967 24853
rect 5717 24848 5967 24850
rect 2466 24792 5320 24810
rect 2405 24790 5320 24792
rect 5717 24792 5722 24848
rect 5778 24792 5906 24848
rect 5962 24792 5967 24848
rect 5717 24790 5967 24792
rect 2405 24787 2471 24790
rect 5717 24787 5783 24790
rect 5901 24787 5967 24790
rect 6085 24850 6151 24853
rect 7465 24850 7531 24853
rect 8017 24850 8083 24853
rect 6085 24848 7068 24850
rect 6085 24792 6090 24848
rect 6146 24792 7068 24848
rect 6085 24790 7068 24792
rect 6085 24787 6151 24790
rect 1393 24714 1459 24717
rect 5625 24716 5691 24717
rect 5574 24714 5580 24716
rect 1393 24712 5320 24714
rect 1393 24656 1398 24712
rect 1454 24656 5320 24712
rect 1393 24654 5320 24656
rect 5534 24654 5580 24714
rect 5644 24712 5691 24716
rect 6862 24714 6868 24716
rect 5686 24656 5691 24712
rect 1393 24651 1459 24654
rect 5260 24581 5320 24654
rect 5574 24652 5580 24654
rect 5644 24652 5691 24656
rect 5625 24651 5691 24652
rect 5812 24654 6868 24714
rect 1526 24516 1532 24580
rect 1596 24578 1602 24580
rect 2037 24578 2103 24581
rect 1596 24576 2103 24578
rect 1596 24520 2042 24576
rect 2098 24520 2103 24576
rect 1596 24518 2103 24520
rect 1596 24516 1602 24518
rect 2037 24515 2103 24518
rect 4700 24516 4706 24580
rect 4770 24578 4776 24580
rect 4770 24518 5136 24578
rect 4770 24516 4776 24518
rect 4318 24512 4634 24513
rect 4318 24448 4324 24512
rect 4388 24448 4404 24512
rect 4468 24448 4484 24512
rect 4548 24448 4564 24512
rect 4628 24448 4634 24512
rect 4318 24447 4634 24448
rect 5076 24445 5136 24518
rect 5257 24576 5323 24581
rect 5257 24520 5262 24576
rect 5318 24520 5323 24576
rect 5257 24515 5323 24520
rect 5441 24578 5507 24581
rect 5812 24578 5872 24654
rect 6862 24652 6868 24654
rect 6932 24652 6938 24716
rect 7008 24714 7068 24790
rect 7465 24848 8083 24850
rect 7465 24792 7470 24848
rect 7526 24792 8022 24848
rect 8078 24792 8083 24848
rect 7465 24790 8083 24792
rect 7465 24787 7531 24790
rect 8017 24787 8083 24790
rect 8569 24714 8635 24717
rect 7008 24712 8635 24714
rect 7008 24656 8574 24712
rect 8630 24656 8635 24712
rect 7008 24654 8635 24656
rect 8569 24651 8635 24654
rect 8702 24652 8708 24716
rect 8772 24714 8778 24716
rect 10041 24714 10107 24717
rect 8772 24712 10107 24714
rect 8772 24656 10046 24712
rect 10102 24656 10107 24712
rect 8772 24654 10107 24656
rect 8772 24652 8778 24654
rect 10041 24651 10107 24654
rect 5441 24576 5872 24578
rect 5441 24520 5446 24576
rect 5502 24520 5872 24576
rect 5441 24518 5872 24520
rect 5441 24515 5507 24518
rect 6126 24516 6132 24580
rect 6196 24578 6202 24580
rect 6453 24578 6519 24581
rect 6196 24576 6519 24578
rect 6196 24520 6458 24576
rect 6514 24520 6519 24576
rect 6196 24518 6519 24520
rect 6196 24516 6202 24518
rect 6453 24515 6519 24518
rect 10718 24512 11034 24513
rect 10718 24448 10724 24512
rect 10788 24448 10804 24512
rect 10868 24448 10884 24512
rect 10948 24448 10964 24512
rect 11028 24448 11034 24512
rect 10718 24447 11034 24448
rect 1761 24442 1827 24445
rect 2037 24442 2103 24445
rect 1761 24440 2103 24442
rect 1761 24384 1766 24440
rect 1822 24384 2042 24440
rect 2098 24384 2103 24440
rect 1761 24382 2103 24384
rect 1761 24379 1827 24382
rect 2037 24379 2103 24382
rect 5073 24442 5139 24445
rect 5717 24444 5783 24445
rect 5206 24442 5212 24444
rect 5073 24440 5212 24442
rect 5073 24384 5078 24440
rect 5134 24384 5212 24440
rect 5073 24382 5212 24384
rect 5073 24379 5139 24382
rect 5206 24380 5212 24382
rect 5276 24380 5282 24444
rect 5717 24442 5764 24444
rect 5672 24440 5764 24442
rect 5672 24384 5722 24440
rect 5672 24382 5764 24384
rect 5717 24380 5764 24382
rect 5828 24380 5834 24444
rect 6126 24380 6132 24444
rect 6196 24442 6202 24444
rect 6545 24442 6611 24445
rect 6196 24440 6611 24442
rect 6196 24384 6550 24440
rect 6606 24384 6611 24440
rect 6196 24382 6611 24384
rect 6196 24380 6202 24382
rect 5717 24379 5783 24380
rect 6545 24379 6611 24382
rect 6913 24442 6979 24445
rect 7046 24442 7052 24444
rect 6913 24440 7052 24442
rect 6913 24384 6918 24440
rect 6974 24384 7052 24440
rect 6913 24382 7052 24384
rect 6913 24379 6979 24382
rect 7046 24380 7052 24382
rect 7116 24380 7122 24444
rect 7373 24442 7439 24445
rect 9213 24442 9279 24445
rect 7373 24440 9279 24442
rect 7373 24384 7378 24440
rect 7434 24384 9218 24440
rect 9274 24384 9279 24440
rect 7373 24382 9279 24384
rect 7373 24379 7439 24382
rect 9213 24379 9279 24382
rect 0 24306 400 24336
rect 1025 24306 1091 24309
rect 0 24304 1091 24306
rect 0 24248 1030 24304
rect 1086 24248 1091 24304
rect 0 24246 1091 24248
rect 0 24216 400 24246
rect 1025 24243 1091 24246
rect 1894 24244 1900 24308
rect 1964 24306 1970 24308
rect 2589 24306 2655 24309
rect 3693 24306 3759 24309
rect 1964 24304 3759 24306
rect 1964 24248 2594 24304
rect 2650 24248 3698 24304
rect 3754 24248 3759 24304
rect 1964 24246 3759 24248
rect 1964 24244 1970 24246
rect 2589 24243 2655 24246
rect 3693 24243 3759 24246
rect 3877 24306 3943 24309
rect 7465 24306 7531 24309
rect 8569 24306 8635 24309
rect 3877 24304 8635 24306
rect 3877 24248 3882 24304
rect 3938 24248 7470 24304
rect 7526 24248 8574 24304
rect 8630 24248 8635 24304
rect 3877 24246 8635 24248
rect 3877 24243 3943 24246
rect 7465 24243 7531 24246
rect 8569 24243 8635 24246
rect 8845 24306 8911 24309
rect 10777 24306 10843 24309
rect 8845 24304 10843 24306
rect 8845 24248 8850 24304
rect 8906 24248 10782 24304
rect 10838 24248 10843 24304
rect 8845 24246 10843 24248
rect 8845 24243 8911 24246
rect 10777 24243 10843 24246
rect 10961 24306 11027 24309
rect 11094 24306 11100 24308
rect 10961 24304 11100 24306
rect 10961 24248 10966 24304
rect 11022 24248 11100 24304
rect 10961 24246 11100 24248
rect 10961 24243 11027 24246
rect 11094 24244 11100 24246
rect 11164 24244 11170 24308
rect 1342 24108 1348 24172
rect 1412 24170 1418 24172
rect 1894 24170 1900 24172
rect 1412 24110 1900 24170
rect 1412 24108 1418 24110
rect 1894 24108 1900 24110
rect 1964 24108 1970 24172
rect 3049 24170 3115 24173
rect 9581 24170 9647 24173
rect 3049 24168 9647 24170
rect 3049 24112 3054 24168
rect 3110 24112 9586 24168
rect 9642 24112 9647 24168
rect 3049 24110 9647 24112
rect 3049 24107 3115 24110
rect 9581 24107 9647 24110
rect 10317 24170 10383 24173
rect 10542 24170 10548 24172
rect 10317 24168 10548 24170
rect 10317 24112 10322 24168
rect 10378 24112 10548 24168
rect 10317 24110 10548 24112
rect 10317 24107 10383 24110
rect 10542 24108 10548 24110
rect 10612 24170 10618 24172
rect 11094 24170 11100 24172
rect 10612 24110 11100 24170
rect 10612 24108 10618 24110
rect 11094 24108 11100 24110
rect 11164 24108 11170 24172
rect 0 24034 400 24064
rect 1301 24034 1367 24037
rect 0 24032 1367 24034
rect 0 23976 1306 24032
rect 1362 23976 1367 24032
rect 0 23974 1367 23976
rect 0 23944 400 23974
rect 1301 23971 1367 23974
rect 4797 24034 4863 24037
rect 6913 24034 6979 24037
rect 7230 24034 7236 24036
rect 4797 24032 7236 24034
rect 4797 23976 4802 24032
rect 4858 23976 6918 24032
rect 6974 23976 7236 24032
rect 4797 23974 7236 23976
rect 4797 23971 4863 23974
rect 6913 23971 6979 23974
rect 7230 23972 7236 23974
rect 7300 23972 7306 24036
rect 7373 24034 7439 24037
rect 8661 24034 8727 24037
rect 8937 24034 9003 24037
rect 9213 24034 9279 24037
rect 7373 24032 8448 24034
rect 7373 23976 7378 24032
rect 7434 23976 8448 24032
rect 7373 23974 8448 23976
rect 7373 23971 7439 23974
rect 3658 23968 3974 23969
rect 3658 23904 3664 23968
rect 3728 23904 3744 23968
rect 3808 23904 3824 23968
rect 3888 23904 3904 23968
rect 3968 23904 3974 23968
rect 3658 23903 3974 23904
rect 8388 23901 8448 23974
rect 8661 24032 9279 24034
rect 8661 23976 8666 24032
rect 8722 23976 8942 24032
rect 8998 23976 9218 24032
rect 9274 23976 9279 24032
rect 8661 23974 9279 23976
rect 8661 23971 8727 23974
rect 8937 23971 9003 23974
rect 9213 23971 9279 23974
rect 9397 24034 9463 24037
rect 9765 24034 9831 24037
rect 9397 24032 9831 24034
rect 9397 23976 9402 24032
rect 9458 23976 9770 24032
rect 9826 23976 9831 24032
rect 9397 23974 9831 23976
rect 9397 23971 9463 23974
rect 9765 23971 9831 23974
rect 10542 23972 10548 24036
rect 10612 24034 10618 24036
rect 10777 24034 10843 24037
rect 10612 24032 10843 24034
rect 10612 23976 10782 24032
rect 10838 23976 10843 24032
rect 10612 23974 10843 23976
rect 10612 23972 10618 23974
rect 10777 23971 10843 23974
rect 10058 23968 10374 23969
rect 10058 23904 10064 23968
rect 10128 23904 10144 23968
rect 10208 23904 10224 23968
rect 10288 23904 10304 23968
rect 10368 23904 10374 23968
rect 10058 23903 10374 23904
rect 933 23898 999 23901
rect 5257 23898 5323 23901
rect 6177 23898 6243 23901
rect 7373 23898 7439 23901
rect 933 23896 3572 23898
rect 933 23840 938 23896
rect 994 23840 3572 23896
rect 933 23838 3572 23840
rect 933 23835 999 23838
rect 0 23762 400 23792
rect 2773 23762 2839 23765
rect 0 23760 2839 23762
rect 0 23704 2778 23760
rect 2834 23704 2839 23760
rect 0 23702 2839 23704
rect 3512 23762 3572 23838
rect 4846 23896 7439 23898
rect 4846 23840 5262 23896
rect 5318 23840 6182 23896
rect 6238 23840 7378 23896
rect 7434 23840 7439 23896
rect 4846 23838 7439 23840
rect 4846 23762 4906 23838
rect 5257 23835 5323 23838
rect 6177 23835 6243 23838
rect 7373 23835 7439 23838
rect 7741 23898 7807 23901
rect 7925 23898 7991 23901
rect 7741 23896 7991 23898
rect 7741 23840 7746 23896
rect 7802 23840 7930 23896
rect 7986 23840 7991 23896
rect 7741 23838 7991 23840
rect 7741 23835 7807 23838
rect 7925 23835 7991 23838
rect 8385 23896 8451 23901
rect 9213 23900 9279 23901
rect 9213 23898 9260 23900
rect 8385 23840 8390 23896
rect 8446 23840 8451 23896
rect 8385 23835 8451 23840
rect 9168 23896 9260 23898
rect 9168 23840 9218 23896
rect 9168 23838 9260 23840
rect 9213 23836 9260 23838
rect 9324 23836 9330 23900
rect 9213 23835 9279 23836
rect 6862 23762 6868 23764
rect 3512 23702 4906 23762
rect 4984 23702 6868 23762
rect 0 23672 400 23702
rect 2773 23699 2839 23702
rect 1158 23564 1164 23628
rect 1228 23626 1234 23628
rect 2497 23626 2563 23629
rect 3601 23626 3667 23629
rect 4984 23626 5044 23702
rect 6862 23700 6868 23702
rect 6932 23700 6938 23764
rect 7046 23700 7052 23764
rect 7116 23762 7122 23764
rect 9029 23762 9095 23765
rect 9438 23762 9444 23764
rect 7116 23702 8908 23762
rect 7116 23700 7122 23702
rect 1228 23624 3667 23626
rect 1228 23568 2502 23624
rect 2558 23568 3606 23624
rect 3662 23568 3667 23624
rect 1228 23566 3667 23568
rect 1228 23564 1234 23566
rect 2497 23563 2563 23566
rect 3601 23563 3667 23566
rect 3880 23566 5044 23626
rect 5625 23626 5691 23629
rect 5625 23624 7114 23626
rect 5625 23568 5630 23624
rect 5686 23568 7114 23624
rect 5625 23566 7114 23568
rect 0 23493 400 23520
rect 0 23488 447 23493
rect 1393 23492 1459 23493
rect 1342 23490 1348 23492
rect 0 23432 386 23488
rect 442 23432 447 23488
rect 0 23427 447 23432
rect 1302 23430 1348 23490
rect 1412 23488 1459 23492
rect 1454 23432 1459 23488
rect 1342 23428 1348 23430
rect 1412 23428 1459 23432
rect 1710 23428 1716 23492
rect 1780 23490 1786 23492
rect 3049 23490 3115 23493
rect 1780 23488 3115 23490
rect 1780 23432 3054 23488
rect 3110 23432 3115 23488
rect 1780 23430 3115 23432
rect 1780 23428 1786 23430
rect 1393 23427 1459 23428
rect 3049 23427 3115 23430
rect 0 23400 400 23427
rect 1710 23292 1716 23356
rect 1780 23354 1786 23356
rect 2078 23354 2084 23356
rect 1780 23294 2084 23354
rect 1780 23292 1786 23294
rect 2078 23292 2084 23294
rect 2148 23292 2154 23356
rect 0 23218 400 23248
rect 841 23218 907 23221
rect 0 23216 907 23218
rect 0 23160 846 23216
rect 902 23160 907 23216
rect 0 23158 907 23160
rect 0 23128 400 23158
rect 841 23155 907 23158
rect 2221 23218 2287 23221
rect 2446 23218 2452 23220
rect 2221 23216 2452 23218
rect 2221 23160 2226 23216
rect 2282 23160 2452 23216
rect 2221 23158 2452 23160
rect 2221 23155 2287 23158
rect 2446 23156 2452 23158
rect 2516 23156 2522 23220
rect 1209 23084 1275 23085
rect 1158 23082 1164 23084
rect 1118 23022 1164 23082
rect 1228 23080 1275 23084
rect 3880 23082 3940 23566
rect 5625 23563 5691 23566
rect 5717 23488 5783 23493
rect 5717 23432 5722 23488
rect 5778 23432 5783 23488
rect 5717 23427 5783 23432
rect 7054 23490 7114 23566
rect 7414 23564 7420 23628
rect 7484 23626 7490 23628
rect 7833 23626 7899 23629
rect 8385 23626 8451 23629
rect 8661 23628 8727 23629
rect 8661 23626 8708 23628
rect 7484 23624 8451 23626
rect 7484 23568 7838 23624
rect 7894 23568 8390 23624
rect 8446 23568 8451 23624
rect 7484 23566 8451 23568
rect 8616 23624 8708 23626
rect 8616 23568 8666 23624
rect 8616 23566 8708 23568
rect 7484 23564 7490 23566
rect 7833 23563 7899 23566
rect 8385 23563 8451 23566
rect 8661 23564 8708 23566
rect 8772 23564 8778 23628
rect 8848 23626 8908 23702
rect 9029 23760 9444 23762
rect 9029 23704 9034 23760
rect 9090 23704 9444 23760
rect 9029 23702 9444 23704
rect 9029 23699 9095 23702
rect 9438 23700 9444 23702
rect 9508 23762 9514 23764
rect 10317 23762 10383 23765
rect 9508 23760 10383 23762
rect 9508 23704 10322 23760
rect 10378 23704 10383 23760
rect 9508 23702 10383 23704
rect 9508 23700 9514 23702
rect 10317 23699 10383 23702
rect 9581 23626 9647 23629
rect 8848 23624 9647 23626
rect 8848 23568 9586 23624
rect 9642 23568 9647 23624
rect 8848 23566 9647 23568
rect 8661 23563 8727 23564
rect 9581 23563 9647 23566
rect 9438 23490 9444 23492
rect 7054 23430 9444 23490
rect 9438 23428 9444 23430
rect 9508 23428 9514 23492
rect 9581 23490 9647 23493
rect 10317 23490 10383 23493
rect 9581 23488 10383 23490
rect 9581 23432 9586 23488
rect 9642 23432 10322 23488
rect 10378 23432 10383 23488
rect 9581 23430 10383 23432
rect 9581 23427 9647 23430
rect 10317 23427 10383 23430
rect 4318 23424 4634 23425
rect 4318 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4634 23424
rect 4318 23359 4634 23360
rect 5720 23354 5780 23427
rect 10718 23424 11034 23425
rect 10718 23360 10724 23424
rect 10788 23360 10804 23424
rect 10868 23360 10884 23424
rect 10948 23360 10964 23424
rect 11028 23360 11034 23424
rect 10718 23359 11034 23360
rect 6085 23354 6151 23357
rect 5720 23352 6151 23354
rect 5720 23296 6090 23352
rect 6146 23296 6151 23352
rect 5720 23294 6151 23296
rect 6085 23291 6151 23294
rect 6269 23354 6335 23357
rect 8201 23354 8267 23357
rect 8886 23354 8892 23356
rect 6269 23352 8892 23354
rect 6269 23296 6274 23352
rect 6330 23296 8206 23352
rect 8262 23296 8892 23352
rect 6269 23294 8892 23296
rect 6269 23291 6335 23294
rect 8201 23291 8267 23294
rect 8886 23292 8892 23294
rect 8956 23292 8962 23356
rect 4429 23218 4495 23221
rect 6862 23218 6868 23220
rect 4429 23216 6056 23218
rect 4429 23160 4434 23216
rect 4490 23184 6056 23216
rect 6180 23184 6868 23218
rect 4490 23160 6868 23184
rect 4429 23158 6868 23160
rect 4429 23155 4495 23158
rect 5996 23124 6240 23158
rect 6862 23156 6868 23158
rect 6932 23156 6938 23220
rect 7230 23156 7236 23220
rect 7300 23218 7306 23220
rect 8201 23218 8267 23221
rect 7300 23216 8267 23218
rect 7300 23160 8206 23216
rect 8262 23160 8267 23216
rect 7300 23158 8267 23160
rect 7300 23156 7306 23158
rect 8201 23155 8267 23158
rect 8518 23156 8524 23220
rect 8588 23218 8594 23220
rect 9029 23218 9095 23221
rect 8588 23216 9095 23218
rect 8588 23160 9034 23216
rect 9090 23160 9095 23216
rect 8588 23158 9095 23160
rect 8588 23156 8594 23158
rect 9029 23155 9095 23158
rect 9397 23218 9463 23221
rect 10133 23218 10199 23221
rect 9397 23216 10199 23218
rect 9397 23160 9402 23216
rect 9458 23160 10138 23216
rect 10194 23160 10199 23216
rect 9397 23158 10199 23160
rect 9397 23155 9463 23158
rect 10133 23155 10199 23158
rect 10685 23218 10751 23221
rect 11094 23218 11100 23220
rect 10685 23216 11100 23218
rect 10685 23160 10690 23216
rect 10746 23160 11100 23216
rect 10685 23158 11100 23160
rect 10685 23155 10751 23158
rect 11094 23156 11100 23158
rect 11164 23156 11170 23220
rect 1270 23024 1275 23080
rect 1158 23020 1164 23022
rect 1228 23020 1275 23024
rect 1209 23019 1275 23020
rect 3512 23022 3940 23082
rect 7281 23082 7347 23085
rect 9949 23082 10015 23085
rect 7281 23080 10015 23082
rect 7281 23024 7286 23080
rect 7342 23024 9954 23080
rect 10010 23024 10015 23080
rect 7281 23022 10015 23024
rect 0 22946 400 22976
rect 933 22946 999 22949
rect 0 22944 999 22946
rect 0 22888 938 22944
rect 994 22888 999 22944
rect 0 22886 999 22888
rect 0 22856 400 22886
rect 933 22883 999 22886
rect 0 22674 400 22704
rect 1669 22674 1735 22677
rect 0 22672 1735 22674
rect 0 22616 1674 22672
rect 1730 22616 1735 22672
rect 0 22614 1735 22616
rect 3512 22674 3572 23022
rect 7281 23019 7347 23022
rect 9949 23019 10015 23022
rect 4102 22884 4108 22948
rect 4172 22946 4178 22948
rect 5349 22946 5415 22949
rect 4172 22944 5415 22946
rect 4172 22888 5354 22944
rect 5410 22888 5415 22944
rect 4172 22886 5415 22888
rect 4172 22884 4178 22886
rect 5349 22883 5415 22886
rect 5901 22946 5967 22949
rect 6821 22946 6887 22949
rect 5901 22944 6887 22946
rect 5901 22888 5906 22944
rect 5962 22888 6826 22944
rect 6882 22888 6887 22944
rect 5901 22886 6887 22888
rect 5901 22883 5967 22886
rect 6821 22883 6887 22886
rect 7414 22884 7420 22948
rect 7484 22946 7490 22948
rect 7782 22946 7788 22948
rect 7484 22886 7788 22946
rect 7484 22884 7490 22886
rect 7782 22884 7788 22886
rect 7852 22884 7858 22948
rect 8150 22884 8156 22948
rect 8220 22946 8226 22948
rect 8518 22946 8524 22948
rect 8220 22886 8524 22946
rect 8220 22884 8226 22886
rect 8518 22884 8524 22886
rect 8588 22884 8594 22948
rect 9305 22946 9371 22949
rect 9438 22946 9444 22948
rect 9305 22944 9444 22946
rect 9305 22888 9310 22944
rect 9366 22888 9444 22944
rect 9305 22886 9444 22888
rect 9305 22883 9371 22886
rect 9438 22884 9444 22886
rect 9508 22884 9514 22948
rect 3658 22880 3974 22881
rect 3658 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3974 22880
rect 3658 22815 3974 22816
rect 10058 22880 10374 22881
rect 10058 22816 10064 22880
rect 10128 22816 10144 22880
rect 10208 22816 10224 22880
rect 10288 22816 10304 22880
rect 10368 22816 10374 22880
rect 10058 22815 10374 22816
rect 4102 22748 4108 22812
rect 4172 22810 4178 22812
rect 4245 22810 4311 22813
rect 4172 22808 4311 22810
rect 4172 22752 4250 22808
rect 4306 22752 4311 22808
rect 4172 22750 4311 22752
rect 4172 22748 4178 22750
rect 4245 22747 4311 22750
rect 5073 22810 5139 22813
rect 9254 22810 9260 22812
rect 5073 22808 9260 22810
rect 5073 22752 5078 22808
rect 5134 22752 9260 22808
rect 5073 22750 9260 22752
rect 5073 22747 5139 22750
rect 9254 22748 9260 22750
rect 9324 22748 9330 22812
rect 3785 22674 3851 22677
rect 3512 22672 3851 22674
rect 3512 22616 3790 22672
rect 3846 22616 3851 22672
rect 3512 22614 3851 22616
rect 0 22584 400 22614
rect 1669 22611 1735 22614
rect 3785 22611 3851 22614
rect 5441 22672 5507 22677
rect 5441 22616 5446 22672
rect 5502 22616 5507 22672
rect 5441 22611 5507 22616
rect 5942 22612 5948 22676
rect 6012 22674 6018 22676
rect 6177 22674 6243 22677
rect 6012 22672 6243 22674
rect 6012 22616 6182 22672
rect 6238 22616 6243 22672
rect 6012 22614 6243 22616
rect 6012 22612 6018 22614
rect 6177 22611 6243 22614
rect 6494 22612 6500 22676
rect 6564 22674 6570 22676
rect 6729 22674 6795 22677
rect 6564 22672 6795 22674
rect 6564 22616 6734 22672
rect 6790 22616 6795 22672
rect 6564 22614 6795 22616
rect 6564 22612 6570 22614
rect 6729 22611 6795 22614
rect 7097 22674 7163 22677
rect 8702 22674 8708 22676
rect 7097 22672 8708 22674
rect 7097 22616 7102 22672
rect 7158 22616 8708 22672
rect 7097 22614 8708 22616
rect 7097 22611 7163 22614
rect 8702 22612 8708 22614
rect 8772 22612 8778 22676
rect 1301 22538 1367 22541
rect 1894 22538 1900 22540
rect 1301 22536 1900 22538
rect 1301 22480 1306 22536
rect 1362 22480 1900 22536
rect 1301 22478 1900 22480
rect 1301 22475 1367 22478
rect 1894 22476 1900 22478
rect 1964 22476 1970 22540
rect 2446 22476 2452 22540
rect 2516 22538 2522 22540
rect 5444 22538 5504 22611
rect 7230 22538 7236 22540
rect 2516 22478 4768 22538
rect 5444 22478 7236 22538
rect 2516 22476 2522 22478
rect 422 22340 428 22404
rect 492 22402 498 22404
rect 933 22402 999 22405
rect 492 22400 999 22402
rect 492 22344 938 22400
rect 994 22344 999 22400
rect 492 22342 999 22344
rect 492 22340 498 22342
rect 933 22339 999 22342
rect 2221 22400 2287 22405
rect 2497 22404 2563 22405
rect 2221 22344 2226 22400
rect 2282 22344 2287 22400
rect 2221 22339 2287 22344
rect 2446 22340 2452 22404
rect 2516 22402 2563 22404
rect 2516 22400 2608 22402
rect 2558 22344 2608 22400
rect 2516 22342 2608 22344
rect 2516 22340 2563 22342
rect 2814 22340 2820 22404
rect 2884 22402 2890 22404
rect 3049 22402 3115 22405
rect 2884 22400 3115 22402
rect 2884 22344 3054 22400
rect 3110 22344 3115 22400
rect 2884 22342 3115 22344
rect 2884 22340 2890 22342
rect 2497 22339 2563 22340
rect 3049 22339 3115 22342
rect 3182 22340 3188 22404
rect 3252 22402 3258 22404
rect 3877 22402 3943 22405
rect 3252 22400 3943 22402
rect 3252 22344 3882 22400
rect 3938 22344 3943 22400
rect 3252 22342 3943 22344
rect 3252 22340 3258 22342
rect 3877 22339 3943 22342
rect 105 22266 171 22269
rect 790 22266 796 22268
rect 105 22264 796 22266
rect 105 22208 110 22264
rect 166 22208 796 22264
rect 105 22206 796 22208
rect 105 22203 171 22206
rect 790 22204 796 22206
rect 860 22204 866 22268
rect 2224 22266 2284 22339
rect 4318 22336 4634 22337
rect 4318 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4634 22336
rect 4318 22271 4634 22272
rect 4708 22269 4768 22478
rect 7230 22476 7236 22478
rect 7300 22538 7306 22540
rect 8569 22538 8635 22541
rect 7300 22536 8635 22538
rect 7300 22480 8574 22536
rect 8630 22480 8635 22536
rect 7300 22478 8635 22480
rect 7300 22476 7306 22478
rect 8569 22475 8635 22478
rect 5206 22340 5212 22404
rect 5276 22402 5282 22404
rect 6729 22402 6795 22405
rect 5276 22400 6795 22402
rect 5276 22344 6734 22400
rect 6790 22344 6795 22400
rect 5276 22342 6795 22344
rect 5276 22340 5282 22342
rect 6729 22339 6795 22342
rect 8150 22340 8156 22404
rect 8220 22402 8226 22404
rect 9121 22402 9187 22405
rect 8220 22400 9187 22402
rect 8220 22344 9126 22400
rect 9182 22344 9187 22400
rect 8220 22342 9187 22344
rect 8220 22340 8226 22342
rect 9121 22339 9187 22342
rect 10718 22336 11034 22337
rect 10718 22272 10724 22336
rect 10788 22272 10804 22336
rect 10868 22272 10884 22336
rect 10948 22272 10964 22336
rect 11028 22272 11034 22336
rect 10718 22271 11034 22272
rect 2497 22266 2563 22269
rect 2224 22264 2563 22266
rect 2224 22208 2502 22264
rect 2558 22208 2563 22264
rect 2224 22206 2563 22208
rect 2497 22203 2563 22206
rect 4705 22264 4771 22269
rect 4705 22208 4710 22264
rect 4766 22208 4771 22264
rect 4705 22203 4771 22208
rect 5257 22266 5323 22269
rect 6494 22266 6500 22268
rect 5257 22264 6500 22266
rect 5257 22208 5262 22264
rect 5318 22208 6500 22264
rect 5257 22206 6500 22208
rect 5257 22203 5323 22206
rect 6494 22204 6500 22206
rect 6564 22266 6570 22268
rect 6637 22266 6703 22269
rect 6564 22264 6703 22266
rect 6564 22208 6642 22264
rect 6698 22208 6703 22264
rect 6564 22206 6703 22208
rect 6564 22204 6570 22206
rect 6637 22203 6703 22206
rect 7097 22266 7163 22269
rect 7741 22266 7807 22269
rect 7097 22264 7807 22266
rect 7097 22208 7102 22264
rect 7158 22208 7746 22264
rect 7802 22208 7807 22264
rect 7097 22206 7807 22208
rect 7097 22203 7163 22206
rect 7741 22203 7807 22206
rect 7925 22266 7991 22269
rect 8753 22266 8819 22269
rect 7925 22264 8819 22266
rect 7925 22208 7930 22264
rect 7986 22208 8758 22264
rect 8814 22208 8819 22264
rect 7925 22206 8819 22208
rect 7925 22203 7991 22206
rect 8753 22203 8819 22206
rect 974 22068 980 22132
rect 1044 22130 1050 22132
rect 2814 22130 2820 22132
rect 1044 22070 2820 22130
rect 1044 22068 1050 22070
rect 2814 22068 2820 22070
rect 2884 22068 2890 22132
rect 4153 22128 4219 22133
rect 4153 22072 4158 22128
rect 4214 22072 4219 22128
rect 4153 22067 4219 22072
rect 4429 22130 4495 22133
rect 7782 22130 7788 22132
rect 4429 22128 7788 22130
rect 4429 22072 4434 22128
rect 4490 22072 7788 22128
rect 4429 22070 7788 22072
rect 4429 22067 4495 22070
rect 7782 22068 7788 22070
rect 7852 22068 7858 22132
rect 8845 22128 8911 22133
rect 8845 22072 8850 22128
rect 8906 22072 8911 22128
rect 8845 22067 8911 22072
rect 3049 21992 3115 21997
rect 3049 21936 3054 21992
rect 3110 21936 3115 21992
rect 3049 21931 3115 21936
rect 4156 21994 4216 22067
rect 5257 21994 5323 21997
rect 5993 21996 6059 21997
rect 5942 21994 5948 21996
rect 4156 21992 5323 21994
rect 4156 21936 5262 21992
rect 5318 21936 5323 21992
rect 4156 21934 5323 21936
rect 5902 21934 5948 21994
rect 6012 21992 6059 21996
rect 6054 21936 6059 21992
rect 5257 21931 5323 21934
rect 5942 21932 5948 21934
rect 6012 21932 6059 21936
rect 5993 21931 6059 21932
rect 6269 21996 6335 21997
rect 6269 21992 6316 21996
rect 6380 21994 6386 21996
rect 6545 21994 6611 21997
rect 6862 21994 6868 21996
rect 6269 21936 6274 21992
rect 6269 21932 6316 21936
rect 6380 21934 6426 21994
rect 6545 21992 6868 21994
rect 6545 21936 6550 21992
rect 6606 21936 6868 21992
rect 6545 21934 6868 21936
rect 6380 21932 6386 21934
rect 6269 21931 6335 21932
rect 6545 21931 6611 21934
rect 6862 21932 6868 21934
rect 6932 21994 6938 21996
rect 7557 21994 7623 21997
rect 8385 21996 8451 21997
rect 8334 21994 8340 21996
rect 6932 21992 7623 21994
rect 6932 21936 7562 21992
rect 7618 21936 7623 21992
rect 6932 21934 7623 21936
rect 8294 21934 8340 21994
rect 8404 21992 8451 21996
rect 8848 21994 8908 22067
rect 8446 21936 8451 21992
rect 6932 21932 6938 21934
rect 7557 21931 7623 21934
rect 8334 21932 8340 21934
rect 8404 21932 8451 21936
rect 8385 21931 8451 21932
rect 8756 21934 8908 21994
rect 9029 21994 9095 21997
rect 9673 21994 9739 21997
rect 9029 21992 9739 21994
rect 9029 21936 9034 21992
rect 9090 21936 9678 21992
rect 9734 21936 9739 21992
rect 9029 21934 9739 21936
rect 3052 21858 3112 21931
rect 3182 21858 3188 21860
rect 3052 21798 3188 21858
rect 3182 21796 3188 21798
rect 3252 21796 3258 21860
rect 4337 21858 4403 21861
rect 8756 21858 8816 21934
rect 9029 21931 9095 21934
rect 9673 21931 9739 21934
rect 4337 21856 8816 21858
rect 4337 21800 4342 21856
rect 4398 21800 8816 21856
rect 4337 21798 8816 21800
rect 4337 21795 4403 21798
rect 9438 21796 9444 21860
rect 9508 21858 9514 21860
rect 9581 21858 9647 21861
rect 10593 21860 10659 21861
rect 10542 21858 10548 21860
rect 9508 21856 9647 21858
rect 9508 21800 9586 21856
rect 9642 21800 9647 21856
rect 9508 21798 9647 21800
rect 10502 21798 10548 21858
rect 10612 21856 10659 21860
rect 10654 21800 10659 21856
rect 9508 21796 9514 21798
rect 9581 21795 9647 21798
rect 10542 21796 10548 21798
rect 10612 21796 10659 21800
rect 10593 21795 10659 21796
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 10058 21792 10374 21793
rect 10058 21728 10064 21792
rect 10128 21728 10144 21792
rect 10208 21728 10224 21792
rect 10288 21728 10304 21792
rect 10368 21728 10374 21792
rect 10058 21727 10374 21728
rect 2589 21722 2655 21725
rect 3049 21722 3115 21725
rect 2589 21720 3115 21722
rect 2589 21664 2594 21720
rect 2650 21664 3054 21720
rect 3110 21664 3115 21720
rect 2589 21662 3115 21664
rect 2589 21659 2655 21662
rect 3049 21659 3115 21662
rect 4337 21722 4403 21725
rect 5165 21722 5231 21725
rect 4337 21720 5231 21722
rect 4337 21664 4342 21720
rect 4398 21664 5170 21720
rect 5226 21664 5231 21720
rect 4337 21662 5231 21664
rect 4337 21659 4403 21662
rect 5165 21659 5231 21662
rect 5441 21722 5507 21725
rect 9397 21722 9463 21725
rect 5441 21720 9463 21722
rect 5441 21664 5446 21720
rect 5502 21664 9402 21720
rect 9458 21664 9463 21720
rect 5441 21662 9463 21664
rect 5441 21659 5507 21662
rect 9397 21659 9463 21662
rect 1393 21586 1459 21589
rect 4061 21586 4127 21589
rect 1393 21584 4127 21586
rect 1393 21528 1398 21584
rect 1454 21528 4066 21584
rect 4122 21528 4127 21584
rect 1393 21526 4127 21528
rect 1393 21523 1459 21526
rect 4061 21523 4127 21526
rect 4337 21586 4403 21589
rect 5574 21586 5580 21588
rect 4337 21584 5580 21586
rect 4337 21528 4342 21584
rect 4398 21528 5580 21584
rect 4337 21526 5580 21528
rect 4337 21523 4403 21526
rect 5574 21524 5580 21526
rect 5644 21586 5650 21588
rect 5993 21586 6059 21589
rect 5644 21584 6059 21586
rect 5644 21528 5998 21584
rect 6054 21528 6059 21584
rect 5644 21526 6059 21528
rect 5644 21524 5650 21526
rect 5993 21523 6059 21526
rect 8201 21586 8267 21589
rect 8334 21586 8340 21588
rect 8201 21584 8340 21586
rect 8201 21528 8206 21584
rect 8262 21528 8340 21584
rect 8201 21526 8340 21528
rect 8201 21523 8267 21526
rect 8334 21524 8340 21526
rect 8404 21524 8410 21588
rect 9029 21586 9095 21589
rect 9213 21586 9279 21589
rect 9673 21586 9739 21589
rect 9029 21584 9279 21586
rect 9029 21528 9034 21584
rect 9090 21528 9218 21584
rect 9274 21528 9279 21584
rect 9029 21526 9279 21528
rect 9029 21523 9095 21526
rect 9213 21523 9279 21526
rect 9630 21584 9739 21586
rect 9630 21528 9678 21584
rect 9734 21528 9739 21584
rect 9630 21523 9739 21528
rect 9806 21524 9812 21588
rect 9876 21586 9882 21588
rect 10542 21586 10548 21588
rect 9876 21526 10548 21586
rect 9876 21524 9882 21526
rect 10542 21524 10548 21526
rect 10612 21524 10618 21588
rect 3141 21450 3207 21453
rect 6821 21450 6887 21453
rect 3141 21448 6887 21450
rect 3141 21392 3146 21448
rect 3202 21392 6826 21448
rect 6882 21392 6887 21448
rect 3141 21390 6887 21392
rect 3141 21387 3207 21390
rect 6821 21387 6887 21390
rect 3233 21314 3299 21317
rect 4061 21314 4127 21317
rect 3233 21312 4127 21314
rect 3233 21256 3238 21312
rect 3294 21256 4066 21312
rect 4122 21256 4127 21312
rect 3233 21254 4127 21256
rect 3233 21251 3299 21254
rect 4061 21251 4127 21254
rect 5349 21314 5415 21317
rect 5901 21314 5967 21317
rect 5349 21312 5967 21314
rect 5349 21256 5354 21312
rect 5410 21256 5906 21312
rect 5962 21256 5967 21312
rect 5349 21254 5967 21256
rect 5349 21251 5415 21254
rect 5901 21251 5967 21254
rect 6269 21314 6335 21317
rect 7189 21314 7255 21317
rect 6269 21312 7255 21314
rect 6269 21256 6274 21312
rect 6330 21256 7194 21312
rect 7250 21256 7255 21312
rect 6269 21254 7255 21256
rect 9630 21314 9690 21523
rect 9765 21314 9831 21317
rect 9630 21312 9831 21314
rect 9630 21256 9770 21312
rect 9826 21256 9831 21312
rect 9630 21254 9831 21256
rect 6269 21251 6335 21254
rect 7189 21251 7255 21254
rect 9765 21251 9831 21254
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 10718 21248 11034 21249
rect 10718 21184 10724 21248
rect 10788 21184 10804 21248
rect 10868 21184 10884 21248
rect 10948 21184 10964 21248
rect 11028 21184 11034 21248
rect 10718 21183 11034 21184
rect 1526 21116 1532 21180
rect 1596 21178 1602 21180
rect 3325 21178 3391 21181
rect 1596 21176 3391 21178
rect 1596 21120 3330 21176
rect 3386 21120 3391 21176
rect 1596 21118 3391 21120
rect 1596 21116 1602 21118
rect 3325 21115 3391 21118
rect 4797 21178 4863 21181
rect 5533 21180 5599 21181
rect 5390 21178 5396 21180
rect 4797 21176 5396 21178
rect 4797 21120 4802 21176
rect 4858 21120 5396 21176
rect 4797 21118 5396 21120
rect 4797 21115 4863 21118
rect 5390 21116 5396 21118
rect 5460 21116 5466 21180
rect 5533 21176 5580 21180
rect 5644 21178 5650 21180
rect 5533 21120 5538 21176
rect 5533 21116 5580 21120
rect 5644 21118 5690 21178
rect 5644 21116 5650 21118
rect 5533 21115 5599 21116
rect 3328 21042 3388 21115
rect 4705 21042 4771 21045
rect 3328 21040 4771 21042
rect 3328 20984 4710 21040
rect 4766 20984 4771 21040
rect 3328 20982 4771 20984
rect 4705 20979 4771 20982
rect 4981 21042 5047 21045
rect 6085 21042 6151 21045
rect 4981 21040 6151 21042
rect 4981 20984 4986 21040
rect 5042 20984 6090 21040
rect 6146 20984 6151 21040
rect 4981 20982 6151 20984
rect 4981 20979 5047 20982
rect 6085 20979 6151 20982
rect 9213 21042 9279 21045
rect 10133 21042 10199 21045
rect 9213 21040 10199 21042
rect 9213 20984 9218 21040
rect 9274 20984 10138 21040
rect 10194 20984 10199 21040
rect 9213 20982 10199 20984
rect 9213 20979 9279 20982
rect 10133 20979 10199 20982
rect 3141 20906 3207 20909
rect 4797 20906 4863 20909
rect 3141 20904 4863 20906
rect 3141 20848 3146 20904
rect 3202 20848 4802 20904
rect 4858 20848 4863 20904
rect 3141 20846 4863 20848
rect 3141 20843 3207 20846
rect 4797 20843 4863 20846
rect 5993 20906 6059 20909
rect 7598 20906 7604 20908
rect 5993 20904 7604 20906
rect 5993 20848 5998 20904
rect 6054 20848 7604 20904
rect 5993 20846 7604 20848
rect 5993 20843 6059 20846
rect 7598 20844 7604 20846
rect 7668 20906 7674 20908
rect 7833 20906 7899 20909
rect 7668 20904 7899 20906
rect 7668 20848 7838 20904
rect 7894 20848 7899 20904
rect 7668 20846 7899 20848
rect 7668 20844 7674 20846
rect 7833 20843 7899 20846
rect 8702 20844 8708 20908
rect 8772 20906 8778 20908
rect 8845 20906 8911 20909
rect 8772 20904 8911 20906
rect 8772 20848 8850 20904
rect 8906 20848 8911 20904
rect 8772 20846 8911 20848
rect 8772 20844 8778 20846
rect 8845 20843 8911 20846
rect 9029 20906 9095 20909
rect 10041 20906 10107 20909
rect 9029 20904 10107 20906
rect 9029 20848 9034 20904
rect 9090 20848 10046 20904
rect 10102 20848 10107 20904
rect 9029 20846 10107 20848
rect 9029 20843 9095 20846
rect 10041 20843 10107 20846
rect 1301 20770 1367 20773
rect 3325 20770 3391 20773
rect 1301 20768 3391 20770
rect 1301 20712 1306 20768
rect 1362 20712 3330 20768
rect 3386 20712 3391 20768
rect 1301 20710 3391 20712
rect 1301 20707 1367 20710
rect 3325 20707 3391 20710
rect 4245 20770 4311 20773
rect 5022 20770 5028 20772
rect 4245 20768 5028 20770
rect 4245 20712 4250 20768
rect 4306 20712 5028 20768
rect 4245 20710 5028 20712
rect 4245 20707 4311 20710
rect 5022 20708 5028 20710
rect 5092 20708 5098 20772
rect 5165 20770 5231 20773
rect 8385 20770 8451 20773
rect 5165 20768 8451 20770
rect 5165 20712 5170 20768
rect 5226 20712 8390 20768
rect 8446 20712 8451 20768
rect 5165 20710 8451 20712
rect 5165 20707 5231 20710
rect 8385 20707 8451 20710
rect 9121 20770 9187 20773
rect 9622 20770 9628 20772
rect 9121 20768 9628 20770
rect 9121 20712 9126 20768
rect 9182 20712 9628 20768
rect 9121 20710 9628 20712
rect 9121 20707 9187 20710
rect 9622 20708 9628 20710
rect 9692 20708 9698 20772
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 10058 20704 10374 20705
rect 10058 20640 10064 20704
rect 10128 20640 10144 20704
rect 10208 20640 10224 20704
rect 10288 20640 10304 20704
rect 10368 20640 10374 20704
rect 10058 20639 10374 20640
rect 974 20572 980 20636
rect 1044 20634 1050 20636
rect 1117 20634 1183 20637
rect 1044 20632 1183 20634
rect 1044 20576 1122 20632
rect 1178 20576 1183 20632
rect 1044 20574 1183 20576
rect 1044 20572 1050 20574
rect 1117 20571 1183 20574
rect 2129 20634 2195 20637
rect 2446 20634 2452 20636
rect 2129 20632 2452 20634
rect 2129 20576 2134 20632
rect 2190 20576 2452 20632
rect 2129 20574 2452 20576
rect 2129 20571 2195 20574
rect 2446 20572 2452 20574
rect 2516 20634 2522 20636
rect 3325 20634 3391 20637
rect 2516 20632 3391 20634
rect 2516 20576 3330 20632
rect 3386 20576 3391 20632
rect 2516 20574 3391 20576
rect 2516 20572 2522 20574
rect 3325 20571 3391 20574
rect 54 20436 60 20500
rect 124 20498 130 20500
rect 1393 20498 1459 20501
rect 124 20496 1459 20498
rect 124 20440 1398 20496
rect 1454 20440 1459 20496
rect 124 20438 1459 20440
rect 124 20436 130 20438
rect 1393 20435 1459 20438
rect 4061 20498 4127 20501
rect 5206 20498 5212 20500
rect 4061 20496 5212 20498
rect 4061 20440 4066 20496
rect 4122 20440 5212 20496
rect 4061 20438 5212 20440
rect 4061 20435 4127 20438
rect 5206 20436 5212 20438
rect 5276 20498 5282 20500
rect 7557 20498 7623 20501
rect 5276 20496 7623 20498
rect 5276 20440 7562 20496
rect 7618 20440 7623 20496
rect 5276 20438 7623 20440
rect 5276 20436 5282 20438
rect 7557 20435 7623 20438
rect 8477 20500 8543 20501
rect 8477 20496 8524 20500
rect 8588 20498 8594 20500
rect 8477 20440 8482 20496
rect 8477 20436 8524 20440
rect 8588 20438 8634 20498
rect 8588 20436 8594 20438
rect 8477 20435 8543 20436
rect 2773 20362 2839 20365
rect 5073 20362 5139 20365
rect 2773 20360 5139 20362
rect 2773 20304 2778 20360
rect 2834 20304 5078 20360
rect 5134 20304 5139 20360
rect 2773 20302 5139 20304
rect 2773 20299 2839 20302
rect 5073 20299 5139 20302
rect 6678 20300 6684 20364
rect 6748 20362 6754 20364
rect 6821 20362 6887 20365
rect 6748 20360 6887 20362
rect 6748 20304 6826 20360
rect 6882 20304 6887 20360
rect 6748 20302 6887 20304
rect 6748 20300 6754 20302
rect 6821 20299 6887 20302
rect 7281 20362 7347 20365
rect 10685 20362 10751 20365
rect 7281 20360 10751 20362
rect 7281 20304 7286 20360
rect 7342 20304 10690 20360
rect 10746 20304 10751 20360
rect 7281 20302 10751 20304
rect 7281 20299 7347 20302
rect 10685 20299 10751 20302
rect 2446 20164 2452 20228
rect 2516 20226 2522 20228
rect 4102 20226 4108 20228
rect 2516 20166 4108 20226
rect 2516 20164 2522 20166
rect 4102 20164 4108 20166
rect 4172 20164 4178 20228
rect 5390 20164 5396 20228
rect 5460 20226 5466 20228
rect 6862 20226 6868 20228
rect 5460 20166 6868 20226
rect 5460 20164 5466 20166
rect 6862 20164 6868 20166
rect 6932 20226 6938 20228
rect 9121 20226 9187 20229
rect 6932 20224 9187 20226
rect 6932 20168 9126 20224
rect 9182 20168 9187 20224
rect 6932 20166 9187 20168
rect 6932 20164 6938 20166
rect 9121 20163 9187 20166
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 10718 20160 11034 20161
rect 10718 20096 10724 20160
rect 10788 20096 10804 20160
rect 10868 20096 10884 20160
rect 10948 20096 10964 20160
rect 11028 20096 11034 20160
rect 10718 20095 11034 20096
rect 5625 20090 5691 20093
rect 5490 20088 5691 20090
rect 5490 20032 5630 20088
rect 5686 20032 5691 20088
rect 5490 20030 5691 20032
rect 2078 19892 2084 19956
rect 2148 19954 2154 19956
rect 2773 19954 2839 19957
rect 2148 19952 2839 19954
rect 2148 19896 2778 19952
rect 2834 19896 2839 19952
rect 2148 19894 2839 19896
rect 2148 19892 2154 19894
rect 2773 19891 2839 19894
rect 4521 19954 4587 19957
rect 5490 19954 5550 20030
rect 5625 20027 5691 20030
rect 6085 20090 6151 20093
rect 6678 20090 6684 20092
rect 6085 20088 6684 20090
rect 6085 20032 6090 20088
rect 6146 20032 6684 20088
rect 6085 20030 6684 20032
rect 6085 20027 6151 20030
rect 6678 20028 6684 20030
rect 6748 20090 6754 20092
rect 7741 20090 7807 20093
rect 6748 20088 7807 20090
rect 6748 20032 7746 20088
rect 7802 20032 7807 20088
rect 6748 20030 7807 20032
rect 6748 20028 6754 20030
rect 7741 20027 7807 20030
rect 4521 19952 5550 19954
rect 4521 19896 4526 19952
rect 4582 19896 5550 19952
rect 4521 19894 5550 19896
rect 5628 19954 5688 20027
rect 7925 19954 7991 19957
rect 5628 19952 7991 19954
rect 5628 19896 7930 19952
rect 7986 19896 7991 19952
rect 5628 19894 7991 19896
rect 4521 19891 4587 19894
rect 7925 19891 7991 19894
rect 3233 19818 3299 19821
rect 5717 19818 5783 19821
rect 6310 19818 6316 19820
rect 3233 19816 6316 19818
rect 3233 19760 3238 19816
rect 3294 19760 5722 19816
rect 5778 19760 6316 19816
rect 3233 19758 6316 19760
rect 3233 19755 3299 19758
rect 5717 19755 5783 19758
rect 6310 19756 6316 19758
rect 6380 19756 6386 19820
rect 4061 19682 4127 19685
rect 5625 19682 5691 19685
rect 6913 19682 6979 19685
rect 4061 19680 6979 19682
rect 4061 19624 4066 19680
rect 4122 19624 5630 19680
rect 5686 19624 6918 19680
rect 6974 19624 6979 19680
rect 4061 19622 6979 19624
rect 4061 19619 4127 19622
rect 5625 19619 5691 19622
rect 6913 19619 6979 19622
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 3658 19551 3974 19552
rect 10058 19616 10374 19617
rect 10058 19552 10064 19616
rect 10128 19552 10144 19616
rect 10208 19552 10224 19616
rect 10288 19552 10304 19616
rect 10368 19552 10374 19616
rect 10058 19551 10374 19552
rect 4981 19546 5047 19549
rect 8661 19546 8727 19549
rect 4981 19544 8727 19546
rect 4981 19488 4986 19544
rect 5042 19488 8666 19544
rect 8722 19488 8727 19544
rect 4981 19486 8727 19488
rect 4981 19483 5047 19486
rect 8661 19483 8727 19486
rect 8886 19484 8892 19548
rect 8956 19546 8962 19548
rect 9121 19546 9187 19549
rect 8956 19544 9187 19546
rect 8956 19488 9126 19544
rect 9182 19488 9187 19544
rect 8956 19486 9187 19488
rect 8956 19484 8962 19486
rect 9121 19483 9187 19486
rect 289 19410 355 19413
rect 3233 19410 3299 19413
rect 5901 19410 5967 19413
rect 289 19408 1410 19410
rect 289 19352 294 19408
rect 350 19352 1410 19408
rect 289 19350 1410 19352
rect 289 19347 355 19350
rect 1350 19277 1410 19350
rect 3233 19408 5967 19410
rect 3233 19352 3238 19408
rect 3294 19352 5906 19408
rect 5962 19352 5967 19408
rect 3233 19350 5967 19352
rect 3233 19347 3299 19350
rect 5901 19347 5967 19350
rect 7046 19348 7052 19412
rect 7116 19410 7122 19412
rect 7649 19410 7715 19413
rect 7116 19408 7715 19410
rect 7116 19352 7654 19408
rect 7710 19352 7715 19408
rect 7116 19350 7715 19352
rect 7116 19348 7122 19350
rect 7649 19347 7715 19350
rect 1350 19272 1459 19277
rect 1350 19216 1398 19272
rect 1454 19216 1459 19272
rect 1350 19214 1459 19216
rect 1393 19211 1459 19214
rect 2630 19212 2636 19276
rect 2700 19274 2706 19276
rect 4337 19274 4403 19277
rect 2700 19272 4403 19274
rect 2700 19216 4342 19272
rect 4398 19216 4403 19272
rect 2700 19214 4403 19216
rect 2700 19212 2706 19214
rect 4337 19211 4403 19214
rect 4521 19274 4587 19277
rect 5533 19274 5599 19277
rect 4521 19272 5599 19274
rect 4521 19216 4526 19272
rect 4582 19216 5538 19272
rect 5594 19216 5599 19272
rect 4521 19214 5599 19216
rect 4521 19211 4587 19214
rect 5533 19211 5599 19214
rect 11237 19276 11303 19277
rect 11237 19272 11284 19276
rect 11348 19274 11354 19276
rect 11237 19216 11242 19272
rect 11237 19212 11284 19216
rect 11348 19214 11394 19274
rect 11348 19212 11354 19214
rect 11237 19211 11303 19212
rect 5625 19138 5691 19141
rect 6310 19138 6316 19140
rect 5625 19136 6316 19138
rect 5625 19080 5630 19136
rect 5686 19080 6316 19136
rect 5625 19078 6316 19080
rect 5625 19075 5691 19078
rect 6310 19076 6316 19078
rect 6380 19076 6386 19140
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 10718 19072 11034 19073
rect 10718 19008 10724 19072
rect 10788 19008 10804 19072
rect 10868 19008 10884 19072
rect 10948 19008 10964 19072
rect 11028 19008 11034 19072
rect 10718 19007 11034 19008
rect 4705 19002 4771 19005
rect 6085 19002 6151 19005
rect 4705 19000 6151 19002
rect 4705 18944 4710 19000
rect 4766 18944 6090 19000
rect 6146 18944 6151 19000
rect 4705 18942 6151 18944
rect 4705 18939 4771 18942
rect 6085 18939 6151 18942
rect 2630 18804 2636 18868
rect 2700 18866 2706 18868
rect 3141 18866 3207 18869
rect 5073 18866 5139 18869
rect 6821 18866 6887 18869
rect 2700 18864 6887 18866
rect 2700 18808 3146 18864
rect 3202 18808 5078 18864
rect 5134 18808 6826 18864
rect 6882 18808 6887 18864
rect 2700 18806 6887 18808
rect 2700 18804 2706 18806
rect 3141 18803 3207 18806
rect 5073 18803 5139 18806
rect 6821 18803 6887 18806
rect 9121 18866 9187 18869
rect 11278 18866 11284 18868
rect 9121 18864 11284 18866
rect 9121 18808 9126 18864
rect 9182 18808 11284 18864
rect 9121 18806 11284 18808
rect 9121 18803 9187 18806
rect 11278 18804 11284 18806
rect 11348 18804 11354 18868
rect 3877 18730 3943 18733
rect 5022 18730 5028 18732
rect 3877 18728 5028 18730
rect 3877 18672 3882 18728
rect 3938 18672 5028 18728
rect 3877 18670 5028 18672
rect 3877 18667 3943 18670
rect 5022 18668 5028 18670
rect 5092 18668 5098 18732
rect 5717 18730 5783 18733
rect 8017 18730 8083 18733
rect 8385 18730 8451 18733
rect 5717 18728 8451 18730
rect 5717 18672 5722 18728
rect 5778 18672 8022 18728
rect 8078 18672 8390 18728
rect 8446 18672 8451 18728
rect 5717 18670 8451 18672
rect 5717 18667 5783 18670
rect 8017 18667 8083 18670
rect 8385 18667 8451 18670
rect 9673 18730 9739 18733
rect 9806 18730 9812 18732
rect 9673 18728 9812 18730
rect 9673 18672 9678 18728
rect 9734 18672 9812 18728
rect 9673 18670 9812 18672
rect 9673 18667 9739 18670
rect 9806 18668 9812 18670
rect 9876 18668 9882 18732
rect 4153 18594 4219 18597
rect 5073 18594 5139 18597
rect 4153 18592 5139 18594
rect 4153 18536 4158 18592
rect 4214 18536 5078 18592
rect 5134 18536 5139 18592
rect 4153 18534 5139 18536
rect 4153 18531 4219 18534
rect 5073 18531 5139 18534
rect 5533 18594 5599 18597
rect 7281 18594 7347 18597
rect 7414 18594 7420 18596
rect 5533 18592 6148 18594
rect 5533 18536 5538 18592
rect 5594 18536 6148 18592
rect 5533 18534 6148 18536
rect 5533 18531 5599 18534
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 6088 18461 6148 18534
rect 7281 18592 7420 18594
rect 7281 18536 7286 18592
rect 7342 18536 7420 18592
rect 7281 18534 7420 18536
rect 7281 18531 7347 18534
rect 7414 18532 7420 18534
rect 7484 18532 7490 18596
rect 8334 18532 8340 18596
rect 8404 18594 8410 18596
rect 9121 18594 9187 18597
rect 8404 18592 9187 18594
rect 8404 18536 9126 18592
rect 9182 18536 9187 18592
rect 8404 18534 9187 18536
rect 8404 18532 8410 18534
rect 9121 18531 9187 18534
rect 10058 18528 10374 18529
rect 10058 18464 10064 18528
rect 10128 18464 10144 18528
rect 10208 18464 10224 18528
rect 10288 18464 10304 18528
rect 10368 18464 10374 18528
rect 10058 18463 10374 18464
rect 4337 18458 4403 18461
rect 4705 18458 4771 18461
rect 4337 18456 4771 18458
rect 4337 18400 4342 18456
rect 4398 18400 4710 18456
rect 4766 18400 4771 18456
rect 4337 18398 4771 18400
rect 4337 18395 4403 18398
rect 4705 18395 4771 18398
rect 5165 18458 5231 18461
rect 5717 18458 5783 18461
rect 5165 18456 5783 18458
rect 5165 18400 5170 18456
rect 5226 18400 5722 18456
rect 5778 18400 5783 18456
rect 5165 18398 5783 18400
rect 5165 18395 5231 18398
rect 5717 18395 5783 18398
rect 6085 18456 6151 18461
rect 6085 18400 6090 18456
rect 6146 18400 6151 18456
rect 6085 18395 6151 18400
rect 6821 18458 6887 18461
rect 7281 18458 7347 18461
rect 8293 18458 8359 18461
rect 6821 18456 8359 18458
rect 6821 18400 6826 18456
rect 6882 18400 7286 18456
rect 7342 18400 8298 18456
rect 8354 18400 8359 18456
rect 6821 18398 8359 18400
rect 6821 18395 6887 18398
rect 7281 18395 7347 18398
rect 8293 18395 8359 18398
rect 4838 18322 4844 18324
rect 3420 18262 4844 18322
rect 3420 18189 3480 18262
rect 4838 18260 4844 18262
rect 4908 18260 4914 18324
rect 5073 18322 5139 18325
rect 5717 18324 5783 18325
rect 5206 18322 5212 18324
rect 5073 18320 5212 18322
rect 5073 18264 5078 18320
rect 5134 18264 5212 18320
rect 5073 18262 5212 18264
rect 5073 18259 5139 18262
rect 5206 18260 5212 18262
rect 5276 18260 5282 18324
rect 5717 18320 5764 18324
rect 5828 18322 5834 18324
rect 7465 18322 7531 18325
rect 7649 18322 7715 18325
rect 11145 18324 11211 18325
rect 11094 18322 11100 18324
rect 5717 18264 5722 18320
rect 5717 18260 5764 18264
rect 5828 18262 5874 18322
rect 6364 18320 7715 18322
rect 6364 18264 7470 18320
rect 7526 18264 7654 18320
rect 7710 18264 7715 18320
rect 6364 18262 7715 18264
rect 11054 18262 11100 18322
rect 11164 18320 11211 18324
rect 11206 18264 11211 18320
rect 5828 18260 5834 18262
rect 5717 18259 5783 18260
rect 3417 18184 3483 18189
rect 3417 18128 3422 18184
rect 3478 18128 3483 18184
rect 3417 18123 3483 18128
rect 4102 18124 4108 18188
rect 4172 18186 4178 18188
rect 4981 18186 5047 18189
rect 4172 18184 5047 18186
rect 4172 18128 4986 18184
rect 5042 18128 5047 18184
rect 4172 18126 5047 18128
rect 4172 18124 4178 18126
rect 4981 18123 5047 18126
rect 5165 18186 5231 18189
rect 5390 18186 5396 18188
rect 5165 18184 5396 18186
rect 5165 18128 5170 18184
rect 5226 18128 5396 18184
rect 5165 18126 5396 18128
rect 5165 18123 5231 18126
rect 5390 18124 5396 18126
rect 5460 18186 5466 18188
rect 5533 18186 5599 18189
rect 5460 18184 5599 18186
rect 5460 18128 5538 18184
rect 5594 18128 5599 18184
rect 5460 18126 5599 18128
rect 5460 18124 5466 18126
rect 5533 18123 5599 18126
rect 5717 18186 5783 18189
rect 6364 18186 6424 18262
rect 7465 18259 7531 18262
rect 7649 18259 7715 18262
rect 11094 18260 11100 18262
rect 11164 18260 11211 18264
rect 11145 18259 11211 18260
rect 5717 18184 6424 18186
rect 5717 18128 5722 18184
rect 5778 18128 6424 18184
rect 5717 18126 6424 18128
rect 6545 18186 6611 18189
rect 6862 18186 6868 18188
rect 6545 18184 6868 18186
rect 6545 18128 6550 18184
rect 6606 18128 6868 18184
rect 6545 18126 6868 18128
rect 5717 18123 5783 18126
rect 6545 18123 6611 18126
rect 6862 18124 6868 18126
rect 6932 18186 6938 18188
rect 7465 18186 7531 18189
rect 7966 18186 7972 18188
rect 6932 18184 7531 18186
rect 6932 18128 7470 18184
rect 7526 18128 7531 18184
rect 6932 18126 7531 18128
rect 6932 18124 6938 18126
rect 7465 18123 7531 18126
rect 7606 18126 7972 18186
rect 657 18052 723 18053
rect 606 18050 612 18052
rect 566 17990 612 18050
rect 676 18048 723 18052
rect 718 17992 723 18048
rect 606 17988 612 17990
rect 676 17988 723 17992
rect 657 17987 723 17988
rect 2405 18050 2471 18053
rect 2814 18050 2820 18052
rect 2405 18048 2820 18050
rect 2405 17992 2410 18048
rect 2466 17992 2820 18048
rect 2405 17990 2820 17992
rect 2405 17987 2471 17990
rect 2814 17988 2820 17990
rect 2884 17988 2890 18052
rect 4797 18048 4863 18053
rect 4797 17992 4802 18048
rect 4858 17992 4863 18048
rect 4797 17987 4863 17992
rect 5022 17988 5028 18052
rect 5092 18050 5098 18052
rect 5165 18050 5231 18053
rect 5092 18048 5231 18050
rect 5092 17992 5170 18048
rect 5226 17992 5231 18048
rect 5092 17990 5231 17992
rect 5092 17988 5098 17990
rect 5165 17987 5231 17990
rect 6545 18050 6611 18053
rect 7606 18050 7666 18126
rect 7966 18124 7972 18126
rect 8036 18124 8042 18188
rect 6545 18048 7666 18050
rect 6545 17992 6550 18048
rect 6606 17992 7666 18048
rect 6545 17990 7666 17992
rect 7741 18050 7807 18053
rect 7925 18050 7991 18053
rect 7741 18048 7991 18050
rect 7741 17992 7746 18048
rect 7802 17992 7930 18048
rect 7986 17992 7991 18048
rect 7741 17990 7991 17992
rect 6545 17987 6611 17990
rect 7741 17987 7807 17990
rect 7925 17987 7991 17990
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 4800 17917 4860 17987
rect 10718 17984 11034 17985
rect 10718 17920 10724 17984
rect 10788 17920 10804 17984
rect 10868 17920 10884 17984
rect 10948 17920 10964 17984
rect 11028 17920 11034 17984
rect 10718 17919 11034 17920
rect 54 17852 60 17916
rect 124 17914 130 17916
rect 1853 17914 1919 17917
rect 124 17912 1919 17914
rect 124 17856 1858 17912
rect 1914 17856 1919 17912
rect 124 17854 1919 17856
rect 124 17852 130 17854
rect 1853 17851 1919 17854
rect 4797 17912 4863 17917
rect 4797 17856 4802 17912
rect 4858 17856 4863 17912
rect 4797 17851 4863 17856
rect 7189 17912 7255 17917
rect 7189 17856 7194 17912
rect 7250 17856 7255 17912
rect 7189 17851 7255 17856
rect 7373 17914 7439 17917
rect 7557 17914 7623 17917
rect 7373 17912 7623 17914
rect 7373 17856 7378 17912
rect 7434 17856 7562 17912
rect 7618 17856 7623 17912
rect 7373 17854 7623 17856
rect 7373 17851 7439 17854
rect 7557 17851 7623 17854
rect 8017 17914 8083 17917
rect 8017 17912 8218 17914
rect 8017 17856 8022 17912
rect 8078 17856 8218 17912
rect 8017 17854 8218 17856
rect 8017 17851 8083 17854
rect 3969 17778 4035 17781
rect 4705 17778 4771 17781
rect 3969 17776 4771 17778
rect 3969 17720 3974 17776
rect 4030 17720 4710 17776
rect 4766 17720 4771 17776
rect 3969 17718 4771 17720
rect 3969 17715 4035 17718
rect 4705 17715 4771 17718
rect 5022 17716 5028 17780
rect 5092 17778 5098 17780
rect 5257 17778 5323 17781
rect 5092 17776 5323 17778
rect 5092 17720 5262 17776
rect 5318 17720 5323 17776
rect 5092 17718 5323 17720
rect 5092 17716 5098 17718
rect 5257 17715 5323 17718
rect 3785 17642 3851 17645
rect 5717 17642 5783 17645
rect 6269 17644 6335 17645
rect 6269 17642 6316 17644
rect 3785 17640 5783 17642
rect 3785 17584 3790 17640
rect 3846 17584 5722 17640
rect 5778 17584 5783 17640
rect 3785 17582 5783 17584
rect 6224 17640 6316 17642
rect 6224 17584 6274 17640
rect 6224 17582 6316 17584
rect 3785 17579 3851 17582
rect 5717 17579 5783 17582
rect 6269 17580 6316 17582
rect 6380 17580 6386 17644
rect 7192 17642 7252 17851
rect 8158 17645 8218 17854
rect 7465 17642 7531 17645
rect 7192 17640 7531 17642
rect 7192 17584 7470 17640
rect 7526 17584 7531 17640
rect 7192 17582 7531 17584
rect 8158 17640 8267 17645
rect 8477 17644 8543 17645
rect 8477 17642 8524 17644
rect 8158 17584 8206 17640
rect 8262 17584 8267 17640
rect 8158 17582 8267 17584
rect 8432 17640 8524 17642
rect 8432 17584 8482 17640
rect 8432 17582 8524 17584
rect 6269 17579 6335 17580
rect 7465 17579 7531 17582
rect 8201 17579 8267 17582
rect 8477 17580 8524 17582
rect 8588 17580 8594 17644
rect 9438 17580 9444 17644
rect 9508 17642 9514 17644
rect 9673 17642 9739 17645
rect 9508 17640 9739 17642
rect 9508 17584 9678 17640
rect 9734 17584 9739 17640
rect 9508 17582 9739 17584
rect 9508 17580 9514 17582
rect 8477 17579 8543 17580
rect 9673 17579 9739 17582
rect 289 17508 355 17509
rect 238 17444 244 17508
rect 308 17506 355 17508
rect 4429 17506 4495 17509
rect 5257 17506 5323 17509
rect 308 17504 400 17506
rect 350 17448 400 17504
rect 308 17446 400 17448
rect 4429 17504 5323 17506
rect 4429 17448 4434 17504
rect 4490 17448 5262 17504
rect 5318 17448 5323 17504
rect 4429 17446 5323 17448
rect 308 17444 355 17446
rect 289 17443 355 17444
rect 4429 17443 4495 17446
rect 5257 17443 5323 17446
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 10058 17440 10374 17441
rect 10058 17376 10064 17440
rect 10128 17376 10144 17440
rect 10208 17376 10224 17440
rect 10288 17376 10304 17440
rect 10368 17376 10374 17440
rect 10058 17375 10374 17376
rect 3417 17368 3483 17373
rect 3417 17312 3422 17368
rect 3478 17312 3483 17368
rect 3417 17307 3483 17312
rect 4797 17370 4863 17373
rect 6269 17370 6335 17373
rect 4797 17368 6335 17370
rect 4797 17312 4802 17368
rect 4858 17312 6274 17368
rect 6330 17312 6335 17368
rect 4797 17310 6335 17312
rect 4797 17307 4863 17310
rect 6269 17307 6335 17310
rect 6637 17370 6703 17373
rect 7557 17370 7623 17373
rect 6637 17368 7623 17370
rect 6637 17312 6642 17368
rect 6698 17312 7562 17368
rect 7618 17312 7623 17368
rect 6637 17310 7623 17312
rect 6637 17307 6703 17310
rect 7557 17307 7623 17310
rect 0 17234 400 17264
rect 933 17234 999 17237
rect 1485 17236 1551 17237
rect 1485 17234 1532 17236
rect 0 17232 999 17234
rect 0 17176 938 17232
rect 994 17176 999 17232
rect 0 17174 999 17176
rect 1440 17232 1532 17234
rect 1440 17176 1490 17232
rect 1440 17174 1532 17176
rect 0 17144 400 17174
rect 933 17171 999 17174
rect 1485 17172 1532 17174
rect 1596 17172 1602 17236
rect 3141 17234 3207 17237
rect 3420 17234 3480 17307
rect 3141 17232 3480 17234
rect 3141 17176 3146 17232
rect 3202 17176 3480 17232
rect 3141 17174 3480 17176
rect 3693 17234 3759 17237
rect 4245 17234 4311 17237
rect 3693 17232 4311 17234
rect 3693 17176 3698 17232
rect 3754 17176 4250 17232
rect 4306 17176 4311 17232
rect 3693 17174 4311 17176
rect 1485 17171 1551 17172
rect 3141 17171 3207 17174
rect 3693 17171 3759 17174
rect 4245 17171 4311 17174
rect 4521 17234 4587 17237
rect 4838 17234 4844 17236
rect 4521 17232 4844 17234
rect 4521 17176 4526 17232
rect 4582 17176 4844 17232
rect 4521 17174 4844 17176
rect 4521 17171 4587 17174
rect 4838 17172 4844 17174
rect 4908 17234 4914 17236
rect 6126 17234 6132 17236
rect 4908 17174 6132 17234
rect 4908 17172 4914 17174
rect 6126 17172 6132 17174
rect 6196 17172 6202 17236
rect 6678 17172 6684 17236
rect 6748 17234 6754 17236
rect 6821 17234 6887 17237
rect 6748 17232 6887 17234
rect 6748 17176 6826 17232
rect 6882 17176 6887 17232
rect 6748 17174 6887 17176
rect 6748 17172 6754 17174
rect 6821 17171 6887 17174
rect 8334 17172 8340 17236
rect 8404 17234 8410 17236
rect 9070 17234 9076 17236
rect 8404 17174 9076 17234
rect 8404 17172 8410 17174
rect 9070 17172 9076 17174
rect 9140 17172 9146 17236
rect 565 17098 631 17101
rect 1342 17098 1348 17100
rect 565 17096 1348 17098
rect 565 17040 570 17096
rect 626 17040 1348 17096
rect 565 17038 1348 17040
rect 565 17035 631 17038
rect 1342 17036 1348 17038
rect 1412 17036 1418 17100
rect 2865 17098 2931 17101
rect 3969 17098 4035 17101
rect 2865 17096 4035 17098
rect 2865 17040 2870 17096
rect 2926 17040 3974 17096
rect 4030 17040 4035 17096
rect 2865 17038 4035 17040
rect 2865 17035 2931 17038
rect 3969 17035 4035 17038
rect 4429 17098 4495 17101
rect 5717 17098 5783 17101
rect 4429 17096 5783 17098
rect 4429 17040 4434 17096
rect 4490 17040 5722 17096
rect 5778 17040 5783 17096
rect 4429 17038 5783 17040
rect 4429 17035 4495 17038
rect 5717 17035 5783 17038
rect 8477 17098 8543 17101
rect 9305 17098 9371 17101
rect 8477 17096 9371 17098
rect 8477 17040 8482 17096
rect 8538 17040 9310 17096
rect 9366 17040 9371 17096
rect 8477 17038 9371 17040
rect 8477 17035 8543 17038
rect 9305 17035 9371 17038
rect 0 16962 400 16992
rect 1117 16962 1183 16965
rect 2681 16964 2747 16965
rect 2630 16962 2636 16964
rect 0 16960 1183 16962
rect 0 16904 1122 16960
rect 1178 16904 1183 16960
rect 0 16902 1183 16904
rect 2590 16902 2636 16962
rect 2700 16962 2747 16964
rect 3785 16962 3851 16965
rect 2700 16960 3851 16962
rect 2742 16904 3790 16960
rect 3846 16904 3851 16960
rect 0 16872 400 16902
rect 1117 16899 1183 16902
rect 2630 16900 2636 16902
rect 2700 16902 3851 16904
rect 2700 16900 2747 16902
rect 2681 16899 2747 16900
rect 3785 16899 3851 16902
rect 4705 16962 4771 16965
rect 6862 16962 6868 16964
rect 4705 16960 6868 16962
rect 4705 16904 4710 16960
rect 4766 16904 6868 16960
rect 4705 16902 6868 16904
rect 4705 16899 4771 16902
rect 6862 16900 6868 16902
rect 6932 16900 6938 16964
rect 8109 16962 8175 16965
rect 8937 16962 9003 16965
rect 9765 16962 9831 16965
rect 8109 16960 9003 16962
rect 8109 16904 8114 16960
rect 8170 16904 8942 16960
rect 8998 16904 9003 16960
rect 8109 16902 9003 16904
rect 8109 16899 8175 16902
rect 8937 16899 9003 16902
rect 9630 16960 9831 16962
rect 9630 16904 9770 16960
rect 9826 16904 9831 16960
rect 9630 16902 9831 16904
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 1117 16826 1183 16829
rect 3366 16826 3372 16828
rect 1117 16824 3372 16826
rect 1117 16768 1122 16824
rect 1178 16768 3372 16824
rect 1117 16766 3372 16768
rect 1117 16763 1183 16766
rect 3366 16764 3372 16766
rect 3436 16764 3442 16828
rect 5441 16826 5507 16829
rect 6821 16826 6887 16829
rect 5441 16824 6887 16826
rect 5441 16768 5446 16824
rect 5502 16768 6826 16824
rect 6882 16768 6887 16824
rect 5441 16766 6887 16768
rect 5441 16763 5507 16766
rect 6821 16763 6887 16766
rect 7598 16764 7604 16828
rect 7668 16826 7674 16828
rect 9254 16826 9260 16828
rect 7668 16766 9260 16826
rect 7668 16764 7674 16766
rect 9254 16764 9260 16766
rect 9324 16764 9330 16828
rect 0 16693 400 16720
rect 9630 16693 9690 16902
rect 9765 16899 9831 16902
rect 10718 16896 11034 16897
rect 10718 16832 10724 16896
rect 10788 16832 10804 16896
rect 10868 16832 10884 16896
rect 10948 16832 10964 16896
rect 11028 16832 11034 16896
rect 10718 16831 11034 16832
rect 0 16688 447 16693
rect 0 16632 386 16688
rect 442 16632 447 16688
rect 0 16627 447 16632
rect 5901 16690 5967 16693
rect 6821 16690 6887 16693
rect 5901 16688 6887 16690
rect 5901 16632 5906 16688
rect 5962 16632 6826 16688
rect 6882 16632 6887 16688
rect 5901 16630 6887 16632
rect 5901 16627 5967 16630
rect 6821 16627 6887 16630
rect 8385 16690 8451 16693
rect 9121 16692 9187 16693
rect 9070 16690 9076 16692
rect 8385 16688 9076 16690
rect 9140 16690 9187 16692
rect 9140 16688 9232 16690
rect 8385 16632 8390 16688
rect 8446 16632 9076 16688
rect 9182 16632 9232 16688
rect 8385 16630 9076 16632
rect 8385 16627 8451 16630
rect 9070 16628 9076 16630
rect 9140 16630 9232 16632
rect 9630 16688 9739 16693
rect 9630 16632 9678 16688
rect 9734 16632 9739 16688
rect 9630 16630 9739 16632
rect 9140 16628 9187 16630
rect 9121 16627 9187 16628
rect 9673 16627 9739 16630
rect 0 16600 400 16627
rect 3877 16554 3943 16557
rect 4705 16554 4771 16557
rect 3877 16552 4771 16554
rect 3877 16496 3882 16552
rect 3938 16496 4710 16552
rect 4766 16496 4771 16552
rect 3877 16494 4771 16496
rect 3877 16491 3943 16494
rect 4705 16491 4771 16494
rect 6361 16554 6427 16557
rect 6545 16554 6611 16557
rect 6361 16552 6611 16554
rect 6361 16496 6366 16552
rect 6422 16496 6550 16552
rect 6606 16496 6611 16552
rect 6361 16494 6611 16496
rect 6361 16491 6427 16494
rect 6545 16491 6611 16494
rect 7230 16492 7236 16556
rect 7300 16554 7306 16556
rect 7925 16554 7991 16557
rect 7300 16552 7991 16554
rect 7300 16496 7930 16552
rect 7986 16496 7991 16552
rect 7300 16494 7991 16496
rect 7300 16492 7306 16494
rect 7925 16491 7991 16494
rect 8886 16492 8892 16556
rect 8956 16554 8962 16556
rect 9397 16554 9463 16557
rect 11237 16554 11303 16557
rect 8956 16552 11303 16554
rect 8956 16496 9402 16552
rect 9458 16496 11242 16552
rect 11298 16496 11303 16552
rect 8956 16494 11303 16496
rect 8956 16492 8962 16494
rect 9397 16491 9463 16494
rect 11237 16491 11303 16494
rect 0 16418 400 16448
rect 790 16418 796 16420
rect 0 16358 796 16418
rect 0 16328 400 16358
rect 790 16356 796 16358
rect 860 16356 866 16420
rect 6637 16418 6703 16421
rect 8702 16418 8708 16420
rect 6637 16416 8708 16418
rect 6637 16360 6642 16416
rect 6698 16360 8708 16416
rect 6637 16358 8708 16360
rect 6637 16355 6703 16358
rect 8702 16356 8708 16358
rect 8772 16356 8778 16420
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 10058 16352 10374 16353
rect 10058 16288 10064 16352
rect 10128 16288 10144 16352
rect 10208 16288 10224 16352
rect 10288 16288 10304 16352
rect 10368 16288 10374 16352
rect 10058 16287 10374 16288
rect 933 16146 999 16149
rect 1710 16146 1716 16148
rect 933 16144 1716 16146
rect 933 16088 938 16144
rect 994 16088 1716 16144
rect 933 16086 1716 16088
rect 933 16083 999 16086
rect 1710 16084 1716 16086
rect 1780 16084 1786 16148
rect 3182 16084 3188 16148
rect 3252 16146 3258 16148
rect 3693 16146 3759 16149
rect 3252 16144 3759 16146
rect 3252 16088 3698 16144
rect 3754 16088 3759 16144
rect 3252 16086 3759 16088
rect 3252 16084 3258 16086
rect 3693 16083 3759 16086
rect 841 15874 907 15877
rect 2998 15874 3004 15876
rect 841 15872 3004 15874
rect 841 15816 846 15872
rect 902 15816 3004 15872
rect 841 15814 3004 15816
rect 841 15811 907 15814
rect 2998 15812 3004 15814
rect 3068 15812 3074 15876
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 10718 15808 11034 15809
rect 10718 15744 10724 15808
rect 10788 15744 10804 15808
rect 10868 15744 10884 15808
rect 10948 15744 10964 15808
rect 11028 15744 11034 15808
rect 10718 15743 11034 15744
rect 8385 15738 8451 15741
rect 9765 15738 9831 15741
rect 8385 15736 9831 15738
rect 8385 15680 8390 15736
rect 8446 15680 9770 15736
rect 9826 15680 9831 15736
rect 8385 15678 9831 15680
rect 8385 15675 8451 15678
rect 9765 15675 9831 15678
rect 2773 15602 2839 15605
rect 8845 15602 8911 15605
rect 2773 15600 8911 15602
rect 2773 15544 2778 15600
rect 2834 15544 8850 15600
rect 8906 15544 8911 15600
rect 2773 15542 8911 15544
rect 2773 15539 2839 15542
rect 8845 15539 8911 15542
rect 7925 15466 7991 15469
rect 8201 15466 8267 15469
rect 8385 15468 8451 15469
rect 7925 15464 8267 15466
rect 7925 15408 7930 15464
rect 7986 15408 8206 15464
rect 8262 15408 8267 15464
rect 7925 15406 8267 15408
rect 7925 15403 7991 15406
rect 8201 15403 8267 15406
rect 8334 15404 8340 15468
rect 8404 15466 8451 15468
rect 10542 15466 10548 15468
rect 8404 15464 8496 15466
rect 8446 15408 8496 15464
rect 8404 15406 8496 15408
rect 9262 15406 10548 15466
rect 8404 15404 8451 15406
rect 8342 15403 8451 15404
rect 5574 15268 5580 15332
rect 5644 15268 5650 15332
rect 6545 15330 6611 15333
rect 8342 15330 8402 15403
rect 9262 15333 9322 15406
rect 10542 15404 10548 15406
rect 10612 15404 10618 15468
rect 6545 15328 8402 15330
rect 6545 15272 6550 15328
rect 6606 15272 8402 15328
rect 6545 15270 8402 15272
rect 9213 15328 9322 15333
rect 9213 15272 9218 15328
rect 9274 15272 9322 15328
rect 9213 15270 9322 15272
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 2221 15196 2287 15197
rect 2221 15194 2268 15196
rect 2176 15192 2268 15194
rect 2176 15136 2226 15192
rect 2176 15134 2268 15136
rect 2221 15132 2268 15134
rect 2332 15132 2338 15196
rect 4102 15132 4108 15196
rect 4172 15194 4178 15196
rect 4245 15194 4311 15197
rect 4172 15192 4311 15194
rect 4172 15136 4250 15192
rect 4306 15136 4311 15192
rect 4172 15134 4311 15136
rect 5582 15194 5642 15268
rect 6545 15267 6611 15270
rect 9213 15267 9279 15270
rect 10058 15264 10374 15265
rect 10058 15200 10064 15264
rect 10128 15200 10144 15264
rect 10208 15200 10224 15264
rect 10288 15200 10304 15264
rect 10368 15200 10374 15264
rect 10058 15199 10374 15200
rect 7557 15194 7623 15197
rect 5582 15192 7623 15194
rect 5582 15136 7562 15192
rect 7618 15136 7623 15192
rect 5582 15134 7623 15136
rect 4172 15132 4178 15134
rect 2221 15131 2287 15132
rect 4245 15131 4311 15134
rect 7557 15131 7623 15134
rect 5942 14996 5948 15060
rect 6012 15058 6018 15060
rect 6085 15058 6151 15061
rect 6012 15056 6151 15058
rect 6012 15000 6090 15056
rect 6146 15000 6151 15056
rect 6012 14998 6151 15000
rect 6012 14996 6018 14998
rect 6085 14995 6151 14998
rect 9254 14996 9260 15060
rect 9324 15058 9330 15060
rect 9397 15058 9463 15061
rect 9324 15056 9463 15058
rect 9324 15000 9402 15056
rect 9458 15000 9463 15056
rect 9324 14998 9463 15000
rect 9324 14996 9330 14998
rect 3969 14922 4035 14925
rect 6637 14922 6703 14925
rect 3969 14920 6703 14922
rect 3969 14864 3974 14920
rect 4030 14864 6642 14920
rect 6698 14864 6703 14920
rect 3969 14862 6703 14864
rect 3969 14859 4035 14862
rect 6637 14859 6703 14862
rect 8569 14922 8635 14925
rect 9262 14922 9322 14996
rect 9397 14995 9463 14998
rect 9622 14996 9628 15060
rect 9692 15058 9698 15060
rect 9949 15058 10015 15061
rect 9692 15056 10015 15058
rect 9692 15000 9954 15056
rect 10010 15000 10015 15056
rect 9692 14998 10015 15000
rect 9692 14996 9698 14998
rect 9949 14995 10015 14998
rect 8569 14920 9322 14922
rect 8569 14864 8574 14920
rect 8630 14864 9322 14920
rect 8569 14862 9322 14864
rect 8569 14859 8635 14862
rect 1761 14786 1827 14789
rect 3877 14786 3943 14789
rect 1761 14784 3943 14786
rect 1761 14728 1766 14784
rect 1822 14728 3882 14784
rect 3938 14728 3943 14784
rect 1761 14726 3943 14728
rect 1761 14723 1827 14726
rect 3877 14723 3943 14726
rect 8753 14786 8819 14789
rect 9581 14786 9647 14789
rect 8753 14784 9647 14786
rect 8753 14728 8758 14784
rect 8814 14728 9586 14784
rect 9642 14728 9647 14784
rect 8753 14726 9647 14728
rect 8753 14723 8819 14726
rect 9581 14723 9647 14726
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 10718 14720 11034 14721
rect 10718 14656 10724 14720
rect 10788 14656 10804 14720
rect 10868 14656 10884 14720
rect 10948 14656 10964 14720
rect 11028 14656 11034 14720
rect 10718 14655 11034 14656
rect 2681 14650 2747 14653
rect 2814 14650 2820 14652
rect 2681 14648 2820 14650
rect 2681 14592 2686 14648
rect 2742 14592 2820 14648
rect 2681 14590 2820 14592
rect 2681 14587 2747 14590
rect 2814 14588 2820 14590
rect 2884 14588 2890 14652
rect 8477 14514 8543 14517
rect 9397 14514 9463 14517
rect 8477 14512 9463 14514
rect 8477 14456 8482 14512
rect 8538 14456 9402 14512
rect 9458 14456 9463 14512
rect 8477 14454 9463 14456
rect 8477 14451 8543 14454
rect 9397 14451 9463 14454
rect 3693 14378 3759 14381
rect 4153 14378 4219 14381
rect 3693 14376 4219 14378
rect 3693 14320 3698 14376
rect 3754 14320 4158 14376
rect 4214 14320 4219 14376
rect 3693 14318 4219 14320
rect 3693 14315 3759 14318
rect 4153 14315 4219 14318
rect 5073 14242 5139 14245
rect 7373 14242 7439 14245
rect 5073 14240 7439 14242
rect 5073 14184 5078 14240
rect 5134 14184 7378 14240
rect 7434 14184 7439 14240
rect 5073 14182 7439 14184
rect 5073 14179 5139 14182
rect 7373 14179 7439 14182
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 10058 14176 10374 14177
rect 10058 14112 10064 14176
rect 10128 14112 10144 14176
rect 10208 14112 10224 14176
rect 10288 14112 10304 14176
rect 10368 14112 10374 14176
rect 10058 14111 10374 14112
rect 3785 13970 3851 13973
rect 5165 13970 5231 13973
rect 3785 13968 5231 13970
rect 3785 13912 3790 13968
rect 3846 13912 5170 13968
rect 5226 13912 5231 13968
rect 3785 13910 5231 13912
rect 3785 13907 3851 13910
rect 5165 13907 5231 13910
rect 8937 13970 9003 13973
rect 9489 13970 9555 13973
rect 8937 13968 9555 13970
rect 8937 13912 8942 13968
rect 8998 13912 9494 13968
rect 9550 13912 9555 13968
rect 8937 13910 9555 13912
rect 8937 13907 9003 13910
rect 9489 13907 9555 13910
rect 1526 13772 1532 13836
rect 1596 13834 1602 13836
rect 1669 13834 1735 13837
rect 1596 13832 1735 13834
rect 1596 13776 1674 13832
rect 1730 13776 1735 13832
rect 1596 13774 1735 13776
rect 1596 13772 1602 13774
rect 1669 13771 1735 13774
rect 3141 13834 3207 13837
rect 4838 13834 4844 13836
rect 3141 13832 4844 13834
rect 3141 13776 3146 13832
rect 3202 13776 4844 13832
rect 3141 13774 4844 13776
rect 3141 13771 3207 13774
rect 4838 13772 4844 13774
rect 4908 13772 4914 13836
rect 2998 13636 3004 13700
rect 3068 13698 3074 13700
rect 3233 13698 3299 13701
rect 3068 13696 3299 13698
rect 3068 13640 3238 13696
rect 3294 13640 3299 13696
rect 3068 13638 3299 13640
rect 3068 13636 3074 13638
rect 3233 13635 3299 13638
rect 7414 13636 7420 13700
rect 7484 13698 7490 13700
rect 7741 13698 7807 13701
rect 7484 13696 7807 13698
rect 7484 13640 7746 13696
rect 7802 13640 7807 13696
rect 7484 13638 7807 13640
rect 7484 13636 7490 13638
rect 7741 13635 7807 13638
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 10718 13632 11034 13633
rect 10718 13568 10724 13632
rect 10788 13568 10804 13632
rect 10868 13568 10884 13632
rect 10948 13568 10964 13632
rect 11028 13568 11034 13632
rect 10718 13567 11034 13568
rect 8109 13562 8175 13565
rect 9438 13562 9444 13564
rect 8109 13560 9444 13562
rect 8109 13504 8114 13560
rect 8170 13504 9444 13560
rect 8109 13502 9444 13504
rect 8109 13499 8175 13502
rect 9438 13500 9444 13502
rect 9508 13500 9514 13564
rect 2865 13428 2931 13429
rect 2814 13426 2820 13428
rect 2738 13366 2820 13426
rect 2884 13426 2931 13428
rect 4337 13426 4403 13429
rect 2884 13424 4403 13426
rect 2926 13368 4342 13424
rect 4398 13368 4403 13424
rect 2814 13364 2820 13366
rect 2884 13366 4403 13368
rect 2884 13364 2931 13366
rect 2865 13363 2931 13364
rect 4337 13363 4403 13366
rect 4889 13426 4955 13429
rect 5022 13426 5028 13428
rect 4889 13424 5028 13426
rect 4889 13368 4894 13424
rect 4950 13368 5028 13424
rect 4889 13366 5028 13368
rect 4889 13363 4955 13366
rect 5022 13364 5028 13366
rect 5092 13364 5098 13428
rect 2957 13290 3023 13293
rect 3233 13290 3299 13293
rect 2957 13288 3299 13290
rect 2957 13232 2962 13288
rect 3018 13232 3238 13288
rect 3294 13232 3299 13288
rect 2957 13230 3299 13232
rect 2957 13227 3023 13230
rect 3233 13227 3299 13230
rect 3049 13154 3115 13157
rect 3325 13154 3391 13157
rect 3049 13152 3391 13154
rect 3049 13096 3054 13152
rect 3110 13096 3330 13152
rect 3386 13096 3391 13152
rect 3049 13094 3391 13096
rect 3049 13091 3115 13094
rect 3325 13091 3391 13094
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 10058 13088 10374 13089
rect 10058 13024 10064 13088
rect 10128 13024 10144 13088
rect 10208 13024 10224 13088
rect 10288 13024 10304 13088
rect 10368 13024 10374 13088
rect 10058 13023 10374 13024
rect 8150 12956 8156 13020
rect 8220 13018 8226 13020
rect 9121 13018 9187 13021
rect 8220 13016 9187 13018
rect 8220 12960 9126 13016
rect 9182 12960 9187 13016
rect 8220 12958 9187 12960
rect 8220 12956 8226 12958
rect 9121 12955 9187 12958
rect 2078 12820 2084 12884
rect 2148 12882 2154 12884
rect 2589 12882 2655 12885
rect 2148 12880 2655 12882
rect 2148 12824 2594 12880
rect 2650 12824 2655 12880
rect 2148 12822 2655 12824
rect 2148 12820 2154 12822
rect 2589 12819 2655 12822
rect 6361 12882 6427 12885
rect 7230 12882 7236 12884
rect 6361 12880 7236 12882
rect 6361 12824 6366 12880
rect 6422 12824 7236 12880
rect 6361 12822 7236 12824
rect 6361 12819 6427 12822
rect 7230 12820 7236 12822
rect 7300 12882 7306 12884
rect 7833 12882 7899 12885
rect 7300 12880 7899 12882
rect 7300 12824 7838 12880
rect 7894 12824 7899 12880
rect 7300 12822 7899 12824
rect 7300 12820 7306 12822
rect 7833 12819 7899 12822
rect 0 12610 400 12640
rect 1209 12610 1275 12613
rect 0 12608 1275 12610
rect 0 12552 1214 12608
rect 1270 12552 1275 12608
rect 0 12550 1275 12552
rect 0 12520 400 12550
rect 1209 12547 1275 12550
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 10718 12544 11034 12545
rect 10718 12480 10724 12544
rect 10788 12480 10804 12544
rect 10868 12480 10884 12544
rect 10948 12480 10964 12544
rect 11028 12480 11034 12544
rect 10718 12479 11034 12480
rect 1853 12474 1919 12477
rect 2681 12474 2747 12477
rect 5073 12474 5139 12477
rect 1853 12472 2747 12474
rect 1853 12416 1858 12472
rect 1914 12416 2686 12472
rect 2742 12416 2747 12472
rect 1853 12414 2747 12416
rect 1853 12411 1919 12414
rect 2681 12411 2747 12414
rect 5030 12472 5139 12474
rect 5030 12416 5078 12472
rect 5134 12416 5139 12472
rect 5030 12411 5139 12416
rect 0 12338 400 12368
rect 749 12338 815 12341
rect 0 12336 815 12338
rect 0 12280 754 12336
rect 810 12280 815 12336
rect 0 12278 815 12280
rect 0 12248 400 12278
rect 749 12275 815 12278
rect 2221 12338 2287 12341
rect 2446 12338 2452 12340
rect 2221 12336 2452 12338
rect 2221 12280 2226 12336
rect 2282 12280 2452 12336
rect 2221 12278 2452 12280
rect 2221 12275 2287 12278
rect 2446 12276 2452 12278
rect 2516 12276 2522 12340
rect 2681 12338 2747 12341
rect 5030 12338 5090 12411
rect 2681 12336 5090 12338
rect 2681 12280 2686 12336
rect 2742 12280 5090 12336
rect 2681 12278 5090 12280
rect 2681 12275 2747 12278
rect 3693 12202 3759 12205
rect 3190 12200 3759 12202
rect 3190 12144 3698 12200
rect 3754 12144 3759 12200
rect 3190 12142 3759 12144
rect 0 12066 400 12096
rect 565 12066 631 12069
rect 0 12064 631 12066
rect 0 12008 570 12064
rect 626 12008 631 12064
rect 0 12006 631 12008
rect 0 11976 400 12006
rect 565 12003 631 12006
rect 1158 12004 1164 12068
rect 1228 12066 1234 12068
rect 1577 12066 1643 12069
rect 1945 12068 2011 12069
rect 1894 12066 1900 12068
rect 1228 12064 1643 12066
rect 1228 12008 1582 12064
rect 1638 12008 1643 12064
rect 1228 12006 1643 12008
rect 1854 12006 1900 12066
rect 1964 12064 2011 12068
rect 2006 12008 2011 12064
rect 1228 12004 1234 12006
rect 1577 12003 1643 12006
rect 1894 12004 1900 12006
rect 1964 12004 2011 12008
rect 1945 12003 2011 12004
rect 2957 12066 3023 12069
rect 3190 12066 3250 12142
rect 3693 12139 3759 12142
rect 4102 12140 4108 12204
rect 4172 12202 4178 12204
rect 4705 12202 4771 12205
rect 8477 12204 8543 12205
rect 8477 12202 8524 12204
rect 4172 12200 4771 12202
rect 4172 12144 4710 12200
rect 4766 12144 4771 12200
rect 4172 12142 4771 12144
rect 8432 12200 8524 12202
rect 8432 12144 8482 12200
rect 8432 12142 8524 12144
rect 4172 12140 4178 12142
rect 4705 12139 4771 12142
rect 8477 12140 8524 12142
rect 8588 12140 8594 12204
rect 8477 12139 8543 12140
rect 2957 12064 3250 12066
rect 2957 12008 2962 12064
rect 3018 12008 3250 12064
rect 2957 12006 3250 12008
rect 8293 12066 8359 12069
rect 8293 12064 8402 12066
rect 8293 12008 8298 12064
rect 8354 12008 8402 12064
rect 2957 12003 3023 12006
rect 8293 12003 8402 12008
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 0 11794 400 11824
rect 8342 11797 8402 12003
rect 10058 12000 10374 12001
rect 10058 11936 10064 12000
rect 10128 11936 10144 12000
rect 10208 11936 10224 12000
rect 10288 11936 10304 12000
rect 10368 11936 10374 12000
rect 10058 11935 10374 11936
rect 2773 11796 2839 11797
rect 974 11794 980 11796
rect 0 11734 980 11794
rect 0 11704 400 11734
rect 974 11732 980 11734
rect 1044 11732 1050 11796
rect 2773 11794 2820 11796
rect 2728 11792 2820 11794
rect 2728 11736 2778 11792
rect 2728 11734 2820 11736
rect 2773 11732 2820 11734
rect 2884 11732 2890 11796
rect 8293 11792 8402 11797
rect 8293 11736 8298 11792
rect 8354 11736 8402 11792
rect 8293 11734 8402 11736
rect 8477 11794 8543 11797
rect 8845 11794 8911 11797
rect 8477 11792 8911 11794
rect 8477 11736 8482 11792
rect 8538 11736 8850 11792
rect 8906 11736 8911 11792
rect 8477 11734 8911 11736
rect 2773 11731 2839 11732
rect 8293 11731 8359 11734
rect 8477 11731 8543 11734
rect 8845 11731 8911 11734
rect 8385 11658 8451 11661
rect 8518 11658 8524 11660
rect 8385 11656 8524 11658
rect 8385 11600 8390 11656
rect 8446 11600 8524 11656
rect 8385 11598 8524 11600
rect 8385 11595 8451 11598
rect 8518 11596 8524 11598
rect 8588 11596 8594 11660
rect 0 11522 400 11552
rect 1485 11522 1551 11525
rect 0 11520 1551 11522
rect 0 11464 1490 11520
rect 1546 11464 1551 11520
rect 0 11462 1551 11464
rect 0 11432 400 11462
rect 1485 11459 1551 11462
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 10718 11456 11034 11457
rect 10718 11392 10724 11456
rect 10788 11392 10804 11456
rect 10868 11392 10884 11456
rect 10948 11392 10964 11456
rect 11028 11392 11034 11456
rect 10718 11391 11034 11392
rect 0 11250 400 11280
rect 1393 11250 1459 11253
rect 0 11248 1459 11250
rect 0 11192 1398 11248
rect 1454 11192 1459 11248
rect 0 11190 1459 11192
rect 0 11160 400 11190
rect 1393 11187 1459 11190
rect 0 10978 400 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 400 10918
rect 1577 10915 1643 10918
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 10058 10912 10374 10913
rect 10058 10848 10064 10912
rect 10128 10848 10144 10912
rect 10208 10848 10224 10912
rect 10288 10848 10304 10912
rect 10368 10848 10374 10912
rect 10058 10847 10374 10848
rect 5625 10570 5691 10573
rect 6545 10570 6611 10573
rect 5625 10568 6611 10570
rect 5625 10512 5630 10568
rect 5686 10512 6550 10568
rect 6606 10512 6611 10568
rect 5625 10510 6611 10512
rect 5625 10507 5691 10510
rect 6545 10507 6611 10510
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 10718 10368 11034 10369
rect 10718 10304 10724 10368
rect 10788 10304 10804 10368
rect 10868 10304 10884 10368
rect 10948 10304 10964 10368
rect 11028 10304 11034 10368
rect 10718 10303 11034 10304
rect 2865 10162 2931 10165
rect 3877 10162 3943 10165
rect 4102 10162 4108 10164
rect 2865 10160 4108 10162
rect 2865 10104 2870 10160
rect 2926 10104 3882 10160
rect 3938 10104 4108 10160
rect 2865 10102 4108 10104
rect 2865 10099 2931 10102
rect 3877 10099 3943 10102
rect 4102 10100 4108 10102
rect 4172 10162 4178 10164
rect 4797 10162 4863 10165
rect 4172 10160 4863 10162
rect 4172 10104 4802 10160
rect 4858 10104 4863 10160
rect 4172 10102 4863 10104
rect 4172 10100 4178 10102
rect 4797 10099 4863 10102
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 10058 9824 10374 9825
rect 10058 9760 10064 9824
rect 10128 9760 10144 9824
rect 10208 9760 10224 9824
rect 10288 9760 10304 9824
rect 10368 9760 10374 9824
rect 10058 9759 10374 9760
rect 9213 9482 9279 9485
rect 11278 9482 11284 9484
rect 9213 9480 11284 9482
rect 9213 9424 9218 9480
rect 9274 9424 11284 9480
rect 9213 9422 11284 9424
rect 9213 9419 9279 9422
rect 11278 9420 11284 9422
rect 11348 9420 11354 9484
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 10718 9280 11034 9281
rect 10718 9216 10724 9280
rect 10788 9216 10804 9280
rect 10868 9216 10884 9280
rect 10948 9216 10964 9280
rect 11028 9216 11034 9280
rect 10718 9215 11034 9216
rect 1945 9074 2011 9077
rect 2078 9074 2084 9076
rect 1945 9072 2084 9074
rect 1945 9016 1950 9072
rect 2006 9016 2084 9072
rect 1945 9014 2084 9016
rect 1945 9011 2011 9014
rect 2078 9012 2084 9014
rect 2148 9012 2154 9076
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 10058 8736 10374 8737
rect 10058 8672 10064 8736
rect 10128 8672 10144 8736
rect 10208 8672 10224 8736
rect 10288 8672 10304 8736
rect 10368 8672 10374 8736
rect 10058 8671 10374 8672
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 10718 8192 11034 8193
rect 10718 8128 10724 8192
rect 10788 8128 10804 8192
rect 10868 8128 10884 8192
rect 10948 8128 10964 8192
rect 11028 8128 11034 8192
rect 10718 8127 11034 8128
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 10058 7648 10374 7649
rect 10058 7584 10064 7648
rect 10128 7584 10144 7648
rect 10208 7584 10224 7648
rect 10288 7584 10304 7648
rect 10368 7584 10374 7648
rect 10058 7583 10374 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 10718 7104 11034 7105
rect 10718 7040 10724 7104
rect 10788 7040 10804 7104
rect 10868 7040 10884 7104
rect 10948 7040 10964 7104
rect 11028 7040 11034 7104
rect 10718 7039 11034 7040
rect 6913 6762 6979 6765
rect 7046 6762 7052 6764
rect 6913 6760 7052 6762
rect 6913 6704 6918 6760
rect 6974 6704 7052 6760
rect 6913 6702 7052 6704
rect 6913 6699 6979 6702
rect 7046 6700 7052 6702
rect 7116 6700 7122 6764
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 10058 6560 10374 6561
rect 10058 6496 10064 6560
rect 10128 6496 10144 6560
rect 10208 6496 10224 6560
rect 10288 6496 10304 6560
rect 10368 6496 10374 6560
rect 10058 6495 10374 6496
rect 3141 6354 3207 6357
rect 3785 6354 3851 6357
rect 3141 6352 3851 6354
rect 3141 6296 3146 6352
rect 3202 6296 3790 6352
rect 3846 6296 3851 6352
rect 3141 6294 3851 6296
rect 3141 6291 3207 6294
rect 3785 6291 3851 6294
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 10718 6016 11034 6017
rect 10718 5952 10724 6016
rect 10788 5952 10804 6016
rect 10868 5952 10884 6016
rect 10948 5952 10964 6016
rect 11028 5952 11034 6016
rect 10718 5951 11034 5952
rect 0 5538 400 5568
rect 657 5538 723 5541
rect 0 5536 723 5538
rect 0 5480 662 5536
rect 718 5480 723 5536
rect 0 5478 723 5480
rect 0 5448 400 5478
rect 657 5475 723 5478
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 10058 5472 10374 5473
rect 10058 5408 10064 5472
rect 10128 5408 10144 5472
rect 10208 5408 10224 5472
rect 10288 5408 10304 5472
rect 10368 5408 10374 5472
rect 10058 5407 10374 5408
rect 0 5269 400 5296
rect 0 5264 447 5269
rect 0 5208 386 5264
rect 442 5208 447 5264
rect 0 5203 447 5208
rect 0 5176 400 5203
rect 0 4997 400 5024
rect 0 4992 447 4997
rect 0 4936 386 4992
rect 442 4936 447 4992
rect 0 4931 447 4936
rect 0 4904 400 4931
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 10718 4928 11034 4929
rect 10718 4864 10724 4928
rect 10788 4864 10804 4928
rect 10868 4864 10884 4928
rect 10948 4864 10964 4928
rect 11028 4864 11034 4928
rect 10718 4863 11034 4864
rect 0 4722 400 4752
rect 606 4722 612 4724
rect 0 4662 612 4722
rect 0 4632 400 4662
rect 606 4660 612 4662
rect 676 4660 682 4724
rect 54 4388 60 4452
rect 124 4450 130 4452
rect 381 4450 447 4453
rect 124 4448 447 4450
rect 124 4392 386 4448
rect 442 4392 447 4448
rect 124 4390 447 4392
rect 124 4388 130 4390
rect 381 4387 447 4390
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 10058 4384 10374 4385
rect 10058 4320 10064 4384
rect 10128 4320 10144 4384
rect 10208 4320 10224 4384
rect 10288 4320 10304 4384
rect 10368 4320 10374 4384
rect 10058 4319 10374 4320
rect 6862 3980 6868 4044
rect 6932 4042 6938 4044
rect 8017 4042 8083 4045
rect 8937 4044 9003 4045
rect 6932 4040 8083 4042
rect 6932 3984 8022 4040
rect 8078 3984 8083 4040
rect 6932 3982 8083 3984
rect 6932 3980 6938 3982
rect 8017 3979 8083 3982
rect 8886 3980 8892 4044
rect 8956 4042 9003 4044
rect 8956 4040 9048 4042
rect 8998 3984 9048 4040
rect 8956 3982 9048 3984
rect 8956 3980 9003 3982
rect 8937 3979 9003 3980
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 10718 3840 11034 3841
rect 10718 3776 10724 3840
rect 10788 3776 10804 3840
rect 10868 3776 10884 3840
rect 10948 3776 10964 3840
rect 11028 3776 11034 3840
rect 10718 3775 11034 3776
rect 9121 3772 9187 3773
rect 9070 3708 9076 3772
rect 9140 3770 9187 3772
rect 9140 3768 9232 3770
rect 9182 3712 9232 3768
rect 9140 3710 9232 3712
rect 9140 3708 9187 3710
rect 9121 3707 9187 3708
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 10058 3296 10374 3297
rect 10058 3232 10064 3296
rect 10128 3232 10144 3296
rect 10208 3232 10224 3296
rect 10288 3232 10304 3296
rect 10368 3232 10374 3296
rect 10058 3231 10374 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 10718 2752 11034 2753
rect 10718 2688 10724 2752
rect 10788 2688 10804 2752
rect 10868 2688 10884 2752
rect 10948 2688 10964 2752
rect 11028 2688 11034 2752
rect 10718 2687 11034 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 10058 2208 10374 2209
rect 10058 2144 10064 2208
rect 10128 2144 10144 2208
rect 10208 2144 10224 2208
rect 10288 2144 10304 2208
rect 10368 2144 10374 2208
rect 10058 2143 10374 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 10718 1664 11034 1665
rect 10718 1600 10724 1664
rect 10788 1600 10804 1664
rect 10868 1600 10884 1664
rect 10948 1600 10964 1664
rect 11028 1600 11034 1664
rect 10718 1599 11034 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 10058 1120 10374 1121
rect 10058 1056 10064 1120
rect 10128 1056 10144 1120
rect 10208 1056 10224 1120
rect 10288 1056 10304 1120
rect 10368 1056 10374 1120
rect 10058 1055 10374 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
rect 10718 576 11034 577
rect 10718 512 10724 576
rect 10788 512 10804 576
rect 10868 512 10884 576
rect 10948 512 10964 576
rect 11028 512 11034 576
rect 10718 511 11034 512
<< via3 >>
rect 980 43556 1044 43620
rect 7788 43616 7852 43620
rect 7788 43560 7802 43616
rect 7802 43560 7852 43616
rect 7788 43556 7852 43560
rect 4324 43004 4388 43008
rect 4324 42948 4328 43004
rect 4328 42948 4384 43004
rect 4384 42948 4388 43004
rect 4324 42944 4388 42948
rect 4404 43004 4468 43008
rect 4404 42948 4408 43004
rect 4408 42948 4464 43004
rect 4464 42948 4468 43004
rect 4404 42944 4468 42948
rect 4484 43004 4548 43008
rect 4484 42948 4488 43004
rect 4488 42948 4544 43004
rect 4544 42948 4548 43004
rect 4484 42944 4548 42948
rect 4564 43004 4628 43008
rect 4564 42948 4568 43004
rect 4568 42948 4624 43004
rect 4624 42948 4628 43004
rect 4564 42944 4628 42948
rect 10724 43004 10788 43008
rect 10724 42948 10728 43004
rect 10728 42948 10784 43004
rect 10784 42948 10788 43004
rect 10724 42944 10788 42948
rect 10804 43004 10868 43008
rect 10804 42948 10808 43004
rect 10808 42948 10864 43004
rect 10864 42948 10868 43004
rect 10804 42944 10868 42948
rect 10884 43004 10948 43008
rect 10884 42948 10888 43004
rect 10888 42948 10944 43004
rect 10944 42948 10948 43004
rect 10884 42944 10948 42948
rect 10964 43004 11028 43008
rect 10964 42948 10968 43004
rect 10968 42948 11024 43004
rect 11024 42948 11028 43004
rect 10964 42944 11028 42948
rect 3664 42460 3728 42464
rect 3664 42404 3668 42460
rect 3668 42404 3724 42460
rect 3724 42404 3728 42460
rect 3664 42400 3728 42404
rect 3744 42460 3808 42464
rect 3744 42404 3748 42460
rect 3748 42404 3804 42460
rect 3804 42404 3808 42460
rect 3744 42400 3808 42404
rect 3824 42460 3888 42464
rect 3824 42404 3828 42460
rect 3828 42404 3884 42460
rect 3884 42404 3888 42460
rect 3824 42400 3888 42404
rect 3904 42460 3968 42464
rect 3904 42404 3908 42460
rect 3908 42404 3964 42460
rect 3964 42404 3968 42460
rect 3904 42400 3968 42404
rect 10064 42460 10128 42464
rect 10064 42404 10068 42460
rect 10068 42404 10124 42460
rect 10124 42404 10128 42460
rect 10064 42400 10128 42404
rect 10144 42460 10208 42464
rect 10144 42404 10148 42460
rect 10148 42404 10204 42460
rect 10204 42404 10208 42460
rect 10144 42400 10208 42404
rect 10224 42460 10288 42464
rect 10224 42404 10228 42460
rect 10228 42404 10284 42460
rect 10284 42404 10288 42460
rect 10224 42400 10288 42404
rect 10304 42460 10368 42464
rect 10304 42404 10308 42460
rect 10308 42404 10364 42460
rect 10364 42404 10368 42460
rect 10304 42400 10368 42404
rect 5580 42196 5644 42260
rect 5212 42060 5276 42124
rect 4324 41916 4388 41920
rect 4324 41860 4328 41916
rect 4328 41860 4384 41916
rect 4384 41860 4388 41916
rect 4324 41856 4388 41860
rect 4404 41916 4468 41920
rect 4404 41860 4408 41916
rect 4408 41860 4464 41916
rect 4464 41860 4468 41916
rect 4404 41856 4468 41860
rect 4484 41916 4548 41920
rect 4484 41860 4488 41916
rect 4488 41860 4544 41916
rect 4544 41860 4548 41916
rect 4484 41856 4548 41860
rect 4564 41916 4628 41920
rect 4564 41860 4568 41916
rect 4568 41860 4624 41916
rect 4624 41860 4628 41916
rect 4564 41856 4628 41860
rect 10724 41916 10788 41920
rect 10724 41860 10728 41916
rect 10728 41860 10784 41916
rect 10784 41860 10788 41916
rect 10724 41856 10788 41860
rect 10804 41916 10868 41920
rect 10804 41860 10808 41916
rect 10808 41860 10864 41916
rect 10864 41860 10868 41916
rect 10804 41856 10868 41860
rect 10884 41916 10948 41920
rect 10884 41860 10888 41916
rect 10888 41860 10944 41916
rect 10944 41860 10948 41916
rect 10884 41856 10948 41860
rect 10964 41916 11028 41920
rect 10964 41860 10968 41916
rect 10968 41860 11024 41916
rect 11024 41860 11028 41916
rect 10964 41856 11028 41860
rect 6684 41712 6748 41716
rect 6684 41656 6698 41712
rect 6698 41656 6748 41712
rect 6684 41652 6748 41656
rect 1164 41576 1228 41580
rect 1164 41520 1178 41576
rect 1178 41520 1228 41576
rect 1164 41516 1228 41520
rect 7972 41380 8036 41444
rect 3664 41372 3728 41376
rect 3664 41316 3668 41372
rect 3668 41316 3724 41372
rect 3724 41316 3728 41372
rect 3664 41312 3728 41316
rect 3744 41372 3808 41376
rect 3744 41316 3748 41372
rect 3748 41316 3804 41372
rect 3804 41316 3808 41372
rect 3744 41312 3808 41316
rect 3824 41372 3888 41376
rect 3824 41316 3828 41372
rect 3828 41316 3884 41372
rect 3884 41316 3888 41372
rect 3824 41312 3888 41316
rect 3904 41372 3968 41376
rect 3904 41316 3908 41372
rect 3908 41316 3964 41372
rect 3964 41316 3968 41372
rect 3904 41312 3968 41316
rect 10064 41372 10128 41376
rect 10064 41316 10068 41372
rect 10068 41316 10124 41372
rect 10124 41316 10128 41372
rect 10064 41312 10128 41316
rect 10144 41372 10208 41376
rect 10144 41316 10148 41372
rect 10148 41316 10204 41372
rect 10204 41316 10208 41372
rect 10144 41312 10208 41316
rect 10224 41372 10288 41376
rect 10224 41316 10228 41372
rect 10228 41316 10284 41372
rect 10284 41316 10288 41372
rect 10224 41312 10288 41316
rect 10304 41372 10368 41376
rect 10304 41316 10308 41372
rect 10308 41316 10364 41372
rect 10364 41316 10368 41372
rect 10304 41312 10368 41316
rect 2636 41108 2700 41172
rect 3372 40972 3436 41036
rect 4324 40828 4388 40832
rect 4324 40772 4328 40828
rect 4328 40772 4384 40828
rect 4384 40772 4388 40828
rect 4324 40768 4388 40772
rect 4404 40828 4468 40832
rect 4404 40772 4408 40828
rect 4408 40772 4464 40828
rect 4464 40772 4468 40828
rect 4404 40768 4468 40772
rect 4484 40828 4548 40832
rect 4484 40772 4488 40828
rect 4488 40772 4544 40828
rect 4544 40772 4548 40828
rect 4484 40768 4548 40772
rect 4564 40828 4628 40832
rect 4564 40772 4568 40828
rect 4568 40772 4624 40828
rect 4624 40772 4628 40828
rect 4564 40768 4628 40772
rect 10724 40828 10788 40832
rect 10724 40772 10728 40828
rect 10728 40772 10784 40828
rect 10784 40772 10788 40828
rect 10724 40768 10788 40772
rect 10804 40828 10868 40832
rect 10804 40772 10808 40828
rect 10808 40772 10864 40828
rect 10864 40772 10868 40828
rect 10804 40768 10868 40772
rect 10884 40828 10948 40832
rect 10884 40772 10888 40828
rect 10888 40772 10944 40828
rect 10944 40772 10948 40828
rect 10884 40768 10948 40772
rect 10964 40828 11028 40832
rect 10964 40772 10968 40828
rect 10968 40772 11024 40828
rect 11024 40772 11028 40828
rect 10964 40768 11028 40772
rect 3664 40284 3728 40288
rect 3664 40228 3668 40284
rect 3668 40228 3724 40284
rect 3724 40228 3728 40284
rect 3664 40224 3728 40228
rect 3744 40284 3808 40288
rect 3744 40228 3748 40284
rect 3748 40228 3804 40284
rect 3804 40228 3808 40284
rect 3744 40224 3808 40228
rect 3824 40284 3888 40288
rect 3824 40228 3828 40284
rect 3828 40228 3884 40284
rect 3884 40228 3888 40284
rect 3824 40224 3888 40228
rect 3904 40284 3968 40288
rect 3904 40228 3908 40284
rect 3908 40228 3964 40284
rect 3964 40228 3968 40284
rect 3904 40224 3968 40228
rect 10064 40284 10128 40288
rect 10064 40228 10068 40284
rect 10068 40228 10124 40284
rect 10124 40228 10128 40284
rect 10064 40224 10128 40228
rect 10144 40284 10208 40288
rect 10144 40228 10148 40284
rect 10148 40228 10204 40284
rect 10204 40228 10208 40284
rect 10144 40224 10208 40228
rect 10224 40284 10288 40288
rect 10224 40228 10228 40284
rect 10228 40228 10284 40284
rect 10284 40228 10288 40284
rect 10224 40224 10288 40228
rect 10304 40284 10368 40288
rect 10304 40228 10308 40284
rect 10308 40228 10364 40284
rect 10364 40228 10368 40284
rect 10304 40224 10368 40228
rect 1900 40156 1964 40220
rect 4844 40156 4908 40220
rect 4108 40020 4172 40084
rect 5948 40020 6012 40084
rect 6500 40020 6564 40084
rect 2084 39884 2148 39948
rect 4324 39740 4388 39744
rect 4324 39684 4328 39740
rect 4328 39684 4384 39740
rect 4384 39684 4388 39740
rect 4324 39680 4388 39684
rect 4404 39740 4468 39744
rect 4404 39684 4408 39740
rect 4408 39684 4464 39740
rect 4464 39684 4468 39740
rect 4404 39680 4468 39684
rect 4484 39740 4548 39744
rect 4484 39684 4488 39740
rect 4488 39684 4544 39740
rect 4544 39684 4548 39740
rect 4484 39680 4548 39684
rect 4564 39740 4628 39744
rect 4564 39684 4568 39740
rect 4568 39684 4624 39740
rect 4624 39684 4628 39740
rect 4564 39680 4628 39684
rect 10724 39740 10788 39744
rect 10724 39684 10728 39740
rect 10728 39684 10784 39740
rect 10784 39684 10788 39740
rect 10724 39680 10788 39684
rect 10804 39740 10868 39744
rect 10804 39684 10808 39740
rect 10808 39684 10864 39740
rect 10864 39684 10868 39740
rect 10804 39680 10868 39684
rect 10884 39740 10948 39744
rect 10884 39684 10888 39740
rect 10888 39684 10944 39740
rect 10944 39684 10948 39740
rect 10884 39680 10948 39684
rect 10964 39740 11028 39744
rect 10964 39684 10968 39740
rect 10968 39684 11024 39740
rect 11024 39684 11028 39740
rect 10964 39680 11028 39684
rect 9444 39612 9508 39676
rect 8340 39476 8404 39540
rect 2084 39340 2148 39404
rect 7604 39340 7668 39404
rect 3664 39196 3728 39200
rect 3664 39140 3668 39196
rect 3668 39140 3724 39196
rect 3724 39140 3728 39196
rect 3664 39136 3728 39140
rect 3744 39196 3808 39200
rect 3744 39140 3748 39196
rect 3748 39140 3804 39196
rect 3804 39140 3808 39196
rect 3744 39136 3808 39140
rect 3824 39196 3888 39200
rect 3824 39140 3828 39196
rect 3828 39140 3884 39196
rect 3884 39140 3888 39196
rect 3824 39136 3888 39140
rect 3904 39196 3968 39200
rect 3904 39140 3908 39196
rect 3908 39140 3964 39196
rect 3964 39140 3968 39196
rect 3904 39136 3968 39140
rect 10064 39196 10128 39200
rect 10064 39140 10068 39196
rect 10068 39140 10124 39196
rect 10124 39140 10128 39196
rect 10064 39136 10128 39140
rect 10144 39196 10208 39200
rect 10144 39140 10148 39196
rect 10148 39140 10204 39196
rect 10204 39140 10208 39196
rect 10144 39136 10208 39140
rect 10224 39196 10288 39200
rect 10224 39140 10228 39196
rect 10228 39140 10284 39196
rect 10284 39140 10288 39196
rect 10224 39136 10288 39140
rect 10304 39196 10368 39200
rect 10304 39140 10308 39196
rect 10308 39140 10364 39196
rect 10364 39140 10368 39196
rect 10304 39136 10368 39140
rect 5028 38660 5092 38724
rect 4324 38652 4388 38656
rect 4324 38596 4328 38652
rect 4328 38596 4384 38652
rect 4384 38596 4388 38652
rect 4324 38592 4388 38596
rect 4404 38652 4468 38656
rect 4404 38596 4408 38652
rect 4408 38596 4464 38652
rect 4464 38596 4468 38652
rect 4404 38592 4468 38596
rect 4484 38652 4548 38656
rect 4484 38596 4488 38652
rect 4488 38596 4544 38652
rect 4544 38596 4548 38652
rect 4484 38592 4548 38596
rect 4564 38652 4628 38656
rect 4564 38596 4568 38652
rect 4568 38596 4624 38652
rect 4624 38596 4628 38652
rect 4564 38592 4628 38596
rect 10724 38652 10788 38656
rect 10724 38596 10728 38652
rect 10728 38596 10784 38652
rect 10784 38596 10788 38652
rect 10724 38592 10788 38596
rect 10804 38652 10868 38656
rect 10804 38596 10808 38652
rect 10808 38596 10864 38652
rect 10864 38596 10868 38652
rect 10804 38592 10868 38596
rect 10884 38652 10948 38656
rect 10884 38596 10888 38652
rect 10888 38596 10944 38652
rect 10944 38596 10948 38652
rect 10884 38592 10948 38596
rect 10964 38652 11028 38656
rect 10964 38596 10968 38652
rect 10968 38596 11024 38652
rect 11024 38596 11028 38652
rect 10964 38592 11028 38596
rect 5580 38388 5644 38452
rect 9076 38448 9140 38452
rect 9076 38392 9126 38448
rect 9126 38392 9140 38448
rect 9076 38388 9140 38392
rect 8524 38312 8588 38316
rect 8524 38256 8538 38312
rect 8538 38256 8588 38312
rect 8524 38252 8588 38256
rect 8708 38312 8772 38316
rect 8708 38256 8758 38312
rect 8758 38256 8772 38312
rect 8708 38252 8772 38256
rect 8156 38116 8220 38180
rect 9260 38116 9324 38180
rect 3664 38108 3728 38112
rect 3664 38052 3668 38108
rect 3668 38052 3724 38108
rect 3724 38052 3728 38108
rect 3664 38048 3728 38052
rect 3744 38108 3808 38112
rect 3744 38052 3748 38108
rect 3748 38052 3804 38108
rect 3804 38052 3808 38108
rect 3744 38048 3808 38052
rect 3824 38108 3888 38112
rect 3824 38052 3828 38108
rect 3828 38052 3884 38108
rect 3884 38052 3888 38108
rect 3824 38048 3888 38052
rect 3904 38108 3968 38112
rect 3904 38052 3908 38108
rect 3908 38052 3964 38108
rect 3964 38052 3968 38108
rect 3904 38048 3968 38052
rect 10064 38108 10128 38112
rect 10064 38052 10068 38108
rect 10068 38052 10124 38108
rect 10124 38052 10128 38108
rect 10064 38048 10128 38052
rect 10144 38108 10208 38112
rect 10144 38052 10148 38108
rect 10148 38052 10204 38108
rect 10204 38052 10208 38108
rect 10144 38048 10208 38052
rect 10224 38108 10288 38112
rect 10224 38052 10228 38108
rect 10228 38052 10284 38108
rect 10284 38052 10288 38108
rect 10224 38048 10288 38052
rect 10304 38108 10368 38112
rect 10304 38052 10308 38108
rect 10308 38052 10364 38108
rect 10364 38052 10368 38108
rect 10304 38048 10368 38052
rect 8892 37980 8956 38044
rect 3372 37844 3436 37908
rect 4324 37564 4388 37568
rect 4324 37508 4328 37564
rect 4328 37508 4384 37564
rect 4384 37508 4388 37564
rect 4324 37504 4388 37508
rect 4404 37564 4468 37568
rect 4404 37508 4408 37564
rect 4408 37508 4464 37564
rect 4464 37508 4468 37564
rect 4404 37504 4468 37508
rect 4484 37564 4548 37568
rect 4484 37508 4488 37564
rect 4488 37508 4544 37564
rect 4544 37508 4548 37564
rect 4484 37504 4548 37508
rect 4564 37564 4628 37568
rect 4564 37508 4568 37564
rect 4568 37508 4624 37564
rect 4624 37508 4628 37564
rect 4564 37504 4628 37508
rect 10724 37564 10788 37568
rect 10724 37508 10728 37564
rect 10728 37508 10784 37564
rect 10784 37508 10788 37564
rect 10724 37504 10788 37508
rect 10804 37564 10868 37568
rect 10804 37508 10808 37564
rect 10808 37508 10864 37564
rect 10864 37508 10868 37564
rect 10804 37504 10868 37508
rect 10884 37564 10948 37568
rect 10884 37508 10888 37564
rect 10888 37508 10944 37564
rect 10944 37508 10948 37564
rect 10884 37504 10948 37508
rect 10964 37564 11028 37568
rect 10964 37508 10968 37564
rect 10968 37508 11024 37564
rect 11024 37508 11028 37564
rect 10964 37504 11028 37508
rect 8524 37496 8588 37500
rect 8524 37440 8538 37496
rect 8538 37440 8588 37496
rect 8524 37436 8588 37440
rect 8892 37436 8956 37500
rect 9444 37436 9508 37500
rect 1348 37300 1412 37364
rect 9260 37164 9324 37228
rect 382 37028 446 37092
rect 5580 37028 5644 37092
rect 8524 37028 8588 37092
rect 3664 37020 3728 37024
rect 3664 36964 3668 37020
rect 3668 36964 3724 37020
rect 3724 36964 3728 37020
rect 3664 36960 3728 36964
rect 3744 37020 3808 37024
rect 3744 36964 3748 37020
rect 3748 36964 3804 37020
rect 3804 36964 3808 37020
rect 3744 36960 3808 36964
rect 3824 37020 3888 37024
rect 3824 36964 3828 37020
rect 3828 36964 3884 37020
rect 3884 36964 3888 37020
rect 3824 36960 3888 36964
rect 3904 37020 3968 37024
rect 3904 36964 3908 37020
rect 3908 36964 3964 37020
rect 3964 36964 3968 37020
rect 3904 36960 3968 36964
rect 10064 37020 10128 37024
rect 10064 36964 10068 37020
rect 10068 36964 10124 37020
rect 10124 36964 10128 37020
rect 10064 36960 10128 36964
rect 10144 37020 10208 37024
rect 10144 36964 10148 37020
rect 10148 36964 10204 37020
rect 10204 36964 10208 37020
rect 10144 36960 10208 36964
rect 10224 37020 10288 37024
rect 10224 36964 10228 37020
rect 10228 36964 10284 37020
rect 10284 36964 10288 37020
rect 10224 36960 10288 36964
rect 10304 37020 10368 37024
rect 10304 36964 10308 37020
rect 10308 36964 10364 37020
rect 10364 36964 10368 37020
rect 10304 36960 10368 36964
rect 5396 36816 5460 36820
rect 5396 36760 5446 36816
rect 5446 36760 5460 36816
rect 5396 36756 5460 36760
rect 6132 36756 6196 36820
rect 8340 36756 8404 36820
rect 4324 36476 4388 36480
rect 4324 36420 4328 36476
rect 4328 36420 4384 36476
rect 4384 36420 4388 36476
rect 4324 36416 4388 36420
rect 4404 36476 4468 36480
rect 4404 36420 4408 36476
rect 4408 36420 4464 36476
rect 4464 36420 4468 36476
rect 4404 36416 4468 36420
rect 4484 36476 4548 36480
rect 4484 36420 4488 36476
rect 4488 36420 4544 36476
rect 4544 36420 4548 36476
rect 4484 36416 4548 36420
rect 4564 36476 4628 36480
rect 4564 36420 4568 36476
rect 4568 36420 4624 36476
rect 4624 36420 4628 36476
rect 4564 36416 4628 36420
rect 10724 36476 10788 36480
rect 10724 36420 10728 36476
rect 10728 36420 10784 36476
rect 10784 36420 10788 36476
rect 10724 36416 10788 36420
rect 10804 36476 10868 36480
rect 10804 36420 10808 36476
rect 10808 36420 10864 36476
rect 10864 36420 10868 36476
rect 10804 36416 10868 36420
rect 10884 36476 10948 36480
rect 10884 36420 10888 36476
rect 10888 36420 10944 36476
rect 10944 36420 10948 36476
rect 10884 36416 10948 36420
rect 10964 36476 11028 36480
rect 10964 36420 10968 36476
rect 10968 36420 11024 36476
rect 11024 36420 11028 36476
rect 10964 36416 11028 36420
rect 3188 36348 3252 36412
rect 9076 36348 9140 36412
rect 4844 36076 4908 36140
rect 9076 35940 9140 36004
rect 3664 35932 3728 35936
rect 3664 35876 3668 35932
rect 3668 35876 3724 35932
rect 3724 35876 3728 35932
rect 3664 35872 3728 35876
rect 3744 35932 3808 35936
rect 3744 35876 3748 35932
rect 3748 35876 3804 35932
rect 3804 35876 3808 35932
rect 3744 35872 3808 35876
rect 3824 35932 3888 35936
rect 3824 35876 3828 35932
rect 3828 35876 3884 35932
rect 3884 35876 3888 35932
rect 3824 35872 3888 35876
rect 3904 35932 3968 35936
rect 3904 35876 3908 35932
rect 3908 35876 3964 35932
rect 3964 35876 3968 35932
rect 3904 35872 3968 35876
rect 10064 35932 10128 35936
rect 10064 35876 10068 35932
rect 10068 35876 10124 35932
rect 10124 35876 10128 35932
rect 10064 35872 10128 35876
rect 10144 35932 10208 35936
rect 10144 35876 10148 35932
rect 10148 35876 10204 35932
rect 10204 35876 10208 35932
rect 10144 35872 10208 35876
rect 10224 35932 10288 35936
rect 10224 35876 10228 35932
rect 10228 35876 10284 35932
rect 10284 35876 10288 35932
rect 10224 35872 10288 35876
rect 10304 35932 10368 35936
rect 10304 35876 10308 35932
rect 10308 35876 10364 35932
rect 10364 35876 10368 35932
rect 10304 35872 10368 35876
rect 8156 35668 8220 35732
rect 7052 35532 7116 35596
rect 4324 35388 4388 35392
rect 4324 35332 4328 35388
rect 4328 35332 4384 35388
rect 4384 35332 4388 35388
rect 4324 35328 4388 35332
rect 4404 35388 4468 35392
rect 4404 35332 4408 35388
rect 4408 35332 4464 35388
rect 4464 35332 4468 35388
rect 4404 35328 4468 35332
rect 4484 35388 4548 35392
rect 4484 35332 4488 35388
rect 4488 35332 4544 35388
rect 4544 35332 4548 35388
rect 4484 35328 4548 35332
rect 4564 35388 4628 35392
rect 4564 35332 4568 35388
rect 4568 35332 4624 35388
rect 4624 35332 4628 35388
rect 4564 35328 4628 35332
rect 10724 35388 10788 35392
rect 10724 35332 10728 35388
rect 10728 35332 10784 35388
rect 10784 35332 10788 35388
rect 10724 35328 10788 35332
rect 10804 35388 10868 35392
rect 10804 35332 10808 35388
rect 10808 35332 10864 35388
rect 10864 35332 10868 35388
rect 10804 35328 10868 35332
rect 10884 35388 10948 35392
rect 10884 35332 10888 35388
rect 10888 35332 10944 35388
rect 10944 35332 10948 35388
rect 10884 35328 10948 35332
rect 10964 35388 11028 35392
rect 10964 35332 10968 35388
rect 10968 35332 11024 35388
rect 11024 35332 11028 35388
rect 10964 35328 11028 35332
rect 428 35124 492 35188
rect 1900 35184 1964 35188
rect 1900 35128 1914 35184
rect 1914 35128 1964 35184
rect 1900 35124 1964 35128
rect 9260 35124 9324 35188
rect 980 34988 1044 35052
rect 5396 34988 5460 35052
rect 2452 34852 2516 34916
rect 7788 34852 7852 34916
rect 3664 34844 3728 34848
rect 3664 34788 3668 34844
rect 3668 34788 3724 34844
rect 3724 34788 3728 34844
rect 3664 34784 3728 34788
rect 3744 34844 3808 34848
rect 3744 34788 3748 34844
rect 3748 34788 3804 34844
rect 3804 34788 3808 34844
rect 3744 34784 3808 34788
rect 3824 34844 3888 34848
rect 3824 34788 3828 34844
rect 3828 34788 3884 34844
rect 3884 34788 3888 34844
rect 3824 34784 3888 34788
rect 3904 34844 3968 34848
rect 3904 34788 3908 34844
rect 3908 34788 3964 34844
rect 3964 34788 3968 34844
rect 3904 34784 3968 34788
rect 10064 34844 10128 34848
rect 10064 34788 10068 34844
rect 10068 34788 10124 34844
rect 10124 34788 10128 34844
rect 10064 34784 10128 34788
rect 10144 34844 10208 34848
rect 10144 34788 10148 34844
rect 10148 34788 10204 34844
rect 10204 34788 10208 34844
rect 10144 34784 10208 34788
rect 10224 34844 10288 34848
rect 10224 34788 10228 34844
rect 10228 34788 10284 34844
rect 10284 34788 10288 34844
rect 10224 34784 10288 34788
rect 10304 34844 10368 34848
rect 10304 34788 10308 34844
rect 10308 34788 10364 34844
rect 10364 34788 10368 34844
rect 10304 34784 10368 34788
rect 1900 34776 1964 34780
rect 1900 34720 1950 34776
rect 1950 34720 1964 34776
rect 1900 34716 1964 34720
rect 4108 34580 4172 34644
rect 4844 34444 4908 34508
rect 5212 34504 5276 34508
rect 5212 34448 5226 34504
rect 5226 34448 5276 34504
rect 5212 34444 5276 34448
rect 8156 34444 8220 34508
rect 8708 34308 8772 34372
rect 4324 34300 4388 34304
rect 4324 34244 4328 34300
rect 4328 34244 4384 34300
rect 4384 34244 4388 34300
rect 4324 34240 4388 34244
rect 4404 34300 4468 34304
rect 4404 34244 4408 34300
rect 4408 34244 4464 34300
rect 4464 34244 4468 34300
rect 4404 34240 4468 34244
rect 4484 34300 4548 34304
rect 4484 34244 4488 34300
rect 4488 34244 4544 34300
rect 4544 34244 4548 34300
rect 4484 34240 4548 34244
rect 4564 34300 4628 34304
rect 4564 34244 4568 34300
rect 4568 34244 4624 34300
rect 4624 34244 4628 34300
rect 4564 34240 4628 34244
rect 10724 34300 10788 34304
rect 10724 34244 10728 34300
rect 10728 34244 10784 34300
rect 10784 34244 10788 34300
rect 10724 34240 10788 34244
rect 10804 34300 10868 34304
rect 10804 34244 10808 34300
rect 10808 34244 10864 34300
rect 10864 34244 10868 34300
rect 10804 34240 10868 34244
rect 10884 34300 10948 34304
rect 10884 34244 10888 34300
rect 10888 34244 10944 34300
rect 10944 34244 10948 34300
rect 10884 34240 10948 34244
rect 10964 34300 11028 34304
rect 10964 34244 10968 34300
rect 10968 34244 11024 34300
rect 11024 34244 11028 34300
rect 10964 34240 11028 34244
rect 3372 34036 3436 34100
rect 5396 34036 5460 34100
rect 7972 34036 8036 34100
rect 10548 33900 10612 33964
rect 3664 33756 3728 33760
rect 3664 33700 3668 33756
rect 3668 33700 3724 33756
rect 3724 33700 3728 33756
rect 3664 33696 3728 33700
rect 3744 33756 3808 33760
rect 3744 33700 3748 33756
rect 3748 33700 3804 33756
rect 3804 33700 3808 33756
rect 3744 33696 3808 33700
rect 3824 33756 3888 33760
rect 3824 33700 3828 33756
rect 3828 33700 3884 33756
rect 3884 33700 3888 33756
rect 3824 33696 3888 33700
rect 3904 33756 3968 33760
rect 3904 33700 3908 33756
rect 3908 33700 3964 33756
rect 3964 33700 3968 33756
rect 3904 33696 3968 33700
rect 10064 33756 10128 33760
rect 10064 33700 10068 33756
rect 10068 33700 10124 33756
rect 10124 33700 10128 33756
rect 10064 33696 10128 33700
rect 10144 33756 10208 33760
rect 10144 33700 10148 33756
rect 10148 33700 10204 33756
rect 10204 33700 10208 33756
rect 10144 33696 10208 33700
rect 10224 33756 10288 33760
rect 10224 33700 10228 33756
rect 10228 33700 10284 33756
rect 10284 33700 10288 33756
rect 10224 33696 10288 33700
rect 10304 33756 10368 33760
rect 10304 33700 10308 33756
rect 10308 33700 10364 33756
rect 10364 33700 10368 33756
rect 10304 33696 10368 33700
rect 9444 33628 9508 33692
rect 7604 33492 7668 33556
rect 8156 33356 8220 33420
rect 1532 33220 1596 33284
rect 3372 33220 3436 33284
rect 4324 33212 4388 33216
rect 4324 33156 4328 33212
rect 4328 33156 4384 33212
rect 4384 33156 4388 33212
rect 4324 33152 4388 33156
rect 4404 33212 4468 33216
rect 4404 33156 4408 33212
rect 4408 33156 4464 33212
rect 4464 33156 4468 33212
rect 4404 33152 4468 33156
rect 4484 33212 4548 33216
rect 4484 33156 4488 33212
rect 4488 33156 4544 33212
rect 4544 33156 4548 33212
rect 4484 33152 4548 33156
rect 4564 33212 4628 33216
rect 4564 33156 4568 33212
rect 4568 33156 4624 33212
rect 4624 33156 4628 33212
rect 4564 33152 4628 33156
rect 2268 33084 2332 33148
rect 6868 33084 6932 33148
rect 7420 33144 7484 33148
rect 10724 33212 10788 33216
rect 10724 33156 10728 33212
rect 10728 33156 10784 33212
rect 10784 33156 10788 33212
rect 10724 33152 10788 33156
rect 10804 33212 10868 33216
rect 10804 33156 10808 33212
rect 10808 33156 10864 33212
rect 10864 33156 10868 33212
rect 10804 33152 10868 33156
rect 10884 33212 10948 33216
rect 10884 33156 10888 33212
rect 10888 33156 10944 33212
rect 10944 33156 10948 33212
rect 10884 33152 10948 33156
rect 10964 33212 11028 33216
rect 10964 33156 10968 33212
rect 10968 33156 11024 33212
rect 11024 33156 11028 33212
rect 10964 33152 11028 33156
rect 7420 33088 7470 33144
rect 7470 33088 7484 33144
rect 7420 33084 7484 33088
rect 980 32948 1044 33012
rect 5764 32676 5828 32740
rect 9076 32676 9140 32740
rect 3664 32668 3728 32672
rect 3664 32612 3668 32668
rect 3668 32612 3724 32668
rect 3724 32612 3728 32668
rect 3664 32608 3728 32612
rect 3744 32668 3808 32672
rect 3744 32612 3748 32668
rect 3748 32612 3804 32668
rect 3804 32612 3808 32668
rect 3744 32608 3808 32612
rect 3824 32668 3888 32672
rect 3824 32612 3828 32668
rect 3828 32612 3884 32668
rect 3884 32612 3888 32668
rect 3824 32608 3888 32612
rect 3904 32668 3968 32672
rect 3904 32612 3908 32668
rect 3908 32612 3964 32668
rect 3964 32612 3968 32668
rect 3904 32608 3968 32612
rect 10064 32668 10128 32672
rect 10064 32612 10068 32668
rect 10068 32612 10124 32668
rect 10124 32612 10128 32668
rect 10064 32608 10128 32612
rect 10144 32668 10208 32672
rect 10144 32612 10148 32668
rect 10148 32612 10204 32668
rect 10204 32612 10208 32668
rect 10144 32608 10208 32612
rect 10224 32668 10288 32672
rect 10224 32612 10228 32668
rect 10228 32612 10284 32668
rect 10284 32612 10288 32668
rect 10224 32608 10288 32612
rect 10304 32668 10368 32672
rect 10304 32612 10308 32668
rect 10308 32612 10364 32668
rect 10364 32612 10368 32668
rect 10304 32608 10368 32612
rect 6132 32600 6196 32604
rect 6132 32544 6182 32600
rect 6182 32544 6196 32600
rect 6132 32540 6196 32544
rect 7972 32600 8036 32604
rect 7972 32544 7986 32600
rect 7986 32544 8036 32600
rect 7972 32540 8036 32544
rect 9076 32540 9140 32604
rect 5580 32404 5644 32468
rect 2268 31920 2332 31924
rect 2268 31864 2318 31920
rect 2318 31864 2332 31920
rect 2268 31860 2332 31864
rect 4324 32124 4388 32128
rect 4324 32068 4328 32124
rect 4328 32068 4384 32124
rect 4384 32068 4388 32124
rect 4324 32064 4388 32068
rect 4404 32124 4468 32128
rect 4404 32068 4408 32124
rect 4408 32068 4464 32124
rect 4464 32068 4468 32124
rect 4404 32064 4468 32068
rect 4484 32124 4548 32128
rect 4484 32068 4488 32124
rect 4488 32068 4544 32124
rect 4544 32068 4548 32124
rect 4484 32064 4548 32068
rect 4564 32124 4628 32128
rect 4564 32068 4568 32124
rect 4568 32068 4624 32124
rect 4624 32068 4628 32124
rect 4564 32064 4628 32068
rect 6868 31996 6932 32060
rect 10724 32124 10788 32128
rect 10724 32068 10728 32124
rect 10728 32068 10784 32124
rect 10784 32068 10788 32124
rect 10724 32064 10788 32068
rect 10804 32124 10868 32128
rect 10804 32068 10808 32124
rect 10808 32068 10864 32124
rect 10864 32068 10868 32124
rect 10804 32064 10868 32068
rect 10884 32124 10948 32128
rect 10884 32068 10888 32124
rect 10888 32068 10944 32124
rect 10944 32068 10948 32124
rect 10884 32064 10948 32068
rect 10964 32124 11028 32128
rect 10964 32068 10968 32124
rect 10968 32068 11024 32124
rect 11024 32068 11028 32124
rect 10964 32064 11028 32068
rect 7788 32056 7852 32060
rect 7788 32000 7802 32056
rect 7802 32000 7852 32056
rect 7788 31996 7852 32000
rect 7972 31996 8036 32060
rect 9076 31996 9140 32060
rect 5212 31724 5276 31788
rect 1716 31648 1780 31652
rect 1716 31592 1766 31648
rect 1766 31592 1780 31648
rect 1716 31588 1780 31592
rect 5764 31588 5828 31652
rect 7420 31724 7484 31788
rect 9076 31648 9140 31652
rect 9076 31592 9126 31648
rect 9126 31592 9140 31648
rect 9076 31588 9140 31592
rect 3664 31580 3728 31584
rect 3664 31524 3668 31580
rect 3668 31524 3724 31580
rect 3724 31524 3728 31580
rect 3664 31520 3728 31524
rect 3744 31580 3808 31584
rect 3744 31524 3748 31580
rect 3748 31524 3804 31580
rect 3804 31524 3808 31580
rect 3744 31520 3808 31524
rect 3824 31580 3888 31584
rect 3824 31524 3828 31580
rect 3828 31524 3884 31580
rect 3884 31524 3888 31580
rect 3824 31520 3888 31524
rect 3904 31580 3968 31584
rect 3904 31524 3908 31580
rect 3908 31524 3964 31580
rect 3964 31524 3968 31580
rect 3904 31520 3968 31524
rect 10064 31580 10128 31584
rect 10064 31524 10068 31580
rect 10068 31524 10124 31580
rect 10124 31524 10128 31580
rect 10064 31520 10128 31524
rect 10144 31580 10208 31584
rect 10144 31524 10148 31580
rect 10148 31524 10204 31580
rect 10204 31524 10208 31580
rect 10144 31520 10208 31524
rect 10224 31580 10288 31584
rect 10224 31524 10228 31580
rect 10228 31524 10284 31580
rect 10284 31524 10288 31580
rect 10224 31520 10288 31524
rect 10304 31580 10368 31584
rect 10304 31524 10308 31580
rect 10308 31524 10364 31580
rect 10364 31524 10368 31580
rect 10304 31520 10368 31524
rect 7788 31452 7852 31516
rect 1532 31316 1596 31380
rect 1716 31104 1780 31108
rect 1716 31048 1766 31104
rect 1766 31048 1780 31104
rect 1716 31044 1780 31048
rect 4324 31036 4388 31040
rect 4324 30980 4328 31036
rect 4328 30980 4384 31036
rect 4384 30980 4388 31036
rect 4324 30976 4388 30980
rect 4404 31036 4468 31040
rect 4404 30980 4408 31036
rect 4408 30980 4464 31036
rect 4464 30980 4468 31036
rect 4404 30976 4468 30980
rect 4484 31036 4548 31040
rect 4484 30980 4488 31036
rect 4488 30980 4544 31036
rect 4544 30980 4548 31036
rect 4484 30976 4548 30980
rect 4564 31036 4628 31040
rect 4564 30980 4568 31036
rect 4568 30980 4624 31036
rect 4624 30980 4628 31036
rect 4564 30976 4628 30980
rect 5580 30908 5644 30972
rect 10724 31036 10788 31040
rect 10724 30980 10728 31036
rect 10728 30980 10784 31036
rect 10784 30980 10788 31036
rect 10724 30976 10788 30980
rect 10804 31036 10868 31040
rect 10804 30980 10808 31036
rect 10808 30980 10864 31036
rect 10864 30980 10868 31036
rect 10804 30976 10868 30980
rect 10884 31036 10948 31040
rect 10884 30980 10888 31036
rect 10888 30980 10944 31036
rect 10944 30980 10948 31036
rect 10884 30976 10948 30980
rect 10964 31036 11028 31040
rect 10964 30980 10968 31036
rect 10968 30980 11024 31036
rect 11024 30980 11028 31036
rect 10964 30976 11028 30980
rect 5580 30772 5644 30836
rect 6500 30772 6564 30836
rect 7420 30772 7484 30836
rect 9628 30636 9692 30700
rect 5764 30500 5828 30564
rect 6500 30560 6564 30564
rect 6500 30504 6550 30560
rect 6550 30504 6564 30560
rect 6500 30500 6564 30504
rect 9812 30500 9876 30564
rect 3664 30492 3728 30496
rect 3664 30436 3668 30492
rect 3668 30436 3724 30492
rect 3724 30436 3728 30492
rect 3664 30432 3728 30436
rect 3744 30492 3808 30496
rect 3744 30436 3748 30492
rect 3748 30436 3804 30492
rect 3804 30436 3808 30492
rect 3744 30432 3808 30436
rect 3824 30492 3888 30496
rect 3824 30436 3828 30492
rect 3828 30436 3884 30492
rect 3884 30436 3888 30492
rect 3824 30432 3888 30436
rect 3904 30492 3968 30496
rect 3904 30436 3908 30492
rect 3908 30436 3964 30492
rect 3964 30436 3968 30492
rect 3904 30432 3968 30436
rect 10064 30492 10128 30496
rect 10064 30436 10068 30492
rect 10068 30436 10124 30492
rect 10124 30436 10128 30492
rect 10064 30432 10128 30436
rect 10144 30492 10208 30496
rect 10144 30436 10148 30492
rect 10148 30436 10204 30492
rect 10204 30436 10208 30492
rect 10144 30432 10208 30436
rect 10224 30492 10288 30496
rect 10224 30436 10228 30492
rect 10228 30436 10284 30492
rect 10284 30436 10288 30492
rect 10224 30432 10288 30436
rect 10304 30492 10368 30496
rect 10304 30436 10308 30492
rect 10308 30436 10364 30492
rect 10364 30436 10368 30492
rect 10304 30432 10368 30436
rect 612 30364 676 30428
rect 1348 30364 1412 30428
rect 4108 30364 4172 30428
rect 6684 30364 6748 30428
rect 2084 30228 2148 30292
rect 2636 30228 2700 30292
rect 5948 30228 6012 30292
rect 7236 30288 7300 30292
rect 7236 30232 7250 30288
rect 7250 30232 7300 30288
rect 7236 30228 7300 30232
rect 9260 30228 9324 30292
rect 5764 30092 5828 30156
rect 7052 29956 7116 30020
rect 4324 29948 4388 29952
rect 4324 29892 4328 29948
rect 4328 29892 4384 29948
rect 4384 29892 4388 29948
rect 4324 29888 4388 29892
rect 4404 29948 4468 29952
rect 4404 29892 4408 29948
rect 4408 29892 4464 29948
rect 4464 29892 4468 29948
rect 4404 29888 4468 29892
rect 4484 29948 4548 29952
rect 4484 29892 4488 29948
rect 4488 29892 4544 29948
rect 4544 29892 4548 29948
rect 4484 29888 4548 29892
rect 4564 29948 4628 29952
rect 4564 29892 4568 29948
rect 4568 29892 4624 29948
rect 4624 29892 4628 29948
rect 4564 29888 4628 29892
rect 2084 29684 2148 29748
rect 2452 29684 2516 29748
rect 3188 29744 3252 29748
rect 3188 29688 3202 29744
rect 3202 29688 3252 29744
rect 3188 29684 3252 29688
rect 244 29548 308 29612
rect 1348 29548 1412 29612
rect 10724 29948 10788 29952
rect 10724 29892 10728 29948
rect 10728 29892 10784 29948
rect 10784 29892 10788 29948
rect 10724 29888 10788 29892
rect 10804 29948 10868 29952
rect 10804 29892 10808 29948
rect 10808 29892 10864 29948
rect 10864 29892 10868 29948
rect 10804 29888 10868 29892
rect 10884 29948 10948 29952
rect 10884 29892 10888 29948
rect 10888 29892 10944 29948
rect 10944 29892 10948 29948
rect 10884 29888 10948 29892
rect 10964 29948 11028 29952
rect 10964 29892 10968 29948
rect 10968 29892 11024 29948
rect 11024 29892 11028 29948
rect 10964 29888 11028 29892
rect 5948 29548 6012 29612
rect 4108 29412 4172 29476
rect 6316 29412 6380 29476
rect 3664 29404 3728 29408
rect 3664 29348 3668 29404
rect 3668 29348 3724 29404
rect 3724 29348 3728 29404
rect 3664 29344 3728 29348
rect 3744 29404 3808 29408
rect 3744 29348 3748 29404
rect 3748 29348 3804 29404
rect 3804 29348 3808 29404
rect 3744 29344 3808 29348
rect 3824 29404 3888 29408
rect 3824 29348 3828 29404
rect 3828 29348 3884 29404
rect 3884 29348 3888 29404
rect 3824 29344 3888 29348
rect 3904 29404 3968 29408
rect 3904 29348 3908 29404
rect 3908 29348 3964 29404
rect 3964 29348 3968 29404
rect 3904 29344 3968 29348
rect 980 29276 1044 29340
rect 4844 29276 4908 29340
rect 10064 29404 10128 29408
rect 10064 29348 10068 29404
rect 10068 29348 10124 29404
rect 10124 29348 10128 29404
rect 10064 29344 10128 29348
rect 10144 29404 10208 29408
rect 10144 29348 10148 29404
rect 10148 29348 10204 29404
rect 10204 29348 10208 29404
rect 10144 29344 10208 29348
rect 10224 29404 10288 29408
rect 10224 29348 10228 29404
rect 10228 29348 10284 29404
rect 10284 29348 10288 29404
rect 10224 29344 10288 29348
rect 10304 29404 10368 29408
rect 10304 29348 10308 29404
rect 10308 29348 10364 29404
rect 10364 29348 10368 29404
rect 10304 29344 10368 29348
rect 2452 29140 2516 29204
rect 3372 29140 3436 29204
rect 4844 29140 4908 29204
rect 5212 29140 5276 29204
rect 1532 29004 1596 29068
rect 2820 29004 2884 29068
rect 9444 29140 9508 29204
rect 7788 29004 7852 29068
rect 8708 29004 8772 29068
rect 796 28732 860 28796
rect 1164 27916 1228 27980
rect 244 27780 308 27844
rect 1164 27780 1228 27844
rect 244 27508 308 27572
rect 3372 28868 3436 28932
rect 5028 28928 5092 28932
rect 5028 28872 5042 28928
rect 5042 28872 5092 28928
rect 5028 28868 5092 28872
rect 4324 28860 4388 28864
rect 4324 28804 4328 28860
rect 4328 28804 4384 28860
rect 4384 28804 4388 28860
rect 4324 28800 4388 28804
rect 4404 28860 4468 28864
rect 4404 28804 4408 28860
rect 4408 28804 4464 28860
rect 4464 28804 4468 28860
rect 4404 28800 4468 28804
rect 4484 28860 4548 28864
rect 4484 28804 4488 28860
rect 4488 28804 4544 28860
rect 4544 28804 4548 28860
rect 4484 28800 4548 28804
rect 4564 28860 4628 28864
rect 4564 28804 4568 28860
rect 4568 28804 4624 28860
rect 4624 28804 4628 28860
rect 4564 28800 4628 28804
rect 2268 28732 2332 28796
rect 2820 28732 2884 28796
rect 4108 28732 4172 28796
rect 6132 28732 6196 28796
rect 10724 28860 10788 28864
rect 10724 28804 10728 28860
rect 10728 28804 10784 28860
rect 10784 28804 10788 28860
rect 10724 28800 10788 28804
rect 10804 28860 10868 28864
rect 10804 28804 10808 28860
rect 10808 28804 10864 28860
rect 10864 28804 10868 28860
rect 10804 28800 10868 28804
rect 10884 28860 10948 28864
rect 10884 28804 10888 28860
rect 10888 28804 10944 28860
rect 10944 28804 10948 28860
rect 10884 28800 10948 28804
rect 10964 28860 11028 28864
rect 10964 28804 10968 28860
rect 10968 28804 11024 28860
rect 11024 28804 11028 28860
rect 10964 28800 11028 28804
rect 6316 28596 6380 28660
rect 3004 28460 3068 28524
rect 3372 28460 3436 28524
rect 4108 28460 4172 28524
rect 7420 28520 7484 28524
rect 7420 28464 7434 28520
rect 7434 28464 7484 28520
rect 7420 28460 7484 28464
rect 2084 28324 2148 28388
rect 2084 28188 2148 28252
rect 3004 28188 3068 28252
rect 3664 28316 3728 28320
rect 3664 28260 3668 28316
rect 3668 28260 3724 28316
rect 3724 28260 3728 28316
rect 3664 28256 3728 28260
rect 3744 28316 3808 28320
rect 3744 28260 3748 28316
rect 3748 28260 3804 28316
rect 3804 28260 3808 28316
rect 3744 28256 3808 28260
rect 3824 28316 3888 28320
rect 3824 28260 3828 28316
rect 3828 28260 3884 28316
rect 3884 28260 3888 28316
rect 3824 28256 3888 28260
rect 3904 28316 3968 28320
rect 3904 28260 3908 28316
rect 3908 28260 3964 28316
rect 3964 28260 3968 28316
rect 3904 28256 3968 28260
rect 6500 28324 6564 28388
rect 10064 28316 10128 28320
rect 10064 28260 10068 28316
rect 10068 28260 10124 28316
rect 10124 28260 10128 28316
rect 10064 28256 10128 28260
rect 10144 28316 10208 28320
rect 10144 28260 10148 28316
rect 10148 28260 10204 28316
rect 10204 28260 10208 28316
rect 10144 28256 10208 28260
rect 10224 28316 10288 28320
rect 10224 28260 10228 28316
rect 10228 28260 10284 28316
rect 10284 28260 10288 28316
rect 10224 28256 10288 28260
rect 10304 28316 10368 28320
rect 10304 28260 10308 28316
rect 10308 28260 10364 28316
rect 10364 28260 10368 28316
rect 10304 28256 10368 28260
rect 6132 28112 6196 28116
rect 6132 28056 6182 28112
rect 6182 28056 6196 28112
rect 6132 28052 6196 28056
rect 3188 27644 3252 27708
rect 8524 27916 8588 27980
rect 10548 27916 10612 27980
rect 4324 27772 4388 27776
rect 4324 27716 4328 27772
rect 4328 27716 4384 27772
rect 4384 27716 4388 27772
rect 4324 27712 4388 27716
rect 4404 27772 4468 27776
rect 4404 27716 4408 27772
rect 4408 27716 4464 27772
rect 4464 27716 4468 27772
rect 4404 27712 4468 27716
rect 4484 27772 4548 27776
rect 4484 27716 4488 27772
rect 4488 27716 4544 27772
rect 4544 27716 4548 27772
rect 4484 27712 4548 27716
rect 4564 27772 4628 27776
rect 4564 27716 4568 27772
rect 4568 27716 4624 27772
rect 4624 27716 4628 27772
rect 4564 27712 4628 27716
rect 10724 27772 10788 27776
rect 10724 27716 10728 27772
rect 10728 27716 10784 27772
rect 10784 27716 10788 27772
rect 10724 27712 10788 27716
rect 10804 27772 10868 27776
rect 10804 27716 10808 27772
rect 10808 27716 10864 27772
rect 10864 27716 10868 27772
rect 10804 27712 10868 27716
rect 10884 27772 10948 27776
rect 10884 27716 10888 27772
rect 10888 27716 10944 27772
rect 10944 27716 10948 27772
rect 10884 27712 10948 27716
rect 10964 27772 11028 27776
rect 10964 27716 10968 27772
rect 10968 27716 11024 27772
rect 11024 27716 11028 27772
rect 10964 27712 11028 27716
rect 7604 27644 7668 27708
rect 612 27372 676 27436
rect 5212 27372 5276 27436
rect 5212 27236 5276 27300
rect 5948 27236 6012 27300
rect 3664 27228 3728 27232
rect 3664 27172 3668 27228
rect 3668 27172 3724 27228
rect 3724 27172 3728 27228
rect 3664 27168 3728 27172
rect 3744 27228 3808 27232
rect 3744 27172 3748 27228
rect 3748 27172 3804 27228
rect 3804 27172 3808 27228
rect 3744 27168 3808 27172
rect 3824 27228 3888 27232
rect 3824 27172 3828 27228
rect 3828 27172 3884 27228
rect 3884 27172 3888 27228
rect 3824 27168 3888 27172
rect 3904 27228 3968 27232
rect 3904 27172 3908 27228
rect 3908 27172 3964 27228
rect 3964 27172 3968 27228
rect 3904 27168 3968 27172
rect 5764 27100 5828 27164
rect 1900 26964 1964 27028
rect 3372 26828 3436 26892
rect 3372 26692 3436 26756
rect 5580 26692 5644 26756
rect 6316 26964 6380 27028
rect 10548 27372 10612 27436
rect 9444 27236 9508 27300
rect 10064 27228 10128 27232
rect 10064 27172 10068 27228
rect 10068 27172 10124 27228
rect 10124 27172 10128 27228
rect 10064 27168 10128 27172
rect 10144 27228 10208 27232
rect 10144 27172 10148 27228
rect 10148 27172 10204 27228
rect 10204 27172 10208 27228
rect 10144 27168 10208 27172
rect 10224 27228 10288 27232
rect 10224 27172 10228 27228
rect 10228 27172 10284 27228
rect 10284 27172 10288 27228
rect 10224 27168 10288 27172
rect 10304 27228 10368 27232
rect 10304 27172 10308 27228
rect 10308 27172 10364 27228
rect 10364 27172 10368 27228
rect 10304 27168 10368 27172
rect 9260 26828 9324 26892
rect 11284 26828 11348 26892
rect 4324 26684 4388 26688
rect 4324 26628 4328 26684
rect 4328 26628 4384 26684
rect 4384 26628 4388 26684
rect 4324 26624 4388 26628
rect 4404 26684 4468 26688
rect 4404 26628 4408 26684
rect 4408 26628 4464 26684
rect 4464 26628 4468 26684
rect 4404 26624 4468 26628
rect 4484 26684 4548 26688
rect 4484 26628 4488 26684
rect 4488 26628 4544 26684
rect 4544 26628 4548 26684
rect 4484 26624 4548 26628
rect 4564 26684 4628 26688
rect 4564 26628 4568 26684
rect 4568 26628 4624 26684
rect 4624 26628 4628 26684
rect 4564 26624 4628 26628
rect 10724 26684 10788 26688
rect 10724 26628 10728 26684
rect 10728 26628 10784 26684
rect 10784 26628 10788 26684
rect 10724 26624 10788 26628
rect 10804 26684 10868 26688
rect 10804 26628 10808 26684
rect 10808 26628 10864 26684
rect 10864 26628 10868 26684
rect 10804 26624 10868 26628
rect 10884 26684 10948 26688
rect 10884 26628 10888 26684
rect 10888 26628 10944 26684
rect 10944 26628 10948 26684
rect 10884 26624 10948 26628
rect 10964 26684 11028 26688
rect 10964 26628 10968 26684
rect 10968 26628 11024 26684
rect 11024 26628 11028 26684
rect 10964 26624 11028 26628
rect 2084 26420 2148 26484
rect 1348 26148 1412 26212
rect 5580 26556 5644 26620
rect 10548 26556 10612 26620
rect 11100 26556 11164 26620
rect 7052 26420 7116 26484
rect 3188 26148 3252 26212
rect 1716 26012 1780 26076
rect 3188 26012 3252 26076
rect 4844 26284 4908 26348
rect 6316 26284 6380 26348
rect 4706 26148 4770 26212
rect 5764 26148 5828 26212
rect 8156 26284 8220 26348
rect 8892 26284 8956 26348
rect 8156 26148 8220 26212
rect 3664 26140 3728 26144
rect 3664 26084 3668 26140
rect 3668 26084 3724 26140
rect 3724 26084 3728 26140
rect 3664 26080 3728 26084
rect 3744 26140 3808 26144
rect 3744 26084 3748 26140
rect 3748 26084 3804 26140
rect 3804 26084 3808 26140
rect 3744 26080 3808 26084
rect 3824 26140 3888 26144
rect 3824 26084 3828 26140
rect 3828 26084 3884 26140
rect 3884 26084 3888 26140
rect 3824 26080 3888 26084
rect 3904 26140 3968 26144
rect 3904 26084 3908 26140
rect 3908 26084 3964 26140
rect 3964 26084 3968 26140
rect 3904 26080 3968 26084
rect 1532 25876 1596 25940
rect 1716 25876 1780 25940
rect 8340 26012 8404 26076
rect 6500 25876 6564 25940
rect 7972 25876 8036 25940
rect 1348 25740 1412 25804
rect 1900 25740 1964 25804
rect 3004 25740 3068 25804
rect 3188 25740 3252 25804
rect 10064 26140 10128 26144
rect 10064 26084 10068 26140
rect 10068 26084 10124 26140
rect 10124 26084 10128 26140
rect 10064 26080 10128 26084
rect 10144 26140 10208 26144
rect 10144 26084 10148 26140
rect 10148 26084 10204 26140
rect 10204 26084 10208 26140
rect 10144 26080 10208 26084
rect 10224 26140 10288 26144
rect 10224 26084 10228 26140
rect 10228 26084 10284 26140
rect 10284 26084 10288 26140
rect 10224 26080 10288 26084
rect 10304 26140 10368 26144
rect 10304 26084 10308 26140
rect 10308 26084 10364 26140
rect 10364 26084 10368 26140
rect 10304 26080 10368 26084
rect 6316 25740 6380 25804
rect 3188 25604 3252 25668
rect 4324 25596 4388 25600
rect 4324 25540 4328 25596
rect 4328 25540 4384 25596
rect 4384 25540 4388 25596
rect 4324 25536 4388 25540
rect 4404 25596 4468 25600
rect 4404 25540 4408 25596
rect 4408 25540 4464 25596
rect 4464 25540 4468 25596
rect 4404 25536 4468 25540
rect 4484 25596 4548 25600
rect 4484 25540 4488 25596
rect 4488 25540 4544 25596
rect 4544 25540 4548 25596
rect 4484 25536 4548 25540
rect 4564 25596 4628 25600
rect 4564 25540 4568 25596
rect 4568 25540 4624 25596
rect 4624 25540 4628 25596
rect 4564 25536 4628 25540
rect 5764 25604 5828 25668
rect 10724 25596 10788 25600
rect 10724 25540 10728 25596
rect 10728 25540 10784 25596
rect 10784 25540 10788 25596
rect 10724 25536 10788 25540
rect 10804 25596 10868 25600
rect 10804 25540 10808 25596
rect 10808 25540 10864 25596
rect 10864 25540 10868 25596
rect 10804 25536 10868 25540
rect 10884 25596 10948 25600
rect 10884 25540 10888 25596
rect 10888 25540 10944 25596
rect 10944 25540 10948 25596
rect 10884 25536 10948 25540
rect 10964 25596 11028 25600
rect 10964 25540 10968 25596
rect 10968 25540 11024 25596
rect 11024 25540 11028 25596
rect 10964 25536 11028 25540
rect 2084 25332 2148 25396
rect 3004 25332 3068 25396
rect 3372 25196 3436 25260
rect 2268 25060 2332 25124
rect 5212 25196 5276 25260
rect 9260 25332 9324 25396
rect 8524 25196 8588 25260
rect 6500 25120 6564 25124
rect 6500 25064 6514 25120
rect 6514 25064 6564 25120
rect 3664 25052 3728 25056
rect 3664 24996 3668 25052
rect 3668 24996 3724 25052
rect 3724 24996 3728 25052
rect 3664 24992 3728 24996
rect 3744 25052 3808 25056
rect 3744 24996 3748 25052
rect 3748 24996 3804 25052
rect 3804 24996 3808 25052
rect 3744 24992 3808 24996
rect 3824 25052 3888 25056
rect 3824 24996 3828 25052
rect 3828 24996 3884 25052
rect 3884 24996 3888 25052
rect 3824 24992 3888 24996
rect 3904 25052 3968 25056
rect 3904 24996 3908 25052
rect 3908 24996 3964 25052
rect 3964 24996 3968 25052
rect 3904 24992 3968 24996
rect 2268 24984 2332 24988
rect 2268 24928 2318 24984
rect 2318 24928 2332 24984
rect 2268 24924 2332 24928
rect 6500 25060 6564 25064
rect 8524 25060 8588 25124
rect 8892 25060 8956 25124
rect 10064 25052 10128 25056
rect 10064 24996 10068 25052
rect 10068 24996 10124 25052
rect 10124 24996 10128 25052
rect 10064 24992 10128 24996
rect 10144 25052 10208 25056
rect 10144 24996 10148 25052
rect 10148 24996 10204 25052
rect 10204 24996 10208 25052
rect 10144 24992 10208 24996
rect 10224 25052 10288 25056
rect 10224 24996 10228 25052
rect 10228 24996 10284 25052
rect 10284 24996 10288 25052
rect 10224 24992 10288 24996
rect 10304 25052 10368 25056
rect 10304 24996 10308 25052
rect 10308 24996 10364 25052
rect 10364 24996 10368 25052
rect 10304 24992 10368 24996
rect 7972 24924 8036 24988
rect 8892 24924 8956 24988
rect 5580 24712 5644 24716
rect 5580 24656 5630 24712
rect 5630 24656 5644 24712
rect 5580 24652 5644 24656
rect 1532 24516 1596 24580
rect 4706 24516 4770 24580
rect 4324 24508 4388 24512
rect 4324 24452 4328 24508
rect 4328 24452 4384 24508
rect 4384 24452 4388 24508
rect 4324 24448 4388 24452
rect 4404 24508 4468 24512
rect 4404 24452 4408 24508
rect 4408 24452 4464 24508
rect 4464 24452 4468 24508
rect 4404 24448 4468 24452
rect 4484 24508 4548 24512
rect 4484 24452 4488 24508
rect 4488 24452 4544 24508
rect 4544 24452 4548 24508
rect 4484 24448 4548 24452
rect 4564 24508 4628 24512
rect 4564 24452 4568 24508
rect 4568 24452 4624 24508
rect 4624 24452 4628 24508
rect 4564 24448 4628 24452
rect 6868 24652 6932 24716
rect 8708 24652 8772 24716
rect 6132 24516 6196 24580
rect 10724 24508 10788 24512
rect 10724 24452 10728 24508
rect 10728 24452 10784 24508
rect 10784 24452 10788 24508
rect 10724 24448 10788 24452
rect 10804 24508 10868 24512
rect 10804 24452 10808 24508
rect 10808 24452 10864 24508
rect 10864 24452 10868 24508
rect 10804 24448 10868 24452
rect 10884 24508 10948 24512
rect 10884 24452 10888 24508
rect 10888 24452 10944 24508
rect 10944 24452 10948 24508
rect 10884 24448 10948 24452
rect 10964 24508 11028 24512
rect 10964 24452 10968 24508
rect 10968 24452 11024 24508
rect 11024 24452 11028 24508
rect 10964 24448 11028 24452
rect 5212 24380 5276 24444
rect 5764 24440 5828 24444
rect 5764 24384 5778 24440
rect 5778 24384 5828 24440
rect 5764 24380 5828 24384
rect 6132 24380 6196 24444
rect 7052 24380 7116 24444
rect 1900 24244 1964 24308
rect 11100 24244 11164 24308
rect 1348 24108 1412 24172
rect 1900 24108 1964 24172
rect 10548 24108 10612 24172
rect 11100 24108 11164 24172
rect 7236 23972 7300 24036
rect 3664 23964 3728 23968
rect 3664 23908 3668 23964
rect 3668 23908 3724 23964
rect 3724 23908 3728 23964
rect 3664 23904 3728 23908
rect 3744 23964 3808 23968
rect 3744 23908 3748 23964
rect 3748 23908 3804 23964
rect 3804 23908 3808 23964
rect 3744 23904 3808 23908
rect 3824 23964 3888 23968
rect 3824 23908 3828 23964
rect 3828 23908 3884 23964
rect 3884 23908 3888 23964
rect 3824 23904 3888 23908
rect 3904 23964 3968 23968
rect 3904 23908 3908 23964
rect 3908 23908 3964 23964
rect 3964 23908 3968 23964
rect 3904 23904 3968 23908
rect 10548 23972 10612 24036
rect 10064 23964 10128 23968
rect 10064 23908 10068 23964
rect 10068 23908 10124 23964
rect 10124 23908 10128 23964
rect 10064 23904 10128 23908
rect 10144 23964 10208 23968
rect 10144 23908 10148 23964
rect 10148 23908 10204 23964
rect 10204 23908 10208 23964
rect 10144 23904 10208 23908
rect 10224 23964 10288 23968
rect 10224 23908 10228 23964
rect 10228 23908 10284 23964
rect 10284 23908 10288 23964
rect 10224 23904 10288 23908
rect 10304 23964 10368 23968
rect 10304 23908 10308 23964
rect 10308 23908 10364 23964
rect 10364 23908 10368 23964
rect 10304 23904 10368 23908
rect 9260 23896 9324 23900
rect 9260 23840 9274 23896
rect 9274 23840 9324 23896
rect 9260 23836 9324 23840
rect 1164 23564 1228 23628
rect 6868 23700 6932 23764
rect 7052 23700 7116 23764
rect 1348 23488 1412 23492
rect 1348 23432 1398 23488
rect 1398 23432 1412 23488
rect 1348 23428 1412 23432
rect 1716 23428 1780 23492
rect 1716 23292 1780 23356
rect 2084 23292 2148 23356
rect 2452 23156 2516 23220
rect 1164 23080 1228 23084
rect 7420 23564 7484 23628
rect 8708 23624 8772 23628
rect 8708 23568 8722 23624
rect 8722 23568 8772 23624
rect 8708 23564 8772 23568
rect 9444 23700 9508 23764
rect 9444 23428 9508 23492
rect 4324 23420 4388 23424
rect 4324 23364 4328 23420
rect 4328 23364 4384 23420
rect 4384 23364 4388 23420
rect 4324 23360 4388 23364
rect 4404 23420 4468 23424
rect 4404 23364 4408 23420
rect 4408 23364 4464 23420
rect 4464 23364 4468 23420
rect 4404 23360 4468 23364
rect 4484 23420 4548 23424
rect 4484 23364 4488 23420
rect 4488 23364 4544 23420
rect 4544 23364 4548 23420
rect 4484 23360 4548 23364
rect 4564 23420 4628 23424
rect 4564 23364 4568 23420
rect 4568 23364 4624 23420
rect 4624 23364 4628 23420
rect 4564 23360 4628 23364
rect 10724 23420 10788 23424
rect 10724 23364 10728 23420
rect 10728 23364 10784 23420
rect 10784 23364 10788 23420
rect 10724 23360 10788 23364
rect 10804 23420 10868 23424
rect 10804 23364 10808 23420
rect 10808 23364 10864 23420
rect 10864 23364 10868 23420
rect 10804 23360 10868 23364
rect 10884 23420 10948 23424
rect 10884 23364 10888 23420
rect 10888 23364 10944 23420
rect 10944 23364 10948 23420
rect 10884 23360 10948 23364
rect 10964 23420 11028 23424
rect 10964 23364 10968 23420
rect 10968 23364 11024 23420
rect 11024 23364 11028 23420
rect 10964 23360 11028 23364
rect 8892 23292 8956 23356
rect 6868 23156 6932 23220
rect 7236 23156 7300 23220
rect 8524 23156 8588 23220
rect 11100 23156 11164 23220
rect 1164 23024 1214 23080
rect 1214 23024 1228 23080
rect 1164 23020 1228 23024
rect 4108 22884 4172 22948
rect 7420 22884 7484 22948
rect 7788 22884 7852 22948
rect 8156 22884 8220 22948
rect 8524 22884 8588 22948
rect 9444 22884 9508 22948
rect 3664 22876 3728 22880
rect 3664 22820 3668 22876
rect 3668 22820 3724 22876
rect 3724 22820 3728 22876
rect 3664 22816 3728 22820
rect 3744 22876 3808 22880
rect 3744 22820 3748 22876
rect 3748 22820 3804 22876
rect 3804 22820 3808 22876
rect 3744 22816 3808 22820
rect 3824 22876 3888 22880
rect 3824 22820 3828 22876
rect 3828 22820 3884 22876
rect 3884 22820 3888 22876
rect 3824 22816 3888 22820
rect 3904 22876 3968 22880
rect 3904 22820 3908 22876
rect 3908 22820 3964 22876
rect 3964 22820 3968 22876
rect 3904 22816 3968 22820
rect 10064 22876 10128 22880
rect 10064 22820 10068 22876
rect 10068 22820 10124 22876
rect 10124 22820 10128 22876
rect 10064 22816 10128 22820
rect 10144 22876 10208 22880
rect 10144 22820 10148 22876
rect 10148 22820 10204 22876
rect 10204 22820 10208 22876
rect 10144 22816 10208 22820
rect 10224 22876 10288 22880
rect 10224 22820 10228 22876
rect 10228 22820 10284 22876
rect 10284 22820 10288 22876
rect 10224 22816 10288 22820
rect 10304 22876 10368 22880
rect 10304 22820 10308 22876
rect 10308 22820 10364 22876
rect 10364 22820 10368 22876
rect 10304 22816 10368 22820
rect 4108 22748 4172 22812
rect 9260 22748 9324 22812
rect 5948 22612 6012 22676
rect 6500 22612 6564 22676
rect 8708 22612 8772 22676
rect 1900 22476 1964 22540
rect 2452 22476 2516 22540
rect 428 22340 492 22404
rect 2452 22400 2516 22404
rect 2452 22344 2502 22400
rect 2502 22344 2516 22400
rect 2452 22340 2516 22344
rect 2820 22340 2884 22404
rect 3188 22340 3252 22404
rect 796 22204 860 22268
rect 4324 22332 4388 22336
rect 4324 22276 4328 22332
rect 4328 22276 4384 22332
rect 4384 22276 4388 22332
rect 4324 22272 4388 22276
rect 4404 22332 4468 22336
rect 4404 22276 4408 22332
rect 4408 22276 4464 22332
rect 4464 22276 4468 22332
rect 4404 22272 4468 22276
rect 4484 22332 4548 22336
rect 4484 22276 4488 22332
rect 4488 22276 4544 22332
rect 4544 22276 4548 22332
rect 4484 22272 4548 22276
rect 4564 22332 4628 22336
rect 4564 22276 4568 22332
rect 4568 22276 4624 22332
rect 4624 22276 4628 22332
rect 4564 22272 4628 22276
rect 7236 22476 7300 22540
rect 5212 22340 5276 22404
rect 8156 22340 8220 22404
rect 10724 22332 10788 22336
rect 10724 22276 10728 22332
rect 10728 22276 10784 22332
rect 10784 22276 10788 22332
rect 10724 22272 10788 22276
rect 10804 22332 10868 22336
rect 10804 22276 10808 22332
rect 10808 22276 10864 22332
rect 10864 22276 10868 22332
rect 10804 22272 10868 22276
rect 10884 22332 10948 22336
rect 10884 22276 10888 22332
rect 10888 22276 10944 22332
rect 10944 22276 10948 22332
rect 10884 22272 10948 22276
rect 10964 22332 11028 22336
rect 10964 22276 10968 22332
rect 10968 22276 11024 22332
rect 11024 22276 11028 22332
rect 10964 22272 11028 22276
rect 6500 22204 6564 22268
rect 980 22068 1044 22132
rect 2820 22068 2884 22132
rect 7788 22068 7852 22132
rect 5948 21992 6012 21996
rect 5948 21936 5998 21992
rect 5998 21936 6012 21992
rect 5948 21932 6012 21936
rect 6316 21992 6380 21996
rect 6316 21936 6330 21992
rect 6330 21936 6380 21992
rect 6316 21932 6380 21936
rect 6868 21932 6932 21996
rect 8340 21992 8404 21996
rect 8340 21936 8390 21992
rect 8390 21936 8404 21992
rect 8340 21932 8404 21936
rect 3188 21796 3252 21860
rect 9444 21796 9508 21860
rect 10548 21856 10612 21860
rect 10548 21800 10598 21856
rect 10598 21800 10612 21856
rect 10548 21796 10612 21800
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 10064 21788 10128 21792
rect 10064 21732 10068 21788
rect 10068 21732 10124 21788
rect 10124 21732 10128 21788
rect 10064 21728 10128 21732
rect 10144 21788 10208 21792
rect 10144 21732 10148 21788
rect 10148 21732 10204 21788
rect 10204 21732 10208 21788
rect 10144 21728 10208 21732
rect 10224 21788 10288 21792
rect 10224 21732 10228 21788
rect 10228 21732 10284 21788
rect 10284 21732 10288 21788
rect 10224 21728 10288 21732
rect 10304 21788 10368 21792
rect 10304 21732 10308 21788
rect 10308 21732 10364 21788
rect 10364 21732 10368 21788
rect 10304 21728 10368 21732
rect 5580 21524 5644 21588
rect 8340 21524 8404 21588
rect 9812 21524 9876 21588
rect 10548 21524 10612 21588
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 10724 21244 10788 21248
rect 10724 21188 10728 21244
rect 10728 21188 10784 21244
rect 10784 21188 10788 21244
rect 10724 21184 10788 21188
rect 10804 21244 10868 21248
rect 10804 21188 10808 21244
rect 10808 21188 10864 21244
rect 10864 21188 10868 21244
rect 10804 21184 10868 21188
rect 10884 21244 10948 21248
rect 10884 21188 10888 21244
rect 10888 21188 10944 21244
rect 10944 21188 10948 21244
rect 10884 21184 10948 21188
rect 10964 21244 11028 21248
rect 10964 21188 10968 21244
rect 10968 21188 11024 21244
rect 11024 21188 11028 21244
rect 10964 21184 11028 21188
rect 1532 21116 1596 21180
rect 5396 21116 5460 21180
rect 5580 21176 5644 21180
rect 5580 21120 5594 21176
rect 5594 21120 5644 21176
rect 5580 21116 5644 21120
rect 7604 20844 7668 20908
rect 8708 20844 8772 20908
rect 5028 20708 5092 20772
rect 9628 20708 9692 20772
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 10064 20700 10128 20704
rect 10064 20644 10068 20700
rect 10068 20644 10124 20700
rect 10124 20644 10128 20700
rect 10064 20640 10128 20644
rect 10144 20700 10208 20704
rect 10144 20644 10148 20700
rect 10148 20644 10204 20700
rect 10204 20644 10208 20700
rect 10144 20640 10208 20644
rect 10224 20700 10288 20704
rect 10224 20644 10228 20700
rect 10228 20644 10284 20700
rect 10284 20644 10288 20700
rect 10224 20640 10288 20644
rect 10304 20700 10368 20704
rect 10304 20644 10308 20700
rect 10308 20644 10364 20700
rect 10364 20644 10368 20700
rect 10304 20640 10368 20644
rect 980 20572 1044 20636
rect 2452 20572 2516 20636
rect 60 20436 124 20500
rect 5212 20436 5276 20500
rect 8524 20496 8588 20500
rect 8524 20440 8538 20496
rect 8538 20440 8588 20496
rect 8524 20436 8588 20440
rect 6684 20300 6748 20364
rect 2452 20164 2516 20228
rect 4108 20164 4172 20228
rect 5396 20164 5460 20228
rect 6868 20164 6932 20228
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 10724 20156 10788 20160
rect 10724 20100 10728 20156
rect 10728 20100 10784 20156
rect 10784 20100 10788 20156
rect 10724 20096 10788 20100
rect 10804 20156 10868 20160
rect 10804 20100 10808 20156
rect 10808 20100 10864 20156
rect 10864 20100 10868 20156
rect 10804 20096 10868 20100
rect 10884 20156 10948 20160
rect 10884 20100 10888 20156
rect 10888 20100 10944 20156
rect 10944 20100 10948 20156
rect 10884 20096 10948 20100
rect 10964 20156 11028 20160
rect 10964 20100 10968 20156
rect 10968 20100 11024 20156
rect 11024 20100 11028 20156
rect 10964 20096 11028 20100
rect 2084 19892 2148 19956
rect 6684 20028 6748 20092
rect 6316 19756 6380 19820
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 10064 19612 10128 19616
rect 10064 19556 10068 19612
rect 10068 19556 10124 19612
rect 10124 19556 10128 19612
rect 10064 19552 10128 19556
rect 10144 19612 10208 19616
rect 10144 19556 10148 19612
rect 10148 19556 10204 19612
rect 10204 19556 10208 19612
rect 10144 19552 10208 19556
rect 10224 19612 10288 19616
rect 10224 19556 10228 19612
rect 10228 19556 10284 19612
rect 10284 19556 10288 19612
rect 10224 19552 10288 19556
rect 10304 19612 10368 19616
rect 10304 19556 10308 19612
rect 10308 19556 10364 19612
rect 10364 19556 10368 19612
rect 10304 19552 10368 19556
rect 8892 19484 8956 19548
rect 7052 19348 7116 19412
rect 2636 19212 2700 19276
rect 11284 19272 11348 19276
rect 11284 19216 11298 19272
rect 11298 19216 11348 19272
rect 11284 19212 11348 19216
rect 6316 19076 6380 19140
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 10724 19068 10788 19072
rect 10724 19012 10728 19068
rect 10728 19012 10784 19068
rect 10784 19012 10788 19068
rect 10724 19008 10788 19012
rect 10804 19068 10868 19072
rect 10804 19012 10808 19068
rect 10808 19012 10864 19068
rect 10864 19012 10868 19068
rect 10804 19008 10868 19012
rect 10884 19068 10948 19072
rect 10884 19012 10888 19068
rect 10888 19012 10944 19068
rect 10944 19012 10948 19068
rect 10884 19008 10948 19012
rect 10964 19068 11028 19072
rect 10964 19012 10968 19068
rect 10968 19012 11024 19068
rect 11024 19012 11028 19068
rect 10964 19008 11028 19012
rect 2636 18804 2700 18868
rect 11284 18804 11348 18868
rect 5028 18668 5092 18732
rect 9812 18668 9876 18732
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 7420 18532 7484 18596
rect 8340 18532 8404 18596
rect 10064 18524 10128 18528
rect 10064 18468 10068 18524
rect 10068 18468 10124 18524
rect 10124 18468 10128 18524
rect 10064 18464 10128 18468
rect 10144 18524 10208 18528
rect 10144 18468 10148 18524
rect 10148 18468 10204 18524
rect 10204 18468 10208 18524
rect 10144 18464 10208 18468
rect 10224 18524 10288 18528
rect 10224 18468 10228 18524
rect 10228 18468 10284 18524
rect 10284 18468 10288 18524
rect 10224 18464 10288 18468
rect 10304 18524 10368 18528
rect 10304 18468 10308 18524
rect 10308 18468 10364 18524
rect 10364 18468 10368 18524
rect 10304 18464 10368 18468
rect 4844 18260 4908 18324
rect 5212 18260 5276 18324
rect 5764 18320 5828 18324
rect 5764 18264 5778 18320
rect 5778 18264 5828 18320
rect 5764 18260 5828 18264
rect 11100 18320 11164 18324
rect 11100 18264 11150 18320
rect 11150 18264 11164 18320
rect 4108 18124 4172 18188
rect 5396 18124 5460 18188
rect 11100 18260 11164 18264
rect 6868 18124 6932 18188
rect 612 18048 676 18052
rect 612 17992 662 18048
rect 662 17992 676 18048
rect 612 17988 676 17992
rect 2820 17988 2884 18052
rect 5028 17988 5092 18052
rect 7972 18124 8036 18188
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 10724 17980 10788 17984
rect 10724 17924 10728 17980
rect 10728 17924 10784 17980
rect 10784 17924 10788 17980
rect 10724 17920 10788 17924
rect 10804 17980 10868 17984
rect 10804 17924 10808 17980
rect 10808 17924 10864 17980
rect 10864 17924 10868 17980
rect 10804 17920 10868 17924
rect 10884 17980 10948 17984
rect 10884 17924 10888 17980
rect 10888 17924 10944 17980
rect 10944 17924 10948 17980
rect 10884 17920 10948 17924
rect 10964 17980 11028 17984
rect 10964 17924 10968 17980
rect 10968 17924 11024 17980
rect 11024 17924 11028 17980
rect 10964 17920 11028 17924
rect 60 17852 124 17916
rect 5028 17716 5092 17780
rect 6316 17640 6380 17644
rect 6316 17584 6330 17640
rect 6330 17584 6380 17640
rect 6316 17580 6380 17584
rect 8524 17640 8588 17644
rect 8524 17584 8538 17640
rect 8538 17584 8588 17640
rect 8524 17580 8588 17584
rect 9444 17580 9508 17644
rect 244 17504 308 17508
rect 244 17448 294 17504
rect 294 17448 308 17504
rect 244 17444 308 17448
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 10064 17436 10128 17440
rect 10064 17380 10068 17436
rect 10068 17380 10124 17436
rect 10124 17380 10128 17436
rect 10064 17376 10128 17380
rect 10144 17436 10208 17440
rect 10144 17380 10148 17436
rect 10148 17380 10204 17436
rect 10204 17380 10208 17436
rect 10144 17376 10208 17380
rect 10224 17436 10288 17440
rect 10224 17380 10228 17436
rect 10228 17380 10284 17436
rect 10284 17380 10288 17436
rect 10224 17376 10288 17380
rect 10304 17436 10368 17440
rect 10304 17380 10308 17436
rect 10308 17380 10364 17436
rect 10364 17380 10368 17436
rect 10304 17376 10368 17380
rect 1532 17232 1596 17236
rect 1532 17176 1546 17232
rect 1546 17176 1596 17232
rect 1532 17172 1596 17176
rect 4844 17172 4908 17236
rect 6132 17172 6196 17236
rect 6684 17172 6748 17236
rect 8340 17172 8404 17236
rect 9076 17172 9140 17236
rect 1348 17036 1412 17100
rect 2636 16960 2700 16964
rect 2636 16904 2686 16960
rect 2686 16904 2700 16960
rect 2636 16900 2700 16904
rect 6868 16900 6932 16964
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 3372 16764 3436 16828
rect 7604 16764 7668 16828
rect 9260 16764 9324 16828
rect 10724 16892 10788 16896
rect 10724 16836 10728 16892
rect 10728 16836 10784 16892
rect 10784 16836 10788 16892
rect 10724 16832 10788 16836
rect 10804 16892 10868 16896
rect 10804 16836 10808 16892
rect 10808 16836 10864 16892
rect 10864 16836 10868 16892
rect 10804 16832 10868 16836
rect 10884 16892 10948 16896
rect 10884 16836 10888 16892
rect 10888 16836 10944 16892
rect 10944 16836 10948 16892
rect 10884 16832 10948 16836
rect 10964 16892 11028 16896
rect 10964 16836 10968 16892
rect 10968 16836 11024 16892
rect 11024 16836 11028 16892
rect 10964 16832 11028 16836
rect 9076 16688 9140 16692
rect 9076 16632 9126 16688
rect 9126 16632 9140 16688
rect 9076 16628 9140 16632
rect 7236 16492 7300 16556
rect 8892 16492 8956 16556
rect 796 16356 860 16420
rect 8708 16356 8772 16420
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 10064 16348 10128 16352
rect 10064 16292 10068 16348
rect 10068 16292 10124 16348
rect 10124 16292 10128 16348
rect 10064 16288 10128 16292
rect 10144 16348 10208 16352
rect 10144 16292 10148 16348
rect 10148 16292 10204 16348
rect 10204 16292 10208 16348
rect 10144 16288 10208 16292
rect 10224 16348 10288 16352
rect 10224 16292 10228 16348
rect 10228 16292 10284 16348
rect 10284 16292 10288 16348
rect 10224 16288 10288 16292
rect 10304 16348 10368 16352
rect 10304 16292 10308 16348
rect 10308 16292 10364 16348
rect 10364 16292 10368 16348
rect 10304 16288 10368 16292
rect 1716 16084 1780 16148
rect 3188 16084 3252 16148
rect 3004 15812 3068 15876
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 10724 15804 10788 15808
rect 10724 15748 10728 15804
rect 10728 15748 10784 15804
rect 10784 15748 10788 15804
rect 10724 15744 10788 15748
rect 10804 15804 10868 15808
rect 10804 15748 10808 15804
rect 10808 15748 10864 15804
rect 10864 15748 10868 15804
rect 10804 15744 10868 15748
rect 10884 15804 10948 15808
rect 10884 15748 10888 15804
rect 10888 15748 10944 15804
rect 10944 15748 10948 15804
rect 10884 15744 10948 15748
rect 10964 15804 11028 15808
rect 10964 15748 10968 15804
rect 10968 15748 11024 15804
rect 11024 15748 11028 15804
rect 10964 15744 11028 15748
rect 8340 15464 8404 15468
rect 8340 15408 8390 15464
rect 8390 15408 8404 15464
rect 8340 15404 8404 15408
rect 5580 15268 5644 15332
rect 10548 15404 10612 15468
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 2268 15192 2332 15196
rect 2268 15136 2282 15192
rect 2282 15136 2332 15192
rect 2268 15132 2332 15136
rect 4108 15132 4172 15196
rect 10064 15260 10128 15264
rect 10064 15204 10068 15260
rect 10068 15204 10124 15260
rect 10124 15204 10128 15260
rect 10064 15200 10128 15204
rect 10144 15260 10208 15264
rect 10144 15204 10148 15260
rect 10148 15204 10204 15260
rect 10204 15204 10208 15260
rect 10144 15200 10208 15204
rect 10224 15260 10288 15264
rect 10224 15204 10228 15260
rect 10228 15204 10284 15260
rect 10284 15204 10288 15260
rect 10224 15200 10288 15204
rect 10304 15260 10368 15264
rect 10304 15204 10308 15260
rect 10308 15204 10364 15260
rect 10364 15204 10368 15260
rect 10304 15200 10368 15204
rect 5948 14996 6012 15060
rect 9260 14996 9324 15060
rect 9628 14996 9692 15060
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 10724 14716 10788 14720
rect 10724 14660 10728 14716
rect 10728 14660 10784 14716
rect 10784 14660 10788 14716
rect 10724 14656 10788 14660
rect 10804 14716 10868 14720
rect 10804 14660 10808 14716
rect 10808 14660 10864 14716
rect 10864 14660 10868 14716
rect 10804 14656 10868 14660
rect 10884 14716 10948 14720
rect 10884 14660 10888 14716
rect 10888 14660 10944 14716
rect 10944 14660 10948 14716
rect 10884 14656 10948 14660
rect 10964 14716 11028 14720
rect 10964 14660 10968 14716
rect 10968 14660 11024 14716
rect 11024 14660 11028 14716
rect 10964 14656 11028 14660
rect 2820 14588 2884 14652
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 10064 14172 10128 14176
rect 10064 14116 10068 14172
rect 10068 14116 10124 14172
rect 10124 14116 10128 14172
rect 10064 14112 10128 14116
rect 10144 14172 10208 14176
rect 10144 14116 10148 14172
rect 10148 14116 10204 14172
rect 10204 14116 10208 14172
rect 10144 14112 10208 14116
rect 10224 14172 10288 14176
rect 10224 14116 10228 14172
rect 10228 14116 10284 14172
rect 10284 14116 10288 14172
rect 10224 14112 10288 14116
rect 10304 14172 10368 14176
rect 10304 14116 10308 14172
rect 10308 14116 10364 14172
rect 10364 14116 10368 14172
rect 10304 14112 10368 14116
rect 1532 13772 1596 13836
rect 4844 13772 4908 13836
rect 3004 13636 3068 13700
rect 7420 13636 7484 13700
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 10724 13628 10788 13632
rect 10724 13572 10728 13628
rect 10728 13572 10784 13628
rect 10784 13572 10788 13628
rect 10724 13568 10788 13572
rect 10804 13628 10868 13632
rect 10804 13572 10808 13628
rect 10808 13572 10864 13628
rect 10864 13572 10868 13628
rect 10804 13568 10868 13572
rect 10884 13628 10948 13632
rect 10884 13572 10888 13628
rect 10888 13572 10944 13628
rect 10944 13572 10948 13628
rect 10884 13568 10948 13572
rect 10964 13628 11028 13632
rect 10964 13572 10968 13628
rect 10968 13572 11024 13628
rect 11024 13572 11028 13628
rect 10964 13568 11028 13572
rect 9444 13500 9508 13564
rect 2820 13424 2884 13428
rect 2820 13368 2870 13424
rect 2870 13368 2884 13424
rect 2820 13364 2884 13368
rect 5028 13364 5092 13428
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 10064 13084 10128 13088
rect 10064 13028 10068 13084
rect 10068 13028 10124 13084
rect 10124 13028 10128 13084
rect 10064 13024 10128 13028
rect 10144 13084 10208 13088
rect 10144 13028 10148 13084
rect 10148 13028 10204 13084
rect 10204 13028 10208 13084
rect 10144 13024 10208 13028
rect 10224 13084 10288 13088
rect 10224 13028 10228 13084
rect 10228 13028 10284 13084
rect 10284 13028 10288 13084
rect 10224 13024 10288 13028
rect 10304 13084 10368 13088
rect 10304 13028 10308 13084
rect 10308 13028 10364 13084
rect 10364 13028 10368 13084
rect 10304 13024 10368 13028
rect 8156 12956 8220 13020
rect 2084 12820 2148 12884
rect 7236 12820 7300 12884
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 10724 12540 10788 12544
rect 10724 12484 10728 12540
rect 10728 12484 10784 12540
rect 10784 12484 10788 12540
rect 10724 12480 10788 12484
rect 10804 12540 10868 12544
rect 10804 12484 10808 12540
rect 10808 12484 10864 12540
rect 10864 12484 10868 12540
rect 10804 12480 10868 12484
rect 10884 12540 10948 12544
rect 10884 12484 10888 12540
rect 10888 12484 10944 12540
rect 10944 12484 10948 12540
rect 10884 12480 10948 12484
rect 10964 12540 11028 12544
rect 10964 12484 10968 12540
rect 10968 12484 11024 12540
rect 11024 12484 11028 12540
rect 10964 12480 11028 12484
rect 2452 12276 2516 12340
rect 1164 12004 1228 12068
rect 1900 12064 1964 12068
rect 1900 12008 1950 12064
rect 1950 12008 1964 12064
rect 1900 12004 1964 12008
rect 4108 12140 4172 12204
rect 8524 12200 8588 12204
rect 8524 12144 8538 12200
rect 8538 12144 8588 12200
rect 8524 12140 8588 12144
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 10064 11996 10128 12000
rect 10064 11940 10068 11996
rect 10068 11940 10124 11996
rect 10124 11940 10128 11996
rect 10064 11936 10128 11940
rect 10144 11996 10208 12000
rect 10144 11940 10148 11996
rect 10148 11940 10204 11996
rect 10204 11940 10208 11996
rect 10144 11936 10208 11940
rect 10224 11996 10288 12000
rect 10224 11940 10228 11996
rect 10228 11940 10284 11996
rect 10284 11940 10288 11996
rect 10224 11936 10288 11940
rect 10304 11996 10368 12000
rect 10304 11940 10308 11996
rect 10308 11940 10364 11996
rect 10364 11940 10368 11996
rect 10304 11936 10368 11940
rect 980 11732 1044 11796
rect 2820 11792 2884 11796
rect 2820 11736 2834 11792
rect 2834 11736 2884 11792
rect 2820 11732 2884 11736
rect 8524 11596 8588 11660
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 10724 11452 10788 11456
rect 10724 11396 10728 11452
rect 10728 11396 10784 11452
rect 10784 11396 10788 11452
rect 10724 11392 10788 11396
rect 10804 11452 10868 11456
rect 10804 11396 10808 11452
rect 10808 11396 10864 11452
rect 10864 11396 10868 11452
rect 10804 11392 10868 11396
rect 10884 11452 10948 11456
rect 10884 11396 10888 11452
rect 10888 11396 10944 11452
rect 10944 11396 10948 11452
rect 10884 11392 10948 11396
rect 10964 11452 11028 11456
rect 10964 11396 10968 11452
rect 10968 11396 11024 11452
rect 11024 11396 11028 11452
rect 10964 11392 11028 11396
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 10064 10908 10128 10912
rect 10064 10852 10068 10908
rect 10068 10852 10124 10908
rect 10124 10852 10128 10908
rect 10064 10848 10128 10852
rect 10144 10908 10208 10912
rect 10144 10852 10148 10908
rect 10148 10852 10204 10908
rect 10204 10852 10208 10908
rect 10144 10848 10208 10852
rect 10224 10908 10288 10912
rect 10224 10852 10228 10908
rect 10228 10852 10284 10908
rect 10284 10852 10288 10908
rect 10224 10848 10288 10852
rect 10304 10908 10368 10912
rect 10304 10852 10308 10908
rect 10308 10852 10364 10908
rect 10364 10852 10368 10908
rect 10304 10848 10368 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 10724 10364 10788 10368
rect 10724 10308 10728 10364
rect 10728 10308 10784 10364
rect 10784 10308 10788 10364
rect 10724 10304 10788 10308
rect 10804 10364 10868 10368
rect 10804 10308 10808 10364
rect 10808 10308 10864 10364
rect 10864 10308 10868 10364
rect 10804 10304 10868 10308
rect 10884 10364 10948 10368
rect 10884 10308 10888 10364
rect 10888 10308 10944 10364
rect 10944 10308 10948 10364
rect 10884 10304 10948 10308
rect 10964 10364 11028 10368
rect 10964 10308 10968 10364
rect 10968 10308 11024 10364
rect 11024 10308 11028 10364
rect 10964 10304 11028 10308
rect 4108 10100 4172 10164
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 10064 9820 10128 9824
rect 10064 9764 10068 9820
rect 10068 9764 10124 9820
rect 10124 9764 10128 9820
rect 10064 9760 10128 9764
rect 10144 9820 10208 9824
rect 10144 9764 10148 9820
rect 10148 9764 10204 9820
rect 10204 9764 10208 9820
rect 10144 9760 10208 9764
rect 10224 9820 10288 9824
rect 10224 9764 10228 9820
rect 10228 9764 10284 9820
rect 10284 9764 10288 9820
rect 10224 9760 10288 9764
rect 10304 9820 10368 9824
rect 10304 9764 10308 9820
rect 10308 9764 10364 9820
rect 10364 9764 10368 9820
rect 10304 9760 10368 9764
rect 11284 9420 11348 9484
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 10724 9276 10788 9280
rect 10724 9220 10728 9276
rect 10728 9220 10784 9276
rect 10784 9220 10788 9276
rect 10724 9216 10788 9220
rect 10804 9276 10868 9280
rect 10804 9220 10808 9276
rect 10808 9220 10864 9276
rect 10864 9220 10868 9276
rect 10804 9216 10868 9220
rect 10884 9276 10948 9280
rect 10884 9220 10888 9276
rect 10888 9220 10944 9276
rect 10944 9220 10948 9276
rect 10884 9216 10948 9220
rect 10964 9276 11028 9280
rect 10964 9220 10968 9276
rect 10968 9220 11024 9276
rect 11024 9220 11028 9276
rect 10964 9216 11028 9220
rect 2084 9012 2148 9076
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 10064 8732 10128 8736
rect 10064 8676 10068 8732
rect 10068 8676 10124 8732
rect 10124 8676 10128 8732
rect 10064 8672 10128 8676
rect 10144 8732 10208 8736
rect 10144 8676 10148 8732
rect 10148 8676 10204 8732
rect 10204 8676 10208 8732
rect 10144 8672 10208 8676
rect 10224 8732 10288 8736
rect 10224 8676 10228 8732
rect 10228 8676 10284 8732
rect 10284 8676 10288 8732
rect 10224 8672 10288 8676
rect 10304 8732 10368 8736
rect 10304 8676 10308 8732
rect 10308 8676 10364 8732
rect 10364 8676 10368 8732
rect 10304 8672 10368 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 10724 8188 10788 8192
rect 10724 8132 10728 8188
rect 10728 8132 10784 8188
rect 10784 8132 10788 8188
rect 10724 8128 10788 8132
rect 10804 8188 10868 8192
rect 10804 8132 10808 8188
rect 10808 8132 10864 8188
rect 10864 8132 10868 8188
rect 10804 8128 10868 8132
rect 10884 8188 10948 8192
rect 10884 8132 10888 8188
rect 10888 8132 10944 8188
rect 10944 8132 10948 8188
rect 10884 8128 10948 8132
rect 10964 8188 11028 8192
rect 10964 8132 10968 8188
rect 10968 8132 11024 8188
rect 11024 8132 11028 8188
rect 10964 8128 11028 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 10064 7644 10128 7648
rect 10064 7588 10068 7644
rect 10068 7588 10124 7644
rect 10124 7588 10128 7644
rect 10064 7584 10128 7588
rect 10144 7644 10208 7648
rect 10144 7588 10148 7644
rect 10148 7588 10204 7644
rect 10204 7588 10208 7644
rect 10144 7584 10208 7588
rect 10224 7644 10288 7648
rect 10224 7588 10228 7644
rect 10228 7588 10284 7644
rect 10284 7588 10288 7644
rect 10224 7584 10288 7588
rect 10304 7644 10368 7648
rect 10304 7588 10308 7644
rect 10308 7588 10364 7644
rect 10364 7588 10368 7644
rect 10304 7584 10368 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 10724 7100 10788 7104
rect 10724 7044 10728 7100
rect 10728 7044 10784 7100
rect 10784 7044 10788 7100
rect 10724 7040 10788 7044
rect 10804 7100 10868 7104
rect 10804 7044 10808 7100
rect 10808 7044 10864 7100
rect 10864 7044 10868 7100
rect 10804 7040 10868 7044
rect 10884 7100 10948 7104
rect 10884 7044 10888 7100
rect 10888 7044 10944 7100
rect 10944 7044 10948 7100
rect 10884 7040 10948 7044
rect 10964 7100 11028 7104
rect 10964 7044 10968 7100
rect 10968 7044 11024 7100
rect 11024 7044 11028 7100
rect 10964 7040 11028 7044
rect 7052 6700 7116 6764
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 10064 6556 10128 6560
rect 10064 6500 10068 6556
rect 10068 6500 10124 6556
rect 10124 6500 10128 6556
rect 10064 6496 10128 6500
rect 10144 6556 10208 6560
rect 10144 6500 10148 6556
rect 10148 6500 10204 6556
rect 10204 6500 10208 6556
rect 10144 6496 10208 6500
rect 10224 6556 10288 6560
rect 10224 6500 10228 6556
rect 10228 6500 10284 6556
rect 10284 6500 10288 6556
rect 10224 6496 10288 6500
rect 10304 6556 10368 6560
rect 10304 6500 10308 6556
rect 10308 6500 10364 6556
rect 10364 6500 10368 6556
rect 10304 6496 10368 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 10724 6012 10788 6016
rect 10724 5956 10728 6012
rect 10728 5956 10784 6012
rect 10784 5956 10788 6012
rect 10724 5952 10788 5956
rect 10804 6012 10868 6016
rect 10804 5956 10808 6012
rect 10808 5956 10864 6012
rect 10864 5956 10868 6012
rect 10804 5952 10868 5956
rect 10884 6012 10948 6016
rect 10884 5956 10888 6012
rect 10888 5956 10944 6012
rect 10944 5956 10948 6012
rect 10884 5952 10948 5956
rect 10964 6012 11028 6016
rect 10964 5956 10968 6012
rect 10968 5956 11024 6012
rect 11024 5956 11028 6012
rect 10964 5952 11028 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 10064 5468 10128 5472
rect 10064 5412 10068 5468
rect 10068 5412 10124 5468
rect 10124 5412 10128 5468
rect 10064 5408 10128 5412
rect 10144 5468 10208 5472
rect 10144 5412 10148 5468
rect 10148 5412 10204 5468
rect 10204 5412 10208 5468
rect 10144 5408 10208 5412
rect 10224 5468 10288 5472
rect 10224 5412 10228 5468
rect 10228 5412 10284 5468
rect 10284 5412 10288 5468
rect 10224 5408 10288 5412
rect 10304 5468 10368 5472
rect 10304 5412 10308 5468
rect 10308 5412 10364 5468
rect 10364 5412 10368 5468
rect 10304 5408 10368 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 10724 4924 10788 4928
rect 10724 4868 10728 4924
rect 10728 4868 10784 4924
rect 10784 4868 10788 4924
rect 10724 4864 10788 4868
rect 10804 4924 10868 4928
rect 10804 4868 10808 4924
rect 10808 4868 10864 4924
rect 10864 4868 10868 4924
rect 10804 4864 10868 4868
rect 10884 4924 10948 4928
rect 10884 4868 10888 4924
rect 10888 4868 10944 4924
rect 10944 4868 10948 4924
rect 10884 4864 10948 4868
rect 10964 4924 11028 4928
rect 10964 4868 10968 4924
rect 10968 4868 11024 4924
rect 11024 4868 11028 4924
rect 10964 4864 11028 4868
rect 612 4660 676 4724
rect 60 4388 124 4452
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 10064 4380 10128 4384
rect 10064 4324 10068 4380
rect 10068 4324 10124 4380
rect 10124 4324 10128 4380
rect 10064 4320 10128 4324
rect 10144 4380 10208 4384
rect 10144 4324 10148 4380
rect 10148 4324 10204 4380
rect 10204 4324 10208 4380
rect 10144 4320 10208 4324
rect 10224 4380 10288 4384
rect 10224 4324 10228 4380
rect 10228 4324 10284 4380
rect 10284 4324 10288 4380
rect 10224 4320 10288 4324
rect 10304 4380 10368 4384
rect 10304 4324 10308 4380
rect 10308 4324 10364 4380
rect 10364 4324 10368 4380
rect 10304 4320 10368 4324
rect 6868 3980 6932 4044
rect 8892 4040 8956 4044
rect 8892 3984 8942 4040
rect 8942 3984 8956 4040
rect 8892 3980 8956 3984
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 10724 3836 10788 3840
rect 10724 3780 10728 3836
rect 10728 3780 10784 3836
rect 10784 3780 10788 3836
rect 10724 3776 10788 3780
rect 10804 3836 10868 3840
rect 10804 3780 10808 3836
rect 10808 3780 10864 3836
rect 10864 3780 10868 3836
rect 10804 3776 10868 3780
rect 10884 3836 10948 3840
rect 10884 3780 10888 3836
rect 10888 3780 10944 3836
rect 10944 3780 10948 3836
rect 10884 3776 10948 3780
rect 10964 3836 11028 3840
rect 10964 3780 10968 3836
rect 10968 3780 11024 3836
rect 11024 3780 11028 3836
rect 10964 3776 11028 3780
rect 9076 3768 9140 3772
rect 9076 3712 9126 3768
rect 9126 3712 9140 3768
rect 9076 3708 9140 3712
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 10064 3292 10128 3296
rect 10064 3236 10068 3292
rect 10068 3236 10124 3292
rect 10124 3236 10128 3292
rect 10064 3232 10128 3236
rect 10144 3292 10208 3296
rect 10144 3236 10148 3292
rect 10148 3236 10204 3292
rect 10204 3236 10208 3292
rect 10144 3232 10208 3236
rect 10224 3292 10288 3296
rect 10224 3236 10228 3292
rect 10228 3236 10284 3292
rect 10284 3236 10288 3292
rect 10224 3232 10288 3236
rect 10304 3292 10368 3296
rect 10304 3236 10308 3292
rect 10308 3236 10364 3292
rect 10364 3236 10368 3292
rect 10304 3232 10368 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 10724 2748 10788 2752
rect 10724 2692 10728 2748
rect 10728 2692 10784 2748
rect 10784 2692 10788 2748
rect 10724 2688 10788 2692
rect 10804 2748 10868 2752
rect 10804 2692 10808 2748
rect 10808 2692 10864 2748
rect 10864 2692 10868 2748
rect 10804 2688 10868 2692
rect 10884 2748 10948 2752
rect 10884 2692 10888 2748
rect 10888 2692 10944 2748
rect 10944 2692 10948 2748
rect 10884 2688 10948 2692
rect 10964 2748 11028 2752
rect 10964 2692 10968 2748
rect 10968 2692 11024 2748
rect 11024 2692 11028 2748
rect 10964 2688 11028 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 10064 2204 10128 2208
rect 10064 2148 10068 2204
rect 10068 2148 10124 2204
rect 10124 2148 10128 2204
rect 10064 2144 10128 2148
rect 10144 2204 10208 2208
rect 10144 2148 10148 2204
rect 10148 2148 10204 2204
rect 10204 2148 10208 2204
rect 10144 2144 10208 2148
rect 10224 2204 10288 2208
rect 10224 2148 10228 2204
rect 10228 2148 10284 2204
rect 10284 2148 10288 2204
rect 10224 2144 10288 2148
rect 10304 2204 10368 2208
rect 10304 2148 10308 2204
rect 10308 2148 10364 2204
rect 10364 2148 10368 2204
rect 10304 2144 10368 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 10724 1660 10788 1664
rect 10724 1604 10728 1660
rect 10728 1604 10784 1660
rect 10784 1604 10788 1660
rect 10724 1600 10788 1604
rect 10804 1660 10868 1664
rect 10804 1604 10808 1660
rect 10808 1604 10864 1660
rect 10864 1604 10868 1660
rect 10804 1600 10868 1604
rect 10884 1660 10948 1664
rect 10884 1604 10888 1660
rect 10888 1604 10944 1660
rect 10944 1604 10948 1660
rect 10884 1600 10948 1604
rect 10964 1660 11028 1664
rect 10964 1604 10968 1660
rect 10968 1604 11024 1660
rect 11024 1604 11028 1660
rect 10964 1600 11028 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 10064 1116 10128 1120
rect 10064 1060 10068 1116
rect 10068 1060 10124 1116
rect 10124 1060 10128 1116
rect 10064 1056 10128 1060
rect 10144 1116 10208 1120
rect 10144 1060 10148 1116
rect 10148 1060 10204 1116
rect 10204 1060 10208 1116
rect 10144 1056 10208 1060
rect 10224 1116 10288 1120
rect 10224 1060 10228 1116
rect 10228 1060 10284 1116
rect 10284 1060 10288 1116
rect 10224 1056 10288 1060
rect 10304 1116 10368 1120
rect 10304 1060 10308 1116
rect 10308 1060 10364 1116
rect 10364 1060 10368 1116
rect 10304 1056 10368 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
rect 10724 572 10788 576
rect 10724 516 10728 572
rect 10728 516 10784 572
rect 10784 516 10788 572
rect 10724 512 10788 516
rect 10804 572 10868 576
rect 10804 516 10808 572
rect 10808 516 10864 572
rect 10864 516 10868 572
rect 10804 512 10868 516
rect 10884 572 10948 576
rect 10884 516 10888 572
rect 10888 516 10944 572
rect 10944 516 10948 572
rect 10884 512 10948 516
rect 10964 572 11028 576
rect 10964 516 10968 572
rect 10968 516 11024 572
rect 11024 516 11028 572
rect 10964 512 11028 516
<< metal4 >>
rect 979 43620 1045 43621
rect 979 43556 980 43620
rect 1044 43556 1045 43620
rect 979 43555 1045 43556
rect 7787 43620 7853 43621
rect 7787 43556 7788 43620
rect 7852 43556 7853 43620
rect 7787 43555 7853 43556
rect 381 37092 447 37093
rect 381 37090 382 37092
rect 62 37030 382 37090
rect 62 20501 122 37030
rect 381 37028 382 37030
rect 446 37028 447 37092
rect 381 37027 447 37028
rect 427 35188 493 35189
rect 427 35124 428 35188
rect 492 35124 493 35188
rect 427 35123 493 35124
rect 243 29612 309 29613
rect 243 29548 244 29612
rect 308 29548 309 29612
rect 243 29547 309 29548
rect 246 27845 306 29547
rect 243 27844 309 27845
rect 243 27780 244 27844
rect 308 27780 309 27844
rect 243 27779 309 27780
rect 243 27572 309 27573
rect 243 27508 244 27572
rect 308 27508 309 27572
rect 243 27507 309 27508
rect 59 20500 125 20501
rect 59 20436 60 20500
rect 124 20436 125 20500
rect 59 20435 125 20436
rect 59 17916 125 17917
rect 59 17852 60 17916
rect 124 17852 125 17916
rect 59 17851 125 17852
rect 62 4453 122 17851
rect 246 17509 306 27507
rect 430 22405 490 35123
rect 982 35053 1042 43555
rect 3656 42464 3976 43024
rect 3656 42400 3664 42464
rect 3728 42400 3744 42464
rect 3808 42400 3824 42464
rect 3888 42400 3904 42464
rect 3968 42400 3976 42464
rect 1163 41580 1229 41581
rect 1163 41516 1164 41580
rect 1228 41516 1229 41580
rect 1163 41515 1229 41516
rect 979 35052 1045 35053
rect 979 34988 980 35052
rect 1044 34988 1045 35052
rect 979 34987 1045 34988
rect 979 33012 1045 33013
rect 979 32948 980 33012
rect 1044 32948 1045 33012
rect 979 32947 1045 32948
rect 611 30428 677 30429
rect 611 30364 612 30428
rect 676 30364 677 30428
rect 611 30363 677 30364
rect 614 27437 674 30363
rect 982 29474 1042 32947
rect 1166 29610 1226 41515
rect 3656 41376 3976 42400
rect 3656 41312 3664 41376
rect 3728 41312 3744 41376
rect 3808 41312 3824 41376
rect 3888 41312 3904 41376
rect 3968 41312 3976 41376
rect 2635 41172 2701 41173
rect 2635 41108 2636 41172
rect 2700 41108 2701 41172
rect 2635 41107 2701 41108
rect 1899 40220 1965 40221
rect 1899 40156 1900 40220
rect 1964 40156 1965 40220
rect 1899 40155 1965 40156
rect 1347 37364 1413 37365
rect 1347 37300 1348 37364
rect 1412 37300 1413 37364
rect 1347 37299 1413 37300
rect 1350 30429 1410 37299
rect 1902 35189 1962 40155
rect 2083 39948 2149 39949
rect 2083 39884 2084 39948
rect 2148 39884 2149 39948
rect 2083 39883 2149 39884
rect 2086 39405 2146 39883
rect 2083 39404 2149 39405
rect 2083 39340 2084 39404
rect 2148 39340 2149 39404
rect 2083 39339 2149 39340
rect 1899 35188 1965 35189
rect 1899 35124 1900 35188
rect 1964 35124 1965 35188
rect 1899 35123 1965 35124
rect 1899 34780 1965 34781
rect 1899 34716 1900 34780
rect 1964 34716 1965 34780
rect 1899 34715 1965 34716
rect 1531 33284 1597 33285
rect 1531 33220 1532 33284
rect 1596 33220 1597 33284
rect 1531 33219 1597 33220
rect 1534 31381 1594 33219
rect 1715 31652 1781 31653
rect 1715 31588 1716 31652
rect 1780 31588 1781 31652
rect 1715 31587 1781 31588
rect 1531 31380 1597 31381
rect 1531 31316 1532 31380
rect 1596 31316 1597 31380
rect 1531 31315 1597 31316
rect 1718 31109 1778 31587
rect 1715 31108 1781 31109
rect 1715 31044 1716 31108
rect 1780 31044 1781 31108
rect 1715 31043 1781 31044
rect 1347 30428 1413 30429
rect 1347 30364 1348 30428
rect 1412 30364 1413 30428
rect 1347 30363 1413 30364
rect 1347 29612 1413 29613
rect 1347 29610 1348 29612
rect 1166 29550 1348 29610
rect 1347 29548 1348 29550
rect 1412 29548 1413 29612
rect 1347 29547 1413 29548
rect 982 29414 1226 29474
rect 979 29340 1045 29341
rect 979 29276 980 29340
rect 1044 29276 1045 29340
rect 979 29275 1045 29276
rect 795 28796 861 28797
rect 795 28732 796 28796
rect 860 28732 861 28796
rect 795 28731 861 28732
rect 611 27436 677 27437
rect 611 27372 612 27436
rect 676 27372 677 27436
rect 611 27371 677 27372
rect 427 22404 493 22405
rect 427 22340 428 22404
rect 492 22340 493 22404
rect 427 22339 493 22340
rect 614 18730 674 27371
rect 798 22269 858 28731
rect 795 22268 861 22269
rect 795 22204 796 22268
rect 860 22204 861 22268
rect 795 22203 861 22204
rect 982 22133 1042 29275
rect 1166 27981 1226 29414
rect 1163 27980 1229 27981
rect 1163 27916 1164 27980
rect 1228 27916 1229 27980
rect 1163 27915 1229 27916
rect 1163 27844 1229 27845
rect 1163 27780 1164 27844
rect 1228 27780 1229 27844
rect 1163 27779 1229 27780
rect 1166 23629 1226 27779
rect 1350 26213 1410 29547
rect 1531 29068 1597 29069
rect 1531 29004 1532 29068
rect 1596 29004 1597 29068
rect 1531 29003 1597 29004
rect 1347 26212 1413 26213
rect 1347 26148 1348 26212
rect 1412 26148 1413 26212
rect 1347 26147 1413 26148
rect 1534 25941 1594 29003
rect 1718 26077 1778 31043
rect 1902 27029 1962 34715
rect 2086 30293 2146 39339
rect 2451 34916 2517 34917
rect 2451 34852 2452 34916
rect 2516 34852 2517 34916
rect 2451 34851 2517 34852
rect 2267 33148 2333 33149
rect 2267 33084 2268 33148
rect 2332 33084 2333 33148
rect 2267 33083 2333 33084
rect 2270 31925 2330 33083
rect 2267 31924 2333 31925
rect 2267 31860 2268 31924
rect 2332 31860 2333 31924
rect 2267 31859 2333 31860
rect 2083 30292 2149 30293
rect 2083 30228 2084 30292
rect 2148 30228 2149 30292
rect 2083 30227 2149 30228
rect 2454 29749 2514 34851
rect 2638 33690 2698 41107
rect 3371 41036 3437 41037
rect 3371 40972 3372 41036
rect 3436 40972 3437 41036
rect 3371 40971 3437 40972
rect 3374 37909 3434 40971
rect 3656 40288 3976 41312
rect 3656 40224 3664 40288
rect 3728 40224 3744 40288
rect 3808 40224 3824 40288
rect 3888 40224 3904 40288
rect 3968 40224 3976 40288
rect 3656 39200 3976 40224
rect 4316 43008 4636 43024
rect 4316 42944 4324 43008
rect 4388 42944 4404 43008
rect 4468 42944 4484 43008
rect 4548 42944 4564 43008
rect 4628 42944 4636 43008
rect 4316 41920 4636 42944
rect 5579 42260 5645 42261
rect 5579 42196 5580 42260
rect 5644 42196 5645 42260
rect 5579 42195 5645 42196
rect 5211 42124 5277 42125
rect 5211 42060 5212 42124
rect 5276 42060 5277 42124
rect 5211 42059 5277 42060
rect 4316 41856 4324 41920
rect 4388 41856 4404 41920
rect 4468 41856 4484 41920
rect 4548 41856 4564 41920
rect 4628 41856 4636 41920
rect 4316 40832 4636 41856
rect 4316 40768 4324 40832
rect 4388 40768 4404 40832
rect 4468 40768 4484 40832
rect 4548 40768 4564 40832
rect 4628 40768 4636 40832
rect 4107 40084 4173 40085
rect 4107 40020 4108 40084
rect 4172 40020 4173 40084
rect 4107 40019 4173 40020
rect 3656 39136 3664 39200
rect 3728 39136 3744 39200
rect 3808 39136 3824 39200
rect 3888 39136 3904 39200
rect 3968 39136 3976 39200
rect 3656 38112 3976 39136
rect 3656 38048 3664 38112
rect 3728 38048 3744 38112
rect 3808 38048 3824 38112
rect 3888 38048 3904 38112
rect 3968 38048 3976 38112
rect 3371 37908 3437 37909
rect 3371 37844 3372 37908
rect 3436 37844 3437 37908
rect 3371 37843 3437 37844
rect 3187 36412 3253 36413
rect 3187 36348 3188 36412
rect 3252 36348 3253 36412
rect 3187 36347 3253 36348
rect 2638 33630 2882 33690
rect 2635 30292 2701 30293
rect 2635 30228 2636 30292
rect 2700 30228 2701 30292
rect 2635 30227 2701 30228
rect 2083 29748 2149 29749
rect 2083 29684 2084 29748
rect 2148 29684 2149 29748
rect 2083 29683 2149 29684
rect 2451 29748 2517 29749
rect 2451 29684 2452 29748
rect 2516 29684 2517 29748
rect 2451 29683 2517 29684
rect 2086 28389 2146 29683
rect 2451 29204 2517 29205
rect 2451 29140 2452 29204
rect 2516 29140 2517 29204
rect 2451 29139 2517 29140
rect 2267 28796 2333 28797
rect 2267 28732 2268 28796
rect 2332 28732 2333 28796
rect 2267 28731 2333 28732
rect 2083 28388 2149 28389
rect 2083 28324 2084 28388
rect 2148 28324 2149 28388
rect 2083 28323 2149 28324
rect 2083 28252 2149 28253
rect 2083 28188 2084 28252
rect 2148 28188 2149 28252
rect 2083 28187 2149 28188
rect 1899 27028 1965 27029
rect 1899 26964 1900 27028
rect 1964 26964 1965 27028
rect 1899 26963 1965 26964
rect 2086 26485 2146 28187
rect 2083 26484 2149 26485
rect 2083 26420 2084 26484
rect 2148 26420 2149 26484
rect 2083 26419 2149 26420
rect 1715 26076 1781 26077
rect 1715 26012 1716 26076
rect 1780 26012 1781 26076
rect 1715 26011 1781 26012
rect 1531 25940 1597 25941
rect 1531 25876 1532 25940
rect 1596 25876 1597 25940
rect 1531 25875 1597 25876
rect 1715 25940 1781 25941
rect 1715 25876 1716 25940
rect 1780 25876 1781 25940
rect 1715 25875 1781 25876
rect 1347 25804 1413 25805
rect 1347 25740 1348 25804
rect 1412 25740 1413 25804
rect 1347 25739 1413 25740
rect 1350 24173 1410 25739
rect 1531 24580 1597 24581
rect 1531 24516 1532 24580
rect 1596 24516 1597 24580
rect 1531 24515 1597 24516
rect 1347 24172 1413 24173
rect 1347 24108 1348 24172
rect 1412 24108 1413 24172
rect 1347 24107 1413 24108
rect 1163 23628 1229 23629
rect 1163 23564 1164 23628
rect 1228 23564 1229 23628
rect 1163 23563 1229 23564
rect 1347 23492 1413 23493
rect 1347 23428 1348 23492
rect 1412 23428 1413 23492
rect 1347 23427 1413 23428
rect 1163 23084 1229 23085
rect 1163 23020 1164 23084
rect 1228 23020 1229 23084
rect 1163 23019 1229 23020
rect 979 22132 1045 22133
rect 979 22068 980 22132
rect 1044 22068 1045 22132
rect 979 22067 1045 22068
rect 979 20636 1045 20637
rect 979 20572 980 20636
rect 1044 20572 1045 20636
rect 979 20571 1045 20572
rect 614 18670 858 18730
rect 611 18052 677 18053
rect 611 17988 612 18052
rect 676 17988 677 18052
rect 611 17987 677 17988
rect 243 17508 309 17509
rect 243 17444 244 17508
rect 308 17444 309 17508
rect 243 17443 309 17444
rect 614 4725 674 17987
rect 798 16421 858 18670
rect 795 16420 861 16421
rect 795 16356 796 16420
rect 860 16356 861 16420
rect 795 16355 861 16356
rect 982 11797 1042 20571
rect 1166 12069 1226 23019
rect 1350 17101 1410 23427
rect 1534 21181 1594 24515
rect 1718 23493 1778 25875
rect 1899 25804 1965 25805
rect 1899 25740 1900 25804
rect 1964 25740 1965 25804
rect 1899 25739 1965 25740
rect 1902 24309 1962 25739
rect 2083 25396 2149 25397
rect 2083 25332 2084 25396
rect 2148 25332 2149 25396
rect 2083 25331 2149 25332
rect 1899 24308 1965 24309
rect 1899 24244 1900 24308
rect 1964 24244 1965 24308
rect 1899 24243 1965 24244
rect 1899 24172 1965 24173
rect 1899 24108 1900 24172
rect 1964 24108 1965 24172
rect 1899 24107 1965 24108
rect 1715 23492 1781 23493
rect 1715 23428 1716 23492
rect 1780 23428 1781 23492
rect 1715 23427 1781 23428
rect 1715 23356 1781 23357
rect 1715 23292 1716 23356
rect 1780 23292 1781 23356
rect 1715 23291 1781 23292
rect 1531 21180 1597 21181
rect 1531 21116 1532 21180
rect 1596 21116 1597 21180
rect 1531 21115 1597 21116
rect 1531 17236 1597 17237
rect 1531 17172 1532 17236
rect 1596 17172 1597 17236
rect 1531 17171 1597 17172
rect 1347 17100 1413 17101
rect 1347 17036 1348 17100
rect 1412 17036 1413 17100
rect 1347 17035 1413 17036
rect 1534 13837 1594 17171
rect 1718 16149 1778 23291
rect 1902 22674 1962 24107
rect 2086 23357 2146 25331
rect 2270 25125 2330 28731
rect 2267 25124 2333 25125
rect 2267 25060 2268 25124
rect 2332 25060 2333 25124
rect 2267 25059 2333 25060
rect 2267 24988 2333 24989
rect 2267 24924 2268 24988
rect 2332 24924 2333 24988
rect 2267 24923 2333 24924
rect 2083 23356 2149 23357
rect 2083 23292 2084 23356
rect 2148 23292 2149 23356
rect 2083 23291 2149 23292
rect 1902 22614 2146 22674
rect 1899 22540 1965 22541
rect 1899 22476 1900 22540
rect 1964 22476 1965 22540
rect 1899 22475 1965 22476
rect 1715 16148 1781 16149
rect 1715 16084 1716 16148
rect 1780 16084 1781 16148
rect 1715 16083 1781 16084
rect 1531 13836 1597 13837
rect 1531 13772 1532 13836
rect 1596 13772 1597 13836
rect 1531 13771 1597 13772
rect 1902 12069 1962 22475
rect 2086 19957 2146 22614
rect 2083 19956 2149 19957
rect 2083 19892 2084 19956
rect 2148 19892 2149 19956
rect 2083 19891 2149 19892
rect 2270 15197 2330 24923
rect 2454 23221 2514 29139
rect 2451 23220 2517 23221
rect 2451 23156 2452 23220
rect 2516 23156 2517 23220
rect 2451 23155 2517 23156
rect 2454 22541 2514 23155
rect 2451 22540 2517 22541
rect 2451 22476 2452 22540
rect 2516 22476 2517 22540
rect 2451 22475 2517 22476
rect 2451 22404 2517 22405
rect 2451 22340 2452 22404
rect 2516 22340 2517 22404
rect 2451 22339 2517 22340
rect 2454 20637 2514 22339
rect 2451 20636 2517 20637
rect 2451 20572 2452 20636
rect 2516 20572 2517 20636
rect 2451 20571 2517 20572
rect 2451 20228 2517 20229
rect 2451 20164 2452 20228
rect 2516 20164 2517 20228
rect 2451 20163 2517 20164
rect 2267 15196 2333 15197
rect 2267 15132 2268 15196
rect 2332 15132 2333 15196
rect 2267 15131 2333 15132
rect 2083 12884 2149 12885
rect 2083 12820 2084 12884
rect 2148 12820 2149 12884
rect 2083 12819 2149 12820
rect 1163 12068 1229 12069
rect 1163 12004 1164 12068
rect 1228 12004 1229 12068
rect 1163 12003 1229 12004
rect 1899 12068 1965 12069
rect 1899 12004 1900 12068
rect 1964 12004 1965 12068
rect 1899 12003 1965 12004
rect 979 11796 1045 11797
rect 979 11732 980 11796
rect 1044 11732 1045 11796
rect 979 11731 1045 11732
rect 2086 9077 2146 12819
rect 2454 12341 2514 20163
rect 2638 19277 2698 30227
rect 2822 29069 2882 33630
rect 3190 29749 3250 36347
rect 3374 34101 3434 37843
rect 3656 37024 3976 38048
rect 3656 36960 3664 37024
rect 3728 36960 3744 37024
rect 3808 36960 3824 37024
rect 3888 36960 3904 37024
rect 3968 36960 3976 37024
rect 3656 35936 3976 36960
rect 3656 35872 3664 35936
rect 3728 35872 3744 35936
rect 3808 35872 3824 35936
rect 3888 35872 3904 35936
rect 3968 35872 3976 35936
rect 3656 34848 3976 35872
rect 3656 34784 3664 34848
rect 3728 34784 3744 34848
rect 3808 34784 3824 34848
rect 3888 34784 3904 34848
rect 3968 34784 3976 34848
rect 3371 34100 3437 34101
rect 3371 34036 3372 34100
rect 3436 34036 3437 34100
rect 3371 34035 3437 34036
rect 3656 33760 3976 34784
rect 4110 34645 4170 40019
rect 4316 39744 4636 40768
rect 4843 40220 4909 40221
rect 4843 40156 4844 40220
rect 4908 40156 4909 40220
rect 4843 40155 4909 40156
rect 4316 39680 4324 39744
rect 4388 39680 4404 39744
rect 4468 39680 4484 39744
rect 4548 39680 4564 39744
rect 4628 39680 4636 39744
rect 4316 38656 4636 39680
rect 4316 38592 4324 38656
rect 4388 38592 4404 38656
rect 4468 38592 4484 38656
rect 4548 38592 4564 38656
rect 4628 38592 4636 38656
rect 4316 37568 4636 38592
rect 4316 37504 4324 37568
rect 4388 37504 4404 37568
rect 4468 37504 4484 37568
rect 4548 37504 4564 37568
rect 4628 37504 4636 37568
rect 4316 36480 4636 37504
rect 4316 36416 4324 36480
rect 4388 36416 4404 36480
rect 4468 36416 4484 36480
rect 4548 36416 4564 36480
rect 4628 36416 4636 36480
rect 4316 35392 4636 36416
rect 4846 36141 4906 40155
rect 5027 38724 5093 38725
rect 5027 38660 5028 38724
rect 5092 38660 5093 38724
rect 5027 38659 5093 38660
rect 4843 36140 4909 36141
rect 4843 36076 4844 36140
rect 4908 36076 4909 36140
rect 4843 36075 4909 36076
rect 4316 35328 4324 35392
rect 4388 35328 4404 35392
rect 4468 35328 4484 35392
rect 4548 35328 4564 35392
rect 4628 35328 4636 35392
rect 4107 34644 4173 34645
rect 4107 34580 4108 34644
rect 4172 34580 4173 34644
rect 4107 34579 4173 34580
rect 3656 33696 3664 33760
rect 3728 33696 3744 33760
rect 3808 33696 3824 33760
rect 3888 33696 3904 33760
rect 3968 33696 3976 33760
rect 3371 33284 3437 33285
rect 3371 33220 3372 33284
rect 3436 33220 3437 33284
rect 3371 33219 3437 33220
rect 3187 29748 3253 29749
rect 3187 29684 3188 29748
rect 3252 29684 3253 29748
rect 3187 29683 3253 29684
rect 3374 29205 3434 33219
rect 3656 32672 3976 33696
rect 3656 32608 3664 32672
rect 3728 32608 3744 32672
rect 3808 32608 3824 32672
rect 3888 32608 3904 32672
rect 3968 32608 3976 32672
rect 3656 31584 3976 32608
rect 3656 31520 3664 31584
rect 3728 31520 3744 31584
rect 3808 31520 3824 31584
rect 3888 31520 3904 31584
rect 3968 31520 3976 31584
rect 3656 30496 3976 31520
rect 3656 30432 3664 30496
rect 3728 30432 3744 30496
rect 3808 30432 3824 30496
rect 3888 30432 3904 30496
rect 3968 30432 3976 30496
rect 3656 29408 3976 30432
rect 4110 30429 4170 34579
rect 4316 34304 4636 35328
rect 4843 34508 4909 34509
rect 4843 34444 4844 34508
rect 4908 34444 4909 34508
rect 4843 34443 4909 34444
rect 4316 34240 4324 34304
rect 4388 34240 4404 34304
rect 4468 34240 4484 34304
rect 4548 34240 4564 34304
rect 4628 34240 4636 34304
rect 4316 33216 4636 34240
rect 4316 33152 4324 33216
rect 4388 33152 4404 33216
rect 4468 33152 4484 33216
rect 4548 33152 4564 33216
rect 4628 33152 4636 33216
rect 4316 32128 4636 33152
rect 4316 32064 4324 32128
rect 4388 32064 4404 32128
rect 4468 32064 4484 32128
rect 4548 32064 4564 32128
rect 4628 32064 4636 32128
rect 4316 31040 4636 32064
rect 4316 30976 4324 31040
rect 4388 30976 4404 31040
rect 4468 30976 4484 31040
rect 4548 30976 4564 31040
rect 4628 30976 4636 31040
rect 4107 30428 4173 30429
rect 4107 30364 4108 30428
rect 4172 30364 4173 30428
rect 4107 30363 4173 30364
rect 4316 29952 4636 30976
rect 4316 29888 4324 29952
rect 4388 29888 4404 29952
rect 4468 29888 4484 29952
rect 4548 29888 4564 29952
rect 4628 29888 4636 29952
rect 4107 29476 4173 29477
rect 4107 29412 4108 29476
rect 4172 29412 4173 29476
rect 4107 29411 4173 29412
rect 3656 29344 3664 29408
rect 3728 29344 3744 29408
rect 3808 29344 3824 29408
rect 3888 29344 3904 29408
rect 3968 29344 3976 29408
rect 3371 29204 3437 29205
rect 3371 29140 3372 29204
rect 3436 29140 3437 29204
rect 3371 29139 3437 29140
rect 2819 29068 2885 29069
rect 2819 29004 2820 29068
rect 2884 29004 2885 29068
rect 2819 29003 2885 29004
rect 3371 28932 3437 28933
rect 3371 28930 3372 28932
rect 3190 28870 3372 28930
rect 2819 28796 2885 28797
rect 2819 28732 2820 28796
rect 2884 28732 2885 28796
rect 2819 28731 2885 28732
rect 2822 22405 2882 28731
rect 3003 28524 3069 28525
rect 3003 28460 3004 28524
rect 3068 28460 3069 28524
rect 3003 28459 3069 28460
rect 3006 28253 3066 28459
rect 3003 28252 3069 28253
rect 3003 28188 3004 28252
rect 3068 28188 3069 28252
rect 3003 28187 3069 28188
rect 3190 27842 3250 28870
rect 3371 28868 3372 28870
rect 3436 28868 3437 28932
rect 3371 28867 3437 28868
rect 3371 28524 3437 28525
rect 3371 28460 3372 28524
rect 3436 28460 3437 28524
rect 3371 28459 3437 28460
rect 3006 27782 3250 27842
rect 3006 25805 3066 27782
rect 3187 27708 3253 27709
rect 3187 27644 3188 27708
rect 3252 27644 3253 27708
rect 3187 27643 3253 27644
rect 3190 26213 3250 27643
rect 3374 26893 3434 28459
rect 3656 28320 3976 29344
rect 4110 28797 4170 29411
rect 4316 28864 4636 29888
rect 4846 29341 4906 34443
rect 4843 29340 4909 29341
rect 4843 29276 4844 29340
rect 4908 29276 4909 29340
rect 4843 29275 4909 29276
rect 4843 29204 4909 29205
rect 4843 29140 4844 29204
rect 4908 29140 4909 29204
rect 4843 29139 4909 29140
rect 4316 28800 4324 28864
rect 4388 28800 4404 28864
rect 4468 28800 4484 28864
rect 4548 28800 4564 28864
rect 4628 28800 4636 28864
rect 4107 28796 4173 28797
rect 4107 28732 4108 28796
rect 4172 28732 4173 28796
rect 4107 28731 4173 28732
rect 4107 28524 4173 28525
rect 4107 28460 4108 28524
rect 4172 28460 4173 28524
rect 4107 28459 4173 28460
rect 3656 28256 3664 28320
rect 3728 28256 3744 28320
rect 3808 28256 3824 28320
rect 3888 28256 3904 28320
rect 3968 28256 3976 28320
rect 3656 27232 3976 28256
rect 3656 27168 3664 27232
rect 3728 27168 3744 27232
rect 3808 27168 3824 27232
rect 3888 27168 3904 27232
rect 3968 27168 3976 27232
rect 3371 26892 3437 26893
rect 3371 26828 3372 26892
rect 3436 26828 3437 26892
rect 3371 26827 3437 26828
rect 3371 26756 3437 26757
rect 3371 26692 3372 26756
rect 3436 26692 3437 26756
rect 3371 26691 3437 26692
rect 3187 26212 3253 26213
rect 3187 26148 3188 26212
rect 3252 26148 3253 26212
rect 3187 26147 3253 26148
rect 3187 26076 3253 26077
rect 3187 26012 3188 26076
rect 3252 26012 3253 26076
rect 3187 26011 3253 26012
rect 3190 25805 3250 26011
rect 3003 25804 3069 25805
rect 3003 25740 3004 25804
rect 3068 25740 3069 25804
rect 3003 25739 3069 25740
rect 3187 25804 3253 25805
rect 3187 25740 3188 25804
rect 3252 25740 3253 25804
rect 3187 25739 3253 25740
rect 3187 25668 3253 25669
rect 3187 25604 3188 25668
rect 3252 25604 3253 25668
rect 3187 25603 3253 25604
rect 3003 25396 3069 25397
rect 3003 25332 3004 25396
rect 3068 25332 3069 25396
rect 3003 25331 3069 25332
rect 2819 22404 2885 22405
rect 2819 22340 2820 22404
rect 2884 22340 2885 22404
rect 2819 22339 2885 22340
rect 2819 22132 2885 22133
rect 2819 22068 2820 22132
rect 2884 22068 2885 22132
rect 2819 22067 2885 22068
rect 2635 19276 2701 19277
rect 2635 19212 2636 19276
rect 2700 19212 2701 19276
rect 2635 19211 2701 19212
rect 2635 18868 2701 18869
rect 2635 18804 2636 18868
rect 2700 18804 2701 18868
rect 2635 18803 2701 18804
rect 2638 16965 2698 18803
rect 2822 18053 2882 22067
rect 2819 18052 2885 18053
rect 2819 17988 2820 18052
rect 2884 17988 2885 18052
rect 2819 17987 2885 17988
rect 2635 16964 2701 16965
rect 2635 16900 2636 16964
rect 2700 16900 2701 16964
rect 2635 16899 2701 16900
rect 3006 16010 3066 25331
rect 3190 22405 3250 25603
rect 3374 25261 3434 26691
rect 3656 26144 3976 27168
rect 3656 26080 3664 26144
rect 3728 26080 3744 26144
rect 3808 26080 3824 26144
rect 3888 26080 3904 26144
rect 3968 26080 3976 26144
rect 3371 25260 3437 25261
rect 3371 25196 3372 25260
rect 3436 25196 3437 25260
rect 3371 25195 3437 25196
rect 3187 22404 3253 22405
rect 3187 22340 3188 22404
rect 3252 22340 3253 22404
rect 3187 22339 3253 22340
rect 3187 21860 3253 21861
rect 3187 21796 3188 21860
rect 3252 21796 3253 21860
rect 3187 21795 3253 21796
rect 3190 16149 3250 21795
rect 3374 16829 3434 25195
rect 3656 25056 3976 26080
rect 3656 24992 3664 25056
rect 3728 24992 3744 25056
rect 3808 24992 3824 25056
rect 3888 24992 3904 25056
rect 3968 24992 3976 25056
rect 3656 23968 3976 24992
rect 3656 23904 3664 23968
rect 3728 23904 3744 23968
rect 3808 23904 3824 23968
rect 3888 23904 3904 23968
rect 3968 23904 3976 23968
rect 3656 22880 3976 23904
rect 4110 22949 4170 28459
rect 4316 27776 4636 28800
rect 4316 27712 4324 27776
rect 4388 27712 4404 27776
rect 4468 27712 4484 27776
rect 4548 27712 4564 27776
rect 4628 27712 4636 27776
rect 4316 26688 4636 27712
rect 4316 26624 4324 26688
rect 4388 26624 4404 26688
rect 4468 26624 4484 26688
rect 4548 26624 4564 26688
rect 4628 26624 4636 26688
rect 4316 25600 4636 26624
rect 4846 26349 4906 29139
rect 5030 29066 5090 38659
rect 5214 34509 5274 42059
rect 5582 38453 5642 42195
rect 6683 41716 6749 41717
rect 6683 41652 6684 41716
rect 6748 41652 6749 41716
rect 6683 41651 6749 41652
rect 6686 41430 6746 41651
rect 6686 41370 6930 41430
rect 5947 40084 6013 40085
rect 5947 40020 5948 40084
rect 6012 40020 6013 40084
rect 5947 40019 6013 40020
rect 6499 40084 6565 40085
rect 6499 40020 6500 40084
rect 6564 40020 6565 40084
rect 6499 40019 6565 40020
rect 5579 38452 5645 38453
rect 5579 38388 5580 38452
rect 5644 38388 5645 38452
rect 5579 38387 5645 38388
rect 5582 37093 5642 38387
rect 5579 37092 5645 37093
rect 5579 37028 5580 37092
rect 5644 37028 5645 37092
rect 5579 37027 5645 37028
rect 5395 36820 5461 36821
rect 5395 36756 5396 36820
rect 5460 36756 5461 36820
rect 5395 36755 5461 36756
rect 5398 35053 5458 36755
rect 5395 35052 5461 35053
rect 5395 34988 5396 35052
rect 5460 34988 5461 35052
rect 5395 34987 5461 34988
rect 5211 34508 5277 34509
rect 5211 34444 5212 34508
rect 5276 34444 5277 34508
rect 5211 34443 5277 34444
rect 5395 34100 5461 34101
rect 5395 34036 5396 34100
rect 5460 34036 5461 34100
rect 5395 34035 5461 34036
rect 5211 31788 5277 31789
rect 5211 31724 5212 31788
rect 5276 31724 5277 31788
rect 5211 31723 5277 31724
rect 5214 29205 5274 31723
rect 5211 29204 5277 29205
rect 5211 29140 5212 29204
rect 5276 29140 5277 29204
rect 5211 29139 5277 29140
rect 5030 29006 5274 29066
rect 5027 28932 5093 28933
rect 5027 28868 5028 28932
rect 5092 28868 5093 28932
rect 5027 28867 5093 28868
rect 4843 26348 4909 26349
rect 4843 26284 4844 26348
rect 4908 26284 4909 26348
rect 4843 26283 4909 26284
rect 4705 26212 4771 26213
rect 4705 26148 4706 26212
rect 4770 26148 4771 26212
rect 4705 26147 4771 26148
rect 4316 25536 4324 25600
rect 4388 25536 4404 25600
rect 4468 25536 4484 25600
rect 4548 25536 4564 25600
rect 4628 25536 4636 25600
rect 4316 24512 4636 25536
rect 4708 24581 4768 26147
rect 4705 24580 4771 24581
rect 4705 24516 4706 24580
rect 4770 24516 4771 24580
rect 4705 24515 4771 24516
rect 4316 24448 4324 24512
rect 4388 24448 4404 24512
rect 4468 24448 4484 24512
rect 4548 24448 4564 24512
rect 4628 24448 4636 24512
rect 4316 23424 4636 24448
rect 4316 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4636 23424
rect 4107 22948 4173 22949
rect 4107 22884 4108 22948
rect 4172 22884 4173 22948
rect 4107 22883 4173 22884
rect 3656 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3976 22880
rect 3656 21792 3976 22816
rect 4107 22812 4173 22813
rect 4107 22748 4108 22812
rect 4172 22748 4173 22812
rect 4107 22747 4173 22748
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 4110 20229 4170 22747
rect 4316 22336 4636 23360
rect 4316 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4636 22336
rect 4316 21248 4636 22272
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4107 20228 4173 20229
rect 4107 20164 4108 20228
rect 4172 20164 4173 20228
rect 4107 20163 4173 20164
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 4316 20160 4636 21184
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4107 18188 4173 18189
rect 4107 18124 4108 18188
rect 4172 18124 4173 18188
rect 4107 18123 4173 18124
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3371 16828 3437 16829
rect 3371 16764 3372 16828
rect 3436 16764 3437 16828
rect 3371 16763 3437 16764
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3187 16148 3253 16149
rect 3187 16084 3188 16148
rect 3252 16084 3253 16148
rect 3187 16083 3253 16084
rect 2822 15950 3066 16010
rect 2822 14653 2882 15950
rect 3003 15876 3069 15877
rect 3003 15812 3004 15876
rect 3068 15812 3069 15876
rect 3003 15811 3069 15812
rect 2819 14652 2885 14653
rect 2819 14588 2820 14652
rect 2884 14588 2885 14652
rect 2819 14587 2885 14588
rect 3006 13701 3066 15811
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 4110 15197 4170 18123
rect 4316 17984 4636 19008
rect 4846 18325 4906 26283
rect 5030 20773 5090 28867
rect 5214 27437 5274 29006
rect 5211 27436 5277 27437
rect 5211 27372 5212 27436
rect 5276 27372 5277 27436
rect 5211 27371 5277 27372
rect 5211 27300 5277 27301
rect 5211 27236 5212 27300
rect 5276 27236 5277 27300
rect 5211 27235 5277 27236
rect 5214 25261 5274 27235
rect 5211 25260 5277 25261
rect 5211 25196 5212 25260
rect 5276 25196 5277 25260
rect 5211 25195 5277 25196
rect 5211 24444 5277 24445
rect 5211 24380 5212 24444
rect 5276 24380 5277 24444
rect 5211 24379 5277 24380
rect 5214 22405 5274 24379
rect 5211 22404 5277 22405
rect 5211 22340 5212 22404
rect 5276 22340 5277 22404
rect 5211 22339 5277 22340
rect 5398 21181 5458 34035
rect 5763 32740 5829 32741
rect 5763 32676 5764 32740
rect 5828 32676 5829 32740
rect 5763 32675 5829 32676
rect 5579 32468 5645 32469
rect 5579 32404 5580 32468
rect 5644 32404 5645 32468
rect 5579 32403 5645 32404
rect 5582 30973 5642 32403
rect 5766 31653 5826 32675
rect 5763 31652 5829 31653
rect 5763 31588 5764 31652
rect 5828 31588 5829 31652
rect 5763 31587 5829 31588
rect 5579 30972 5645 30973
rect 5579 30908 5580 30972
rect 5644 30908 5645 30972
rect 5579 30907 5645 30908
rect 5579 30836 5645 30837
rect 5579 30772 5580 30836
rect 5644 30772 5645 30836
rect 5579 30771 5645 30772
rect 5582 26757 5642 30771
rect 5766 30565 5826 31587
rect 5763 30564 5829 30565
rect 5763 30500 5764 30564
rect 5828 30500 5829 30564
rect 5763 30499 5829 30500
rect 5950 30293 6010 40019
rect 6131 36820 6197 36821
rect 6131 36756 6132 36820
rect 6196 36756 6197 36820
rect 6131 36755 6197 36756
rect 6134 32605 6194 36755
rect 6131 32604 6197 32605
rect 6131 32540 6132 32604
rect 6196 32540 6197 32604
rect 6131 32539 6197 32540
rect 5947 30292 6013 30293
rect 5947 30228 5948 30292
rect 6012 30228 6013 30292
rect 5947 30227 6013 30228
rect 5763 30156 5829 30157
rect 5763 30092 5764 30156
rect 5828 30092 5829 30156
rect 5763 30091 5829 30092
rect 5766 27165 5826 30091
rect 5950 29613 6010 30227
rect 5947 29612 6013 29613
rect 5947 29548 5948 29612
rect 6012 29548 6013 29612
rect 5947 29547 6013 29548
rect 6134 28797 6194 32539
rect 6502 30837 6562 40019
rect 6870 38670 6930 41370
rect 7603 39404 7669 39405
rect 7603 39340 7604 39404
rect 7668 39340 7669 39404
rect 7603 39339 7669 39340
rect 6870 38610 7298 38670
rect 7051 35596 7117 35597
rect 7051 35532 7052 35596
rect 7116 35532 7117 35596
rect 7051 35531 7117 35532
rect 6867 33148 6933 33149
rect 6867 33084 6868 33148
rect 6932 33084 6933 33148
rect 6867 33083 6933 33084
rect 6870 32061 6930 33083
rect 6867 32060 6933 32061
rect 6867 31996 6868 32060
rect 6932 31996 6933 32060
rect 6867 31995 6933 31996
rect 7054 31770 7114 35531
rect 6870 31710 7114 31770
rect 6499 30836 6565 30837
rect 6499 30772 6500 30836
rect 6564 30772 6565 30836
rect 6499 30771 6565 30772
rect 6499 30564 6565 30565
rect 6499 30500 6500 30564
rect 6564 30500 6565 30564
rect 6499 30499 6565 30500
rect 6315 29476 6381 29477
rect 6315 29412 6316 29476
rect 6380 29412 6381 29476
rect 6315 29411 6381 29412
rect 6131 28796 6197 28797
rect 6131 28732 6132 28796
rect 6196 28732 6197 28796
rect 6131 28731 6197 28732
rect 6318 28661 6378 29411
rect 6315 28660 6381 28661
rect 6315 28596 6316 28660
rect 6380 28596 6381 28660
rect 6315 28595 6381 28596
rect 6131 28116 6197 28117
rect 6131 28052 6132 28116
rect 6196 28052 6197 28116
rect 6131 28051 6197 28052
rect 5947 27300 6013 27301
rect 5947 27236 5948 27300
rect 6012 27236 6013 27300
rect 5947 27235 6013 27236
rect 5763 27164 5829 27165
rect 5763 27100 5764 27164
rect 5828 27100 5829 27164
rect 5763 27099 5829 27100
rect 5579 26756 5645 26757
rect 5579 26692 5580 26756
rect 5644 26692 5645 26756
rect 5579 26691 5645 26692
rect 5579 26620 5645 26621
rect 5579 26556 5580 26620
rect 5644 26556 5645 26620
rect 5579 26555 5645 26556
rect 5582 24850 5642 26555
rect 5763 26212 5829 26213
rect 5763 26148 5764 26212
rect 5828 26148 5829 26212
rect 5763 26147 5829 26148
rect 5766 25669 5826 26147
rect 5763 25668 5829 25669
rect 5763 25604 5764 25668
rect 5828 25604 5829 25668
rect 5763 25603 5829 25604
rect 5582 24790 5780 24850
rect 5579 24716 5645 24717
rect 5579 24652 5580 24716
rect 5644 24652 5645 24716
rect 5720 24714 5780 24790
rect 5720 24654 5826 24714
rect 5579 24651 5645 24652
rect 5582 21589 5642 24651
rect 5766 24445 5826 24654
rect 5763 24444 5829 24445
rect 5763 24380 5764 24444
rect 5828 24380 5829 24444
rect 5763 24379 5829 24380
rect 5950 22677 6010 27235
rect 6134 24581 6194 28051
rect 6318 27029 6378 28595
rect 6502 28389 6562 30499
rect 6683 30428 6749 30429
rect 6683 30364 6684 30428
rect 6748 30364 6749 30428
rect 6683 30363 6749 30364
rect 6499 28388 6565 28389
rect 6499 28324 6500 28388
rect 6564 28324 6565 28388
rect 6499 28323 6565 28324
rect 6315 27028 6381 27029
rect 6315 26964 6316 27028
rect 6380 26964 6381 27028
rect 6315 26963 6381 26964
rect 6315 26348 6381 26349
rect 6315 26284 6316 26348
rect 6380 26284 6381 26348
rect 6315 26283 6381 26284
rect 6318 25805 6378 26283
rect 6502 25941 6562 28323
rect 6499 25940 6565 25941
rect 6499 25876 6500 25940
rect 6564 25876 6565 25940
rect 6499 25875 6565 25876
rect 6315 25804 6381 25805
rect 6315 25740 6316 25804
rect 6380 25740 6381 25804
rect 6315 25739 6381 25740
rect 6131 24580 6197 24581
rect 6131 24516 6132 24580
rect 6196 24516 6197 24580
rect 6131 24515 6197 24516
rect 6131 24444 6197 24445
rect 6131 24380 6132 24444
rect 6196 24380 6197 24444
rect 6131 24379 6197 24380
rect 5947 22676 6013 22677
rect 5947 22612 5948 22676
rect 6012 22612 6013 22676
rect 5947 22611 6013 22612
rect 6134 22538 6194 24379
rect 5766 22478 6194 22538
rect 5579 21588 5645 21589
rect 5579 21524 5580 21588
rect 5644 21524 5645 21588
rect 5579 21523 5645 21524
rect 5395 21180 5461 21181
rect 5395 21116 5396 21180
rect 5460 21116 5461 21180
rect 5395 21115 5461 21116
rect 5579 21180 5645 21181
rect 5579 21116 5580 21180
rect 5644 21116 5645 21180
rect 5579 21115 5645 21116
rect 5027 20772 5093 20773
rect 5027 20708 5028 20772
rect 5092 20708 5093 20772
rect 5027 20707 5093 20708
rect 5030 18733 5090 20707
rect 5211 20500 5277 20501
rect 5211 20436 5212 20500
rect 5276 20436 5277 20500
rect 5211 20435 5277 20436
rect 5027 18732 5093 18733
rect 5027 18668 5028 18732
rect 5092 18668 5093 18732
rect 5027 18667 5093 18668
rect 4843 18324 4909 18325
rect 4843 18260 4844 18324
rect 4908 18260 4909 18324
rect 4843 18259 4909 18260
rect 5030 18053 5090 18667
rect 5214 18325 5274 20435
rect 5395 20228 5461 20229
rect 5395 20164 5396 20228
rect 5460 20164 5461 20228
rect 5395 20163 5461 20164
rect 5211 18324 5277 18325
rect 5211 18260 5212 18324
rect 5276 18260 5277 18324
rect 5211 18259 5277 18260
rect 5398 18189 5458 20163
rect 5395 18188 5461 18189
rect 5395 18124 5396 18188
rect 5460 18124 5461 18188
rect 5395 18123 5461 18124
rect 5027 18052 5093 18053
rect 5027 17988 5028 18052
rect 5092 17988 5093 18052
rect 5027 17987 5093 17988
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 5027 17780 5093 17781
rect 5027 17716 5028 17780
rect 5092 17716 5093 17780
rect 5027 17715 5093 17716
rect 4843 17236 4909 17237
rect 4843 17172 4844 17236
rect 4908 17172 4909 17236
rect 4843 17171 4909 17172
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4107 15196 4173 15197
rect 4107 15132 4108 15196
rect 4172 15132 4173 15196
rect 4107 15131 4173 15132
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3003 13700 3069 13701
rect 3003 13636 3004 13700
rect 3068 13636 3069 13700
rect 3003 13635 3069 13636
rect 2819 13428 2885 13429
rect 2819 13364 2820 13428
rect 2884 13364 2885 13428
rect 2819 13363 2885 13364
rect 2451 12340 2517 12341
rect 2451 12276 2452 12340
rect 2516 12276 2517 12340
rect 2451 12275 2517 12276
rect 2822 11797 2882 13363
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4846 13837 4906 17171
rect 4843 13836 4909 13837
rect 4843 13772 4844 13836
rect 4908 13772 4909 13836
rect 4843 13771 4909 13772
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 5030 13429 5090 17715
rect 5582 15333 5642 21115
rect 5766 18325 5826 22478
rect 6318 21997 6378 25739
rect 6499 25124 6565 25125
rect 6499 25060 6500 25124
rect 6564 25060 6565 25124
rect 6499 25059 6565 25060
rect 6502 22677 6562 25059
rect 6499 22676 6565 22677
rect 6499 22612 6500 22676
rect 6564 22612 6565 22676
rect 6499 22611 6565 22612
rect 6499 22268 6565 22269
rect 6499 22204 6500 22268
rect 6564 22204 6565 22268
rect 6499 22203 6565 22204
rect 5947 21996 6013 21997
rect 5947 21932 5948 21996
rect 6012 21932 6013 21996
rect 5947 21931 6013 21932
rect 6315 21996 6381 21997
rect 6315 21932 6316 21996
rect 6380 21932 6381 21996
rect 6315 21931 6381 21932
rect 5763 18324 5829 18325
rect 5763 18260 5764 18324
rect 5828 18260 5829 18324
rect 5763 18259 5829 18260
rect 5579 15332 5645 15333
rect 5579 15268 5580 15332
rect 5644 15268 5645 15332
rect 5579 15267 5645 15268
rect 5950 15061 6010 21931
rect 6502 20498 6562 22203
rect 6318 20438 6562 20498
rect 6318 19821 6378 20438
rect 6686 20365 6746 30363
rect 6870 24717 6930 31710
rect 7238 30293 7298 38610
rect 7606 33557 7666 39339
rect 7790 34917 7850 43555
rect 10056 42464 10376 43024
rect 10056 42400 10064 42464
rect 10128 42400 10144 42464
rect 10208 42400 10224 42464
rect 10288 42400 10304 42464
rect 10368 42400 10376 42464
rect 7971 41444 8037 41445
rect 7971 41380 7972 41444
rect 8036 41380 8037 41444
rect 7971 41379 8037 41380
rect 7787 34916 7853 34917
rect 7787 34852 7788 34916
rect 7852 34852 7853 34916
rect 7787 34851 7853 34852
rect 7974 34101 8034 41379
rect 10056 41376 10376 42400
rect 10056 41312 10064 41376
rect 10128 41312 10144 41376
rect 10208 41312 10224 41376
rect 10288 41312 10304 41376
rect 10368 41312 10376 41376
rect 10056 40288 10376 41312
rect 10056 40224 10064 40288
rect 10128 40224 10144 40288
rect 10208 40224 10224 40288
rect 10288 40224 10304 40288
rect 10368 40224 10376 40288
rect 9443 39676 9509 39677
rect 9443 39612 9444 39676
rect 9508 39612 9509 39676
rect 9443 39611 9509 39612
rect 8339 39540 8405 39541
rect 8339 39476 8340 39540
rect 8404 39476 8405 39540
rect 8339 39475 8405 39476
rect 8155 38180 8221 38181
rect 8155 38116 8156 38180
rect 8220 38116 8221 38180
rect 8155 38115 8221 38116
rect 8158 35733 8218 38115
rect 8342 36821 8402 39475
rect 9075 38452 9141 38453
rect 9075 38388 9076 38452
rect 9140 38388 9141 38452
rect 9075 38387 9141 38388
rect 8523 38316 8589 38317
rect 8523 38252 8524 38316
rect 8588 38252 8589 38316
rect 8523 38251 8589 38252
rect 8707 38316 8773 38317
rect 8707 38252 8708 38316
rect 8772 38252 8773 38316
rect 8707 38251 8773 38252
rect 8526 37501 8586 38251
rect 8523 37500 8589 37501
rect 8523 37436 8524 37500
rect 8588 37436 8589 37500
rect 8523 37435 8589 37436
rect 8523 37092 8589 37093
rect 8523 37028 8524 37092
rect 8588 37028 8589 37092
rect 8523 37027 8589 37028
rect 8339 36820 8405 36821
rect 8339 36756 8340 36820
rect 8404 36756 8405 36820
rect 8339 36755 8405 36756
rect 8155 35732 8221 35733
rect 8155 35668 8156 35732
rect 8220 35668 8221 35732
rect 8155 35667 8221 35668
rect 8155 34508 8221 34509
rect 8155 34444 8156 34508
rect 8220 34444 8221 34508
rect 8155 34443 8221 34444
rect 7971 34100 8037 34101
rect 7971 34036 7972 34100
rect 8036 34036 8037 34100
rect 7971 34035 8037 34036
rect 7603 33556 7669 33557
rect 7603 33492 7604 33556
rect 7668 33492 7669 33556
rect 7603 33491 7669 33492
rect 8158 33421 8218 34443
rect 8155 33420 8221 33421
rect 8155 33356 8156 33420
rect 8220 33356 8221 33420
rect 8155 33355 8221 33356
rect 7419 33148 7485 33149
rect 7419 33084 7420 33148
rect 7484 33084 7485 33148
rect 7419 33083 7485 33084
rect 7422 31789 7482 33083
rect 7971 32604 8037 32605
rect 7971 32540 7972 32604
rect 8036 32540 8037 32604
rect 7971 32539 8037 32540
rect 7974 32061 8034 32539
rect 7787 32060 7853 32061
rect 7787 31996 7788 32060
rect 7852 31996 7853 32060
rect 7787 31995 7853 31996
rect 7971 32060 8037 32061
rect 7971 31996 7972 32060
rect 8036 31996 8037 32060
rect 7971 31995 8037 31996
rect 7419 31788 7485 31789
rect 7419 31724 7420 31788
rect 7484 31724 7485 31788
rect 7419 31723 7485 31724
rect 7790 31517 7850 31995
rect 8158 31770 8218 33355
rect 8526 31770 8586 37027
rect 8710 34373 8770 38251
rect 8891 38044 8957 38045
rect 8891 37980 8892 38044
rect 8956 37980 8957 38044
rect 8891 37979 8957 37980
rect 8894 37501 8954 37979
rect 8891 37500 8957 37501
rect 8891 37436 8892 37500
rect 8956 37436 8957 37500
rect 8891 37435 8957 37436
rect 9078 36413 9138 38387
rect 9259 38180 9325 38181
rect 9259 38116 9260 38180
rect 9324 38116 9325 38180
rect 9259 38115 9325 38116
rect 9262 37229 9322 38115
rect 9446 37501 9506 39611
rect 10056 39200 10376 40224
rect 10056 39136 10064 39200
rect 10128 39136 10144 39200
rect 10208 39136 10224 39200
rect 10288 39136 10304 39200
rect 10368 39136 10376 39200
rect 10056 38112 10376 39136
rect 10056 38048 10064 38112
rect 10128 38048 10144 38112
rect 10208 38048 10224 38112
rect 10288 38048 10304 38112
rect 10368 38048 10376 38112
rect 9443 37500 9509 37501
rect 9443 37436 9444 37500
rect 9508 37436 9509 37500
rect 9443 37435 9509 37436
rect 9259 37228 9325 37229
rect 9259 37164 9260 37228
rect 9324 37164 9325 37228
rect 9259 37163 9325 37164
rect 10056 37024 10376 38048
rect 10056 36960 10064 37024
rect 10128 36960 10144 37024
rect 10208 36960 10224 37024
rect 10288 36960 10304 37024
rect 10368 36960 10376 37024
rect 9075 36412 9141 36413
rect 9075 36348 9076 36412
rect 9140 36348 9141 36412
rect 9075 36347 9141 36348
rect 9075 36004 9141 36005
rect 9075 35940 9076 36004
rect 9140 35940 9141 36004
rect 9075 35939 9141 35940
rect 8707 34372 8773 34373
rect 8707 34308 8708 34372
rect 8772 34308 8773 34372
rect 8707 34307 8773 34308
rect 9078 32741 9138 35939
rect 10056 35936 10376 36960
rect 10056 35872 10064 35936
rect 10128 35872 10144 35936
rect 10208 35872 10224 35936
rect 10288 35872 10304 35936
rect 10368 35872 10376 35936
rect 9259 35188 9325 35189
rect 9259 35124 9260 35188
rect 9324 35124 9325 35188
rect 9259 35123 9325 35124
rect 9075 32740 9141 32741
rect 9075 32676 9076 32740
rect 9140 32676 9141 32740
rect 9075 32675 9141 32676
rect 9075 32604 9141 32605
rect 9075 32540 9076 32604
rect 9140 32540 9141 32604
rect 9075 32539 9141 32540
rect 9078 32061 9138 32539
rect 9075 32060 9141 32061
rect 9075 31996 9076 32060
rect 9140 31996 9141 32060
rect 9075 31995 9141 31996
rect 7974 31710 8218 31770
rect 8342 31710 8586 31770
rect 7787 31516 7853 31517
rect 7787 31452 7788 31516
rect 7852 31452 7853 31516
rect 7787 31451 7853 31452
rect 7419 30836 7485 30837
rect 7419 30772 7420 30836
rect 7484 30772 7485 30836
rect 7419 30771 7485 30772
rect 7235 30292 7301 30293
rect 7235 30228 7236 30292
rect 7300 30228 7301 30292
rect 7235 30227 7301 30228
rect 7051 30020 7117 30021
rect 7051 29956 7052 30020
rect 7116 29956 7117 30020
rect 7051 29955 7117 29956
rect 7054 26485 7114 29955
rect 7422 29610 7482 30771
rect 7238 29550 7482 29610
rect 7051 26484 7117 26485
rect 7051 26420 7052 26484
rect 7116 26420 7117 26484
rect 7051 26419 7117 26420
rect 6867 24716 6933 24717
rect 6867 24652 6868 24716
rect 6932 24652 6933 24716
rect 6867 24651 6933 24652
rect 7054 24445 7114 26419
rect 7051 24444 7117 24445
rect 7051 24380 7052 24444
rect 7116 24380 7117 24444
rect 7051 24379 7117 24380
rect 7238 24170 7298 29550
rect 7787 29068 7853 29069
rect 7787 29004 7788 29068
rect 7852 29004 7853 29068
rect 7787 29003 7853 29004
rect 7419 28524 7485 28525
rect 7419 28460 7420 28524
rect 7484 28460 7485 28524
rect 7419 28459 7485 28460
rect 6870 24110 7298 24170
rect 6870 23765 6930 24110
rect 7235 24036 7301 24037
rect 7235 23972 7236 24036
rect 7300 23972 7301 24036
rect 7235 23971 7301 23972
rect 6867 23764 6933 23765
rect 6867 23700 6868 23764
rect 6932 23700 6933 23764
rect 6867 23699 6933 23700
rect 7051 23764 7117 23765
rect 7051 23700 7052 23764
rect 7116 23700 7117 23764
rect 7051 23699 7117 23700
rect 6867 23220 6933 23221
rect 6867 23156 6868 23220
rect 6932 23218 6933 23220
rect 7054 23218 7114 23699
rect 7238 23221 7298 23971
rect 7422 23629 7482 28459
rect 7603 27708 7669 27709
rect 7603 27644 7604 27708
rect 7668 27644 7669 27708
rect 7603 27643 7669 27644
rect 7419 23628 7485 23629
rect 7419 23564 7420 23628
rect 7484 23564 7485 23628
rect 7419 23563 7485 23564
rect 6932 23158 7114 23218
rect 7235 23220 7301 23221
rect 6932 23156 6933 23158
rect 6867 23155 6933 23156
rect 7235 23156 7236 23220
rect 7300 23156 7301 23220
rect 7235 23155 7301 23156
rect 7419 22948 7485 22949
rect 7419 22946 7420 22948
rect 7054 22886 7420 22946
rect 6867 21996 6933 21997
rect 6867 21932 6868 21996
rect 6932 21932 6933 21996
rect 6867 21931 6933 21932
rect 6683 20364 6749 20365
rect 6683 20362 6684 20364
rect 6502 20302 6684 20362
rect 6315 19820 6381 19821
rect 6315 19756 6316 19820
rect 6380 19756 6381 19820
rect 6315 19755 6381 19756
rect 6502 19350 6562 20302
rect 6683 20300 6684 20302
rect 6748 20300 6749 20364
rect 6683 20299 6749 20300
rect 6686 20208 6746 20299
rect 6870 20229 6930 21931
rect 6867 20228 6933 20229
rect 6867 20164 6868 20228
rect 6932 20164 6933 20228
rect 6867 20163 6933 20164
rect 6683 20092 6749 20093
rect 6683 20028 6684 20092
rect 6748 20028 6749 20092
rect 6683 20027 6749 20028
rect 6134 19290 6562 19350
rect 6134 17237 6194 19290
rect 6315 19140 6381 19141
rect 6315 19076 6316 19140
rect 6380 19076 6381 19140
rect 6315 19075 6381 19076
rect 6318 17645 6378 19075
rect 6315 17644 6381 17645
rect 6315 17580 6316 17644
rect 6380 17580 6381 17644
rect 6315 17579 6381 17580
rect 6686 17237 6746 20027
rect 7054 19682 7114 22886
rect 7419 22884 7420 22886
rect 7484 22884 7485 22948
rect 7419 22883 7485 22884
rect 7235 22540 7301 22541
rect 7235 22476 7236 22540
rect 7300 22476 7301 22540
rect 7235 22475 7301 22476
rect 6870 19622 7114 19682
rect 6870 18189 6930 19622
rect 7051 19412 7117 19413
rect 7051 19348 7052 19412
rect 7116 19348 7117 19412
rect 7051 19347 7117 19348
rect 6867 18188 6933 18189
rect 6867 18124 6868 18188
rect 6932 18124 6933 18188
rect 6867 18123 6933 18124
rect 6131 17236 6197 17237
rect 6131 17172 6132 17236
rect 6196 17172 6197 17236
rect 6131 17171 6197 17172
rect 6683 17236 6749 17237
rect 6683 17172 6684 17236
rect 6748 17172 6749 17236
rect 6683 17171 6749 17172
rect 6867 16964 6933 16965
rect 6867 16900 6868 16964
rect 6932 16900 6933 16964
rect 6867 16899 6933 16900
rect 5947 15060 6013 15061
rect 5947 14996 5948 15060
rect 6012 14996 6013 15060
rect 5947 14995 6013 14996
rect 5027 13428 5093 13429
rect 5027 13364 5028 13428
rect 5092 13364 5093 13428
rect 5027 13363 5093 13364
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4107 12204 4173 12205
rect 4107 12140 4108 12204
rect 4172 12140 4173 12204
rect 4107 12139 4173 12140
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 2819 11796 2885 11797
rect 2819 11732 2820 11796
rect 2884 11732 2885 11796
rect 2819 11731 2885 11732
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 4110 10165 4170 12139
rect 4316 11456 4636 12480
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4107 10164 4173 10165
rect 4107 10100 4108 10164
rect 4172 10100 4173 10164
rect 4107 10099 4173 10100
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 2083 9076 2149 9077
rect 2083 9012 2084 9076
rect 2148 9012 2149 9076
rect 2083 9011 2149 9012
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 611 4724 677 4725
rect 611 4660 612 4724
rect 676 4660 677 4724
rect 611 4659 677 4660
rect 59 4452 125 4453
rect 59 4388 60 4452
rect 124 4388 125 4452
rect 59 4387 125 4388
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 6870 4045 6930 16899
rect 7054 6765 7114 19347
rect 7238 16557 7298 22475
rect 7606 20909 7666 27643
rect 7790 22949 7850 29003
rect 7974 25941 8034 31710
rect 8342 30970 8402 31710
rect 9075 31652 9141 31653
rect 9075 31588 9076 31652
rect 9140 31588 9141 31652
rect 9075 31587 9141 31588
rect 8158 30910 8402 30970
rect 8158 26349 8218 30910
rect 8707 29068 8773 29069
rect 8707 29004 8708 29068
rect 8772 29004 8773 29068
rect 8707 29003 8773 29004
rect 8523 27980 8589 27981
rect 8523 27916 8524 27980
rect 8588 27916 8589 27980
rect 8523 27915 8589 27916
rect 8155 26348 8221 26349
rect 8155 26284 8156 26348
rect 8220 26284 8221 26348
rect 8155 26283 8221 26284
rect 8155 26212 8221 26213
rect 8155 26148 8156 26212
rect 8220 26148 8221 26212
rect 8155 26147 8221 26148
rect 7971 25940 8037 25941
rect 7971 25876 7972 25940
rect 8036 25876 8037 25940
rect 7971 25875 8037 25876
rect 7971 24988 8037 24989
rect 7971 24924 7972 24988
rect 8036 24924 8037 24988
rect 7971 24923 8037 24924
rect 7787 22948 7853 22949
rect 7787 22884 7788 22948
rect 7852 22884 7853 22948
rect 7787 22883 7853 22884
rect 7787 22132 7853 22133
rect 7787 22068 7788 22132
rect 7852 22068 7853 22132
rect 7787 22067 7853 22068
rect 7603 20908 7669 20909
rect 7603 20844 7604 20908
rect 7668 20844 7669 20908
rect 7603 20843 7669 20844
rect 7790 19350 7850 22067
rect 7606 19290 7850 19350
rect 7419 18596 7485 18597
rect 7419 18532 7420 18596
rect 7484 18532 7485 18596
rect 7419 18531 7485 18532
rect 7235 16556 7301 16557
rect 7235 16492 7236 16556
rect 7300 16492 7301 16556
rect 7235 16491 7301 16492
rect 7238 12885 7298 16491
rect 7422 13701 7482 18531
rect 7606 16829 7666 19290
rect 7974 18189 8034 24923
rect 8158 22949 8218 26147
rect 8339 26076 8405 26077
rect 8339 26012 8340 26076
rect 8404 26012 8405 26076
rect 8339 26011 8405 26012
rect 8155 22948 8221 22949
rect 8155 22884 8156 22948
rect 8220 22884 8221 22948
rect 8155 22883 8221 22884
rect 8155 22404 8221 22405
rect 8155 22340 8156 22404
rect 8220 22340 8221 22404
rect 8155 22339 8221 22340
rect 7971 18188 8037 18189
rect 7971 18124 7972 18188
rect 8036 18124 8037 18188
rect 7971 18123 8037 18124
rect 7603 16828 7669 16829
rect 7603 16764 7604 16828
rect 7668 16764 7669 16828
rect 7603 16763 7669 16764
rect 7419 13700 7485 13701
rect 7419 13636 7420 13700
rect 7484 13636 7485 13700
rect 7419 13635 7485 13636
rect 8158 13021 8218 22339
rect 8342 21997 8402 26011
rect 8526 25261 8586 27915
rect 8523 25260 8589 25261
rect 8523 25196 8524 25260
rect 8588 25196 8589 25260
rect 8523 25195 8589 25196
rect 8523 25124 8589 25125
rect 8523 25060 8524 25124
rect 8588 25060 8589 25124
rect 8523 25059 8589 25060
rect 8526 23221 8586 25059
rect 8710 24717 8770 29003
rect 8891 26348 8957 26349
rect 8891 26284 8892 26348
rect 8956 26284 8957 26348
rect 8891 26283 8957 26284
rect 8894 25125 8954 26283
rect 8891 25124 8957 25125
rect 8891 25060 8892 25124
rect 8956 25060 8957 25124
rect 8891 25059 8957 25060
rect 8891 24988 8957 24989
rect 8891 24924 8892 24988
rect 8956 24924 8957 24988
rect 8891 24923 8957 24924
rect 8707 24716 8773 24717
rect 8707 24652 8708 24716
rect 8772 24652 8773 24716
rect 8707 24651 8773 24652
rect 8710 23629 8770 24651
rect 8707 23628 8773 23629
rect 8707 23564 8708 23628
rect 8772 23564 8773 23628
rect 8707 23563 8773 23564
rect 8894 23490 8954 24923
rect 8710 23430 8954 23490
rect 8523 23220 8589 23221
rect 8523 23156 8524 23220
rect 8588 23156 8589 23220
rect 8523 23155 8589 23156
rect 8523 22948 8589 22949
rect 8523 22884 8524 22948
rect 8588 22884 8589 22948
rect 8523 22883 8589 22884
rect 8339 21996 8405 21997
rect 8339 21932 8340 21996
rect 8404 21932 8405 21996
rect 8339 21931 8405 21932
rect 8339 21588 8405 21589
rect 8339 21524 8340 21588
rect 8404 21524 8405 21588
rect 8339 21523 8405 21524
rect 8342 18597 8402 21523
rect 8526 20501 8586 22883
rect 8710 22677 8770 23430
rect 8891 23356 8957 23357
rect 8891 23292 8892 23356
rect 8956 23292 8957 23356
rect 8891 23291 8957 23292
rect 8707 22676 8773 22677
rect 8707 22612 8708 22676
rect 8772 22612 8773 22676
rect 8707 22611 8773 22612
rect 8707 20908 8773 20909
rect 8707 20844 8708 20908
rect 8772 20844 8773 20908
rect 8707 20843 8773 20844
rect 8523 20500 8589 20501
rect 8523 20436 8524 20500
rect 8588 20436 8589 20500
rect 8523 20435 8589 20436
rect 8339 18596 8405 18597
rect 8339 18532 8340 18596
rect 8404 18532 8405 18596
rect 8339 18531 8405 18532
rect 8523 17644 8589 17645
rect 8523 17580 8524 17644
rect 8588 17580 8589 17644
rect 8523 17579 8589 17580
rect 8339 17236 8405 17237
rect 8339 17172 8340 17236
rect 8404 17172 8405 17236
rect 8339 17171 8405 17172
rect 8342 15469 8402 17171
rect 8339 15468 8405 15469
rect 8339 15404 8340 15468
rect 8404 15404 8405 15468
rect 8339 15403 8405 15404
rect 8155 13020 8221 13021
rect 8155 12956 8156 13020
rect 8220 12956 8221 13020
rect 8155 12955 8221 12956
rect 7235 12884 7301 12885
rect 7235 12820 7236 12884
rect 7300 12820 7301 12884
rect 7235 12819 7301 12820
rect 8526 12205 8586 17579
rect 8710 16421 8770 20843
rect 8894 19549 8954 23291
rect 8891 19548 8957 19549
rect 8891 19484 8892 19548
rect 8956 19484 8957 19548
rect 8891 19483 8957 19484
rect 9078 17237 9138 31587
rect 9262 30293 9322 35123
rect 10056 34848 10376 35872
rect 10056 34784 10064 34848
rect 10128 34784 10144 34848
rect 10208 34784 10224 34848
rect 10288 34784 10304 34848
rect 10368 34784 10376 34848
rect 10056 33760 10376 34784
rect 10716 43008 11036 43024
rect 10716 42944 10724 43008
rect 10788 42944 10804 43008
rect 10868 42944 10884 43008
rect 10948 42944 10964 43008
rect 11028 42944 11036 43008
rect 10716 41920 11036 42944
rect 10716 41856 10724 41920
rect 10788 41856 10804 41920
rect 10868 41856 10884 41920
rect 10948 41856 10964 41920
rect 11028 41856 11036 41920
rect 10716 40832 11036 41856
rect 10716 40768 10724 40832
rect 10788 40768 10804 40832
rect 10868 40768 10884 40832
rect 10948 40768 10964 40832
rect 11028 40768 11036 40832
rect 10716 39744 11036 40768
rect 10716 39680 10724 39744
rect 10788 39680 10804 39744
rect 10868 39680 10884 39744
rect 10948 39680 10964 39744
rect 11028 39680 11036 39744
rect 10716 38656 11036 39680
rect 10716 38592 10724 38656
rect 10788 38592 10804 38656
rect 10868 38592 10884 38656
rect 10948 38592 10964 38656
rect 11028 38592 11036 38656
rect 10716 37568 11036 38592
rect 10716 37504 10724 37568
rect 10788 37504 10804 37568
rect 10868 37504 10884 37568
rect 10948 37504 10964 37568
rect 11028 37504 11036 37568
rect 10716 36480 11036 37504
rect 10716 36416 10724 36480
rect 10788 36416 10804 36480
rect 10868 36416 10884 36480
rect 10948 36416 10964 36480
rect 11028 36416 11036 36480
rect 10716 35392 11036 36416
rect 10716 35328 10724 35392
rect 10788 35328 10804 35392
rect 10868 35328 10884 35392
rect 10948 35328 10964 35392
rect 11028 35328 11036 35392
rect 10716 34304 11036 35328
rect 10716 34240 10724 34304
rect 10788 34240 10804 34304
rect 10868 34240 10884 34304
rect 10948 34240 10964 34304
rect 11028 34240 11036 34304
rect 10547 33964 10613 33965
rect 10547 33900 10548 33964
rect 10612 33900 10613 33964
rect 10547 33899 10613 33900
rect 10056 33696 10064 33760
rect 10128 33696 10144 33760
rect 10208 33696 10224 33760
rect 10288 33696 10304 33760
rect 10368 33696 10376 33760
rect 9443 33692 9509 33693
rect 9443 33628 9444 33692
rect 9508 33628 9509 33692
rect 9443 33627 9509 33628
rect 9259 30292 9325 30293
rect 9259 30228 9260 30292
rect 9324 30228 9325 30292
rect 9259 30227 9325 30228
rect 9446 29205 9506 33627
rect 10056 32672 10376 33696
rect 10056 32608 10064 32672
rect 10128 32608 10144 32672
rect 10208 32608 10224 32672
rect 10288 32608 10304 32672
rect 10368 32608 10376 32672
rect 10056 31584 10376 32608
rect 10056 31520 10064 31584
rect 10128 31520 10144 31584
rect 10208 31520 10224 31584
rect 10288 31520 10304 31584
rect 10368 31520 10376 31584
rect 9627 30700 9693 30701
rect 9627 30636 9628 30700
rect 9692 30636 9693 30700
rect 9627 30635 9693 30636
rect 9443 29204 9509 29205
rect 9443 29140 9444 29204
rect 9508 29140 9509 29204
rect 9443 29139 9509 29140
rect 9443 27300 9509 27301
rect 9443 27236 9444 27300
rect 9508 27236 9509 27300
rect 9443 27235 9509 27236
rect 9259 26892 9325 26893
rect 9259 26828 9260 26892
rect 9324 26828 9325 26892
rect 9259 26827 9325 26828
rect 9262 25397 9322 26827
rect 9259 25396 9325 25397
rect 9259 25332 9260 25396
rect 9324 25332 9325 25396
rect 9259 25331 9325 25332
rect 9259 23900 9325 23901
rect 9259 23836 9260 23900
rect 9324 23836 9325 23900
rect 9259 23835 9325 23836
rect 9262 22813 9322 23835
rect 9446 23765 9506 27235
rect 9443 23764 9509 23765
rect 9443 23700 9444 23764
rect 9508 23700 9509 23764
rect 9443 23699 9509 23700
rect 9443 23492 9509 23493
rect 9443 23428 9444 23492
rect 9508 23428 9509 23492
rect 9443 23427 9509 23428
rect 9446 22949 9506 23427
rect 9443 22948 9509 22949
rect 9443 22884 9444 22948
rect 9508 22884 9509 22948
rect 9443 22883 9509 22884
rect 9259 22812 9325 22813
rect 9259 22748 9260 22812
rect 9324 22748 9325 22812
rect 9259 22747 9325 22748
rect 9262 21858 9322 22747
rect 9443 21860 9509 21861
rect 9443 21858 9444 21860
rect 9262 21798 9444 21858
rect 9443 21796 9444 21798
rect 9508 21796 9509 21860
rect 9443 21795 9509 21796
rect 9446 17645 9506 21795
rect 9630 21450 9690 30635
rect 9811 30564 9877 30565
rect 9811 30500 9812 30564
rect 9876 30500 9877 30564
rect 9811 30499 9877 30500
rect 9814 21589 9874 30499
rect 10056 30496 10376 31520
rect 10056 30432 10064 30496
rect 10128 30432 10144 30496
rect 10208 30432 10224 30496
rect 10288 30432 10304 30496
rect 10368 30432 10376 30496
rect 10056 29408 10376 30432
rect 10056 29344 10064 29408
rect 10128 29344 10144 29408
rect 10208 29344 10224 29408
rect 10288 29344 10304 29408
rect 10368 29344 10376 29408
rect 10056 28320 10376 29344
rect 10056 28256 10064 28320
rect 10128 28256 10144 28320
rect 10208 28256 10224 28320
rect 10288 28256 10304 28320
rect 10368 28256 10376 28320
rect 10056 27232 10376 28256
rect 10550 27981 10610 33899
rect 10716 33216 11036 34240
rect 10716 33152 10724 33216
rect 10788 33152 10804 33216
rect 10868 33152 10884 33216
rect 10948 33152 10964 33216
rect 11028 33152 11036 33216
rect 10716 32128 11036 33152
rect 10716 32064 10724 32128
rect 10788 32064 10804 32128
rect 10868 32064 10884 32128
rect 10948 32064 10964 32128
rect 11028 32064 11036 32128
rect 10716 31040 11036 32064
rect 10716 30976 10724 31040
rect 10788 30976 10804 31040
rect 10868 30976 10884 31040
rect 10948 30976 10964 31040
rect 11028 30976 11036 31040
rect 10716 29952 11036 30976
rect 10716 29888 10724 29952
rect 10788 29888 10804 29952
rect 10868 29888 10884 29952
rect 10948 29888 10964 29952
rect 11028 29888 11036 29952
rect 10716 28864 11036 29888
rect 10716 28800 10724 28864
rect 10788 28800 10804 28864
rect 10868 28800 10884 28864
rect 10948 28800 10964 28864
rect 11028 28800 11036 28864
rect 10547 27980 10613 27981
rect 10547 27916 10548 27980
rect 10612 27916 10613 27980
rect 10547 27915 10613 27916
rect 10716 27776 11036 28800
rect 10716 27712 10724 27776
rect 10788 27712 10804 27776
rect 10868 27712 10884 27776
rect 10948 27712 10964 27776
rect 11028 27712 11036 27776
rect 10547 27436 10613 27437
rect 10547 27372 10548 27436
rect 10612 27372 10613 27436
rect 10547 27371 10613 27372
rect 10056 27168 10064 27232
rect 10128 27168 10144 27232
rect 10208 27168 10224 27232
rect 10288 27168 10304 27232
rect 10368 27168 10376 27232
rect 10056 26144 10376 27168
rect 10550 26621 10610 27371
rect 10716 26688 11036 27712
rect 11283 26892 11349 26893
rect 11283 26828 11284 26892
rect 11348 26828 11349 26892
rect 11283 26827 11349 26828
rect 10716 26624 10724 26688
rect 10788 26624 10804 26688
rect 10868 26624 10884 26688
rect 10948 26624 10964 26688
rect 11028 26624 11036 26688
rect 10547 26620 10613 26621
rect 10547 26556 10548 26620
rect 10612 26556 10613 26620
rect 10547 26555 10613 26556
rect 10056 26080 10064 26144
rect 10128 26080 10144 26144
rect 10208 26080 10224 26144
rect 10288 26080 10304 26144
rect 10368 26080 10376 26144
rect 10056 25056 10376 26080
rect 10056 24992 10064 25056
rect 10128 24992 10144 25056
rect 10208 24992 10224 25056
rect 10288 24992 10304 25056
rect 10368 24992 10376 25056
rect 10056 23968 10376 24992
rect 10550 24173 10610 26555
rect 10716 25600 11036 26624
rect 11099 26620 11165 26621
rect 11099 26556 11100 26620
rect 11164 26556 11165 26620
rect 11099 26555 11165 26556
rect 10716 25536 10724 25600
rect 10788 25536 10804 25600
rect 10868 25536 10884 25600
rect 10948 25536 10964 25600
rect 11028 25536 11036 25600
rect 10716 24512 11036 25536
rect 10716 24448 10724 24512
rect 10788 24448 10804 24512
rect 10868 24448 10884 24512
rect 10948 24448 10964 24512
rect 11028 24448 11036 24512
rect 10547 24172 10613 24173
rect 10547 24108 10548 24172
rect 10612 24108 10613 24172
rect 10547 24107 10613 24108
rect 10547 24036 10613 24037
rect 10547 23972 10548 24036
rect 10612 23972 10613 24036
rect 10547 23971 10613 23972
rect 10056 23904 10064 23968
rect 10128 23904 10144 23968
rect 10208 23904 10224 23968
rect 10288 23904 10304 23968
rect 10368 23904 10376 23968
rect 10056 22880 10376 23904
rect 10056 22816 10064 22880
rect 10128 22816 10144 22880
rect 10208 22816 10224 22880
rect 10288 22816 10304 22880
rect 10368 22816 10376 22880
rect 10056 21792 10376 22816
rect 10550 21861 10610 23971
rect 10716 23424 11036 24448
rect 11102 24309 11162 26555
rect 11099 24308 11165 24309
rect 11099 24244 11100 24308
rect 11164 24244 11165 24308
rect 11099 24243 11165 24244
rect 11099 24172 11165 24173
rect 11099 24108 11100 24172
rect 11164 24108 11165 24172
rect 11099 24107 11165 24108
rect 10716 23360 10724 23424
rect 10788 23360 10804 23424
rect 10868 23360 10884 23424
rect 10948 23360 10964 23424
rect 11028 23360 11036 23424
rect 10716 22336 11036 23360
rect 11102 23221 11162 24107
rect 11099 23220 11165 23221
rect 11099 23156 11100 23220
rect 11164 23156 11165 23220
rect 11099 23155 11165 23156
rect 10716 22272 10724 22336
rect 10788 22272 10804 22336
rect 10868 22272 10884 22336
rect 10948 22272 10964 22336
rect 11028 22272 11036 22336
rect 10547 21860 10613 21861
rect 10547 21796 10548 21860
rect 10612 21796 10613 21860
rect 10547 21795 10613 21796
rect 10056 21728 10064 21792
rect 10128 21728 10144 21792
rect 10208 21728 10224 21792
rect 10288 21728 10304 21792
rect 10368 21728 10376 21792
rect 9811 21588 9877 21589
rect 9811 21524 9812 21588
rect 9876 21524 9877 21588
rect 9811 21523 9877 21524
rect 9630 21390 9874 21450
rect 9627 20772 9693 20773
rect 9627 20708 9628 20772
rect 9692 20708 9693 20772
rect 9627 20707 9693 20708
rect 9443 17644 9509 17645
rect 9443 17580 9444 17644
rect 9508 17580 9509 17644
rect 9443 17579 9509 17580
rect 9075 17236 9141 17237
rect 9075 17172 9076 17236
rect 9140 17172 9141 17236
rect 9075 17171 9141 17172
rect 9259 16828 9325 16829
rect 9259 16764 9260 16828
rect 9324 16764 9325 16828
rect 9259 16763 9325 16764
rect 9075 16692 9141 16693
rect 9075 16628 9076 16692
rect 9140 16628 9141 16692
rect 9075 16627 9141 16628
rect 8891 16556 8957 16557
rect 8891 16492 8892 16556
rect 8956 16492 8957 16556
rect 8891 16491 8957 16492
rect 8707 16420 8773 16421
rect 8707 16356 8708 16420
rect 8772 16356 8773 16420
rect 8707 16355 8773 16356
rect 8523 12204 8589 12205
rect 8523 12140 8524 12204
rect 8588 12140 8589 12204
rect 8523 12139 8589 12140
rect 8526 11661 8586 12139
rect 8523 11660 8589 11661
rect 8523 11596 8524 11660
rect 8588 11596 8589 11660
rect 8523 11595 8589 11596
rect 7051 6764 7117 6765
rect 7051 6700 7052 6764
rect 7116 6700 7117 6764
rect 7051 6699 7117 6700
rect 8894 4045 8954 16491
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 8891 4044 8957 4045
rect 8891 3980 8892 4044
rect 8956 3980 8957 4044
rect 8891 3979 8957 3980
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 9078 3773 9138 16627
rect 9262 15061 9322 16763
rect 9259 15060 9325 15061
rect 9259 14996 9260 15060
rect 9324 14996 9325 15060
rect 9259 14995 9325 14996
rect 9446 13565 9506 17579
rect 9630 15061 9690 20707
rect 9814 18733 9874 21390
rect 10056 20704 10376 21728
rect 10547 21588 10613 21589
rect 10547 21524 10548 21588
rect 10612 21524 10613 21588
rect 10547 21523 10613 21524
rect 10056 20640 10064 20704
rect 10128 20640 10144 20704
rect 10208 20640 10224 20704
rect 10288 20640 10304 20704
rect 10368 20640 10376 20704
rect 10056 19616 10376 20640
rect 10056 19552 10064 19616
rect 10128 19552 10144 19616
rect 10208 19552 10224 19616
rect 10288 19552 10304 19616
rect 10368 19552 10376 19616
rect 9811 18732 9877 18733
rect 9811 18668 9812 18732
rect 9876 18668 9877 18732
rect 9811 18667 9877 18668
rect 10056 18528 10376 19552
rect 10056 18464 10064 18528
rect 10128 18464 10144 18528
rect 10208 18464 10224 18528
rect 10288 18464 10304 18528
rect 10368 18464 10376 18528
rect 10056 17440 10376 18464
rect 10056 17376 10064 17440
rect 10128 17376 10144 17440
rect 10208 17376 10224 17440
rect 10288 17376 10304 17440
rect 10368 17376 10376 17440
rect 10056 16352 10376 17376
rect 10056 16288 10064 16352
rect 10128 16288 10144 16352
rect 10208 16288 10224 16352
rect 10288 16288 10304 16352
rect 10368 16288 10376 16352
rect 10056 15264 10376 16288
rect 10550 15469 10610 21523
rect 10716 21248 11036 22272
rect 10716 21184 10724 21248
rect 10788 21184 10804 21248
rect 10868 21184 10884 21248
rect 10948 21184 10964 21248
rect 11028 21184 11036 21248
rect 10716 20160 11036 21184
rect 10716 20096 10724 20160
rect 10788 20096 10804 20160
rect 10868 20096 10884 20160
rect 10948 20096 10964 20160
rect 11028 20096 11036 20160
rect 10716 19072 11036 20096
rect 10716 19008 10724 19072
rect 10788 19008 10804 19072
rect 10868 19008 10884 19072
rect 10948 19008 10964 19072
rect 11028 19008 11036 19072
rect 10716 17984 11036 19008
rect 11102 18325 11162 23155
rect 11286 19277 11346 26827
rect 11283 19276 11349 19277
rect 11283 19212 11284 19276
rect 11348 19212 11349 19276
rect 11283 19211 11349 19212
rect 11283 18868 11349 18869
rect 11283 18804 11284 18868
rect 11348 18804 11349 18868
rect 11283 18803 11349 18804
rect 11099 18324 11165 18325
rect 11099 18260 11100 18324
rect 11164 18260 11165 18324
rect 11099 18259 11165 18260
rect 10716 17920 10724 17984
rect 10788 17920 10804 17984
rect 10868 17920 10884 17984
rect 10948 17920 10964 17984
rect 11028 17920 11036 17984
rect 10716 16896 11036 17920
rect 10716 16832 10724 16896
rect 10788 16832 10804 16896
rect 10868 16832 10884 16896
rect 10948 16832 10964 16896
rect 11028 16832 11036 16896
rect 10716 15808 11036 16832
rect 10716 15744 10724 15808
rect 10788 15744 10804 15808
rect 10868 15744 10884 15808
rect 10948 15744 10964 15808
rect 11028 15744 11036 15808
rect 10547 15468 10613 15469
rect 10547 15404 10548 15468
rect 10612 15404 10613 15468
rect 10547 15403 10613 15404
rect 10056 15200 10064 15264
rect 10128 15200 10144 15264
rect 10208 15200 10224 15264
rect 10288 15200 10304 15264
rect 10368 15200 10376 15264
rect 9627 15060 9693 15061
rect 9627 14996 9628 15060
rect 9692 14996 9693 15060
rect 9627 14995 9693 14996
rect 10056 14176 10376 15200
rect 10056 14112 10064 14176
rect 10128 14112 10144 14176
rect 10208 14112 10224 14176
rect 10288 14112 10304 14176
rect 10368 14112 10376 14176
rect 9443 13564 9509 13565
rect 9443 13500 9444 13564
rect 9508 13500 9509 13564
rect 9443 13499 9509 13500
rect 10056 13088 10376 14112
rect 10056 13024 10064 13088
rect 10128 13024 10144 13088
rect 10208 13024 10224 13088
rect 10288 13024 10304 13088
rect 10368 13024 10376 13088
rect 10056 12000 10376 13024
rect 10056 11936 10064 12000
rect 10128 11936 10144 12000
rect 10208 11936 10224 12000
rect 10288 11936 10304 12000
rect 10368 11936 10376 12000
rect 10056 10912 10376 11936
rect 10056 10848 10064 10912
rect 10128 10848 10144 10912
rect 10208 10848 10224 10912
rect 10288 10848 10304 10912
rect 10368 10848 10376 10912
rect 10056 9824 10376 10848
rect 10056 9760 10064 9824
rect 10128 9760 10144 9824
rect 10208 9760 10224 9824
rect 10288 9760 10304 9824
rect 10368 9760 10376 9824
rect 10056 8736 10376 9760
rect 10056 8672 10064 8736
rect 10128 8672 10144 8736
rect 10208 8672 10224 8736
rect 10288 8672 10304 8736
rect 10368 8672 10376 8736
rect 10056 7648 10376 8672
rect 10056 7584 10064 7648
rect 10128 7584 10144 7648
rect 10208 7584 10224 7648
rect 10288 7584 10304 7648
rect 10368 7584 10376 7648
rect 10056 6560 10376 7584
rect 10056 6496 10064 6560
rect 10128 6496 10144 6560
rect 10208 6496 10224 6560
rect 10288 6496 10304 6560
rect 10368 6496 10376 6560
rect 10056 5472 10376 6496
rect 10056 5408 10064 5472
rect 10128 5408 10144 5472
rect 10208 5408 10224 5472
rect 10288 5408 10304 5472
rect 10368 5408 10376 5472
rect 10056 4384 10376 5408
rect 10056 4320 10064 4384
rect 10128 4320 10144 4384
rect 10208 4320 10224 4384
rect 10288 4320 10304 4384
rect 10368 4320 10376 4384
rect 9075 3772 9141 3773
rect 9075 3708 9076 3772
rect 9140 3708 9141 3772
rect 9075 3707 9141 3708
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
rect 10056 3296 10376 4320
rect 10056 3232 10064 3296
rect 10128 3232 10144 3296
rect 10208 3232 10224 3296
rect 10288 3232 10304 3296
rect 10368 3232 10376 3296
rect 10056 2208 10376 3232
rect 10056 2144 10064 2208
rect 10128 2144 10144 2208
rect 10208 2144 10224 2208
rect 10288 2144 10304 2208
rect 10368 2144 10376 2208
rect 10056 1120 10376 2144
rect 10056 1056 10064 1120
rect 10128 1056 10144 1120
rect 10208 1056 10224 1120
rect 10288 1056 10304 1120
rect 10368 1056 10376 1120
rect 10056 496 10376 1056
rect 10716 14720 11036 15744
rect 10716 14656 10724 14720
rect 10788 14656 10804 14720
rect 10868 14656 10884 14720
rect 10948 14656 10964 14720
rect 11028 14656 11036 14720
rect 10716 13632 11036 14656
rect 10716 13568 10724 13632
rect 10788 13568 10804 13632
rect 10868 13568 10884 13632
rect 10948 13568 10964 13632
rect 11028 13568 11036 13632
rect 10716 12544 11036 13568
rect 10716 12480 10724 12544
rect 10788 12480 10804 12544
rect 10868 12480 10884 12544
rect 10948 12480 10964 12544
rect 11028 12480 11036 12544
rect 10716 11456 11036 12480
rect 10716 11392 10724 11456
rect 10788 11392 10804 11456
rect 10868 11392 10884 11456
rect 10948 11392 10964 11456
rect 11028 11392 11036 11456
rect 10716 10368 11036 11392
rect 10716 10304 10724 10368
rect 10788 10304 10804 10368
rect 10868 10304 10884 10368
rect 10948 10304 10964 10368
rect 11028 10304 11036 10368
rect 10716 9280 11036 10304
rect 11286 9485 11346 18803
rect 11283 9484 11349 9485
rect 11283 9420 11284 9484
rect 11348 9420 11349 9484
rect 11283 9419 11349 9420
rect 10716 9216 10724 9280
rect 10788 9216 10804 9280
rect 10868 9216 10884 9280
rect 10948 9216 10964 9280
rect 11028 9216 11036 9280
rect 10716 8192 11036 9216
rect 10716 8128 10724 8192
rect 10788 8128 10804 8192
rect 10868 8128 10884 8192
rect 10948 8128 10964 8192
rect 11028 8128 11036 8192
rect 10716 7104 11036 8128
rect 10716 7040 10724 7104
rect 10788 7040 10804 7104
rect 10868 7040 10884 7104
rect 10948 7040 10964 7104
rect 11028 7040 11036 7104
rect 10716 6016 11036 7040
rect 10716 5952 10724 6016
rect 10788 5952 10804 6016
rect 10868 5952 10884 6016
rect 10948 5952 10964 6016
rect 11028 5952 11036 6016
rect 10716 4928 11036 5952
rect 10716 4864 10724 4928
rect 10788 4864 10804 4928
rect 10868 4864 10884 4928
rect 10948 4864 10964 4928
rect 11028 4864 11036 4928
rect 10716 3840 11036 4864
rect 10716 3776 10724 3840
rect 10788 3776 10804 3840
rect 10868 3776 10884 3840
rect 10948 3776 10964 3840
rect 11028 3776 11036 3840
rect 10716 2752 11036 3776
rect 10716 2688 10724 2752
rect 10788 2688 10804 2752
rect 10868 2688 10884 2752
rect 10948 2688 10964 2752
rect 11028 2688 11036 2752
rect 10716 1664 11036 2688
rect 10716 1600 10724 1664
rect 10788 1600 10804 1664
rect 10868 1600 10884 1664
rect 10948 1600 10964 1664
rect 11028 1600 11036 1664
rect 10716 576 11036 1600
rect 10716 512 10724 576
rect 10788 512 10804 576
rect 10868 512 10884 576
rect 10948 512 10964 576
rect 11028 512 11036 576
rect 10716 496 11036 512
use sky130_fd_sc_hd__inv_2  _0824_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform -1 0 5704 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1757695336
transform -1 0 6900 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1757695336
transform -1 0 5612 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1757695336
transform -1 0 3588 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1757695336
transform -1 0 6900 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1757695336
transform 1 0 8648 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1757695336
transform 1 0 3036 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1757695336
transform -1 0 8464 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1757695336
transform 1 0 5428 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1757695336
transform -1 0 8648 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1757695336
transform -1 0 4140 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1757695336
transform -1 0 6624 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1757695336
transform 1 0 5796 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1757695336
transform -1 0 5704 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0838_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 1 0 5796 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5060 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0840_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4600 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0841_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5796 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4784 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_2  _0843_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4692 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0844_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 3404 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 1723858470
transform 1 0 2852 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 1723858470
transform 1 0 3220 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0847_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1104 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0849_
timestamp 1723858470
transform -1 0 3680 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1757695336
transform 1 0 920 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0851_
timestamp 1723858470
transform 1 0 1380 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0852_
timestamp 1723858470
transform 1 0 920 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0853_
timestamp 1723858470
transform -1 0 7728 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6808 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7452 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0856_
timestamp 1723858470
transform 1 0 5336 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6808 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 1 0 3220 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3956 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 1 0 4232 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0861_
timestamp 1757695336
transform 1 0 5060 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0862_
timestamp 1757695336
transform 1 0 2668 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 1 0 3496 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 2852 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _0865_
timestamp 1723858470
transform 1 0 1472 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1723858470
transform 1 0 5612 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0867_
timestamp 1723858470
transform 1 0 5796 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp 1757695336
transform 1 0 6256 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1723858470
transform -1 0 6256 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0870_
timestamp 1723858470
transform -1 0 7268 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1757695336
transform 1 0 5152 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0872_
timestamp 1723858470
transform 1 0 9016 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0873_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9476 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0874_
timestamp 1757695336
transform 1 0 3680 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0875_
timestamp 1723858470
transform 1 0 5244 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0876_
timestamp 1757695336
transform -1 0 6072 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0877_
timestamp 1757695336
transform -1 0 5612 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 1723858470
transform 1 0 7820 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0879_
timestamp 1723858470
transform 1 0 3680 0 -1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0880_
timestamp 1757695336
transform 1 0 7268 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1757695336
transform -1 0 5704 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0882_
timestamp 1757695336
transform -1 0 4232 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1723858470
transform 1 0 5796 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1723858470
transform -1 0 8188 0 1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0885_
timestamp 1757695336
transform 1 0 8372 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7728 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0887_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6532 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0888_
timestamp 1757695336
transform 1 0 8096 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0889_
timestamp 1757695336
transform -1 0 8004 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0890_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8096 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1723858470
transform -1 0 6992 0 1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0892_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6532 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0893_
timestamp 1723858470
transform 1 0 5796 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_2  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4876 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_4  _0895_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7176 0 1 41888
box -38 -48 1418 592
use sky130_fd_sc_hd__o21ai_2  _0896_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7176 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0897_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8004 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__a211oi_1  _0898_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7820 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0899_
timestamp 1757695336
transform 1 0 8004 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0900_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9108 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0901_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9108 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 1757695336
transform -1 0 8280 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0903_
timestamp 1723858470
transform 1 0 7820 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0904_
timestamp 1757695336
transform -1 0 5704 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0905_
timestamp 1723858470
transform 1 0 6072 0 1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _0906_
timestamp 1723858470
transform 1 0 6440 0 1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1723858470
transform 1 0 7360 0 1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1757695336
transform -1 0 8924 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0909_
timestamp 1723858470
transform 1 0 8372 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0910_
timestamp 1757695336
transform 1 0 6348 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0911_
timestamp 1723858470
transform 1 0 6900 0 -1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0912_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10396 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9292 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _0914_
timestamp 1723858470
transform -1 0 7452 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__or3b_1  _0915_
timestamp 1723858470
transform -1 0 8648 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7544 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _0917_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8096 0 -1 41888
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _0918_
timestamp 1723858470
transform 1 0 5244 0 1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0919_
timestamp 1757695336
transform 1 0 828 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0920_
timestamp 1723858470
transform 1 0 5796 0 -1 40800
box -38 -48 1234 592
use sky130_fd_sc_hd__or3b_1  _0921_
timestamp 1723858470
transform 1 0 6624 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0922_
timestamp 1723858470
transform 1 0 6900 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0923_
timestamp 1723858470
transform 1 0 5520 0 1 40800
box -38 -48 1234 592
use sky130_fd_sc_hd__or3b_1  _0924_
timestamp 1723858470
transform 1 0 6072 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0925_
timestamp 1723858470
transform -1 0 7452 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0926_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7268 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6808 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5612 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6164 0 -1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__nand2_1  _0930_
timestamp 1757695336
transform -1 0 8280 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1723858470
transform 1 0 5244 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1757695336
transform -1 0 7912 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0933_
timestamp 1757695336
transform 1 0 4968 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7452 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1757695336
transform -1 0 8556 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0936_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3220 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _0937_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3128 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0938_
timestamp 1757695336
transform -1 0 10856 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 1723858470
transform -1 0 9200 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0940_
timestamp 1757695336
transform -1 0 9568 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1723858470
transform -1 0 9292 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0942_
timestamp 1757695336
transform -1 0 10488 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1723858470
transform 1 0 8740 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0944_
timestamp 1757695336
transform -1 0 10856 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0945_
timestamp 1723858470
transform 1 0 10304 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _0946_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3220 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1757695336
transform -1 0 3128 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1723858470
transform 1 0 4416 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0949_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8372 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0950_
timestamp 1723858470
transform -1 0 8280 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0951_
timestamp 1757695336
transform -1 0 6808 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8924 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0953_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9384 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0954_
timestamp 1757695336
transform -1 0 3128 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0955_
timestamp 1723858470
transform 1 0 6532 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0956_
timestamp 1723858470
transform 1 0 5152 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _0957_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1196 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _0958_
timestamp 1723858470
transform 1 0 2300 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0959_
timestamp 1723858470
transform -1 0 4876 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0960_
timestamp 1723858470
transform 1 0 3220 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0961_
timestamp 1723858470
transform -1 0 10580 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9660 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0963_
timestamp 1757695336
transform -1 0 10120 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0964_
timestamp 1723858470
transform 1 0 10028 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0965_
timestamp 1723858470
transform -1 0 10764 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0966_
timestamp 1757695336
transform 1 0 10580 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0967_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4600 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0968_
timestamp 1723858470
transform 1 0 3956 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_4  _0969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4232 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__xnor2_1  _0970_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9844 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0971_
timestamp 1723858470
transform 1 0 9108 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0972_
timestamp 1757695336
transform 1 0 9752 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1723858470
transform 1 0 9936 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 1757695336
transform -1 0 10672 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0975_
timestamp 1723858470
transform -1 0 10856 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0976_
timestamp 1723858470
transform -1 0 10212 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0977_
timestamp 1723858470
transform -1 0 10396 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _0978_
timestamp 1723858470
transform -1 0 9384 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_2  _0979_
timestamp 1723858470
transform 1 0 6072 0 1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__a22o_1  _0980_
timestamp 1723858470
transform -1 0 7268 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0981_
timestamp 1723858470
transform 1 0 6164 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0982_
timestamp 1723858470
transform 1 0 5796 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0983_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4968 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0984_
timestamp 1723858470
transform 1 0 4692 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0985_
timestamp 1723858470
transform 1 0 2300 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _0986_
timestamp 1723858470
transform 1 0 1196 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _0987_
timestamp 1723858470
transform 1 0 1748 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0988_
timestamp 1723858470
transform -1 0 5060 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0989_
timestamp 1723858470
transform 1 0 2208 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0990_
timestamp 1723858470
transform 1 0 9384 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0991_
timestamp 1723858470
transform 1 0 9200 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0992_
timestamp 1723858470
transform -1 0 10672 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0993_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 10212 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0994_
timestamp 1723858470
transform 1 0 9660 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0995_
timestamp 1723858470
transform -1 0 10028 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0996_
timestamp 1723858470
transform 1 0 9936 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0997_
timestamp 1723858470
transform 1 0 9292 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0998_
timestamp 1723858470
transform -1 0 9936 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1757695336
transform -1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1000_
timestamp 1723858470
transform 1 0 9384 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1001_
timestamp 1757695336
transform 1 0 9568 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1002_
timestamp 1723858470
transform -1 0 10396 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1003_
timestamp 1757695336
transform -1 0 10764 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1004_
timestamp 1723858470
transform 1 0 10028 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1005_
timestamp 1757695336
transform 1 0 9844 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1723858470
transform 1 0 10396 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1757695336
transform -1 0 10396 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1008_
timestamp 1757695336
transform -1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1009_
timestamp 1723858470
transform 1 0 9568 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1010_
timestamp 1757695336
transform -1 0 10672 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1011_
timestamp 1723858470
transform -1 0 10672 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1012_
timestamp 1723858470
transform -1 0 10396 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1013_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9292 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1014_
timestamp 1723858470
transform 1 0 5888 0 -1 28832
box -38 -48 1694 592
use sky130_fd_sc_hd__o22a_1  _1015_
timestamp 1723858470
transform 1 0 5704 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1016_
timestamp 1723858470
transform -1 0 5704 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1017_
timestamp 1723858470
transform 1 0 4784 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1018_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4784 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1019_
timestamp 1757695336
transform -1 0 5336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1020_
timestamp 1723858470
transform 1 0 3404 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1021_
timestamp 1723858470
transform 1 0 1840 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1022_
timestamp 1723858470
transform 1 0 1196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1023_
timestamp 1723858470
transform 1 0 2392 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1024_
timestamp 1723858470
transform -1 0 5060 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1025_
timestamp 1723858470
transform 1 0 3220 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1026_
timestamp 1757695336
transform 1 0 7912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1027_
timestamp 1723858470
transform -1 0 7268 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1028_
timestamp 1723858470
transform 1 0 7820 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1029_
timestamp 1723858470
transform 1 0 9936 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1030_
timestamp 1723858470
transform 1 0 8648 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1031_
timestamp 1723858470
transform 1 0 8740 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1032_
timestamp 1723858470
transform -1 0 10672 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1033_
timestamp 1723858470
transform 1 0 9292 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1757695336
transform 1 0 8924 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1035_
timestamp 1723858470
transform -1 0 9660 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1036_
timestamp 1723858470
transform -1 0 9568 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1037_
timestamp 1723858470
transform -1 0 9016 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1038_
timestamp 1723858470
transform 1 0 9016 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1039_
timestamp 1723858470
transform 1 0 10120 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1040_
timestamp 1723858470
transform -1 0 10580 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1041_
timestamp 1757695336
transform 1 0 10580 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1042_
timestamp 1757695336
transform -1 0 10580 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1043_
timestamp 1723858470
transform 1 0 9844 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1044_
timestamp 1723858470
transform 1 0 9476 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1045_
timestamp 1757695336
transform 1 0 10580 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1046_
timestamp 1723858470
transform 1 0 9568 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1047_
timestamp 1723858470
transform 1 0 9200 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1048_
timestamp 1723858470
transform 1 0 8648 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_2  _1049_
timestamp 1723858470
transform 1 0 4416 0 1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__o22a_1  _1050_
timestamp 1723858470
transform 1 0 6256 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1051_
timestamp 1723858470
transform -1 0 5796 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1052_
timestamp 1723858470
transform 1 0 4784 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1053_
timestamp 1757695336
transform -1 0 4784 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1054_
timestamp 1723858470
transform 1 0 4692 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1055_
timestamp 1723858470
transform 1 0 3588 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1056_
timestamp 1723858470
transform 1 0 2300 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1057_
timestamp 1723858470
transform 1 0 1196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1058_
timestamp 1723858470
transform 1 0 2300 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1723858470
transform -1 0 4600 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1060_
timestamp 1723858470
transform 1 0 2852 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1061_
timestamp 1723858470
transform -1 0 7544 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1062_
timestamp 1723858470
transform 1 0 5520 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1063_
timestamp 1723858470
transform 1 0 6532 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1064_
timestamp 1723858470
transform 1 0 7820 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1065_
timestamp 1723858470
transform -1 0 8280 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1066_
timestamp 1723858470
transform 1 0 7176 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1067_
timestamp 1723858470
transform -1 0 9660 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _1068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8372 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1069_
timestamp 1723858470
transform -1 0 8188 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1070_
timestamp 1723858470
transform -1 0 9844 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1071_
timestamp 1757695336
transform 1 0 7820 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1072_
timestamp 1723858470
transform 1 0 8372 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1073_
timestamp 1723858470
transform 1 0 8832 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1074_
timestamp 1757695336
transform 1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1075_
timestamp 1723858470
transform 1 0 9568 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1076_
timestamp 1723858470
transform 1 0 9844 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1077_
timestamp 1757695336
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 1723858470
transform 1 0 10028 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1079_
timestamp 1757695336
transform -1 0 10856 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1080_
timestamp 1723858470
transform -1 0 10304 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1081_
timestamp 1723858470
transform -1 0 10212 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1082_
timestamp 1757695336
transform 1 0 10304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1083_
timestamp 1723858470
transform 1 0 9292 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1084_
timestamp 1723858470
transform 1 0 8740 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1085_
timestamp 1723858470
transform 1 0 8372 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_2  _1086_
timestamp 1723858470
transform 1 0 4692 0 1 26656
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1087_
timestamp 1723858470
transform 1 0 6900 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1088_
timestamp 1723858470
transform 1 0 7268 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1089_
timestamp 1757695336
transform 1 0 7636 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1090_
timestamp 1723858470
transform -1 0 8004 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1723858470
transform -1 0 7820 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1723858470
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1093_
timestamp 1723858470
transform 1 0 1012 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1094_
timestamp 1723858470
transform 1 0 1196 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1095_
timestamp 1723858470
transform -1 0 4600 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1723858470
transform -1 0 3404 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1097_
timestamp 1723858470
transform 1 0 828 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1098_
timestamp 1723858470
transform -1 0 4600 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1099_
timestamp 1723858470
transform -1 0 4968 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1100_
timestamp 1723858470
transform 1 0 4600 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1101_
timestamp 1723858470
transform -1 0 6532 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1102_
timestamp 1757695336
transform -1 0 5704 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1103_
timestamp 1723858470
transform 1 0 5796 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1104_
timestamp 1723858470
transform 1 0 7544 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1105_
timestamp 1723858470
transform 1 0 7176 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1106_
timestamp 1723858470
transform 1 0 6716 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1107_
timestamp 1723858470
transform 1 0 7084 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1108_
timestamp 1723858470
transform 1 0 7820 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1109_
timestamp 1723858470
transform -1 0 8740 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1110_
timestamp 1723858470
transform -1 0 8280 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1111_
timestamp 1723858470
transform -1 0 9936 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1112_
timestamp 1757695336
transform 1 0 9936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1113_
timestamp 1757695336
transform -1 0 8740 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1114_
timestamp 1723858470
transform 1 0 10212 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1115_
timestamp 1723858470
transform -1 0 9568 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1116_
timestamp 1757695336
transform -1 0 8280 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1117_
timestamp 1723858470
transform 1 0 7452 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1118_
timestamp 1723858470
transform -1 0 7360 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1119_
timestamp 1723858470
transform -1 0 6992 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1120_
timestamp 1723858470
transform -1 0 5428 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _1121_
timestamp 1723858470
transform 1 0 3220 0 1 28832
box -38 -48 1694 592
use sky130_fd_sc_hd__o22a_1  _1122_
timestamp 1723858470
transform 1 0 5060 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1123_
timestamp 1723858470
transform 1 0 3220 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1124_
timestamp 1723858470
transform -1 0 4600 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1125_
timestamp 1757695336
transform 1 0 4692 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1126_
timestamp 1723858470
transform 1 0 4048 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1127_
timestamp 1723858470
transform 1 0 2392 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1128_
timestamp 1723858470
transform 1 0 2392 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1129_
timestamp 1723858470
transform 1 0 1196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1130_
timestamp 1723858470
transform 1 0 2576 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1131_
timestamp 1723858470
transform -1 0 2392 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1132_
timestamp 1723858470
transform -1 0 2576 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1133_
timestamp 1723858470
transform -1 0 3128 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1134_
timestamp 1723858470
transform 1 0 920 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1135_
timestamp 1723858470
transform 1 0 1932 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1136_
timestamp 1723858470
transform -1 0 4324 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1723858470
transform 1 0 3312 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1138_
timestamp 1723858470
transform 1 0 3312 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _1139_
timestamp 1723858470
transform 1 0 4600 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1140_
timestamp 1723858470
transform 1 0 4692 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1141_
timestamp 1723858470
transform -1 0 5612 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1142_
timestamp 1723858470
transform -1 0 4876 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1143_
timestamp 1723858470
transform -1 0 6992 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1144_
timestamp 1757695336
transform 1 0 4508 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1145_
timestamp 1723858470
transform 1 0 5704 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1146_
timestamp 1757695336
transform 1 0 4324 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1147_
timestamp 1723858470
transform 1 0 5060 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1148_
timestamp 1757695336
transform -1 0 6716 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1149_
timestamp 1723858470
transform 1 0 4600 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1150_
timestamp 1757695336
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1151_
timestamp 1723858470
transform 1 0 8740 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1152_
timestamp 1723858470
transform 1 0 5060 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1153_
timestamp 1723858470
transform -1 0 6440 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1154_
timestamp 1723858470
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_2  _1155_
timestamp 1723858470
transform 1 0 2944 0 -1 29920
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1156_
timestamp 1723858470
transform 1 0 5060 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1157_
timestamp 1723858470
transform -1 0 5060 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1158_
timestamp 1723858470
transform 1 0 4600 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1159_
timestamp 1723858470
transform 1 0 4324 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1160_
timestamp 1723858470
transform 1 0 3588 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1161_
timestamp 1723858470
transform 1 0 2300 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1162_
timestamp 1723858470
transform 1 0 1472 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _1163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 1840 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1164_
timestamp 1757695336
transform -1 0 2116 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1723858470
transform -1 0 1288 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1166_
timestamp 1723858470
transform 1 0 828 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1167_
timestamp 1723858470
transform 1 0 1564 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1168_
timestamp 1723858470
transform 1 0 1472 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1169_
timestamp 1723858470
transform 1 0 920 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1170_
timestamp 1723858470
transform 1 0 1288 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1171_
timestamp 1723858470
transform 1 0 3772 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1172_
timestamp 1723858470
transform 1 0 3772 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1173_
timestamp 1723858470
transform -1 0 2852 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1174_
timestamp 1723858470
transform -1 0 5152 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1175_
timestamp 1723858470
transform 1 0 2484 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1176_
timestamp 1723858470
transform 1 0 5152 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1177_
timestamp 1723858470
transform 1 0 1840 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1178_
timestamp 1723858470
transform 1 0 3128 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1179_
timestamp 1723858470
transform 1 0 3220 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1180_
timestamp 1723858470
transform -1 0 4508 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1181_
timestamp 1723858470
transform 1 0 3404 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1723858470
transform -1 0 3036 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1183_
timestamp 1757695336
transform 1 0 4324 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1184_
timestamp 1723858470
transform -1 0 5428 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1185_
timestamp 1723858470
transform -1 0 5428 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1186_
timestamp 1723858470
transform 1 0 3680 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1187_
timestamp 1757695336
transform 1 0 7544 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1188_
timestamp 1723858470
transform -1 0 4692 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1189_
timestamp 1723858470
transform -1 0 5152 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1190_
timestamp 1723858470
transform 1 0 3220 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1191_
timestamp 1757695336
transform 1 0 2300 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1192_
timestamp 1723858470
transform 1 0 2392 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1193_
timestamp 1723858470
transform 1 0 828 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1194_
timestamp 1723858470
transform 1 0 2300 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1195_
timestamp 1723858470
transform -1 0 2300 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _1196_
timestamp 1723858470
transform -1 0 5336 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1197_
timestamp 1723858470
transform -1 0 9200 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1198_
timestamp 1723858470
transform 1 0 8372 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1199_
timestamp 1723858470
transform -1 0 7728 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1200_
timestamp 1757695336
transform -1 0 5704 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1201_
timestamp 1723858470
transform 1 0 7268 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1202_
timestamp 1723858470
transform 1 0 8096 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1203_
timestamp 1723858470
transform 1 0 7176 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1204_
timestamp 1723858470
transform -1 0 7912 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1205_
timestamp 1723858470
transform 1 0 5796 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _1206_
timestamp 1723858470
transform 1 0 1196 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1207_
timestamp 1757695336
transform -1 0 8648 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1208_
timestamp 1757695336
transform 1 0 10304 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1723858470
transform 1 0 9844 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _1210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10212 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1211_
timestamp 1723858470
transform 1 0 9476 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1723858470
transform -1 0 10212 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1213_
timestamp 1723858470
transform -1 0 9568 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1214_
timestamp 1723858470
transform -1 0 8832 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1215_
timestamp 1723858470
transform -1 0 10028 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1216_
timestamp 1723858470
transform 1 0 8464 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1217_
timestamp 1723858470
transform 1 0 8832 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _1218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8832 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1219_
timestamp 1723858470
transform 1 0 8096 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1723858470
transform -1 0 6348 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1221_
timestamp 1723858470
transform 1 0 6808 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1222_
timestamp 1723858470
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1223_
timestamp 1723858470
transform 1 0 7636 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1224_
timestamp 1723858470
transform 1 0 6440 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1225_
timestamp 1723858470
transform 1 0 4140 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1226_
timestamp 1723858470
transform 1 0 1932 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2484 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1228_
timestamp 1723858470
transform -1 0 8464 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1229_
timestamp 1723858470
transform -1 0 9844 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1230_
timestamp 1723858470
transform 1 0 8832 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1231_
timestamp 1723858470
transform -1 0 10672 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1723858470
transform -1 0 9752 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1233_
timestamp 1723858470
transform -1 0 8740 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1234_
timestamp 1757695336
transform 1 0 8740 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1235_
timestamp 1757695336
transform -1 0 8188 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1236_
timestamp 1723858470
transform -1 0 8740 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1237_
timestamp 1723858470
transform 1 0 8372 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1238_
timestamp 1723858470
transform 1 0 9660 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1239_
timestamp 1723858470
transform 1 0 8924 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1240_
timestamp 1723858470
transform 1 0 8648 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1241_
timestamp 1723858470
transform 1 0 8096 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1242_
timestamp 1723858470
transform -1 0 8280 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1243_
timestamp 1723858470
transform -1 0 7912 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1244_
timestamp 1723858470
transform 1 0 6992 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1245_
timestamp 1723858470
transform -1 0 9384 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1246_
timestamp 1723858470
transform 1 0 6348 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1247_
timestamp 1723858470
transform 1 0 2300 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1248_
timestamp 1723858470
transform -1 0 2852 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1249_
timestamp 1723858470
transform -1 0 1748 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1250_
timestamp 1723858470
transform 1 0 7360 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1251_
timestamp 1723858470
transform 1 0 8464 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1252_
timestamp 1757695336
transform 1 0 6624 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1253_
timestamp 1723858470
transform -1 0 7544 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1254_
timestamp 1723858470
transform 1 0 6624 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1255_
timestamp 1757695336
transform 1 0 7728 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1723858470
transform 1 0 6992 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1257_
timestamp 1757695336
transform 1 0 7452 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1258_
timestamp 1757695336
transform -1 0 5704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1259_
timestamp 1723858470
transform -1 0 6992 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1260_
timestamp 1757695336
transform -1 0 5980 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1261_
timestamp 1723858470
transform 1 0 7544 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1262_
timestamp 1723858470
transform 1 0 6348 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1263_
timestamp 1757695336
transform 1 0 7268 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1264_
timestamp 1723858470
transform 1 0 6716 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1265_
timestamp 1723858470
transform 1 0 6532 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1266_
timestamp 1723858470
transform 1 0 6164 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1723858470
transform -1 0 7360 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1268_
timestamp 1723858470
transform 1 0 6900 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1269_
timestamp 1723858470
transform 1 0 7360 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1270_
timestamp 1723858470
transform 1 0 8188 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1271_
timestamp 1723858470
transform 1 0 5888 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1272_
timestamp 1723858470
transform 1 0 3128 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1273_
timestamp 1723858470
transform 1 0 1288 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1274_
timestamp 1723858470
transform -1 0 1472 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1275_
timestamp 1723858470
transform 1 0 6072 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1276_
timestamp 1723858470
transform 1 0 5428 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1277_
timestamp 1723858470
transform 1 0 5336 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1278_
timestamp 1723858470
transform -1 0 6624 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1723858470
transform -1 0 6440 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1280_
timestamp 1723858470
transform 1 0 4324 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1281_
timestamp 1757695336
transform -1 0 5060 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 1757695336
transform 1 0 5152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1283_
timestamp 1723858470
transform 1 0 5980 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1284_
timestamp 1723858470
transform 1 0 4692 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1285_
timestamp 1723858470
transform 1 0 5796 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1286_
timestamp 1723858470
transform -1 0 5704 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1287_
timestamp 1723858470
transform -1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1288_
timestamp 1723858470
transform -1 0 6532 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1289_
timestamp 1723858470
transform -1 0 6900 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1290_
timestamp 1723858470
transform 1 0 6440 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1291_
timestamp 1723858470
transform 1 0 6348 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1292_
timestamp 1723858470
transform 1 0 7084 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1293_
timestamp 1723858470
transform 1 0 5796 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1294_
timestamp 1723858470
transform 1 0 3128 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1295_
timestamp 1723858470
transform 1 0 1564 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1296_
timestamp 1723858470
transform -1 0 1564 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1297_
timestamp 1757695336
transform -1 0 5152 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1298_
timestamp 1723858470
transform 1 0 4968 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1299_
timestamp 1757695336
transform 1 0 3036 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1300_
timestamp 1723858470
transform 1 0 3864 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1301_
timestamp 1757695336
transform -1 0 4600 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1302_
timestamp 1723858470
transform 1 0 3680 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1303_
timestamp 1757695336
transform 1 0 3220 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1304_
timestamp 1723858470
transform 1 0 3772 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1305_
timestamp 1757695336
transform -1 0 4324 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1306_
timestamp 1723858470
transform 1 0 4416 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1307_
timestamp 1723858470
transform 1 0 3772 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1308_
timestamp 1757695336
transform 1 0 4784 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1309_
timestamp 1723858470
transform -1 0 4784 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1311_
timestamp 1723858470
transform 1 0 3312 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1312_
timestamp 1723858470
transform 1 0 4692 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1313_
timestamp 1723858470
transform -1 0 5060 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1314_
timestamp 1723858470
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1315_
timestamp 1723858470
transform 1 0 2484 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1316_
timestamp 1723858470
transform 1 0 2300 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1317_
timestamp 1723858470
transform 1 0 1656 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _1318_
timestamp 1723858470
transform 1 0 1012 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1319_
timestamp 1723858470
transform -1 0 4692 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1320_
timestamp 1723858470
transform -1 0 5704 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1321_
timestamp 1757695336
transform 1 0 3588 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1322_
timestamp 1723858470
transform 1 0 3312 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1323_
timestamp 1757695336
transform -1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1324_
timestamp 1723858470
transform 1 0 1380 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1325_
timestamp 1757695336
transform -1 0 2668 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1326_
timestamp 1723858470
transform 1 0 1932 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1327_
timestamp 1757695336
transform -1 0 2668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1723858470
transform 1 0 1932 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1329_
timestamp 1757695336
transform -1 0 2944 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1330_
timestamp 1723858470
transform 1 0 3496 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1331_
timestamp 1723858470
transform 1 0 2024 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1332_
timestamp 1757695336
transform 1 0 3772 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1333_
timestamp 1723858470
transform 1 0 3220 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1334_
timestamp 1723858470
transform 1 0 2668 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1335_
timestamp 1723858470
transform 1 0 3496 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1336_
timestamp 1723858470
transform 1 0 2852 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1337_
timestamp 1723858470
transform 1 0 5796 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1338_
timestamp 1757695336
transform -1 0 5520 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1339_
timestamp 1757695336
transform -1 0 3496 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1340_
timestamp 1723858470
transform -1 0 3312 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1341_
timestamp 1723858470
transform 1 0 3220 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1342_
timestamp 1723858470
transform 1 0 1196 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1343_
timestamp 1757695336
transform 1 0 2576 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1344_
timestamp 1723858470
transform 1 0 2944 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1345_
timestamp 1723858470
transform 1 0 1840 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1346_
timestamp 1723858470
transform -1 0 1932 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1347_
timestamp 1723858470
transform 1 0 1840 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1348_
timestamp 1723858470
transform 1 0 1012 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1349_
timestamp 1723858470
transform 1 0 1196 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1350_
timestamp 1723858470
transform 1 0 1380 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1351_
timestamp 1757695336
transform -1 0 1932 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1352_
timestamp 1723858470
transform -1 0 3128 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1353_
timestamp 1723858470
transform 1 0 1932 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _1354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3036 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1355_
timestamp 1757695336
transform 1 0 2852 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1356_
timestamp 1723858470
transform 1 0 4784 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1357_
timestamp 1723858470
transform -1 0 4784 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1358_
timestamp 1723858470
transform 1 0 4416 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1359_
timestamp 1723858470
transform 1 0 2300 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1360_
timestamp 1723858470
transform 1 0 2024 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1361_
timestamp 1723858470
transform 1 0 1288 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1362_
timestamp 1723858470
transform 1 0 8740 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1363_
timestamp 1723858470
transform 1 0 8372 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1364_
timestamp 1757695336
transform -1 0 9200 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1365_
timestamp 1723858470
transform 1 0 8648 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1366_
timestamp 1757695336
transform -1 0 9752 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1367_
timestamp 1723858470
transform -1 0 9476 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1368_
timestamp 1757695336
transform 1 0 7636 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1369_
timestamp 1757695336
transform 1 0 7268 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1370_
timestamp 1723858470
transform 1 0 8372 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1371_
timestamp 1757695336
transform 1 0 9200 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1372_
timestamp 1723858470
transform 1 0 9108 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1373_
timestamp 1723858470
transform 1 0 9108 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1374_
timestamp 1723858470
transform 1 0 8648 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1375_
timestamp 1723858470
transform -1 0 4968 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1376_
timestamp 1723858470
transform 1 0 8372 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1377_
timestamp 1723858470
transform -1 0 8096 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1378_
timestamp 1723858470
transform -1 0 8280 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1379_
timestamp 1723858470
transform -1 0 7268 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1380_
timestamp 1723858470
transform 1 0 5152 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1381_
timestamp 1723858470
transform 1 0 1196 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1382_
timestamp 1757695336
transform 1 0 6624 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1383_
timestamp 1723858470
transform -1 0 6716 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1384_
timestamp 1757695336
transform -1 0 8648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1385_
timestamp 1723858470
transform -1 0 8280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1386_
timestamp 1723858470
transform 1 0 7084 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1387_
timestamp 1723858470
transform 1 0 7176 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1388_
timestamp 1723858470
transform -1 0 8096 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1389_
timestamp 1723858470
transform 1 0 7820 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1390_
timestamp 1723858470
transform 1 0 9016 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1391_
timestamp 1757695336
transform -1 0 9016 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1723858470
transform 1 0 7820 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1393_
timestamp 1723858470
transform 1 0 8372 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1394_
timestamp 1723858470
transform 1 0 7820 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1395_
timestamp 1723858470
transform 1 0 7268 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1396_
timestamp 1723858470
transform -1 0 6808 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1397_
timestamp 1723858470
transform 1 0 7084 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1398_
timestamp 1723858470
transform 1 0 6072 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1399_
timestamp 1723858470
transform 1 0 5336 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1400_
timestamp 1723858470
transform -1 0 6532 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1401_
timestamp 1723858470
transform 1 0 5060 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1402_
timestamp 1723858470
transform 1 0 2300 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1403_
timestamp 1723858470
transform 1 0 1196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1404_
timestamp 1757695336
transform -1 0 7176 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1405_
timestamp 1723858470
transform 1 0 5980 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1406_
timestamp 1757695336
transform -1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1407_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6716 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1408_
timestamp 1723858470
transform 1 0 6348 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1409_
timestamp 1723858470
transform 1 0 7268 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1410_
timestamp 1723858470
transform -1 0 7452 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1411_
timestamp 1723858470
transform 1 0 6348 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1412_
timestamp 1723858470
transform 1 0 6808 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1413_
timestamp 1757695336
transform 1 0 8096 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1414_
timestamp 1723858470
transform 1 0 7544 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1415_
timestamp 1723858470
transform 1 0 6992 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1416_
timestamp 1723858470
transform 1 0 5796 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1417_
timestamp 1723858470
transform 1 0 6256 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1418_
timestamp 1757695336
transform -1 0 9200 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1419_
timestamp 1723858470
transform -1 0 7452 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1420_
timestamp 1723858470
transform -1 0 8004 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1421_
timestamp 1723858470
transform 1 0 2576 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1422_
timestamp 1723858470
transform 1 0 1472 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _1423_
timestamp 1723858470
transform -1 0 1840 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1424_
timestamp 1723858470
transform 1 0 4324 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1425_
timestamp 1757695336
transform -1 0 4876 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1426_
timestamp 1757695336
transform -1 0 5060 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1427_
timestamp 1723858470
transform 1 0 5796 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1428_
timestamp 1723858470
transform 1 0 5060 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1429_
timestamp 1723858470
transform 1 0 4968 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1430_
timestamp 1723858470
transform -1 0 6348 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1431_
timestamp 1723858470
transform 1 0 5428 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1432_
timestamp 1723858470
transform 1 0 6440 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1433_
timestamp 1723858470
transform -1 0 6440 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1434_
timestamp 1757695336
transform -1 0 6164 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1435_
timestamp 1723858470
transform 1 0 5336 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1436_
timestamp 1723858470
transform 1 0 5336 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1437_
timestamp 1723858470
transform 1 0 6440 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1438_
timestamp 1723858470
transform -1 0 7360 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1439_
timestamp 1723858470
transform 1 0 5796 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1440_
timestamp 1723858470
transform -1 0 6164 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1441_
timestamp 1723858470
transform 1 0 4784 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1442_
timestamp 1723858470
transform 1 0 2300 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1443_
timestamp 1723858470
transform 1 0 1196 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1444_
timestamp 1723858470
transform 1 0 4876 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1445_
timestamp 1723858470
transform 1 0 2300 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1446_
timestamp 1723858470
transform -1 0 4232 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1447_
timestamp 1723858470
transform 1 0 3312 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1448_
timestamp 1723858470
transform 1 0 3220 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1449_
timestamp 1723858470
transform 1 0 4324 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1450_
timestamp 1757695336
transform -1 0 3036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1451_
timestamp 1723858470
transform 1 0 3404 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1452_
timestamp 1757695336
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1453_
timestamp 1723858470
transform 1 0 3036 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1454_
timestamp 1723858470
transform 1 0 3680 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1455_
timestamp 1723858470
transform 1 0 5152 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1456_
timestamp 1723858470
transform 1 0 5796 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1457_
timestamp 1723858470
transform -1 0 6256 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1458_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5796 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1459_
timestamp 1723858470
transform 1 0 5612 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1460_
timestamp 1723858470
transform 1 0 3680 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1461_
timestamp 1723858470
transform -1 0 2116 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1462_
timestamp 1723858470
transform 1 0 1196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1463_
timestamp 1723858470
transform 1 0 2760 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1464_
timestamp 1723858470
transform -1 0 2668 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1465_
timestamp 1723858470
transform -1 0 1840 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1466_
timestamp 1723858470
transform -1 0 1288 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1467_
timestamp 1723858470
transform 1 0 1288 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1468_
timestamp 1757695336
transform -1 0 1472 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1469_
timestamp 1723858470
transform 1 0 1748 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1470_
timestamp 1757695336
transform -1 0 3036 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1471_
timestamp 1723858470
transform -1 0 3772 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1472_
timestamp 1723858470
transform 1 0 1472 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1473_
timestamp 1723858470
transform 1 0 2116 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1474_
timestamp 1723858470
transform -1 0 3772 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1475_
timestamp 1723858470
transform 1 0 3036 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1476_
timestamp 1723858470
transform 1 0 4140 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1477_
timestamp 1723858470
transform -1 0 4692 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1478_
timestamp 1723858470
transform -1 0 3588 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1479_
timestamp 1723858470
transform -1 0 3864 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1480_
timestamp 1723858470
transform -1 0 5336 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1481_
timestamp 1723858470
transform -1 0 2852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1482_
timestamp 1723858470
transform 1 0 828 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1483_
timestamp 1723858470
transform 1 0 1196 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _1484_
timestamp 1723858470
transform 1 0 1748 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1485_
timestamp 1723858470
transform -1 0 2300 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1486_
timestamp 1723858470
transform 1 0 1196 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1487_
timestamp 1723858470
transform 1 0 1840 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1488_
timestamp 1723858470
transform -1 0 3128 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1489_
timestamp 1723858470
transform 1 0 2116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1490_
timestamp 1723858470
transform 1 0 3680 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1491_
timestamp 1723858470
transform -1 0 4508 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1492_
timestamp 1723858470
transform 1 0 3220 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1493_
timestamp 1723858470
transform 1 0 2392 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1494_
timestamp 1723858470
transform 1 0 2576 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1495_
timestamp 1723858470
transform -1 0 2668 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1496_
timestamp 1723858470
transform 1 0 3772 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1497_
timestamp 1723858470
transform 1 0 1196 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1498_
timestamp 1723858470
transform 1 0 2484 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1499_
timestamp 1723858470
transform 1 0 1656 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _1500_
timestamp 1723858470
transform -1 0 5060 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1501_
timestamp 1757695336
transform 1 0 2484 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1502_
timestamp 1757695336
transform -1 0 2484 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1503_
timestamp 1723858470
transform 1 0 828 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1504_
timestamp 1723858470
transform 1 0 1472 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1505_
timestamp 1757695336
transform 1 0 3036 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1506_
timestamp 1723858470
transform 1 0 1196 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1507_
timestamp 1723858470
transform -1 0 3128 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1508_
timestamp 1723858470
transform -1 0 2300 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 1723858470
transform -1 0 3956 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1510_
timestamp 1723858470
transform -1 0 4416 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1511_
timestamp 1723858470
transform 1 0 828 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1512_
timestamp 1723858470
transform -1 0 3036 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1513_
timestamp 1757695336
transform 1 0 828 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1514_
timestamp 1723858470
transform 1 0 3220 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1515_
timestamp 1723858470
transform 1 0 828 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1516_
timestamp 1723858470
transform -1 0 2300 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _1517_
timestamp 1723858470
transform 1 0 1012 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1518_
timestamp 1723858470
transform 1 0 4232 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1519_
timestamp 1723858470
transform 1 0 3496 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1520_
timestamp 1723858470
transform 1 0 1932 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1723858470
transform -1 0 2852 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 1723858470
transform 1 0 1380 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1523_
timestamp 1723858470
transform 1 0 8648 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1524_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9936 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1525_
timestamp 1723858470
transform 1 0 8096 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1526_
timestamp 1723858470
transform -1 0 9752 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1527_
timestamp 1723858470
transform -1 0 10672 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1528_
timestamp 1723858470
transform -1 0 8280 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1529_
timestamp 1723858470
transform 1 0 6992 0 1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1530_
timestamp 1723858470
transform 1 0 9016 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1531_
timestamp 1757695336
transform -1 0 9200 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1532_
timestamp 1723858470
transform 1 0 8280 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1533_
timestamp 1723858470
transform 1 0 9936 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8372 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1535_
timestamp 1723858470
transform -1 0 8188 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1536_
timestamp 1723858470
transform -1 0 10212 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1537_
timestamp 1723858470
transform 1 0 6624 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _1538_
timestamp 1723858470
transform -1 0 9200 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1539_
timestamp 1723858470
transform 1 0 7360 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1540_
timestamp 1723858470
transform 1 0 7636 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1541_
timestamp 1723858470
transform -1 0 9384 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1542_
timestamp 1723858470
transform 1 0 8372 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1543_
timestamp 1723858470
transform -1 0 6440 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1544_
timestamp 1723858470
transform -1 0 1380 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1545_
timestamp 1723858470
transform -1 0 5704 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1546_
timestamp 1723858470
transform 1 0 6348 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1547_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8740 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1548_
timestamp 1723858470
transform 1 0 6992 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1549_
timestamp 1757695336
transform -1 0 8648 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1550_
timestamp 1723858470
transform 1 0 6992 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1551_
timestamp 1757695336
transform -1 0 10856 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1552_
timestamp 1723858470
transform 1 0 8096 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1553_
timestamp 1757695336
transform -1 0 7176 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1554_
timestamp 1723858470
transform 1 0 8556 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1555_
timestamp 1723858470
transform 1 0 9200 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1556_
timestamp 1723858470
transform -1 0 9200 0 1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1557_
timestamp 1723858470
transform 1 0 9200 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1558_
timestamp 1723858470
transform -1 0 10120 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1559_
timestamp 1757695336
transform -1 0 8648 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1560_
timestamp 1723858470
transform 1 0 8924 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1561_
timestamp 1723858470
transform -1 0 10580 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1562_
timestamp 1723858470
transform 1 0 9108 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1563_
timestamp 1723858470
transform -1 0 10672 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1564_
timestamp 1723858470
transform 1 0 10028 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1565_
timestamp 1723858470
transform 1 0 9384 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1566_
timestamp 1757695336
transform -1 0 5152 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1567_
timestamp 1723858470
transform 1 0 10120 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1568_
timestamp 1723858470
transform -1 0 10488 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1569_
timestamp 1723858470
transform 1 0 8740 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1570_
timestamp 1757695336
transform -1 0 3128 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1571_
timestamp 1723858470
transform -1 0 9292 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1572_
timestamp 1723858470
transform -1 0 8648 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1573_
timestamp 1723858470
transform 1 0 6992 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1574_
timestamp 1723858470
transform 1 0 8004 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1575_
timestamp 1723858470
transform -1 0 8740 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1576_
timestamp 1723858470
transform -1 0 8004 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1577_
timestamp 1757695336
transform -1 0 6716 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1578_
timestamp 1723858470
transform 1 0 6624 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1579_
timestamp 1723858470
transform 1 0 5612 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6256 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1581_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6900 0 -1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1582_
timestamp 1723858470
transform -1 0 7728 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1583_
timestamp 1723858470
transform 1 0 5888 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1584_
timestamp 1723858470
transform -1 0 6992 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1585_
timestamp 1723858470
transform 1 0 7728 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1586_
timestamp 1723858470
transform 1 0 7728 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1587_
timestamp 1723858470
transform 1 0 5980 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1588_
timestamp 1723858470
transform -1 0 5980 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1589_
timestamp 1723858470
transform 1 0 3864 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1590_
timestamp 1723858470
transform 1 0 828 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1591_
timestamp 1723858470
transform 1 0 1380 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1592_
timestamp 1723858470
transform 1 0 5152 0 1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _1593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4508 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1594_
timestamp 1723858470
transform -1 0 3956 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1595_
timestamp 1723858470
transform 1 0 4508 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1596_
timestamp 1723858470
transform 1 0 4508 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1597_
timestamp 1723858470
transform -1 0 5704 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1598_
timestamp 1723858470
transform 1 0 4232 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1599_
timestamp 1723858470
transform -1 0 6072 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1600_
timestamp 1723858470
transform 1 0 4232 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1601_
timestamp 1723858470
transform 1 0 4784 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1602_
timestamp 1723858470
transform 1 0 5796 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1603_
timestamp 1723858470
transform 1 0 3404 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1604_
timestamp 1723858470
transform 1 0 4140 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1605_
timestamp 1723858470
transform 1 0 1656 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1606_
timestamp 1723858470
transform 1 0 4048 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1723858470
transform 1 0 8372 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1608_
timestamp 1723858470
transform -1 0 3680 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp 1723858470
transform -1 0 1656 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1610_
timestamp 1723858470
transform 1 0 4876 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1611_
timestamp 1723858470
transform 1 0 8188 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1612_
timestamp 1723858470
transform -1 0 10764 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8280 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1614_
timestamp 1723858470
transform 1 0 8740 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1615_
timestamp 1723858470
transform 1 0 8280 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1616_
timestamp 1757695336
transform 1 0 10488 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1617_
timestamp 1723858470
transform 1 0 9844 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1618_
timestamp 1723858470
transform 1 0 9200 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1619_
timestamp 1723858470
transform -1 0 8280 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1620_
timestamp 1723858470
transform 1 0 9660 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1621_
timestamp 1723858470
transform -1 0 9200 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1622_
timestamp 1723858470
transform 1 0 9016 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1623_
timestamp 1723858470
transform -1 0 9108 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1624_
timestamp 1723858470
transform -1 0 8280 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1625_
timestamp 1723858470
transform 1 0 8372 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1626_
timestamp 1723858470
transform 1 0 8372 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1627_
timestamp 1757695336
transform 1 0 7912 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1628_
timestamp 1723858470
transform -1 0 9936 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1629_
timestamp 1723858470
transform 1 0 7268 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1630_
timestamp 1723858470
transform -1 0 7452 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1631_
timestamp 1723858470
transform 1 0 6532 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1632_
timestamp 1723858470
transform 1 0 3312 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1633_
timestamp 1723858470
transform 1 0 2392 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1634_
timestamp 1723858470
transform 1 0 3404 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1635_
timestamp 1723858470
transform 1 0 2208 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1636_
timestamp 1757695336
transform -1 0 2392 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1637_
timestamp 1723858470
transform -1 0 3680 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1638_
timestamp 1723858470
transform -1 0 3312 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1639_
timestamp 1723858470
transform -1 0 2668 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1640_
timestamp 1723858470
transform 1 0 2484 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1641_
timestamp 1723858470
transform 1 0 1104 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1642_
timestamp 1723858470
transform 1 0 1196 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1643_
timestamp 1723858470
transform -1 0 2208 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _1644_
timestamp 1723858470
transform -1 0 1932 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1645_
timestamp 1723858470
transform 1 0 8832 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1646_
timestamp 1723858470
transform 1 0 9292 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1647_
timestamp 1723858470
transform -1 0 10672 0 1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1648_
timestamp 1723858470
transform -1 0 10764 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1649_
timestamp 1723858470
transform -1 0 10580 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1650_
timestamp 1757695336
transform 1 0 10580 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1651_
timestamp 1723858470
transform 1 0 9752 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1652_
timestamp 1723858470
transform 1 0 9108 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1653_
timestamp 1723858470
transform 1 0 10396 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1654_
timestamp 1723858470
transform -1 0 10396 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1655_
timestamp 1723858470
transform -1 0 3588 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1656_
timestamp 1723858470
transform -1 0 4140 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1657_
timestamp 1723858470
transform 1 0 3588 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1658_
timestamp 1723858470
transform 1 0 1380 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1659_
timestamp 1723858470
transform 1 0 2760 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1660_
timestamp 1723858470
transform 1 0 1380 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1661_
timestamp 1757695336
transform -1 0 3496 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1662_
timestamp 1723858470
transform -1 0 1472 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1663_
timestamp 1723858470
transform 1 0 2484 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1664_
timestamp 1723858470
transform 1 0 920 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1665_
timestamp 1723858470
transform -1 0 2944 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1666_
timestamp 1757695336
transform 1 0 2852 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1667_
timestamp 1723858470
transform -1 0 3128 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1668_
timestamp 1723858470
transform 1 0 920 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _1669_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3864 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1670_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1012 0 -1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1671_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1196 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1723858470
transform 1 0 2116 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1673_
timestamp 1723858470
transform 1 0 3128 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1674_
timestamp 1723858470
transform 1 0 1288 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1675_
timestamp 1723858470
transform -1 0 2760 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1723858470
transform 1 0 1288 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1723858470
transform -1 0 7176 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1723858470
transform 1 0 8648 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1679_
timestamp 1723858470
transform -1 0 10856 0 -1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1723858470
transform 1 0 9384 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1723858470
transform 1 0 9200 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1723858470
transform 1 0 9384 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1683_
timestamp 1723858470
transform 1 0 9292 0 1 40800
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1684_
timestamp 1723858470
transform 1 0 8648 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1685_
timestamp 1723858470
transform -1 0 10120 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1686_
timestamp 1723858470
transform 1 0 8372 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1687_
timestamp 1723858470
transform -1 0 8280 0 1 40800
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1688_
timestamp 1723858470
transform -1 0 7268 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1723858470
transform 1 0 4324 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1723858470
transform 1 0 3956 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1723858470
transform 1 0 3956 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1723858470
transform -1 0 5520 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1723858470
transform 1 0 3772 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1723858470
transform 1 0 3680 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1723858470
transform 1 0 3680 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1723858470
transform -1 0 5060 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1723858470
transform 1 0 9384 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1723858470
transform -1 0 10856 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1723858470
transform 1 0 9200 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1700_
timestamp 1723858470
transform 1 0 9384 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1701_
timestamp 1723858470
transform 1 0 9016 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1702_
timestamp 1723858470
transform -1 0 9476 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1723858470
transform 1 0 6532 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1723858470
transform 1 0 3772 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1723858470
transform -1 0 4324 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1723858470
transform -1 0 3128 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1723858470
transform 1 0 1012 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1723858470
transform 1 0 1840 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1723858470
transform 1 0 1380 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1723858470
transform 1 0 1472 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1723858470
transform 1 0 1656 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1723858470
transform 1 0 1564 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1723858470
transform 1 0 1656 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1723858470
transform -1 0 10856 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1723858470
transform -1 0 10396 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1723858470
transform -1 0 10580 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1723858470
transform -1 0 10856 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1723858470
transform -1 0 10212 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1723858470
transform 1 0 3772 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1723858470
transform -1 0 2300 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1723858470
transform 1 0 920 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1723858470
transform 1 0 2392 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1723858470
transform 1 0 3220 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1723858470
transform 1 0 1288 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1725_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 1656 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1726_
timestamp 1723858470
transform -1 0 1656 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1727_
timestamp 1723858470
transform -1 0 2024 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1728_
timestamp 1723858470
transform -1 0 1196 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1729_
timestamp 1723858470
transform -1 0 1196 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1730_
timestamp 1723858470
transform 1 0 1840 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1731_
timestamp 1723858470
transform -1 0 1380 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1732_
timestamp 1723858470
transform 1 0 2760 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1733_
timestamp 1723858470
transform -1 0 1196 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1734_
timestamp 1723858470
transform -1 0 1196 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1735_
timestamp 1723858470
transform -1 0 1380 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1736_
timestamp 1723858470
transform 1 0 2760 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1737_
timestamp 1723858470
transform 1 0 2300 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1738_
timestamp 1723858470
transform 1 0 1932 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1739_
timestamp 1723858470
transform 1 0 3220 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1740_
timestamp 1723858470
transform -1 0 1196 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1741_
timestamp 1723858470
transform -1 0 1288 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1742_
timestamp 1723858470
transform -1 0 1288 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1743_
timestamp 1723858470
transform -1 0 1564 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7636 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1723858470
transform 1 0 8464 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1723858470
transform 1 0 8372 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1723858470
transform -1 0 5152 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1723858470
transform -1 0 5428 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_8  clkload0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8464 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__clkinvlp_4  clkload1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8280 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  clkload2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3220 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  fanout10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7452 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 1723858470
transform -1 0 4968 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1723858470
transform 1 0 6532 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1723858470
transform 1 0 8372 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8096 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout16
timestamp 1723858470
transform 1 0 8280 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1723858470
transform -1 0 8096 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7176 0 1 24480
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1723858470
transform 1 0 8832 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1723858470
transform 1 0 6164 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1723858470
transform -1 0 3128 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1723858470
transform 1 0 5796 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1723858470
transform -1 0 2576 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1723858470
transform 1 0 1104 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1723858470
transform 1 0 828 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1723858470
transform 1 0 8372 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1723858470
transform -1 0 5704 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout28
timestamp 1723858470
transform 1 0 4968 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1723858470
transform 1 0 2300 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1723858470
transform 1 0 9476 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1723858470
transform -1 0 1472 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 1723858470
transform -1 0 1196 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1723858470
transform -1 0 8004 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 1723858470
transform 1 0 10212 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 1723858470
transform -1 0 4324 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1723858470
transform 1 0 7636 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp 1723858470
transform 1 0 2944 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1723858470
transform 1 0 9292 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 1723858470
transform 1 0 10396 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout40
timestamp 1723858470
transform -1 0 8372 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 1723858470
transform 1 0 6716 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1723858470
transform 1 0 9384 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1723858470
transform -1 0 8096 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1723858470
transform -1 0 3680 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1723858470
transform -1 0 1196 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 1723858470
transform 1 0 5336 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1723858470
transform 1 0 5244 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp 1723858470
transform 1 0 828 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1723858470
transform -1 0 2300 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1723858470
transform 1 0 3036 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1723858470
transform -1 0 1748 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1723858470
transform 1 0 7176 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp 1723858470
transform -1 0 5888 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout54
timestamp 1723858470
transform 1 0 10028 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1723858470
transform -1 0 3772 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp 1723858470
transform -1 0 9108 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 1723858470
transform -1 0 9108 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout58
timestamp 1723858470
transform 1 0 10396 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 1723858470
transform 1 0 10212 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 1723858470
transform 1 0 8372 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 1723858470
transform 1 0 7912 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout62
timestamp 1723858470
transform -1 0 8740 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout63
timestamp 1723858470
transform -1 0 10028 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout64
timestamp 1723858470
transform -1 0 8740 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout65
timestamp 1723858470
transform -1 0 7820 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 1723858470
transform 1 0 3220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp 1723858470
transform -1 0 4692 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout68
timestamp 1723858470
transform -1 0 4416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 1723858470
transform 1 0 8280 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 1723858470
transform 1 0 7728 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp 1723858470
transform -1 0 9200 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout72
timestamp 1723858470
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 1723858470
transform 1 0 10488 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp 1723858470
transform 1 0 9476 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp 1723858470
transform -1 0 9476 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 1723858470
transform -1 0 10120 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout77
timestamp 1723858470
transform -1 0 10856 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp 1723858470
transform -1 0 8280 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp 1723858470
transform -1 0 8188 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 1723858470
transform 1 0 10488 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout81
timestamp 1723858470
transform 1 0 1012 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp 1723858470
transform 1 0 3220 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 1723858470
transform 1 0 5244 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout84
timestamp 1723858470
transform 1 0 9844 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout85
timestamp 1723858470
transform 1 0 8004 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout86 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8004 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout87
timestamp 1723858470
transform -1 0 10856 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout88
timestamp 1723858470
transform 1 0 7912 0 1 39712
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1723858470
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34
timestamp 1723858470
transform 1 0 3680 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4784 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5520 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1723858470
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1723858470
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1723858470
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1723858470
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1723858470
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1723858470
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1723858470
transform 1 0 1932 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_45
timestamp 1723858470
transform 1 0 4692 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1723858470
transform 1 0 5428 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1723858470
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1723858470
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1723858470
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1723858470
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1723858470
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 828 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1723858470
transform 1 0 3220 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_51
timestamp 1723858470
transform 1 0 5244 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_63
timestamp 1723858470
transform 1 0 6348 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_72
timestamp 1723858470
transform 1 0 7176 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1723858470
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_94
timestamp 1723858470
transform 1 0 9200 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_106
timestamp 1723858470
transform 1 0 10304 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1723858470
transform 1 0 828 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1723858470
transform 1 0 3312 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_42
timestamp 1723858470
transform 1 0 4416 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1723858470
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1723858470
transform 1 0 5796 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_102
timestamp 1723858470
transform 1 0 9936 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1723858470
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1723858470
transform 1 0 828 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_33
timestamp 1723858470
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1723858470
transform 1 0 4692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_59
timestamp 1723858470
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_67
timestamp 1723858470
transform 1 0 6716 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_75
timestamp 1723858470
transform 1 0 7452 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1723858470
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp 1723858470
transform 1 0 1932 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1723858470
transform 1 0 2668 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1723858470
transform 1 0 3036 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_35
timestamp 1723858470
transform 1 0 3772 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_67
timestamp 1723858470
transform 1 0 6716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_101
timestamp 1723858470
transform 1 0 9844 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1723858470
transform 1 0 10580 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1723858470
transform 1 0 828 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_61
timestamp 1723858470
transform 1 0 6164 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_65
timestamp 1723858470
transform 1 0 6532 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_70
timestamp 1723858470
transform 1 0 6992 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_78
timestamp 1723858470
transform 1 0 7728 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1723858470
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1723858470
transform 1 0 8372 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_105
timestamp 1723858470
transform 1 0 10212 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_111
timestamp 1723858470
transform 1 0 10764 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_40
timestamp 1723858470
transform 1 0 4232 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1723858470
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1723858470
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_69
timestamp 1723858470
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_78
timestamp 1723858470
transform 1 0 7728 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_89
timestamp 1723858470
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1723858470
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1723858470
transform 1 0 828 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1723858470
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1723858470
transform 1 0 2668 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1723858470
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_36
timestamp 1723858470
transform 1 0 3864 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp 1723858470
transform 1 0 4600 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_75
timestamp 1723858470
transform 1 0 7452 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1723858470
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_111
timestamp 1723858470
transform 1 0 10764 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1723858470
transform 1 0 828 0 -1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1723858470
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1723858470
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1723858470
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1723858470
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_64
timestamp 1723858470
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_84
timestamp 1723858470
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_92
timestamp 1723858470
transform 1 0 9016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1723858470
transform 1 0 828 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1723858470
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1723858470
transform 1 0 2484 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1723858470
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_38
timestamp 1723858470
transform 1 0 4048 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_49
timestamp 1723858470
transform 1 0 5060 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_58
timestamp 1723858470
transform 1 0 5888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1723858470
transform 1 0 7360 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1723858470
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1723858470
transform 1 0 8372 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_95
timestamp 1723858470
transform 1 0 9292 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_107
timestamp 1723858470
transform 1 0 10396 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_111
timestamp 1723858470
transform 1 0 10764 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1723858470
transform 1 0 828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_85
timestamp 1723858470
transform 1 0 8372 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1723858470
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_101
timestamp 1723858470
transform 1 0 9844 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1723858470
transform 1 0 10580 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1723858470
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1723858470
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_36
timestamp 1723858470
transform 1 0 3864 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_47
timestamp 1723858470
transform 1 0 4876 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_51
timestamp 1723858470
transform 1 0 5244 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_64
timestamp 1723858470
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1723858470
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1723858470
transform 1 0 8372 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_109
timestamp 1723858470
transform 1 0 10580 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1723858470
transform 1 0 828 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1723858470
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1723858470
transform 1 0 2668 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_35
timestamp 1723858470
transform 1 0 3772 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1723858470
transform 1 0 4876 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1723858470
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1723858470
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_61
timestamp 1723858470
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1723858470
transform 1 0 828 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1723858470
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_17
timestamp 1723858470
transform 1 0 2116 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1723858470
transform 1 0 2852 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_29
timestamp 1723858470
transform 1 0 3220 0 1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_40
timestamp 1723858470
transform 1 0 4232 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_52
timestamp 1723858470
transform 1 0 5336 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_64
timestamp 1723858470
transform 1 0 6440 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_70
timestamp 1723858470
transform 1 0 6992 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_78
timestamp 1723858470
transform 1 0 7728 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_92
timestamp 1723858470
transform 1 0 9016 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1723858470
transform 1 0 828 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1723858470
transform 1 0 1196 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_23
timestamp 1723858470
transform 1 0 2668 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1723858470
transform 1 0 5060 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1723858470
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1723858470
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1723858470
transform 1 0 6900 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_86
timestamp 1723858470
transform 1 0 8464 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_100
timestamp 1723858470
transform 1 0 9752 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1723858470
transform 1 0 828 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1723858470
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1723858470
transform 1 0 3220 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_60
timestamp 1723858470
transform 1 0 6072 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_69
timestamp 1723858470
transform 1 0 6900 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1723858470
transform 1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_99
timestamp 1723858470
transform 1 0 9660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1723858470
transform 1 0 10396 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1723858470
transform 1 0 10764 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1723858470
transform 1 0 828 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_20
timestamp 1723858470
transform 1 0 2392 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_26
timestamp 1723858470
transform 1 0 2944 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_44
timestamp 1723858470
transform 1 0 4600 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1723858470
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_64
timestamp 1723858470
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_76
timestamp 1723858470
transform 1 0 7544 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_95
timestamp 1723858470
transform 1 0 9292 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1723858470
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1723858470
transform 1 0 828 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1723858470
transform 1 0 2668 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1723858470
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1723858470
transform 1 0 3220 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_33
timestamp 1723858470
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_41
timestamp 1723858470
transform 1 0 4324 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_47
timestamp 1723858470
transform 1 0 4876 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_52
timestamp 1723858470
transform 1 0 5336 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1723858470
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1723858470
transform 1 0 8372 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_94
timestamp 1723858470
transform 1 0 9200 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_101
timestamp 1723858470
transform 1 0 9844 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_109
timestamp 1723858470
transform 1 0 10580 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1723858470
transform 1 0 828 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1723858470
transform 1 0 1564 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_28
timestamp 1723858470
transform 1 0 3128 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_49
timestamp 1723858470
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1723858470
transform 1 0 6256 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_70
timestamp 1723858470
transform 1 0 6992 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1723858470
transform 1 0 8096 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1723858470
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_97
timestamp 1723858470
transform 1 0 9476 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1723858470
transform 1 0 10396 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1723858470
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1723858470
transform 1 0 828 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1723858470
transform 1 0 1196 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_16
timestamp 1723858470
transform 1 0 2024 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1723858470
transform 1 0 2852 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_38
timestamp 1723858470
transform 1 0 4048 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_50
timestamp 1723858470
transform 1 0 5152 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_62
timestamp 1723858470
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1723858470
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_76
timestamp 1723858470
transform 1 0 7544 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_100
timestamp 1723858470
transform 1 0 9752 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1723858470
transform 1 0 828 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1723858470
transform 1 0 1196 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_12
timestamp 1723858470
transform 1 0 1656 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_37
timestamp 1723858470
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1723858470
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1723858470
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_64
timestamp 1723858470
transform 1 0 6440 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1723858470
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_92
timestamp 1723858470
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1723858470
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1723858470
transform 1 0 828 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_17
timestamp 1723858470
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1723858470
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_92
timestamp 1723858470
transform 1 0 9016 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_110
timestamp 1723858470
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1723858470
transform 1 0 828 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_17
timestamp 1723858470
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_25
timestamp 1723858470
transform 1 0 2852 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_36
timestamp 1723858470
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1723858470
transform 1 0 5152 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 1723858470
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_73
timestamp 1723858470
transform 1 0 7268 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_83
timestamp 1723858470
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_89
timestamp 1723858470
transform 1 0 8740 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_97
timestamp 1723858470
transform 1 0 9476 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1723858470
transform 1 0 10580 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1723858470
transform 1 0 828 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_11
timestamp 1723858470
transform 1 0 1564 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1723858470
transform 1 0 3220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_37
timestamp 1723858470
transform 1 0 3956 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1723858470
transform 1 0 5244 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1723858470
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1723858470
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1723858470
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1723858470
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1723858470
transform 1 0 8372 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_103
timestamp 1723858470
transform 1 0 10028 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_111
timestamp 1723858470
transform 1 0 10764 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1723858470
transform 1 0 828 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1723858470
transform 1 0 1196 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1723858470
transform 1 0 1932 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_42
timestamp 1723858470
transform 1 0 4416 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_52
timestamp 1723858470
transform 1 0 5336 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1723858470
transform 1 0 10580 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1723858470
transform 1 0 828 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 1723858470
transform 1 0 3220 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_39
timestamp 1723858470
transform 1 0 4140 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_43
timestamp 1723858470
transform 1 0 4508 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_55
timestamp 1723858470
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1723858470
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_111
timestamp 1723858470
transform 1 0 10764 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1723858470
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1723858470
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_38
timestamp 1723858470
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1723858470
transform 1 0 4968 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1723858470
transform 1 0 5796 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_69
timestamp 1723858470
transform 1 0 6900 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1723858470
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1723858470
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1723858470
transform 1 0 828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_17
timestamp 1723858470
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_48
timestamp 1723858470
transform 1 0 4968 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_60
timestamp 1723858470
transform 1 0 6072 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_72
timestamp 1723858470
transform 1 0 7176 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_104
timestamp 1723858470
transform 1 0 10120 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1723858470
transform 1 0 828 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp 1723858470
transform 1 0 2300 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1723858470
transform 1 0 5428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_79
timestamp 1723858470
transform 1 0 7820 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_86
timestamp 1723858470
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1723858470
transform 1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1723858470
transform 1 0 828 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1723858470
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_54
timestamp 1723858470
transform 1 0 5520 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_62
timestamp 1723858470
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_81
timestamp 1723858470
transform 1 0 8004 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1723858470
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_94
timestamp 1723858470
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1723858470
transform 1 0 828 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_90
timestamp 1723858470
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_99
timestamp 1723858470
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1723858470
transform 1 0 10120 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1723858470
transform 1 0 828 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1723858470
transform 1 0 2852 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_50
timestamp 1723858470
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1723858470
transform 1 0 7912 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1723858470
transform 1 0 8372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 1723858470
transform 1 0 10396 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_111
timestamp 1723858470
transform 1 0 10764 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_31
timestamp 1723858470
transform 1 0 3404 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1723858470
transform 1 0 5336 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1723858470
transform 1 0 5796 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1723858470
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_74
timestamp 1723858470
transform 1 0 7360 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_78
timestamp 1723858470
transform 1 0 7728 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_86
timestamp 1723858470
transform 1 0 8464 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp 1723858470
transform 1 0 2852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_44
timestamp 1723858470
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_61
timestamp 1723858470
transform 1 0 6164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1723858470
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1723858470
transform 1 0 8372 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_110
timestamp 1723858470
transform 1 0 10672 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1723858470
transform 1 0 828 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_19
timestamp 1723858470
transform 1 0 2300 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1723858470
transform 1 0 5612 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp 1723858470
transform 1 0 5796 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_89
timestamp 1723858470
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_94
timestamp 1723858470
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_98
timestamp 1723858470
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1723858470
transform 1 0 10212 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1723858470
transform 1 0 10764 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1723858470
transform 1 0 828 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_25
timestamp 1723858470
transform 1 0 2852 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_35
timestamp 1723858470
transform 1 0 3772 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_56
timestamp 1723858470
transform 1 0 5704 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1723858470
transform 1 0 8004 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_94
timestamp 1723858470
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_110
timestamp 1723858470
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1723858470
transform 1 0 828 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_7
timestamp 1723858470
transform 1 0 1196 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_80
timestamp 1723858470
transform 1 0 7912 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_88
timestamp 1723858470
transform 1 0 8648 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1723858470
transform 1 0 10304 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1723858470
transform 1 0 828 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_55
timestamp 1723858470
transform 1 0 5612 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_89
timestamp 1723858470
transform 1 0 8740 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_103
timestamp 1723858470
transform 1 0 10028 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_111
timestamp 1723858470
transform 1 0 10764 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1723858470
transform 1 0 828 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_81
timestamp 1723858470
transform 1 0 8004 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1723858470
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_36
timestamp 1723858470
transform 1 0 3864 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_56
timestamp 1723858470
transform 1 0 5704 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1723858470
transform 1 0 8188 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_96
timestamp 1723858470
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_25
timestamp 1723858470
transform 1 0 2852 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1723858470
transform 1 0 5612 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_85
timestamp 1723858470
transform 1 0 8372 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_107
timestamp 1723858470
transform 1 0 10396 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1723858470
transform 1 0 10764 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1723858470
transform 1 0 828 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1723858470
transform 1 0 2852 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_35
timestamp 1723858470
transform 1 0 3772 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_54
timestamp 1723858470
transform 1 0 5520 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1723858470
transform 1 0 8096 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_104
timestamp 1723858470
transform 1 0 10120 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_111
timestamp 1723858470
transform 1 0 10764 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1723858470
transform 1 0 828 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_47
timestamp 1723858470
transform 1 0 4876 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_66
timestamp 1723858470
transform 1 0 6624 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_71
timestamp 1723858470
transform 1 0 7084 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_96
timestamp 1723858470
transform 1 0 9384 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1723858470
transform 1 0 828 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_14
timestamp 1723858470
transform 1 0 1840 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1723858470
transform 1 0 3036 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_41
timestamp 1723858470
transform 1 0 4324 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_56
timestamp 1723858470
transform 1 0 5704 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_95
timestamp 1723858470
transform 1 0 9292 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_25
timestamp 1723858470
transform 1 0 2852 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_32
timestamp 1723858470
transform 1 0 3496 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_63
timestamp 1723858470
transform 1 0 6348 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1723858470
transform 1 0 9660 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_103
timestamp 1723858470
transform 1 0 10028 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_19
timestamp 1723858470
transform 1 0 2300 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1723858470
transform 1 0 3036 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_36
timestamp 1723858470
transform 1 0 3864 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1723858470
transform 1 0 8096 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 1723858470
transform 1 0 8372 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_111
timestamp 1723858470
transform 1 0 10764 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_24
timestamp 1723858470
transform 1 0 2760 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_73
timestamp 1723858470
transform 1 0 7268 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_84
timestamp 1723858470
transform 1 0 8280 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_98
timestamp 1723858470
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1723858470
transform 1 0 10764 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1723858470
transform 1 0 8096 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_27
timestamp 1723858470
transform 1 0 3036 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_60
timestamp 1723858470
transform 1 0 6072 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_79
timestamp 1723858470
transform 1 0 7820 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1723858470
transform 1 0 10672 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_41
timestamp 1723858470
transform 1 0 4324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_78
timestamp 1723858470
transform 1 0 7728 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_101
timestamp 1723858470
transform 1 0 9844 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_110
timestamp 1723858470
transform 1 0 10672 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_57
timestamp 1723858470
transform 1 0 5796 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1723858470
transform 1 0 10764 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_53
timestamp 1723858470
transform 1 0 5428 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_75
timestamp 1723858470
transform 1 0 7452 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_65
timestamp 1723858470
transform 1 0 6532 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_80
timestamp 1723858470
transform 1 0 7912 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1723858470
transform 1 0 828 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_32
timestamp 1723858470
transform 1 0 3496 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_40
timestamp 1723858470
transform 1 0 4232 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_75
timestamp 1723858470
transform 1 0 7452 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_110
timestamp 1723858470
transform 1 0 10672 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1723858470
transform 1 0 828 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_67
timestamp 1723858470
transform 1 0 6716 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_3
timestamp 1723858470
transform 1 0 828 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_78
timestamp 1723858470
transform 1 0 7728 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_111
timestamp 1723858470
transform 1 0 10764 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_3
timestamp 1723858470
transform 1 0 828 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1723858470
transform 1 0 10764 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1723858470
transform 1 0 2944 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_78
timestamp 1723858470
transform 1 0 7728 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_19
timestamp 1723858470
transform 1 0 2300 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_31
timestamp 1723858470
transform 1 0 3404 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_46
timestamp 1723858470
transform 1 0 4784 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1723858470
transform 1 0 5612 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_69
timestamp 1723858470
transform 1 0 6900 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_3
timestamp 1723858470
transform 1 0 828 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_13
timestamp 1723858470
transform 1 0 1748 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_29
timestamp 1723858470
transform 1 0 3220 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_41
timestamp 1723858470
transform 1 0 4324 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp 1723858470
transform 1 0 9108 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_101
timestamp 1723858470
transform 1 0 9844 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_111
timestamp 1723858470
transform 1 0 10764 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1723858470
transform 1 0 828 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_7
timestamp 1723858470
transform 1 0 1196 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_25
timestamp 1723858470
transform 1 0 2852 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_45
timestamp 1723858470
transform 1 0 4692 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_73
timestamp 1723858470
transform 1 0 7268 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_93
timestamp 1723858470
transform 1 0 9108 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1723858470
transform 1 0 10764 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_55
timestamp 1723858470
transform 1 0 5612 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_72
timestamp 1723858470
transform 1 0 7176 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_79
timestamp 1723858470
transform 1 0 7820 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_104
timestamp 1723858470
transform 1 0 10120 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1723858470
transform 1 0 828 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1723858470
transform 1 0 5612 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_57
timestamp 1723858470
transform 1 0 5796 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_65
timestamp 1723858470
transform 1 0 6532 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_93
timestamp 1723858470
transform 1 0 9108 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1723858470
transform 1 0 2944 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_29
timestamp 1723858470
transform 1 0 3220 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1723858470
transform 1 0 8188 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_88
timestamp 1723858470
transform 1 0 8648 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1723858470
transform 1 0 10764 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1723858470
transform 1 0 828 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_31
timestamp 1723858470
transform 1 0 3404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_3
timestamp 1723858470
transform 1 0 828 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp 1723858470
transform 1 0 2944 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_3
timestamp 1723858470
transform 1 0 828 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_76
timestamp 1723858470
transform 1 0 7544 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1723858470
transform 1 0 10672 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_7
timestamp 1723858470
transform 1 0 1196 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_23
timestamp 1723858470
transform 1 0 2668 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_38
timestamp 1723858470
transform 1 0 4048 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_49
timestamp 1723858470
transform 1 0 5060 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_64
timestamp 1723858470
transform 1 0 6440 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_75
timestamp 1723858470
transform 1 0 7452 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_102
timestamp 1723858470
transform 1 0 9936 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_3
timestamp 1723858470
transform 1 0 828 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_30
timestamp 1723858470
transform 1 0 3312 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_54
timestamp 1723858470
transform 1 0 5520 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_66
timestamp 1723858470
transform 1 0 6624 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_100
timestamp 1723858470
transform 1 0 9752 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_34
timestamp 1723858470
transform 1 0 3680 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_51
timestamp 1723858470
transform 1 0 5244 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_66
timestamp 1723858470
transform 1 0 6624 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1723858470
transform 1 0 8188 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_110
timestamp 1723858470
transform 1 0 10672 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1723858470
transform 1 0 828 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_15
timestamp 1723858470
transform 1 0 1932 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_33
timestamp 1723858470
transform 1 0 3588 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_65
timestamp 1723858470
transform 1 0 6532 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1723858470
transform 1 0 828 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1723858470
transform 1 0 3036 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_29
timestamp 1723858470
transform 1 0 3220 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_95
timestamp 1723858470
transform 1 0 9292 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1723858470
transform 1 0 828 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_33
timestamp 1723858470
transform 1 0 3588 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_85
timestamp 1723858470
transform 1 0 8372 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_3
timestamp 1723858470
transform 1 0 828 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_24
timestamp 1723858470
transform 1 0 2760 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_50
timestamp 1723858470
transform 1 0 5152 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_104
timestamp 1723858470
transform 1 0 10120 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1723858470
transform 1 0 10672 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_3
timestamp 1723858470
transform 1 0 828 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_101
timestamp 1723858470
transform 1 0 9844 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_110
timestamp 1723858470
transform 1 0 10672 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1723858470
transform 1 0 828 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_71
timestamp 1723858470
transform 1 0 7084 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_83
timestamp 1723858470
transform 1 0 8188 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_102
timestamp 1723858470
transform 1 0 9936 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 3036 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1723858470
transform -1 0 6440 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1723858470
transform -1 0 5704 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1723858470
transform -1 0 5796 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1723858470
transform -1 0 4784 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1723858470
transform -1 0 4048 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1723858470
transform 1 0 3312 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1723858470
transform -1 0 6624 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1723858470
transform -1 0 7268 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1723858470
transform 1 0 3220 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1723858470
transform -1 0 7912 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1723858470
transform -1 0 6532 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1723858470
transform 1 0 3588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1723858470
transform -1 0 10856 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1723858470
transform 1 0 3128 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1723858470
transform 1 0 3220 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1723858470
transform -1 0 10672 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1723858470
transform 1 0 10120 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5336 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1723858470
transform 1 0 7268 0 -1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1723858470
transform -1 0 6164 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1723858470
transform 1 0 6164 0 -1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1723858470
transform -1 0 10856 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1723858470
transform -1 0 5520 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1723858470
transform -1 0 3128 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1723858470
transform 1 0 3956 0 -1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1723858470
transform -1 0 3128 0 -1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_78
timestamp 1723858470
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1723858470
transform -1 0 11132 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_79
timestamp 1723858470
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1723858470
transform -1 0 11132 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_80
timestamp 1723858470
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1723858470
transform -1 0 11132 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_81
timestamp 1723858470
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1723858470
transform -1 0 11132 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_82
timestamp 1723858470
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1723858470
transform -1 0 11132 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_83
timestamp 1723858470
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1723858470
transform -1 0 11132 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_84
timestamp 1723858470
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1723858470
transform -1 0 11132 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_85
timestamp 1723858470
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1723858470
transform -1 0 11132 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_86
timestamp 1723858470
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1723858470
transform -1 0 11132 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_87
timestamp 1723858470
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1723858470
transform -1 0 11132 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_88
timestamp 1723858470
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1723858470
transform -1 0 11132 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_89
timestamp 1723858470
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1723858470
transform -1 0 11132 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_90
timestamp 1723858470
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1723858470
transform -1 0 11132 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_91
timestamp 1723858470
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1723858470
transform -1 0 11132 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_92
timestamp 1723858470
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1723858470
transform -1 0 11132 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_93
timestamp 1723858470
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1723858470
transform -1 0 11132 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_94
timestamp 1723858470
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1723858470
transform -1 0 11132 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_95
timestamp 1723858470
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1723858470
transform -1 0 11132 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_96
timestamp 1723858470
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1723858470
transform -1 0 11132 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_97
timestamp 1723858470
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1723858470
transform -1 0 11132 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_98
timestamp 1723858470
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1723858470
transform -1 0 11132 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_99
timestamp 1723858470
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1723858470
transform -1 0 11132 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_100
timestamp 1723858470
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1723858470
transform -1 0 11132 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_101
timestamp 1723858470
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1723858470
transform -1 0 11132 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_102
timestamp 1723858470
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1723858470
transform -1 0 11132 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_103
timestamp 1723858470
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1723858470
transform -1 0 11132 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_104
timestamp 1723858470
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1723858470
transform -1 0 11132 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_105
timestamp 1723858470
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1723858470
transform -1 0 11132 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_106
timestamp 1723858470
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1723858470
transform -1 0 11132 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_107
timestamp 1723858470
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1723858470
transform -1 0 11132 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_108
timestamp 1723858470
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1723858470
transform -1 0 11132 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_109
timestamp 1723858470
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1723858470
transform -1 0 11132 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_110
timestamp 1723858470
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1723858470
transform -1 0 11132 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_111
timestamp 1723858470
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1723858470
transform -1 0 11132 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_112
timestamp 1723858470
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1723858470
transform -1 0 11132 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_113
timestamp 1723858470
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1723858470
transform -1 0 11132 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_114
timestamp 1723858470
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1723858470
transform -1 0 11132 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_115
timestamp 1723858470
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1723858470
transform -1 0 11132 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_116
timestamp 1723858470
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1723858470
transform -1 0 11132 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_117
timestamp 1723858470
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1723858470
transform -1 0 11132 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_118
timestamp 1723858470
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1723858470
transform -1 0 11132 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_119
timestamp 1723858470
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1723858470
transform -1 0 11132 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_120
timestamp 1723858470
transform 1 0 552 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1723858470
transform -1 0 11132 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_121
timestamp 1723858470
transform 1 0 552 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1723858470
transform -1 0 11132 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_122
timestamp 1723858470
transform 1 0 552 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1723858470
transform -1 0 11132 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_123
timestamp 1723858470
transform 1 0 552 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1723858470
transform -1 0 11132 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_124
timestamp 1723858470
transform 1 0 552 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1723858470
transform -1 0 11132 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_125
timestamp 1723858470
transform 1 0 552 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1723858470
transform -1 0 11132 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_126
timestamp 1723858470
transform 1 0 552 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1723858470
transform -1 0 11132 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_127
timestamp 1723858470
transform 1 0 552 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1723858470
transform -1 0 11132 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_128
timestamp 1723858470
transform 1 0 552 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1723858470
transform -1 0 11132 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_129
timestamp 1723858470
transform 1 0 552 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1723858470
transform -1 0 11132 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_130
timestamp 1723858470
transform 1 0 552 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1723858470
transform -1 0 11132 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_131
timestamp 1723858470
transform 1 0 552 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1723858470
transform -1 0 11132 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_132
timestamp 1723858470
transform 1 0 552 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1723858470
transform -1 0 11132 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_133
timestamp 1723858470
transform 1 0 552 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1723858470
transform -1 0 11132 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_134
timestamp 1723858470
transform 1 0 552 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1723858470
transform -1 0 11132 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_135
timestamp 1723858470
transform 1 0 552 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1723858470
transform -1 0 11132 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_136
timestamp 1723858470
transform 1 0 552 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1723858470
transform -1 0 11132 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_137
timestamp 1723858470
transform 1 0 552 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1723858470
transform -1 0 11132 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_138
timestamp 1723858470
transform 1 0 552 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1723858470
transform -1 0 11132 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_139
timestamp 1723858470
transform 1 0 552 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1723858470
transform -1 0 11132 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_140
timestamp 1723858470
transform 1 0 552 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1723858470
transform -1 0 11132 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_141
timestamp 1723858470
transform 1 0 552 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1723858470
transform -1 0 11132 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_142
timestamp 1723858470
transform 1 0 552 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1723858470
transform -1 0 11132 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_143
timestamp 1723858470
transform 1 0 552 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1723858470
transform -1 0 11132 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_144
timestamp 1723858470
transform 1 0 552 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1723858470
transform -1 0 11132 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_145
timestamp 1723858470
transform 1 0 552 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1723858470
transform -1 0 11132 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_146
timestamp 1723858470
transform 1 0 552 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1723858470
transform -1 0 11132 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_147
timestamp 1723858470
transform 1 0 552 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 1723858470
transform -1 0 11132 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_148
timestamp 1723858470
transform 1 0 552 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 1723858470
transform -1 0 11132 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_149
timestamp 1723858470
transform 1 0 552 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 1723858470
transform -1 0 11132 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_150
timestamp 1723858470
transform 1 0 552 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 1723858470
transform -1 0 11132 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_151
timestamp 1723858470
transform 1 0 552 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 1723858470
transform -1 0 11132 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_152
timestamp 1723858470
transform 1 0 552 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 1723858470
transform -1 0 11132 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_153
timestamp 1723858470
transform 1 0 552 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 1723858470
transform -1 0 11132 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_154
timestamp 1723858470
transform 1 0 552 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 1723858470
transform -1 0 11132 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_155
timestamp 1723858470
transform 1 0 552 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 1723858470
transform -1 0 11132 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_156 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_157
timestamp 1757695336
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_158
timestamp 1757695336
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_159
timestamp 1757695336
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_160
timestamp 1757695336
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_161
timestamp 1757695336
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_162
timestamp 1757695336
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_163
timestamp 1757695336
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_164
timestamp 1757695336
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_165
timestamp 1757695336
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_166
timestamp 1757695336
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_167
timestamp 1757695336
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_168
timestamp 1757695336
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_169
timestamp 1757695336
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_170
timestamp 1757695336
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_171
timestamp 1757695336
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_172
timestamp 1757695336
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_173
timestamp 1757695336
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_174
timestamp 1757695336
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_175
timestamp 1757695336
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_176
timestamp 1757695336
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_177
timestamp 1757695336
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_178
timestamp 1757695336
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_179
timestamp 1757695336
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_180
timestamp 1757695336
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_181
timestamp 1757695336
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_182
timestamp 1757695336
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_183
timestamp 1757695336
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1757695336
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1757695336
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_186
timestamp 1757695336
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1757695336
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1757695336
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1757695336
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_190
timestamp 1757695336
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_191
timestamp 1757695336
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_192
timestamp 1757695336
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_193
timestamp 1757695336
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_194
timestamp 1757695336
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_195
timestamp 1757695336
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_196
timestamp 1757695336
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_197
timestamp 1757695336
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_198
timestamp 1757695336
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_199
timestamp 1757695336
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_200
timestamp 1757695336
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_201
timestamp 1757695336
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_202
timestamp 1757695336
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_203
timestamp 1757695336
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_204
timestamp 1757695336
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_205
timestamp 1757695336
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_206
timestamp 1757695336
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_207
timestamp 1757695336
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_208
timestamp 1757695336
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_209
timestamp 1757695336
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_210
timestamp 1757695336
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_211
timestamp 1757695336
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_212
timestamp 1757695336
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_213
timestamp 1757695336
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_214
timestamp 1757695336
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_215
timestamp 1757695336
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_216
timestamp 1757695336
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_217
timestamp 1757695336
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_218
timestamp 1757695336
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_219
timestamp 1757695336
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_220
timestamp 1757695336
transform 1 0 3128 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_221
timestamp 1757695336
transform 1 0 8280 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_222
timestamp 1757695336
transform 1 0 5704 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_223
timestamp 1757695336
transform 1 0 3128 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_224
timestamp 1757695336
transform 1 0 8280 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_225
timestamp 1757695336
transform 1 0 5704 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_226
timestamp 1757695336
transform 1 0 3128 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_227
timestamp 1757695336
transform 1 0 8280 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_228
timestamp 1757695336
transform 1 0 5704 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_229
timestamp 1757695336
transform 1 0 3128 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_230
timestamp 1757695336
transform 1 0 8280 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_231
timestamp 1757695336
transform 1 0 5704 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_232
timestamp 1757695336
transform 1 0 3128 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_233
timestamp 1757695336
transform 1 0 8280 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_234
timestamp 1757695336
transform 1 0 5704 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_235
timestamp 1757695336
transform 1 0 3128 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_236
timestamp 1757695336
transform 1 0 8280 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_237
timestamp 1757695336
transform 1 0 5704 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_238
timestamp 1757695336
transform 1 0 3128 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_239
timestamp 1757695336
transform 1 0 8280 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_240
timestamp 1757695336
transform 1 0 5704 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_241
timestamp 1757695336
transform 1 0 3128 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_242
timestamp 1757695336
transform 1 0 8280 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_243
timestamp 1757695336
transform 1 0 5704 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_244
timestamp 1757695336
transform 1 0 3128 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_245
timestamp 1757695336
transform 1 0 8280 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_246
timestamp 1757695336
transform 1 0 5704 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_247
timestamp 1757695336
transform 1 0 3128 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_248
timestamp 1757695336
transform 1 0 8280 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_249
timestamp 1757695336
transform 1 0 5704 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_250
timestamp 1757695336
transform 1 0 3128 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_251
timestamp 1757695336
transform 1 0 8280 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_252
timestamp 1757695336
transform 1 0 5704 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_253
timestamp 1757695336
transform 1 0 3128 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_254
timestamp 1757695336
transform 1 0 8280 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_255
timestamp 1757695336
transform 1 0 5704 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_256
timestamp 1757695336
transform 1 0 3128 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_257
timestamp 1757695336
transform 1 0 8280 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_258
timestamp 1757695336
transform 1 0 5704 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_259
timestamp 1757695336
transform 1 0 3128 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_260
timestamp 1757695336
transform 1 0 8280 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_261
timestamp 1757695336
transform 1 0 5704 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_262
timestamp 1757695336
transform 1 0 3128 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_263
timestamp 1757695336
transform 1 0 8280 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_264
timestamp 1757695336
transform 1 0 5704 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_265
timestamp 1757695336
transform 1 0 3128 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_266
timestamp 1757695336
transform 1 0 8280 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_267
timestamp 1757695336
transform 1 0 5704 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_268
timestamp 1757695336
transform 1 0 3128 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_269
timestamp 1757695336
transform 1 0 8280 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_270
timestamp 1757695336
transform 1 0 5704 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_271
timestamp 1757695336
transform 1 0 3128 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_272
timestamp 1757695336
transform 1 0 8280 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_273
timestamp 1757695336
transform 1 0 3128 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_274
timestamp 1757695336
transform 1 0 5704 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_275
timestamp 1757695336
transform 1 0 8280 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire12
timestamp 1723858470
transform 1 0 6072 0 1 28832
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 11704 400 11824 0 FreeSans 600 0 0 0 B[0]
port 1 nsew
flabel metal3 s 0 11976 400 12096 0 FreeSans 600 0 0 0 B[1]
port 2 nsew
flabel metal3 s 0 12248 400 12368 0 FreeSans 600 0 0 0 B[2]
port 3 nsew
flabel metal3 s 0 12520 400 12640 0 FreeSans 600 0 0 0 B[3]
port 4 nsew
flabel metal3 s 0 5448 400 5568 0 FreeSans 600 0 0 0 B[4]
port 5 nsew
flabel metal3 s 0 5176 400 5296 0 FreeSans 600 0 0 0 B[5]
port 6 nsew
flabel metal3 s 0 4904 400 5024 0 FreeSans 600 0 0 0 B[6]
port 7 nsew
flabel metal3 s 0 4632 400 4752 0 FreeSans 600 0 0 0 B[7]
port 8 nsew
flabel metal3 s 0 11432 400 11552 0 FreeSans 600 0 0 0 Bbias[0]
port 9 nsew
flabel metal3 s 0 11160 400 11280 0 FreeSans 600 0 0 0 Bbias[1]
port 10 nsew
flabel metal3 s 0 10888 400 11008 0 FreeSans 600 0 0 0 Bbias[2]
port 11 nsew
flabel metal3 s 0 23400 400 23520 0 FreeSans 600 0 0 0 G[0]
port 12 nsew
flabel metal3 s 0 23672 400 23792 0 FreeSans 600 0 0 0 G[1]
port 13 nsew
flabel metal3 s 0 23944 400 24064 0 FreeSans 600 0 0 0 G[2]
port 14 nsew
flabel metal3 s 0 24216 400 24336 0 FreeSans 600 0 0 0 G[3]
port 15 nsew
flabel metal3 s 0 17144 400 17264 0 FreeSans 600 0 0 0 G[4]
port 16 nsew
flabel metal3 s 0 16872 400 16992 0 FreeSans 600 0 0 0 G[5]
port 17 nsew
flabel metal3 s 0 16600 400 16720 0 FreeSans 600 0 0 0 G[6]
port 18 nsew
flabel metal3 s 0 16328 400 16448 0 FreeSans 600 0 0 0 G[7]
port 19 nsew
flabel metal3 s 0 23128 400 23248 0 FreeSans 600 0 0 0 Gbias[0]
port 20 nsew
flabel metal3 s 0 22856 400 22976 0 FreeSans 600 0 0 0 Gbias[1]
port 21 nsew
flabel metal3 s 0 22584 400 22704 0 FreeSans 600 0 0 0 Gbias[2]
port 22 nsew
flabel metal3 s 0 36184 400 36304 0 FreeSans 600 0 0 0 R[0]
port 23 nsew
flabel metal3 s 0 36456 400 36576 0 FreeSans 600 0 0 0 R[1]
port 24 nsew
flabel metal3 s 0 36728 400 36848 0 FreeSans 600 0 0 0 R[2]
port 25 nsew
flabel metal3 s 0 37000 400 37120 0 FreeSans 600 0 0 0 R[3]
port 26 nsew
flabel metal3 s 0 28840 400 28960 0 FreeSans 600 0 0 0 R[4]
port 27 nsew
flabel metal3 s 0 28568 400 28688 0 FreeSans 600 0 0 0 R[5]
port 28 nsew
flabel metal3 s 0 28296 400 28416 0 FreeSans 600 0 0 0 R[6]
port 29 nsew
flabel metal3 s 0 28024 400 28144 0 FreeSans 600 0 0 0 R[7]
port 30 nsew
flabel metal3 s 0 34824 400 34944 0 FreeSans 600 0 0 0 Rbias[0]
port 31 nsew
flabel metal3 s 0 34552 400 34672 0 FreeSans 600 0 0 0 Rbias[1]
port 32 nsew
flabel metal3 s 0 34280 400 34400 0 FreeSans 600 0 0 0 Rbias[2]
port 33 nsew
flabel metal4 s 10716 496 11036 43024 0 FreeSans 2400 90 0 0 VGND
port 34 nsew
flabel metal4 s 4316 496 4636 43024 0 FreeSans 2400 90 0 0 VGND
port 34 nsew
flabel metal4 s 10056 496 10376 43024 0 FreeSans 2400 90 0 0 VPWR
port 35 nsew
flabel metal4 s 3656 496 3976 43024 0 FreeSans 2400 90 0 0 VPWR
port 35 nsew
flabel metal2 s 8298 43500 8354 43900 0 FreeSans 280 90 0 0 clk
port 36 nsew
flabel metal2 s 8850 43500 8906 43900 0 FreeSans 280 90 0 0 ena
port 37 nsew
flabel metal2 s 7746 43500 7802 43900 0 FreeSans 280 90 0 0 rst_n
port 38 nsew
flabel metal2 s 7194 43500 7250 43900 0 FreeSans 280 90 0 0 ui_in[0]
port 39 nsew
flabel metal2 s 6642 43500 6698 43900 0 FreeSans 280 90 0 0 ui_in[1]
port 40 nsew
flabel metal2 s 6090 43500 6146 43900 0 FreeSans 280 90 0 0 ui_in[2]
port 41 nsew
flabel metal2 s 5538 43500 5594 43900 0 FreeSans 280 90 0 0 ui_in[3]
port 42 nsew
flabel metal2 s 4986 43500 5042 43900 0 FreeSans 280 90 0 0 ui_in[4]
port 43 nsew
flabel metal2 s 4434 43500 4490 43900 0 FreeSans 280 90 0 0 ui_in[5]
port 44 nsew
flabel metal2 s 3882 43500 3938 43900 0 FreeSans 280 90 0 0 ui_in[6]
port 45 nsew
flabel metal2 s 3330 43500 3386 43900 0 FreeSans 280 90 0 0 ui_in[7]
port 46 nsew
flabel metal2 s 1674 43500 1730 43900 0 FreeSans 280 90 0 0 uio_in2
port 47 nsew
flabel metal2 s 1122 43500 1178 43900 0 FreeSans 280 90 0 0 uio_in3
port 48 nsew
flabel metal2 s 570 43500 626 43900 0 FreeSans 280 90 0 0 uio_in4
port 49 nsew
flabel metal3 s 0 39448 400 39568 0 FreeSans 600 0 0 0 uio_out[0]
port 50 nsew
flabel metal3 s 0 39176 400 39296 0 FreeSans 600 0 0 0 uio_out[1]
port 51 nsew
flabel metal3 s 0 41624 400 41744 0 FreeSans 600 0 0 0 uo_out[0]
port 52 nsew
flabel metal3 s 0 41352 400 41472 0 FreeSans 600 0 0 0 uo_out[1]
port 53 nsew
flabel metal3 s 0 41080 400 41200 0 FreeSans 600 0 0 0 uo_out[2]
port 54 nsew
flabel metal3 s 0 40808 400 40928 0 FreeSans 600 0 0 0 uo_out[3]
port 55 nsew
flabel metal3 s 0 40536 400 40656 0 FreeSans 600 0 0 0 uo_out[4]
port 56 nsew
flabel metal3 s 0 40264 400 40384 0 FreeSans 600 0 0 0 uo_out[5]
port 57 nsew
flabel metal3 s 0 39992 400 40112 0 FreeSans 600 0 0 0 uo_out[6]
port 58 nsew
flabel metal3 s 0 39720 400 39840 0 FreeSans 600 0 0 0 uo_out[7]
port 59 nsew
<< properties >>
string FIXED_BBOX 0 0 11400 43900
string GDS_END 3477402
string GDS_FILE ../gds/controller_wrapper.gds
string GDS_START 582034
<< end >>
