magic
tech sky130A
timestamp 1762784779
<< metal1 >>
rect 450 220 468 232
rect 843 220 861 232
rect 1236 220 1254 232
rect 1629 220 1647 232
rect 2022 220 2040 232
rect 2415 220 2433 232
rect 2808 220 2826 232
rect 3201 220 3219 232
rect 3594 220 3612 232
rect 3987 220 4005 232
rect 4380 220 4398 232
rect 4773 220 4791 232
rect 5166 220 5184 232
rect 5559 220 5577 232
rect 5952 220 5970 232
<< metal2 >>
rect -28 188 407 202
rect -28 -44 407 -30
<< metal3 >>
rect 0 213 30 243
rect 173 213 217 243
rect 726 213 756 243
<< metal4 >>
rect 6640 7 6681 48
use icellwrap  XIC[0]
timestamp 1762784779
transform 1 0 393 0 1 0
box 0 -55 393 243
use icellwrap  XIC[1]
timestamp 1762784779
transform 1 0 786 0 1 0
box 0 -55 393 243
use icellwrap  XIC[2]
timestamp 1762784779
transform 1 0 1179 0 1 0
box 0 -55 393 243
use icellwrap  XIC[3]
timestamp 1762784779
transform 1 0 1572 0 1 0
box 0 -55 393 243
use icellwrap  XIC[4]
timestamp 1762784779
transform 1 0 1965 0 1 0
box 0 -55 393 243
use icellwrap  XIC[5]
timestamp 1762784779
transform 1 0 2358 0 1 0
box 0 -55 393 243
use icellwrap  XIC[6]
timestamp 1762784779
transform 1 0 2751 0 1 0
box 0 -55 393 243
use icellwrap  XIC[7]
timestamp 1762784779
transform 1 0 3144 0 1 0
box 0 -55 393 243
use icellwrap  XIC[8]
timestamp 1762784779
transform 1 0 3537 0 1 0
box 0 -55 393 243
use icellwrap  XIC[9]
timestamp 1762784779
transform 1 0 3930 0 1 0
box 0 -55 393 243
use icellwrap  XIC[10]
timestamp 1762784779
transform 1 0 4323 0 1 0
box 0 -55 393 243
use icellwrap  XIC[11]
timestamp 1762784779
transform 1 0 4716 0 1 0
box 0 -55 393 243
use icellwrap  XIC[12]
timestamp 1762784779
transform 1 0 5109 0 1 0
box 0 -55 393 243
use icellwrap  XIC[13]
timestamp 1762784779
transform 1 0 5502 0 1 0
box 0 -55 393 243
use icellwrap  XIC[14]
timestamp 1762784779
transform 1 0 5895 0 1 0
box 0 -55 393 243
use icellwrapfinal  XIC_15
timestamp 1762784779
transform 1 0 6288 0 1 0
box 0 -47 393 243
use icellwrapdummy  XIC_dummy_left
timestamp 1762784779
transform 1 0 0 0 1 0
box 0 -4 393 243
use icellwrapdummy  XIC_dummy_right
timestamp 1762784779
transform 1 0 6681 0 1 0
box 0 -4 393 243
<< labels >>
flabel metal2 -28 188 -14 202 0 FreeSans 40 0 0 0 Rn
port 0 nsew
flabel metal2 -28 -44 -14 -30 0 FreeSans 40 0 0 0 Sn
port 1 nsew
flabel metal3 0 220 30 232 0 FreeSans 48 0 0 0 VPWR
port 2 nsew
flabel metal3 173 220 217 232 0 FreeSans 48 0 0 0 VGND
port 3 nsew
flabel metal4 6640 7 6681 48 0 FreeSans 48 0 0 0 Iout
port 4 nsew
flabel metal3 726 220 756 232 0 FreeSans 48 0 0 0 Vbias
port 5 nsew
flabel metal1 450 220 468 232 0 FreeSans 40 0 0 0 Cn[0]
port 6 nsew
flabel metal1 843 220 861 232 0 FreeSans 40 0 0 0 Cn[1]
port 7 nsew
flabel metal1 1236 220 1254 232 0 FreeSans 40 0 0 0 Cn[2]
port 8 nsew
flabel metal1 1629 220 1647 232 0 FreeSans 40 0 0 0 Cn[3]
port 9 nsew
flabel metal1 2022 220 2040 232 0 FreeSans 40 0 0 0 Cn[4]
port 10 nsew
flabel metal1 2415 220 2433 232 0 FreeSans 40 0 0 0 Cn[5]
port 11 nsew
flabel metal1 2808 220 2826 232 0 FreeSans 40 0 0 0 Cn[6]
port 12 nsew
flabel metal1 3201 220 3219 232 0 FreeSans 40 0 0 0 Cn[7]
port 13 nsew
flabel metal1 3594 220 3612 232 0 FreeSans 40 0 0 0 Cn[8]
port 14 nsew
flabel metal1 3987 220 4005 232 0 FreeSans 40 0 0 0 Cn[9]
port 15 nsew
flabel metal1 4380 220 4398 232 0 FreeSans 40 0 0 0 Cn[10]
port 17 nsew
flabel metal1 4773 220 4791 232 0 FreeSans 40 0 0 0 Cn[11]
port 18 nsew
flabel metal1 5166 220 5184 232 0 FreeSans 40 0 0 0 Cn[12]
port 19 nsew
flabel metal1 5559 220 5577 232 0 FreeSans 40 0 0 0 Cn[13]
port 20 nsew
flabel metal1 5952 220 5970 232 0 FreeSans 40 0 0 0 Cn[14]
port 21 nsew
<< properties >>
string FIXED_BBOX 0 0 7074 232
<< end >>
